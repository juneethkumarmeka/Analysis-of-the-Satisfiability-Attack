module basic_1500_15000_2000_3_levels_5xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10004,N_10006,N_10007,N_10008,N_10009,N_10010,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10029,N_10030,N_10031,N_10032,N_10035,N_10037,N_10038,N_10040,N_10042,N_10043,N_10044,N_10045,N_10047,N_10048,N_10049,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10072,N_10073,N_10074,N_10076,N_10077,N_10078,N_10079,N_10080,N_10082,N_10083,N_10084,N_10085,N_10086,N_10088,N_10089,N_10090,N_10092,N_10093,N_10094,N_10095,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10126,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10164,N_10165,N_10168,N_10169,N_10170,N_10171,N_10173,N_10174,N_10175,N_10176,N_10177,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10194,N_10195,N_10196,N_10197,N_10199,N_10200,N_10201,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10228,N_10229,N_10230,N_10232,N_10233,N_10235,N_10236,N_10237,N_10238,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10280,N_10281,N_10283,N_10284,N_10285,N_10286,N_10287,N_10289,N_10290,N_10291,N_10294,N_10295,N_10296,N_10297,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10331,N_10332,N_10334,N_10337,N_10339,N_10340,N_10342,N_10343,N_10345,N_10346,N_10348,N_10349,N_10350,N_10352,N_10354,N_10355,N_10357,N_10358,N_10359,N_10360,N_10362,N_10363,N_10364,N_10365,N_10366,N_10368,N_10369,N_10370,N_10371,N_10373,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10393,N_10395,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10404,N_10405,N_10406,N_10407,N_10408,N_10410,N_10411,N_10412,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10422,N_10423,N_10424,N_10425,N_10427,N_10428,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10450,N_10452,N_10453,N_10455,N_10456,N_10457,N_10459,N_10461,N_10462,N_10464,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10496,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10523,N_10525,N_10526,N_10528,N_10531,N_10533,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10551,N_10552,N_10553,N_10554,N_10555,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10566,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10577,N_10579,N_10580,N_10581,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10609,N_10610,N_10612,N_10613,N_10615,N_10616,N_10617,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10629,N_10630,N_10631,N_10632,N_10633,N_10635,N_10636,N_10637,N_10640,N_10642,N_10643,N_10644,N_10645,N_10647,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10657,N_10658,N_10659,N_10660,N_10661,N_10663,N_10664,N_10667,N_10668,N_10669,N_10671,N_10672,N_10673,N_10675,N_10676,N_10677,N_10678,N_10679,N_10681,N_10682,N_10683,N_10684,N_10686,N_10688,N_10689,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10715,N_10716,N_10717,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10727,N_10728,N_10732,N_10733,N_10735,N_10737,N_10738,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10763,N_10764,N_10766,N_10767,N_10768,N_10769,N_10771,N_10772,N_10773,N_10774,N_10775,N_10779,N_10780,N_10782,N_10783,N_10784,N_10786,N_10787,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10819,N_10821,N_10822,N_10823,N_10824,N_10825,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10839,N_10840,N_10841,N_10842,N_10844,N_10845,N_10846,N_10847,N_10848,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10859,N_10860,N_10861,N_10862,N_10863,N_10865,N_10866,N_10867,N_10868,N_10870,N_10871,N_10872,N_10873,N_10875,N_10878,N_10879,N_10880,N_10883,N_10884,N_10885,N_10887,N_10888,N_10889,N_10890,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10901,N_10902,N_10903,N_10905,N_10906,N_10907,N_10908,N_10910,N_10911,N_10912,N_10913,N_10914,N_10917,N_10919,N_10920,N_10921,N_10922,N_10924,N_10925,N_10926,N_10928,N_10931,N_10933,N_10934,N_10935,N_10936,N_10937,N_10940,N_10941,N_10942,N_10943,N_10944,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10964,N_10965,N_10966,N_10967,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11003,N_11004,N_11006,N_11008,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11018,N_11019,N_11020,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11031,N_11032,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11056,N_11058,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11074,N_11075,N_11076,N_11077,N_11078,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11087,N_11091,N_11092,N_11093,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11108,N_11109,N_11110,N_11111,N_11112,N_11114,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11125,N_11126,N_11128,N_11129,N_11130,N_11132,N_11133,N_11136,N_11138,N_11139,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11157,N_11158,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11173,N_11174,N_11175,N_11178,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11247,N_11248,N_11252,N_11253,N_11254,N_11256,N_11258,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11273,N_11274,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11296,N_11297,N_11298,N_11300,N_11301,N_11302,N_11303,N_11306,N_11307,N_11308,N_11309,N_11310,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11331,N_11332,N_11333,N_11334,N_11335,N_11337,N_11338,N_11339,N_11341,N_11343,N_11344,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11370,N_11371,N_11373,N_11374,N_11375,N_11376,N_11377,N_11379,N_11382,N_11383,N_11384,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11405,N_11408,N_11409,N_11412,N_11413,N_11414,N_11415,N_11416,N_11418,N_11419,N_11420,N_11421,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11434,N_11435,N_11437,N_11438,N_11441,N_11442,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11463,N_11465,N_11468,N_11469,N_11470,N_11471,N_11473,N_11474,N_11476,N_11477,N_11478,N_11479,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11490,N_11492,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11512,N_11513,N_11514,N_11515,N_11516,N_11518,N_11520,N_11522,N_11523,N_11525,N_11526,N_11527,N_11528,N_11530,N_11531,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11560,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11575,N_11576,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11593,N_11594,N_11595,N_11596,N_11597,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11608,N_11609,N_11610,N_11611,N_11613,N_11614,N_11615,N_11618,N_11619,N_11620,N_11622,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11631,N_11632,N_11633,N_11635,N_11636,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11648,N_11649,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11686,N_11687,N_11688,N_11690,N_11691,N_11693,N_11694,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11753,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11765,N_11766,N_11767,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11809,N_11810,N_11811,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11828,N_11830,N_11831,N_11832,N_11835,N_11837,N_11838,N_11839,N_11840,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11861,N_11862,N_11864,N_11865,N_11866,N_11867,N_11868,N_11871,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11880,N_11881,N_11882,N_11884,N_11886,N_11887,N_11888,N_11891,N_11892,N_11894,N_11896,N_11897,N_11898,N_11899,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11910,N_11912,N_11913,N_11914,N_11915,N_11916,N_11918,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11932,N_11933,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11987,N_11988,N_11989,N_11991,N_11992,N_11994,N_11995,N_11996,N_11997,N_12000,N_12001,N_12002,N_12003,N_12005,N_12006,N_12007,N_12008,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12022,N_12024,N_12025,N_12026,N_12027,N_12030,N_12031,N_12033,N_12034,N_12035,N_12037,N_12038,N_12039,N_12040,N_12043,N_12044,N_12045,N_12046,N_12047,N_12049,N_12050,N_12051,N_12053,N_12054,N_12055,N_12056,N_12057,N_12059,N_12060,N_12061,N_12062,N_12063,N_12065,N_12066,N_12067,N_12068,N_12070,N_12071,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12084,N_12086,N_12087,N_12088,N_12089,N_12091,N_12092,N_12094,N_12095,N_12096,N_12102,N_12103,N_12104,N_12105,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12123,N_12124,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12154,N_12156,N_12158,N_12159,N_12160,N_12161,N_12162,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12185,N_12186,N_12187,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12202,N_12204,N_12205,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12217,N_12218,N_12219,N_12221,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12236,N_12237,N_12240,N_12241,N_12242,N_12243,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12257,N_12258,N_12259,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12289,N_12290,N_12291,N_12293,N_12294,N_12295,N_12297,N_12298,N_12299,N_12300,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12309,N_12310,N_12311,N_12312,N_12313,N_12315,N_12317,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12372,N_12373,N_12375,N_12376,N_12377,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12398,N_12399,N_12400,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12411,N_12413,N_12414,N_12415,N_12417,N_12418,N_12419,N_12422,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12433,N_12436,N_12437,N_12440,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12459,N_12460,N_12461,N_12462,N_12463,N_12465,N_12466,N_12467,N_12469,N_12470,N_12472,N_12474,N_12475,N_12476,N_12477,N_12478,N_12481,N_12482,N_12483,N_12485,N_12486,N_12488,N_12489,N_12491,N_12493,N_12494,N_12495,N_12497,N_12498,N_12500,N_12501,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12515,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12538,N_12540,N_12542,N_12543,N_12544,N_12546,N_12547,N_12548,N_12551,N_12552,N_12554,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12564,N_12565,N_12566,N_12567,N_12568,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12580,N_12581,N_12582,N_12583,N_12585,N_12586,N_12587,N_12590,N_12591,N_12592,N_12594,N_12595,N_12596,N_12598,N_12599,N_12601,N_12602,N_12604,N_12606,N_12609,N_12610,N_12611,N_12613,N_12614,N_12615,N_12617,N_12618,N_12619,N_12620,N_12622,N_12623,N_12624,N_12625,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12635,N_12636,N_12638,N_12639,N_12640,N_12641,N_12643,N_12644,N_12645,N_12646,N_12647,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12677,N_12678,N_12680,N_12681,N_12682,N_12683,N_12685,N_12687,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12699,N_12700,N_12701,N_12702,N_12704,N_12705,N_12706,N_12707,N_12708,N_12710,N_12711,N_12712,N_12714,N_12715,N_12716,N_12718,N_12720,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12732,N_12733,N_12734,N_12735,N_12737,N_12738,N_12739,N_12741,N_12742,N_12743,N_12744,N_12746,N_12747,N_12748,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12764,N_12767,N_12768,N_12770,N_12771,N_12772,N_12773,N_12774,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12802,N_12803,N_12807,N_12808,N_12809,N_12811,N_12812,N_12814,N_12815,N_12816,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12828,N_12829,N_12831,N_12832,N_12833,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12844,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12857,N_12858,N_12860,N_12861,N_12862,N_12863,N_12867,N_12869,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12881,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12912,N_12913,N_12915,N_12917,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12926,N_12928,N_12929,N_12930,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12950,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12987,N_12988,N_12989,N_12990,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13006,N_13007,N_13008,N_13009,N_13010,N_13012,N_13014,N_13016,N_13018,N_13019,N_13020,N_13021,N_13023,N_13024,N_13025,N_13026,N_13028,N_13029,N_13031,N_13033,N_13034,N_13035,N_13036,N_13038,N_13039,N_13040,N_13041,N_13042,N_13044,N_13046,N_13049,N_13051,N_13053,N_13055,N_13056,N_13057,N_13059,N_13061,N_13062,N_13063,N_13064,N_13065,N_13067,N_13069,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13088,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13104,N_13105,N_13106,N_13107,N_13108,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13119,N_13120,N_13121,N_13122,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13131,N_13132,N_13133,N_13135,N_13137,N_13138,N_13139,N_13141,N_13142,N_13143,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13154,N_13155,N_13156,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13166,N_13168,N_13169,N_13170,N_13171,N_13173,N_13174,N_13175,N_13176,N_13177,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13186,N_13187,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13201,N_13203,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13220,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13232,N_13233,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13269,N_13270,N_13271,N_13272,N_13273,N_13275,N_13276,N_13278,N_13279,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13289,N_13290,N_13291,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13308,N_13310,N_13311,N_13312,N_13313,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13324,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13341,N_13342,N_13344,N_13345,N_13346,N_13348,N_13349,N_13351,N_13352,N_13353,N_13354,N_13355,N_13357,N_13358,N_13359,N_13361,N_13362,N_13364,N_13365,N_13366,N_13368,N_13369,N_13370,N_13373,N_13374,N_13377,N_13379,N_13380,N_13381,N_13383,N_13384,N_13385,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13410,N_13411,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13452,N_13453,N_13454,N_13455,N_13457,N_13458,N_13459,N_13461,N_13462,N_13463,N_13464,N_13465,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13489,N_13490,N_13492,N_13495,N_13496,N_13497,N_13498,N_13503,N_13504,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13514,N_13515,N_13517,N_13518,N_13519,N_13520,N_13521,N_13523,N_13524,N_13527,N_13528,N_13529,N_13531,N_13532,N_13533,N_13535,N_13536,N_13537,N_13538,N_13540,N_13542,N_13543,N_13544,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13559,N_13560,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13583,N_13584,N_13585,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13608,N_13609,N_13610,N_13611,N_13612,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13657,N_13659,N_13660,N_13662,N_13663,N_13665,N_13667,N_13668,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13685,N_13686,N_13687,N_13688,N_13689,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13705,N_13706,N_13707,N_13708,N_13709,N_13711,N_13712,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13728,N_13729,N_13730,N_13731,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13740,N_13741,N_13742,N_13743,N_13745,N_13746,N_13748,N_13749,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13759,N_13760,N_13761,N_13762,N_13764,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13781,N_13782,N_13785,N_13787,N_13789,N_13791,N_13792,N_13793,N_13794,N_13797,N_13799,N_13800,N_13801,N_13805,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13817,N_13818,N_13819,N_13821,N_13822,N_13823,N_13824,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13835,N_13837,N_13838,N_13839,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13853,N_13855,N_13856,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13877,N_13878,N_13879,N_13880,N_13881,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13894,N_13895,N_13896,N_13898,N_13900,N_13901,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13937,N_13938,N_13939,N_13941,N_13942,N_13945,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13956,N_13957,N_13958,N_13959,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13993,N_13995,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14032,N_14033,N_14035,N_14037,N_14038,N_14039,N_14041,N_14042,N_14043,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14055,N_14059,N_14060,N_14062,N_14068,N_14070,N_14071,N_14072,N_14073,N_14074,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14093,N_14095,N_14096,N_14098,N_14099,N_14100,N_14101,N_14102,N_14104,N_14105,N_14106,N_14107,N_14108,N_14110,N_14111,N_14114,N_14115,N_14116,N_14117,N_14119,N_14121,N_14123,N_14125,N_14126,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14143,N_14144,N_14145,N_14146,N_14148,N_14150,N_14151,N_14153,N_14155,N_14157,N_14158,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14170,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14180,N_14181,N_14183,N_14184,N_14185,N_14186,N_14188,N_14189,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14199,N_14200,N_14201,N_14202,N_14203,N_14205,N_14207,N_14208,N_14209,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14228,N_14230,N_14231,N_14232,N_14233,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14243,N_14245,N_14246,N_14247,N_14248,N_14250,N_14251,N_14252,N_14253,N_14254,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14279,N_14280,N_14283,N_14284,N_14285,N_14286,N_14287,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14303,N_14305,N_14307,N_14308,N_14309,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14350,N_14351,N_14352,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14363,N_14364,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14381,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14398,N_14400,N_14402,N_14403,N_14404,N_14405,N_14406,N_14408,N_14409,N_14410,N_14411,N_14412,N_14415,N_14416,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14427,N_14428,N_14431,N_14432,N_14433,N_14434,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14446,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14464,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14478,N_14479,N_14480,N_14481,N_14482,N_14484,N_14485,N_14486,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14541,N_14542,N_14543,N_14544,N_14546,N_14547,N_14549,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14562,N_14564,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14586,N_14587,N_14588,N_14590,N_14591,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14605,N_14606,N_14607,N_14608,N_14609,N_14611,N_14613,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14623,N_14624,N_14625,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14637,N_14638,N_14640,N_14642,N_14643,N_14644,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14662,N_14663,N_14666,N_14667,N_14669,N_14670,N_14671,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14687,N_14688,N_14690,N_14691,N_14692,N_14693,N_14694,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14713,N_14714,N_14717,N_14718,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14737,N_14739,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14749,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14762,N_14763,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14846,N_14847,N_14848,N_14851,N_14852,N_14853,N_14854,N_14855,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14868,N_14869,N_14871,N_14872,N_14873,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14901,N_14903,N_14905,N_14906,N_14907,N_14909,N_14910,N_14911,N_14912,N_14914,N_14915,N_14916,N_14918,N_14919,N_14926,N_14927,N_14928,N_14929,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14940,N_14941,N_14944,N_14945,N_14946,N_14948,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14966,N_14967,N_14968,N_14970,N_14971,N_14972,N_14975,N_14976,N_14977,N_14978,N_14979,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14990,N_14991,N_14992,N_14994,N_14995,N_14996,N_14997,N_14998;
and U0 (N_0,In_513,In_374);
or U1 (N_1,In_1085,In_1090);
xnor U2 (N_2,In_427,In_1118);
or U3 (N_3,In_70,In_1391);
nor U4 (N_4,In_307,In_1218);
and U5 (N_5,In_1277,In_821);
and U6 (N_6,In_1246,In_633);
nor U7 (N_7,In_900,In_1358);
or U8 (N_8,In_792,In_1234);
or U9 (N_9,In_1484,In_781);
nand U10 (N_10,In_772,In_1288);
and U11 (N_11,In_1333,In_7);
and U12 (N_12,In_66,In_688);
nor U13 (N_13,In_118,In_1212);
nand U14 (N_14,In_1461,In_619);
and U15 (N_15,In_1350,In_1481);
or U16 (N_16,In_62,In_135);
or U17 (N_17,In_730,In_644);
or U18 (N_18,In_1167,In_1449);
and U19 (N_19,In_973,In_13);
nor U20 (N_20,In_1458,In_1279);
xor U21 (N_21,In_388,In_317);
nor U22 (N_22,In_1198,In_966);
nand U23 (N_23,In_1448,In_731);
and U24 (N_24,In_941,In_691);
nand U25 (N_25,In_915,In_261);
nor U26 (N_26,In_764,In_113);
xor U27 (N_27,In_1187,In_657);
nand U28 (N_28,In_313,In_970);
or U29 (N_29,In_27,In_1154);
or U30 (N_30,In_642,In_1462);
or U31 (N_31,In_373,In_123);
and U32 (N_32,In_447,In_446);
and U33 (N_33,In_1248,In_82);
and U34 (N_34,In_1250,In_942);
or U35 (N_35,In_304,In_1438);
or U36 (N_36,In_521,In_311);
and U37 (N_37,In_1347,In_293);
or U38 (N_38,In_1425,In_822);
or U39 (N_39,In_160,In_1128);
or U40 (N_40,In_334,In_574);
nand U41 (N_41,In_473,In_628);
nor U42 (N_42,In_766,In_178);
nand U43 (N_43,In_981,In_605);
and U44 (N_44,In_59,In_616);
or U45 (N_45,In_734,In_341);
nand U46 (N_46,In_924,In_486);
nand U47 (N_47,In_880,In_1326);
and U48 (N_48,In_958,In_1026);
nor U49 (N_49,In_319,In_149);
or U50 (N_50,In_1343,In_1173);
or U51 (N_51,In_1002,In_523);
and U52 (N_52,In_1321,In_272);
or U53 (N_53,In_1238,In_623);
xor U54 (N_54,In_357,In_1328);
and U55 (N_55,In_434,In_1144);
and U56 (N_56,In_1372,In_286);
nand U57 (N_57,In_1088,In_409);
xor U58 (N_58,In_443,In_945);
nor U59 (N_59,In_692,In_569);
or U60 (N_60,In_1202,In_1394);
and U61 (N_61,In_283,In_469);
or U62 (N_62,In_856,In_454);
or U63 (N_63,In_218,In_253);
nor U64 (N_64,In_77,In_423);
and U65 (N_65,In_1311,In_663);
and U66 (N_66,In_1264,In_1183);
nor U67 (N_67,In_700,In_445);
nor U68 (N_68,In_535,In_1254);
or U69 (N_69,In_216,In_618);
or U70 (N_70,In_868,In_639);
nor U71 (N_71,In_690,In_796);
and U72 (N_72,In_338,In_1188);
xor U73 (N_73,In_277,In_548);
or U74 (N_74,In_359,In_1072);
nand U75 (N_75,In_193,In_1431);
nor U76 (N_76,In_479,In_685);
xor U77 (N_77,In_1101,In_879);
xor U78 (N_78,In_170,In_546);
nand U79 (N_79,In_115,In_1359);
nand U80 (N_80,In_94,In_1171);
or U81 (N_81,In_957,In_570);
or U82 (N_82,In_380,In_3);
nand U83 (N_83,In_827,In_793);
nand U84 (N_84,In_1256,In_1435);
or U85 (N_85,In_527,In_1368);
or U86 (N_86,In_1061,In_1217);
or U87 (N_87,In_763,In_1447);
and U88 (N_88,In_816,In_207);
nand U89 (N_89,In_624,In_251);
or U90 (N_90,In_383,In_1012);
nor U91 (N_91,In_1080,In_750);
or U92 (N_92,In_844,In_1339);
or U93 (N_93,In_1293,In_1180);
nor U94 (N_94,In_516,In_534);
nor U95 (N_95,In_1089,In_976);
nand U96 (N_96,In_202,In_774);
and U97 (N_97,In_353,In_1204);
nor U98 (N_98,In_839,In_835);
or U99 (N_99,In_408,In_531);
and U100 (N_100,In_1142,In_1139);
and U101 (N_101,In_1262,In_820);
and U102 (N_102,In_1352,In_591);
xor U103 (N_103,In_626,In_1330);
or U104 (N_104,In_354,In_122);
and U105 (N_105,In_1236,In_213);
and U106 (N_106,In_168,In_808);
nor U107 (N_107,In_404,In_348);
or U108 (N_108,In_972,In_194);
or U109 (N_109,In_549,In_309);
or U110 (N_110,In_906,In_950);
or U111 (N_111,In_1141,In_459);
and U112 (N_112,In_250,In_603);
nor U113 (N_113,In_73,In_166);
nor U114 (N_114,In_1243,In_853);
nor U115 (N_115,In_268,In_977);
and U116 (N_116,In_1093,In_422);
nand U117 (N_117,In_920,In_1498);
or U118 (N_118,In_930,In_1299);
or U119 (N_119,In_502,In_1056);
and U120 (N_120,In_867,In_372);
or U121 (N_121,In_1344,In_622);
or U122 (N_122,In_347,In_1361);
or U123 (N_123,In_953,In_98);
nor U124 (N_124,In_866,In_1166);
nand U125 (N_125,In_705,In_992);
xnor U126 (N_126,In_1396,In_478);
or U127 (N_127,In_1209,In_485);
nor U128 (N_128,In_556,In_226);
nor U129 (N_129,In_1062,In_833);
or U130 (N_130,In_785,In_499);
nor U131 (N_131,In_684,In_607);
or U132 (N_132,In_775,In_698);
nand U133 (N_133,In_1115,In_1224);
nor U134 (N_134,In_524,In_955);
and U135 (N_135,In_1024,In_749);
xnor U136 (N_136,In_42,In_89);
nand U137 (N_137,In_1332,In_420);
nor U138 (N_138,In_183,In_1038);
or U139 (N_139,In_1245,In_1068);
and U140 (N_140,In_389,In_16);
nand U141 (N_141,In_416,In_124);
and U142 (N_142,In_761,In_1457);
and U143 (N_143,In_725,In_1278);
nand U144 (N_144,In_25,In_142);
nor U145 (N_145,In_236,In_858);
nor U146 (N_146,In_169,In_503);
and U147 (N_147,In_703,In_71);
xnor U148 (N_148,In_767,In_1406);
and U149 (N_149,In_1110,In_285);
and U150 (N_150,In_1478,In_40);
and U151 (N_151,In_184,In_629);
or U152 (N_152,In_1374,In_428);
nand U153 (N_153,In_1466,In_24);
nand U154 (N_154,In_289,In_1420);
or U155 (N_155,In_1156,In_1369);
or U156 (N_156,In_810,In_511);
nand U157 (N_157,In_1137,In_162);
nand U158 (N_158,In_215,In_577);
or U159 (N_159,In_545,In_1413);
or U160 (N_160,In_819,In_448);
nand U161 (N_161,In_1009,In_246);
nor U162 (N_162,In_681,In_753);
nand U163 (N_163,In_130,In_431);
or U164 (N_164,In_18,In_864);
nand U165 (N_165,In_457,In_733);
and U166 (N_166,In_580,In_266);
or U167 (N_167,In_862,In_247);
or U168 (N_168,In_803,In_831);
nand U169 (N_169,In_212,In_846);
nand U170 (N_170,In_498,In_490);
or U171 (N_171,In_1222,In_86);
nand U172 (N_172,In_112,In_871);
and U173 (N_173,In_177,In_911);
nand U174 (N_174,In_219,In_63);
and U175 (N_175,In_996,In_191);
nor U176 (N_176,In_1162,In_223);
xnor U177 (N_177,In_196,In_1240);
nand U178 (N_178,In_717,In_658);
nor U179 (N_179,In_1006,In_5);
or U180 (N_180,In_1289,In_401);
nor U181 (N_181,In_384,In_225);
or U182 (N_182,In_1302,In_652);
nor U183 (N_183,In_176,In_252);
nor U184 (N_184,In_1336,In_295);
nand U185 (N_185,In_1237,In_325);
nand U186 (N_186,In_558,In_949);
and U187 (N_187,In_415,In_107);
nor U188 (N_188,In_460,In_1312);
and U189 (N_189,In_974,In_1303);
and U190 (N_190,In_903,In_1407);
and U191 (N_191,In_33,In_852);
nor U192 (N_192,In_520,In_878);
nor U193 (N_193,In_640,In_1261);
nor U194 (N_194,In_921,In_345);
or U195 (N_195,In_762,In_786);
or U196 (N_196,In_83,In_1091);
nor U197 (N_197,In_195,In_1170);
and U198 (N_198,In_989,In_1395);
nor U199 (N_199,In_1231,In_807);
nor U200 (N_200,In_1244,In_678);
nor U201 (N_201,In_1003,In_897);
xor U202 (N_202,In_901,In_886);
xnor U203 (N_203,In_12,In_34);
nor U204 (N_204,In_994,In_1184);
nor U205 (N_205,In_262,In_744);
and U206 (N_206,In_328,In_1376);
nand U207 (N_207,In_614,In_943);
nor U208 (N_208,In_494,In_1015);
or U209 (N_209,In_185,In_155);
or U210 (N_210,In_197,In_68);
or U211 (N_211,In_1393,In_952);
and U212 (N_212,In_541,In_776);
nand U213 (N_213,In_392,In_602);
and U214 (N_214,In_1228,In_1260);
or U215 (N_215,In_590,In_528);
nand U216 (N_216,In_413,In_889);
and U217 (N_217,In_1356,In_1185);
or U218 (N_218,In_982,In_257);
nor U219 (N_219,In_896,In_1463);
nand U220 (N_220,In_229,In_116);
xor U221 (N_221,In_1161,In_760);
or U222 (N_222,In_563,In_376);
or U223 (N_223,In_1086,In_584);
nor U224 (N_224,In_399,In_1113);
nand U225 (N_225,In_665,In_530);
nand U226 (N_226,In_505,In_1028);
nand U227 (N_227,In_1355,In_364);
or U228 (N_228,In_397,In_1386);
nand U229 (N_229,In_1121,In_153);
nand U230 (N_230,In_566,In_1410);
or U231 (N_231,In_1308,In_164);
nand U232 (N_232,In_128,In_1223);
or U233 (N_233,In_114,In_517);
and U234 (N_234,In_1114,In_332);
or U235 (N_235,In_84,In_260);
and U236 (N_236,In_661,In_1098);
nand U237 (N_237,In_296,In_795);
nand U238 (N_238,In_1189,In_1083);
nand U239 (N_239,In_1415,In_206);
or U240 (N_240,In_904,In_961);
nand U241 (N_241,In_189,In_145);
and U242 (N_242,In_363,In_38);
xnor U243 (N_243,In_55,In_47);
nor U244 (N_244,In_403,In_547);
nand U245 (N_245,In_1153,In_1010);
nand U246 (N_246,In_440,In_1268);
and U247 (N_247,In_385,In_15);
xnor U248 (N_248,In_1408,In_927);
nor U249 (N_249,In_529,In_641);
and U250 (N_250,In_631,In_694);
or U251 (N_251,In_342,In_146);
nor U252 (N_252,In_248,In_242);
and U253 (N_253,In_706,In_1047);
nor U254 (N_254,In_429,In_1424);
xnor U255 (N_255,In_532,In_693);
and U256 (N_256,In_1030,In_276);
nor U257 (N_257,In_1078,In_1342);
nand U258 (N_258,In_1349,In_233);
nand U259 (N_259,In_497,In_165);
or U260 (N_260,In_314,In_504);
or U261 (N_261,In_1283,In_41);
or U262 (N_262,In_1033,In_424);
or U263 (N_263,In_1437,In_710);
nor U264 (N_264,In_870,In_96);
nor U265 (N_265,In_540,In_1469);
nand U266 (N_266,In_1317,In_278);
nor U267 (N_267,In_57,In_1057);
or U268 (N_268,In_533,In_1247);
or U269 (N_269,In_1270,In_1058);
nor U270 (N_270,In_888,In_1474);
or U271 (N_271,In_208,In_849);
nor U272 (N_272,In_842,In_680);
nor U273 (N_273,In_809,In_724);
or U274 (N_274,In_74,In_635);
nor U275 (N_275,In_368,In_1436);
xnor U276 (N_276,In_35,In_1096);
nor U277 (N_277,In_337,In_1337);
xor U278 (N_278,In_1042,In_1453);
or U279 (N_279,In_1398,In_653);
or U280 (N_280,In_453,In_723);
or U281 (N_281,In_539,In_349);
nor U282 (N_282,In_425,In_192);
and U283 (N_283,In_627,In_1272);
nand U284 (N_284,In_418,In_525);
nand U285 (N_285,In_1150,In_139);
nor U286 (N_286,In_1271,In_959);
or U287 (N_287,In_1233,In_370);
and U288 (N_288,In_1133,In_1132);
nor U289 (N_289,In_615,In_1476);
nor U290 (N_290,In_270,In_95);
xnor U291 (N_291,In_1120,In_264);
xor U292 (N_292,In_76,In_991);
nor U293 (N_293,In_50,In_979);
xor U294 (N_294,In_674,In_600);
or U295 (N_295,In_769,In_971);
nand U296 (N_296,In_1488,In_1370);
or U297 (N_297,In_472,In_620);
and U298 (N_298,In_1206,In_571);
xor U299 (N_299,In_1384,In_1215);
nand U300 (N_300,In_765,In_210);
nor U301 (N_301,In_656,In_136);
nor U302 (N_302,In_891,In_294);
and U303 (N_303,In_393,In_1340);
and U304 (N_304,In_85,In_567);
nor U305 (N_305,In_609,In_1490);
or U306 (N_306,In_152,In_412);
nand U307 (N_307,In_1004,In_72);
nor U308 (N_308,In_1059,In_175);
and U309 (N_309,In_414,In_1387);
nand U310 (N_310,In_1036,In_352);
and U311 (N_311,In_1414,In_829);
xor U312 (N_312,In_737,In_675);
or U313 (N_313,In_1404,In_893);
or U314 (N_314,In_1275,In_65);
nor U315 (N_315,In_391,In_964);
and U316 (N_316,In_721,In_1473);
xor U317 (N_317,In_265,In_514);
xnor U318 (N_318,In_882,In_1446);
xnor U319 (N_319,In_667,In_779);
nand U320 (N_320,In_797,In_1050);
nor U321 (N_321,In_437,In_1242);
nand U322 (N_322,In_1373,In_1338);
nor U323 (N_323,In_1354,In_1251);
or U324 (N_324,In_303,In_1158);
or U325 (N_325,In_1266,In_316);
nand U326 (N_326,In_1296,In_1160);
nor U327 (N_327,In_103,In_147);
xor U328 (N_328,In_845,In_1419);
nor U329 (N_329,In_969,In_69);
and U330 (N_330,In_1172,In_117);
nand U331 (N_331,In_946,In_787);
and U332 (N_332,In_638,In_1140);
or U333 (N_333,In_477,In_1152);
or U334 (N_334,In_1131,In_1031);
nor U335 (N_335,In_90,In_788);
xnor U336 (N_336,In_1040,In_824);
nand U337 (N_337,In_1220,In_1427);
nand U338 (N_338,In_406,In_944);
and U339 (N_339,In_426,In_306);
nor U340 (N_340,In_435,In_919);
and U341 (N_341,In_1151,In_884);
nor U342 (N_342,In_840,In_1046);
and U343 (N_343,In_1100,In_492);
or U344 (N_344,In_259,In_1138);
and U345 (N_345,In_967,In_553);
and U346 (N_346,In_975,In_1147);
nand U347 (N_347,In_284,In_1210);
nand U348 (N_348,In_1200,In_452);
nand U349 (N_349,In_463,In_1329);
nand U350 (N_350,In_1442,In_489);
or U351 (N_351,In_782,In_993);
or U352 (N_352,In_410,In_127);
and U353 (N_353,In_402,In_679);
and U354 (N_354,In_758,In_1403);
and U355 (N_355,In_557,In_757);
and U356 (N_356,In_481,In_1092);
nor U357 (N_357,In_1322,In_910);
and U358 (N_358,In_608,In_432);
or U359 (N_359,In_918,In_986);
nor U360 (N_360,In_669,In_713);
and U361 (N_361,In_814,In_588);
xor U362 (N_362,In_654,In_1315);
and U363 (N_363,In_1495,In_327);
and U364 (N_364,In_1134,In_411);
or U365 (N_365,In_1399,In_214);
nor U366 (N_366,In_379,In_682);
nor U367 (N_367,In_17,In_565);
and U368 (N_368,In_855,In_173);
nand U369 (N_369,In_1014,In_230);
or U370 (N_370,In_720,In_220);
nor U371 (N_371,In_315,In_171);
or U372 (N_372,In_67,In_417);
xor U373 (N_373,In_222,In_450);
or U374 (N_374,In_37,In_1380);
nor U375 (N_375,In_909,In_1418);
and U376 (N_376,In_436,In_507);
or U377 (N_377,In_655,In_1105);
nor U378 (N_378,In_1194,In_395);
and U379 (N_379,In_279,In_672);
nor U380 (N_380,In_677,In_58);
nor U381 (N_381,In_646,In_887);
nand U382 (N_382,In_912,In_1323);
or U383 (N_383,In_1411,In_156);
and U384 (N_384,In_823,In_121);
or U385 (N_385,In_643,In_709);
or U386 (N_386,In_351,In_28);
nand U387 (N_387,In_1084,In_108);
or U388 (N_388,In_1367,In_1005);
or U389 (N_389,In_649,In_1087);
nand U390 (N_390,In_1346,In_1345);
xnor U391 (N_391,In_1168,In_1081);
xor U392 (N_392,In_589,In_456);
or U393 (N_393,In_1023,In_960);
and U394 (N_394,In_228,In_818);
and U395 (N_395,In_267,In_1227);
nand U396 (N_396,In_466,In_200);
nand U397 (N_397,In_1017,In_275);
nand U398 (N_398,In_1280,In_441);
and U399 (N_399,In_1269,In_234);
or U400 (N_400,In_102,In_1477);
or U401 (N_401,In_990,In_741);
and U402 (N_402,In_1039,In_125);
nand U403 (N_403,In_894,In_1318);
nand U404 (N_404,In_468,In_1021);
and U405 (N_405,In_1381,In_770);
or U406 (N_406,In_1428,In_1309);
nand U407 (N_407,In_825,In_487);
and U408 (N_408,In_39,In_759);
nand U409 (N_409,In_1129,In_863);
xnor U410 (N_410,In_369,In_1310);
nand U411 (N_411,In_722,In_1348);
and U412 (N_412,In_1255,In_340);
nand U413 (N_413,In_873,In_465);
nor U414 (N_414,In_997,In_872);
or U415 (N_415,In_963,In_1281);
and U416 (N_416,In_1365,In_581);
and U417 (N_417,In_1252,In_716);
and U418 (N_418,In_339,In_1000);
nor U419 (N_419,In_97,In_890);
and U420 (N_420,In_604,In_687);
nor U421 (N_421,In_31,In_1433);
or U422 (N_422,In_597,In_300);
nand U423 (N_423,In_1067,In_1402);
and U424 (N_424,In_1383,In_1274);
xor U425 (N_425,In_1298,In_606);
nand U426 (N_426,In_1095,In_1470);
or U427 (N_427,In_292,In_695);
or U428 (N_428,In_1287,In_1079);
nor U429 (N_429,In_555,In_36);
nor U430 (N_430,In_1127,In_790);
nand U431 (N_431,In_1364,In_1363);
nor U432 (N_432,In_815,In_1108);
and U433 (N_433,In_881,In_198);
nand U434 (N_434,In_1226,In_1123);
nand U435 (N_435,In_1066,In_613);
or U436 (N_436,In_596,In_1094);
and U437 (N_437,In_784,In_282);
xor U438 (N_438,In_923,In_45);
nor U439 (N_439,In_205,In_582);
or U440 (N_440,In_199,In_458);
nand U441 (N_441,In_1016,In_748);
and U442 (N_442,In_1456,In_1122);
or U443 (N_443,In_718,In_544);
xnor U444 (N_444,In_54,In_1439);
or U445 (N_445,In_1052,In_1430);
and U446 (N_446,In_907,In_154);
and U447 (N_447,In_670,In_780);
and U448 (N_448,In_902,In_1148);
or U449 (N_449,In_877,In_594);
and U450 (N_450,In_980,In_1136);
or U451 (N_451,In_471,In_249);
nor U452 (N_452,In_204,In_1479);
nand U453 (N_453,In_256,In_1064);
nand U454 (N_454,In_711,In_916);
or U455 (N_455,In_728,In_995);
nand U456 (N_456,In_579,In_151);
or U457 (N_457,In_1082,In_484);
nand U458 (N_458,In_1316,In_999);
nand U459 (N_459,In_1450,In_929);
nor U460 (N_460,In_1065,In_601);
xnor U461 (N_461,In_1019,In_1103);
nor U462 (N_462,In_1008,In_983);
nand U463 (N_463,In_885,In_132);
xor U464 (N_464,In_1035,In_962);
nand U465 (N_465,In_1195,In_52);
nand U466 (N_466,In_578,In_801);
and U467 (N_467,In_648,In_461);
nand U468 (N_468,In_1011,In_64);
and U469 (N_469,In_933,In_636);
and U470 (N_470,In_719,In_1265);
nor U471 (N_471,In_1022,In_612);
nor U472 (N_472,In_1119,In_48);
nand U473 (N_473,In_131,In_1051);
or U474 (N_474,In_1032,In_1273);
or U475 (N_475,In_181,In_1441);
and U476 (N_476,In_1371,In_1491);
and U477 (N_477,In_805,In_271);
xnor U478 (N_478,In_280,In_1106);
nand U479 (N_479,In_305,In_671);
or U480 (N_480,In_617,In_1175);
and U481 (N_481,In_522,In_143);
and U482 (N_482,In_1480,In_751);
nand U483 (N_483,In_1196,In_60);
and U484 (N_484,In_1135,In_985);
nor U485 (N_485,In_1104,In_287);
nor U486 (N_486,In_263,In_1186);
nand U487 (N_487,In_798,In_576);
nor U488 (N_488,In_433,In_1494);
xnor U489 (N_489,In_830,In_1054);
nand U490 (N_490,In_150,In_1241);
and U491 (N_491,In_662,In_905);
nor U492 (N_492,In_331,In_1276);
xor U493 (N_493,In_1385,In_1063);
nand U494 (N_494,In_925,In_137);
or U495 (N_495,In_355,In_396);
or U496 (N_496,In_133,In_947);
or U497 (N_497,In_794,In_875);
xnor U498 (N_498,In_93,In_449);
or U499 (N_499,In_157,In_1178);
or U500 (N_500,In_1468,In_1163);
nor U501 (N_501,In_804,In_1258);
or U502 (N_502,In_1125,In_939);
and U503 (N_503,In_1499,In_1282);
or U504 (N_504,In_1191,In_358);
or U505 (N_505,In_398,In_381);
xnor U506 (N_506,In_938,In_187);
and U507 (N_507,In_366,In_847);
and U508 (N_508,In_1305,In_543);
nand U509 (N_509,In_274,In_421);
and U510 (N_510,In_756,In_1044);
xnor U511 (N_511,In_771,In_299);
and U512 (N_512,In_928,In_1048);
or U513 (N_513,In_464,In_811);
nor U514 (N_514,In_174,In_651);
nor U515 (N_515,In_1177,In_298);
xnor U516 (N_516,In_1357,In_932);
and U517 (N_517,In_712,In_518);
nor U518 (N_518,In_482,In_686);
and U519 (N_519,In_568,In_630);
nor U520 (N_520,In_75,In_80);
and U521 (N_521,In_159,In_1213);
and U522 (N_522,In_488,In_1143);
nor U523 (N_523,In_632,In_1146);
nor U524 (N_524,In_1327,In_237);
nor U525 (N_525,In_474,In_1029);
nor U526 (N_526,In_1405,In_1300);
and U527 (N_527,In_550,In_321);
and U528 (N_528,In_1165,In_10);
or U529 (N_529,In_735,In_1257);
xor U530 (N_530,In_650,In_335);
or U531 (N_531,In_451,In_29);
nand U532 (N_532,In_1130,In_324);
nand U533 (N_533,In_46,In_1295);
nor U534 (N_534,In_752,In_1203);
nor U535 (N_535,In_826,In_180);
or U536 (N_536,In_745,In_167);
or U537 (N_537,In_583,In_702);
and U538 (N_538,In_110,In_258);
nand U539 (N_539,In_129,In_1263);
nand U540 (N_540,In_519,In_561);
xor U541 (N_541,In_813,In_800);
and U542 (N_542,In_49,In_14);
or U543 (N_543,In_1360,In_1306);
nor U544 (N_544,In_1117,In_1214);
nor U545 (N_545,In_1197,In_111);
xor U546 (N_546,In_708,In_243);
xnor U547 (N_547,In_739,In_297);
nand U548 (N_548,In_978,In_405);
and U549 (N_549,In_344,In_1335);
nand U550 (N_550,In_23,In_323);
nand U551 (N_551,In_1116,In_119);
or U552 (N_552,In_508,In_343);
nor U553 (N_553,In_1077,In_965);
or U554 (N_554,In_1045,In_1409);
xnor U555 (N_555,In_951,In_850);
nor U556 (N_556,In_865,In_1390);
or U557 (N_557,In_1205,In_1199);
and U558 (N_558,In_740,In_318);
or U559 (N_559,In_56,In_1400);
and U560 (N_560,In_231,In_386);
nor U561 (N_561,In_281,In_11);
or U562 (N_562,In_689,In_360);
nor U563 (N_563,In_908,In_1070);
or U564 (N_564,In_1465,In_1102);
nand U565 (N_565,In_1334,In_1076);
nor U566 (N_566,In_746,In_1467);
or U567 (N_567,In_876,In_874);
and U568 (N_568,In_747,In_1451);
or U569 (N_569,In_1176,In_1464);
nand U570 (N_570,In_812,In_9);
xnor U571 (N_571,In_475,In_956);
and U572 (N_572,In_537,In_1471);
and U573 (N_573,In_144,In_483);
xor U574 (N_574,In_696,In_51);
nor U575 (N_575,In_1331,In_91);
and U576 (N_576,In_1320,In_572);
or U577 (N_577,In_1232,In_559);
and U578 (N_578,In_1294,In_736);
or U579 (N_579,In_1182,In_515);
nand U580 (N_580,In_462,In_387);
or U581 (N_581,In_592,In_937);
and U582 (N_582,In_1307,In_1181);
or U583 (N_583,In_444,In_754);
nand U584 (N_584,In_241,In_1290);
and U585 (N_585,In_350,In_1392);
nand U586 (N_586,In_140,In_1164);
or U587 (N_587,In_1107,In_859);
and U588 (N_588,In_138,In_610);
nor U589 (N_589,In_729,In_322);
xnor U590 (N_590,In_1018,In_1043);
nor U591 (N_591,In_697,In_1455);
nand U592 (N_592,In_1483,In_560);
or U593 (N_593,In_922,In_1207);
or U594 (N_594,In_586,In_1037);
or U595 (N_595,In_1055,In_1482);
nand U596 (N_596,In_496,In_676);
and U597 (N_597,In_704,In_637);
or U598 (N_598,In_1487,In_126);
nor U599 (N_599,In_998,In_1001);
nand U600 (N_600,In_738,In_244);
nand U601 (N_601,In_573,In_509);
and U602 (N_602,In_1362,In_668);
or U603 (N_603,In_954,In_913);
xor U604 (N_604,In_356,In_491);
xnor U605 (N_605,In_659,In_1378);
nand U606 (N_606,In_1074,In_493);
and U607 (N_607,In_288,In_1313);
or U608 (N_608,In_914,In_1301);
nand U609 (N_609,In_1060,In_371);
and U610 (N_610,In_892,In_1219);
nor U611 (N_611,In_777,In_455);
or U612 (N_612,In_1126,In_120);
or U613 (N_613,In_1292,In_320);
or U614 (N_614,In_1239,In_538);
xor U615 (N_615,In_148,In_1155);
nand U616 (N_616,In_161,In_81);
nor U617 (N_617,In_470,In_1422);
nor U618 (N_618,In_1109,In_1025);
or U619 (N_619,In_239,In_848);
nand U620 (N_620,In_203,In_837);
or U621 (N_621,In_841,In_326);
and U622 (N_622,In_476,In_227);
and U623 (N_623,In_1049,In_715);
xor U624 (N_624,In_598,In_1149);
xnor U625 (N_625,In_1073,In_211);
xor U626 (N_626,In_430,In_832);
nor U627 (N_627,In_1253,In_883);
or U628 (N_628,In_141,In_789);
or U629 (N_629,In_1099,In_238);
nand U630 (N_630,In_1111,In_926);
nand U631 (N_631,In_1440,In_361);
xnor U632 (N_632,In_20,In_714);
or U633 (N_633,In_1179,In_273);
nor U634 (N_634,In_727,In_799);
nand U635 (N_635,In_467,In_1034);
nor U636 (N_636,In_743,In_302);
xnor U637 (N_637,In_917,In_1351);
nand U638 (N_638,In_1053,In_0);
nand U639 (N_639,In_1225,In_1235);
and U640 (N_640,In_1443,In_1174);
or U641 (N_641,In_1284,In_179);
nand U642 (N_642,In_828,In_88);
and U643 (N_643,In_346,In_1434);
and U644 (N_644,In_22,In_1460);
and U645 (N_645,In_61,In_699);
nor U646 (N_646,In_898,In_382);
nor U647 (N_647,In_101,In_1401);
nand U648 (N_648,In_1211,In_1485);
nor U649 (N_649,In_1421,In_21);
nor U650 (N_650,In_480,In_1013);
xnor U651 (N_651,In_1267,In_1454);
and U652 (N_652,In_899,In_394);
nand U653 (N_653,In_1159,In_254);
nand U654 (N_654,In_1426,In_1020);
nand U655 (N_655,In_1097,In_755);
nand U656 (N_656,In_634,In_109);
or U657 (N_657,In_1324,In_4);
nor U658 (N_658,In_43,In_312);
and U659 (N_659,In_269,In_984);
nor U660 (N_660,In_768,In_329);
or U661 (N_661,In_1221,In_1366);
or U662 (N_662,In_1297,In_645);
nand U663 (N_663,In_1375,In_595);
nor U664 (N_664,In_1382,In_611);
nor U665 (N_665,In_336,In_78);
nor U666 (N_666,In_773,In_536);
xor U667 (N_667,In_26,In_1259);
nand U668 (N_668,In_512,In_1389);
or U669 (N_669,In_778,In_1472);
nor U670 (N_670,In_987,In_948);
and U671 (N_671,In_1497,In_333);
or U672 (N_672,In_224,In_1041);
nor U673 (N_673,In_562,In_500);
nor U674 (N_674,In_660,In_1412);
nor U675 (N_675,In_378,In_1397);
and U676 (N_676,In_575,In_742);
nor U677 (N_677,In_19,In_1314);
and U678 (N_678,In_968,In_843);
or U679 (N_679,In_510,In_495);
nand U680 (N_680,In_407,In_1192);
nor U681 (N_681,In_106,In_931);
nor U682 (N_682,In_1291,In_1075);
nor U683 (N_683,In_666,In_188);
nand U684 (N_684,In_201,In_1353);
nor U685 (N_685,In_100,In_940);
nor U686 (N_686,In_701,In_30);
or U687 (N_687,In_1190,In_1377);
xnor U688 (N_688,In_390,In_1249);
nand U689 (N_689,In_1452,In_625);
xnor U690 (N_690,In_310,In_1475);
or U691 (N_691,In_158,In_209);
nor U692 (N_692,In_186,In_587);
xor U693 (N_693,In_836,In_1445);
or U694 (N_694,In_365,In_1489);
and U695 (N_695,In_673,In_1124);
or U696 (N_696,In_104,In_301);
or U697 (N_697,In_621,In_190);
nor U698 (N_698,In_564,In_935);
and U699 (N_699,In_1071,In_308);
or U700 (N_700,In_1157,In_182);
nand U701 (N_701,In_163,In_593);
nor U702 (N_702,In_1208,In_367);
or U703 (N_703,In_1379,In_647);
xnor U704 (N_704,In_79,In_1341);
xor U705 (N_705,In_1027,In_1423);
and U706 (N_706,In_1319,In_664);
nor U707 (N_707,In_1007,In_857);
and U708 (N_708,In_683,In_8);
or U709 (N_709,In_1486,In_552);
and U710 (N_710,In_419,In_439);
and U711 (N_711,In_2,In_860);
nand U712 (N_712,In_330,In_1432);
nor U713 (N_713,In_1193,In_134);
nor U714 (N_714,In_438,In_1286);
nor U715 (N_715,In_1304,In_988);
nand U716 (N_716,In_377,In_1325);
nand U717 (N_717,In_291,In_53);
and U718 (N_718,In_442,In_936);
nand U719 (N_719,In_554,In_44);
or U720 (N_720,In_217,In_1169);
nand U721 (N_721,In_221,In_1216);
and U722 (N_722,In_87,In_1429);
and U723 (N_723,In_934,In_1493);
or U724 (N_724,In_726,In_105);
and U725 (N_725,In_806,In_172);
and U726 (N_726,In_895,In_1416);
xnor U727 (N_727,In_32,In_838);
or U728 (N_728,In_240,In_400);
nand U729 (N_729,In_1459,In_1);
nor U730 (N_730,In_1230,In_551);
and U731 (N_731,In_1417,In_99);
nor U732 (N_732,In_1201,In_585);
or U733 (N_733,In_362,In_599);
nor U734 (N_734,In_802,In_1145);
nand U735 (N_735,In_834,In_1112);
and U736 (N_736,In_92,In_707);
nor U737 (N_737,In_783,In_232);
nor U738 (N_738,In_869,In_817);
nor U739 (N_739,In_542,In_1492);
xor U740 (N_740,In_245,In_1496);
nor U741 (N_741,In_854,In_1285);
nand U742 (N_742,In_290,In_526);
nand U743 (N_743,In_255,In_501);
or U744 (N_744,In_791,In_1388);
and U745 (N_745,In_235,In_732);
and U746 (N_746,In_1069,In_1444);
nand U747 (N_747,In_375,In_506);
nor U748 (N_748,In_6,In_851);
or U749 (N_749,In_861,In_1229);
nor U750 (N_750,In_345,In_67);
nand U751 (N_751,In_1423,In_941);
nand U752 (N_752,In_1241,In_303);
nor U753 (N_753,In_933,In_771);
nand U754 (N_754,In_19,In_821);
or U755 (N_755,In_139,In_175);
nand U756 (N_756,In_1070,In_668);
nor U757 (N_757,In_417,In_697);
nor U758 (N_758,In_1333,In_1327);
nor U759 (N_759,In_1318,In_1362);
nand U760 (N_760,In_723,In_210);
xnor U761 (N_761,In_718,In_271);
or U762 (N_762,In_1276,In_973);
nor U763 (N_763,In_1211,In_884);
or U764 (N_764,In_288,In_803);
and U765 (N_765,In_1441,In_465);
xor U766 (N_766,In_1465,In_209);
nand U767 (N_767,In_182,In_554);
nor U768 (N_768,In_391,In_430);
nor U769 (N_769,In_229,In_171);
or U770 (N_770,In_1346,In_507);
and U771 (N_771,In_417,In_235);
nor U772 (N_772,In_1357,In_1130);
nand U773 (N_773,In_1262,In_129);
nor U774 (N_774,In_833,In_516);
xnor U775 (N_775,In_836,In_477);
nor U776 (N_776,In_115,In_1354);
or U777 (N_777,In_17,In_1369);
and U778 (N_778,In_939,In_832);
or U779 (N_779,In_1052,In_250);
nor U780 (N_780,In_1212,In_483);
nor U781 (N_781,In_1463,In_1064);
xnor U782 (N_782,In_244,In_781);
and U783 (N_783,In_188,In_1436);
and U784 (N_784,In_145,In_486);
nor U785 (N_785,In_214,In_1496);
nand U786 (N_786,In_304,In_1406);
and U787 (N_787,In_1051,In_261);
nor U788 (N_788,In_1495,In_11);
and U789 (N_789,In_1031,In_1321);
and U790 (N_790,In_903,In_1415);
nand U791 (N_791,In_686,In_1361);
nand U792 (N_792,In_772,In_416);
nand U793 (N_793,In_455,In_339);
and U794 (N_794,In_645,In_1258);
or U795 (N_795,In_987,In_508);
nor U796 (N_796,In_1124,In_1308);
nand U797 (N_797,In_609,In_194);
and U798 (N_798,In_1362,In_913);
or U799 (N_799,In_1456,In_700);
and U800 (N_800,In_477,In_110);
or U801 (N_801,In_242,In_1429);
and U802 (N_802,In_1252,In_554);
and U803 (N_803,In_392,In_368);
or U804 (N_804,In_527,In_272);
or U805 (N_805,In_1199,In_1484);
or U806 (N_806,In_803,In_194);
and U807 (N_807,In_363,In_1230);
nand U808 (N_808,In_1429,In_1021);
nor U809 (N_809,In_108,In_1407);
and U810 (N_810,In_1230,In_923);
or U811 (N_811,In_45,In_392);
nor U812 (N_812,In_723,In_1171);
nand U813 (N_813,In_96,In_1072);
nand U814 (N_814,In_667,In_942);
nand U815 (N_815,In_1183,In_1239);
nor U816 (N_816,In_357,In_110);
nand U817 (N_817,In_806,In_453);
or U818 (N_818,In_1288,In_491);
or U819 (N_819,In_126,In_233);
nor U820 (N_820,In_94,In_1208);
nand U821 (N_821,In_995,In_84);
and U822 (N_822,In_1020,In_618);
xor U823 (N_823,In_1464,In_1381);
or U824 (N_824,In_566,In_1329);
or U825 (N_825,In_868,In_1214);
nor U826 (N_826,In_782,In_280);
nor U827 (N_827,In_139,In_419);
or U828 (N_828,In_225,In_1320);
and U829 (N_829,In_761,In_1365);
or U830 (N_830,In_132,In_1078);
nand U831 (N_831,In_629,In_1304);
xor U832 (N_832,In_417,In_956);
nand U833 (N_833,In_1351,In_808);
xnor U834 (N_834,In_772,In_421);
nand U835 (N_835,In_573,In_1457);
nor U836 (N_836,In_133,In_1342);
and U837 (N_837,In_891,In_1064);
xor U838 (N_838,In_1229,In_254);
xor U839 (N_839,In_225,In_591);
nand U840 (N_840,In_93,In_758);
nor U841 (N_841,In_646,In_633);
xor U842 (N_842,In_918,In_1081);
and U843 (N_843,In_1002,In_467);
or U844 (N_844,In_774,In_899);
and U845 (N_845,In_644,In_173);
or U846 (N_846,In_1359,In_1111);
xor U847 (N_847,In_97,In_204);
xor U848 (N_848,In_998,In_1097);
xor U849 (N_849,In_1042,In_1117);
and U850 (N_850,In_1001,In_359);
nand U851 (N_851,In_1206,In_434);
nor U852 (N_852,In_446,In_1483);
nand U853 (N_853,In_1089,In_662);
or U854 (N_854,In_53,In_855);
xnor U855 (N_855,In_430,In_964);
nand U856 (N_856,In_1176,In_1118);
or U857 (N_857,In_861,In_491);
and U858 (N_858,In_443,In_635);
and U859 (N_859,In_557,In_395);
nand U860 (N_860,In_595,In_97);
or U861 (N_861,In_505,In_835);
xor U862 (N_862,In_1367,In_1056);
and U863 (N_863,In_230,In_179);
and U864 (N_864,In_127,In_1453);
nand U865 (N_865,In_909,In_979);
and U866 (N_866,In_967,In_1001);
or U867 (N_867,In_978,In_1072);
or U868 (N_868,In_720,In_1459);
and U869 (N_869,In_46,In_435);
nand U870 (N_870,In_1003,In_991);
nor U871 (N_871,In_450,In_833);
nor U872 (N_872,In_427,In_898);
or U873 (N_873,In_773,In_1167);
and U874 (N_874,In_949,In_1190);
nor U875 (N_875,In_646,In_237);
or U876 (N_876,In_863,In_1373);
nand U877 (N_877,In_579,In_619);
and U878 (N_878,In_738,In_75);
or U879 (N_879,In_1409,In_288);
and U880 (N_880,In_255,In_621);
or U881 (N_881,In_600,In_192);
nor U882 (N_882,In_942,In_1310);
nand U883 (N_883,In_598,In_443);
and U884 (N_884,In_931,In_1304);
nand U885 (N_885,In_568,In_1009);
or U886 (N_886,In_516,In_543);
xnor U887 (N_887,In_204,In_193);
or U888 (N_888,In_1241,In_400);
nand U889 (N_889,In_1309,In_176);
nand U890 (N_890,In_1333,In_1024);
nand U891 (N_891,In_243,In_892);
nor U892 (N_892,In_838,In_285);
nand U893 (N_893,In_1398,In_759);
and U894 (N_894,In_1222,In_1411);
or U895 (N_895,In_1223,In_776);
and U896 (N_896,In_529,In_564);
nand U897 (N_897,In_1174,In_151);
nand U898 (N_898,In_1110,In_368);
and U899 (N_899,In_927,In_339);
or U900 (N_900,In_851,In_767);
xor U901 (N_901,In_820,In_602);
nor U902 (N_902,In_962,In_364);
or U903 (N_903,In_846,In_514);
and U904 (N_904,In_1387,In_1448);
nand U905 (N_905,In_329,In_340);
or U906 (N_906,In_683,In_1168);
and U907 (N_907,In_1493,In_1451);
nor U908 (N_908,In_143,In_1345);
nand U909 (N_909,In_1194,In_754);
and U910 (N_910,In_246,In_1357);
nand U911 (N_911,In_1001,In_239);
or U912 (N_912,In_1336,In_1389);
xnor U913 (N_913,In_39,In_1402);
nor U914 (N_914,In_1076,In_111);
nand U915 (N_915,In_919,In_953);
nand U916 (N_916,In_1256,In_1174);
xor U917 (N_917,In_1206,In_708);
nor U918 (N_918,In_358,In_188);
nand U919 (N_919,In_1042,In_1039);
nand U920 (N_920,In_1055,In_1427);
nand U921 (N_921,In_625,In_423);
and U922 (N_922,In_1109,In_951);
or U923 (N_923,In_17,In_612);
or U924 (N_924,In_117,In_1027);
or U925 (N_925,In_1227,In_318);
nand U926 (N_926,In_182,In_277);
or U927 (N_927,In_711,In_1242);
or U928 (N_928,In_840,In_388);
or U929 (N_929,In_126,In_376);
and U930 (N_930,In_1270,In_447);
or U931 (N_931,In_430,In_1164);
nand U932 (N_932,In_285,In_963);
nand U933 (N_933,In_1010,In_1435);
or U934 (N_934,In_1008,In_283);
and U935 (N_935,In_521,In_668);
nor U936 (N_936,In_34,In_1457);
nand U937 (N_937,In_349,In_407);
or U938 (N_938,In_1429,In_951);
and U939 (N_939,In_163,In_1452);
and U940 (N_940,In_525,In_1036);
and U941 (N_941,In_159,In_325);
and U942 (N_942,In_1064,In_1213);
nand U943 (N_943,In_161,In_1011);
and U944 (N_944,In_46,In_69);
nand U945 (N_945,In_1348,In_168);
and U946 (N_946,In_1182,In_1042);
nand U947 (N_947,In_559,In_943);
nor U948 (N_948,In_396,In_216);
nor U949 (N_949,In_834,In_982);
nor U950 (N_950,In_994,In_105);
nor U951 (N_951,In_1223,In_1234);
nor U952 (N_952,In_686,In_868);
or U953 (N_953,In_549,In_1369);
nand U954 (N_954,In_1008,In_21);
nor U955 (N_955,In_304,In_1462);
nor U956 (N_956,In_521,In_24);
and U957 (N_957,In_1182,In_737);
nand U958 (N_958,In_587,In_467);
nor U959 (N_959,In_1412,In_914);
or U960 (N_960,In_1093,In_367);
and U961 (N_961,In_501,In_1283);
nand U962 (N_962,In_463,In_433);
and U963 (N_963,In_318,In_1244);
nand U964 (N_964,In_1150,In_49);
nand U965 (N_965,In_889,In_382);
and U966 (N_966,In_649,In_561);
nor U967 (N_967,In_1452,In_1021);
and U968 (N_968,In_1163,In_1365);
and U969 (N_969,In_829,In_1187);
and U970 (N_970,In_54,In_1441);
nor U971 (N_971,In_879,In_357);
or U972 (N_972,In_428,In_11);
nor U973 (N_973,In_1291,In_632);
nor U974 (N_974,In_766,In_301);
nand U975 (N_975,In_474,In_118);
nand U976 (N_976,In_945,In_466);
or U977 (N_977,In_1247,In_475);
nor U978 (N_978,In_1181,In_1217);
xor U979 (N_979,In_996,In_826);
nor U980 (N_980,In_1182,In_273);
nor U981 (N_981,In_853,In_358);
nand U982 (N_982,In_642,In_1437);
or U983 (N_983,In_943,In_635);
nor U984 (N_984,In_879,In_1379);
or U985 (N_985,In_319,In_104);
or U986 (N_986,In_598,In_947);
or U987 (N_987,In_948,In_1393);
nor U988 (N_988,In_273,In_1152);
nor U989 (N_989,In_1104,In_1274);
nand U990 (N_990,In_704,In_1497);
and U991 (N_991,In_1001,In_513);
and U992 (N_992,In_1416,In_1181);
or U993 (N_993,In_7,In_1228);
nor U994 (N_994,In_428,In_1138);
nor U995 (N_995,In_1013,In_1159);
nor U996 (N_996,In_1170,In_753);
nand U997 (N_997,In_725,In_1142);
or U998 (N_998,In_508,In_697);
or U999 (N_999,In_175,In_153);
nor U1000 (N_1000,In_669,In_831);
and U1001 (N_1001,In_618,In_748);
nor U1002 (N_1002,In_423,In_721);
nand U1003 (N_1003,In_141,In_410);
and U1004 (N_1004,In_162,In_810);
or U1005 (N_1005,In_430,In_471);
nor U1006 (N_1006,In_990,In_473);
nand U1007 (N_1007,In_1441,In_699);
xor U1008 (N_1008,In_780,In_906);
nand U1009 (N_1009,In_416,In_1349);
or U1010 (N_1010,In_246,In_811);
and U1011 (N_1011,In_1396,In_1250);
xnor U1012 (N_1012,In_657,In_1419);
or U1013 (N_1013,In_668,In_859);
or U1014 (N_1014,In_418,In_772);
or U1015 (N_1015,In_478,In_1096);
or U1016 (N_1016,In_71,In_358);
nand U1017 (N_1017,In_912,In_737);
nand U1018 (N_1018,In_259,In_1275);
xnor U1019 (N_1019,In_1075,In_338);
and U1020 (N_1020,In_49,In_1403);
nor U1021 (N_1021,In_1194,In_35);
and U1022 (N_1022,In_761,In_330);
nor U1023 (N_1023,In_1063,In_1047);
and U1024 (N_1024,In_108,In_1080);
xnor U1025 (N_1025,In_277,In_1481);
and U1026 (N_1026,In_1308,In_355);
xor U1027 (N_1027,In_0,In_645);
nor U1028 (N_1028,In_317,In_599);
and U1029 (N_1029,In_320,In_664);
nor U1030 (N_1030,In_259,In_582);
or U1031 (N_1031,In_938,In_508);
and U1032 (N_1032,In_774,In_1428);
and U1033 (N_1033,In_481,In_1257);
nor U1034 (N_1034,In_799,In_942);
xnor U1035 (N_1035,In_1019,In_440);
nor U1036 (N_1036,In_776,In_833);
and U1037 (N_1037,In_978,In_1134);
or U1038 (N_1038,In_958,In_1126);
nand U1039 (N_1039,In_197,In_1286);
nor U1040 (N_1040,In_804,In_1185);
nor U1041 (N_1041,In_1313,In_590);
and U1042 (N_1042,In_267,In_526);
and U1043 (N_1043,In_948,In_959);
or U1044 (N_1044,In_1346,In_1465);
and U1045 (N_1045,In_1207,In_1292);
and U1046 (N_1046,In_934,In_1060);
nor U1047 (N_1047,In_635,In_332);
nor U1048 (N_1048,In_499,In_836);
and U1049 (N_1049,In_1382,In_1048);
nor U1050 (N_1050,In_1150,In_955);
and U1051 (N_1051,In_624,In_148);
and U1052 (N_1052,In_775,In_680);
or U1053 (N_1053,In_845,In_824);
or U1054 (N_1054,In_1045,In_1395);
nand U1055 (N_1055,In_1136,In_956);
or U1056 (N_1056,In_850,In_148);
nand U1057 (N_1057,In_1389,In_796);
nand U1058 (N_1058,In_1187,In_972);
and U1059 (N_1059,In_202,In_1401);
nand U1060 (N_1060,In_579,In_585);
nand U1061 (N_1061,In_1310,In_890);
and U1062 (N_1062,In_19,In_951);
nor U1063 (N_1063,In_221,In_756);
nand U1064 (N_1064,In_1437,In_1046);
or U1065 (N_1065,In_984,In_540);
nor U1066 (N_1066,In_865,In_873);
or U1067 (N_1067,In_1324,In_221);
or U1068 (N_1068,In_1491,In_852);
nand U1069 (N_1069,In_442,In_796);
nand U1070 (N_1070,In_440,In_570);
xnor U1071 (N_1071,In_1274,In_1115);
nor U1072 (N_1072,In_793,In_612);
xor U1073 (N_1073,In_1300,In_413);
and U1074 (N_1074,In_16,In_1392);
nand U1075 (N_1075,In_873,In_891);
or U1076 (N_1076,In_119,In_454);
and U1077 (N_1077,In_94,In_1324);
nor U1078 (N_1078,In_1127,In_118);
or U1079 (N_1079,In_941,In_1029);
or U1080 (N_1080,In_1275,In_208);
nand U1081 (N_1081,In_632,In_1422);
nor U1082 (N_1082,In_1277,In_1496);
or U1083 (N_1083,In_1312,In_922);
and U1084 (N_1084,In_989,In_9);
nand U1085 (N_1085,In_1371,In_1399);
and U1086 (N_1086,In_457,In_1497);
and U1087 (N_1087,In_250,In_998);
or U1088 (N_1088,In_1425,In_925);
nand U1089 (N_1089,In_1254,In_804);
xnor U1090 (N_1090,In_342,In_516);
and U1091 (N_1091,In_779,In_229);
and U1092 (N_1092,In_1383,In_86);
and U1093 (N_1093,In_289,In_465);
or U1094 (N_1094,In_481,In_99);
nand U1095 (N_1095,In_1154,In_1487);
and U1096 (N_1096,In_1142,In_1129);
xor U1097 (N_1097,In_1017,In_1225);
nand U1098 (N_1098,In_851,In_1448);
nand U1099 (N_1099,In_1048,In_1150);
or U1100 (N_1100,In_594,In_1148);
xnor U1101 (N_1101,In_1106,In_1349);
and U1102 (N_1102,In_819,In_143);
and U1103 (N_1103,In_624,In_1401);
or U1104 (N_1104,In_213,In_1027);
and U1105 (N_1105,In_383,In_1063);
nor U1106 (N_1106,In_1040,In_1383);
or U1107 (N_1107,In_360,In_589);
or U1108 (N_1108,In_228,In_1253);
or U1109 (N_1109,In_224,In_488);
nor U1110 (N_1110,In_838,In_1302);
nor U1111 (N_1111,In_1275,In_1490);
or U1112 (N_1112,In_1424,In_519);
and U1113 (N_1113,In_2,In_392);
nor U1114 (N_1114,In_606,In_100);
and U1115 (N_1115,In_1359,In_61);
nand U1116 (N_1116,In_1075,In_115);
nand U1117 (N_1117,In_444,In_909);
and U1118 (N_1118,In_1226,In_157);
nand U1119 (N_1119,In_802,In_243);
and U1120 (N_1120,In_960,In_314);
and U1121 (N_1121,In_62,In_168);
and U1122 (N_1122,In_1018,In_871);
nor U1123 (N_1123,In_1327,In_1231);
and U1124 (N_1124,In_726,In_249);
and U1125 (N_1125,In_1116,In_710);
nand U1126 (N_1126,In_1439,In_80);
nand U1127 (N_1127,In_939,In_839);
nor U1128 (N_1128,In_873,In_541);
nor U1129 (N_1129,In_760,In_1319);
and U1130 (N_1130,In_731,In_863);
or U1131 (N_1131,In_1356,In_500);
or U1132 (N_1132,In_81,In_365);
or U1133 (N_1133,In_760,In_523);
nor U1134 (N_1134,In_1065,In_231);
nand U1135 (N_1135,In_847,In_1408);
or U1136 (N_1136,In_1322,In_705);
nor U1137 (N_1137,In_1229,In_295);
and U1138 (N_1138,In_96,In_1483);
xnor U1139 (N_1139,In_1110,In_731);
and U1140 (N_1140,In_1423,In_972);
and U1141 (N_1141,In_828,In_520);
or U1142 (N_1142,In_118,In_1439);
nand U1143 (N_1143,In_194,In_1482);
nand U1144 (N_1144,In_559,In_197);
nand U1145 (N_1145,In_463,In_1315);
nor U1146 (N_1146,In_92,In_525);
and U1147 (N_1147,In_632,In_519);
and U1148 (N_1148,In_885,In_721);
nor U1149 (N_1149,In_938,In_832);
or U1150 (N_1150,In_1464,In_796);
or U1151 (N_1151,In_1398,In_54);
xnor U1152 (N_1152,In_364,In_628);
nand U1153 (N_1153,In_925,In_1363);
nand U1154 (N_1154,In_1058,In_815);
xor U1155 (N_1155,In_532,In_272);
xnor U1156 (N_1156,In_1487,In_475);
and U1157 (N_1157,In_391,In_302);
or U1158 (N_1158,In_240,In_56);
and U1159 (N_1159,In_634,In_538);
or U1160 (N_1160,In_607,In_792);
nor U1161 (N_1161,In_1125,In_180);
nor U1162 (N_1162,In_622,In_780);
nor U1163 (N_1163,In_873,In_737);
or U1164 (N_1164,In_511,In_1276);
and U1165 (N_1165,In_293,In_285);
nor U1166 (N_1166,In_792,In_1463);
and U1167 (N_1167,In_837,In_1488);
xnor U1168 (N_1168,In_167,In_272);
xor U1169 (N_1169,In_904,In_168);
xor U1170 (N_1170,In_861,In_1070);
and U1171 (N_1171,In_55,In_433);
nor U1172 (N_1172,In_62,In_1061);
nand U1173 (N_1173,In_257,In_631);
nand U1174 (N_1174,In_472,In_475);
nand U1175 (N_1175,In_1273,In_162);
nor U1176 (N_1176,In_438,In_726);
xnor U1177 (N_1177,In_1285,In_601);
nor U1178 (N_1178,In_466,In_562);
nand U1179 (N_1179,In_761,In_1413);
nor U1180 (N_1180,In_232,In_553);
and U1181 (N_1181,In_1166,In_889);
nor U1182 (N_1182,In_270,In_1168);
or U1183 (N_1183,In_12,In_267);
or U1184 (N_1184,In_744,In_1248);
nor U1185 (N_1185,In_591,In_1127);
nand U1186 (N_1186,In_1355,In_768);
xor U1187 (N_1187,In_128,In_515);
nand U1188 (N_1188,In_1067,In_1145);
and U1189 (N_1189,In_1492,In_424);
nand U1190 (N_1190,In_1396,In_629);
or U1191 (N_1191,In_1027,In_338);
and U1192 (N_1192,In_40,In_732);
and U1193 (N_1193,In_566,In_1353);
xor U1194 (N_1194,In_194,In_1456);
or U1195 (N_1195,In_512,In_659);
and U1196 (N_1196,In_388,In_681);
and U1197 (N_1197,In_455,In_1151);
nor U1198 (N_1198,In_806,In_631);
nor U1199 (N_1199,In_1083,In_957);
nand U1200 (N_1200,In_932,In_287);
nand U1201 (N_1201,In_269,In_819);
or U1202 (N_1202,In_458,In_83);
and U1203 (N_1203,In_638,In_288);
nor U1204 (N_1204,In_1476,In_914);
nand U1205 (N_1205,In_1045,In_927);
nand U1206 (N_1206,In_743,In_423);
and U1207 (N_1207,In_983,In_1464);
xor U1208 (N_1208,In_641,In_374);
nor U1209 (N_1209,In_523,In_416);
nor U1210 (N_1210,In_654,In_640);
and U1211 (N_1211,In_849,In_778);
nor U1212 (N_1212,In_939,In_1109);
and U1213 (N_1213,In_317,In_541);
nor U1214 (N_1214,In_1146,In_966);
nand U1215 (N_1215,In_23,In_1331);
nand U1216 (N_1216,In_131,In_1404);
nand U1217 (N_1217,In_662,In_1477);
or U1218 (N_1218,In_590,In_1075);
or U1219 (N_1219,In_556,In_1088);
nor U1220 (N_1220,In_502,In_660);
and U1221 (N_1221,In_1017,In_1278);
nand U1222 (N_1222,In_1269,In_1313);
nand U1223 (N_1223,In_13,In_831);
or U1224 (N_1224,In_55,In_788);
or U1225 (N_1225,In_32,In_453);
nand U1226 (N_1226,In_69,In_1070);
nand U1227 (N_1227,In_472,In_30);
nand U1228 (N_1228,In_690,In_1491);
nand U1229 (N_1229,In_750,In_24);
and U1230 (N_1230,In_681,In_1233);
nor U1231 (N_1231,In_57,In_289);
nor U1232 (N_1232,In_676,In_27);
nor U1233 (N_1233,In_16,In_392);
nand U1234 (N_1234,In_313,In_1051);
nor U1235 (N_1235,In_762,In_1059);
nand U1236 (N_1236,In_1207,In_0);
and U1237 (N_1237,In_1441,In_515);
xor U1238 (N_1238,In_639,In_107);
nand U1239 (N_1239,In_485,In_609);
or U1240 (N_1240,In_628,In_875);
or U1241 (N_1241,In_1368,In_499);
xor U1242 (N_1242,In_223,In_974);
and U1243 (N_1243,In_924,In_964);
nor U1244 (N_1244,In_40,In_70);
or U1245 (N_1245,In_1184,In_38);
nand U1246 (N_1246,In_149,In_1198);
or U1247 (N_1247,In_485,In_153);
and U1248 (N_1248,In_629,In_178);
and U1249 (N_1249,In_426,In_947);
nand U1250 (N_1250,In_349,In_137);
nor U1251 (N_1251,In_1182,In_1350);
xor U1252 (N_1252,In_548,In_1123);
or U1253 (N_1253,In_1406,In_1203);
and U1254 (N_1254,In_40,In_1129);
nand U1255 (N_1255,In_49,In_1378);
or U1256 (N_1256,In_712,In_970);
nand U1257 (N_1257,In_206,In_702);
nand U1258 (N_1258,In_660,In_640);
nand U1259 (N_1259,In_79,In_530);
or U1260 (N_1260,In_952,In_135);
or U1261 (N_1261,In_174,In_548);
nor U1262 (N_1262,In_457,In_79);
xnor U1263 (N_1263,In_470,In_906);
nor U1264 (N_1264,In_378,In_982);
or U1265 (N_1265,In_1443,In_361);
or U1266 (N_1266,In_888,In_319);
nor U1267 (N_1267,In_209,In_1244);
nor U1268 (N_1268,In_89,In_1167);
and U1269 (N_1269,In_1444,In_1351);
or U1270 (N_1270,In_724,In_168);
and U1271 (N_1271,In_442,In_1247);
nand U1272 (N_1272,In_354,In_463);
nor U1273 (N_1273,In_1018,In_903);
and U1274 (N_1274,In_543,In_1035);
and U1275 (N_1275,In_1418,In_568);
xnor U1276 (N_1276,In_691,In_1324);
or U1277 (N_1277,In_1402,In_1031);
or U1278 (N_1278,In_1437,In_951);
xnor U1279 (N_1279,In_65,In_956);
xor U1280 (N_1280,In_787,In_625);
nor U1281 (N_1281,In_279,In_474);
and U1282 (N_1282,In_423,In_1094);
and U1283 (N_1283,In_1240,In_283);
nor U1284 (N_1284,In_68,In_471);
nor U1285 (N_1285,In_39,In_1231);
xnor U1286 (N_1286,In_300,In_1103);
nor U1287 (N_1287,In_855,In_31);
and U1288 (N_1288,In_727,In_1141);
and U1289 (N_1289,In_448,In_1197);
nor U1290 (N_1290,In_500,In_1025);
or U1291 (N_1291,In_1135,In_152);
nor U1292 (N_1292,In_267,In_1279);
or U1293 (N_1293,In_479,In_933);
or U1294 (N_1294,In_73,In_1208);
nor U1295 (N_1295,In_270,In_575);
nor U1296 (N_1296,In_1080,In_678);
and U1297 (N_1297,In_793,In_819);
xnor U1298 (N_1298,In_1133,In_993);
nor U1299 (N_1299,In_148,In_326);
nand U1300 (N_1300,In_449,In_21);
nand U1301 (N_1301,In_1313,In_1381);
nor U1302 (N_1302,In_203,In_781);
nor U1303 (N_1303,In_483,In_227);
nor U1304 (N_1304,In_949,In_553);
nor U1305 (N_1305,In_1099,In_478);
or U1306 (N_1306,In_1081,In_959);
and U1307 (N_1307,In_1362,In_673);
and U1308 (N_1308,In_744,In_1168);
or U1309 (N_1309,In_752,In_44);
nand U1310 (N_1310,In_1163,In_350);
nand U1311 (N_1311,In_1260,In_743);
nor U1312 (N_1312,In_1354,In_1224);
nor U1313 (N_1313,In_1305,In_1005);
nor U1314 (N_1314,In_1272,In_256);
nand U1315 (N_1315,In_1214,In_1229);
and U1316 (N_1316,In_681,In_812);
nand U1317 (N_1317,In_75,In_349);
and U1318 (N_1318,In_1361,In_1483);
xor U1319 (N_1319,In_248,In_240);
and U1320 (N_1320,In_1326,In_1293);
and U1321 (N_1321,In_1204,In_1160);
nand U1322 (N_1322,In_62,In_980);
nand U1323 (N_1323,In_483,In_1469);
and U1324 (N_1324,In_831,In_1265);
nand U1325 (N_1325,In_32,In_1176);
or U1326 (N_1326,In_212,In_1239);
nor U1327 (N_1327,In_1421,In_138);
xnor U1328 (N_1328,In_886,In_986);
and U1329 (N_1329,In_483,In_137);
nand U1330 (N_1330,In_534,In_1418);
nand U1331 (N_1331,In_271,In_771);
nand U1332 (N_1332,In_263,In_1024);
nand U1333 (N_1333,In_1247,In_509);
nor U1334 (N_1334,In_1268,In_733);
and U1335 (N_1335,In_510,In_103);
and U1336 (N_1336,In_606,In_249);
nand U1337 (N_1337,In_660,In_1152);
or U1338 (N_1338,In_1132,In_872);
or U1339 (N_1339,In_705,In_1089);
nor U1340 (N_1340,In_502,In_1008);
nor U1341 (N_1341,In_887,In_763);
and U1342 (N_1342,In_390,In_388);
nor U1343 (N_1343,In_769,In_302);
and U1344 (N_1344,In_318,In_1235);
nand U1345 (N_1345,In_418,In_1360);
and U1346 (N_1346,In_1207,In_716);
xnor U1347 (N_1347,In_264,In_124);
or U1348 (N_1348,In_1384,In_145);
or U1349 (N_1349,In_164,In_1333);
nor U1350 (N_1350,In_427,In_406);
and U1351 (N_1351,In_268,In_416);
nand U1352 (N_1352,In_1069,In_1097);
and U1353 (N_1353,In_1479,In_460);
and U1354 (N_1354,In_1113,In_1090);
and U1355 (N_1355,In_728,In_563);
and U1356 (N_1356,In_1154,In_49);
nand U1357 (N_1357,In_1309,In_803);
or U1358 (N_1358,In_1458,In_914);
nor U1359 (N_1359,In_688,In_1107);
nor U1360 (N_1360,In_1293,In_1105);
nor U1361 (N_1361,In_1459,In_514);
nand U1362 (N_1362,In_1032,In_1061);
nor U1363 (N_1363,In_1162,In_345);
or U1364 (N_1364,In_143,In_433);
nand U1365 (N_1365,In_1282,In_1365);
or U1366 (N_1366,In_1008,In_252);
xnor U1367 (N_1367,In_27,In_488);
nor U1368 (N_1368,In_916,In_695);
nor U1369 (N_1369,In_859,In_1240);
or U1370 (N_1370,In_60,In_253);
nor U1371 (N_1371,In_153,In_499);
and U1372 (N_1372,In_1347,In_687);
or U1373 (N_1373,In_465,In_1167);
or U1374 (N_1374,In_476,In_222);
or U1375 (N_1375,In_819,In_679);
and U1376 (N_1376,In_76,In_727);
or U1377 (N_1377,In_1141,In_1336);
xnor U1378 (N_1378,In_365,In_1417);
and U1379 (N_1379,In_1162,In_36);
nor U1380 (N_1380,In_879,In_1449);
and U1381 (N_1381,In_342,In_1230);
or U1382 (N_1382,In_400,In_531);
xor U1383 (N_1383,In_40,In_578);
xor U1384 (N_1384,In_1079,In_956);
nand U1385 (N_1385,In_507,In_132);
xnor U1386 (N_1386,In_1364,In_1080);
xnor U1387 (N_1387,In_1197,In_389);
or U1388 (N_1388,In_719,In_255);
and U1389 (N_1389,In_526,In_20);
nor U1390 (N_1390,In_905,In_1119);
and U1391 (N_1391,In_266,In_642);
or U1392 (N_1392,In_242,In_783);
nor U1393 (N_1393,In_1208,In_1035);
nor U1394 (N_1394,In_1235,In_181);
nor U1395 (N_1395,In_575,In_58);
or U1396 (N_1396,In_512,In_162);
or U1397 (N_1397,In_112,In_530);
nor U1398 (N_1398,In_106,In_608);
and U1399 (N_1399,In_1384,In_888);
nand U1400 (N_1400,In_501,In_704);
or U1401 (N_1401,In_80,In_354);
nor U1402 (N_1402,In_403,In_1046);
and U1403 (N_1403,In_180,In_1421);
and U1404 (N_1404,In_597,In_1129);
or U1405 (N_1405,In_351,In_477);
or U1406 (N_1406,In_991,In_448);
nor U1407 (N_1407,In_769,In_568);
nand U1408 (N_1408,In_747,In_1003);
nand U1409 (N_1409,In_1229,In_12);
xnor U1410 (N_1410,In_750,In_74);
or U1411 (N_1411,In_24,In_269);
nand U1412 (N_1412,In_1112,In_673);
or U1413 (N_1413,In_350,In_639);
or U1414 (N_1414,In_787,In_1244);
and U1415 (N_1415,In_310,In_382);
nand U1416 (N_1416,In_1402,In_285);
nor U1417 (N_1417,In_1214,In_138);
or U1418 (N_1418,In_664,In_598);
nand U1419 (N_1419,In_1443,In_228);
and U1420 (N_1420,In_187,In_790);
nand U1421 (N_1421,In_345,In_597);
nor U1422 (N_1422,In_124,In_537);
nand U1423 (N_1423,In_916,In_349);
and U1424 (N_1424,In_316,In_476);
or U1425 (N_1425,In_502,In_437);
and U1426 (N_1426,In_990,In_499);
or U1427 (N_1427,In_926,In_227);
nand U1428 (N_1428,In_1296,In_520);
nor U1429 (N_1429,In_344,In_264);
nand U1430 (N_1430,In_180,In_224);
and U1431 (N_1431,In_142,In_435);
and U1432 (N_1432,In_528,In_483);
and U1433 (N_1433,In_1000,In_979);
or U1434 (N_1434,In_19,In_431);
or U1435 (N_1435,In_166,In_1408);
nor U1436 (N_1436,In_836,In_823);
nor U1437 (N_1437,In_1497,In_817);
and U1438 (N_1438,In_1255,In_701);
or U1439 (N_1439,In_1283,In_435);
or U1440 (N_1440,In_1083,In_71);
nand U1441 (N_1441,In_1384,In_882);
xor U1442 (N_1442,In_756,In_326);
nor U1443 (N_1443,In_1346,In_85);
and U1444 (N_1444,In_908,In_234);
xnor U1445 (N_1445,In_783,In_447);
nand U1446 (N_1446,In_494,In_595);
and U1447 (N_1447,In_848,In_466);
nor U1448 (N_1448,In_622,In_1121);
or U1449 (N_1449,In_1224,In_774);
nand U1450 (N_1450,In_15,In_169);
or U1451 (N_1451,In_1363,In_903);
or U1452 (N_1452,In_246,In_1444);
nor U1453 (N_1453,In_72,In_865);
or U1454 (N_1454,In_625,In_63);
nand U1455 (N_1455,In_1085,In_1089);
xnor U1456 (N_1456,In_1045,In_377);
and U1457 (N_1457,In_594,In_1005);
nand U1458 (N_1458,In_484,In_593);
or U1459 (N_1459,In_398,In_1338);
nor U1460 (N_1460,In_1225,In_1162);
xor U1461 (N_1461,In_167,In_1306);
nand U1462 (N_1462,In_625,In_890);
and U1463 (N_1463,In_545,In_1412);
nand U1464 (N_1464,In_400,In_148);
xnor U1465 (N_1465,In_404,In_393);
nor U1466 (N_1466,In_386,In_842);
xor U1467 (N_1467,In_1000,In_1469);
nand U1468 (N_1468,In_205,In_834);
or U1469 (N_1469,In_6,In_253);
and U1470 (N_1470,In_670,In_1315);
nand U1471 (N_1471,In_317,In_338);
nor U1472 (N_1472,In_827,In_973);
nand U1473 (N_1473,In_947,In_908);
nand U1474 (N_1474,In_847,In_915);
nand U1475 (N_1475,In_1056,In_30);
nand U1476 (N_1476,In_1182,In_910);
and U1477 (N_1477,In_72,In_1021);
nor U1478 (N_1478,In_332,In_341);
and U1479 (N_1479,In_197,In_1373);
nor U1480 (N_1480,In_101,In_1448);
and U1481 (N_1481,In_1041,In_296);
or U1482 (N_1482,In_642,In_350);
nor U1483 (N_1483,In_1317,In_717);
nand U1484 (N_1484,In_983,In_239);
or U1485 (N_1485,In_64,In_75);
or U1486 (N_1486,In_254,In_1456);
nand U1487 (N_1487,In_67,In_1221);
or U1488 (N_1488,In_443,In_385);
and U1489 (N_1489,In_1370,In_70);
xnor U1490 (N_1490,In_1112,In_248);
and U1491 (N_1491,In_288,In_1137);
and U1492 (N_1492,In_592,In_1330);
nor U1493 (N_1493,In_1392,In_239);
or U1494 (N_1494,In_1034,In_26);
or U1495 (N_1495,In_1216,In_1415);
nor U1496 (N_1496,In_1070,In_255);
nor U1497 (N_1497,In_869,In_527);
nand U1498 (N_1498,In_1212,In_686);
and U1499 (N_1499,In_117,In_845);
nand U1500 (N_1500,In_553,In_929);
nor U1501 (N_1501,In_1248,In_655);
or U1502 (N_1502,In_1336,In_29);
or U1503 (N_1503,In_949,In_230);
nor U1504 (N_1504,In_606,In_1306);
nand U1505 (N_1505,In_794,In_1281);
and U1506 (N_1506,In_13,In_217);
xnor U1507 (N_1507,In_468,In_105);
nor U1508 (N_1508,In_906,In_1477);
or U1509 (N_1509,In_1387,In_90);
nand U1510 (N_1510,In_784,In_1263);
nor U1511 (N_1511,In_778,In_795);
and U1512 (N_1512,In_734,In_1401);
nor U1513 (N_1513,In_919,In_1263);
and U1514 (N_1514,In_1075,In_1217);
or U1515 (N_1515,In_181,In_917);
nor U1516 (N_1516,In_210,In_155);
and U1517 (N_1517,In_1287,In_533);
nor U1518 (N_1518,In_650,In_1068);
nor U1519 (N_1519,In_1464,In_638);
xor U1520 (N_1520,In_819,In_645);
xor U1521 (N_1521,In_666,In_471);
xor U1522 (N_1522,In_655,In_328);
nor U1523 (N_1523,In_867,In_231);
and U1524 (N_1524,In_300,In_3);
or U1525 (N_1525,In_364,In_1010);
xnor U1526 (N_1526,In_1297,In_595);
nor U1527 (N_1527,In_1116,In_1330);
or U1528 (N_1528,In_1231,In_830);
nor U1529 (N_1529,In_166,In_836);
or U1530 (N_1530,In_1299,In_61);
xor U1531 (N_1531,In_517,In_268);
and U1532 (N_1532,In_1076,In_135);
and U1533 (N_1533,In_216,In_831);
or U1534 (N_1534,In_1342,In_644);
and U1535 (N_1535,In_936,In_923);
and U1536 (N_1536,In_785,In_960);
xor U1537 (N_1537,In_196,In_949);
or U1538 (N_1538,In_952,In_1446);
or U1539 (N_1539,In_315,In_296);
or U1540 (N_1540,In_662,In_152);
nand U1541 (N_1541,In_29,In_368);
nand U1542 (N_1542,In_959,In_826);
nor U1543 (N_1543,In_1253,In_1125);
and U1544 (N_1544,In_1260,In_250);
and U1545 (N_1545,In_552,In_953);
nand U1546 (N_1546,In_684,In_1177);
and U1547 (N_1547,In_1025,In_505);
nor U1548 (N_1548,In_167,In_942);
nor U1549 (N_1549,In_759,In_329);
nand U1550 (N_1550,In_1126,In_578);
nand U1551 (N_1551,In_154,In_914);
and U1552 (N_1552,In_354,In_1041);
nand U1553 (N_1553,In_600,In_341);
nand U1554 (N_1554,In_522,In_981);
or U1555 (N_1555,In_943,In_631);
nand U1556 (N_1556,In_357,In_900);
and U1557 (N_1557,In_21,In_1494);
nand U1558 (N_1558,In_724,In_273);
or U1559 (N_1559,In_972,In_507);
and U1560 (N_1560,In_532,In_140);
and U1561 (N_1561,In_453,In_537);
and U1562 (N_1562,In_1356,In_506);
nand U1563 (N_1563,In_1371,In_541);
and U1564 (N_1564,In_881,In_1364);
nor U1565 (N_1565,In_1434,In_309);
or U1566 (N_1566,In_770,In_26);
or U1567 (N_1567,In_1007,In_61);
or U1568 (N_1568,In_424,In_543);
nor U1569 (N_1569,In_1162,In_1332);
nor U1570 (N_1570,In_18,In_185);
nor U1571 (N_1571,In_668,In_630);
or U1572 (N_1572,In_947,In_282);
and U1573 (N_1573,In_1251,In_1285);
nor U1574 (N_1574,In_445,In_457);
or U1575 (N_1575,In_1120,In_1197);
or U1576 (N_1576,In_146,In_1297);
and U1577 (N_1577,In_730,In_885);
nand U1578 (N_1578,In_1129,In_516);
xor U1579 (N_1579,In_620,In_351);
or U1580 (N_1580,In_90,In_1038);
xnor U1581 (N_1581,In_576,In_612);
nand U1582 (N_1582,In_887,In_96);
xor U1583 (N_1583,In_475,In_194);
or U1584 (N_1584,In_671,In_877);
and U1585 (N_1585,In_1278,In_1465);
or U1586 (N_1586,In_1253,In_317);
or U1587 (N_1587,In_1478,In_1150);
xor U1588 (N_1588,In_998,In_928);
nor U1589 (N_1589,In_865,In_1435);
nand U1590 (N_1590,In_266,In_747);
nand U1591 (N_1591,In_921,In_32);
or U1592 (N_1592,In_249,In_1375);
nand U1593 (N_1593,In_667,In_1239);
nor U1594 (N_1594,In_1397,In_1348);
nand U1595 (N_1595,In_1145,In_1350);
and U1596 (N_1596,In_478,In_379);
and U1597 (N_1597,In_500,In_951);
and U1598 (N_1598,In_860,In_1471);
or U1599 (N_1599,In_1224,In_1088);
xor U1600 (N_1600,In_827,In_296);
nor U1601 (N_1601,In_133,In_372);
and U1602 (N_1602,In_967,In_1329);
nand U1603 (N_1603,In_76,In_443);
and U1604 (N_1604,In_1465,In_569);
nand U1605 (N_1605,In_1192,In_1486);
nor U1606 (N_1606,In_1327,In_216);
nor U1607 (N_1607,In_1355,In_457);
nor U1608 (N_1608,In_1449,In_1218);
nand U1609 (N_1609,In_804,In_889);
or U1610 (N_1610,In_928,In_1059);
or U1611 (N_1611,In_95,In_914);
or U1612 (N_1612,In_224,In_107);
or U1613 (N_1613,In_436,In_101);
or U1614 (N_1614,In_752,In_1398);
xnor U1615 (N_1615,In_522,In_221);
xnor U1616 (N_1616,In_1290,In_1350);
xnor U1617 (N_1617,In_19,In_459);
or U1618 (N_1618,In_182,In_629);
or U1619 (N_1619,In_1191,In_1351);
nor U1620 (N_1620,In_12,In_1198);
nand U1621 (N_1621,In_1180,In_740);
and U1622 (N_1622,In_1286,In_750);
nor U1623 (N_1623,In_642,In_519);
and U1624 (N_1624,In_167,In_1439);
xor U1625 (N_1625,In_144,In_597);
or U1626 (N_1626,In_78,In_387);
or U1627 (N_1627,In_869,In_823);
nor U1628 (N_1628,In_702,In_981);
and U1629 (N_1629,In_50,In_747);
or U1630 (N_1630,In_743,In_576);
nand U1631 (N_1631,In_784,In_96);
nand U1632 (N_1632,In_509,In_1315);
and U1633 (N_1633,In_667,In_607);
nor U1634 (N_1634,In_1428,In_136);
nand U1635 (N_1635,In_349,In_834);
xnor U1636 (N_1636,In_1498,In_1145);
nor U1637 (N_1637,In_1392,In_1223);
and U1638 (N_1638,In_313,In_635);
xnor U1639 (N_1639,In_238,In_891);
nor U1640 (N_1640,In_942,In_1442);
or U1641 (N_1641,In_434,In_1322);
and U1642 (N_1642,In_1036,In_420);
or U1643 (N_1643,In_999,In_1189);
and U1644 (N_1644,In_141,In_941);
nor U1645 (N_1645,In_5,In_837);
or U1646 (N_1646,In_1066,In_376);
and U1647 (N_1647,In_467,In_63);
nand U1648 (N_1648,In_688,In_110);
and U1649 (N_1649,In_1453,In_612);
and U1650 (N_1650,In_3,In_1196);
xnor U1651 (N_1651,In_471,In_362);
or U1652 (N_1652,In_1108,In_1227);
nor U1653 (N_1653,In_1026,In_599);
nand U1654 (N_1654,In_553,In_431);
or U1655 (N_1655,In_14,In_322);
and U1656 (N_1656,In_184,In_73);
and U1657 (N_1657,In_1075,In_881);
and U1658 (N_1658,In_343,In_770);
or U1659 (N_1659,In_3,In_906);
nand U1660 (N_1660,In_961,In_1264);
and U1661 (N_1661,In_1153,In_283);
xnor U1662 (N_1662,In_1441,In_502);
and U1663 (N_1663,In_845,In_420);
and U1664 (N_1664,In_419,In_688);
or U1665 (N_1665,In_1147,In_32);
nand U1666 (N_1666,In_1238,In_1425);
nor U1667 (N_1667,In_141,In_475);
nor U1668 (N_1668,In_729,In_1060);
or U1669 (N_1669,In_421,In_1171);
and U1670 (N_1670,In_319,In_91);
nor U1671 (N_1671,In_389,In_733);
or U1672 (N_1672,In_1299,In_818);
nor U1673 (N_1673,In_97,In_1446);
nor U1674 (N_1674,In_914,In_1254);
nand U1675 (N_1675,In_271,In_567);
or U1676 (N_1676,In_930,In_594);
nand U1677 (N_1677,In_807,In_1338);
and U1678 (N_1678,In_1159,In_1313);
nand U1679 (N_1679,In_36,In_119);
nor U1680 (N_1680,In_986,In_1253);
nand U1681 (N_1681,In_1349,In_1149);
and U1682 (N_1682,In_163,In_436);
and U1683 (N_1683,In_227,In_567);
and U1684 (N_1684,In_1042,In_806);
or U1685 (N_1685,In_786,In_1229);
or U1686 (N_1686,In_352,In_165);
xnor U1687 (N_1687,In_1290,In_1264);
nor U1688 (N_1688,In_1029,In_442);
xor U1689 (N_1689,In_675,In_937);
xor U1690 (N_1690,In_699,In_1348);
and U1691 (N_1691,In_1359,In_1196);
nand U1692 (N_1692,In_1299,In_995);
or U1693 (N_1693,In_295,In_50);
nand U1694 (N_1694,In_1284,In_1340);
xnor U1695 (N_1695,In_275,In_300);
nand U1696 (N_1696,In_649,In_470);
xor U1697 (N_1697,In_1382,In_966);
and U1698 (N_1698,In_977,In_636);
or U1699 (N_1699,In_1449,In_1153);
nor U1700 (N_1700,In_1138,In_1337);
nor U1701 (N_1701,In_22,In_227);
nor U1702 (N_1702,In_948,In_763);
or U1703 (N_1703,In_993,In_669);
and U1704 (N_1704,In_434,In_1121);
nand U1705 (N_1705,In_1338,In_422);
or U1706 (N_1706,In_1180,In_240);
and U1707 (N_1707,In_512,In_1415);
nor U1708 (N_1708,In_153,In_1210);
or U1709 (N_1709,In_266,In_75);
xor U1710 (N_1710,In_1129,In_936);
nand U1711 (N_1711,In_977,In_1087);
xnor U1712 (N_1712,In_855,In_1284);
and U1713 (N_1713,In_222,In_1448);
nor U1714 (N_1714,In_1465,In_205);
or U1715 (N_1715,In_1109,In_852);
or U1716 (N_1716,In_201,In_1406);
and U1717 (N_1717,In_1420,In_185);
or U1718 (N_1718,In_119,In_444);
nand U1719 (N_1719,In_1368,In_410);
and U1720 (N_1720,In_556,In_1362);
nand U1721 (N_1721,In_1035,In_1013);
nor U1722 (N_1722,In_188,In_592);
nor U1723 (N_1723,In_652,In_1295);
and U1724 (N_1724,In_72,In_1131);
or U1725 (N_1725,In_1119,In_1430);
or U1726 (N_1726,In_727,In_1355);
or U1727 (N_1727,In_374,In_1075);
nor U1728 (N_1728,In_737,In_1458);
nand U1729 (N_1729,In_233,In_1148);
nand U1730 (N_1730,In_699,In_159);
nor U1731 (N_1731,In_96,In_82);
or U1732 (N_1732,In_1495,In_1424);
nand U1733 (N_1733,In_1494,In_488);
and U1734 (N_1734,In_1188,In_1343);
or U1735 (N_1735,In_1,In_1463);
nor U1736 (N_1736,In_480,In_291);
or U1737 (N_1737,In_98,In_458);
xor U1738 (N_1738,In_570,In_558);
or U1739 (N_1739,In_832,In_1367);
or U1740 (N_1740,In_368,In_476);
or U1741 (N_1741,In_1130,In_1047);
and U1742 (N_1742,In_917,In_609);
nor U1743 (N_1743,In_954,In_445);
and U1744 (N_1744,In_380,In_524);
and U1745 (N_1745,In_630,In_817);
nand U1746 (N_1746,In_189,In_314);
nand U1747 (N_1747,In_1016,In_1092);
or U1748 (N_1748,In_253,In_1255);
xnor U1749 (N_1749,In_725,In_314);
xor U1750 (N_1750,In_697,In_1142);
or U1751 (N_1751,In_1212,In_971);
and U1752 (N_1752,In_884,In_187);
nand U1753 (N_1753,In_430,In_694);
and U1754 (N_1754,In_171,In_744);
nand U1755 (N_1755,In_913,In_1483);
nor U1756 (N_1756,In_1458,In_729);
nor U1757 (N_1757,In_1042,In_1191);
and U1758 (N_1758,In_1116,In_1421);
and U1759 (N_1759,In_107,In_1005);
nor U1760 (N_1760,In_1095,In_950);
or U1761 (N_1761,In_518,In_1199);
and U1762 (N_1762,In_214,In_472);
nor U1763 (N_1763,In_1199,In_1221);
and U1764 (N_1764,In_732,In_848);
nor U1765 (N_1765,In_210,In_345);
or U1766 (N_1766,In_457,In_1207);
or U1767 (N_1767,In_807,In_427);
xor U1768 (N_1768,In_451,In_758);
or U1769 (N_1769,In_1121,In_932);
or U1770 (N_1770,In_1175,In_36);
nand U1771 (N_1771,In_1440,In_293);
nand U1772 (N_1772,In_1132,In_624);
nor U1773 (N_1773,In_521,In_937);
or U1774 (N_1774,In_27,In_682);
nand U1775 (N_1775,In_578,In_863);
and U1776 (N_1776,In_66,In_55);
nand U1777 (N_1777,In_1122,In_1411);
and U1778 (N_1778,In_109,In_119);
and U1779 (N_1779,In_146,In_1232);
and U1780 (N_1780,In_446,In_1076);
nor U1781 (N_1781,In_1243,In_266);
xnor U1782 (N_1782,In_744,In_1435);
xor U1783 (N_1783,In_1271,In_1417);
or U1784 (N_1784,In_857,In_1091);
nand U1785 (N_1785,In_1298,In_405);
or U1786 (N_1786,In_1283,In_408);
nor U1787 (N_1787,In_290,In_1048);
xor U1788 (N_1788,In_412,In_312);
xor U1789 (N_1789,In_252,In_830);
and U1790 (N_1790,In_1150,In_702);
nor U1791 (N_1791,In_620,In_1421);
or U1792 (N_1792,In_1408,In_701);
xnor U1793 (N_1793,In_1006,In_28);
nor U1794 (N_1794,In_980,In_349);
xnor U1795 (N_1795,In_878,In_872);
nor U1796 (N_1796,In_454,In_1098);
and U1797 (N_1797,In_890,In_299);
nand U1798 (N_1798,In_1292,In_833);
and U1799 (N_1799,In_1045,In_252);
nor U1800 (N_1800,In_1467,In_267);
and U1801 (N_1801,In_866,In_876);
xor U1802 (N_1802,In_699,In_1100);
xor U1803 (N_1803,In_1244,In_393);
xor U1804 (N_1804,In_766,In_24);
nand U1805 (N_1805,In_1246,In_1223);
xor U1806 (N_1806,In_663,In_399);
or U1807 (N_1807,In_1116,In_727);
nand U1808 (N_1808,In_798,In_1388);
or U1809 (N_1809,In_92,In_1181);
and U1810 (N_1810,In_191,In_33);
and U1811 (N_1811,In_927,In_562);
nand U1812 (N_1812,In_184,In_244);
nor U1813 (N_1813,In_499,In_563);
and U1814 (N_1814,In_1342,In_912);
xor U1815 (N_1815,In_515,In_411);
nor U1816 (N_1816,In_359,In_321);
xnor U1817 (N_1817,In_939,In_1323);
nor U1818 (N_1818,In_716,In_1278);
nor U1819 (N_1819,In_1468,In_1332);
or U1820 (N_1820,In_929,In_979);
nand U1821 (N_1821,In_339,In_399);
or U1822 (N_1822,In_851,In_1080);
nand U1823 (N_1823,In_855,In_973);
xnor U1824 (N_1824,In_1416,In_1203);
nand U1825 (N_1825,In_933,In_576);
or U1826 (N_1826,In_1305,In_1465);
nand U1827 (N_1827,In_161,In_1452);
and U1828 (N_1828,In_592,In_1239);
nand U1829 (N_1829,In_800,In_868);
or U1830 (N_1830,In_755,In_415);
nor U1831 (N_1831,In_1453,In_1256);
or U1832 (N_1832,In_774,In_826);
or U1833 (N_1833,In_325,In_1387);
and U1834 (N_1834,In_760,In_1195);
or U1835 (N_1835,In_153,In_908);
and U1836 (N_1836,In_1411,In_319);
and U1837 (N_1837,In_904,In_1153);
nand U1838 (N_1838,In_966,In_364);
nand U1839 (N_1839,In_1430,In_1467);
and U1840 (N_1840,In_1420,In_427);
or U1841 (N_1841,In_346,In_1119);
or U1842 (N_1842,In_396,In_340);
and U1843 (N_1843,In_1190,In_732);
xor U1844 (N_1844,In_1145,In_338);
nand U1845 (N_1845,In_882,In_946);
nor U1846 (N_1846,In_714,In_239);
nand U1847 (N_1847,In_727,In_709);
nor U1848 (N_1848,In_17,In_340);
xor U1849 (N_1849,In_300,In_683);
nor U1850 (N_1850,In_870,In_1287);
and U1851 (N_1851,In_796,In_650);
and U1852 (N_1852,In_59,In_1130);
and U1853 (N_1853,In_623,In_87);
nor U1854 (N_1854,In_1307,In_922);
or U1855 (N_1855,In_1056,In_749);
and U1856 (N_1856,In_1365,In_1040);
and U1857 (N_1857,In_1228,In_145);
nand U1858 (N_1858,In_294,In_1170);
nand U1859 (N_1859,In_346,In_991);
or U1860 (N_1860,In_84,In_1454);
or U1861 (N_1861,In_528,In_795);
or U1862 (N_1862,In_552,In_509);
and U1863 (N_1863,In_357,In_804);
nor U1864 (N_1864,In_612,In_167);
nand U1865 (N_1865,In_1053,In_746);
nand U1866 (N_1866,In_956,In_921);
nor U1867 (N_1867,In_1391,In_1447);
nand U1868 (N_1868,In_846,In_731);
nor U1869 (N_1869,In_858,In_710);
or U1870 (N_1870,In_1346,In_362);
and U1871 (N_1871,In_68,In_1495);
or U1872 (N_1872,In_1463,In_16);
nand U1873 (N_1873,In_1470,In_1080);
or U1874 (N_1874,In_184,In_139);
and U1875 (N_1875,In_859,In_1307);
xor U1876 (N_1876,In_815,In_363);
nor U1877 (N_1877,In_768,In_1121);
and U1878 (N_1878,In_1016,In_484);
nor U1879 (N_1879,In_832,In_1454);
nor U1880 (N_1880,In_1006,In_1353);
and U1881 (N_1881,In_691,In_1495);
nor U1882 (N_1882,In_118,In_895);
xnor U1883 (N_1883,In_792,In_827);
xnor U1884 (N_1884,In_969,In_1460);
xnor U1885 (N_1885,In_1163,In_1475);
or U1886 (N_1886,In_923,In_203);
nor U1887 (N_1887,In_102,In_1396);
xnor U1888 (N_1888,In_566,In_828);
and U1889 (N_1889,In_1293,In_1216);
nand U1890 (N_1890,In_1277,In_1253);
or U1891 (N_1891,In_60,In_145);
nand U1892 (N_1892,In_1151,In_653);
or U1893 (N_1893,In_1002,In_705);
nand U1894 (N_1894,In_1027,In_280);
nor U1895 (N_1895,In_570,In_1250);
nand U1896 (N_1896,In_1308,In_1206);
nand U1897 (N_1897,In_63,In_459);
and U1898 (N_1898,In_82,In_1234);
or U1899 (N_1899,In_52,In_841);
nand U1900 (N_1900,In_1456,In_1013);
or U1901 (N_1901,In_474,In_1050);
nand U1902 (N_1902,In_1291,In_1356);
and U1903 (N_1903,In_1411,In_890);
nand U1904 (N_1904,In_52,In_1401);
and U1905 (N_1905,In_990,In_399);
nor U1906 (N_1906,In_952,In_272);
nor U1907 (N_1907,In_529,In_1449);
and U1908 (N_1908,In_70,In_1334);
or U1909 (N_1909,In_1365,In_1453);
nand U1910 (N_1910,In_1056,In_907);
or U1911 (N_1911,In_236,In_169);
nor U1912 (N_1912,In_466,In_1231);
xnor U1913 (N_1913,In_336,In_1324);
and U1914 (N_1914,In_884,In_1265);
nor U1915 (N_1915,In_267,In_796);
nand U1916 (N_1916,In_1198,In_693);
and U1917 (N_1917,In_393,In_1368);
nor U1918 (N_1918,In_109,In_434);
or U1919 (N_1919,In_403,In_1058);
nor U1920 (N_1920,In_938,In_632);
and U1921 (N_1921,In_1057,In_1341);
or U1922 (N_1922,In_450,In_265);
nor U1923 (N_1923,In_535,In_469);
and U1924 (N_1924,In_398,In_568);
and U1925 (N_1925,In_725,In_16);
and U1926 (N_1926,In_44,In_1366);
nor U1927 (N_1927,In_83,In_1083);
xor U1928 (N_1928,In_613,In_934);
xor U1929 (N_1929,In_918,In_513);
nor U1930 (N_1930,In_1054,In_802);
and U1931 (N_1931,In_965,In_94);
nand U1932 (N_1932,In_1092,In_361);
or U1933 (N_1933,In_921,In_254);
nand U1934 (N_1934,In_782,In_941);
and U1935 (N_1935,In_204,In_523);
and U1936 (N_1936,In_1431,In_767);
and U1937 (N_1937,In_1277,In_346);
nor U1938 (N_1938,In_277,In_284);
or U1939 (N_1939,In_432,In_709);
nand U1940 (N_1940,In_576,In_1314);
and U1941 (N_1941,In_1280,In_544);
nand U1942 (N_1942,In_413,In_1212);
or U1943 (N_1943,In_98,In_548);
nor U1944 (N_1944,In_55,In_198);
nor U1945 (N_1945,In_109,In_216);
xnor U1946 (N_1946,In_902,In_1374);
and U1947 (N_1947,In_1388,In_896);
or U1948 (N_1948,In_1158,In_276);
nor U1949 (N_1949,In_897,In_1091);
nor U1950 (N_1950,In_219,In_253);
nor U1951 (N_1951,In_464,In_626);
or U1952 (N_1952,In_291,In_805);
nor U1953 (N_1953,In_366,In_257);
nor U1954 (N_1954,In_1380,In_191);
and U1955 (N_1955,In_95,In_392);
nor U1956 (N_1956,In_117,In_799);
nand U1957 (N_1957,In_138,In_1335);
and U1958 (N_1958,In_1308,In_668);
and U1959 (N_1959,In_1053,In_167);
nor U1960 (N_1960,In_510,In_1227);
nand U1961 (N_1961,In_137,In_1066);
nor U1962 (N_1962,In_543,In_838);
and U1963 (N_1963,In_1399,In_264);
and U1964 (N_1964,In_883,In_825);
nor U1965 (N_1965,In_855,In_898);
nor U1966 (N_1966,In_876,In_1262);
and U1967 (N_1967,In_592,In_489);
or U1968 (N_1968,In_542,In_373);
or U1969 (N_1969,In_413,In_573);
xor U1970 (N_1970,In_664,In_46);
and U1971 (N_1971,In_423,In_76);
nor U1972 (N_1972,In_27,In_964);
nand U1973 (N_1973,In_186,In_1435);
and U1974 (N_1974,In_641,In_381);
nor U1975 (N_1975,In_1214,In_422);
or U1976 (N_1976,In_1227,In_0);
or U1977 (N_1977,In_507,In_1266);
nand U1978 (N_1978,In_857,In_1353);
and U1979 (N_1979,In_181,In_1272);
and U1980 (N_1980,In_1253,In_976);
nand U1981 (N_1981,In_778,In_338);
nand U1982 (N_1982,In_17,In_559);
nor U1983 (N_1983,In_873,In_1301);
or U1984 (N_1984,In_272,In_1153);
nand U1985 (N_1985,In_476,In_902);
nor U1986 (N_1986,In_456,In_1303);
nand U1987 (N_1987,In_287,In_519);
or U1988 (N_1988,In_67,In_128);
nor U1989 (N_1989,In_1229,In_91);
and U1990 (N_1990,In_1379,In_640);
and U1991 (N_1991,In_1303,In_116);
nor U1992 (N_1992,In_848,In_668);
or U1993 (N_1993,In_1003,In_791);
or U1994 (N_1994,In_154,In_147);
nor U1995 (N_1995,In_1054,In_523);
and U1996 (N_1996,In_1302,In_940);
and U1997 (N_1997,In_996,In_314);
and U1998 (N_1998,In_212,In_1160);
xnor U1999 (N_1999,In_1082,In_1178);
nor U2000 (N_2000,In_693,In_1395);
nor U2001 (N_2001,In_612,In_1261);
nor U2002 (N_2002,In_410,In_783);
nor U2003 (N_2003,In_1475,In_47);
nor U2004 (N_2004,In_318,In_1475);
nor U2005 (N_2005,In_742,In_493);
and U2006 (N_2006,In_83,In_708);
or U2007 (N_2007,In_247,In_1383);
nand U2008 (N_2008,In_625,In_952);
nor U2009 (N_2009,In_427,In_153);
nand U2010 (N_2010,In_1134,In_1064);
nor U2011 (N_2011,In_25,In_973);
nor U2012 (N_2012,In_25,In_1360);
nor U2013 (N_2013,In_56,In_1492);
nand U2014 (N_2014,In_1308,In_768);
or U2015 (N_2015,In_1026,In_1066);
nand U2016 (N_2016,In_484,In_927);
or U2017 (N_2017,In_1016,In_623);
nor U2018 (N_2018,In_1431,In_665);
nor U2019 (N_2019,In_208,In_677);
nor U2020 (N_2020,In_1201,In_165);
nor U2021 (N_2021,In_521,In_726);
nor U2022 (N_2022,In_952,In_831);
nand U2023 (N_2023,In_705,In_655);
nand U2024 (N_2024,In_203,In_663);
nor U2025 (N_2025,In_460,In_443);
nand U2026 (N_2026,In_680,In_905);
and U2027 (N_2027,In_1365,In_731);
and U2028 (N_2028,In_656,In_1482);
nor U2029 (N_2029,In_287,In_1026);
and U2030 (N_2030,In_825,In_735);
and U2031 (N_2031,In_437,In_80);
and U2032 (N_2032,In_286,In_1490);
or U2033 (N_2033,In_52,In_1367);
xor U2034 (N_2034,In_62,In_506);
nand U2035 (N_2035,In_685,In_0);
xor U2036 (N_2036,In_883,In_1260);
xor U2037 (N_2037,In_347,In_1415);
nand U2038 (N_2038,In_601,In_879);
nand U2039 (N_2039,In_623,In_662);
nand U2040 (N_2040,In_349,In_496);
or U2041 (N_2041,In_1391,In_685);
or U2042 (N_2042,In_1341,In_775);
and U2043 (N_2043,In_709,In_313);
or U2044 (N_2044,In_1052,In_1207);
and U2045 (N_2045,In_1092,In_248);
and U2046 (N_2046,In_608,In_1221);
nand U2047 (N_2047,In_1259,In_1456);
xor U2048 (N_2048,In_934,In_711);
and U2049 (N_2049,In_821,In_574);
or U2050 (N_2050,In_956,In_287);
or U2051 (N_2051,In_1055,In_483);
or U2052 (N_2052,In_609,In_1420);
or U2053 (N_2053,In_606,In_373);
or U2054 (N_2054,In_890,In_197);
or U2055 (N_2055,In_147,In_1177);
or U2056 (N_2056,In_1161,In_262);
or U2057 (N_2057,In_936,In_749);
or U2058 (N_2058,In_494,In_469);
and U2059 (N_2059,In_255,In_510);
xnor U2060 (N_2060,In_1283,In_62);
or U2061 (N_2061,In_89,In_1493);
nor U2062 (N_2062,In_1311,In_992);
nand U2063 (N_2063,In_150,In_1117);
nor U2064 (N_2064,In_1247,In_160);
nand U2065 (N_2065,In_203,In_892);
nor U2066 (N_2066,In_260,In_594);
and U2067 (N_2067,In_1126,In_683);
nand U2068 (N_2068,In_629,In_824);
nor U2069 (N_2069,In_8,In_625);
nand U2070 (N_2070,In_971,In_274);
xnor U2071 (N_2071,In_716,In_1176);
and U2072 (N_2072,In_570,In_329);
nor U2073 (N_2073,In_1013,In_909);
nor U2074 (N_2074,In_244,In_734);
nor U2075 (N_2075,In_1338,In_910);
nor U2076 (N_2076,In_97,In_144);
and U2077 (N_2077,In_216,In_1117);
xnor U2078 (N_2078,In_1289,In_791);
and U2079 (N_2079,In_767,In_1380);
and U2080 (N_2080,In_479,In_1334);
nand U2081 (N_2081,In_1457,In_1367);
nor U2082 (N_2082,In_892,In_760);
and U2083 (N_2083,In_1326,In_18);
or U2084 (N_2084,In_1315,In_1094);
nor U2085 (N_2085,In_230,In_1190);
nor U2086 (N_2086,In_1433,In_260);
nand U2087 (N_2087,In_1184,In_349);
nand U2088 (N_2088,In_1497,In_864);
nand U2089 (N_2089,In_158,In_1187);
and U2090 (N_2090,In_775,In_1458);
or U2091 (N_2091,In_350,In_808);
xnor U2092 (N_2092,In_949,In_1142);
or U2093 (N_2093,In_642,In_381);
nor U2094 (N_2094,In_533,In_1356);
or U2095 (N_2095,In_593,In_50);
nor U2096 (N_2096,In_1382,In_1223);
nor U2097 (N_2097,In_1317,In_1386);
nand U2098 (N_2098,In_829,In_1474);
nor U2099 (N_2099,In_600,In_959);
nor U2100 (N_2100,In_634,In_1264);
or U2101 (N_2101,In_660,In_1099);
nand U2102 (N_2102,In_767,In_1456);
nor U2103 (N_2103,In_822,In_957);
nor U2104 (N_2104,In_1354,In_713);
xnor U2105 (N_2105,In_361,In_885);
nand U2106 (N_2106,In_1312,In_399);
nor U2107 (N_2107,In_353,In_682);
nand U2108 (N_2108,In_905,In_938);
nand U2109 (N_2109,In_369,In_779);
or U2110 (N_2110,In_210,In_1386);
nand U2111 (N_2111,In_381,In_537);
nor U2112 (N_2112,In_366,In_355);
nand U2113 (N_2113,In_1095,In_501);
and U2114 (N_2114,In_882,In_601);
nand U2115 (N_2115,In_223,In_535);
nand U2116 (N_2116,In_8,In_682);
xnor U2117 (N_2117,In_763,In_1057);
xor U2118 (N_2118,In_651,In_61);
and U2119 (N_2119,In_1251,In_95);
and U2120 (N_2120,In_686,In_570);
nand U2121 (N_2121,In_374,In_94);
and U2122 (N_2122,In_555,In_197);
nand U2123 (N_2123,In_450,In_1168);
nor U2124 (N_2124,In_1485,In_981);
nor U2125 (N_2125,In_1376,In_225);
xnor U2126 (N_2126,In_906,In_331);
nor U2127 (N_2127,In_621,In_811);
nand U2128 (N_2128,In_507,In_430);
nor U2129 (N_2129,In_796,In_975);
and U2130 (N_2130,In_532,In_786);
nand U2131 (N_2131,In_1004,In_322);
nor U2132 (N_2132,In_1175,In_241);
xor U2133 (N_2133,In_451,In_660);
and U2134 (N_2134,In_109,In_1370);
nor U2135 (N_2135,In_351,In_645);
nand U2136 (N_2136,In_1279,In_786);
and U2137 (N_2137,In_509,In_732);
or U2138 (N_2138,In_78,In_391);
and U2139 (N_2139,In_1156,In_1222);
and U2140 (N_2140,In_918,In_913);
and U2141 (N_2141,In_751,In_1270);
nor U2142 (N_2142,In_1448,In_1130);
and U2143 (N_2143,In_252,In_832);
and U2144 (N_2144,In_185,In_395);
and U2145 (N_2145,In_639,In_528);
xnor U2146 (N_2146,In_270,In_548);
nor U2147 (N_2147,In_1033,In_505);
and U2148 (N_2148,In_300,In_910);
or U2149 (N_2149,In_1180,In_1452);
and U2150 (N_2150,In_181,In_1379);
and U2151 (N_2151,In_1001,In_1057);
nor U2152 (N_2152,In_1309,In_767);
or U2153 (N_2153,In_385,In_491);
nor U2154 (N_2154,In_572,In_561);
or U2155 (N_2155,In_1265,In_1422);
or U2156 (N_2156,In_819,In_671);
nand U2157 (N_2157,In_1144,In_87);
nor U2158 (N_2158,In_252,In_174);
and U2159 (N_2159,In_707,In_1066);
or U2160 (N_2160,In_799,In_1424);
xnor U2161 (N_2161,In_682,In_561);
and U2162 (N_2162,In_533,In_306);
xor U2163 (N_2163,In_733,In_978);
and U2164 (N_2164,In_1064,In_989);
nand U2165 (N_2165,In_587,In_892);
nor U2166 (N_2166,In_552,In_106);
nand U2167 (N_2167,In_985,In_645);
and U2168 (N_2168,In_22,In_720);
nand U2169 (N_2169,In_432,In_56);
or U2170 (N_2170,In_837,In_525);
nor U2171 (N_2171,In_613,In_201);
nor U2172 (N_2172,In_807,In_1272);
and U2173 (N_2173,In_477,In_197);
nor U2174 (N_2174,In_294,In_1371);
nand U2175 (N_2175,In_205,In_484);
nand U2176 (N_2176,In_318,In_1327);
or U2177 (N_2177,In_563,In_363);
and U2178 (N_2178,In_680,In_930);
nand U2179 (N_2179,In_1426,In_156);
xor U2180 (N_2180,In_224,In_263);
nand U2181 (N_2181,In_399,In_623);
and U2182 (N_2182,In_1410,In_74);
and U2183 (N_2183,In_1204,In_112);
and U2184 (N_2184,In_567,In_651);
nor U2185 (N_2185,In_659,In_1256);
and U2186 (N_2186,In_8,In_1183);
and U2187 (N_2187,In_1126,In_168);
and U2188 (N_2188,In_1387,In_990);
nor U2189 (N_2189,In_83,In_1302);
nor U2190 (N_2190,In_1001,In_752);
nand U2191 (N_2191,In_1431,In_1071);
nand U2192 (N_2192,In_275,In_725);
and U2193 (N_2193,In_248,In_352);
nor U2194 (N_2194,In_92,In_1178);
or U2195 (N_2195,In_1454,In_1277);
and U2196 (N_2196,In_1133,In_647);
and U2197 (N_2197,In_1471,In_260);
nand U2198 (N_2198,In_328,In_382);
and U2199 (N_2199,In_1228,In_394);
and U2200 (N_2200,In_907,In_225);
or U2201 (N_2201,In_655,In_576);
nand U2202 (N_2202,In_322,In_1272);
and U2203 (N_2203,In_729,In_142);
and U2204 (N_2204,In_1461,In_59);
xnor U2205 (N_2205,In_1100,In_183);
or U2206 (N_2206,In_959,In_417);
nand U2207 (N_2207,In_1437,In_1164);
nor U2208 (N_2208,In_418,In_1404);
and U2209 (N_2209,In_297,In_275);
nand U2210 (N_2210,In_435,In_1435);
nand U2211 (N_2211,In_1273,In_1389);
and U2212 (N_2212,In_921,In_1221);
and U2213 (N_2213,In_209,In_1341);
nor U2214 (N_2214,In_601,In_461);
and U2215 (N_2215,In_601,In_733);
or U2216 (N_2216,In_245,In_573);
nor U2217 (N_2217,In_163,In_641);
or U2218 (N_2218,In_215,In_170);
and U2219 (N_2219,In_1144,In_1114);
nor U2220 (N_2220,In_206,In_124);
or U2221 (N_2221,In_94,In_159);
xnor U2222 (N_2222,In_942,In_900);
and U2223 (N_2223,In_602,In_1312);
nor U2224 (N_2224,In_872,In_912);
nand U2225 (N_2225,In_854,In_1323);
nor U2226 (N_2226,In_551,In_972);
nand U2227 (N_2227,In_911,In_534);
nand U2228 (N_2228,In_1067,In_670);
nor U2229 (N_2229,In_138,In_119);
or U2230 (N_2230,In_471,In_454);
or U2231 (N_2231,In_1064,In_844);
xor U2232 (N_2232,In_1161,In_1166);
nand U2233 (N_2233,In_667,In_29);
nor U2234 (N_2234,In_304,In_572);
and U2235 (N_2235,In_302,In_1294);
nor U2236 (N_2236,In_1032,In_657);
and U2237 (N_2237,In_1458,In_47);
and U2238 (N_2238,In_379,In_739);
nand U2239 (N_2239,In_1141,In_410);
xnor U2240 (N_2240,In_450,In_425);
or U2241 (N_2241,In_50,In_196);
and U2242 (N_2242,In_1420,In_541);
nand U2243 (N_2243,In_1165,In_806);
or U2244 (N_2244,In_1468,In_1000);
nand U2245 (N_2245,In_968,In_794);
or U2246 (N_2246,In_173,In_745);
nand U2247 (N_2247,In_1190,In_263);
xor U2248 (N_2248,In_1144,In_1191);
or U2249 (N_2249,In_344,In_148);
or U2250 (N_2250,In_600,In_680);
and U2251 (N_2251,In_552,In_423);
nand U2252 (N_2252,In_461,In_619);
nor U2253 (N_2253,In_904,In_985);
xnor U2254 (N_2254,In_0,In_112);
nor U2255 (N_2255,In_970,In_1174);
nand U2256 (N_2256,In_699,In_993);
nor U2257 (N_2257,In_1010,In_1137);
nand U2258 (N_2258,In_825,In_831);
and U2259 (N_2259,In_1376,In_102);
nor U2260 (N_2260,In_178,In_295);
xnor U2261 (N_2261,In_698,In_906);
and U2262 (N_2262,In_826,In_699);
and U2263 (N_2263,In_1294,In_1190);
nor U2264 (N_2264,In_1441,In_812);
or U2265 (N_2265,In_370,In_1098);
and U2266 (N_2266,In_834,In_1332);
nor U2267 (N_2267,In_329,In_15);
nor U2268 (N_2268,In_244,In_1080);
and U2269 (N_2269,In_1173,In_1404);
xor U2270 (N_2270,In_102,In_1252);
and U2271 (N_2271,In_885,In_524);
nand U2272 (N_2272,In_645,In_1279);
and U2273 (N_2273,In_463,In_444);
nand U2274 (N_2274,In_140,In_132);
xor U2275 (N_2275,In_957,In_520);
and U2276 (N_2276,In_1360,In_630);
or U2277 (N_2277,In_381,In_88);
or U2278 (N_2278,In_328,In_106);
nor U2279 (N_2279,In_977,In_174);
nand U2280 (N_2280,In_417,In_1043);
and U2281 (N_2281,In_894,In_59);
and U2282 (N_2282,In_444,In_259);
or U2283 (N_2283,In_582,In_18);
nand U2284 (N_2284,In_1431,In_1328);
or U2285 (N_2285,In_1408,In_290);
nor U2286 (N_2286,In_843,In_280);
nor U2287 (N_2287,In_997,In_777);
nand U2288 (N_2288,In_1173,In_557);
nor U2289 (N_2289,In_1225,In_1210);
nand U2290 (N_2290,In_707,In_577);
nand U2291 (N_2291,In_298,In_406);
xor U2292 (N_2292,In_1241,In_396);
or U2293 (N_2293,In_1016,In_457);
nand U2294 (N_2294,In_1143,In_696);
or U2295 (N_2295,In_1341,In_968);
nand U2296 (N_2296,In_620,In_1263);
and U2297 (N_2297,In_213,In_968);
nor U2298 (N_2298,In_1078,In_103);
nor U2299 (N_2299,In_447,In_1140);
nor U2300 (N_2300,In_508,In_855);
nor U2301 (N_2301,In_1198,In_558);
or U2302 (N_2302,In_1275,In_517);
nor U2303 (N_2303,In_849,In_215);
nor U2304 (N_2304,In_775,In_1207);
and U2305 (N_2305,In_14,In_1226);
or U2306 (N_2306,In_70,In_175);
xnor U2307 (N_2307,In_614,In_1216);
nand U2308 (N_2308,In_579,In_1104);
and U2309 (N_2309,In_748,In_847);
nor U2310 (N_2310,In_393,In_558);
nor U2311 (N_2311,In_88,In_871);
and U2312 (N_2312,In_896,In_1185);
and U2313 (N_2313,In_91,In_1242);
nand U2314 (N_2314,In_1402,In_583);
nor U2315 (N_2315,In_295,In_1239);
or U2316 (N_2316,In_1314,In_449);
nor U2317 (N_2317,In_544,In_114);
and U2318 (N_2318,In_248,In_1363);
or U2319 (N_2319,In_1056,In_832);
or U2320 (N_2320,In_681,In_903);
or U2321 (N_2321,In_1401,In_818);
or U2322 (N_2322,In_186,In_1304);
or U2323 (N_2323,In_959,In_1403);
and U2324 (N_2324,In_660,In_454);
xor U2325 (N_2325,In_67,In_152);
nor U2326 (N_2326,In_1259,In_598);
nor U2327 (N_2327,In_287,In_1280);
nor U2328 (N_2328,In_328,In_711);
and U2329 (N_2329,In_1316,In_884);
xnor U2330 (N_2330,In_1071,In_498);
nand U2331 (N_2331,In_676,In_58);
or U2332 (N_2332,In_743,In_1208);
or U2333 (N_2333,In_96,In_473);
and U2334 (N_2334,In_163,In_1127);
and U2335 (N_2335,In_1475,In_683);
or U2336 (N_2336,In_1391,In_304);
nand U2337 (N_2337,In_1143,In_699);
nand U2338 (N_2338,In_1450,In_1326);
nor U2339 (N_2339,In_1067,In_765);
or U2340 (N_2340,In_678,In_1445);
or U2341 (N_2341,In_725,In_829);
nor U2342 (N_2342,In_1035,In_103);
or U2343 (N_2343,In_526,In_81);
or U2344 (N_2344,In_85,In_167);
nor U2345 (N_2345,In_1429,In_56);
nand U2346 (N_2346,In_1377,In_580);
and U2347 (N_2347,In_1289,In_888);
and U2348 (N_2348,In_252,In_1475);
and U2349 (N_2349,In_1023,In_582);
and U2350 (N_2350,In_648,In_147);
and U2351 (N_2351,In_1373,In_1052);
or U2352 (N_2352,In_530,In_643);
or U2353 (N_2353,In_843,In_50);
or U2354 (N_2354,In_707,In_695);
nand U2355 (N_2355,In_355,In_972);
and U2356 (N_2356,In_897,In_1487);
xor U2357 (N_2357,In_186,In_414);
and U2358 (N_2358,In_488,In_330);
or U2359 (N_2359,In_1006,In_808);
nand U2360 (N_2360,In_1045,In_456);
and U2361 (N_2361,In_1423,In_614);
nor U2362 (N_2362,In_785,In_999);
or U2363 (N_2363,In_1135,In_204);
and U2364 (N_2364,In_453,In_1397);
nand U2365 (N_2365,In_1203,In_411);
or U2366 (N_2366,In_310,In_1469);
or U2367 (N_2367,In_679,In_706);
xnor U2368 (N_2368,In_995,In_110);
or U2369 (N_2369,In_526,In_683);
or U2370 (N_2370,In_363,In_913);
nand U2371 (N_2371,In_965,In_1480);
nor U2372 (N_2372,In_1487,In_256);
nor U2373 (N_2373,In_539,In_248);
nor U2374 (N_2374,In_314,In_149);
or U2375 (N_2375,In_529,In_1160);
or U2376 (N_2376,In_129,In_1317);
nor U2377 (N_2377,In_992,In_1101);
nand U2378 (N_2378,In_523,In_409);
or U2379 (N_2379,In_687,In_96);
and U2380 (N_2380,In_72,In_1149);
or U2381 (N_2381,In_513,In_1321);
or U2382 (N_2382,In_274,In_1219);
and U2383 (N_2383,In_1360,In_1448);
or U2384 (N_2384,In_1104,In_357);
or U2385 (N_2385,In_268,In_967);
xor U2386 (N_2386,In_380,In_208);
xor U2387 (N_2387,In_478,In_1361);
and U2388 (N_2388,In_1106,In_116);
nor U2389 (N_2389,In_821,In_1446);
nor U2390 (N_2390,In_316,In_910);
nor U2391 (N_2391,In_1052,In_1120);
and U2392 (N_2392,In_522,In_1227);
nand U2393 (N_2393,In_1049,In_644);
nand U2394 (N_2394,In_578,In_80);
nand U2395 (N_2395,In_1436,In_366);
and U2396 (N_2396,In_1383,In_1050);
and U2397 (N_2397,In_842,In_1059);
and U2398 (N_2398,In_1062,In_278);
nand U2399 (N_2399,In_614,In_1467);
nand U2400 (N_2400,In_1142,In_1107);
nor U2401 (N_2401,In_1054,In_293);
nor U2402 (N_2402,In_1418,In_1015);
and U2403 (N_2403,In_875,In_1420);
nor U2404 (N_2404,In_204,In_1400);
or U2405 (N_2405,In_129,In_1310);
and U2406 (N_2406,In_825,In_519);
or U2407 (N_2407,In_1172,In_627);
nand U2408 (N_2408,In_595,In_1093);
xnor U2409 (N_2409,In_662,In_430);
nor U2410 (N_2410,In_149,In_756);
nor U2411 (N_2411,In_468,In_635);
nand U2412 (N_2412,In_730,In_1387);
xnor U2413 (N_2413,In_102,In_487);
and U2414 (N_2414,In_1227,In_327);
xor U2415 (N_2415,In_1346,In_1045);
and U2416 (N_2416,In_1078,In_93);
and U2417 (N_2417,In_1451,In_409);
xor U2418 (N_2418,In_314,In_597);
nand U2419 (N_2419,In_1095,In_377);
nor U2420 (N_2420,In_196,In_268);
nor U2421 (N_2421,In_811,In_1112);
nor U2422 (N_2422,In_497,In_446);
or U2423 (N_2423,In_606,In_310);
nor U2424 (N_2424,In_457,In_801);
xor U2425 (N_2425,In_511,In_721);
and U2426 (N_2426,In_1374,In_1008);
and U2427 (N_2427,In_1063,In_1425);
nor U2428 (N_2428,In_1277,In_636);
nand U2429 (N_2429,In_452,In_146);
nor U2430 (N_2430,In_1107,In_563);
nor U2431 (N_2431,In_492,In_314);
nand U2432 (N_2432,In_173,In_612);
nor U2433 (N_2433,In_803,In_484);
nor U2434 (N_2434,In_2,In_89);
or U2435 (N_2435,In_404,In_740);
nor U2436 (N_2436,In_261,In_976);
xnor U2437 (N_2437,In_1086,In_137);
nand U2438 (N_2438,In_1478,In_663);
xor U2439 (N_2439,In_386,In_481);
xnor U2440 (N_2440,In_1463,In_853);
and U2441 (N_2441,In_948,In_764);
nor U2442 (N_2442,In_911,In_261);
and U2443 (N_2443,In_687,In_54);
or U2444 (N_2444,In_831,In_344);
or U2445 (N_2445,In_313,In_1106);
and U2446 (N_2446,In_453,In_324);
nand U2447 (N_2447,In_657,In_936);
nand U2448 (N_2448,In_829,In_89);
nand U2449 (N_2449,In_150,In_336);
and U2450 (N_2450,In_99,In_1164);
or U2451 (N_2451,In_585,In_949);
nand U2452 (N_2452,In_366,In_1055);
nor U2453 (N_2453,In_617,In_581);
and U2454 (N_2454,In_21,In_771);
and U2455 (N_2455,In_879,In_1015);
xor U2456 (N_2456,In_1338,In_112);
nand U2457 (N_2457,In_1016,In_1241);
and U2458 (N_2458,In_395,In_117);
or U2459 (N_2459,In_1222,In_849);
nor U2460 (N_2460,In_1411,In_1118);
or U2461 (N_2461,In_1043,In_1028);
and U2462 (N_2462,In_1125,In_614);
or U2463 (N_2463,In_3,In_360);
or U2464 (N_2464,In_216,In_1313);
and U2465 (N_2465,In_511,In_938);
and U2466 (N_2466,In_564,In_439);
or U2467 (N_2467,In_254,In_418);
nand U2468 (N_2468,In_693,In_397);
nand U2469 (N_2469,In_976,In_822);
and U2470 (N_2470,In_838,In_502);
and U2471 (N_2471,In_293,In_854);
nand U2472 (N_2472,In_639,In_839);
and U2473 (N_2473,In_546,In_1474);
nor U2474 (N_2474,In_1336,In_779);
nor U2475 (N_2475,In_924,In_748);
xnor U2476 (N_2476,In_823,In_1489);
nor U2477 (N_2477,In_926,In_617);
nand U2478 (N_2478,In_46,In_262);
and U2479 (N_2479,In_914,In_497);
or U2480 (N_2480,In_1139,In_1128);
and U2481 (N_2481,In_606,In_999);
or U2482 (N_2482,In_765,In_1414);
or U2483 (N_2483,In_1117,In_939);
and U2484 (N_2484,In_503,In_293);
nand U2485 (N_2485,In_1316,In_979);
or U2486 (N_2486,In_1284,In_1225);
nor U2487 (N_2487,In_156,In_136);
or U2488 (N_2488,In_1464,In_677);
nand U2489 (N_2489,In_553,In_544);
or U2490 (N_2490,In_682,In_120);
nand U2491 (N_2491,In_1489,In_143);
or U2492 (N_2492,In_547,In_500);
and U2493 (N_2493,In_597,In_1018);
and U2494 (N_2494,In_902,In_1205);
and U2495 (N_2495,In_916,In_400);
and U2496 (N_2496,In_834,In_443);
nand U2497 (N_2497,In_211,In_1025);
or U2498 (N_2498,In_1482,In_61);
xnor U2499 (N_2499,In_936,In_45);
and U2500 (N_2500,In_429,In_350);
nor U2501 (N_2501,In_754,In_656);
nor U2502 (N_2502,In_814,In_1251);
or U2503 (N_2503,In_621,In_32);
nor U2504 (N_2504,In_1127,In_992);
nand U2505 (N_2505,In_67,In_914);
and U2506 (N_2506,In_1477,In_1256);
or U2507 (N_2507,In_278,In_1049);
xor U2508 (N_2508,In_403,In_744);
nor U2509 (N_2509,In_1204,In_1085);
nor U2510 (N_2510,In_74,In_554);
or U2511 (N_2511,In_1085,In_1209);
or U2512 (N_2512,In_21,In_795);
nor U2513 (N_2513,In_159,In_744);
nor U2514 (N_2514,In_111,In_958);
and U2515 (N_2515,In_850,In_107);
nand U2516 (N_2516,In_330,In_812);
nand U2517 (N_2517,In_95,In_523);
nand U2518 (N_2518,In_1133,In_1293);
nor U2519 (N_2519,In_370,In_789);
and U2520 (N_2520,In_1482,In_462);
xor U2521 (N_2521,In_844,In_184);
and U2522 (N_2522,In_1084,In_177);
nor U2523 (N_2523,In_1167,In_254);
and U2524 (N_2524,In_906,In_239);
nor U2525 (N_2525,In_1254,In_140);
nand U2526 (N_2526,In_1446,In_462);
or U2527 (N_2527,In_347,In_1338);
xor U2528 (N_2528,In_775,In_530);
and U2529 (N_2529,In_321,In_1092);
or U2530 (N_2530,In_870,In_441);
and U2531 (N_2531,In_264,In_988);
and U2532 (N_2532,In_882,In_1456);
or U2533 (N_2533,In_195,In_1397);
or U2534 (N_2534,In_363,In_820);
nor U2535 (N_2535,In_423,In_5);
nor U2536 (N_2536,In_148,In_1118);
or U2537 (N_2537,In_1014,In_1349);
nand U2538 (N_2538,In_1062,In_628);
nand U2539 (N_2539,In_366,In_662);
nand U2540 (N_2540,In_884,In_976);
nand U2541 (N_2541,In_862,In_1268);
nor U2542 (N_2542,In_1013,In_1135);
nand U2543 (N_2543,In_729,In_290);
or U2544 (N_2544,In_93,In_566);
and U2545 (N_2545,In_569,In_1009);
nor U2546 (N_2546,In_1140,In_1249);
and U2547 (N_2547,In_542,In_425);
nand U2548 (N_2548,In_534,In_892);
or U2549 (N_2549,In_276,In_310);
xor U2550 (N_2550,In_1278,In_753);
nor U2551 (N_2551,In_1168,In_857);
nand U2552 (N_2552,In_426,In_1315);
nor U2553 (N_2553,In_1269,In_1085);
nor U2554 (N_2554,In_1008,In_1184);
or U2555 (N_2555,In_951,In_22);
and U2556 (N_2556,In_456,In_1386);
or U2557 (N_2557,In_551,In_557);
nand U2558 (N_2558,In_105,In_752);
xor U2559 (N_2559,In_1362,In_983);
and U2560 (N_2560,In_215,In_100);
and U2561 (N_2561,In_1473,In_932);
and U2562 (N_2562,In_501,In_683);
or U2563 (N_2563,In_1427,In_597);
nor U2564 (N_2564,In_151,In_692);
and U2565 (N_2565,In_258,In_1069);
nor U2566 (N_2566,In_296,In_582);
nor U2567 (N_2567,In_1442,In_416);
xnor U2568 (N_2568,In_843,In_180);
nor U2569 (N_2569,In_564,In_719);
nor U2570 (N_2570,In_896,In_1034);
nand U2571 (N_2571,In_1250,In_867);
and U2572 (N_2572,In_1494,In_616);
and U2573 (N_2573,In_1418,In_425);
nand U2574 (N_2574,In_859,In_631);
nand U2575 (N_2575,In_253,In_886);
xor U2576 (N_2576,In_1014,In_535);
xor U2577 (N_2577,In_440,In_253);
and U2578 (N_2578,In_223,In_470);
nor U2579 (N_2579,In_1381,In_206);
xor U2580 (N_2580,In_887,In_1264);
nand U2581 (N_2581,In_963,In_673);
nand U2582 (N_2582,In_350,In_374);
nand U2583 (N_2583,In_1001,In_315);
xnor U2584 (N_2584,In_1103,In_775);
or U2585 (N_2585,In_95,In_790);
nor U2586 (N_2586,In_623,In_232);
or U2587 (N_2587,In_59,In_387);
nor U2588 (N_2588,In_1330,In_418);
and U2589 (N_2589,In_1173,In_520);
nand U2590 (N_2590,In_526,In_877);
nand U2591 (N_2591,In_207,In_1355);
xnor U2592 (N_2592,In_997,In_1420);
nand U2593 (N_2593,In_1327,In_717);
or U2594 (N_2594,In_61,In_1456);
nor U2595 (N_2595,In_403,In_393);
nand U2596 (N_2596,In_711,In_1023);
nand U2597 (N_2597,In_14,In_631);
and U2598 (N_2598,In_1362,In_878);
or U2599 (N_2599,In_1383,In_728);
nand U2600 (N_2600,In_191,In_1277);
nand U2601 (N_2601,In_1018,In_1095);
and U2602 (N_2602,In_705,In_1240);
and U2603 (N_2603,In_197,In_1491);
nand U2604 (N_2604,In_303,In_648);
nor U2605 (N_2605,In_1143,In_225);
nand U2606 (N_2606,In_647,In_838);
nor U2607 (N_2607,In_927,In_734);
nand U2608 (N_2608,In_232,In_644);
nor U2609 (N_2609,In_1363,In_1397);
xor U2610 (N_2610,In_433,In_303);
nor U2611 (N_2611,In_1335,In_767);
nor U2612 (N_2612,In_1106,In_312);
nor U2613 (N_2613,In_1058,In_587);
or U2614 (N_2614,In_545,In_213);
and U2615 (N_2615,In_895,In_888);
and U2616 (N_2616,In_865,In_1315);
nand U2617 (N_2617,In_1170,In_1490);
nand U2618 (N_2618,In_1041,In_774);
and U2619 (N_2619,In_1066,In_110);
xnor U2620 (N_2620,In_445,In_419);
nand U2621 (N_2621,In_849,In_1204);
or U2622 (N_2622,In_302,In_1319);
or U2623 (N_2623,In_1300,In_535);
and U2624 (N_2624,In_453,In_319);
and U2625 (N_2625,In_1170,In_987);
nand U2626 (N_2626,In_792,In_474);
nor U2627 (N_2627,In_1122,In_713);
nor U2628 (N_2628,In_1290,In_958);
or U2629 (N_2629,In_1384,In_105);
nor U2630 (N_2630,In_1200,In_464);
and U2631 (N_2631,In_113,In_952);
and U2632 (N_2632,In_9,In_1016);
nand U2633 (N_2633,In_687,In_1440);
xnor U2634 (N_2634,In_1083,In_324);
and U2635 (N_2635,In_555,In_1407);
nand U2636 (N_2636,In_345,In_946);
nand U2637 (N_2637,In_405,In_1344);
and U2638 (N_2638,In_190,In_939);
nor U2639 (N_2639,In_802,In_683);
nor U2640 (N_2640,In_1072,In_1234);
nor U2641 (N_2641,In_988,In_368);
and U2642 (N_2642,In_659,In_375);
xor U2643 (N_2643,In_1336,In_1349);
nand U2644 (N_2644,In_1010,In_749);
nand U2645 (N_2645,In_348,In_1340);
and U2646 (N_2646,In_131,In_1219);
or U2647 (N_2647,In_22,In_616);
nor U2648 (N_2648,In_734,In_299);
nand U2649 (N_2649,In_109,In_743);
and U2650 (N_2650,In_393,In_566);
or U2651 (N_2651,In_930,In_1017);
nand U2652 (N_2652,In_1404,In_954);
nor U2653 (N_2653,In_909,In_1473);
xor U2654 (N_2654,In_1101,In_279);
or U2655 (N_2655,In_506,In_689);
nand U2656 (N_2656,In_1314,In_1302);
or U2657 (N_2657,In_1031,In_498);
and U2658 (N_2658,In_927,In_1341);
and U2659 (N_2659,In_895,In_498);
xor U2660 (N_2660,In_457,In_114);
or U2661 (N_2661,In_1144,In_1023);
or U2662 (N_2662,In_765,In_1386);
nor U2663 (N_2663,In_1142,In_61);
nand U2664 (N_2664,In_1462,In_826);
and U2665 (N_2665,In_78,In_1141);
nor U2666 (N_2666,In_1110,In_668);
xor U2667 (N_2667,In_1230,In_1387);
or U2668 (N_2668,In_1353,In_762);
nand U2669 (N_2669,In_440,In_1494);
nand U2670 (N_2670,In_954,In_713);
nor U2671 (N_2671,In_521,In_865);
or U2672 (N_2672,In_77,In_420);
or U2673 (N_2673,In_410,In_891);
or U2674 (N_2674,In_929,In_495);
or U2675 (N_2675,In_72,In_628);
or U2676 (N_2676,In_1327,In_1100);
and U2677 (N_2677,In_142,In_494);
or U2678 (N_2678,In_277,In_1180);
and U2679 (N_2679,In_1424,In_375);
or U2680 (N_2680,In_387,In_1327);
nand U2681 (N_2681,In_602,In_233);
nor U2682 (N_2682,In_306,In_1027);
nor U2683 (N_2683,In_55,In_1158);
nand U2684 (N_2684,In_719,In_291);
or U2685 (N_2685,In_687,In_1421);
and U2686 (N_2686,In_231,In_71);
and U2687 (N_2687,In_1179,In_1238);
nand U2688 (N_2688,In_1004,In_1470);
nand U2689 (N_2689,In_839,In_1343);
nand U2690 (N_2690,In_795,In_1198);
or U2691 (N_2691,In_671,In_1435);
xnor U2692 (N_2692,In_176,In_1410);
and U2693 (N_2693,In_385,In_665);
nand U2694 (N_2694,In_512,In_853);
or U2695 (N_2695,In_809,In_933);
or U2696 (N_2696,In_1317,In_281);
nand U2697 (N_2697,In_944,In_1077);
nand U2698 (N_2698,In_1,In_739);
or U2699 (N_2699,In_632,In_293);
xor U2700 (N_2700,In_263,In_1030);
and U2701 (N_2701,In_232,In_745);
nor U2702 (N_2702,In_156,In_1165);
or U2703 (N_2703,In_415,In_1019);
nand U2704 (N_2704,In_1072,In_950);
nor U2705 (N_2705,In_1453,In_1447);
nor U2706 (N_2706,In_1314,In_1082);
and U2707 (N_2707,In_1115,In_611);
and U2708 (N_2708,In_552,In_138);
and U2709 (N_2709,In_1139,In_978);
or U2710 (N_2710,In_73,In_37);
xnor U2711 (N_2711,In_184,In_663);
nor U2712 (N_2712,In_222,In_424);
nand U2713 (N_2713,In_1346,In_670);
or U2714 (N_2714,In_189,In_83);
nor U2715 (N_2715,In_755,In_308);
nand U2716 (N_2716,In_751,In_316);
and U2717 (N_2717,In_335,In_908);
and U2718 (N_2718,In_795,In_928);
or U2719 (N_2719,In_1357,In_634);
nand U2720 (N_2720,In_1139,In_1349);
and U2721 (N_2721,In_998,In_799);
and U2722 (N_2722,In_1353,In_1387);
nand U2723 (N_2723,In_957,In_687);
nand U2724 (N_2724,In_1115,In_294);
and U2725 (N_2725,In_487,In_360);
and U2726 (N_2726,In_1091,In_149);
nor U2727 (N_2727,In_882,In_239);
nor U2728 (N_2728,In_421,In_615);
or U2729 (N_2729,In_873,In_1096);
and U2730 (N_2730,In_215,In_0);
nor U2731 (N_2731,In_1321,In_1209);
xnor U2732 (N_2732,In_205,In_1291);
xnor U2733 (N_2733,In_64,In_1463);
nor U2734 (N_2734,In_381,In_824);
xnor U2735 (N_2735,In_1246,In_46);
nor U2736 (N_2736,In_340,In_843);
nand U2737 (N_2737,In_92,In_1100);
and U2738 (N_2738,In_619,In_1326);
nor U2739 (N_2739,In_321,In_1301);
or U2740 (N_2740,In_1372,In_1033);
nand U2741 (N_2741,In_1229,In_1448);
nor U2742 (N_2742,In_992,In_666);
nand U2743 (N_2743,In_160,In_701);
and U2744 (N_2744,In_1037,In_964);
and U2745 (N_2745,In_981,In_492);
nand U2746 (N_2746,In_1274,In_1474);
or U2747 (N_2747,In_1092,In_731);
or U2748 (N_2748,In_290,In_697);
and U2749 (N_2749,In_355,In_21);
and U2750 (N_2750,In_718,In_1328);
or U2751 (N_2751,In_1284,In_349);
nor U2752 (N_2752,In_1142,In_846);
nand U2753 (N_2753,In_288,In_1262);
or U2754 (N_2754,In_1362,In_431);
nand U2755 (N_2755,In_198,In_1132);
or U2756 (N_2756,In_658,In_569);
nand U2757 (N_2757,In_716,In_731);
nand U2758 (N_2758,In_821,In_363);
or U2759 (N_2759,In_1074,In_1264);
and U2760 (N_2760,In_1479,In_720);
nand U2761 (N_2761,In_1046,In_925);
and U2762 (N_2762,In_946,In_1380);
nor U2763 (N_2763,In_1286,In_1033);
nand U2764 (N_2764,In_967,In_589);
nand U2765 (N_2765,In_1383,In_1217);
nor U2766 (N_2766,In_1363,In_1009);
nor U2767 (N_2767,In_447,In_329);
and U2768 (N_2768,In_826,In_773);
or U2769 (N_2769,In_611,In_1167);
nand U2770 (N_2770,In_729,In_25);
and U2771 (N_2771,In_25,In_150);
and U2772 (N_2772,In_900,In_1070);
nor U2773 (N_2773,In_227,In_337);
or U2774 (N_2774,In_701,In_1379);
xnor U2775 (N_2775,In_8,In_651);
nor U2776 (N_2776,In_1439,In_733);
xnor U2777 (N_2777,In_1108,In_1080);
nand U2778 (N_2778,In_1155,In_98);
nand U2779 (N_2779,In_610,In_691);
nand U2780 (N_2780,In_908,In_418);
or U2781 (N_2781,In_1102,In_844);
or U2782 (N_2782,In_890,In_175);
xor U2783 (N_2783,In_498,In_810);
nor U2784 (N_2784,In_1080,In_700);
or U2785 (N_2785,In_391,In_1059);
and U2786 (N_2786,In_9,In_1139);
nand U2787 (N_2787,In_224,In_971);
and U2788 (N_2788,In_31,In_26);
or U2789 (N_2789,In_909,In_1334);
and U2790 (N_2790,In_635,In_597);
nand U2791 (N_2791,In_36,In_1090);
nor U2792 (N_2792,In_314,In_266);
or U2793 (N_2793,In_562,In_1391);
nor U2794 (N_2794,In_847,In_1155);
nor U2795 (N_2795,In_1304,In_68);
nand U2796 (N_2796,In_595,In_838);
and U2797 (N_2797,In_192,In_1049);
nand U2798 (N_2798,In_1071,In_1440);
nand U2799 (N_2799,In_121,In_386);
xnor U2800 (N_2800,In_812,In_740);
or U2801 (N_2801,In_933,In_1295);
nor U2802 (N_2802,In_628,In_1199);
xnor U2803 (N_2803,In_3,In_892);
or U2804 (N_2804,In_1471,In_633);
or U2805 (N_2805,In_947,In_1186);
and U2806 (N_2806,In_1201,In_1350);
nand U2807 (N_2807,In_627,In_543);
or U2808 (N_2808,In_539,In_609);
xor U2809 (N_2809,In_873,In_907);
and U2810 (N_2810,In_1423,In_199);
and U2811 (N_2811,In_998,In_1339);
and U2812 (N_2812,In_247,In_93);
nor U2813 (N_2813,In_1426,In_1116);
or U2814 (N_2814,In_380,In_646);
or U2815 (N_2815,In_678,In_0);
or U2816 (N_2816,In_353,In_1391);
nand U2817 (N_2817,In_536,In_1190);
nor U2818 (N_2818,In_302,In_274);
or U2819 (N_2819,In_855,In_594);
xor U2820 (N_2820,In_894,In_544);
or U2821 (N_2821,In_1329,In_835);
or U2822 (N_2822,In_979,In_969);
and U2823 (N_2823,In_483,In_842);
nand U2824 (N_2824,In_483,In_814);
nor U2825 (N_2825,In_396,In_768);
nand U2826 (N_2826,In_219,In_999);
nor U2827 (N_2827,In_152,In_1362);
nand U2828 (N_2828,In_1163,In_704);
and U2829 (N_2829,In_290,In_583);
or U2830 (N_2830,In_967,In_728);
or U2831 (N_2831,In_768,In_89);
xor U2832 (N_2832,In_566,In_1181);
or U2833 (N_2833,In_884,In_41);
or U2834 (N_2834,In_613,In_797);
nand U2835 (N_2835,In_45,In_1105);
and U2836 (N_2836,In_1447,In_1093);
nor U2837 (N_2837,In_1018,In_484);
or U2838 (N_2838,In_177,In_1145);
nand U2839 (N_2839,In_43,In_856);
and U2840 (N_2840,In_758,In_748);
or U2841 (N_2841,In_538,In_642);
or U2842 (N_2842,In_1454,In_589);
or U2843 (N_2843,In_1109,In_1472);
xnor U2844 (N_2844,In_690,In_1411);
nor U2845 (N_2845,In_508,In_895);
nand U2846 (N_2846,In_1262,In_925);
or U2847 (N_2847,In_881,In_1297);
or U2848 (N_2848,In_670,In_1007);
nand U2849 (N_2849,In_257,In_1462);
nand U2850 (N_2850,In_1131,In_1241);
and U2851 (N_2851,In_353,In_717);
or U2852 (N_2852,In_74,In_686);
nor U2853 (N_2853,In_1497,In_1413);
and U2854 (N_2854,In_395,In_97);
nor U2855 (N_2855,In_974,In_713);
xor U2856 (N_2856,In_539,In_800);
nor U2857 (N_2857,In_1432,In_145);
nand U2858 (N_2858,In_864,In_938);
xnor U2859 (N_2859,In_894,In_996);
nand U2860 (N_2860,In_529,In_1147);
nand U2861 (N_2861,In_39,In_17);
or U2862 (N_2862,In_58,In_1067);
nand U2863 (N_2863,In_798,In_498);
or U2864 (N_2864,In_609,In_1173);
or U2865 (N_2865,In_835,In_949);
xor U2866 (N_2866,In_840,In_695);
or U2867 (N_2867,In_617,In_1323);
and U2868 (N_2868,In_1015,In_674);
nor U2869 (N_2869,In_151,In_762);
or U2870 (N_2870,In_1282,In_284);
nand U2871 (N_2871,In_698,In_1238);
or U2872 (N_2872,In_581,In_1298);
and U2873 (N_2873,In_1214,In_1333);
or U2874 (N_2874,In_634,In_1401);
nand U2875 (N_2875,In_536,In_897);
nand U2876 (N_2876,In_167,In_605);
or U2877 (N_2877,In_937,In_607);
nand U2878 (N_2878,In_1180,In_411);
or U2879 (N_2879,In_35,In_1155);
and U2880 (N_2880,In_1382,In_1395);
nand U2881 (N_2881,In_355,In_980);
nor U2882 (N_2882,In_1112,In_1294);
or U2883 (N_2883,In_1416,In_724);
and U2884 (N_2884,In_1151,In_932);
and U2885 (N_2885,In_789,In_598);
nand U2886 (N_2886,In_413,In_929);
and U2887 (N_2887,In_515,In_1091);
nand U2888 (N_2888,In_978,In_1119);
nand U2889 (N_2889,In_583,In_864);
and U2890 (N_2890,In_314,In_421);
nand U2891 (N_2891,In_1420,In_358);
and U2892 (N_2892,In_833,In_257);
or U2893 (N_2893,In_453,In_171);
nand U2894 (N_2894,In_1307,In_1489);
and U2895 (N_2895,In_1100,In_668);
nor U2896 (N_2896,In_245,In_1470);
and U2897 (N_2897,In_49,In_179);
or U2898 (N_2898,In_53,In_710);
or U2899 (N_2899,In_908,In_475);
or U2900 (N_2900,In_600,In_799);
and U2901 (N_2901,In_578,In_1312);
nand U2902 (N_2902,In_435,In_461);
nand U2903 (N_2903,In_884,In_1245);
nor U2904 (N_2904,In_152,In_822);
or U2905 (N_2905,In_1490,In_392);
and U2906 (N_2906,In_340,In_1460);
nand U2907 (N_2907,In_492,In_1001);
nor U2908 (N_2908,In_648,In_361);
and U2909 (N_2909,In_48,In_687);
nand U2910 (N_2910,In_1232,In_1378);
nor U2911 (N_2911,In_1322,In_655);
and U2912 (N_2912,In_741,In_996);
and U2913 (N_2913,In_806,In_1190);
and U2914 (N_2914,In_197,In_842);
or U2915 (N_2915,In_466,In_1039);
nor U2916 (N_2916,In_466,In_528);
nand U2917 (N_2917,In_777,In_659);
and U2918 (N_2918,In_776,In_848);
and U2919 (N_2919,In_1088,In_454);
nor U2920 (N_2920,In_614,In_441);
and U2921 (N_2921,In_1110,In_1363);
or U2922 (N_2922,In_345,In_1414);
and U2923 (N_2923,In_381,In_1140);
or U2924 (N_2924,In_532,In_1252);
nand U2925 (N_2925,In_799,In_1460);
nor U2926 (N_2926,In_288,In_806);
nor U2927 (N_2927,In_495,In_532);
and U2928 (N_2928,In_732,In_1303);
and U2929 (N_2929,In_1364,In_864);
and U2930 (N_2930,In_408,In_61);
or U2931 (N_2931,In_1153,In_1314);
and U2932 (N_2932,In_208,In_483);
nand U2933 (N_2933,In_1352,In_505);
and U2934 (N_2934,In_97,In_302);
nor U2935 (N_2935,In_783,In_595);
nor U2936 (N_2936,In_588,In_772);
and U2937 (N_2937,In_1056,In_745);
nand U2938 (N_2938,In_64,In_1408);
nor U2939 (N_2939,In_947,In_110);
or U2940 (N_2940,In_432,In_255);
nand U2941 (N_2941,In_1334,In_362);
and U2942 (N_2942,In_609,In_1102);
and U2943 (N_2943,In_135,In_1143);
and U2944 (N_2944,In_896,In_1030);
or U2945 (N_2945,In_765,In_38);
nor U2946 (N_2946,In_1481,In_146);
or U2947 (N_2947,In_674,In_1241);
nor U2948 (N_2948,In_11,In_1429);
nand U2949 (N_2949,In_606,In_940);
nand U2950 (N_2950,In_1087,In_999);
nand U2951 (N_2951,In_1131,In_970);
nand U2952 (N_2952,In_272,In_309);
and U2953 (N_2953,In_354,In_1272);
nor U2954 (N_2954,In_596,In_706);
and U2955 (N_2955,In_1459,In_869);
or U2956 (N_2956,In_520,In_325);
or U2957 (N_2957,In_794,In_115);
nand U2958 (N_2958,In_538,In_654);
nand U2959 (N_2959,In_207,In_960);
or U2960 (N_2960,In_174,In_36);
nor U2961 (N_2961,In_1080,In_1185);
nor U2962 (N_2962,In_33,In_1098);
xor U2963 (N_2963,In_1040,In_113);
and U2964 (N_2964,In_1027,In_1167);
or U2965 (N_2965,In_560,In_1300);
or U2966 (N_2966,In_99,In_1150);
and U2967 (N_2967,In_102,In_902);
nor U2968 (N_2968,In_1443,In_318);
or U2969 (N_2969,In_1311,In_1061);
nand U2970 (N_2970,In_943,In_1201);
or U2971 (N_2971,In_1100,In_1290);
nor U2972 (N_2972,In_775,In_499);
nand U2973 (N_2973,In_771,In_651);
or U2974 (N_2974,In_511,In_519);
and U2975 (N_2975,In_392,In_178);
nand U2976 (N_2976,In_436,In_766);
or U2977 (N_2977,In_16,In_1298);
or U2978 (N_2978,In_139,In_47);
or U2979 (N_2979,In_1048,In_605);
nor U2980 (N_2980,In_1178,In_1168);
and U2981 (N_2981,In_7,In_984);
nor U2982 (N_2982,In_888,In_438);
or U2983 (N_2983,In_1323,In_23);
and U2984 (N_2984,In_387,In_929);
and U2985 (N_2985,In_561,In_945);
xor U2986 (N_2986,In_171,In_728);
nor U2987 (N_2987,In_696,In_469);
or U2988 (N_2988,In_1034,In_1372);
nor U2989 (N_2989,In_897,In_374);
nor U2990 (N_2990,In_342,In_123);
nand U2991 (N_2991,In_992,In_630);
nand U2992 (N_2992,In_488,In_207);
nand U2993 (N_2993,In_213,In_139);
nand U2994 (N_2994,In_1306,In_1087);
or U2995 (N_2995,In_903,In_224);
nand U2996 (N_2996,In_1425,In_476);
and U2997 (N_2997,In_842,In_947);
or U2998 (N_2998,In_88,In_62);
nor U2999 (N_2999,In_268,In_1206);
and U3000 (N_3000,In_988,In_1306);
and U3001 (N_3001,In_884,In_1);
nand U3002 (N_3002,In_1029,In_899);
or U3003 (N_3003,In_591,In_1074);
xor U3004 (N_3004,In_908,In_1462);
and U3005 (N_3005,In_634,In_716);
nand U3006 (N_3006,In_349,In_91);
nor U3007 (N_3007,In_892,In_123);
or U3008 (N_3008,In_198,In_16);
nand U3009 (N_3009,In_533,In_671);
or U3010 (N_3010,In_714,In_293);
and U3011 (N_3011,In_244,In_406);
nor U3012 (N_3012,In_44,In_140);
nand U3013 (N_3013,In_853,In_872);
nand U3014 (N_3014,In_362,In_29);
xor U3015 (N_3015,In_19,In_523);
nand U3016 (N_3016,In_1002,In_158);
nand U3017 (N_3017,In_96,In_451);
xor U3018 (N_3018,In_687,In_571);
nand U3019 (N_3019,In_1138,In_227);
and U3020 (N_3020,In_767,In_586);
nor U3021 (N_3021,In_1138,In_1335);
nand U3022 (N_3022,In_650,In_38);
nor U3023 (N_3023,In_1131,In_680);
and U3024 (N_3024,In_307,In_315);
and U3025 (N_3025,In_570,In_283);
or U3026 (N_3026,In_820,In_1026);
xnor U3027 (N_3027,In_20,In_689);
or U3028 (N_3028,In_11,In_599);
nor U3029 (N_3029,In_531,In_262);
nand U3030 (N_3030,In_347,In_814);
or U3031 (N_3031,In_393,In_435);
xor U3032 (N_3032,In_667,In_1288);
xor U3033 (N_3033,In_394,In_1083);
nor U3034 (N_3034,In_724,In_1338);
and U3035 (N_3035,In_733,In_1025);
and U3036 (N_3036,In_1494,In_97);
nand U3037 (N_3037,In_856,In_561);
nand U3038 (N_3038,In_1437,In_1125);
nand U3039 (N_3039,In_684,In_769);
nor U3040 (N_3040,In_554,In_700);
nor U3041 (N_3041,In_457,In_215);
and U3042 (N_3042,In_680,In_991);
and U3043 (N_3043,In_1308,In_1113);
and U3044 (N_3044,In_213,In_367);
nor U3045 (N_3045,In_1389,In_871);
and U3046 (N_3046,In_940,In_1093);
nor U3047 (N_3047,In_970,In_224);
nand U3048 (N_3048,In_1213,In_997);
nor U3049 (N_3049,In_333,In_465);
nand U3050 (N_3050,In_1265,In_826);
and U3051 (N_3051,In_1139,In_89);
nor U3052 (N_3052,In_465,In_467);
xnor U3053 (N_3053,In_1171,In_1475);
xor U3054 (N_3054,In_1080,In_408);
and U3055 (N_3055,In_886,In_1216);
and U3056 (N_3056,In_1251,In_618);
and U3057 (N_3057,In_227,In_1430);
nand U3058 (N_3058,In_1017,In_971);
nand U3059 (N_3059,In_1187,In_1247);
nand U3060 (N_3060,In_171,In_299);
nand U3061 (N_3061,In_61,In_360);
and U3062 (N_3062,In_69,In_812);
and U3063 (N_3063,In_795,In_517);
nand U3064 (N_3064,In_619,In_1142);
xor U3065 (N_3065,In_929,In_1333);
nor U3066 (N_3066,In_1467,In_601);
and U3067 (N_3067,In_737,In_685);
xor U3068 (N_3068,In_435,In_172);
or U3069 (N_3069,In_189,In_1024);
xnor U3070 (N_3070,In_1065,In_1314);
or U3071 (N_3071,In_1177,In_61);
or U3072 (N_3072,In_244,In_38);
nand U3073 (N_3073,In_1146,In_352);
xnor U3074 (N_3074,In_260,In_1405);
nor U3075 (N_3075,In_120,In_1129);
xnor U3076 (N_3076,In_1316,In_1280);
and U3077 (N_3077,In_581,In_423);
or U3078 (N_3078,In_1113,In_274);
nor U3079 (N_3079,In_207,In_470);
nor U3080 (N_3080,In_891,In_692);
or U3081 (N_3081,In_1096,In_988);
nand U3082 (N_3082,In_852,In_1250);
and U3083 (N_3083,In_357,In_551);
and U3084 (N_3084,In_18,In_1293);
nand U3085 (N_3085,In_1205,In_994);
xor U3086 (N_3086,In_106,In_1191);
nor U3087 (N_3087,In_456,In_971);
or U3088 (N_3088,In_932,In_697);
or U3089 (N_3089,In_74,In_172);
or U3090 (N_3090,In_1380,In_627);
nor U3091 (N_3091,In_1435,In_123);
nand U3092 (N_3092,In_449,In_619);
nand U3093 (N_3093,In_34,In_919);
and U3094 (N_3094,In_861,In_322);
and U3095 (N_3095,In_830,In_1317);
xnor U3096 (N_3096,In_720,In_324);
or U3097 (N_3097,In_1030,In_914);
nor U3098 (N_3098,In_464,In_580);
nand U3099 (N_3099,In_691,In_1310);
nand U3100 (N_3100,In_116,In_301);
nor U3101 (N_3101,In_1460,In_556);
and U3102 (N_3102,In_1358,In_878);
nor U3103 (N_3103,In_1350,In_1247);
nand U3104 (N_3104,In_396,In_1208);
and U3105 (N_3105,In_1068,In_92);
or U3106 (N_3106,In_171,In_721);
nand U3107 (N_3107,In_943,In_1471);
nor U3108 (N_3108,In_1180,In_0);
nand U3109 (N_3109,In_518,In_297);
and U3110 (N_3110,In_902,In_1391);
and U3111 (N_3111,In_875,In_984);
nor U3112 (N_3112,In_913,In_397);
nor U3113 (N_3113,In_124,In_1013);
or U3114 (N_3114,In_228,In_250);
xor U3115 (N_3115,In_242,In_1295);
and U3116 (N_3116,In_832,In_879);
nor U3117 (N_3117,In_683,In_950);
xor U3118 (N_3118,In_1171,In_1437);
nand U3119 (N_3119,In_1107,In_1001);
and U3120 (N_3120,In_470,In_181);
or U3121 (N_3121,In_990,In_504);
and U3122 (N_3122,In_1475,In_888);
or U3123 (N_3123,In_505,In_109);
nand U3124 (N_3124,In_61,In_453);
nand U3125 (N_3125,In_212,In_966);
and U3126 (N_3126,In_569,In_1462);
nor U3127 (N_3127,In_786,In_1282);
or U3128 (N_3128,In_791,In_454);
nand U3129 (N_3129,In_1306,In_26);
nor U3130 (N_3130,In_608,In_1176);
or U3131 (N_3131,In_258,In_1096);
xnor U3132 (N_3132,In_896,In_1467);
nor U3133 (N_3133,In_888,In_25);
xnor U3134 (N_3134,In_1219,In_359);
nor U3135 (N_3135,In_1451,In_494);
and U3136 (N_3136,In_229,In_1250);
or U3137 (N_3137,In_491,In_1297);
nor U3138 (N_3138,In_163,In_779);
or U3139 (N_3139,In_653,In_90);
and U3140 (N_3140,In_1152,In_395);
nor U3141 (N_3141,In_132,In_1371);
or U3142 (N_3142,In_630,In_1002);
and U3143 (N_3143,In_1190,In_1490);
nor U3144 (N_3144,In_761,In_853);
nand U3145 (N_3145,In_1380,In_392);
and U3146 (N_3146,In_933,In_886);
or U3147 (N_3147,In_1146,In_195);
nand U3148 (N_3148,In_538,In_1485);
and U3149 (N_3149,In_41,In_350);
nand U3150 (N_3150,In_185,In_1080);
nor U3151 (N_3151,In_1179,In_1210);
or U3152 (N_3152,In_894,In_642);
nand U3153 (N_3153,In_952,In_832);
and U3154 (N_3154,In_1412,In_863);
nor U3155 (N_3155,In_142,In_927);
nand U3156 (N_3156,In_1123,In_301);
and U3157 (N_3157,In_1060,In_1368);
and U3158 (N_3158,In_287,In_584);
or U3159 (N_3159,In_621,In_558);
nor U3160 (N_3160,In_1325,In_694);
nand U3161 (N_3161,In_640,In_375);
and U3162 (N_3162,In_733,In_522);
nor U3163 (N_3163,In_1415,In_1399);
nand U3164 (N_3164,In_740,In_269);
or U3165 (N_3165,In_1423,In_1360);
nand U3166 (N_3166,In_1022,In_437);
nand U3167 (N_3167,In_841,In_1000);
nand U3168 (N_3168,In_1438,In_1480);
or U3169 (N_3169,In_137,In_734);
xnor U3170 (N_3170,In_1282,In_792);
xnor U3171 (N_3171,In_130,In_1249);
nand U3172 (N_3172,In_1237,In_123);
and U3173 (N_3173,In_678,In_312);
and U3174 (N_3174,In_1041,In_1229);
and U3175 (N_3175,In_199,In_1492);
and U3176 (N_3176,In_1490,In_1325);
xor U3177 (N_3177,In_691,In_1085);
or U3178 (N_3178,In_1030,In_1048);
nor U3179 (N_3179,In_620,In_1046);
nand U3180 (N_3180,In_32,In_704);
nor U3181 (N_3181,In_1177,In_46);
nor U3182 (N_3182,In_1271,In_1345);
or U3183 (N_3183,In_334,In_1385);
and U3184 (N_3184,In_1488,In_607);
or U3185 (N_3185,In_1261,In_886);
or U3186 (N_3186,In_310,In_220);
nor U3187 (N_3187,In_1417,In_1035);
and U3188 (N_3188,In_327,In_1190);
and U3189 (N_3189,In_116,In_766);
and U3190 (N_3190,In_608,In_1492);
nand U3191 (N_3191,In_524,In_527);
and U3192 (N_3192,In_768,In_1480);
and U3193 (N_3193,In_523,In_898);
nor U3194 (N_3194,In_1295,In_148);
nand U3195 (N_3195,In_307,In_351);
nor U3196 (N_3196,In_705,In_1163);
or U3197 (N_3197,In_294,In_1135);
and U3198 (N_3198,In_413,In_730);
nor U3199 (N_3199,In_159,In_297);
nor U3200 (N_3200,In_1190,In_1162);
or U3201 (N_3201,In_367,In_1197);
nand U3202 (N_3202,In_408,In_70);
and U3203 (N_3203,In_171,In_1022);
nand U3204 (N_3204,In_1339,In_494);
and U3205 (N_3205,In_11,In_24);
and U3206 (N_3206,In_597,In_944);
and U3207 (N_3207,In_106,In_213);
nand U3208 (N_3208,In_1493,In_715);
or U3209 (N_3209,In_105,In_115);
nor U3210 (N_3210,In_1410,In_388);
xnor U3211 (N_3211,In_112,In_1167);
xor U3212 (N_3212,In_124,In_1281);
nand U3213 (N_3213,In_974,In_915);
or U3214 (N_3214,In_317,In_1236);
nor U3215 (N_3215,In_523,In_152);
nor U3216 (N_3216,In_831,In_455);
xnor U3217 (N_3217,In_1262,In_466);
nor U3218 (N_3218,In_534,In_834);
or U3219 (N_3219,In_1165,In_648);
nand U3220 (N_3220,In_1046,In_1130);
nand U3221 (N_3221,In_815,In_1190);
nand U3222 (N_3222,In_251,In_925);
and U3223 (N_3223,In_423,In_1070);
nor U3224 (N_3224,In_1478,In_854);
nor U3225 (N_3225,In_395,In_828);
nand U3226 (N_3226,In_942,In_905);
nor U3227 (N_3227,In_945,In_1199);
nand U3228 (N_3228,In_780,In_295);
nor U3229 (N_3229,In_564,In_418);
nand U3230 (N_3230,In_127,In_833);
or U3231 (N_3231,In_937,In_1126);
or U3232 (N_3232,In_1221,In_181);
nor U3233 (N_3233,In_413,In_988);
nor U3234 (N_3234,In_1355,In_560);
nand U3235 (N_3235,In_130,In_738);
or U3236 (N_3236,In_283,In_272);
xnor U3237 (N_3237,In_1058,In_225);
xnor U3238 (N_3238,In_2,In_1193);
nand U3239 (N_3239,In_1302,In_1325);
or U3240 (N_3240,In_365,In_1061);
and U3241 (N_3241,In_350,In_401);
and U3242 (N_3242,In_1475,In_61);
xor U3243 (N_3243,In_385,In_68);
xnor U3244 (N_3244,In_1274,In_512);
xnor U3245 (N_3245,In_99,In_159);
and U3246 (N_3246,In_607,In_1021);
nor U3247 (N_3247,In_295,In_422);
xnor U3248 (N_3248,In_322,In_451);
nand U3249 (N_3249,In_1289,In_224);
nand U3250 (N_3250,In_575,In_815);
and U3251 (N_3251,In_1399,In_1044);
nor U3252 (N_3252,In_213,In_366);
nor U3253 (N_3253,In_329,In_1351);
and U3254 (N_3254,In_1342,In_1343);
or U3255 (N_3255,In_1405,In_596);
or U3256 (N_3256,In_1471,In_669);
or U3257 (N_3257,In_706,In_1418);
nand U3258 (N_3258,In_2,In_630);
nand U3259 (N_3259,In_145,In_700);
or U3260 (N_3260,In_491,In_822);
and U3261 (N_3261,In_914,In_1307);
and U3262 (N_3262,In_711,In_385);
nor U3263 (N_3263,In_1108,In_715);
xnor U3264 (N_3264,In_1120,In_285);
and U3265 (N_3265,In_460,In_503);
xor U3266 (N_3266,In_986,In_358);
nor U3267 (N_3267,In_1098,In_800);
and U3268 (N_3268,In_495,In_1026);
and U3269 (N_3269,In_638,In_1279);
xnor U3270 (N_3270,In_1154,In_780);
nand U3271 (N_3271,In_1168,In_903);
xnor U3272 (N_3272,In_336,In_321);
nand U3273 (N_3273,In_19,In_232);
nand U3274 (N_3274,In_713,In_1288);
and U3275 (N_3275,In_705,In_1078);
and U3276 (N_3276,In_949,In_645);
nand U3277 (N_3277,In_399,In_381);
or U3278 (N_3278,In_1071,In_609);
or U3279 (N_3279,In_604,In_1300);
nor U3280 (N_3280,In_294,In_748);
and U3281 (N_3281,In_655,In_1357);
nor U3282 (N_3282,In_911,In_353);
and U3283 (N_3283,In_453,In_855);
nand U3284 (N_3284,In_1158,In_212);
or U3285 (N_3285,In_557,In_1451);
and U3286 (N_3286,In_637,In_1430);
nand U3287 (N_3287,In_1136,In_1139);
and U3288 (N_3288,In_1156,In_1317);
nand U3289 (N_3289,In_59,In_169);
and U3290 (N_3290,In_1396,In_1459);
and U3291 (N_3291,In_414,In_109);
and U3292 (N_3292,In_771,In_818);
and U3293 (N_3293,In_266,In_285);
and U3294 (N_3294,In_1483,In_94);
nand U3295 (N_3295,In_709,In_933);
xor U3296 (N_3296,In_1368,In_407);
nor U3297 (N_3297,In_386,In_1045);
nor U3298 (N_3298,In_419,In_812);
or U3299 (N_3299,In_1056,In_830);
nand U3300 (N_3300,In_227,In_1158);
xor U3301 (N_3301,In_1175,In_1217);
or U3302 (N_3302,In_1003,In_1011);
nor U3303 (N_3303,In_1014,In_1067);
xnor U3304 (N_3304,In_1084,In_145);
xor U3305 (N_3305,In_1157,In_1118);
nand U3306 (N_3306,In_1003,In_849);
xor U3307 (N_3307,In_886,In_445);
nand U3308 (N_3308,In_748,In_1396);
nor U3309 (N_3309,In_741,In_1195);
or U3310 (N_3310,In_692,In_244);
xnor U3311 (N_3311,In_881,In_252);
and U3312 (N_3312,In_415,In_1267);
nand U3313 (N_3313,In_1210,In_1272);
or U3314 (N_3314,In_897,In_154);
or U3315 (N_3315,In_975,In_723);
nor U3316 (N_3316,In_598,In_1339);
nand U3317 (N_3317,In_389,In_980);
xnor U3318 (N_3318,In_1107,In_1389);
or U3319 (N_3319,In_1331,In_10);
or U3320 (N_3320,In_1201,In_363);
nand U3321 (N_3321,In_1364,In_431);
or U3322 (N_3322,In_1097,In_1489);
xnor U3323 (N_3323,In_800,In_94);
and U3324 (N_3324,In_1306,In_1185);
nor U3325 (N_3325,In_482,In_1200);
or U3326 (N_3326,In_934,In_1497);
nand U3327 (N_3327,In_1055,In_771);
or U3328 (N_3328,In_334,In_786);
nor U3329 (N_3329,In_21,In_311);
and U3330 (N_3330,In_1019,In_1008);
nor U3331 (N_3331,In_421,In_1375);
nand U3332 (N_3332,In_1210,In_503);
and U3333 (N_3333,In_1417,In_1324);
and U3334 (N_3334,In_664,In_334);
nand U3335 (N_3335,In_563,In_25);
nor U3336 (N_3336,In_977,In_263);
xor U3337 (N_3337,In_363,In_774);
nand U3338 (N_3338,In_451,In_1308);
xnor U3339 (N_3339,In_1038,In_684);
nand U3340 (N_3340,In_98,In_623);
or U3341 (N_3341,In_431,In_366);
and U3342 (N_3342,In_1381,In_624);
nand U3343 (N_3343,In_1313,In_540);
or U3344 (N_3344,In_681,In_1418);
or U3345 (N_3345,In_521,In_941);
nor U3346 (N_3346,In_275,In_404);
and U3347 (N_3347,In_1262,In_1258);
or U3348 (N_3348,In_1421,In_377);
or U3349 (N_3349,In_487,In_1204);
nand U3350 (N_3350,In_1493,In_153);
nand U3351 (N_3351,In_564,In_1241);
or U3352 (N_3352,In_973,In_550);
or U3353 (N_3353,In_892,In_575);
nand U3354 (N_3354,In_835,In_1384);
nand U3355 (N_3355,In_1415,In_1219);
nand U3356 (N_3356,In_1297,In_889);
nand U3357 (N_3357,In_1345,In_811);
nand U3358 (N_3358,In_1322,In_1242);
nor U3359 (N_3359,In_665,In_955);
nor U3360 (N_3360,In_1129,In_96);
and U3361 (N_3361,In_1362,In_1441);
xor U3362 (N_3362,In_523,In_534);
nand U3363 (N_3363,In_776,In_1282);
or U3364 (N_3364,In_879,In_151);
or U3365 (N_3365,In_1111,In_743);
nand U3366 (N_3366,In_515,In_955);
nor U3367 (N_3367,In_843,In_38);
nor U3368 (N_3368,In_518,In_254);
nor U3369 (N_3369,In_580,In_1010);
nand U3370 (N_3370,In_1097,In_1217);
nand U3371 (N_3371,In_931,In_508);
xnor U3372 (N_3372,In_1002,In_758);
nand U3373 (N_3373,In_8,In_922);
nor U3374 (N_3374,In_834,In_954);
nand U3375 (N_3375,In_910,In_157);
and U3376 (N_3376,In_1029,In_1348);
nor U3377 (N_3377,In_572,In_1300);
and U3378 (N_3378,In_344,In_622);
nand U3379 (N_3379,In_435,In_32);
nor U3380 (N_3380,In_135,In_1463);
or U3381 (N_3381,In_374,In_1065);
xnor U3382 (N_3382,In_286,In_1440);
nor U3383 (N_3383,In_1064,In_1446);
and U3384 (N_3384,In_332,In_1110);
or U3385 (N_3385,In_48,In_741);
or U3386 (N_3386,In_39,In_447);
nand U3387 (N_3387,In_1278,In_790);
and U3388 (N_3388,In_7,In_63);
and U3389 (N_3389,In_1143,In_241);
nand U3390 (N_3390,In_797,In_760);
or U3391 (N_3391,In_117,In_477);
or U3392 (N_3392,In_371,In_276);
or U3393 (N_3393,In_299,In_666);
nand U3394 (N_3394,In_328,In_994);
and U3395 (N_3395,In_408,In_893);
nand U3396 (N_3396,In_678,In_169);
nand U3397 (N_3397,In_142,In_820);
nand U3398 (N_3398,In_81,In_742);
or U3399 (N_3399,In_1361,In_998);
or U3400 (N_3400,In_215,In_610);
or U3401 (N_3401,In_297,In_1211);
nor U3402 (N_3402,In_893,In_1371);
or U3403 (N_3403,In_1364,In_1117);
or U3404 (N_3404,In_558,In_996);
nand U3405 (N_3405,In_1148,In_1019);
nor U3406 (N_3406,In_571,In_1263);
xnor U3407 (N_3407,In_1112,In_998);
and U3408 (N_3408,In_832,In_1168);
nor U3409 (N_3409,In_413,In_435);
or U3410 (N_3410,In_912,In_511);
nand U3411 (N_3411,In_441,In_865);
and U3412 (N_3412,In_112,In_525);
nor U3413 (N_3413,In_446,In_1104);
xnor U3414 (N_3414,In_434,In_1408);
and U3415 (N_3415,In_641,In_672);
and U3416 (N_3416,In_1247,In_1210);
and U3417 (N_3417,In_511,In_505);
nand U3418 (N_3418,In_401,In_1045);
xor U3419 (N_3419,In_83,In_717);
or U3420 (N_3420,In_615,In_905);
xnor U3421 (N_3421,In_291,In_717);
and U3422 (N_3422,In_403,In_1431);
and U3423 (N_3423,In_991,In_1156);
nand U3424 (N_3424,In_784,In_179);
xor U3425 (N_3425,In_436,In_1203);
nand U3426 (N_3426,In_975,In_578);
nor U3427 (N_3427,In_593,In_714);
or U3428 (N_3428,In_108,In_1259);
nor U3429 (N_3429,In_497,In_1274);
and U3430 (N_3430,In_1293,In_429);
nand U3431 (N_3431,In_1484,In_559);
nor U3432 (N_3432,In_993,In_1122);
nor U3433 (N_3433,In_623,In_945);
xnor U3434 (N_3434,In_989,In_173);
nand U3435 (N_3435,In_228,In_1001);
and U3436 (N_3436,In_904,In_1128);
nand U3437 (N_3437,In_455,In_925);
nor U3438 (N_3438,In_122,In_551);
nor U3439 (N_3439,In_1424,In_120);
and U3440 (N_3440,In_276,In_1080);
and U3441 (N_3441,In_621,In_1432);
or U3442 (N_3442,In_935,In_329);
and U3443 (N_3443,In_817,In_1456);
nand U3444 (N_3444,In_331,In_556);
and U3445 (N_3445,In_445,In_618);
and U3446 (N_3446,In_960,In_1051);
nor U3447 (N_3447,In_1268,In_819);
or U3448 (N_3448,In_512,In_882);
nand U3449 (N_3449,In_509,In_489);
and U3450 (N_3450,In_458,In_1382);
and U3451 (N_3451,In_813,In_73);
or U3452 (N_3452,In_986,In_286);
or U3453 (N_3453,In_964,In_1052);
and U3454 (N_3454,In_860,In_283);
and U3455 (N_3455,In_397,In_361);
and U3456 (N_3456,In_354,In_560);
nor U3457 (N_3457,In_43,In_1196);
nand U3458 (N_3458,In_1296,In_1024);
and U3459 (N_3459,In_655,In_938);
nand U3460 (N_3460,In_367,In_119);
or U3461 (N_3461,In_403,In_804);
nor U3462 (N_3462,In_1411,In_1320);
nor U3463 (N_3463,In_271,In_528);
nor U3464 (N_3464,In_458,In_110);
or U3465 (N_3465,In_326,In_808);
and U3466 (N_3466,In_1160,In_527);
nor U3467 (N_3467,In_516,In_864);
xor U3468 (N_3468,In_91,In_562);
or U3469 (N_3469,In_412,In_90);
xor U3470 (N_3470,In_999,In_652);
nor U3471 (N_3471,In_271,In_25);
nor U3472 (N_3472,In_231,In_128);
nor U3473 (N_3473,In_466,In_244);
nor U3474 (N_3474,In_700,In_1052);
or U3475 (N_3475,In_1077,In_707);
or U3476 (N_3476,In_1268,In_260);
nor U3477 (N_3477,In_968,In_1108);
and U3478 (N_3478,In_920,In_1256);
and U3479 (N_3479,In_659,In_1289);
or U3480 (N_3480,In_724,In_969);
xnor U3481 (N_3481,In_761,In_1158);
nand U3482 (N_3482,In_72,In_757);
nand U3483 (N_3483,In_406,In_524);
nor U3484 (N_3484,In_900,In_1159);
or U3485 (N_3485,In_1413,In_1202);
nand U3486 (N_3486,In_1166,In_1347);
and U3487 (N_3487,In_485,In_1078);
or U3488 (N_3488,In_799,In_875);
or U3489 (N_3489,In_864,In_777);
or U3490 (N_3490,In_821,In_352);
and U3491 (N_3491,In_982,In_954);
or U3492 (N_3492,In_106,In_1035);
and U3493 (N_3493,In_998,In_1274);
nand U3494 (N_3494,In_1406,In_436);
nand U3495 (N_3495,In_664,In_178);
and U3496 (N_3496,In_506,In_857);
and U3497 (N_3497,In_543,In_829);
nor U3498 (N_3498,In_772,In_24);
and U3499 (N_3499,In_779,In_681);
nand U3500 (N_3500,In_946,In_135);
and U3501 (N_3501,In_1136,In_847);
nand U3502 (N_3502,In_841,In_290);
nor U3503 (N_3503,In_233,In_225);
nor U3504 (N_3504,In_802,In_1282);
or U3505 (N_3505,In_557,In_952);
nor U3506 (N_3506,In_487,In_1425);
nor U3507 (N_3507,In_1244,In_1384);
and U3508 (N_3508,In_334,In_1185);
or U3509 (N_3509,In_568,In_334);
or U3510 (N_3510,In_163,In_206);
nand U3511 (N_3511,In_664,In_280);
and U3512 (N_3512,In_490,In_1064);
and U3513 (N_3513,In_467,In_1013);
nand U3514 (N_3514,In_954,In_354);
and U3515 (N_3515,In_1109,In_1394);
or U3516 (N_3516,In_812,In_1051);
or U3517 (N_3517,In_901,In_580);
and U3518 (N_3518,In_636,In_357);
and U3519 (N_3519,In_1360,In_1032);
or U3520 (N_3520,In_1477,In_253);
nand U3521 (N_3521,In_768,In_750);
nor U3522 (N_3522,In_190,In_367);
or U3523 (N_3523,In_1025,In_996);
or U3524 (N_3524,In_553,In_1354);
nor U3525 (N_3525,In_1292,In_52);
and U3526 (N_3526,In_692,In_752);
and U3527 (N_3527,In_1252,In_754);
and U3528 (N_3528,In_1283,In_392);
nand U3529 (N_3529,In_213,In_428);
xor U3530 (N_3530,In_1321,In_1090);
or U3531 (N_3531,In_710,In_335);
xnor U3532 (N_3532,In_107,In_661);
and U3533 (N_3533,In_433,In_264);
nor U3534 (N_3534,In_649,In_1385);
nor U3535 (N_3535,In_712,In_51);
nor U3536 (N_3536,In_131,In_247);
and U3537 (N_3537,In_47,In_1442);
nand U3538 (N_3538,In_36,In_316);
and U3539 (N_3539,In_889,In_1196);
and U3540 (N_3540,In_463,In_720);
nor U3541 (N_3541,In_782,In_975);
nor U3542 (N_3542,In_230,In_706);
nor U3543 (N_3543,In_1168,In_711);
and U3544 (N_3544,In_560,In_78);
or U3545 (N_3545,In_29,In_1419);
nor U3546 (N_3546,In_314,In_1340);
nand U3547 (N_3547,In_309,In_1112);
nor U3548 (N_3548,In_673,In_160);
or U3549 (N_3549,In_207,In_304);
or U3550 (N_3550,In_1399,In_1333);
nand U3551 (N_3551,In_380,In_1141);
nor U3552 (N_3552,In_1253,In_475);
and U3553 (N_3553,In_370,In_1206);
nor U3554 (N_3554,In_878,In_706);
nand U3555 (N_3555,In_109,In_1200);
nor U3556 (N_3556,In_324,In_167);
or U3557 (N_3557,In_994,In_146);
or U3558 (N_3558,In_819,In_473);
nor U3559 (N_3559,In_910,In_552);
nor U3560 (N_3560,In_906,In_1119);
and U3561 (N_3561,In_81,In_390);
and U3562 (N_3562,In_1087,In_295);
nor U3563 (N_3563,In_1287,In_1165);
and U3564 (N_3564,In_1209,In_1055);
nand U3565 (N_3565,In_288,In_764);
and U3566 (N_3566,In_204,In_1319);
nand U3567 (N_3567,In_366,In_354);
and U3568 (N_3568,In_1005,In_1444);
and U3569 (N_3569,In_614,In_1480);
nand U3570 (N_3570,In_831,In_397);
or U3571 (N_3571,In_590,In_344);
nand U3572 (N_3572,In_1493,In_1259);
nor U3573 (N_3573,In_732,In_683);
and U3574 (N_3574,In_868,In_599);
or U3575 (N_3575,In_531,In_1491);
nand U3576 (N_3576,In_696,In_604);
nor U3577 (N_3577,In_46,In_1470);
xor U3578 (N_3578,In_1030,In_1436);
nor U3579 (N_3579,In_617,In_689);
xnor U3580 (N_3580,In_965,In_414);
nand U3581 (N_3581,In_1108,In_1259);
nor U3582 (N_3582,In_1162,In_226);
nor U3583 (N_3583,In_377,In_257);
or U3584 (N_3584,In_1143,In_1492);
or U3585 (N_3585,In_1143,In_771);
or U3586 (N_3586,In_452,In_511);
and U3587 (N_3587,In_851,In_1451);
nand U3588 (N_3588,In_346,In_1201);
and U3589 (N_3589,In_251,In_368);
xnor U3590 (N_3590,In_1239,In_1348);
and U3591 (N_3591,In_1327,In_273);
nor U3592 (N_3592,In_805,In_52);
or U3593 (N_3593,In_972,In_1090);
or U3594 (N_3594,In_1284,In_764);
and U3595 (N_3595,In_681,In_956);
xor U3596 (N_3596,In_1264,In_541);
and U3597 (N_3597,In_316,In_199);
and U3598 (N_3598,In_1168,In_1112);
nand U3599 (N_3599,In_466,In_1264);
and U3600 (N_3600,In_1230,In_539);
or U3601 (N_3601,In_229,In_818);
nand U3602 (N_3602,In_1304,In_892);
nand U3603 (N_3603,In_455,In_536);
nor U3604 (N_3604,In_1,In_1358);
nor U3605 (N_3605,In_202,In_504);
xor U3606 (N_3606,In_718,In_15);
or U3607 (N_3607,In_70,In_258);
nor U3608 (N_3608,In_835,In_212);
or U3609 (N_3609,In_1483,In_1367);
and U3610 (N_3610,In_385,In_674);
or U3611 (N_3611,In_392,In_316);
nor U3612 (N_3612,In_1007,In_1331);
nor U3613 (N_3613,In_287,In_382);
or U3614 (N_3614,In_1043,In_861);
and U3615 (N_3615,In_589,In_1486);
or U3616 (N_3616,In_898,In_1424);
nand U3617 (N_3617,In_458,In_1118);
xnor U3618 (N_3618,In_223,In_984);
nand U3619 (N_3619,In_155,In_96);
nand U3620 (N_3620,In_456,In_893);
or U3621 (N_3621,In_1077,In_1237);
nand U3622 (N_3622,In_161,In_459);
nand U3623 (N_3623,In_1113,In_1401);
nand U3624 (N_3624,In_382,In_782);
and U3625 (N_3625,In_1189,In_202);
nand U3626 (N_3626,In_447,In_1081);
nand U3627 (N_3627,In_972,In_1020);
xor U3628 (N_3628,In_294,In_179);
nor U3629 (N_3629,In_835,In_1257);
or U3630 (N_3630,In_1198,In_565);
xor U3631 (N_3631,In_867,In_609);
xor U3632 (N_3632,In_162,In_832);
nand U3633 (N_3633,In_941,In_1205);
or U3634 (N_3634,In_637,In_1025);
or U3635 (N_3635,In_876,In_148);
nand U3636 (N_3636,In_689,In_933);
and U3637 (N_3637,In_1178,In_320);
nand U3638 (N_3638,In_899,In_448);
nor U3639 (N_3639,In_957,In_1153);
and U3640 (N_3640,In_1284,In_1358);
and U3641 (N_3641,In_697,In_1397);
and U3642 (N_3642,In_661,In_924);
nor U3643 (N_3643,In_1212,In_1048);
and U3644 (N_3644,In_1016,In_547);
and U3645 (N_3645,In_889,In_550);
or U3646 (N_3646,In_346,In_380);
nand U3647 (N_3647,In_1261,In_189);
and U3648 (N_3648,In_262,In_779);
and U3649 (N_3649,In_602,In_1392);
or U3650 (N_3650,In_223,In_822);
or U3651 (N_3651,In_193,In_202);
and U3652 (N_3652,In_1149,In_982);
xor U3653 (N_3653,In_926,In_932);
and U3654 (N_3654,In_1318,In_1004);
and U3655 (N_3655,In_457,In_7);
and U3656 (N_3656,In_93,In_1121);
or U3657 (N_3657,In_594,In_392);
nand U3658 (N_3658,In_1203,In_1394);
nand U3659 (N_3659,In_601,In_841);
and U3660 (N_3660,In_877,In_813);
nor U3661 (N_3661,In_412,In_1053);
and U3662 (N_3662,In_742,In_9);
and U3663 (N_3663,In_1273,In_1122);
nor U3664 (N_3664,In_218,In_893);
nor U3665 (N_3665,In_36,In_901);
and U3666 (N_3666,In_852,In_1338);
and U3667 (N_3667,In_684,In_335);
nor U3668 (N_3668,In_491,In_840);
nor U3669 (N_3669,In_119,In_1298);
or U3670 (N_3670,In_161,In_896);
nor U3671 (N_3671,In_1442,In_1435);
xnor U3672 (N_3672,In_1140,In_1498);
xnor U3673 (N_3673,In_616,In_949);
xor U3674 (N_3674,In_688,In_354);
or U3675 (N_3675,In_501,In_1476);
nor U3676 (N_3676,In_1406,In_1278);
nand U3677 (N_3677,In_622,In_61);
and U3678 (N_3678,In_1031,In_1343);
nand U3679 (N_3679,In_57,In_56);
nand U3680 (N_3680,In_853,In_1129);
xnor U3681 (N_3681,In_450,In_1143);
nor U3682 (N_3682,In_319,In_600);
nand U3683 (N_3683,In_384,In_712);
xnor U3684 (N_3684,In_817,In_406);
nand U3685 (N_3685,In_259,In_1370);
nor U3686 (N_3686,In_1306,In_120);
or U3687 (N_3687,In_1454,In_839);
and U3688 (N_3688,In_715,In_23);
and U3689 (N_3689,In_856,In_936);
or U3690 (N_3690,In_1184,In_390);
and U3691 (N_3691,In_1279,In_1264);
and U3692 (N_3692,In_792,In_1389);
or U3693 (N_3693,In_1151,In_1203);
or U3694 (N_3694,In_783,In_1033);
nand U3695 (N_3695,In_542,In_148);
and U3696 (N_3696,In_1055,In_685);
xor U3697 (N_3697,In_105,In_1193);
nor U3698 (N_3698,In_722,In_1329);
nor U3699 (N_3699,In_85,In_1189);
xor U3700 (N_3700,In_637,In_124);
nor U3701 (N_3701,In_868,In_115);
and U3702 (N_3702,In_1189,In_1235);
nor U3703 (N_3703,In_717,In_1383);
or U3704 (N_3704,In_668,In_549);
nor U3705 (N_3705,In_350,In_135);
nand U3706 (N_3706,In_658,In_914);
nand U3707 (N_3707,In_580,In_828);
nor U3708 (N_3708,In_1345,In_321);
and U3709 (N_3709,In_174,In_1094);
or U3710 (N_3710,In_851,In_668);
nand U3711 (N_3711,In_1478,In_508);
or U3712 (N_3712,In_1402,In_1004);
nor U3713 (N_3713,In_888,In_1304);
or U3714 (N_3714,In_1423,In_1345);
or U3715 (N_3715,In_1252,In_0);
and U3716 (N_3716,In_613,In_1266);
nand U3717 (N_3717,In_646,In_669);
nand U3718 (N_3718,In_607,In_230);
or U3719 (N_3719,In_1355,In_502);
or U3720 (N_3720,In_1456,In_1472);
or U3721 (N_3721,In_591,In_344);
xor U3722 (N_3722,In_411,In_489);
or U3723 (N_3723,In_764,In_1050);
nor U3724 (N_3724,In_159,In_769);
and U3725 (N_3725,In_213,In_923);
nand U3726 (N_3726,In_479,In_1391);
nor U3727 (N_3727,In_815,In_1012);
nand U3728 (N_3728,In_806,In_266);
or U3729 (N_3729,In_446,In_808);
xor U3730 (N_3730,In_875,In_411);
nor U3731 (N_3731,In_557,In_1434);
xor U3732 (N_3732,In_71,In_497);
nor U3733 (N_3733,In_1408,In_797);
xor U3734 (N_3734,In_567,In_370);
and U3735 (N_3735,In_1115,In_1328);
or U3736 (N_3736,In_1343,In_490);
and U3737 (N_3737,In_588,In_1391);
and U3738 (N_3738,In_772,In_265);
nor U3739 (N_3739,In_896,In_831);
and U3740 (N_3740,In_865,In_1289);
and U3741 (N_3741,In_250,In_1079);
nor U3742 (N_3742,In_1147,In_400);
or U3743 (N_3743,In_483,In_1321);
nand U3744 (N_3744,In_962,In_343);
or U3745 (N_3745,In_854,In_1359);
xnor U3746 (N_3746,In_571,In_1307);
and U3747 (N_3747,In_150,In_189);
xor U3748 (N_3748,In_471,In_885);
nor U3749 (N_3749,In_1236,In_1209);
nand U3750 (N_3750,In_1261,In_742);
or U3751 (N_3751,In_488,In_344);
nor U3752 (N_3752,In_1197,In_469);
or U3753 (N_3753,In_954,In_346);
nor U3754 (N_3754,In_1057,In_478);
or U3755 (N_3755,In_1401,In_1160);
nand U3756 (N_3756,In_929,In_1395);
xor U3757 (N_3757,In_1212,In_508);
nor U3758 (N_3758,In_1106,In_571);
or U3759 (N_3759,In_1060,In_54);
nor U3760 (N_3760,In_517,In_636);
nor U3761 (N_3761,In_1038,In_565);
nand U3762 (N_3762,In_607,In_35);
nor U3763 (N_3763,In_583,In_1112);
or U3764 (N_3764,In_1407,In_1131);
nand U3765 (N_3765,In_947,In_1441);
xor U3766 (N_3766,In_421,In_710);
nand U3767 (N_3767,In_702,In_223);
and U3768 (N_3768,In_499,In_600);
nor U3769 (N_3769,In_636,In_1291);
and U3770 (N_3770,In_557,In_1494);
nor U3771 (N_3771,In_371,In_1123);
xor U3772 (N_3772,In_791,In_609);
or U3773 (N_3773,In_758,In_1023);
or U3774 (N_3774,In_1378,In_1418);
nor U3775 (N_3775,In_331,In_458);
nor U3776 (N_3776,In_343,In_272);
nor U3777 (N_3777,In_882,In_793);
nand U3778 (N_3778,In_482,In_526);
xnor U3779 (N_3779,In_389,In_877);
or U3780 (N_3780,In_552,In_4);
or U3781 (N_3781,In_510,In_779);
nand U3782 (N_3782,In_27,In_818);
or U3783 (N_3783,In_1014,In_257);
and U3784 (N_3784,In_126,In_752);
nand U3785 (N_3785,In_654,In_509);
nand U3786 (N_3786,In_1330,In_598);
nand U3787 (N_3787,In_435,In_1251);
nor U3788 (N_3788,In_477,In_797);
nor U3789 (N_3789,In_1136,In_701);
nor U3790 (N_3790,In_1455,In_260);
nor U3791 (N_3791,In_1259,In_81);
nand U3792 (N_3792,In_1452,In_175);
or U3793 (N_3793,In_31,In_1299);
nor U3794 (N_3794,In_732,In_1239);
nor U3795 (N_3795,In_850,In_63);
or U3796 (N_3796,In_1028,In_1124);
xnor U3797 (N_3797,In_883,In_21);
nor U3798 (N_3798,In_466,In_599);
xnor U3799 (N_3799,In_265,In_1018);
or U3800 (N_3800,In_655,In_1204);
and U3801 (N_3801,In_746,In_653);
nand U3802 (N_3802,In_880,In_1123);
and U3803 (N_3803,In_1284,In_995);
nand U3804 (N_3804,In_578,In_1166);
nand U3805 (N_3805,In_1025,In_788);
nor U3806 (N_3806,In_1360,In_248);
and U3807 (N_3807,In_94,In_24);
nand U3808 (N_3808,In_912,In_251);
and U3809 (N_3809,In_1057,In_653);
nor U3810 (N_3810,In_825,In_888);
and U3811 (N_3811,In_775,In_1336);
nand U3812 (N_3812,In_305,In_1321);
nor U3813 (N_3813,In_466,In_1001);
or U3814 (N_3814,In_383,In_1478);
or U3815 (N_3815,In_506,In_765);
and U3816 (N_3816,In_633,In_1319);
and U3817 (N_3817,In_68,In_1094);
nand U3818 (N_3818,In_1280,In_1493);
and U3819 (N_3819,In_1221,In_667);
nand U3820 (N_3820,In_904,In_186);
nor U3821 (N_3821,In_429,In_240);
nand U3822 (N_3822,In_495,In_701);
xnor U3823 (N_3823,In_1446,In_1380);
and U3824 (N_3824,In_1205,In_500);
nor U3825 (N_3825,In_1425,In_635);
xor U3826 (N_3826,In_1128,In_1005);
and U3827 (N_3827,In_998,In_1406);
nor U3828 (N_3828,In_201,In_530);
nand U3829 (N_3829,In_1042,In_1294);
nor U3830 (N_3830,In_1030,In_1271);
nor U3831 (N_3831,In_117,In_880);
nand U3832 (N_3832,In_823,In_284);
xnor U3833 (N_3833,In_386,In_954);
and U3834 (N_3834,In_1013,In_86);
and U3835 (N_3835,In_330,In_601);
nand U3836 (N_3836,In_988,In_1195);
and U3837 (N_3837,In_956,In_646);
and U3838 (N_3838,In_77,In_460);
nor U3839 (N_3839,In_974,In_1491);
nor U3840 (N_3840,In_1300,In_1125);
nor U3841 (N_3841,In_1245,In_336);
or U3842 (N_3842,In_1463,In_1150);
nor U3843 (N_3843,In_1218,In_1340);
nor U3844 (N_3844,In_633,In_930);
or U3845 (N_3845,In_898,In_407);
nand U3846 (N_3846,In_1087,In_454);
nor U3847 (N_3847,In_13,In_1208);
nand U3848 (N_3848,In_474,In_1163);
nand U3849 (N_3849,In_1335,In_738);
nand U3850 (N_3850,In_218,In_1272);
and U3851 (N_3851,In_1466,In_1057);
nor U3852 (N_3852,In_1334,In_840);
nor U3853 (N_3853,In_553,In_274);
and U3854 (N_3854,In_622,In_623);
nand U3855 (N_3855,In_360,In_268);
nor U3856 (N_3856,In_806,In_642);
nand U3857 (N_3857,In_248,In_1379);
nor U3858 (N_3858,In_520,In_1370);
and U3859 (N_3859,In_1361,In_893);
nor U3860 (N_3860,In_1015,In_1292);
and U3861 (N_3861,In_950,In_675);
nand U3862 (N_3862,In_117,In_204);
nand U3863 (N_3863,In_1000,In_280);
nor U3864 (N_3864,In_1088,In_603);
xor U3865 (N_3865,In_482,In_966);
nor U3866 (N_3866,In_904,In_756);
nor U3867 (N_3867,In_819,In_0);
nor U3868 (N_3868,In_1035,In_1099);
or U3869 (N_3869,In_716,In_432);
xnor U3870 (N_3870,In_1224,In_213);
xnor U3871 (N_3871,In_1454,In_1442);
nor U3872 (N_3872,In_643,In_406);
nor U3873 (N_3873,In_968,In_298);
nand U3874 (N_3874,In_819,In_771);
xnor U3875 (N_3875,In_11,In_1441);
nor U3876 (N_3876,In_1277,In_18);
nor U3877 (N_3877,In_377,In_450);
or U3878 (N_3878,In_791,In_383);
xnor U3879 (N_3879,In_680,In_1280);
xor U3880 (N_3880,In_288,In_1015);
nor U3881 (N_3881,In_462,In_406);
nand U3882 (N_3882,In_1427,In_880);
nand U3883 (N_3883,In_912,In_750);
nand U3884 (N_3884,In_514,In_614);
nand U3885 (N_3885,In_1307,In_1420);
nand U3886 (N_3886,In_1462,In_952);
nand U3887 (N_3887,In_25,In_638);
or U3888 (N_3888,In_1405,In_1403);
and U3889 (N_3889,In_156,In_654);
and U3890 (N_3890,In_1162,In_1389);
nand U3891 (N_3891,In_766,In_341);
nand U3892 (N_3892,In_311,In_340);
nor U3893 (N_3893,In_802,In_654);
nor U3894 (N_3894,In_487,In_736);
nand U3895 (N_3895,In_1477,In_172);
nand U3896 (N_3896,In_1093,In_1202);
xnor U3897 (N_3897,In_44,In_226);
nor U3898 (N_3898,In_86,In_553);
and U3899 (N_3899,In_1345,In_1112);
xor U3900 (N_3900,In_972,In_787);
or U3901 (N_3901,In_576,In_504);
or U3902 (N_3902,In_647,In_39);
or U3903 (N_3903,In_572,In_141);
and U3904 (N_3904,In_74,In_763);
or U3905 (N_3905,In_969,In_232);
and U3906 (N_3906,In_1250,In_1126);
or U3907 (N_3907,In_954,In_457);
or U3908 (N_3908,In_1360,In_229);
nand U3909 (N_3909,In_364,In_670);
and U3910 (N_3910,In_2,In_244);
or U3911 (N_3911,In_1170,In_948);
and U3912 (N_3912,In_892,In_819);
xor U3913 (N_3913,In_1391,In_1077);
nand U3914 (N_3914,In_197,In_598);
or U3915 (N_3915,In_1004,In_112);
and U3916 (N_3916,In_587,In_51);
nor U3917 (N_3917,In_948,In_729);
and U3918 (N_3918,In_338,In_631);
nand U3919 (N_3919,In_1139,In_178);
or U3920 (N_3920,In_571,In_624);
nand U3921 (N_3921,In_594,In_283);
nand U3922 (N_3922,In_80,In_1058);
or U3923 (N_3923,In_583,In_1343);
or U3924 (N_3924,In_863,In_1116);
or U3925 (N_3925,In_461,In_242);
and U3926 (N_3926,In_659,In_266);
nor U3927 (N_3927,In_1124,In_628);
xor U3928 (N_3928,In_197,In_405);
nor U3929 (N_3929,In_329,In_511);
or U3930 (N_3930,In_738,In_91);
nor U3931 (N_3931,In_445,In_530);
or U3932 (N_3932,In_1142,In_499);
nand U3933 (N_3933,In_1359,In_1490);
and U3934 (N_3934,In_827,In_682);
nand U3935 (N_3935,In_1065,In_525);
or U3936 (N_3936,In_575,In_150);
nor U3937 (N_3937,In_953,In_856);
nand U3938 (N_3938,In_119,In_867);
nand U3939 (N_3939,In_1145,In_23);
nor U3940 (N_3940,In_519,In_1103);
or U3941 (N_3941,In_264,In_521);
and U3942 (N_3942,In_1218,In_1167);
and U3943 (N_3943,In_1171,In_1321);
xnor U3944 (N_3944,In_735,In_1336);
nor U3945 (N_3945,In_1196,In_648);
nor U3946 (N_3946,In_716,In_262);
nand U3947 (N_3947,In_258,In_886);
and U3948 (N_3948,In_409,In_699);
and U3949 (N_3949,In_578,In_1330);
nand U3950 (N_3950,In_1126,In_1444);
and U3951 (N_3951,In_347,In_75);
or U3952 (N_3952,In_1006,In_730);
and U3953 (N_3953,In_1422,In_187);
nor U3954 (N_3954,In_92,In_292);
or U3955 (N_3955,In_199,In_612);
nor U3956 (N_3956,In_1479,In_961);
and U3957 (N_3957,In_624,In_750);
nand U3958 (N_3958,In_916,In_1175);
nor U3959 (N_3959,In_531,In_175);
nor U3960 (N_3960,In_1344,In_1220);
nand U3961 (N_3961,In_593,In_980);
or U3962 (N_3962,In_1359,In_1066);
xnor U3963 (N_3963,In_1034,In_926);
and U3964 (N_3964,In_415,In_133);
and U3965 (N_3965,In_708,In_55);
and U3966 (N_3966,In_1373,In_602);
and U3967 (N_3967,In_1166,In_288);
and U3968 (N_3968,In_513,In_416);
and U3969 (N_3969,In_597,In_48);
xor U3970 (N_3970,In_1008,In_1174);
nand U3971 (N_3971,In_183,In_843);
xnor U3972 (N_3972,In_1118,In_883);
and U3973 (N_3973,In_837,In_136);
nor U3974 (N_3974,In_917,In_332);
and U3975 (N_3975,In_892,In_170);
nand U3976 (N_3976,In_366,In_151);
xnor U3977 (N_3977,In_69,In_905);
xor U3978 (N_3978,In_432,In_140);
or U3979 (N_3979,In_575,In_476);
and U3980 (N_3980,In_427,In_1039);
or U3981 (N_3981,In_399,In_894);
nand U3982 (N_3982,In_676,In_402);
nand U3983 (N_3983,In_799,In_1219);
and U3984 (N_3984,In_836,In_1031);
nand U3985 (N_3985,In_353,In_883);
and U3986 (N_3986,In_1118,In_942);
and U3987 (N_3987,In_1103,In_885);
xor U3988 (N_3988,In_518,In_299);
and U3989 (N_3989,In_391,In_1457);
nor U3990 (N_3990,In_1160,In_815);
or U3991 (N_3991,In_1470,In_1460);
or U3992 (N_3992,In_373,In_741);
nor U3993 (N_3993,In_455,In_1024);
and U3994 (N_3994,In_810,In_958);
nand U3995 (N_3995,In_436,In_866);
nand U3996 (N_3996,In_68,In_60);
and U3997 (N_3997,In_918,In_71);
or U3998 (N_3998,In_399,In_1453);
and U3999 (N_3999,In_400,In_960);
nand U4000 (N_4000,In_46,In_1016);
or U4001 (N_4001,In_464,In_67);
and U4002 (N_4002,In_1001,In_163);
xor U4003 (N_4003,In_888,In_409);
or U4004 (N_4004,In_1461,In_281);
nor U4005 (N_4005,In_274,In_1204);
and U4006 (N_4006,In_697,In_1410);
and U4007 (N_4007,In_563,In_975);
xor U4008 (N_4008,In_789,In_497);
and U4009 (N_4009,In_33,In_178);
or U4010 (N_4010,In_143,In_167);
or U4011 (N_4011,In_1151,In_851);
nor U4012 (N_4012,In_298,In_886);
nor U4013 (N_4013,In_451,In_749);
and U4014 (N_4014,In_625,In_663);
xnor U4015 (N_4015,In_53,In_34);
or U4016 (N_4016,In_1413,In_639);
nand U4017 (N_4017,In_291,In_964);
and U4018 (N_4018,In_330,In_798);
xnor U4019 (N_4019,In_848,In_368);
and U4020 (N_4020,In_1101,In_1279);
or U4021 (N_4021,In_727,In_807);
xnor U4022 (N_4022,In_1213,In_634);
and U4023 (N_4023,In_37,In_581);
and U4024 (N_4024,In_236,In_1416);
and U4025 (N_4025,In_1262,In_967);
nor U4026 (N_4026,In_858,In_1006);
or U4027 (N_4027,In_335,In_1038);
nor U4028 (N_4028,In_576,In_1334);
and U4029 (N_4029,In_953,In_505);
or U4030 (N_4030,In_547,In_231);
or U4031 (N_4031,In_39,In_903);
and U4032 (N_4032,In_68,In_353);
and U4033 (N_4033,In_220,In_841);
and U4034 (N_4034,In_137,In_568);
or U4035 (N_4035,In_986,In_461);
and U4036 (N_4036,In_369,In_184);
xnor U4037 (N_4037,In_1188,In_1227);
nor U4038 (N_4038,In_320,In_963);
or U4039 (N_4039,In_434,In_1209);
nor U4040 (N_4040,In_154,In_871);
and U4041 (N_4041,In_950,In_1058);
nand U4042 (N_4042,In_941,In_513);
xor U4043 (N_4043,In_776,In_75);
or U4044 (N_4044,In_87,In_51);
nor U4045 (N_4045,In_642,In_937);
nor U4046 (N_4046,In_814,In_428);
nand U4047 (N_4047,In_315,In_195);
and U4048 (N_4048,In_883,In_1093);
nor U4049 (N_4049,In_687,In_1260);
and U4050 (N_4050,In_1077,In_1379);
nand U4051 (N_4051,In_1490,In_1413);
nand U4052 (N_4052,In_581,In_294);
and U4053 (N_4053,In_1154,In_1495);
or U4054 (N_4054,In_859,In_1195);
nand U4055 (N_4055,In_917,In_528);
and U4056 (N_4056,In_379,In_781);
and U4057 (N_4057,In_60,In_187);
or U4058 (N_4058,In_1024,In_109);
nor U4059 (N_4059,In_973,In_571);
xor U4060 (N_4060,In_1441,In_428);
nor U4061 (N_4061,In_1218,In_1307);
or U4062 (N_4062,In_1106,In_244);
nor U4063 (N_4063,In_380,In_191);
nand U4064 (N_4064,In_110,In_776);
or U4065 (N_4065,In_237,In_211);
and U4066 (N_4066,In_1397,In_512);
nand U4067 (N_4067,In_1414,In_1057);
or U4068 (N_4068,In_769,In_503);
and U4069 (N_4069,In_329,In_358);
nor U4070 (N_4070,In_663,In_113);
nand U4071 (N_4071,In_295,In_261);
xnor U4072 (N_4072,In_1269,In_1346);
xnor U4073 (N_4073,In_1141,In_182);
nand U4074 (N_4074,In_1350,In_1040);
nand U4075 (N_4075,In_1366,In_614);
xnor U4076 (N_4076,In_1420,In_971);
or U4077 (N_4077,In_17,In_366);
nand U4078 (N_4078,In_330,In_286);
nand U4079 (N_4079,In_334,In_942);
and U4080 (N_4080,In_973,In_53);
xnor U4081 (N_4081,In_1219,In_1272);
nor U4082 (N_4082,In_638,In_497);
nor U4083 (N_4083,In_1411,In_459);
nor U4084 (N_4084,In_252,In_937);
or U4085 (N_4085,In_1158,In_461);
and U4086 (N_4086,In_1169,In_607);
xor U4087 (N_4087,In_912,In_1191);
nand U4088 (N_4088,In_16,In_1465);
nand U4089 (N_4089,In_846,In_956);
nor U4090 (N_4090,In_1008,In_213);
nor U4091 (N_4091,In_477,In_962);
nand U4092 (N_4092,In_781,In_1013);
nand U4093 (N_4093,In_349,In_725);
and U4094 (N_4094,In_731,In_859);
or U4095 (N_4095,In_585,In_522);
nor U4096 (N_4096,In_669,In_710);
nand U4097 (N_4097,In_443,In_174);
nor U4098 (N_4098,In_1286,In_709);
or U4099 (N_4099,In_1108,In_1218);
nand U4100 (N_4100,In_125,In_1308);
and U4101 (N_4101,In_997,In_960);
and U4102 (N_4102,In_659,In_353);
nor U4103 (N_4103,In_918,In_187);
or U4104 (N_4104,In_1223,In_502);
nor U4105 (N_4105,In_1226,In_1182);
and U4106 (N_4106,In_549,In_1032);
xnor U4107 (N_4107,In_157,In_394);
nor U4108 (N_4108,In_787,In_193);
nor U4109 (N_4109,In_1197,In_622);
and U4110 (N_4110,In_379,In_438);
xor U4111 (N_4111,In_538,In_389);
or U4112 (N_4112,In_1221,In_955);
nor U4113 (N_4113,In_254,In_523);
nand U4114 (N_4114,In_706,In_614);
nor U4115 (N_4115,In_187,In_955);
nand U4116 (N_4116,In_788,In_686);
nand U4117 (N_4117,In_15,In_305);
and U4118 (N_4118,In_944,In_1478);
nor U4119 (N_4119,In_404,In_504);
or U4120 (N_4120,In_1111,In_10);
nor U4121 (N_4121,In_1473,In_522);
nand U4122 (N_4122,In_123,In_1097);
and U4123 (N_4123,In_50,In_539);
and U4124 (N_4124,In_567,In_172);
xnor U4125 (N_4125,In_758,In_691);
or U4126 (N_4126,In_57,In_1340);
and U4127 (N_4127,In_1342,In_925);
nand U4128 (N_4128,In_474,In_546);
and U4129 (N_4129,In_890,In_228);
or U4130 (N_4130,In_722,In_898);
nor U4131 (N_4131,In_473,In_776);
nand U4132 (N_4132,In_622,In_825);
and U4133 (N_4133,In_1169,In_263);
nor U4134 (N_4134,In_1465,In_793);
and U4135 (N_4135,In_87,In_1170);
or U4136 (N_4136,In_1,In_820);
nor U4137 (N_4137,In_640,In_1058);
nor U4138 (N_4138,In_131,In_569);
or U4139 (N_4139,In_66,In_474);
or U4140 (N_4140,In_127,In_426);
and U4141 (N_4141,In_1008,In_169);
nand U4142 (N_4142,In_248,In_140);
or U4143 (N_4143,In_1012,In_411);
and U4144 (N_4144,In_584,In_66);
nand U4145 (N_4145,In_306,In_663);
nor U4146 (N_4146,In_1314,In_940);
or U4147 (N_4147,In_693,In_1483);
nand U4148 (N_4148,In_1349,In_1371);
xor U4149 (N_4149,In_266,In_624);
or U4150 (N_4150,In_1037,In_939);
or U4151 (N_4151,In_881,In_1312);
nor U4152 (N_4152,In_394,In_1341);
nand U4153 (N_4153,In_911,In_124);
or U4154 (N_4154,In_1232,In_1255);
nor U4155 (N_4155,In_1443,In_710);
nor U4156 (N_4156,In_486,In_897);
or U4157 (N_4157,In_388,In_1142);
nand U4158 (N_4158,In_137,In_333);
and U4159 (N_4159,In_675,In_1027);
nor U4160 (N_4160,In_1292,In_684);
nor U4161 (N_4161,In_1370,In_1061);
nor U4162 (N_4162,In_1420,In_575);
nand U4163 (N_4163,In_1256,In_46);
xnor U4164 (N_4164,In_745,In_564);
nand U4165 (N_4165,In_1185,In_907);
and U4166 (N_4166,In_1393,In_1283);
nand U4167 (N_4167,In_176,In_1332);
or U4168 (N_4168,In_269,In_123);
nor U4169 (N_4169,In_1417,In_35);
or U4170 (N_4170,In_855,In_608);
and U4171 (N_4171,In_732,In_1434);
xnor U4172 (N_4172,In_554,In_838);
or U4173 (N_4173,In_928,In_1370);
nand U4174 (N_4174,In_1172,In_1235);
or U4175 (N_4175,In_640,In_875);
nand U4176 (N_4176,In_609,In_1114);
nor U4177 (N_4177,In_35,In_1086);
nand U4178 (N_4178,In_289,In_1075);
or U4179 (N_4179,In_153,In_100);
nor U4180 (N_4180,In_693,In_844);
or U4181 (N_4181,In_230,In_158);
or U4182 (N_4182,In_146,In_858);
nand U4183 (N_4183,In_608,In_327);
and U4184 (N_4184,In_775,In_393);
or U4185 (N_4185,In_937,In_567);
nor U4186 (N_4186,In_492,In_1204);
and U4187 (N_4187,In_1064,In_817);
nor U4188 (N_4188,In_405,In_1405);
or U4189 (N_4189,In_1286,In_765);
nand U4190 (N_4190,In_927,In_475);
or U4191 (N_4191,In_804,In_555);
nor U4192 (N_4192,In_1307,In_1237);
or U4193 (N_4193,In_271,In_1178);
and U4194 (N_4194,In_1246,In_620);
and U4195 (N_4195,In_1252,In_322);
nand U4196 (N_4196,In_770,In_693);
nand U4197 (N_4197,In_1099,In_1388);
and U4198 (N_4198,In_1176,In_802);
and U4199 (N_4199,In_1466,In_1038);
and U4200 (N_4200,In_1019,In_350);
or U4201 (N_4201,In_1302,In_754);
and U4202 (N_4202,In_1460,In_633);
or U4203 (N_4203,In_614,In_1446);
and U4204 (N_4204,In_584,In_750);
or U4205 (N_4205,In_1142,In_601);
nand U4206 (N_4206,In_82,In_895);
and U4207 (N_4207,In_353,In_1061);
nand U4208 (N_4208,In_23,In_161);
and U4209 (N_4209,In_1394,In_502);
nor U4210 (N_4210,In_1105,In_390);
or U4211 (N_4211,In_329,In_857);
nand U4212 (N_4212,In_336,In_1287);
or U4213 (N_4213,In_956,In_313);
and U4214 (N_4214,In_767,In_1097);
and U4215 (N_4215,In_421,In_554);
nand U4216 (N_4216,In_274,In_33);
nor U4217 (N_4217,In_204,In_971);
nand U4218 (N_4218,In_1485,In_59);
and U4219 (N_4219,In_1038,In_784);
or U4220 (N_4220,In_113,In_120);
and U4221 (N_4221,In_682,In_1177);
nor U4222 (N_4222,In_1048,In_1405);
and U4223 (N_4223,In_858,In_103);
nand U4224 (N_4224,In_1209,In_768);
nor U4225 (N_4225,In_950,In_938);
and U4226 (N_4226,In_899,In_575);
and U4227 (N_4227,In_421,In_823);
or U4228 (N_4228,In_1005,In_700);
xnor U4229 (N_4229,In_449,In_178);
or U4230 (N_4230,In_357,In_1050);
and U4231 (N_4231,In_1303,In_726);
nor U4232 (N_4232,In_980,In_1025);
and U4233 (N_4233,In_438,In_1207);
nand U4234 (N_4234,In_1378,In_1216);
nor U4235 (N_4235,In_488,In_43);
nand U4236 (N_4236,In_422,In_20);
or U4237 (N_4237,In_1174,In_1152);
nor U4238 (N_4238,In_848,In_1419);
nand U4239 (N_4239,In_1220,In_163);
nor U4240 (N_4240,In_992,In_865);
nor U4241 (N_4241,In_368,In_331);
and U4242 (N_4242,In_1022,In_590);
and U4243 (N_4243,In_435,In_443);
or U4244 (N_4244,In_1480,In_177);
nor U4245 (N_4245,In_1138,In_1060);
and U4246 (N_4246,In_282,In_1225);
and U4247 (N_4247,In_1117,In_1102);
xor U4248 (N_4248,In_194,In_934);
nand U4249 (N_4249,In_1145,In_298);
nand U4250 (N_4250,In_145,In_420);
nand U4251 (N_4251,In_225,In_470);
nand U4252 (N_4252,In_1214,In_894);
nand U4253 (N_4253,In_1173,In_1178);
nand U4254 (N_4254,In_1482,In_824);
nand U4255 (N_4255,In_1214,In_1284);
or U4256 (N_4256,In_1496,In_1068);
and U4257 (N_4257,In_652,In_1004);
and U4258 (N_4258,In_455,In_1161);
nand U4259 (N_4259,In_1474,In_691);
and U4260 (N_4260,In_1296,In_558);
and U4261 (N_4261,In_196,In_1107);
nor U4262 (N_4262,In_564,In_727);
or U4263 (N_4263,In_499,In_706);
or U4264 (N_4264,In_1479,In_484);
xnor U4265 (N_4265,In_330,In_281);
nand U4266 (N_4266,In_35,In_74);
and U4267 (N_4267,In_1270,In_1458);
or U4268 (N_4268,In_719,In_778);
nand U4269 (N_4269,In_1360,In_245);
nand U4270 (N_4270,In_161,In_816);
and U4271 (N_4271,In_1118,In_153);
nor U4272 (N_4272,In_5,In_470);
nand U4273 (N_4273,In_63,In_522);
xnor U4274 (N_4274,In_1366,In_1447);
and U4275 (N_4275,In_179,In_138);
nand U4276 (N_4276,In_938,In_233);
nor U4277 (N_4277,In_670,In_1206);
nor U4278 (N_4278,In_548,In_638);
nor U4279 (N_4279,In_45,In_1325);
nor U4280 (N_4280,In_1190,In_1138);
nand U4281 (N_4281,In_907,In_362);
or U4282 (N_4282,In_842,In_981);
nor U4283 (N_4283,In_1253,In_1409);
nor U4284 (N_4284,In_621,In_55);
nand U4285 (N_4285,In_1431,In_1189);
or U4286 (N_4286,In_1447,In_1369);
and U4287 (N_4287,In_1175,In_198);
and U4288 (N_4288,In_244,In_837);
and U4289 (N_4289,In_1354,In_1305);
nand U4290 (N_4290,In_597,In_439);
and U4291 (N_4291,In_766,In_1319);
or U4292 (N_4292,In_710,In_737);
or U4293 (N_4293,In_387,In_1030);
and U4294 (N_4294,In_1437,In_930);
nand U4295 (N_4295,In_1253,In_328);
nor U4296 (N_4296,In_697,In_623);
and U4297 (N_4297,In_190,In_505);
xnor U4298 (N_4298,In_1388,In_1465);
xnor U4299 (N_4299,In_134,In_696);
nand U4300 (N_4300,In_655,In_302);
nor U4301 (N_4301,In_620,In_851);
nand U4302 (N_4302,In_949,In_499);
nand U4303 (N_4303,In_988,In_215);
nor U4304 (N_4304,In_239,In_799);
xnor U4305 (N_4305,In_992,In_27);
or U4306 (N_4306,In_847,In_646);
nand U4307 (N_4307,In_577,In_703);
nor U4308 (N_4308,In_510,In_307);
and U4309 (N_4309,In_1153,In_672);
nand U4310 (N_4310,In_1381,In_104);
nand U4311 (N_4311,In_1203,In_1043);
nor U4312 (N_4312,In_788,In_115);
or U4313 (N_4313,In_496,In_947);
nor U4314 (N_4314,In_77,In_1108);
and U4315 (N_4315,In_422,In_239);
and U4316 (N_4316,In_843,In_1247);
or U4317 (N_4317,In_782,In_973);
and U4318 (N_4318,In_556,In_34);
or U4319 (N_4319,In_1209,In_506);
and U4320 (N_4320,In_19,In_1316);
nand U4321 (N_4321,In_1242,In_327);
or U4322 (N_4322,In_731,In_312);
nand U4323 (N_4323,In_1394,In_1182);
nand U4324 (N_4324,In_535,In_1130);
nor U4325 (N_4325,In_817,In_362);
nor U4326 (N_4326,In_1096,In_1378);
or U4327 (N_4327,In_539,In_775);
or U4328 (N_4328,In_514,In_1397);
or U4329 (N_4329,In_1343,In_568);
and U4330 (N_4330,In_483,In_540);
and U4331 (N_4331,In_910,In_597);
or U4332 (N_4332,In_298,In_367);
nor U4333 (N_4333,In_272,In_41);
nand U4334 (N_4334,In_995,In_45);
xnor U4335 (N_4335,In_953,In_524);
nor U4336 (N_4336,In_352,In_259);
or U4337 (N_4337,In_831,In_1428);
nor U4338 (N_4338,In_567,In_457);
nand U4339 (N_4339,In_162,In_519);
and U4340 (N_4340,In_570,In_731);
and U4341 (N_4341,In_859,In_1054);
and U4342 (N_4342,In_939,In_43);
or U4343 (N_4343,In_1139,In_1183);
nand U4344 (N_4344,In_1127,In_371);
nor U4345 (N_4345,In_182,In_519);
nand U4346 (N_4346,In_25,In_1423);
nor U4347 (N_4347,In_1215,In_1303);
and U4348 (N_4348,In_518,In_378);
nand U4349 (N_4349,In_416,In_30);
and U4350 (N_4350,In_1475,In_951);
nand U4351 (N_4351,In_974,In_1495);
xnor U4352 (N_4352,In_805,In_765);
xor U4353 (N_4353,In_301,In_900);
nor U4354 (N_4354,In_1000,In_1306);
nand U4355 (N_4355,In_1260,In_1262);
nand U4356 (N_4356,In_257,In_733);
and U4357 (N_4357,In_1216,In_290);
or U4358 (N_4358,In_755,In_64);
xor U4359 (N_4359,In_682,In_1487);
or U4360 (N_4360,In_140,In_346);
and U4361 (N_4361,In_251,In_775);
and U4362 (N_4362,In_553,In_722);
nand U4363 (N_4363,In_1434,In_1068);
nor U4364 (N_4364,In_1070,In_1268);
nor U4365 (N_4365,In_1444,In_531);
nor U4366 (N_4366,In_44,In_16);
nor U4367 (N_4367,In_1394,In_1447);
nor U4368 (N_4368,In_504,In_1185);
or U4369 (N_4369,In_209,In_1420);
nand U4370 (N_4370,In_58,In_828);
nand U4371 (N_4371,In_913,In_460);
and U4372 (N_4372,In_941,In_258);
or U4373 (N_4373,In_1316,In_346);
xnor U4374 (N_4374,In_1104,In_870);
and U4375 (N_4375,In_47,In_320);
or U4376 (N_4376,In_708,In_365);
nor U4377 (N_4377,In_86,In_683);
nand U4378 (N_4378,In_668,In_1343);
nand U4379 (N_4379,In_719,In_1366);
and U4380 (N_4380,In_694,In_126);
and U4381 (N_4381,In_180,In_345);
nand U4382 (N_4382,In_1002,In_874);
or U4383 (N_4383,In_968,In_1300);
nand U4384 (N_4384,In_1299,In_218);
or U4385 (N_4385,In_288,In_1312);
and U4386 (N_4386,In_1276,In_62);
nor U4387 (N_4387,In_930,In_239);
and U4388 (N_4388,In_789,In_593);
nor U4389 (N_4389,In_1401,In_755);
nand U4390 (N_4390,In_615,In_449);
and U4391 (N_4391,In_282,In_287);
nand U4392 (N_4392,In_932,In_1107);
nand U4393 (N_4393,In_1287,In_763);
and U4394 (N_4394,In_572,In_579);
or U4395 (N_4395,In_998,In_1400);
or U4396 (N_4396,In_676,In_918);
nand U4397 (N_4397,In_353,In_1337);
nand U4398 (N_4398,In_233,In_670);
nor U4399 (N_4399,In_982,In_45);
or U4400 (N_4400,In_1288,In_920);
nor U4401 (N_4401,In_744,In_343);
nor U4402 (N_4402,In_237,In_222);
nand U4403 (N_4403,In_1366,In_971);
nor U4404 (N_4404,In_1496,In_829);
nor U4405 (N_4405,In_137,In_504);
nor U4406 (N_4406,In_132,In_1384);
and U4407 (N_4407,In_52,In_641);
nor U4408 (N_4408,In_42,In_14);
or U4409 (N_4409,In_203,In_1439);
or U4410 (N_4410,In_593,In_1161);
nor U4411 (N_4411,In_504,In_1241);
nor U4412 (N_4412,In_1438,In_991);
nand U4413 (N_4413,In_1216,In_918);
nor U4414 (N_4414,In_58,In_335);
nor U4415 (N_4415,In_731,In_1300);
and U4416 (N_4416,In_1171,In_136);
and U4417 (N_4417,In_317,In_1218);
nand U4418 (N_4418,In_303,In_155);
nor U4419 (N_4419,In_722,In_314);
and U4420 (N_4420,In_895,In_1176);
nand U4421 (N_4421,In_593,In_462);
nand U4422 (N_4422,In_1086,In_503);
or U4423 (N_4423,In_1309,In_143);
or U4424 (N_4424,In_886,In_730);
or U4425 (N_4425,In_886,In_407);
xnor U4426 (N_4426,In_791,In_150);
nor U4427 (N_4427,In_543,In_643);
and U4428 (N_4428,In_935,In_1035);
xor U4429 (N_4429,In_1400,In_907);
and U4430 (N_4430,In_19,In_481);
or U4431 (N_4431,In_459,In_1271);
nor U4432 (N_4432,In_1226,In_1092);
nand U4433 (N_4433,In_722,In_231);
nand U4434 (N_4434,In_789,In_848);
and U4435 (N_4435,In_1398,In_959);
or U4436 (N_4436,In_1312,In_15);
xor U4437 (N_4437,In_383,In_1499);
nand U4438 (N_4438,In_1453,In_368);
or U4439 (N_4439,In_315,In_593);
and U4440 (N_4440,In_1212,In_1200);
and U4441 (N_4441,In_1399,In_128);
nand U4442 (N_4442,In_1322,In_13);
nand U4443 (N_4443,In_585,In_1008);
nor U4444 (N_4444,In_546,In_862);
nand U4445 (N_4445,In_1051,In_585);
nand U4446 (N_4446,In_217,In_69);
nand U4447 (N_4447,In_682,In_1426);
xor U4448 (N_4448,In_981,In_310);
and U4449 (N_4449,In_25,In_306);
and U4450 (N_4450,In_799,In_360);
or U4451 (N_4451,In_1198,In_404);
nand U4452 (N_4452,In_669,In_1167);
nand U4453 (N_4453,In_160,In_909);
nand U4454 (N_4454,In_830,In_590);
or U4455 (N_4455,In_1390,In_1072);
or U4456 (N_4456,In_786,In_504);
nand U4457 (N_4457,In_251,In_1324);
xnor U4458 (N_4458,In_1122,In_27);
nor U4459 (N_4459,In_355,In_597);
nor U4460 (N_4460,In_114,In_1366);
xor U4461 (N_4461,In_1405,In_252);
nand U4462 (N_4462,In_1416,In_1146);
nand U4463 (N_4463,In_676,In_1002);
and U4464 (N_4464,In_1078,In_589);
xnor U4465 (N_4465,In_406,In_563);
or U4466 (N_4466,In_1261,In_176);
nor U4467 (N_4467,In_911,In_783);
nor U4468 (N_4468,In_59,In_3);
nand U4469 (N_4469,In_854,In_218);
nor U4470 (N_4470,In_421,In_1265);
nor U4471 (N_4471,In_1375,In_950);
nand U4472 (N_4472,In_922,In_612);
nand U4473 (N_4473,In_1448,In_1239);
nor U4474 (N_4474,In_691,In_626);
or U4475 (N_4475,In_772,In_1211);
or U4476 (N_4476,In_1066,In_1382);
nand U4477 (N_4477,In_86,In_393);
nand U4478 (N_4478,In_964,In_449);
nor U4479 (N_4479,In_9,In_269);
and U4480 (N_4480,In_280,In_1219);
nand U4481 (N_4481,In_1031,In_13);
or U4482 (N_4482,In_210,In_869);
xor U4483 (N_4483,In_938,In_405);
nor U4484 (N_4484,In_1225,In_619);
or U4485 (N_4485,In_1284,In_1078);
nor U4486 (N_4486,In_864,In_1265);
or U4487 (N_4487,In_59,In_742);
nor U4488 (N_4488,In_854,In_145);
nor U4489 (N_4489,In_1235,In_1264);
nor U4490 (N_4490,In_502,In_1244);
or U4491 (N_4491,In_1341,In_125);
nand U4492 (N_4492,In_602,In_1063);
or U4493 (N_4493,In_1439,In_1069);
nor U4494 (N_4494,In_424,In_1484);
nand U4495 (N_4495,In_811,In_205);
or U4496 (N_4496,In_1207,In_515);
nor U4497 (N_4497,In_1233,In_167);
nor U4498 (N_4498,In_920,In_1242);
or U4499 (N_4499,In_206,In_404);
nor U4500 (N_4500,In_1398,In_412);
nand U4501 (N_4501,In_1468,In_1302);
xnor U4502 (N_4502,In_609,In_65);
or U4503 (N_4503,In_1460,In_449);
nor U4504 (N_4504,In_1206,In_973);
nand U4505 (N_4505,In_81,In_1494);
and U4506 (N_4506,In_314,In_863);
or U4507 (N_4507,In_539,In_747);
nor U4508 (N_4508,In_781,In_804);
xnor U4509 (N_4509,In_261,In_95);
nor U4510 (N_4510,In_604,In_647);
nand U4511 (N_4511,In_72,In_237);
nor U4512 (N_4512,In_718,In_1154);
and U4513 (N_4513,In_1232,In_1055);
nand U4514 (N_4514,In_1122,In_0);
or U4515 (N_4515,In_519,In_508);
nand U4516 (N_4516,In_1194,In_117);
nand U4517 (N_4517,In_38,In_951);
nand U4518 (N_4518,In_913,In_461);
nor U4519 (N_4519,In_37,In_1188);
nor U4520 (N_4520,In_990,In_764);
and U4521 (N_4521,In_615,In_485);
xnor U4522 (N_4522,In_676,In_1385);
or U4523 (N_4523,In_506,In_1075);
xnor U4524 (N_4524,In_203,In_930);
nand U4525 (N_4525,In_826,In_32);
or U4526 (N_4526,In_431,In_1061);
or U4527 (N_4527,In_292,In_43);
nor U4528 (N_4528,In_774,In_880);
xnor U4529 (N_4529,In_1436,In_710);
nor U4530 (N_4530,In_846,In_843);
and U4531 (N_4531,In_1293,In_982);
nor U4532 (N_4532,In_430,In_13);
nor U4533 (N_4533,In_347,In_186);
nand U4534 (N_4534,In_789,In_957);
nand U4535 (N_4535,In_125,In_1155);
or U4536 (N_4536,In_545,In_862);
or U4537 (N_4537,In_1067,In_400);
or U4538 (N_4538,In_1425,In_193);
and U4539 (N_4539,In_29,In_1002);
and U4540 (N_4540,In_1267,In_394);
nand U4541 (N_4541,In_59,In_325);
nand U4542 (N_4542,In_603,In_392);
and U4543 (N_4543,In_824,In_457);
or U4544 (N_4544,In_748,In_1351);
and U4545 (N_4545,In_451,In_1390);
and U4546 (N_4546,In_407,In_193);
and U4547 (N_4547,In_252,In_545);
xor U4548 (N_4548,In_814,In_473);
nand U4549 (N_4549,In_1031,In_1040);
nor U4550 (N_4550,In_999,In_35);
or U4551 (N_4551,In_666,In_482);
and U4552 (N_4552,In_201,In_325);
nand U4553 (N_4553,In_815,In_30);
nor U4554 (N_4554,In_721,In_987);
nor U4555 (N_4555,In_1031,In_302);
and U4556 (N_4556,In_608,In_1005);
or U4557 (N_4557,In_410,In_1288);
nor U4558 (N_4558,In_1206,In_562);
and U4559 (N_4559,In_660,In_203);
nor U4560 (N_4560,In_915,In_1136);
nand U4561 (N_4561,In_28,In_1345);
or U4562 (N_4562,In_218,In_1259);
or U4563 (N_4563,In_1012,In_260);
or U4564 (N_4564,In_1456,In_1329);
nand U4565 (N_4565,In_549,In_253);
nor U4566 (N_4566,In_1118,In_1075);
nand U4567 (N_4567,In_104,In_353);
nand U4568 (N_4568,In_67,In_997);
and U4569 (N_4569,In_990,In_886);
nor U4570 (N_4570,In_224,In_460);
or U4571 (N_4571,In_121,In_1391);
nand U4572 (N_4572,In_1100,In_304);
nor U4573 (N_4573,In_660,In_218);
nor U4574 (N_4574,In_1003,In_377);
or U4575 (N_4575,In_1307,In_740);
nand U4576 (N_4576,In_407,In_759);
and U4577 (N_4577,In_646,In_1473);
nor U4578 (N_4578,In_141,In_62);
and U4579 (N_4579,In_121,In_967);
or U4580 (N_4580,In_1057,In_911);
or U4581 (N_4581,In_66,In_29);
nor U4582 (N_4582,In_281,In_1157);
nand U4583 (N_4583,In_752,In_1023);
and U4584 (N_4584,In_22,In_124);
nor U4585 (N_4585,In_720,In_219);
or U4586 (N_4586,In_1467,In_1088);
and U4587 (N_4587,In_648,In_633);
and U4588 (N_4588,In_1254,In_899);
and U4589 (N_4589,In_1277,In_751);
and U4590 (N_4590,In_643,In_1295);
nand U4591 (N_4591,In_834,In_177);
or U4592 (N_4592,In_830,In_35);
or U4593 (N_4593,In_688,In_2);
nand U4594 (N_4594,In_1480,In_850);
or U4595 (N_4595,In_817,In_137);
and U4596 (N_4596,In_971,In_196);
nor U4597 (N_4597,In_694,In_1009);
or U4598 (N_4598,In_141,In_512);
nor U4599 (N_4599,In_1490,In_133);
or U4600 (N_4600,In_12,In_644);
and U4601 (N_4601,In_447,In_75);
and U4602 (N_4602,In_680,In_1411);
nor U4603 (N_4603,In_375,In_1109);
nor U4604 (N_4604,In_303,In_1445);
and U4605 (N_4605,In_1448,In_965);
nor U4606 (N_4606,In_421,In_359);
xnor U4607 (N_4607,In_129,In_1266);
nor U4608 (N_4608,In_1150,In_410);
and U4609 (N_4609,In_384,In_455);
nand U4610 (N_4610,In_1237,In_1452);
nor U4611 (N_4611,In_1187,In_445);
nor U4612 (N_4612,In_76,In_1300);
and U4613 (N_4613,In_691,In_1292);
nor U4614 (N_4614,In_1385,In_1290);
nand U4615 (N_4615,In_395,In_394);
and U4616 (N_4616,In_64,In_1044);
xor U4617 (N_4617,In_981,In_1180);
or U4618 (N_4618,In_470,In_653);
and U4619 (N_4619,In_550,In_128);
nand U4620 (N_4620,In_2,In_554);
nor U4621 (N_4621,In_1204,In_33);
xor U4622 (N_4622,In_546,In_985);
nor U4623 (N_4623,In_487,In_283);
nor U4624 (N_4624,In_35,In_1295);
or U4625 (N_4625,In_1462,In_206);
nor U4626 (N_4626,In_207,In_832);
xnor U4627 (N_4627,In_1366,In_926);
or U4628 (N_4628,In_594,In_554);
or U4629 (N_4629,In_569,In_628);
nand U4630 (N_4630,In_669,In_132);
xor U4631 (N_4631,In_445,In_648);
nand U4632 (N_4632,In_354,In_1383);
and U4633 (N_4633,In_481,In_1055);
or U4634 (N_4634,In_418,In_504);
or U4635 (N_4635,In_668,In_949);
nand U4636 (N_4636,In_614,In_1442);
nor U4637 (N_4637,In_125,In_895);
and U4638 (N_4638,In_1046,In_1112);
nand U4639 (N_4639,In_687,In_1060);
nand U4640 (N_4640,In_1171,In_666);
and U4641 (N_4641,In_346,In_531);
nand U4642 (N_4642,In_213,In_1140);
or U4643 (N_4643,In_982,In_690);
and U4644 (N_4644,In_1418,In_533);
or U4645 (N_4645,In_66,In_976);
and U4646 (N_4646,In_981,In_1417);
and U4647 (N_4647,In_1307,In_413);
and U4648 (N_4648,In_1308,In_426);
nor U4649 (N_4649,In_556,In_1348);
or U4650 (N_4650,In_1087,In_1197);
nand U4651 (N_4651,In_104,In_667);
and U4652 (N_4652,In_868,In_104);
nand U4653 (N_4653,In_395,In_466);
nand U4654 (N_4654,In_122,In_892);
and U4655 (N_4655,In_1499,In_577);
xnor U4656 (N_4656,In_434,In_1475);
and U4657 (N_4657,In_311,In_1347);
or U4658 (N_4658,In_603,In_1096);
nor U4659 (N_4659,In_1110,In_1189);
or U4660 (N_4660,In_1217,In_233);
or U4661 (N_4661,In_1105,In_654);
or U4662 (N_4662,In_1173,In_1010);
or U4663 (N_4663,In_742,In_496);
or U4664 (N_4664,In_1069,In_1440);
or U4665 (N_4665,In_355,In_504);
and U4666 (N_4666,In_406,In_610);
and U4667 (N_4667,In_74,In_1442);
nand U4668 (N_4668,In_719,In_386);
nand U4669 (N_4669,In_820,In_412);
and U4670 (N_4670,In_1008,In_1153);
or U4671 (N_4671,In_343,In_824);
or U4672 (N_4672,In_889,In_1247);
and U4673 (N_4673,In_452,In_1482);
xor U4674 (N_4674,In_335,In_1376);
nand U4675 (N_4675,In_896,In_934);
and U4676 (N_4676,In_1201,In_1022);
nand U4677 (N_4677,In_1191,In_246);
or U4678 (N_4678,In_731,In_1463);
nand U4679 (N_4679,In_1367,In_115);
nor U4680 (N_4680,In_12,In_601);
and U4681 (N_4681,In_86,In_172);
nor U4682 (N_4682,In_1131,In_1337);
xnor U4683 (N_4683,In_1485,In_873);
or U4684 (N_4684,In_21,In_764);
or U4685 (N_4685,In_683,In_1203);
nor U4686 (N_4686,In_241,In_321);
nand U4687 (N_4687,In_1122,In_756);
nand U4688 (N_4688,In_766,In_1082);
or U4689 (N_4689,In_1089,In_711);
or U4690 (N_4690,In_1371,In_1460);
nand U4691 (N_4691,In_1488,In_3);
nand U4692 (N_4692,In_19,In_323);
nor U4693 (N_4693,In_115,In_580);
nor U4694 (N_4694,In_61,In_818);
nor U4695 (N_4695,In_1107,In_591);
or U4696 (N_4696,In_580,In_13);
or U4697 (N_4697,In_612,In_573);
nor U4698 (N_4698,In_807,In_1003);
nand U4699 (N_4699,In_1258,In_1136);
and U4700 (N_4700,In_681,In_337);
nand U4701 (N_4701,In_56,In_1260);
nand U4702 (N_4702,In_1494,In_539);
nand U4703 (N_4703,In_1147,In_1325);
or U4704 (N_4704,In_603,In_23);
or U4705 (N_4705,In_588,In_245);
nand U4706 (N_4706,In_1459,In_108);
xor U4707 (N_4707,In_387,In_84);
nor U4708 (N_4708,In_793,In_939);
or U4709 (N_4709,In_1255,In_1497);
or U4710 (N_4710,In_184,In_733);
xnor U4711 (N_4711,In_849,In_596);
nand U4712 (N_4712,In_264,In_300);
nand U4713 (N_4713,In_773,In_687);
nand U4714 (N_4714,In_770,In_224);
or U4715 (N_4715,In_62,In_246);
or U4716 (N_4716,In_347,In_85);
or U4717 (N_4717,In_1405,In_66);
nor U4718 (N_4718,In_1363,In_429);
or U4719 (N_4719,In_207,In_229);
xnor U4720 (N_4720,In_491,In_392);
or U4721 (N_4721,In_679,In_797);
and U4722 (N_4722,In_834,In_974);
nor U4723 (N_4723,In_1269,In_149);
nand U4724 (N_4724,In_291,In_1121);
nor U4725 (N_4725,In_1198,In_217);
nor U4726 (N_4726,In_1218,In_1014);
or U4727 (N_4727,In_621,In_517);
nor U4728 (N_4728,In_1240,In_830);
nor U4729 (N_4729,In_1210,In_992);
or U4730 (N_4730,In_507,In_133);
and U4731 (N_4731,In_347,In_1376);
or U4732 (N_4732,In_1404,In_112);
or U4733 (N_4733,In_156,In_1039);
nor U4734 (N_4734,In_628,In_1365);
nand U4735 (N_4735,In_308,In_447);
nor U4736 (N_4736,In_624,In_490);
and U4737 (N_4737,In_1468,In_1116);
and U4738 (N_4738,In_1200,In_748);
or U4739 (N_4739,In_237,In_102);
nor U4740 (N_4740,In_1118,In_1036);
and U4741 (N_4741,In_1061,In_1044);
nand U4742 (N_4742,In_278,In_207);
and U4743 (N_4743,In_1004,In_467);
nand U4744 (N_4744,In_156,In_491);
and U4745 (N_4745,In_911,In_397);
and U4746 (N_4746,In_388,In_220);
or U4747 (N_4747,In_1432,In_151);
and U4748 (N_4748,In_184,In_566);
and U4749 (N_4749,In_848,In_1400);
xor U4750 (N_4750,In_590,In_580);
and U4751 (N_4751,In_348,In_799);
nor U4752 (N_4752,In_633,In_190);
nand U4753 (N_4753,In_1417,In_165);
nor U4754 (N_4754,In_58,In_255);
or U4755 (N_4755,In_557,In_1143);
xor U4756 (N_4756,In_580,In_1297);
and U4757 (N_4757,In_733,In_1092);
nand U4758 (N_4758,In_366,In_827);
nor U4759 (N_4759,In_813,In_1288);
or U4760 (N_4760,In_466,In_420);
and U4761 (N_4761,In_704,In_467);
nand U4762 (N_4762,In_529,In_582);
nand U4763 (N_4763,In_26,In_613);
nor U4764 (N_4764,In_13,In_1085);
nand U4765 (N_4765,In_943,In_1372);
and U4766 (N_4766,In_1403,In_767);
xor U4767 (N_4767,In_1160,In_239);
nand U4768 (N_4768,In_48,In_635);
or U4769 (N_4769,In_514,In_1285);
and U4770 (N_4770,In_575,In_126);
nand U4771 (N_4771,In_272,In_678);
or U4772 (N_4772,In_238,In_1192);
or U4773 (N_4773,In_80,In_216);
nand U4774 (N_4774,In_1326,In_1028);
nor U4775 (N_4775,In_1399,In_693);
and U4776 (N_4776,In_736,In_466);
xnor U4777 (N_4777,In_1336,In_1216);
nand U4778 (N_4778,In_1016,In_760);
or U4779 (N_4779,In_1421,In_224);
xor U4780 (N_4780,In_34,In_15);
or U4781 (N_4781,In_920,In_1100);
and U4782 (N_4782,In_1056,In_1150);
or U4783 (N_4783,In_318,In_530);
nor U4784 (N_4784,In_754,In_759);
xor U4785 (N_4785,In_1314,In_779);
nor U4786 (N_4786,In_1266,In_96);
and U4787 (N_4787,In_579,In_52);
or U4788 (N_4788,In_1387,In_1403);
nand U4789 (N_4789,In_1120,In_801);
xor U4790 (N_4790,In_1312,In_519);
or U4791 (N_4791,In_156,In_690);
nand U4792 (N_4792,In_1472,In_378);
nor U4793 (N_4793,In_49,In_1239);
nand U4794 (N_4794,In_613,In_1477);
nor U4795 (N_4795,In_1228,In_1004);
or U4796 (N_4796,In_873,In_430);
or U4797 (N_4797,In_1030,In_330);
nand U4798 (N_4798,In_959,In_433);
or U4799 (N_4799,In_413,In_8);
xnor U4800 (N_4800,In_1245,In_1483);
nor U4801 (N_4801,In_49,In_455);
or U4802 (N_4802,In_768,In_876);
nand U4803 (N_4803,In_582,In_395);
nor U4804 (N_4804,In_1009,In_434);
or U4805 (N_4805,In_509,In_864);
nand U4806 (N_4806,In_908,In_1193);
and U4807 (N_4807,In_504,In_761);
nor U4808 (N_4808,In_1211,In_192);
and U4809 (N_4809,In_1066,In_37);
nand U4810 (N_4810,In_1193,In_613);
or U4811 (N_4811,In_418,In_1221);
nand U4812 (N_4812,In_714,In_282);
xnor U4813 (N_4813,In_259,In_541);
nor U4814 (N_4814,In_250,In_0);
nor U4815 (N_4815,In_729,In_270);
nor U4816 (N_4816,In_1306,In_124);
nand U4817 (N_4817,In_398,In_809);
or U4818 (N_4818,In_99,In_1395);
nor U4819 (N_4819,In_1385,In_730);
or U4820 (N_4820,In_1330,In_824);
xor U4821 (N_4821,In_759,In_1160);
xor U4822 (N_4822,In_362,In_482);
nor U4823 (N_4823,In_1415,In_776);
nor U4824 (N_4824,In_749,In_356);
and U4825 (N_4825,In_772,In_335);
and U4826 (N_4826,In_1041,In_903);
nor U4827 (N_4827,In_365,In_1211);
nand U4828 (N_4828,In_883,In_1196);
xor U4829 (N_4829,In_263,In_546);
or U4830 (N_4830,In_756,In_574);
nand U4831 (N_4831,In_1045,In_1105);
nand U4832 (N_4832,In_1032,In_776);
or U4833 (N_4833,In_953,In_44);
and U4834 (N_4834,In_641,In_596);
nor U4835 (N_4835,In_942,In_43);
nand U4836 (N_4836,In_630,In_1078);
xor U4837 (N_4837,In_1474,In_1027);
or U4838 (N_4838,In_136,In_417);
and U4839 (N_4839,In_31,In_808);
and U4840 (N_4840,In_596,In_1298);
or U4841 (N_4841,In_182,In_821);
or U4842 (N_4842,In_35,In_1418);
or U4843 (N_4843,In_60,In_1297);
nor U4844 (N_4844,In_765,In_359);
xnor U4845 (N_4845,In_608,In_32);
and U4846 (N_4846,In_588,In_846);
nor U4847 (N_4847,In_867,In_1456);
nor U4848 (N_4848,In_665,In_1305);
or U4849 (N_4849,In_1455,In_1043);
nor U4850 (N_4850,In_1041,In_1158);
nand U4851 (N_4851,In_577,In_648);
and U4852 (N_4852,In_889,In_877);
nand U4853 (N_4853,In_5,In_938);
nor U4854 (N_4854,In_128,In_944);
nor U4855 (N_4855,In_1218,In_312);
nand U4856 (N_4856,In_1125,In_513);
nand U4857 (N_4857,In_44,In_640);
xor U4858 (N_4858,In_757,In_412);
and U4859 (N_4859,In_322,In_369);
nor U4860 (N_4860,In_64,In_764);
and U4861 (N_4861,In_275,In_929);
nand U4862 (N_4862,In_562,In_1388);
xor U4863 (N_4863,In_136,In_1300);
or U4864 (N_4864,In_992,In_1295);
and U4865 (N_4865,In_331,In_1320);
nand U4866 (N_4866,In_1111,In_949);
xnor U4867 (N_4867,In_7,In_127);
or U4868 (N_4868,In_1236,In_1074);
nor U4869 (N_4869,In_248,In_1370);
nand U4870 (N_4870,In_93,In_24);
or U4871 (N_4871,In_247,In_121);
nand U4872 (N_4872,In_1235,In_469);
nand U4873 (N_4873,In_4,In_719);
and U4874 (N_4874,In_1029,In_1212);
or U4875 (N_4875,In_659,In_837);
or U4876 (N_4876,In_379,In_561);
or U4877 (N_4877,In_354,In_189);
or U4878 (N_4878,In_1191,In_677);
and U4879 (N_4879,In_1254,In_1379);
and U4880 (N_4880,In_638,In_1125);
and U4881 (N_4881,In_77,In_36);
or U4882 (N_4882,In_67,In_1204);
and U4883 (N_4883,In_686,In_101);
and U4884 (N_4884,In_1175,In_389);
and U4885 (N_4885,In_1101,In_495);
or U4886 (N_4886,In_880,In_883);
and U4887 (N_4887,In_655,In_202);
xnor U4888 (N_4888,In_787,In_1091);
and U4889 (N_4889,In_1392,In_1072);
and U4890 (N_4890,In_547,In_162);
nand U4891 (N_4891,In_60,In_204);
nand U4892 (N_4892,In_1430,In_519);
nor U4893 (N_4893,In_1252,In_1265);
nand U4894 (N_4894,In_44,In_375);
or U4895 (N_4895,In_934,In_542);
nor U4896 (N_4896,In_779,In_558);
nor U4897 (N_4897,In_683,In_1009);
nor U4898 (N_4898,In_488,In_1474);
or U4899 (N_4899,In_221,In_1280);
nand U4900 (N_4900,In_1186,In_1254);
nor U4901 (N_4901,In_12,In_919);
nor U4902 (N_4902,In_105,In_1302);
and U4903 (N_4903,In_847,In_1183);
or U4904 (N_4904,In_898,In_839);
nand U4905 (N_4905,In_55,In_503);
and U4906 (N_4906,In_895,In_590);
or U4907 (N_4907,In_972,In_1102);
and U4908 (N_4908,In_106,In_4);
and U4909 (N_4909,In_86,In_1319);
or U4910 (N_4910,In_194,In_1293);
xor U4911 (N_4911,In_618,In_355);
and U4912 (N_4912,In_1341,In_1349);
and U4913 (N_4913,In_1143,In_1473);
xor U4914 (N_4914,In_1268,In_65);
nor U4915 (N_4915,In_1021,In_904);
and U4916 (N_4916,In_881,In_295);
nand U4917 (N_4917,In_1227,In_1434);
nand U4918 (N_4918,In_1335,In_62);
nor U4919 (N_4919,In_500,In_391);
nand U4920 (N_4920,In_804,In_220);
xnor U4921 (N_4921,In_415,In_1045);
or U4922 (N_4922,In_414,In_276);
and U4923 (N_4923,In_1383,In_1024);
or U4924 (N_4924,In_523,In_101);
xor U4925 (N_4925,In_656,In_1064);
nand U4926 (N_4926,In_722,In_965);
nor U4927 (N_4927,In_370,In_172);
nand U4928 (N_4928,In_269,In_1215);
xor U4929 (N_4929,In_1344,In_473);
and U4930 (N_4930,In_216,In_426);
nand U4931 (N_4931,In_659,In_991);
and U4932 (N_4932,In_1435,In_802);
nand U4933 (N_4933,In_1057,In_179);
and U4934 (N_4934,In_1258,In_362);
nor U4935 (N_4935,In_944,In_1236);
or U4936 (N_4936,In_1420,In_377);
and U4937 (N_4937,In_1377,In_178);
nor U4938 (N_4938,In_1084,In_339);
nor U4939 (N_4939,In_744,In_1244);
and U4940 (N_4940,In_925,In_948);
nand U4941 (N_4941,In_1038,In_626);
or U4942 (N_4942,In_863,In_543);
xnor U4943 (N_4943,In_468,In_1225);
nand U4944 (N_4944,In_850,In_1448);
nor U4945 (N_4945,In_758,In_533);
nand U4946 (N_4946,In_767,In_96);
nor U4947 (N_4947,In_1453,In_548);
or U4948 (N_4948,In_629,In_1102);
nor U4949 (N_4949,In_1372,In_256);
xnor U4950 (N_4950,In_951,In_525);
nand U4951 (N_4951,In_401,In_1125);
nor U4952 (N_4952,In_227,In_618);
or U4953 (N_4953,In_1434,In_344);
nor U4954 (N_4954,In_1126,In_765);
and U4955 (N_4955,In_1485,In_290);
nor U4956 (N_4956,In_949,In_1435);
and U4957 (N_4957,In_1422,In_754);
nand U4958 (N_4958,In_1246,In_456);
or U4959 (N_4959,In_1298,In_1182);
or U4960 (N_4960,In_1277,In_1218);
and U4961 (N_4961,In_216,In_562);
nand U4962 (N_4962,In_1468,In_128);
or U4963 (N_4963,In_833,In_198);
and U4964 (N_4964,In_624,In_1175);
or U4965 (N_4965,In_1054,In_846);
nand U4966 (N_4966,In_927,In_476);
or U4967 (N_4967,In_735,In_706);
or U4968 (N_4968,In_815,In_1425);
and U4969 (N_4969,In_311,In_539);
nor U4970 (N_4970,In_1251,In_901);
nor U4971 (N_4971,In_485,In_1411);
or U4972 (N_4972,In_391,In_1005);
nand U4973 (N_4973,In_89,In_505);
or U4974 (N_4974,In_1091,In_1448);
nor U4975 (N_4975,In_1458,In_922);
nand U4976 (N_4976,In_646,In_1091);
xor U4977 (N_4977,In_1484,In_197);
nor U4978 (N_4978,In_1450,In_1453);
and U4979 (N_4979,In_918,In_299);
or U4980 (N_4980,In_1437,In_1187);
xor U4981 (N_4981,In_480,In_341);
or U4982 (N_4982,In_709,In_509);
and U4983 (N_4983,In_619,In_1440);
nor U4984 (N_4984,In_808,In_173);
and U4985 (N_4985,In_148,In_8);
or U4986 (N_4986,In_1008,In_305);
nor U4987 (N_4987,In_75,In_1312);
and U4988 (N_4988,In_1442,In_4);
and U4989 (N_4989,In_1104,In_771);
and U4990 (N_4990,In_1084,In_1363);
and U4991 (N_4991,In_456,In_767);
and U4992 (N_4992,In_1255,In_794);
or U4993 (N_4993,In_1379,In_163);
or U4994 (N_4994,In_1028,In_1468);
or U4995 (N_4995,In_931,In_786);
and U4996 (N_4996,In_594,In_531);
nand U4997 (N_4997,In_840,In_841);
nor U4998 (N_4998,In_1142,In_624);
nor U4999 (N_4999,In_77,In_1205);
nand U5000 (N_5000,N_3131,N_3270);
xnor U5001 (N_5001,N_1445,N_3438);
nor U5002 (N_5002,N_2495,N_1657);
xor U5003 (N_5003,N_4093,N_2591);
xor U5004 (N_5004,N_3931,N_1463);
and U5005 (N_5005,N_4723,N_1794);
or U5006 (N_5006,N_3196,N_2075);
xor U5007 (N_5007,N_4806,N_1414);
nand U5008 (N_5008,N_1387,N_1641);
and U5009 (N_5009,N_3732,N_4190);
xnor U5010 (N_5010,N_2066,N_3762);
or U5011 (N_5011,N_4519,N_699);
nor U5012 (N_5012,N_1655,N_4758);
nand U5013 (N_5013,N_4145,N_1780);
nand U5014 (N_5014,N_4702,N_1553);
and U5015 (N_5015,N_1732,N_2359);
and U5016 (N_5016,N_4315,N_2839);
and U5017 (N_5017,N_3200,N_2767);
nand U5018 (N_5018,N_2830,N_2453);
and U5019 (N_5019,N_3437,N_3230);
and U5020 (N_5020,N_3203,N_4938);
and U5021 (N_5021,N_342,N_4631);
or U5022 (N_5022,N_1072,N_2563);
and U5023 (N_5023,N_1049,N_515);
nand U5024 (N_5024,N_2211,N_2817);
nand U5025 (N_5025,N_3633,N_4);
nand U5026 (N_5026,N_4694,N_2514);
nand U5027 (N_5027,N_1244,N_54);
or U5028 (N_5028,N_4414,N_2366);
and U5029 (N_5029,N_2794,N_21);
and U5030 (N_5030,N_615,N_2479);
and U5031 (N_5031,N_3764,N_2291);
nor U5032 (N_5032,N_622,N_3686);
nor U5033 (N_5033,N_190,N_4900);
nand U5034 (N_5034,N_4784,N_4704);
nand U5035 (N_5035,N_597,N_87);
or U5036 (N_5036,N_1186,N_4061);
xor U5037 (N_5037,N_3356,N_2086);
nand U5038 (N_5038,N_1385,N_3706);
or U5039 (N_5039,N_4304,N_1480);
nor U5040 (N_5040,N_3249,N_655);
nand U5041 (N_5041,N_726,N_800);
and U5042 (N_5042,N_1682,N_4248);
and U5043 (N_5043,N_1241,N_4720);
and U5044 (N_5044,N_4110,N_2678);
nor U5045 (N_5045,N_72,N_4790);
nand U5046 (N_5046,N_2009,N_976);
nand U5047 (N_5047,N_78,N_3174);
or U5048 (N_5048,N_4889,N_4818);
nand U5049 (N_5049,N_3986,N_1420);
nor U5050 (N_5050,N_2543,N_3545);
nor U5051 (N_5051,N_2094,N_1129);
nand U5052 (N_5052,N_3665,N_1520);
nand U5053 (N_5053,N_4284,N_2599);
nand U5054 (N_5054,N_658,N_2774);
or U5055 (N_5055,N_3508,N_4976);
xnor U5056 (N_5056,N_1995,N_3004);
or U5057 (N_5057,N_4984,N_1524);
and U5058 (N_5058,N_39,N_3096);
nor U5059 (N_5059,N_2071,N_3324);
and U5060 (N_5060,N_4430,N_3195);
or U5061 (N_5061,N_1119,N_4876);
and U5062 (N_5062,N_1774,N_3483);
nor U5063 (N_5063,N_3370,N_508);
nand U5064 (N_5064,N_486,N_2402);
nor U5065 (N_5065,N_4004,N_867);
nor U5066 (N_5066,N_4579,N_775);
and U5067 (N_5067,N_34,N_1556);
xor U5068 (N_5068,N_2455,N_2552);
nand U5069 (N_5069,N_466,N_2301);
or U5070 (N_5070,N_4402,N_1474);
and U5071 (N_5071,N_4461,N_3868);
nand U5072 (N_5072,N_2899,N_3977);
and U5073 (N_5073,N_3962,N_745);
or U5074 (N_5074,N_1006,N_1018);
and U5075 (N_5075,N_3002,N_2056);
or U5076 (N_5076,N_2281,N_29);
or U5077 (N_5077,N_1433,N_246);
and U5078 (N_5078,N_2815,N_1290);
nor U5079 (N_5079,N_654,N_2909);
nor U5080 (N_5080,N_4051,N_3472);
nor U5081 (N_5081,N_3458,N_4059);
and U5082 (N_5082,N_3973,N_3617);
or U5083 (N_5083,N_1191,N_4003);
xnor U5084 (N_5084,N_1711,N_4874);
and U5085 (N_5085,N_4858,N_3759);
or U5086 (N_5086,N_4592,N_4877);
nor U5087 (N_5087,N_1260,N_1882);
nor U5088 (N_5088,N_4026,N_2620);
xnor U5089 (N_5089,N_4320,N_4305);
nand U5090 (N_5090,N_963,N_2554);
nand U5091 (N_5091,N_2354,N_563);
nand U5092 (N_5092,N_2394,N_3202);
or U5093 (N_5093,N_1771,N_2714);
and U5094 (N_5094,N_2348,N_1784);
or U5095 (N_5095,N_1533,N_1775);
nor U5096 (N_5096,N_1997,N_631);
nand U5097 (N_5097,N_1605,N_2446);
nor U5098 (N_5098,N_3295,N_2014);
nand U5099 (N_5099,N_4030,N_1615);
nor U5100 (N_5100,N_3741,N_3276);
and U5101 (N_5101,N_1267,N_4306);
nand U5102 (N_5102,N_3242,N_2340);
and U5103 (N_5103,N_3021,N_3591);
and U5104 (N_5104,N_1717,N_4184);
nand U5105 (N_5105,N_103,N_1261);
nand U5106 (N_5106,N_871,N_3014);
or U5107 (N_5107,N_973,N_785);
nor U5108 (N_5108,N_4431,N_2061);
or U5109 (N_5109,N_101,N_3898);
nor U5110 (N_5110,N_3996,N_4355);
or U5111 (N_5111,N_3907,N_4892);
xnor U5112 (N_5112,N_3079,N_4880);
nor U5113 (N_5113,N_3226,N_2537);
or U5114 (N_5114,N_4395,N_4528);
and U5115 (N_5115,N_1767,N_4389);
nand U5116 (N_5116,N_3811,N_3392);
and U5117 (N_5117,N_375,N_2936);
nor U5118 (N_5118,N_3779,N_2037);
nand U5119 (N_5119,N_3045,N_2046);
nand U5120 (N_5120,N_231,N_2755);
and U5121 (N_5121,N_3170,N_4041);
and U5122 (N_5122,N_4529,N_3068);
and U5123 (N_5123,N_4071,N_2533);
and U5124 (N_5124,N_4244,N_299);
or U5125 (N_5125,N_4820,N_3780);
xnor U5126 (N_5126,N_3336,N_1522);
or U5127 (N_5127,N_1800,N_3103);
xnor U5128 (N_5128,N_4252,N_2523);
or U5129 (N_5129,N_2991,N_4356);
or U5130 (N_5130,N_520,N_71);
xnor U5131 (N_5131,N_3168,N_2186);
and U5132 (N_5132,N_2797,N_4985);
nor U5133 (N_5133,N_1280,N_363);
and U5134 (N_5134,N_1663,N_1406);
nand U5135 (N_5135,N_2931,N_4478);
nand U5136 (N_5136,N_1589,N_4640);
nand U5137 (N_5137,N_860,N_4846);
xor U5138 (N_5138,N_3445,N_683);
nor U5139 (N_5139,N_3711,N_192);
and U5140 (N_5140,N_707,N_2146);
or U5141 (N_5141,N_3217,N_3708);
nand U5142 (N_5142,N_58,N_1078);
nor U5143 (N_5143,N_3109,N_4118);
or U5144 (N_5144,N_3668,N_4031);
xor U5145 (N_5145,N_894,N_4235);
xor U5146 (N_5146,N_801,N_2841);
nor U5147 (N_5147,N_1617,N_3638);
and U5148 (N_5148,N_2639,N_853);
and U5149 (N_5149,N_1360,N_3085);
or U5150 (N_5150,N_1301,N_971);
nor U5151 (N_5151,N_2886,N_915);
xor U5152 (N_5152,N_3468,N_1506);
nand U5153 (N_5153,N_3790,N_2);
nand U5154 (N_5154,N_730,N_585);
and U5155 (N_5155,N_3658,N_1240);
nand U5156 (N_5156,N_3705,N_1408);
or U5157 (N_5157,N_1745,N_1176);
nand U5158 (N_5158,N_2214,N_2199);
nor U5159 (N_5159,N_438,N_1332);
nor U5160 (N_5160,N_3024,N_2885);
nor U5161 (N_5161,N_4780,N_2278);
nor U5162 (N_5162,N_2303,N_1528);
nand U5163 (N_5163,N_1237,N_529);
and U5164 (N_5164,N_4522,N_4368);
nand U5165 (N_5165,N_1144,N_470);
nand U5166 (N_5166,N_1600,N_282);
nand U5167 (N_5167,N_2665,N_3173);
nor U5168 (N_5168,N_756,N_4617);
and U5169 (N_5169,N_3802,N_4432);
nor U5170 (N_5170,N_4307,N_846);
nand U5171 (N_5171,N_4839,N_2357);
and U5172 (N_5172,N_580,N_4762);
nand U5173 (N_5173,N_3225,N_1935);
and U5174 (N_5174,N_420,N_290);
nand U5175 (N_5175,N_2655,N_4745);
or U5176 (N_5176,N_2487,N_1287);
nor U5177 (N_5177,N_530,N_3894);
nand U5178 (N_5178,N_145,N_2541);
nor U5179 (N_5179,N_532,N_2522);
nand U5180 (N_5180,N_857,N_1121);
and U5181 (N_5181,N_869,N_3729);
and U5182 (N_5182,N_904,N_4721);
and U5183 (N_5183,N_2410,N_1491);
xor U5184 (N_5184,N_2145,N_3435);
xor U5185 (N_5185,N_63,N_2089);
xnor U5186 (N_5186,N_874,N_168);
nand U5187 (N_5187,N_4209,N_980);
nor U5188 (N_5188,N_3541,N_613);
nand U5189 (N_5189,N_1854,N_447);
or U5190 (N_5190,N_999,N_310);
nand U5191 (N_5191,N_4486,N_4840);
and U5192 (N_5192,N_3001,N_3123);
nor U5193 (N_5193,N_2188,N_2994);
nor U5194 (N_5194,N_4805,N_1976);
nand U5195 (N_5195,N_2265,N_2945);
nand U5196 (N_5196,N_2047,N_1544);
xnor U5197 (N_5197,N_4753,N_2898);
xor U5198 (N_5198,N_2632,N_2738);
nand U5199 (N_5199,N_1590,N_4379);
nand U5200 (N_5200,N_4114,N_2651);
xnor U5201 (N_5201,N_4958,N_2234);
nand U5202 (N_5202,N_1943,N_4300);
nand U5203 (N_5203,N_3743,N_4772);
nand U5204 (N_5204,N_4002,N_979);
nor U5205 (N_5205,N_2571,N_1094);
nand U5206 (N_5206,N_2822,N_1559);
nand U5207 (N_5207,N_653,N_3308);
nand U5208 (N_5208,N_1737,N_3925);
nand U5209 (N_5209,N_3426,N_1369);
and U5210 (N_5210,N_3506,N_1132);
or U5211 (N_5211,N_3467,N_479);
nor U5212 (N_5212,N_3179,N_3129);
nor U5213 (N_5213,N_2572,N_2165);
and U5214 (N_5214,N_33,N_2102);
or U5215 (N_5215,N_4154,N_2360);
and U5216 (N_5216,N_1727,N_3423);
nor U5217 (N_5217,N_1405,N_4448);
and U5218 (N_5218,N_4352,N_4278);
or U5219 (N_5219,N_2198,N_1469);
and U5220 (N_5220,N_1424,N_942);
and U5221 (N_5221,N_4401,N_1623);
or U5222 (N_5222,N_1877,N_3219);
and U5223 (N_5223,N_1541,N_457);
nand U5224 (N_5224,N_2283,N_1333);
nand U5225 (N_5225,N_2613,N_2203);
nand U5226 (N_5226,N_2713,N_4345);
nor U5227 (N_5227,N_3262,N_3728);
nand U5228 (N_5228,N_4783,N_3239);
nand U5229 (N_5229,N_3212,N_4919);
nand U5230 (N_5230,N_2733,N_4761);
nand U5231 (N_5231,N_3836,N_189);
and U5232 (N_5232,N_4654,N_1439);
nand U5233 (N_5233,N_2229,N_1248);
and U5234 (N_5234,N_1157,N_329);
nand U5235 (N_5235,N_2793,N_2010);
or U5236 (N_5236,N_1123,N_3788);
nor U5237 (N_5237,N_1878,N_4104);
or U5238 (N_5238,N_461,N_2317);
xor U5239 (N_5239,N_2057,N_3293);
or U5240 (N_5240,N_76,N_1743);
nand U5241 (N_5241,N_2459,N_3703);
or U5242 (N_5242,N_1869,N_4664);
and U5243 (N_5243,N_56,N_2473);
nor U5244 (N_5244,N_3756,N_1308);
nor U5245 (N_5245,N_119,N_4211);
nor U5246 (N_5246,N_810,N_374);
or U5247 (N_5247,N_1105,N_1550);
or U5248 (N_5248,N_687,N_2378);
nand U5249 (N_5249,N_1453,N_3151);
and U5250 (N_5250,N_3187,N_1977);
xor U5251 (N_5251,N_3882,N_2718);
and U5252 (N_5252,N_3930,N_3035);
or U5253 (N_5253,N_3067,N_1136);
or U5254 (N_5254,N_638,N_2395);
nand U5255 (N_5255,N_284,N_1223);
and U5256 (N_5256,N_1493,N_3422);
xor U5257 (N_5257,N_1970,N_4511);
or U5258 (N_5258,N_4498,N_3229);
nor U5259 (N_5259,N_4347,N_127);
nand U5260 (N_5260,N_3012,N_3715);
and U5261 (N_5261,N_4527,N_4972);
or U5262 (N_5262,N_4491,N_698);
or U5263 (N_5263,N_4400,N_3030);
or U5264 (N_5264,N_817,N_3121);
and U5265 (N_5265,N_3440,N_155);
or U5266 (N_5266,N_3522,N_808);
nor U5267 (N_5267,N_309,N_4020);
nor U5268 (N_5268,N_1959,N_1749);
or U5269 (N_5269,N_3888,N_3403);
nand U5270 (N_5270,N_4800,N_2518);
nand U5271 (N_5271,N_1835,N_4497);
and U5272 (N_5272,N_1650,N_4586);
or U5273 (N_5273,N_1838,N_3433);
nand U5274 (N_5274,N_1195,N_3318);
nor U5275 (N_5275,N_2386,N_998);
and U5276 (N_5276,N_300,N_901);
or U5277 (N_5277,N_2083,N_826);
and U5278 (N_5278,N_3702,N_1020);
nand U5279 (N_5279,N_4436,N_3512);
nor U5280 (N_5280,N_1687,N_94);
or U5281 (N_5281,N_3495,N_4397);
or U5282 (N_5282,N_3555,N_4968);
nand U5283 (N_5283,N_126,N_4339);
xnor U5284 (N_5284,N_1591,N_4999);
nor U5285 (N_5285,N_803,N_3290);
nand U5286 (N_5286,N_3010,N_4099);
nor U5287 (N_5287,N_2058,N_4923);
xor U5288 (N_5288,N_2197,N_4655);
or U5289 (N_5289,N_3935,N_2008);
nand U5290 (N_5290,N_889,N_1677);
nor U5291 (N_5291,N_3338,N_334);
or U5292 (N_5292,N_4973,N_1305);
nand U5293 (N_5293,N_3525,N_3590);
or U5294 (N_5294,N_1972,N_1486);
nor U5295 (N_5295,N_3951,N_4821);
and U5296 (N_5296,N_3439,N_665);
or U5297 (N_5297,N_1418,N_4731);
or U5298 (N_5298,N_2418,N_4204);
nor U5299 (N_5299,N_3709,N_2421);
nor U5300 (N_5300,N_1887,N_2493);
xor U5301 (N_5301,N_956,N_11);
nand U5302 (N_5302,N_2013,N_4692);
xor U5303 (N_5303,N_747,N_1504);
or U5304 (N_5304,N_1725,N_1907);
or U5305 (N_5305,N_3287,N_3415);
or U5306 (N_5306,N_3650,N_688);
or U5307 (N_5307,N_620,N_1404);
and U5308 (N_5308,N_2673,N_1523);
nor U5309 (N_5309,N_1025,N_462);
nor U5310 (N_5310,N_4964,N_1461);
or U5311 (N_5311,N_4180,N_4130);
nand U5312 (N_5312,N_4263,N_4213);
or U5313 (N_5313,N_1850,N_3223);
and U5314 (N_5314,N_2765,N_908);
and U5315 (N_5315,N_82,N_749);
or U5316 (N_5316,N_1434,N_4610);
nor U5317 (N_5317,N_332,N_1194);
and U5318 (N_5318,N_2576,N_2468);
and U5319 (N_5319,N_2350,N_427);
and U5320 (N_5320,N_3569,N_1697);
or U5321 (N_5321,N_2808,N_3774);
nand U5322 (N_5322,N_2245,N_771);
nor U5323 (N_5323,N_629,N_2049);
and U5324 (N_5324,N_4690,N_3858);
and U5325 (N_5325,N_3358,N_1546);
nor U5326 (N_5326,N_2926,N_344);
nor U5327 (N_5327,N_1001,N_4273);
or U5328 (N_5328,N_368,N_985);
nand U5329 (N_5329,N_2215,N_414);
nor U5330 (N_5330,N_2568,N_444);
and U5331 (N_5331,N_2825,N_2752);
nor U5332 (N_5332,N_1627,N_4802);
nand U5333 (N_5333,N_2757,N_798);
nor U5334 (N_5334,N_2085,N_2741);
or U5335 (N_5335,N_1302,N_4878);
nand U5336 (N_5336,N_1307,N_4728);
nand U5337 (N_5337,N_1295,N_3886);
and U5338 (N_5338,N_1656,N_848);
nor U5339 (N_5339,N_1505,N_718);
or U5340 (N_5340,N_575,N_291);
and U5341 (N_5341,N_4303,N_4633);
or U5342 (N_5342,N_3821,N_4779);
and U5343 (N_5343,N_2759,N_2954);
nand U5344 (N_5344,N_1510,N_2393);
nor U5345 (N_5345,N_2477,N_4903);
and U5346 (N_5346,N_3165,N_2087);
or U5347 (N_5347,N_1188,N_1823);
nand U5348 (N_5348,N_2849,N_3602);
or U5349 (N_5349,N_2528,N_2411);
and U5350 (N_5350,N_2963,N_1350);
or U5351 (N_5351,N_4649,N_1905);
nor U5352 (N_5352,N_3000,N_4713);
and U5353 (N_5353,N_4082,N_4293);
nor U5354 (N_5354,N_2905,N_3310);
and U5355 (N_5355,N_1938,N_635);
nand U5356 (N_5356,N_647,N_1017);
xnor U5357 (N_5357,N_451,N_648);
nand U5358 (N_5358,N_4008,N_4852);
nor U5359 (N_5359,N_4010,N_579);
nor U5360 (N_5360,N_19,N_257);
and U5361 (N_5361,N_4064,N_693);
and U5362 (N_5362,N_411,N_1185);
nand U5363 (N_5363,N_3965,N_2730);
nand U5364 (N_5364,N_2476,N_1688);
or U5365 (N_5365,N_206,N_2790);
nand U5366 (N_5366,N_3427,N_1968);
or U5367 (N_5367,N_1104,N_1777);
nor U5368 (N_5368,N_366,N_2792);
nor U5369 (N_5369,N_1916,N_4440);
or U5370 (N_5370,N_1093,N_2124);
and U5371 (N_5371,N_4788,N_1450);
nand U5372 (N_5372,N_1353,N_2645);
nand U5373 (N_5373,N_4993,N_150);
nor U5374 (N_5374,N_1011,N_1376);
nand U5375 (N_5375,N_4374,N_704);
nand U5376 (N_5376,N_1828,N_3059);
or U5377 (N_5377,N_4754,N_3274);
and U5378 (N_5378,N_4358,N_204);
nand U5379 (N_5379,N_2436,N_4137);
nor U5380 (N_5380,N_1639,N_1359);
nand U5381 (N_5381,N_2195,N_151);
xnor U5382 (N_5382,N_4542,N_4768);
nor U5383 (N_5383,N_1648,N_3317);
or U5384 (N_5384,N_1824,N_1515);
nand U5385 (N_5385,N_3847,N_3871);
xor U5386 (N_5386,N_1028,N_1014);
and U5387 (N_5387,N_171,N_4019);
and U5388 (N_5388,N_1631,N_2968);
xor U5389 (N_5389,N_968,N_2525);
nand U5390 (N_5390,N_1162,N_50);
and U5391 (N_5391,N_4626,N_3610);
or U5392 (N_5392,N_4891,N_2427);
nand U5393 (N_5393,N_3379,N_3950);
xnor U5394 (N_5394,N_2966,N_1091);
or U5395 (N_5395,N_4726,N_4144);
and U5396 (N_5396,N_4441,N_2840);
and U5397 (N_5397,N_3843,N_201);
and U5398 (N_5398,N_158,N_361);
or U5399 (N_5399,N_3425,N_509);
and U5400 (N_5400,N_1137,N_3716);
nand U5401 (N_5401,N_3016,N_2212);
nand U5402 (N_5402,N_370,N_3253);
nand U5403 (N_5403,N_2458,N_4865);
or U5404 (N_5404,N_858,N_3354);
nor U5405 (N_5405,N_4333,N_3606);
nor U5406 (N_5406,N_4171,N_4613);
xor U5407 (N_5407,N_3803,N_3044);
xnor U5408 (N_5408,N_2220,N_2464);
nor U5409 (N_5409,N_4058,N_3201);
nor U5410 (N_5410,N_3353,N_2433);
and U5411 (N_5411,N_3106,N_3988);
or U5412 (N_5412,N_662,N_1785);
and U5413 (N_5413,N_61,N_1757);
or U5414 (N_5414,N_3837,N_3971);
and U5415 (N_5415,N_3688,N_1399);
or U5416 (N_5416,N_849,N_3361);
and U5417 (N_5417,N_1833,N_3775);
nand U5418 (N_5418,N_1348,N_4424);
and U5419 (N_5419,N_1354,N_809);
nand U5420 (N_5420,N_1716,N_3752);
and U5421 (N_5421,N_2520,N_3550);
nor U5422 (N_5422,N_2798,N_3322);
nand U5423 (N_5423,N_526,N_1994);
nor U5424 (N_5424,N_4237,N_3833);
nor U5425 (N_5425,N_3450,N_97);
or U5426 (N_5426,N_1042,N_3535);
xor U5427 (N_5427,N_4123,N_3940);
or U5428 (N_5428,N_1135,N_2486);
and U5429 (N_5429,N_1696,N_2654);
and U5430 (N_5430,N_4111,N_4457);
nand U5431 (N_5431,N_2590,N_3020);
nor U5432 (N_5432,N_3527,N_397);
nand U5433 (N_5433,N_727,N_2248);
or U5434 (N_5434,N_3405,N_728);
and U5435 (N_5435,N_298,N_1320);
nor U5436 (N_5436,N_1457,N_1552);
nor U5437 (N_5437,N_2895,N_129);
or U5438 (N_5438,N_2893,N_2007);
nor U5439 (N_5439,N_1343,N_2600);
and U5440 (N_5440,N_4134,N_425);
xnor U5441 (N_5441,N_3357,N_469);
and U5442 (N_5442,N_1181,N_4264);
nor U5443 (N_5443,N_3875,N_731);
nand U5444 (N_5444,N_4513,N_1558);
or U5445 (N_5445,N_4125,N_2469);
and U5446 (N_5446,N_177,N_2305);
and U5447 (N_5447,N_3747,N_584);
and U5448 (N_5448,N_3529,N_3490);
and U5449 (N_5449,N_2163,N_2630);
and U5450 (N_5450,N_1671,N_2351);
or U5451 (N_5451,N_4098,N_1204);
nor U5452 (N_5452,N_3320,N_3629);
and U5453 (N_5453,N_98,N_4944);
nand U5454 (N_5454,N_141,N_3777);
or U5455 (N_5455,N_765,N_2930);
or U5456 (N_5456,N_634,N_138);
or U5457 (N_5457,N_67,N_2999);
and U5458 (N_5458,N_3853,N_3404);
nand U5459 (N_5459,N_2597,N_1391);
and U5460 (N_5460,N_4420,N_3974);
nand U5461 (N_5461,N_3880,N_981);
xnor U5462 (N_5462,N_4219,N_561);
nand U5463 (N_5463,N_1703,N_851);
nor U5464 (N_5464,N_824,N_3690);
nand U5465 (N_5465,N_1090,N_4142);
nand U5466 (N_5466,N_557,N_2423);
nand U5467 (N_5467,N_4712,N_2890);
nand U5468 (N_5468,N_4666,N_666);
or U5469 (N_5469,N_689,N_467);
and U5470 (N_5470,N_14,N_1529);
nand U5471 (N_5471,N_4539,N_4062);
nor U5472 (N_5472,N_234,N_4764);
or U5473 (N_5473,N_1815,N_340);
or U5474 (N_5474,N_1294,N_64);
nand U5475 (N_5475,N_3341,N_1724);
nor U5476 (N_5476,N_705,N_4991);
or U5477 (N_5477,N_2055,N_287);
nand U5478 (N_5478,N_3934,N_3194);
nor U5479 (N_5479,N_4158,N_4047);
nand U5480 (N_5480,N_540,N_4087);
or U5481 (N_5481,N_2609,N_3180);
nand U5482 (N_5482,N_237,N_571);
nor U5483 (N_5483,N_1429,N_4568);
or U5484 (N_5484,N_3749,N_4054);
or U5485 (N_5485,N_1791,N_4868);
and U5486 (N_5486,N_4587,N_610);
xor U5487 (N_5487,N_3135,N_3351);
and U5488 (N_5488,N_1951,N_4599);
nand U5489 (N_5489,N_4635,N_2135);
nand U5490 (N_5490,N_4727,N_1560);
nor U5491 (N_5491,N_4129,N_1079);
nand U5492 (N_5492,N_1371,N_1939);
nor U5493 (N_5493,N_2318,N_3723);
nand U5494 (N_5494,N_891,N_2851);
or U5495 (N_5495,N_2346,N_4826);
nor U5496 (N_5496,N_754,N_1067);
or U5497 (N_5497,N_3663,N_4052);
or U5498 (N_5498,N_1608,N_2863);
nor U5499 (N_5499,N_4479,N_3546);
nand U5500 (N_5500,N_709,N_3247);
nor U5501 (N_5501,N_1044,N_10);
or U5502 (N_5502,N_2388,N_553);
and U5503 (N_5503,N_1489,N_3725);
xnor U5504 (N_5504,N_1728,N_3984);
or U5505 (N_5505,N_4165,N_1415);
xor U5506 (N_5506,N_1860,N_3386);
and U5507 (N_5507,N_3693,N_1957);
nor U5508 (N_5508,N_4733,N_3921);
nor U5509 (N_5509,N_1146,N_1084);
xor U5510 (N_5510,N_4823,N_3205);
nor U5511 (N_5511,N_2619,N_1945);
or U5512 (N_5512,N_2638,N_814);
and U5513 (N_5513,N_4810,N_2080);
nor U5514 (N_5514,N_1233,N_3534);
nand U5515 (N_5515,N_2196,N_2799);
or U5516 (N_5516,N_2550,N_3264);
or U5517 (N_5517,N_3186,N_3049);
xnor U5518 (N_5518,N_1148,N_3822);
nand U5519 (N_5519,N_369,N_2431);
nor U5520 (N_5520,N_2784,N_2553);
xnor U5521 (N_5521,N_1825,N_2623);
nand U5522 (N_5522,N_3607,N_182);
nand U5523 (N_5523,N_3687,N_2297);
nor U5524 (N_5524,N_3250,N_4824);
or U5525 (N_5525,N_3678,N_1582);
nand U5526 (N_5526,N_116,N_1534);
or U5527 (N_5527,N_3497,N_2882);
and U5528 (N_5528,N_65,N_2961);
nand U5529 (N_5529,N_3664,N_153);
nor U5530 (N_5530,N_1834,N_1595);
or U5531 (N_5531,N_3443,N_1885);
nand U5532 (N_5532,N_4905,N_733);
and U5533 (N_5533,N_3899,N_788);
and U5534 (N_5534,N_2239,N_1087);
nand U5535 (N_5535,N_1936,N_4842);
nor U5536 (N_5536,N_1875,N_18);
or U5537 (N_5537,N_1499,N_4700);
or U5538 (N_5538,N_2462,N_4926);
nor U5539 (N_5539,N_3070,N_2972);
nand U5540 (N_5540,N_167,N_4815);
and U5541 (N_5541,N_4977,N_1043);
nand U5542 (N_5542,N_4243,N_518);
and U5543 (N_5543,N_4998,N_3887);
or U5544 (N_5544,N_1427,N_3018);
and U5545 (N_5545,N_389,N_3909);
or U5546 (N_5546,N_2024,N_3161);
nor U5547 (N_5547,N_233,N_2096);
nor U5548 (N_5548,N_2530,N_463);
and U5549 (N_5549,N_627,N_842);
xnor U5550 (N_5550,N_4541,N_2309);
nor U5551 (N_5551,N_3549,N_3034);
nand U5552 (N_5552,N_3388,N_3643);
nand U5553 (N_5553,N_1681,N_1518);
nor U5554 (N_5554,N_4228,N_3207);
nand U5555 (N_5555,N_1019,N_989);
and U5556 (N_5556,N_3855,N_3713);
and U5557 (N_5557,N_2745,N_1401);
nand U5558 (N_5558,N_2923,N_1900);
nor U5559 (N_5559,N_4898,N_1754);
xor U5560 (N_5560,N_1390,N_3592);
nand U5561 (N_5561,N_488,N_174);
and U5562 (N_5562,N_3051,N_3300);
and U5563 (N_5563,N_3417,N_1293);
nand U5564 (N_5564,N_4854,N_3265);
nand U5565 (N_5565,N_2712,N_4857);
and U5566 (N_5566,N_4113,N_997);
nor U5567 (N_5567,N_474,N_2472);
xor U5568 (N_5568,N_2842,N_4384);
or U5569 (N_5569,N_2956,N_2589);
and U5570 (N_5570,N_724,N_333);
nor U5571 (N_5571,N_3772,N_2077);
or U5572 (N_5572,N_1960,N_512);
xor U5573 (N_5573,N_268,N_3145);
and U5574 (N_5574,N_533,N_1419);
xor U5575 (N_5575,N_2336,N_4547);
or U5576 (N_5576,N_1973,N_4995);
or U5577 (N_5577,N_1967,N_3028);
nand U5578 (N_5578,N_3209,N_3227);
nand U5579 (N_5579,N_2137,N_4909);
and U5580 (N_5580,N_566,N_224);
and U5581 (N_5581,N_2578,N_4932);
nand U5582 (N_5582,N_949,N_4835);
nand U5583 (N_5583,N_596,N_4254);
or U5584 (N_5584,N_768,N_3050);
xnor U5585 (N_5585,N_667,N_3614);
or U5586 (N_5586,N_3133,N_962);
or U5587 (N_5587,N_4658,N_1587);
and U5588 (N_5588,N_426,N_3041);
or U5589 (N_5589,N_789,N_4936);
and U5590 (N_5590,N_2110,N_4531);
or U5591 (N_5591,N_2692,N_110);
nor U5592 (N_5592,N_1481,N_1041);
or U5593 (N_5593,N_3040,N_4848);
nand U5594 (N_5594,N_1760,N_3306);
or U5595 (N_5595,N_852,N_1618);
and U5596 (N_5596,N_3444,N_3138);
and U5597 (N_5597,N_4767,N_4094);
and U5598 (N_5598,N_617,N_4079);
nand U5599 (N_5599,N_829,N_4483);
and U5600 (N_5600,N_2329,N_1127);
or U5601 (N_5601,N_4560,N_1397);
or U5602 (N_5602,N_758,N_4927);
or U5603 (N_5603,N_2570,N_2756);
nor U5604 (N_5604,N_1452,N_2501);
or U5605 (N_5605,N_2917,N_4272);
or U5606 (N_5606,N_4170,N_497);
nand U5607 (N_5607,N_2152,N_4773);
nand U5608 (N_5608,N_1769,N_933);
nor U5609 (N_5609,N_2015,N_336);
xor U5610 (N_5610,N_134,N_2032);
and U5611 (N_5611,N_4670,N_4730);
nor U5612 (N_5612,N_3999,N_3789);
xnor U5613 (N_5613,N_3846,N_484);
or U5614 (N_5614,N_3446,N_2277);
nand U5615 (N_5615,N_837,N_4390);
and U5616 (N_5616,N_2213,N_407);
nand U5617 (N_5617,N_3543,N_352);
and U5618 (N_5618,N_587,N_4139);
or U5619 (N_5619,N_2123,N_2716);
nor U5620 (N_5620,N_3504,N_4629);
or U5621 (N_5621,N_4322,N_66);
and U5622 (N_5622,N_2770,N_4477);
and U5623 (N_5623,N_3296,N_592);
or U5624 (N_5624,N_1830,N_2976);
nor U5625 (N_5625,N_4540,N_2857);
nor U5626 (N_5626,N_1392,N_3241);
nand U5627 (N_5627,N_4574,N_162);
xnor U5628 (N_5628,N_4943,N_593);
nand U5629 (N_5629,N_107,N_3862);
or U5630 (N_5630,N_4023,N_2452);
nor U5631 (N_5631,N_4231,N_1064);
nand U5632 (N_5632,N_3738,N_2241);
nor U5633 (N_5633,N_604,N_4510);
and U5634 (N_5634,N_3190,N_1458);
or U5635 (N_5635,N_1265,N_4706);
or U5636 (N_5636,N_3416,N_4897);
nor U5637 (N_5637,N_385,N_3726);
nand U5638 (N_5638,N_822,N_294);
nand U5639 (N_5639,N_1662,N_230);
nor U5640 (N_5640,N_3657,N_4434);
nand U5641 (N_5641,N_4980,N_4904);
and U5642 (N_5642,N_930,N_750);
nor U5643 (N_5643,N_2547,N_844);
or U5644 (N_5644,N_327,N_2867);
and U5645 (N_5645,N_1161,N_4565);
xnor U5646 (N_5646,N_4827,N_4752);
and U5647 (N_5647,N_2475,N_1352);
and U5648 (N_5648,N_4869,N_1196);
nand U5649 (N_5649,N_476,N_4716);
or U5650 (N_5650,N_186,N_909);
nand U5651 (N_5651,N_3486,N_4705);
and U5652 (N_5652,N_1753,N_1150);
nand U5653 (N_5653,N_2492,N_3507);
xnor U5654 (N_5654,N_559,N_820);
or U5655 (N_5655,N_4425,N_3961);
or U5656 (N_5656,N_4176,N_4367);
and U5657 (N_5657,N_4299,N_4669);
and U5658 (N_5658,N_415,N_328);
nor U5659 (N_5659,N_3914,N_2485);
nor U5660 (N_5660,N_4268,N_1013);
and U5661 (N_5661,N_1829,N_547);
nand U5662 (N_5662,N_51,N_1660);
and U5663 (N_5663,N_1981,N_3441);
and U5664 (N_5664,N_3755,N_1066);
and U5665 (N_5665,N_2302,N_1263);
and U5666 (N_5666,N_2928,N_3719);
nor U5667 (N_5667,N_4006,N_89);
nor U5668 (N_5668,N_1047,N_4822);
nand U5669 (N_5669,N_2675,N_3231);
or U5670 (N_5670,N_3114,N_478);
and U5671 (N_5671,N_2043,N_111);
nand U5672 (N_5672,N_3567,N_2624);
nand U5673 (N_5673,N_825,N_2751);
nor U5674 (N_5674,N_4867,N_4015);
nand U5675 (N_5675,N_62,N_4899);
and U5676 (N_5676,N_2816,N_4186);
nand U5677 (N_5677,N_1355,N_79);
nand U5678 (N_5678,N_4933,N_1893);
or U5679 (N_5679,N_1004,N_2540);
nand U5680 (N_5680,N_1184,N_1050);
or U5681 (N_5681,N_3710,N_4269);
nor U5682 (N_5682,N_84,N_3063);
or U5683 (N_5683,N_2521,N_3);
xor U5684 (N_5684,N_4353,N_969);
and U5685 (N_5685,N_3348,N_4362);
nand U5686 (N_5686,N_1721,N_3037);
nor U5687 (N_5687,N_978,N_195);
nand U5688 (N_5688,N_1908,N_30);
nor U5689 (N_5689,N_3816,N_2256);
and U5690 (N_5690,N_1152,N_1107);
xnor U5691 (N_5691,N_1535,N_2240);
and U5692 (N_5692,N_3783,N_4057);
or U5693 (N_5693,N_4619,N_2557);
and U5694 (N_5694,N_1827,N_4189);
nand U5695 (N_5695,N_4505,N_365);
and U5696 (N_5696,N_3505,N_2430);
and U5697 (N_5697,N_2821,N_223);
nor U5698 (N_5698,N_4240,N_161);
and U5699 (N_5699,N_73,N_148);
nor U5700 (N_5700,N_2527,N_2993);
xor U5701 (N_5701,N_1565,N_1021);
or U5702 (N_5702,N_767,N_485);
nand U5703 (N_5703,N_2753,N_3148);
xnor U5704 (N_5704,N_2736,N_3681);
xor U5705 (N_5705,N_4021,N_4466);
nand U5706 (N_5706,N_4538,N_1564);
nand U5707 (N_5707,N_2254,N_603);
xnor U5708 (N_5708,N_3839,N_3573);
nor U5709 (N_5709,N_4794,N_4066);
nor U5710 (N_5710,N_4591,N_1852);
nor U5711 (N_5711,N_1543,N_2631);
xnor U5712 (N_5712,N_1106,N_1599);
xnor U5713 (N_5713,N_1820,N_2125);
or U5714 (N_5714,N_3481,N_2182);
nor U5715 (N_5715,N_3434,N_4551);
nand U5716 (N_5716,N_398,N_4523);
and U5717 (N_5717,N_212,N_2327);
and U5718 (N_5718,N_0,N_1992);
nand U5719 (N_5719,N_4703,N_4060);
xor U5720 (N_5720,N_2616,N_1058);
nor U5721 (N_5721,N_1081,N_797);
nand U5722 (N_5722,N_884,N_2134);
nor U5723 (N_5723,N_3260,N_1625);
and U5724 (N_5724,N_695,N_3334);
nand U5725 (N_5725,N_3454,N_1451);
nor U5726 (N_5726,N_4022,N_4437);
and U5727 (N_5727,N_2596,N_3397);
or U5728 (N_5728,N_1467,N_286);
or U5729 (N_5729,N_1507,N_4411);
nand U5730 (N_5730,N_3863,N_1189);
nand U5731 (N_5731,N_3804,N_4922);
and U5732 (N_5732,N_4009,N_4501);
nor U5733 (N_5733,N_2506,N_3944);
and U5734 (N_5734,N_4224,N_3594);
nor U5735 (N_5735,N_1156,N_3391);
xor U5736 (N_5736,N_1033,N_4952);
nand U5737 (N_5737,N_4916,N_1653);
and U5738 (N_5738,N_4677,N_818);
and U5739 (N_5739,N_1430,N_1776);
and U5740 (N_5740,N_3627,N_4101);
or U5741 (N_5741,N_2708,N_1568);
or U5742 (N_5742,N_4970,N_3585);
and U5743 (N_5743,N_3099,N_737);
nand U5744 (N_5744,N_3473,N_2874);
nand U5745 (N_5745,N_2727,N_4807);
nand U5746 (N_5746,N_4955,N_1551);
nor U5747 (N_5747,N_660,N_2776);
and U5748 (N_5748,N_4796,N_1708);
nor U5749 (N_5749,N_1578,N_68);
nor U5750 (N_5750,N_682,N_2659);
nand U5751 (N_5751,N_833,N_4996);
or U5752 (N_5752,N_1077,N_3993);
xnor U5753 (N_5753,N_717,N_4756);
nor U5754 (N_5754,N_3166,N_2382);
xnor U5755 (N_5755,N_4966,N_661);
or U5756 (N_5756,N_3136,N_377);
nand U5757 (N_5757,N_811,N_1069);
and U5758 (N_5758,N_2621,N_2422);
and U5759 (N_5759,N_3092,N_3142);
or U5760 (N_5760,N_1063,N_3583);
and U5761 (N_5761,N_178,N_1665);
nand U5762 (N_5762,N_490,N_1250);
nand U5763 (N_5763,N_1659,N_2385);
nor U5764 (N_5764,N_3410,N_4350);
nor U5765 (N_5765,N_17,N_3408);
nand U5766 (N_5766,N_2149,N_630);
or U5767 (N_5767,N_400,N_3767);
nand U5768 (N_5768,N_1795,N_565);
and U5769 (N_5769,N_378,N_4236);
or U5770 (N_5770,N_628,N_4349);
and U5771 (N_5771,N_4533,N_452);
nand U5772 (N_5772,N_2883,N_2761);
nor U5773 (N_5773,N_2612,N_3778);
nor U5774 (N_5774,N_4910,N_3536);
or U5775 (N_5775,N_261,N_4467);
and U5776 (N_5776,N_3998,N_4883);
or U5777 (N_5777,N_1046,N_2403);
nand U5778 (N_5778,N_4684,N_3885);
nand U5779 (N_5779,N_1271,N_3125);
and U5780 (N_5780,N_3412,N_2155);
nand U5781 (N_5781,N_536,N_3091);
nand U5782 (N_5782,N_2463,N_1155);
or U5783 (N_5783,N_4311,N_1246);
nand U5784 (N_5784,N_2583,N_1837);
nor U5785 (N_5785,N_690,N_2132);
nor U5786 (N_5786,N_399,N_4630);
and U5787 (N_5787,N_1039,N_2503);
and U5788 (N_5788,N_455,N_2078);
nand U5789 (N_5789,N_4083,N_2070);
or U5790 (N_5790,N_4100,N_1763);
xor U5791 (N_5791,N_2467,N_4855);
nor U5792 (N_5792,N_537,N_2175);
nand U5793 (N_5793,N_376,N_714);
xnor U5794 (N_5794,N_2769,N_3197);
or U5795 (N_5795,N_1314,N_2293);
nand U5796 (N_5796,N_1363,N_1756);
nand U5797 (N_5797,N_3172,N_4645);
and U5798 (N_5798,N_2875,N_710);
or U5799 (N_5799,N_1984,N_1863);
and U5800 (N_5800,N_2811,N_3331);
xnor U5801 (N_5801,N_3552,N_3520);
xnor U5802 (N_5802,N_3208,N_3644);
xnor U5803 (N_5803,N_3584,N_4346);
or U5804 (N_5804,N_2286,N_2549);
nand U5805 (N_5805,N_3224,N_3307);
and U5806 (N_5806,N_405,N_1462);
nor U5807 (N_5807,N_4405,N_4881);
nor U5808 (N_5808,N_220,N_2176);
nor U5809 (N_5809,N_4161,N_3677);
xor U5810 (N_5810,N_2036,N_318);
and U5811 (N_5811,N_1607,N_3329);
nor U5812 (N_5812,N_1235,N_4175);
and U5813 (N_5813,N_3600,N_1300);
and U5814 (N_5814,N_2957,N_200);
nor U5815 (N_5815,N_2369,N_4971);
and U5816 (N_5816,N_1262,N_1685);
nand U5817 (N_5817,N_4597,N_4404);
nand U5818 (N_5818,N_2405,N_2113);
or U5819 (N_5819,N_3869,N_4575);
nand U5820 (N_5820,N_1483,N_1848);
nand U5821 (N_5821,N_3489,N_2919);
nand U5822 (N_5822,N_1464,N_3587);
nor U5823 (N_5823,N_1423,N_80);
or U5824 (N_5824,N_2903,N_2151);
or U5825 (N_5825,N_1575,N_4335);
and U5826 (N_5826,N_460,N_3928);
nand U5827 (N_5827,N_45,N_4476);
nor U5828 (N_5828,N_4124,N_2499);
nor U5829 (N_5829,N_88,N_772);
or U5830 (N_5830,N_2389,N_2807);
or U5831 (N_5831,N_2038,N_2512);
or U5832 (N_5832,N_2448,N_950);
or U5833 (N_5833,N_2688,N_3315);
nor U5834 (N_5834,N_4732,N_23);
nor U5835 (N_5835,N_1247,N_1253);
nor U5836 (N_5836,N_626,N_2383);
nand U5837 (N_5837,N_4678,N_1095);
nand U5838 (N_5838,N_1531,N_1841);
nand U5839 (N_5839,N_834,N_1256);
nand U5840 (N_5840,N_3061,N_1374);
nand U5841 (N_5841,N_778,N_226);
or U5842 (N_5842,N_2587,N_4429);
nand U5843 (N_5843,N_3911,N_140);
nor U5844 (N_5844,N_951,N_3316);
nand U5845 (N_5845,N_4832,N_3808);
and U5846 (N_5846,N_2236,N_401);
nor U5847 (N_5847,N_2737,N_1492);
nor U5848 (N_5848,N_4750,N_3689);
or U5849 (N_5849,N_3903,N_770);
xnor U5850 (N_5850,N_3447,N_3337);
nor U5851 (N_5851,N_549,N_1937);
and U5852 (N_5852,N_2345,N_1853);
or U5853 (N_5853,N_4086,N_3471);
nand U5854 (N_5854,N_1570,N_353);
nor U5855 (N_5855,N_4660,N_424);
or U5856 (N_5856,N_3345,N_3156);
and U5857 (N_5857,N_2819,N_1811);
and U5858 (N_5858,N_3060,N_4325);
nand U5859 (N_5859,N_1683,N_1990);
nand U5860 (N_5860,N_4391,N_473);
nor U5861 (N_5861,N_1200,N_4044);
nor U5862 (N_5862,N_2826,N_3854);
nor U5863 (N_5863,N_1016,N_3233);
nand U5864 (N_5864,N_591,N_3107);
or U5865 (N_5865,N_3511,N_4085);
or U5866 (N_5866,N_4838,N_1779);
or U5867 (N_5867,N_146,N_3760);
and U5868 (N_5868,N_3344,N_4081);
nand U5869 (N_5869,N_1901,N_673);
and U5870 (N_5870,N_306,N_1891);
xor U5871 (N_5871,N_4187,N_1484);
and U5872 (N_5872,N_4978,N_27);
or U5873 (N_5873,N_4122,N_2838);
nand U5874 (N_5874,N_3576,N_4191);
or U5875 (N_5875,N_2667,N_3769);
and U5876 (N_5876,N_4174,N_4407);
or U5877 (N_5877,N_1712,N_1134);
xor U5878 (N_5878,N_4913,N_1428);
and U5879 (N_5879,N_118,N_4571);
or U5880 (N_5880,N_3181,N_4296);
and U5881 (N_5881,N_4210,N_4281);
or U5882 (N_5882,N_595,N_131);
or U5883 (N_5883,N_3612,N_2892);
or U5884 (N_5884,N_4337,N_546);
and U5885 (N_5885,N_3496,N_2268);
and U5886 (N_5886,N_2526,N_203);
or U5887 (N_5887,N_3349,N_3442);
nand U5888 (N_5888,N_3118,N_4557);
and U5889 (N_5889,N_3642,N_3319);
nor U5890 (N_5890,N_3963,N_4831);
nand U5891 (N_5891,N_1865,N_2233);
and U5892 (N_5892,N_3178,N_4331);
nor U5893 (N_5893,N_2744,N_2646);
nand U5894 (N_5894,N_3022,N_4521);
nand U5895 (N_5895,N_528,N_4930);
nor U5896 (N_5896,N_2407,N_3604);
nor U5897 (N_5897,N_3309,N_3380);
nand U5898 (N_5898,N_1844,N_4546);
nor U5899 (N_5899,N_910,N_1097);
nor U5900 (N_5900,N_2136,N_2607);
nor U5901 (N_5901,N_4105,N_2228);
nor U5902 (N_5902,N_643,N_1548);
nand U5903 (N_5903,N_4661,N_1193);
nor U5904 (N_5904,N_1773,N_341);
nor U5905 (N_5905,N_3124,N_1198);
xnor U5906 (N_5906,N_3683,N_1488);
or U5907 (N_5907,N_1169,N_3691);
xor U5908 (N_5908,N_1259,N_4534);
and U5909 (N_5909,N_1221,N_3758);
and U5910 (N_5910,N_459,N_4065);
or U5911 (N_5911,N_511,N_2387);
nand U5912 (N_5912,N_3485,N_2998);
or U5913 (N_5913,N_1298,N_1494);
xor U5914 (N_5914,N_3817,N_4201);
and U5915 (N_5915,N_2661,N_228);
and U5916 (N_5916,N_3730,N_1668);
nand U5917 (N_5917,N_81,N_906);
nand U5918 (N_5918,N_2150,N_3969);
nor U5919 (N_5919,N_882,N_321);
nand U5920 (N_5920,N_1251,N_208);
and U5921 (N_5921,N_2347,N_1213);
and U5922 (N_5922,N_3013,N_1593);
nor U5923 (N_5923,N_144,N_3791);
nor U5924 (N_5924,N_3382,N_4514);
nor U5925 (N_5925,N_120,N_1735);
nor U5926 (N_5926,N_2494,N_2342);
and U5927 (N_5927,N_3189,N_4452);
nand U5928 (N_5928,N_2352,N_4589);
nor U5929 (N_5929,N_242,N_2629);
nand U5930 (N_5930,N_2480,N_404);
and U5931 (N_5931,N_4027,N_4492);
nor U5932 (N_5932,N_330,N_762);
or U5933 (N_5933,N_4225,N_83);
and U5934 (N_5934,N_1112,N_1277);
xnor U5935 (N_5935,N_2471,N_2795);
xnor U5936 (N_5936,N_986,N_1502);
nor U5937 (N_5937,N_3182,N_59);
nand U5938 (N_5938,N_2204,N_213);
nand U5939 (N_5939,N_4493,N_539);
xnor U5940 (N_5940,N_1782,N_746);
nor U5941 (N_5941,N_879,N_996);
nand U5942 (N_5942,N_572,N_964);
and U5943 (N_5943,N_632,N_3786);
and U5944 (N_5944,N_4146,N_2534);
and U5945 (N_5945,N_449,N_3659);
nor U5946 (N_5946,N_251,N_3154);
xor U5947 (N_5947,N_4343,N_836);
nor U5948 (N_5948,N_4398,N_570);
nor U5949 (N_5949,N_360,N_1979);
nor U5950 (N_5950,N_1918,N_3347);
nand U5951 (N_5951,N_2974,N_2615);
nand U5952 (N_5952,N_4295,N_3457);
or U5953 (N_5953,N_4894,N_552);
nor U5954 (N_5954,N_3897,N_4844);
and U5955 (N_5955,N_3221,N_2035);
nand U5956 (N_5956,N_3826,N_2970);
and U5957 (N_5957,N_4247,N_1996);
or U5958 (N_5958,N_4873,N_3488);
nor U5959 (N_5959,N_2754,N_692);
and U5960 (N_5960,N_4965,N_672);
nand U5961 (N_5961,N_4206,N_3393);
xor U5962 (N_5962,N_2742,N_1895);
nand U5963 (N_5963,N_3360,N_703);
and U5964 (N_5964,N_1056,N_3521);
xor U5965 (N_5965,N_2420,N_888);
xnor U5966 (N_5966,N_4786,N_2164);
nor U5967 (N_5967,N_2725,N_3537);
nand U5968 (N_5968,N_4173,N_3915);
nor U5969 (N_5969,N_1917,N_804);
and U5970 (N_5970,N_4622,N_3983);
nor U5971 (N_5971,N_3848,N_3724);
xor U5972 (N_5972,N_4037,N_4506);
or U5973 (N_5973,N_3213,N_786);
or U5974 (N_5974,N_4843,N_2016);
nand U5975 (N_5975,N_2562,N_1375);
nand U5976 (N_5976,N_3981,N_137);
nand U5977 (N_5977,N_1864,N_3680);
or U5978 (N_5978,N_4717,N_406);
nor U5979 (N_5979,N_3104,N_2332);
or U5980 (N_5980,N_2674,N_783);
nand U5981 (N_5981,N_560,N_991);
nor U5982 (N_5982,N_3990,N_4797);
and U5983 (N_5983,N_2937,N_1216);
nand U5984 (N_5984,N_4267,N_594);
or U5985 (N_5985,N_3325,N_914);
and U5986 (N_5986,N_154,N_4691);
xor U5987 (N_5987,N_1646,N_4378);
and U5988 (N_5988,N_899,N_937);
and U5989 (N_5989,N_4707,N_1588);
nand U5990 (N_5990,N_863,N_3418);
nor U5991 (N_5991,N_2679,N_1372);
xnor U5992 (N_5992,N_433,N_2235);
nand U5993 (N_5993,N_43,N_1822);
or U5994 (N_5994,N_2996,N_364);
nand U5995 (N_5995,N_4324,N_1160);
nor U5996 (N_5996,N_4882,N_335);
and U5997 (N_5997,N_160,N_2988);
and U5998 (N_5998,N_4341,N_1931);
nor U5999 (N_5999,N_612,N_3362);
or U6000 (N_6000,N_4077,N_2331);
or U6001 (N_6001,N_621,N_4612);
or U6002 (N_6002,N_4724,N_3770);
and U6003 (N_6003,N_37,N_880);
xor U6004 (N_6004,N_446,N_1126);
and U6005 (N_6005,N_616,N_922);
or U6006 (N_6006,N_4604,N_2894);
and U6007 (N_6007,N_845,N_1283);
nor U6008 (N_6008,N_3076,N_4851);
xnor U6009 (N_6009,N_3987,N_1942);
or U6010 (N_6010,N_2680,N_734);
or U6011 (N_6011,N_955,N_3798);
nand U6012 (N_6012,N_2415,N_957);
nor U6013 (N_6013,N_3183,N_3841);
or U6014 (N_6014,N_3255,N_3776);
nor U6015 (N_6015,N_2445,N_403);
and U6016 (N_6016,N_1858,N_3093);
nor U6017 (N_6017,N_1425,N_1630);
nor U6018 (N_6018,N_2099,N_881);
nand U6019 (N_6019,N_3487,N_3849);
or U6020 (N_6020,N_4960,N_4776);
xor U6021 (N_6021,N_4007,N_868);
and U6022 (N_6022,N_198,N_4109);
and U6023 (N_6023,N_1624,N_948);
nor U6024 (N_6024,N_2948,N_123);
nand U6025 (N_6025,N_4266,N_1638);
nand U6026 (N_6026,N_516,N_1120);
nor U6027 (N_6027,N_1566,N_954);
nor U6028 (N_6028,N_3696,N_3806);
xnor U6029 (N_6029,N_4484,N_2967);
nand U6030 (N_6030,N_1813,N_3626);
and U6031 (N_6031,N_4676,N_4537);
nor U6032 (N_6032,N_3376,N_4447);
and U6033 (N_6033,N_3455,N_4298);
and U6034 (N_6034,N_2582,N_4091);
or U6035 (N_6035,N_2603,N_1470);
nand U6036 (N_6036,N_2489,N_3618);
nor U6037 (N_6037,N_4326,N_1143);
nand U6038 (N_6038,N_3978,N_1498);
nor U6039 (N_6039,N_2870,N_827);
nand U6040 (N_6040,N_3876,N_2260);
and U6041 (N_6041,N_475,N_3796);
and U6042 (N_6042,N_2935,N_3460);
and U6043 (N_6043,N_1629,N_202);
and U6044 (N_6044,N_4169,N_4451);
nor U6045 (N_6045,N_1103,N_1540);
or U6046 (N_6046,N_3889,N_3860);
nor U6047 (N_6047,N_2172,N_3548);
or U6048 (N_6048,N_1245,N_3967);
nor U6049 (N_6049,N_3956,N_2425);
or U6050 (N_6050,N_3343,N_1762);
nand U6051 (N_6051,N_3082,N_1384);
nand U6052 (N_6052,N_4785,N_1116);
and U6053 (N_6053,N_4866,N_3267);
and U6054 (N_6054,N_4673,N_2454);
or U6055 (N_6055,N_510,N_3785);
or U6056 (N_6056,N_2173,N_988);
and U6057 (N_6057,N_525,N_1920);
and U6058 (N_6058,N_538,N_3704);
and U6059 (N_6059,N_450,N_4159);
nand U6060 (N_6060,N_1651,N_1209);
nor U6061 (N_6061,N_4653,N_3134);
xor U6062 (N_6062,N_4198,N_4569);
or U6063 (N_6063,N_1242,N_383);
xor U6064 (N_6064,N_3008,N_2059);
and U6065 (N_6065,N_967,N_1924);
nand U6066 (N_6066,N_3672,N_3339);
xnor U6067 (N_6067,N_2995,N_4628);
or U6068 (N_6068,N_2556,N_2084);
and U6069 (N_6069,N_807,N_2381);
and U6070 (N_6070,N_2801,N_1386);
or U6071 (N_6071,N_4314,N_4561);
or U6072 (N_6072,N_2288,N_2953);
and U6073 (N_6073,N_2726,N_3740);
nand U6074 (N_6074,N_4380,N_100);
nand U6075 (N_6075,N_3748,N_285);
nand U6076 (N_6076,N_70,N_1890);
nor U6077 (N_6077,N_3763,N_668);
nand U6078 (N_6078,N_1154,N_2311);
nor U6079 (N_6079,N_3595,N_1930);
nand U6080 (N_6080,N_590,N_2649);
nand U6081 (N_6081,N_2595,N_2129);
nand U6082 (N_6082,N_2986,N_4489);
nand U6083 (N_6083,N_3158,N_4366);
xor U6084 (N_6084,N_1131,N_2735);
or U6085 (N_6085,N_2147,N_3177);
nor U6086 (N_6086,N_480,N_2392);
or U6087 (N_6087,N_295,N_3952);
nor U6088 (N_6088,N_4163,N_3494);
nand U6089 (N_6089,N_3069,N_3574);
and U6090 (N_6090,N_4594,N_4018);
nand U6091 (N_6091,N_4422,N_2610);
and U6092 (N_6092,N_1086,N_2441);
and U6093 (N_6093,N_934,N_4544);
and U6094 (N_6094,N_1000,N_1296);
nor U6095 (N_6095,N_1585,N_2672);
nand U6096 (N_6096,N_3113,N_1179);
nand U6097 (N_6097,N_2030,N_2693);
or U6098 (N_6098,N_2115,N_3246);
nand U6099 (N_6099,N_885,N_172);
nand U6100 (N_6100,N_3143,N_2729);
nor U6101 (N_6101,N_3739,N_2456);
or U6102 (N_6102,N_1983,N_1946);
nand U6103 (N_6103,N_4562,N_4446);
and U6104 (N_6104,N_2300,N_2888);
and U6105 (N_6105,N_793,N_1928);
or U6106 (N_6106,N_4602,N_4739);
or U6107 (N_6107,N_4131,N_2710);
and U6108 (N_6108,N_4621,N_4609);
and U6109 (N_6109,N_2728,N_3620);
xor U6110 (N_6110,N_494,N_4994);
and U6111 (N_6111,N_4743,N_1965);
nor U6112 (N_6112,N_2190,N_3801);
nand U6113 (N_6113,N_4517,N_2747);
or U6114 (N_6114,N_4443,N_4572);
and U6115 (N_6115,N_1007,N_4357);
and U6116 (N_6116,N_4636,N_2739);
nand U6117 (N_6117,N_941,N_3185);
and U6118 (N_6118,N_3352,N_3144);
nand U6119 (N_6119,N_1174,N_2802);
nor U6120 (N_6120,N_3110,N_2273);
and U6121 (N_6121,N_2955,N_4803);
and U6122 (N_6122,N_1597,N_4249);
xor U6123 (N_6123,N_2555,N_2965);
nor U6124 (N_6124,N_4499,N_3697);
and U6125 (N_6125,N_3972,N_3538);
nor U6126 (N_6126,N_1964,N_850);
and U6127 (N_6127,N_3799,N_3893);
and U6128 (N_6128,N_2809,N_841);
or U6129 (N_6129,N_2192,N_2466);
nor U6130 (N_6130,N_2429,N_2940);
nor U6131 (N_6131,N_777,N_244);
and U6132 (N_6132,N_4507,N_2320);
nand U6133 (N_6133,N_1602,N_164);
nand U6134 (N_6134,N_2031,N_2275);
or U6135 (N_6135,N_3286,N_4312);
xnor U6136 (N_6136,N_1206,N_1652);
and U6137 (N_6137,N_1909,N_1036);
xor U6138 (N_6138,N_1083,N_3701);
and U6139 (N_6139,N_4214,N_2546);
nand U6140 (N_6140,N_663,N_3282);
or U6141 (N_6141,N_4072,N_2984);
or U6142 (N_6142,N_1679,N_409);
nor U6143 (N_6143,N_4119,N_1299);
and U6144 (N_6144,N_4270,N_605);
xor U6145 (N_6145,N_453,N_3551);
or U6146 (N_6146,N_2542,N_180);
nor U6147 (N_6147,N_4600,N_4675);
or U6148 (N_6148,N_3258,N_2921);
nand U6149 (N_6149,N_2997,N_1219);
nor U6150 (N_6150,N_2262,N_1707);
and U6151 (N_6151,N_2060,N_2845);
or U6152 (N_6152,N_1024,N_3510);
and U6153 (N_6153,N_2105,N_795);
xnor U6154 (N_6154,N_347,N_1197);
and U6155 (N_6155,N_77,N_2442);
nand U6156 (N_6156,N_618,N_739);
nand U6157 (N_6157,N_4962,N_995);
nor U6158 (N_6158,N_2681,N_4957);
or U6159 (N_6159,N_2664,N_1140);
nor U6160 (N_6160,N_3364,N_6);
and U6161 (N_6161,N_4526,N_3033);
xor U6162 (N_6162,N_1734,N_3399);
xnor U6163 (N_6163,N_7,N_802);
nor U6164 (N_6164,N_3052,N_2160);
and U6165 (N_6165,N_4833,N_1022);
and U6166 (N_6166,N_3005,N_3751);
xor U6167 (N_6167,N_4799,N_355);
or U6168 (N_6168,N_4014,N_1306);
nor U6169 (N_6169,N_1557,N_2927);
nor U6170 (N_6170,N_3132,N_3305);
xnor U6171 (N_6171,N_3029,N_2292);
or U6172 (N_6172,N_3355,N_4409);
xnor U6173 (N_6173,N_4013,N_4042);
nor U6174 (N_6174,N_556,N_1159);
and U6175 (N_6175,N_1643,N_173);
nor U6176 (N_6176,N_1922,N_1485);
and U6177 (N_6177,N_4986,N_1172);
and U6178 (N_6178,N_2181,N_1109);
or U6179 (N_6179,N_4769,N_1098);
or U6180 (N_6180,N_1910,N_4570);
nand U6181 (N_6181,N_2284,N_4403);
xnor U6182 (N_6182,N_4979,N_578);
or U6183 (N_6183,N_4260,N_4813);
and U6184 (N_6184,N_831,N_4416);
nand U6185 (N_6185,N_1913,N_1874);
or U6186 (N_6186,N_4067,N_1586);
and U6187 (N_6187,N_3640,N_521);
nor U6188 (N_6188,N_413,N_606);
or U6189 (N_6189,N_2244,N_905);
or U6190 (N_6190,N_2504,N_4045);
nand U6191 (N_6191,N_1340,N_4290);
or U6192 (N_6192,N_3367,N_392);
nor U6193 (N_6193,N_1,N_1826);
and U6194 (N_6194,N_1923,N_1437);
and U6195 (N_6195,N_1759,N_4474);
nor U6196 (N_6196,N_1701,N_2914);
nor U6197 (N_6197,N_1700,N_2295);
nand U6198 (N_6198,N_4698,N_2153);
nand U6199 (N_6199,N_588,N_3065);
nand U6200 (N_6200,N_764,N_4286);
nor U6201 (N_6201,N_913,N_1426);
or U6202 (N_6202,N_928,N_2622);
xor U6203 (N_6203,N_4160,N_1934);
and U6204 (N_6204,N_2139,N_685);
or U6205 (N_6205,N_2911,N_2896);
nand U6206 (N_6206,N_1377,N_2161);
nand U6207 (N_6207,N_743,N_4396);
or U6208 (N_6208,N_1514,N_987);
or U6209 (N_6209,N_2447,N_4024);
and U6210 (N_6210,N_4089,N_1449);
or U6211 (N_6211,N_2465,N_1899);
or U6212 (N_6212,N_1921,N_1059);
nand U6213 (N_6213,N_4468,N_4755);
and U6214 (N_6214,N_1988,N_4634);
and U6215 (N_6215,N_3523,N_2938);
xor U6216 (N_6216,N_541,N_1698);
nand U6217 (N_6217,N_2307,N_501);
nor U6218 (N_6218,N_4742,N_3609);
nand U6219 (N_6219,N_2304,N_932);
or U6220 (N_6220,N_3167,N_898);
nand U6221 (N_6221,N_4048,N_395);
xor U6222 (N_6222,N_1611,N_1501);
and U6223 (N_6223,N_812,N_1412);
or U6224 (N_6224,N_4862,N_3240);
nor U6225 (N_6225,N_1124,N_1096);
or U6226 (N_6226,N_1888,N_4342);
nor U6227 (N_6227,N_2498,N_4076);
and U6228 (N_6228,N_3765,N_1319);
xnor U6229 (N_6229,N_1847,N_1628);
xor U6230 (N_6230,N_3533,N_2315);
nand U6231 (N_6231,N_3160,N_2835);
xor U6232 (N_6232,N_1288,N_1581);
xnor U6233 (N_6233,N_3588,N_2969);
and U6234 (N_6234,N_1859,N_3831);
nor U6235 (N_6235,N_670,N_2925);
nand U6236 (N_6236,N_1266,N_1948);
nand U6237 (N_6237,N_4473,N_4220);
or U6238 (N_6238,N_1539,N_2538);
nand U6239 (N_6239,N_96,N_1592);
and U6240 (N_6240,N_4354,N_1941);
or U6241 (N_6241,N_442,N_1211);
and U6242 (N_6242,N_921,N_2362);
or U6243 (N_6243,N_393,N_2398);
or U6244 (N_6244,N_4226,N_2251);
nand U6245 (N_6245,N_3120,N_3312);
xnor U6246 (N_6246,N_279,N_4543);
nor U6247 (N_6247,N_36,N_4287);
and U6248 (N_6248,N_3211,N_3895);
xor U6249 (N_6249,N_4879,N_2368);
nor U6250 (N_6250,N_873,N_3924);
xnor U6251 (N_6251,N_165,N_4274);
nand U6252 (N_6252,N_712,N_779);
nand U6253 (N_6253,N_3966,N_886);
nor U6254 (N_6254,N_2724,N_421);
nor U6255 (N_6255,N_4737,N_3902);
and U6256 (N_6256,N_1252,N_1766);
nor U6257 (N_6257,N_4530,N_4795);
and U6258 (N_6258,N_243,N_1114);
and U6259 (N_6259,N_2230,N_3753);
or U6260 (N_6260,N_2567,N_15);
or U6261 (N_6261,N_3159,N_3245);
nor U6262 (N_6262,N_2690,N_1167);
nor U6263 (N_6263,N_386,N_2847);
nand U6264 (N_6264,N_1403,N_975);
nor U6265 (N_6265,N_3193,N_861);
xor U6266 (N_6266,N_2162,N_1634);
nor U6267 (N_6267,N_1468,N_2529);
and U6268 (N_6268,N_3311,N_1576);
nand U6269 (N_6269,N_170,N_1876);
nand U6270 (N_6270,N_3997,N_4455);
or U6271 (N_6271,N_577,N_4853);
and U6272 (N_6272,N_2108,N_2280);
nand U6273 (N_6273,N_3402,N_4415);
or U6274 (N_6274,N_2946,N_1699);
nand U6275 (N_6275,N_3861,N_2025);
and U6276 (N_6276,N_2272,N_702);
and U6277 (N_6277,N_4856,N_3127);
or U6278 (N_6278,N_3941,N_163);
or U6279 (N_6279,N_2029,N_4212);
or U6280 (N_6280,N_1459,N_2484);
nand U6281 (N_6281,N_2438,N_4017);
nand U6282 (N_6282,N_16,N_215);
nand U6283 (N_6283,N_1616,N_2698);
nor U6284 (N_6284,N_4941,N_2048);
or U6285 (N_6285,N_938,N_4908);
or U6286 (N_6286,N_1733,N_4369);
nand U6287 (N_6287,N_1201,N_2650);
nor U6288 (N_6288,N_2633,N_3692);
nor U6289 (N_6289,N_3616,N_1455);
and U6290 (N_6290,N_2326,N_4195);
nor U6291 (N_6291,N_308,N_3026);
or U6292 (N_6292,N_3636,N_3248);
nor U6293 (N_6293,N_4642,N_821);
and U6294 (N_6294,N_3400,N_3163);
or U6295 (N_6295,N_3908,N_3807);
and U6296 (N_6296,N_1614,N_4330);
nand U6297 (N_6297,N_1806,N_1139);
and U6298 (N_6298,N_3232,N_1440);
and U6299 (N_6299,N_2748,N_1142);
and U6300 (N_6300,N_3047,N_719);
or U6301 (N_6301,N_2253,N_531);
nand U6302 (N_6302,N_2177,N_4614);
nor U6303 (N_6303,N_4738,N_3832);
and U6304 (N_6304,N_715,N_2594);
nand U6305 (N_6305,N_2803,N_1870);
xnor U6306 (N_6306,N_1023,N_2062);
nand U6307 (N_6307,N_2889,N_4262);
nor U6308 (N_6308,N_1862,N_4792);
or U6309 (N_6309,N_4178,N_1473);
nor U6310 (N_6310,N_1861,N_2140);
nor U6311 (N_6311,N_2723,N_2167);
and U6312 (N_6312,N_562,N_4963);
nand U6313 (N_6313,N_3064,N_4392);
and U6314 (N_6314,N_4584,N_2992);
nor U6315 (N_6315,N_4423,N_117);
and U6316 (N_6316,N_524,N_4308);
and U6317 (N_6317,N_2270,N_417);
and U6318 (N_6318,N_3695,N_1005);
or U6319 (N_6319,N_925,N_3813);
xor U6320 (N_6320,N_1730,N_3712);
or U6321 (N_6321,N_581,N_2374);
or U6322 (N_6322,N_4132,N_907);
nor U6323 (N_6323,N_741,N_1075);
xor U6324 (N_6324,N_3707,N_1236);
xor U6325 (N_6325,N_464,N_4328);
nand U6326 (N_6326,N_3820,N_315);
nor U6327 (N_6327,N_792,N_1871);
or U6328 (N_6328,N_1224,N_4112);
nor U6329 (N_6329,N_892,N_3641);
or U6330 (N_6330,N_3840,N_3155);
and U6331 (N_6331,N_4620,N_3086);
nand U6332 (N_6332,N_4884,N_1227);
or U6333 (N_6333,N_3630,N_1845);
nor U6334 (N_6334,N_854,N_4234);
nand U6335 (N_6335,N_53,N_2412);
nand U6336 (N_6336,N_1819,N_91);
or U6337 (N_6337,N_2532,N_354);
nor U6338 (N_6338,N_3873,N_1856);
nor U6339 (N_6339,N_1220,N_2019);
or U6340 (N_6340,N_4981,N_4208);
xor U6341 (N_6341,N_2536,N_4836);
nor U6342 (N_6342,N_3528,N_4472);
xor U6343 (N_6343,N_4096,N_3075);
nand U6344 (N_6344,N_301,N_263);
and U6345 (N_6345,N_1866,N_1092);
nand U6346 (N_6346,N_2205,N_1952);
and U6347 (N_6347,N_1621,N_468);
nand U6348 (N_6348,N_4251,N_4120);
nand U6349 (N_6349,N_4817,N_2685);
or U6350 (N_6350,N_4582,N_4135);
nand U6351 (N_6351,N_3474,N_1803);
nor U6352 (N_6352,N_760,N_840);
or U6353 (N_6353,N_1380,N_2287);
nand U6354 (N_6354,N_2246,N_3323);
and U6355 (N_6355,N_2559,N_4386);
or U6356 (N_6356,N_2343,N_3768);
nand U6357 (N_6357,N_919,N_1282);
nand U6358 (N_6358,N_4406,N_2618);
or U6359 (N_6359,N_729,N_1770);
and U6360 (N_6360,N_3851,N_1739);
nor U6361 (N_6361,N_1324,N_1032);
or U6362 (N_6362,N_4363,N_4417);
and U6363 (N_6363,N_3015,N_3036);
or U6364 (N_6364,N_2837,N_790);
or U6365 (N_6365,N_2432,N_396);
nand U6366 (N_6366,N_1765,N_1279);
or U6367 (N_6367,N_3901,N_4859);
nand U6368 (N_6368,N_2298,N_1573);
or U6369 (N_6369,N_4734,N_4088);
nand U6370 (N_6370,N_761,N_1894);
nand U6371 (N_6371,N_3621,N_1170);
nand U6372 (N_6372,N_4956,N_4781);
or U6373 (N_6373,N_3039,N_2095);
or U6374 (N_6374,N_4313,N_781);
nand U6375 (N_6375,N_1448,N_4408);
nor U6376 (N_6376,N_1212,N_1747);
nand U6377 (N_6377,N_4722,N_3645);
xnor U6378 (N_6378,N_350,N_4292);
nand U6379 (N_6379,N_1304,N_3582);
nor U6380 (N_6380,N_1230,N_1311);
nand U6381 (N_6381,N_4194,N_2126);
and U6382 (N_6382,N_2168,N_2643);
or U6383 (N_6383,N_4793,N_2044);
and U6384 (N_6384,N_4168,N_2832);
nor U6385 (N_6385,N_3175,N_583);
nand U6386 (N_6386,N_3292,N_2247);
and U6387 (N_6387,N_4227,N_1225);
and U6388 (N_6388,N_720,N_649);
nand U6389 (N_6389,N_1215,N_281);
xnor U6390 (N_6390,N_1264,N_4638);
or U6391 (N_6391,N_3396,N_3943);
or U6392 (N_6392,N_3667,N_2565);
and U6393 (N_6393,N_2813,N_1672);
nor U6394 (N_6394,N_4394,N_2859);
nand U6395 (N_6395,N_1476,N_3926);
and U6396 (N_6396,N_4681,N_1082);
and U6397 (N_6397,N_1647,N_3302);
xnor U6398 (N_6398,N_4185,N_1574);
or U6399 (N_6399,N_2789,N_1818);
and U6400 (N_6400,N_2605,N_259);
and U6401 (N_6401,N_4156,N_952);
nor U6402 (N_6402,N_297,N_3575);
and U6403 (N_6403,N_3878,N_1187);
nor U6404 (N_6404,N_2079,N_3942);
xnor U6405 (N_6405,N_343,N_3809);
nor U6406 (N_6406,N_2358,N_4808);
nor U6407 (N_6407,N_1555,N_2943);
or U6408 (N_6408,N_2878,N_2636);
nor U6409 (N_6409,N_3326,N_2981);
nand U6410 (N_6410,N_2232,N_1626);
nand U6411 (N_6411,N_1787,N_519);
or U6412 (N_6412,N_2166,N_3646);
nor U6413 (N_6413,N_3547,N_2020);
xnor U6414 (N_6414,N_4829,N_337);
or U6415 (N_6415,N_2148,N_41);
and U6416 (N_6416,N_351,N_2450);
nand U6417 (N_6417,N_2296,N_766);
nand U6418 (N_6418,N_2625,N_4701);
and U6419 (N_6419,N_348,N_326);
and U6420 (N_6420,N_2922,N_272);
nor U6421 (N_6421,N_388,N_3628);
nand U6422 (N_6422,N_1750,N_49);
or U6423 (N_6423,N_4126,N_3923);
nor U6424 (N_6424,N_1421,N_2451);
nor U6425 (N_6425,N_1675,N_3912);
and U6426 (N_6426,N_1567,N_2022);
nand U6427 (N_6427,N_1117,N_3373);
or U6428 (N_6428,N_1465,N_1270);
xnor U6429 (N_6429,N_4500,N_3500);
and U6430 (N_6430,N_4931,N_1999);
and U6431 (N_6431,N_3829,N_3669);
xor U6432 (N_6432,N_2913,N_4049);
and U6433 (N_6433,N_197,N_611);
nor U6434 (N_6434,N_1892,N_2092);
nor U6435 (N_6435,N_448,N_3283);
nand U6436 (N_6436,N_2428,N_2592);
nand U6437 (N_6437,N_677,N_3649);
nor U6438 (N_6438,N_4811,N_3666);
and U6439 (N_6439,N_3519,N_633);
nand U6440 (N_6440,N_4651,N_4845);
and U6441 (N_6441,N_1966,N_3919);
or U6442 (N_6442,N_4445,N_4950);
or U6443 (N_6443,N_1471,N_1755);
nor U6444 (N_6444,N_1317,N_1410);
nor U6445 (N_6445,N_1030,N_2671);
nor U6446 (N_6446,N_1178,N_1812);
nand U6447 (N_6447,N_2617,N_3540);
nand U6448 (N_6448,N_1349,N_3544);
xor U6449 (N_6449,N_2341,N_953);
and U6450 (N_6450,N_2339,N_1998);
and U6451 (N_6451,N_4959,N_3513);
nand U6452 (N_6452,N_567,N_3478);
or U6453 (N_6453,N_324,N_1373);
xnor U6454 (N_6454,N_4239,N_1801);
and U6455 (N_6455,N_1325,N_2910);
or U6456 (N_6456,N_74,N_2731);
nor U6457 (N_6457,N_4929,N_2224);
nand U6458 (N_6458,N_1321,N_1183);
and U6459 (N_6459,N_1214,N_2053);
nand U6460 (N_6460,N_2040,N_1689);
xor U6461 (N_6461,N_4809,N_4907);
nor U6462 (N_6462,N_4297,N_2904);
or U6463 (N_6463,N_2435,N_3359);
or U6464 (N_6464,N_3560,N_3792);
nand U6465 (N_6465,N_2109,N_4685);
and U6466 (N_6466,N_1789,N_4623);
nand U6467 (N_6467,N_2322,N_1368);
nor U6468 (N_6468,N_2691,N_2098);
nor U6469 (N_6469,N_2920,N_4334);
nor U6470 (N_6470,N_3371,N_3559);
xor U6471 (N_6471,N_2141,N_4583);
nor U6472 (N_6472,N_1741,N_664);
and U6473 (N_6473,N_744,N_235);
nor U6474 (N_6474,N_1855,N_1532);
nor U6475 (N_6475,N_4309,N_4596);
nand U6476 (N_6476,N_381,N_3596);
and U6477 (N_6477,N_3637,N_2531);
nor U6478 (N_6478,N_3579,N_1537);
and U6479 (N_6479,N_2773,N_1192);
nand U6480 (N_6480,N_1443,N_2470);
nor U6481 (N_6481,N_1719,N_1932);
nand U6482 (N_6482,N_1173,N_4261);
or U6483 (N_6483,N_2510,N_3927);
xor U6484 (N_6484,N_1243,N_3979);
nor U6485 (N_6485,N_1254,N_4495);
or U6486 (N_6486,N_1517,N_3797);
and U6487 (N_6487,N_757,N_3259);
nor U6488 (N_6488,N_1151,N_4070);
nand U6489 (N_6489,N_3256,N_3782);
nor U6490 (N_6490,N_373,N_4442);
nand U6491 (N_6491,N_3970,N_193);
xor U6492 (N_6492,N_4150,N_507);
nand U6493 (N_6493,N_543,N_4387);
or U6494 (N_6494,N_1417,N_4935);
and U6495 (N_6495,N_1516,N_2884);
nor U6496 (N_6496,N_2990,N_2000);
and U6497 (N_6497,N_502,N_3470);
and U6498 (N_6498,N_2858,N_1278);
xnor U6499 (N_6499,N_2154,N_2788);
xnor U6500 (N_6500,N_428,N_218);
nand U6501 (N_6501,N_4925,N_408);
nand U6502 (N_6502,N_3297,N_1435);
or U6503 (N_6503,N_4863,N_3453);
nand U6504 (N_6504,N_2185,N_555);
or U6505 (N_6505,N_576,N_4011);
nand U6506 (N_6506,N_1706,N_835);
nor U6507 (N_6507,N_691,N_4332);
and U6508 (N_6508,N_3675,N_2574);
or U6509 (N_6509,N_1411,N_2413);
nand U6510 (N_6510,N_249,N_3346);
nor U6511 (N_6511,N_4992,N_358);
nor U6512 (N_6512,N_384,N_4912);
or U6513 (N_6513,N_3327,N_3285);
and U6514 (N_6514,N_4205,N_3043);
nand U6515 (N_6515,N_69,N_250);
xnor U6516 (N_6516,N_2142,N_4682);
or U6517 (N_6517,N_4555,N_2226);
and U6518 (N_6518,N_3955,N_2111);
and U6519 (N_6519,N_2127,N_92);
and U6520 (N_6520,N_4257,N_4648);
nand U6521 (N_6521,N_4207,N_4012);
and U6522 (N_6522,N_3694,N_1133);
nor U6523 (N_6523,N_2952,N_3727);
nor U6524 (N_6524,N_3268,N_1684);
nand U6525 (N_6525,N_2267,N_38);
nor U6526 (N_6526,N_4108,N_2027);
nor U6527 (N_6527,N_2635,N_3562);
nor U6528 (N_6528,N_4864,N_697);
and U6529 (N_6529,N_2780,N_1149);
xor U6530 (N_6530,N_1926,N_2717);
nor U6531 (N_6531,N_550,N_3866);
and U6532 (N_6532,N_2760,N_2579);
xor U6533 (N_6533,N_4657,N_4545);
and U6534 (N_6534,N_2397,N_3652);
nand U6535 (N_6535,N_4715,N_2860);
xnor U6536 (N_6536,N_1088,N_3291);
and U6537 (N_6537,N_156,N_1478);
or U6538 (N_6538,N_2045,N_2854);
or U6539 (N_6539,N_3684,N_3518);
and U6540 (N_6540,N_652,N_4920);
nor U6541 (N_6541,N_4650,N_2707);
or U6542 (N_6542,N_3685,N_3491);
nand U6543 (N_6543,N_2314,N_4464);
nand U6544 (N_6544,N_2419,N_3112);
nor U6545 (N_6545,N_1068,N_1713);
or U6546 (N_6546,N_4182,N_4453);
nor U6547 (N_6547,N_2178,N_2872);
and U6548 (N_6548,N_1272,N_32);
nand U6549 (N_6549,N_4639,N_3188);
or U6550 (N_6550,N_3771,N_1367);
or U6551 (N_6551,N_1331,N_4318);
and U6552 (N_6552,N_568,N_1805);
or U6553 (N_6553,N_85,N_1122);
nor U6554 (N_6554,N_1906,N_1693);
xnor U6555 (N_6555,N_3218,N_1836);
nor U6556 (N_6556,N_3088,N_4046);
nand U6557 (N_6557,N_1040,N_1034);
or U6558 (N_6558,N_2695,N_4301);
or U6559 (N_6559,N_1318,N_4157);
and U6560 (N_6560,N_1883,N_3964);
or U6561 (N_6561,N_2384,N_4896);
or U6562 (N_6562,N_3149,N_372);
nor U6563 (N_6563,N_3884,N_1676);
or U6564 (N_6564,N_3139,N_2065);
nand U6565 (N_6565,N_2871,N_1163);
nor U6566 (N_6566,N_2380,N_740);
xor U6567 (N_6567,N_2001,N_496);
and U6568 (N_6568,N_2982,N_646);
xor U6569 (N_6569,N_240,N_4812);
nor U6570 (N_6570,N_4162,N_316);
nand U6571 (N_6571,N_3655,N_4177);
nand U6572 (N_6572,N_2496,N_2732);
and U6573 (N_6573,N_13,N_1635);
and U6574 (N_6574,N_3128,N_2474);
nor U6575 (N_6575,N_3084,N_2082);
and U6576 (N_6576,N_46,N_681);
and U6577 (N_6577,N_4556,N_2764);
and U6578 (N_6578,N_675,N_847);
nand U6579 (N_6579,N_2640,N_1678);
and U6580 (N_6580,N_2054,N_2491);
nand U6581 (N_6581,N_903,N_2131);
xor U6582 (N_6582,N_3053,N_12);
nand U6583 (N_6583,N_959,N_1337);
nor U6584 (N_6584,N_2325,N_1345);
nand U6585 (N_6585,N_3284,N_2606);
nor U6586 (N_6586,N_4428,N_4814);
or U6587 (N_6587,N_1839,N_4074);
and U6588 (N_6588,N_4861,N_4725);
xnor U6589 (N_6589,N_4688,N_2355);
nand U6590 (N_6590,N_4323,N_4482);
nor U6591 (N_6591,N_3032,N_3932);
or U6592 (N_6592,N_443,N_1400);
nor U6593 (N_6593,N_4199,N_3936);
nor U6594 (N_6594,N_3814,N_4593);
or U6595 (N_6595,N_1258,N_2734);
and U6596 (N_6596,N_4719,N_3081);
nor U6597 (N_6597,N_4412,N_2608);
and U6598 (N_6598,N_614,N_1338);
nand U6599 (N_6599,N_1527,N_256);
nor U6600 (N_6600,N_2042,N_4729);
nand U6601 (N_6601,N_2950,N_3428);
and U6602 (N_6602,N_2971,N_3671);
or U6603 (N_6603,N_3484,N_3289);
nor U6604 (N_6604,N_216,N_656);
nand U6605 (N_6605,N_253,N_52);
nand U6606 (N_6606,N_912,N_569);
and U6607 (N_6607,N_4652,N_2012);
and U6608 (N_6608,N_3865,N_2306);
or U6609 (N_6609,N_1074,N_102);
or U6610 (N_6610,N_1268,N_4238);
nand U6611 (N_6611,N_441,N_1519);
nand U6612 (N_6612,N_1207,N_280);
or U6613 (N_6613,N_780,N_3119);
nor U6614 (N_6614,N_4834,N_3874);
nor U6615 (N_6615,N_1255,N_1026);
nor U6616 (N_6616,N_3105,N_3006);
nor U6617 (N_6617,N_1561,N_1202);
or U6618 (N_6618,N_4418,N_3586);
xor U6619 (N_6619,N_435,N_4924);
nor U6620 (N_6620,N_247,N_4276);
xor U6621 (N_6621,N_2844,N_4893);
or U6622 (N_6622,N_4709,N_229);
and U6623 (N_6623,N_3870,N_4687);
nand U6624 (N_6624,N_4143,N_1569);
and U6625 (N_6625,N_3406,N_2763);
and U6626 (N_6626,N_498,N_1199);
nor U6627 (N_6627,N_2614,N_1065);
nor U6628 (N_6628,N_1362,N_112);
nor U6629 (N_6629,N_2517,N_3206);
nor U6630 (N_6630,N_3989,N_2786);
or U6631 (N_6631,N_3572,N_3111);
nand U6632 (N_6632,N_2694,N_3515);
and U6633 (N_6633,N_816,N_4850);
nor U6634 (N_6634,N_3381,N_2337);
nor U6635 (N_6635,N_274,N_4787);
nor U6636 (N_6636,N_1334,N_3954);
or U6637 (N_6637,N_412,N_2989);
nor U6638 (N_6638,N_402,N_4870);
nor U6639 (N_6639,N_3216,N_2577);
and U6640 (N_6640,N_3023,N_2509);
xor U6641 (N_6641,N_1138,N_4256);
or U6642 (N_6642,N_322,N_1993);
nand U6643 (N_6643,N_3456,N_1731);
nor U6644 (N_6644,N_2081,N_3913);
or U6645 (N_6645,N_1456,N_3905);
nor U6646 (N_6646,N_2983,N_2836);
xor U6647 (N_6647,N_3199,N_4990);
xnor U6648 (N_6648,N_4034,N_95);
xnor U6649 (N_6649,N_1342,N_4951);
and U6650 (N_6650,N_2686,N_1545);
or U6651 (N_6651,N_551,N_3631);
and U6652 (N_6652,N_514,N_2338);
xor U6653 (N_6653,N_456,N_3670);
nand U6654 (N_6654,N_1335,N_935);
nor U6655 (N_6655,N_4271,N_4778);
nand U6656 (N_6656,N_3108,N_90);
nor U6657 (N_6657,N_3784,N_4028);
and U6658 (N_6658,N_3856,N_911);
xor U6659 (N_6659,N_607,N_4686);
nand U6660 (N_6660,N_3835,N_3342);
nor U6661 (N_6661,N_679,N_1361);
nand U6662 (N_6662,N_1166,N_2778);
or U6663 (N_6663,N_4828,N_1940);
nand U6664 (N_6664,N_1809,N_1431);
and U6665 (N_6665,N_4193,N_723);
nand U6666 (N_6666,N_3673,N_4885);
and U6667 (N_6667,N_2408,N_2222);
nor U6668 (N_6668,N_3891,N_4766);
and U6669 (N_6669,N_1330,N_4552);
and U6670 (N_6670,N_640,N_1274);
nand U6671 (N_6671,N_454,N_169);
nor U6672 (N_6672,N_1723,N_2143);
nor U6673 (N_6673,N_3994,N_3328);
xor U6674 (N_6674,N_3280,N_3299);
and U6675 (N_6675,N_1284,N_2138);
and U6676 (N_6676,N_2644,N_132);
nand U6677 (N_6677,N_1383,N_214);
nor U6678 (N_6678,N_4327,N_725);
nor U6679 (N_6679,N_2865,N_4939);
or U6680 (N_6680,N_4080,N_147);
or U6681 (N_6681,N_2611,N_3660);
or U6682 (N_6682,N_2334,N_866);
and U6683 (N_6683,N_4830,N_273);
and U6684 (N_6684,N_2900,N_175);
xnor U6685 (N_6685,N_542,N_2687);
nand U6686 (N_6686,N_1709,N_3054);
xnor U6687 (N_6687,N_4740,N_4383);
nand U6688 (N_6688,N_2028,N_4152);
nor U6689 (N_6689,N_3599,N_3845);
and U6690 (N_6690,N_1530,N_3398);
and U6691 (N_6691,N_2323,N_958);
or U6692 (N_6692,N_924,N_2271);
and U6693 (N_6693,N_2663,N_2934);
and U6694 (N_6694,N_574,N_3530);
and U6695 (N_6695,N_149,N_4765);
and U6696 (N_6696,N_694,N_1164);
and U6697 (N_6697,N_241,N_2703);
or U6698 (N_6698,N_1868,N_3805);
nor U6699 (N_6699,N_4974,N_819);
or U6700 (N_6700,N_4393,N_4288);
nand U6701 (N_6701,N_4559,N_4735);
and U6702 (N_6702,N_929,N_1554);
nor U6703 (N_6703,N_3734,N_4969);
and U6704 (N_6704,N_918,N_3823);
or U6705 (N_6705,N_3157,N_3570);
or U6706 (N_6706,N_2584,N_936);
or U6707 (N_6707,N_711,N_2424);
and U6708 (N_6708,N_2701,N_1210);
nor U6709 (N_6709,N_3215,N_3421);
nand U6710 (N_6710,N_2416,N_751);
and U6711 (N_6711,N_1633,N_2187);
nand U6712 (N_6712,N_1482,N_4576);
and U6713 (N_6713,N_1466,N_2824);
and U6714 (N_6714,N_4791,N_434);
and U6715 (N_6715,N_2782,N_1057);
and U6716 (N_6716,N_3275,N_4748);
nor U6717 (N_6717,N_3766,N_534);
or U6718 (N_6718,N_2598,N_1792);
or U6719 (N_6719,N_2316,N_1583);
or U6720 (N_6720,N_1432,N_3647);
xor U6721 (N_6721,N_678,N_307);
nand U6722 (N_6722,N_2255,N_1441);
nor U6723 (N_6723,N_3252,N_896);
or U6724 (N_6724,N_2202,N_2103);
and U6725 (N_6725,N_4643,N_4192);
or U6726 (N_6726,N_319,N_601);
or U6727 (N_6727,N_2781,N_2702);
nor U6728 (N_6728,N_1915,N_1810);
nand U6729 (N_6729,N_1323,N_1880);
nor U6730 (N_6730,N_1010,N_2864);
xnor U6731 (N_6731,N_390,N_3137);
and U6732 (N_6732,N_4246,N_4090);
or U6733 (N_6733,N_2682,N_346);
nand U6734 (N_6734,N_495,N_993);
nand U6735 (N_6735,N_1536,N_875);
or U6736 (N_6736,N_4644,N_2985);
xor U6737 (N_6737,N_430,N_1110);
xnor U6738 (N_6738,N_4961,N_4895);
xnor U6739 (N_6739,N_1804,N_722);
nand U6740 (N_6740,N_1477,N_940);
nor U6741 (N_6741,N_4338,N_3827);
or U6742 (N_6742,N_2560,N_3603);
nand U6743 (N_6743,N_4095,N_3721);
nand U6744 (N_6744,N_2257,N_1842);
nand U6745 (N_6745,N_254,N_3089);
nand U6746 (N_6746,N_1673,N_4535);
nor U6747 (N_6747,N_2918,N_2791);
and U6748 (N_6748,N_3613,N_972);
nor U6749 (N_6749,N_1987,N_232);
and U6750 (N_6750,N_1100,N_4188);
nor U6751 (N_6751,N_416,N_3502);
nand U6752 (N_6752,N_4696,N_1637);
or U6753 (N_6753,N_2873,N_1778);
or U6754 (N_6754,N_2777,N_4317);
or U6755 (N_6755,N_4953,N_742);
nand U6756 (N_6756,N_674,N_31);
and U6757 (N_6757,N_3890,N_3385);
and U6758 (N_6758,N_194,N_966);
and U6759 (N_6759,N_1797,N_4983);
nand U6760 (N_6760,N_3071,N_2201);
nor U6761 (N_6761,N_4601,N_2076);
nor U6762 (N_6762,N_916,N_895);
or U6763 (N_6763,N_2170,N_3623);
and U6764 (N_6764,N_1793,N_2225);
or U6765 (N_6765,N_3746,N_2328);
or U6766 (N_6766,N_1402,N_4413);
xnor U6767 (N_6767,N_544,N_4463);
nand U6768 (N_6768,N_4804,N_3509);
nor U6769 (N_6769,N_493,N_738);
or U6770 (N_6770,N_2231,N_1577);
nor U6771 (N_6771,N_2400,N_152);
and U6772 (N_6772,N_4078,N_1726);
nor U6773 (N_6773,N_1808,N_492);
or U6774 (N_6774,N_440,N_2647);
nand U6775 (N_6775,N_1969,N_3881);
and U6776 (N_6776,N_1396,N_1238);
nor U6777 (N_6777,N_3333,N_657);
and U6778 (N_6778,N_1667,N_4775);
or U6779 (N_6779,N_806,N_1579);
and U6780 (N_6780,N_491,N_2740);
nor U6781 (N_6781,N_3859,N_4456);
xnor U6782 (N_6782,N_1071,N_736);
nand U6783 (N_6783,N_1327,N_2783);
and U6784 (N_6784,N_2804,N_1339);
xnor U6785 (N_6785,N_4550,N_2481);
nand U6786 (N_6786,N_1009,N_642);
or U6787 (N_6787,N_2299,N_1912);
or U6788 (N_6788,N_2848,N_2206);
xor U6789 (N_6789,N_3581,N_4954);
nand U6790 (N_6790,N_2121,N_3332);
nor U6791 (N_6791,N_1048,N_2026);
nand U6792 (N_6792,N_939,N_1817);
nor U6793 (N_6793,N_3717,N_3384);
nand U6794 (N_6794,N_3263,N_4918);
and U6795 (N_6795,N_1974,N_1985);
or U6796 (N_6796,N_4241,N_3661);
nand U6797 (N_6797,N_183,N_2208);
and U6798 (N_6798,N_2876,N_2558);
nand U6799 (N_6799,N_2217,N_608);
or U6800 (N_6800,N_3288,N_3564);
and U6801 (N_6801,N_3598,N_3214);
or U6802 (N_6802,N_4915,N_3220);
or U6803 (N_6803,N_2683,N_4435);
and U6804 (N_6804,N_3828,N_4841);
nand U6805 (N_6805,N_3313,N_4469);
nor U6806 (N_6806,N_3273,N_1645);
and U6807 (N_6807,N_3593,N_93);
nor U6808 (N_6808,N_2916,N_1407);
or U6809 (N_6809,N_3857,N_4365);
nor U6810 (N_6810,N_2157,N_4223);
and U6811 (N_6811,N_2227,N_4616);
and U6812 (N_6812,N_3842,N_4605);
xnor U6813 (N_6813,N_4496,N_4860);
nand U6814 (N_6814,N_4668,N_3007);
nor U6815 (N_6815,N_2907,N_130);
nor U6816 (N_6816,N_4763,N_4203);
nand U6817 (N_6817,N_4632,N_114);
or U6818 (N_6818,N_2365,N_2933);
xnor U6819 (N_6819,N_4871,N_40);
nand U6820 (N_6820,N_3100,N_2189);
or U6821 (N_6821,N_3493,N_4471);
and U6822 (N_6822,N_4336,N_227);
nor U6823 (N_6823,N_3818,N_3147);
nor U6824 (N_6824,N_1788,N_2444);
and U6825 (N_6825,N_4117,N_4502);
xor U6826 (N_6826,N_3877,N_1897);
or U6827 (N_6827,N_3281,N_4439);
and U6828 (N_6828,N_1925,N_1963);
nand U6829 (N_6829,N_2373,N_4454);
nor U6830 (N_6830,N_3236,N_166);
nand U6831 (N_6831,N_8,N_2564);
nand U6832 (N_6832,N_696,N_4348);
and U6833 (N_6833,N_3949,N_3169);
and U6834 (N_6834,N_4092,N_623);
xnor U6835 (N_6835,N_3073,N_3411);
and U6836 (N_6836,N_805,N_2133);
and U6837 (N_6837,N_1388,N_2119);
or U6838 (N_6838,N_1798,N_1329);
and U6839 (N_6839,N_2519,N_4216);
xnor U6840 (N_6840,N_1886,N_2850);
nand U6841 (N_6841,N_2580,N_1085);
nor U6842 (N_6842,N_1099,N_1394);
or U6843 (N_6843,N_293,N_1508);
or U6844 (N_6844,N_2947,N_1393);
nor U6845 (N_6845,N_4172,N_1596);
xor U6846 (N_6846,N_3794,N_2705);
nand U6847 (N_6847,N_431,N_513);
and U6848 (N_6848,N_3027,N_4798);
or U6849 (N_6849,N_4121,N_4359);
and U6850 (N_6850,N_2101,N_2483);
or U6851 (N_6851,N_4388,N_506);
or U6852 (N_6852,N_4470,N_830);
nand U6853 (N_6853,N_4321,N_701);
nand U6854 (N_6854,N_4218,N_2720);
or U6855 (N_6855,N_1889,N_1748);
and U6856 (N_6856,N_3462,N_1490);
xor U6857 (N_6857,N_784,N_2746);
nor U6858 (N_6858,N_1783,N_4656);
or U6859 (N_6859,N_1060,N_275);
nand U6860 (N_6860,N_3377,N_4921);
and U6861 (N_6861,N_3720,N_2353);
or U6862 (N_6862,N_3184,N_2697);
nor U6863 (N_6863,N_2805,N_3204);
and U6864 (N_6864,N_2932,N_5);
nor U6865 (N_6865,N_1054,N_4351);
nand U6866 (N_6866,N_2758,N_379);
or U6867 (N_6867,N_3150,N_3864);
or U6868 (N_6868,N_2067,N_3003);
nand U6869 (N_6869,N_1171,N_3083);
nor U6870 (N_6870,N_598,N_1442);
nor U6871 (N_6871,N_3553,N_2648);
nor U6872 (N_6872,N_3272,N_3048);
or U6873 (N_6873,N_108,N_2426);
and U6874 (N_6874,N_1902,N_1947);
nand U6875 (N_6875,N_1273,N_4370);
nand U6876 (N_6876,N_3387,N_26);
nor U6877 (N_6877,N_3171,N_2980);
or U6878 (N_6878,N_1378,N_2586);
xnor U6879 (N_6879,N_2210,N_1816);
xnor U6880 (N_6880,N_1190,N_394);
nor U6881 (N_6881,N_42,N_2391);
and U6882 (N_6882,N_3745,N_2721);
or U6883 (N_6883,N_2908,N_3368);
nor U6884 (N_6884,N_1125,N_926);
and U6885 (N_6885,N_1715,N_3314);
nor U6886 (N_6886,N_304,N_3369);
and U6887 (N_6887,N_4595,N_1898);
or U6888 (N_6888,N_1740,N_3565);
nor U6889 (N_6889,N_2117,N_1598);
or U6890 (N_6890,N_1720,N_4520);
or U6891 (N_6891,N_3191,N_3736);
nor U6892 (N_6892,N_2313,N_3917);
xnor U6893 (N_6893,N_1115,N_4611);
or U6894 (N_6894,N_1500,N_4699);
xnor U6895 (N_6895,N_4283,N_3019);
nand U6896 (N_6896,N_2569,N_4771);
xnor U6897 (N_6897,N_2901,N_1736);
nor U6898 (N_6898,N_1275,N_4481);
or U6899 (N_6899,N_3087,N_1341);
and U6900 (N_6900,N_2064,N_2535);
nor U6901 (N_6901,N_252,N_3566);
and U6902 (N_6902,N_60,N_1955);
xor U6903 (N_6903,N_3235,N_3480);
and U6904 (N_6904,N_2052,N_3465);
or U6905 (N_6905,N_1644,N_2828);
and U6906 (N_6906,N_3906,N_3674);
nor U6907 (N_6907,N_2122,N_4055);
nor U6908 (N_6908,N_4967,N_1704);
nor U6909 (N_6909,N_4360,N_4710);
nor U6910 (N_6910,N_3464,N_3459);
nor U6911 (N_6911,N_1130,N_1843);
nor U6912 (N_6912,N_4618,N_210);
nor U6913 (N_6913,N_3304,N_1971);
nor U6914 (N_6914,N_4548,N_3900);
and U6915 (N_6915,N_917,N_2796);
and U6916 (N_6916,N_4075,N_1764);
nor U6917 (N_6917,N_1702,N_3679);
nand U6918 (N_6918,N_3554,N_2881);
or U6919 (N_6919,N_2684,N_1680);
and U6920 (N_6920,N_716,N_2074);
and U6921 (N_6921,N_292,N_135);
or U6922 (N_6922,N_2180,N_2021);
and U6923 (N_6923,N_1073,N_4603);
and U6924 (N_6924,N_3294,N_4736);
nand U6925 (N_6925,N_2588,N_4233);
and U6926 (N_6926,N_1422,N_2434);
nor U6927 (N_6927,N_2093,N_3757);
and U6928 (N_6928,N_312,N_4888);
nand U6929 (N_6929,N_283,N_1975);
and U6930 (N_6930,N_636,N_3340);
nor U6931 (N_6931,N_1381,N_651);
or U6932 (N_6932,N_1497,N_4789);
nor U6933 (N_6933,N_2371,N_4068);
nor U6934 (N_6934,N_4016,N_3773);
nand U6935 (N_6935,N_4982,N_445);
nand U6936 (N_6936,N_3735,N_1601);
nor U6937 (N_6937,N_432,N_1351);
and U6938 (N_6938,N_296,N_1080);
or U6939 (N_6939,N_1322,N_4508);
xor U6940 (N_6940,N_2709,N_961);
xor U6941 (N_6941,N_4133,N_517);
nand U6942 (N_6942,N_391,N_589);
or U6943 (N_6943,N_3975,N_945);
or U6944 (N_6944,N_2775,N_4302);
and U6945 (N_6945,N_225,N_2401);
and U6946 (N_6946,N_721,N_4816);
or U6947 (N_6947,N_1076,N_28);
or U6948 (N_6948,N_3742,N_637);
and U6949 (N_6949,N_1606,N_3976);
and U6950 (N_6950,N_3761,N_2261);
or U6951 (N_6951,N_331,N_4149);
and U6952 (N_6952,N_4607,N_1594);
nor U6953 (N_6953,N_1849,N_2073);
nor U6954 (N_6954,N_1661,N_2548);
or U6955 (N_6955,N_500,N_753);
or U6956 (N_6956,N_1446,N_3733);
and U6957 (N_6957,N_3953,N_1089);
xor U6958 (N_6958,N_3366,N_2634);
and U6959 (N_6959,N_644,N_4050);
xnor U6960 (N_6960,N_3390,N_3407);
nand U6961 (N_6961,N_222,N_184);
or U6962 (N_6962,N_2171,N_2666);
nand U6963 (N_6963,N_4641,N_2072);
nor U6964 (N_6964,N_4329,N_2439);
or U6965 (N_6965,N_3648,N_1389);
or U6966 (N_6966,N_2308,N_893);
nor U6967 (N_6967,N_1454,N_2575);
xor U6968 (N_6968,N_2349,N_1495);
or U6969 (N_6969,N_4563,N_4711);
nand U6970 (N_6970,N_2097,N_2696);
nand U6971 (N_6971,N_923,N_2829);
nor U6972 (N_6972,N_2852,N_1986);
and U6973 (N_6973,N_3254,N_4285);
nand U6974 (N_6974,N_1310,N_1831);
nor U6975 (N_6975,N_2855,N_2689);
or U6976 (N_6976,N_3409,N_1285);
or U6977 (N_6977,N_2294,N_732);
or U6978 (N_6978,N_1027,N_1158);
nor U6979 (N_6979,N_3277,N_2285);
or U6980 (N_6980,N_2004,N_1249);
and U6981 (N_6981,N_4421,N_1447);
nand U6982 (N_6982,N_2238,N_3501);
nor U6983 (N_6983,N_270,N_1584);
xor U6984 (N_6984,N_2877,N_2906);
nand U6985 (N_6985,N_3146,N_122);
or U6986 (N_6986,N_44,N_2449);
nand U6987 (N_6987,N_3960,N_823);
or U6988 (N_6988,N_1950,N_946);
nor U6989 (N_6989,N_1153,N_2252);
or U6990 (N_6990,N_419,N_4782);
nor U6991 (N_6991,N_4128,N_2818);
or U6992 (N_6992,N_2677,N_1686);
nand U6993 (N_6993,N_813,N_3363);
nand U6994 (N_6994,N_266,N_3561);
nand U6995 (N_6995,N_680,N_1070);
nand U6996 (N_6996,N_3257,N_1379);
or U6997 (N_6997,N_1444,N_3011);
or U6998 (N_6998,N_2772,N_3516);
or U6999 (N_6999,N_4825,N_4215);
xnor U7000 (N_7000,N_1003,N_2593);
nor U7001 (N_7001,N_4679,N_289);
nand U7002 (N_7002,N_3556,N_4230);
nand U7003 (N_7003,N_4039,N_1291);
or U7004 (N_7004,N_2515,N_4032);
and U7005 (N_7005,N_1881,N_4937);
nand U7006 (N_7006,N_3499,N_3662);
nor U7007 (N_7007,N_4364,N_1802);
nor U7008 (N_7008,N_1953,N_2662);
or U7009 (N_7009,N_2942,N_4480);
nand U7010 (N_7010,N_219,N_1761);
xor U7011 (N_7011,N_2258,N_639);
nor U7012 (N_7012,N_1475,N_4444);
or U7013 (N_7013,N_3234,N_2396);
xnor U7014 (N_7014,N_35,N_2128);
and U7015 (N_7015,N_624,N_2363);
or U7016 (N_7016,N_3269,N_2379);
nor U7017 (N_7017,N_380,N_2660);
xnor U7018 (N_7018,N_2869,N_3968);
and U7019 (N_7019,N_599,N_1145);
or U7020 (N_7020,N_2939,N_221);
nor U7021 (N_7021,N_990,N_4036);
nor U7022 (N_7022,N_2130,N_3557);
nor U7023 (N_7023,N_1692,N_2104);
or U7024 (N_7024,N_1927,N_4138);
nor U7025 (N_7025,N_115,N_3424);
and U7026 (N_7026,N_196,N_387);
or U7027 (N_7027,N_139,N_1872);
xnor U7028 (N_7028,N_2209,N_2276);
xnor U7029 (N_7029,N_1956,N_1670);
and U7030 (N_7030,N_314,N_99);
nand U7031 (N_7031,N_2193,N_55);
or U7032 (N_7032,N_4532,N_2902);
nor U7033 (N_7033,N_3503,N_105);
nor U7034 (N_7034,N_2959,N_2573);
nand U7035 (N_7035,N_3531,N_2114);
nand U7036 (N_7036,N_142,N_2879);
xnor U7037 (N_7037,N_4987,N_2144);
or U7038 (N_7038,N_920,N_1714);
nand U7039 (N_7039,N_3754,N_2039);
or U7040 (N_7040,N_1911,N_3389);
nor U7041 (N_7041,N_3517,N_992);
nand U7042 (N_7042,N_3055,N_1180);
nand U7043 (N_7043,N_2372,N_3436);
or U7044 (N_7044,N_1562,N_489);
and U7045 (N_7045,N_2958,N_3795);
and U7046 (N_7046,N_1669,N_1370);
xnor U7047 (N_7047,N_176,N_125);
nor U7048 (N_7048,N_236,N_4197);
and U7049 (N_7049,N_4310,N_2068);
xnor U7050 (N_7050,N_3992,N_600);
and U7051 (N_7051,N_1636,N_3098);
nor U7052 (N_7052,N_3482,N_890);
or U7053 (N_7053,N_3237,N_2106);
nor U7054 (N_7054,N_436,N_106);
nand U7055 (N_7055,N_776,N_2179);
or U7056 (N_7056,N_3982,N_3568);
and U7057 (N_7057,N_2159,N_2063);
and U7058 (N_7058,N_4741,N_2768);
or U7059 (N_7059,N_1228,N_1512);
or U7060 (N_7060,N_3524,N_2642);
and U7061 (N_7061,N_4770,N_3395);
nor U7062 (N_7062,N_4250,N_4475);
nor U7063 (N_7063,N_75,N_4801);
and U7064 (N_7064,N_2704,N_239);
nor U7065 (N_7065,N_2041,N_3700);
nor U7066 (N_7066,N_4259,N_4849);
nand U7067 (N_7067,N_1053,N_2460);
or U7068 (N_7068,N_2806,N_2194);
nand U7069 (N_7069,N_3101,N_1052);
or U7070 (N_7070,N_4659,N_4147);
or U7071 (N_7071,N_1460,N_4819);
and U7072 (N_7072,N_4381,N_1051);
or U7073 (N_7073,N_1851,N_4371);
and U7074 (N_7074,N_4554,N_872);
nor U7075 (N_7075,N_311,N_3244);
or U7076 (N_7076,N_245,N_4516);
nor U7077 (N_7077,N_4615,N_2259);
or U7078 (N_7078,N_4375,N_4837);
and U7079 (N_7079,N_3152,N_2330);
nor U7080 (N_7080,N_1538,N_2237);
or U7081 (N_7081,N_1867,N_4989);
nand U7082 (N_7082,N_2539,N_317);
nand U7083 (N_7083,N_3958,N_410);
or U7084 (N_7084,N_3922,N_1729);
nor U7085 (N_7085,N_1549,N_2833);
nand U7086 (N_7086,N_1572,N_4141);
nor U7087 (N_7087,N_2216,N_3350);
nand U7088 (N_7088,N_1525,N_4581);
nor U7089 (N_7089,N_1168,N_2266);
nor U7090 (N_7090,N_477,N_3141);
or U7091 (N_7091,N_20,N_143);
and U7092 (N_7092,N_1772,N_2502);
and U7093 (N_7093,N_3615,N_3038);
xor U7094 (N_7094,N_1055,N_1954);
or U7095 (N_7095,N_345,N_2585);
or U7096 (N_7096,N_4515,N_944);
nand U7097 (N_7097,N_3122,N_3192);
and U7098 (N_7098,N_199,N_1061);
nor U7099 (N_7099,N_2443,N_4005);
nor U7100 (N_7100,N_191,N_3589);
nor U7101 (N_7101,N_700,N_1177);
nand U7102 (N_7102,N_1919,N_1128);
and U7103 (N_7103,N_2091,N_4590);
or U7104 (N_7104,N_4667,N_4377);
and U7105 (N_7105,N_4316,N_1062);
nand U7106 (N_7106,N_3301,N_3072);
nor U7107 (N_7107,N_815,N_862);
and U7108 (N_7108,N_1547,N_3844);
nand U7109 (N_7109,N_267,N_4056);
or U7110 (N_7110,N_4040,N_2375);
and U7111 (N_7111,N_3985,N_1286);
nor U7112 (N_7112,N_3017,N_4549);
or U7113 (N_7113,N_4751,N_602);
nand U7114 (N_7114,N_2200,N_2376);
nor U7115 (N_7115,N_4148,N_3243);
nor U7116 (N_7116,N_2051,N_523);
or U7117 (N_7117,N_3126,N_1029);
nor U7118 (N_7118,N_4553,N_3608);
nand U7119 (N_7119,N_3153,N_2279);
and U7120 (N_7120,N_2715,N_4934);
nand U7121 (N_7121,N_3991,N_2377);
nand U7122 (N_7122,N_4536,N_2887);
nand U7123 (N_7123,N_1316,N_2880);
nand U7124 (N_7124,N_1758,N_3116);
nand U7125 (N_7125,N_3651,N_3896);
xor U7126 (N_7126,N_2787,N_2264);
or U7127 (N_7127,N_4255,N_4115);
or U7128 (N_7128,N_1226,N_3046);
nor U7129 (N_7129,N_2866,N_4509);
nand U7130 (N_7130,N_3838,N_582);
and U7131 (N_7131,N_3431,N_1395);
nand U7132 (N_7132,N_3946,N_1297);
nand U7133 (N_7133,N_586,N_2856);
or U7134 (N_7134,N_4564,N_2561);
or U7135 (N_7135,N_4084,N_4627);
nor U7136 (N_7136,N_4680,N_2069);
nor U7137 (N_7137,N_2511,N_4102);
nand U7138 (N_7138,N_977,N_3374);
and U7139 (N_7139,N_458,N_4949);
nor U7140 (N_7140,N_2861,N_1511);
nor U7141 (N_7141,N_865,N_3077);
and U7142 (N_7142,N_4847,N_260);
xnor U7143 (N_7143,N_1722,N_2743);
nor U7144 (N_7144,N_4167,N_3948);
nor U7145 (N_7145,N_887,N_4242);
and U7146 (N_7146,N_3892,N_4419);
nor U7147 (N_7147,N_4490,N_3883);
and U7148 (N_7148,N_769,N_4487);
and U7149 (N_7149,N_4872,N_1542);
or U7150 (N_7150,N_4258,N_4503);
and U7151 (N_7151,N_3879,N_1413);
and U7152 (N_7152,N_3078,N_349);
xor U7153 (N_7153,N_2700,N_900);
nand U7154 (N_7154,N_856,N_4663);
and U7155 (N_7155,N_48,N_2812);
or U7156 (N_7156,N_3939,N_3420);
or U7157 (N_7157,N_3867,N_1111);
or U7158 (N_7158,N_2034,N_359);
nand U7159 (N_7159,N_4232,N_1840);
or U7160 (N_7160,N_794,N_983);
nor U7161 (N_7161,N_1664,N_3625);
nor U7162 (N_7162,N_970,N_4063);
and U7163 (N_7163,N_2749,N_4674);
nand U7164 (N_7164,N_1982,N_870);
and U7165 (N_7165,N_1364,N_3514);
or U7166 (N_7166,N_4164,N_3477);
nor U7167 (N_7167,N_2002,N_4073);
and U7168 (N_7168,N_1347,N_4155);
or U7169 (N_7169,N_4340,N_4749);
or U7170 (N_7170,N_2823,N_883);
or U7171 (N_7171,N_2282,N_1944);
or U7172 (N_7172,N_124,N_3850);
nor U7173 (N_7173,N_4671,N_3266);
and U7174 (N_7174,N_1991,N_3676);
and U7175 (N_7175,N_2699,N_1205);
nand U7176 (N_7176,N_2641,N_1768);
nor U7177 (N_7177,N_548,N_1814);
and U7178 (N_7178,N_2668,N_1904);
nor U7179 (N_7179,N_1269,N_2831);
xnor U7180 (N_7180,N_2274,N_1229);
nand U7181 (N_7181,N_773,N_3682);
xnor U7182 (N_7182,N_2221,N_708);
or U7183 (N_7183,N_1612,N_2669);
and U7184 (N_7184,N_859,N_3176);
nand U7185 (N_7185,N_3303,N_3929);
nand U7186 (N_7186,N_1978,N_2169);
xnor U7187 (N_7187,N_2242,N_2478);
nor U7188 (N_7188,N_4222,N_1509);
nand U7189 (N_7189,N_4997,N_2088);
or U7190 (N_7190,N_2370,N_2941);
or U7191 (N_7191,N_2978,N_4200);
or U7192 (N_7192,N_4229,N_1832);
nand U7193 (N_7193,N_3094,N_3938);
nor U7194 (N_7194,N_159,N_1234);
or U7195 (N_7195,N_320,N_2545);
or U7196 (N_7196,N_1008,N_2290);
or U7197 (N_7197,N_4153,N_3632);
and U7198 (N_7198,N_2853,N_4399);
or U7199 (N_7199,N_3793,N_2676);
nand U7200 (N_7200,N_3025,N_2333);
or U7201 (N_7201,N_2929,N_3271);
nand U7202 (N_7202,N_1603,N_2107);
and U7203 (N_7203,N_4759,N_3429);
or U7204 (N_7204,N_3162,N_1786);
xor U7205 (N_7205,N_2156,N_3056);
and U7206 (N_7206,N_1690,N_4588);
or U7207 (N_7207,N_4975,N_1231);
nor U7208 (N_7208,N_4426,N_4136);
nor U7209 (N_7209,N_4689,N_1289);
xnor U7210 (N_7210,N_313,N_1358);
nor U7211 (N_7211,N_3699,N_752);
or U7212 (N_7212,N_3920,N_1313);
or U7213 (N_7213,N_2006,N_136);
or U7214 (N_7214,N_4458,N_2461);
nor U7215 (N_7215,N_3611,N_4265);
and U7216 (N_7216,N_24,N_3744);
nor U7217 (N_7217,N_1141,N_3102);
nor U7218 (N_7218,N_3466,N_1642);
and U7219 (N_7219,N_1742,N_57);
or U7220 (N_7220,N_185,N_3463);
or U7221 (N_7221,N_4947,N_104);
or U7222 (N_7222,N_4697,N_4940);
nor U7223 (N_7223,N_3080,N_994);
nor U7224 (N_7224,N_2335,N_4097);
and U7225 (N_7225,N_3918,N_429);
xor U7226 (N_7226,N_2524,N_4906);
nor U7227 (N_7227,N_1281,N_4433);
and U7228 (N_7228,N_1929,N_1012);
and U7229 (N_7229,N_4518,N_4718);
or U7230 (N_7230,N_465,N_982);
xor U7231 (N_7231,N_3365,N_927);
and U7232 (N_7232,N_686,N_3261);
nand U7233 (N_7233,N_3394,N_1479);
and U7234 (N_7234,N_2409,N_1217);
nand U7235 (N_7235,N_1884,N_121);
nand U7236 (N_7236,N_1416,N_2223);
and U7237 (N_7237,N_4196,N_4221);
nand U7238 (N_7238,N_4427,N_4646);
and U7239 (N_7239,N_1257,N_3578);
or U7240 (N_7240,N_554,N_4106);
nor U7241 (N_7241,N_4746,N_4282);
nor U7242 (N_7242,N_3815,N_706);
and U7243 (N_7243,N_325,N_4025);
and U7244 (N_7244,N_2174,N_1175);
or U7245 (N_7245,N_2324,N_3539);
or U7246 (N_7246,N_669,N_4202);
or U7247 (N_7247,N_3210,N_423);
nand U7248 (N_7248,N_759,N_1961);
and U7249 (N_7249,N_362,N_2120);
nor U7250 (N_7250,N_2356,N_2319);
and U7251 (N_7251,N_25,N_3622);
and U7252 (N_7252,N_3819,N_2960);
nand U7253 (N_7253,N_2250,N_188);
or U7254 (N_7254,N_2488,N_1790);
nand U7255 (N_7255,N_625,N_2505);
nor U7256 (N_7256,N_181,N_4567);
nand U7257 (N_7257,N_276,N_2987);
nand U7258 (N_7258,N_877,N_439);
or U7259 (N_7259,N_4757,N_265);
xnor U7260 (N_7260,N_2118,N_1654);
nor U7261 (N_7261,N_211,N_3824);
xor U7262 (N_7262,N_3279,N_1222);
or U7263 (N_7263,N_4946,N_4361);
or U7264 (N_7264,N_1239,N_855);
nand U7265 (N_7265,N_2269,N_2843);
or U7266 (N_7266,N_573,N_2361);
and U7267 (N_7267,N_864,N_4382);
or U7268 (N_7268,N_4637,N_4449);
nor U7269 (N_7269,N_4945,N_3654);
or U7270 (N_7270,N_3476,N_1746);
nand U7271 (N_7271,N_2023,N_2785);
and U7272 (N_7272,N_3781,N_4462);
nor U7273 (N_7273,N_2112,N_503);
and U7274 (N_7274,N_4000,N_1807);
or U7275 (N_7275,N_2207,N_1203);
nor U7276 (N_7276,N_3140,N_1751);
nor U7277 (N_7277,N_3580,N_3330);
nand U7278 (N_7278,N_2604,N_843);
or U7279 (N_7279,N_356,N_1694);
nand U7280 (N_7280,N_1336,N_1526);
nand U7281 (N_7281,N_2191,N_1356);
nand U7282 (N_7282,N_209,N_1619);
nand U7283 (N_7283,N_2868,N_4693);
nor U7284 (N_7284,N_3130,N_3452);
nand U7285 (N_7285,N_1503,N_2810);
nor U7286 (N_7286,N_47,N_207);
xor U7287 (N_7287,N_3449,N_2011);
nand U7288 (N_7288,N_483,N_3624);
nor U7289 (N_7289,N_3731,N_258);
xor U7290 (N_7290,N_1398,N_3031);
nor U7291 (N_7291,N_2289,N_3378);
and U7292 (N_7292,N_422,N_3800);
nand U7293 (N_7293,N_2482,N_271);
nor U7294 (N_7294,N_1873,N_1101);
nand U7295 (N_7295,N_382,N_4887);
and U7296 (N_7296,N_4217,N_2862);
nor U7297 (N_7297,N_4914,N_3718);
or U7298 (N_7298,N_2915,N_2658);
or U7299 (N_7299,N_2652,N_4662);
or U7300 (N_7300,N_4029,N_3074);
nand U7301 (N_7301,N_3042,N_3115);
nand U7302 (N_7302,N_3750,N_2513);
xor U7303 (N_7303,N_2949,N_504);
nand U7304 (N_7304,N_2719,N_4573);
xnor U7305 (N_7305,N_277,N_3959);
and U7306 (N_7306,N_650,N_619);
nor U7307 (N_7307,N_1609,N_4279);
and U7308 (N_7308,N_2602,N_4580);
or U7309 (N_7309,N_4410,N_302);
or U7310 (N_7310,N_1744,N_2973);
or U7311 (N_7311,N_4001,N_2399);
xor U7312 (N_7312,N_2508,N_4566);
or U7313 (N_7313,N_2566,N_1962);
nand U7314 (N_7314,N_2404,N_799);
and U7315 (N_7315,N_3830,N_2977);
xnor U7316 (N_7316,N_3095,N_748);
nand U7317 (N_7317,N_1879,N_179);
or U7318 (N_7318,N_4598,N_1799);
xor U7319 (N_7319,N_1031,N_1513);
nand U7320 (N_7320,N_128,N_2414);
nand U7321 (N_7321,N_2218,N_4485);
or U7322 (N_7322,N_2249,N_1276);
nand U7323 (N_7323,N_4525,N_1857);
nand U7324 (N_7324,N_3577,N_3980);
and U7325 (N_7325,N_3635,N_2033);
xor U7326 (N_7326,N_2100,N_4577);
nor U7327 (N_7327,N_3639,N_2762);
nand U7328 (N_7328,N_4053,N_1118);
nor U7329 (N_7329,N_3451,N_4033);
nor U7330 (N_7330,N_1208,N_2653);
and U7331 (N_7331,N_1695,N_2516);
xnor U7332 (N_7332,N_1436,N_3164);
xnor U7333 (N_7333,N_3947,N_471);
nor U7334 (N_7334,N_2779,N_1357);
nor U7335 (N_7335,N_2551,N_897);
nand U7336 (N_7336,N_1903,N_3825);
xnor U7337 (N_7337,N_2722,N_1344);
nand U7338 (N_7338,N_4886,N_3492);
or U7339 (N_7339,N_4488,N_974);
and U7340 (N_7340,N_3945,N_1896);
or U7341 (N_7341,N_262,N_3714);
nor U7342 (N_7342,N_4140,N_3526);
nand U7343 (N_7343,N_4151,N_2310);
and U7344 (N_7344,N_481,N_1232);
xnor U7345 (N_7345,N_4558,N_2944);
nor U7346 (N_7346,N_2951,N_1620);
and U7347 (N_7347,N_943,N_22);
nand U7348 (N_7348,N_4043,N_4917);
or U7349 (N_7349,N_3542,N_4524);
nor U7350 (N_7350,N_2924,N_255);
xor U7351 (N_7351,N_1666,N_2183);
or U7352 (N_7352,N_4683,N_2627);
nand U7353 (N_7353,N_1563,N_4450);
nand U7354 (N_7354,N_2706,N_4504);
nor U7355 (N_7355,N_2601,N_4624);
and U7356 (N_7356,N_3605,N_371);
or U7357 (N_7357,N_2834,N_1610);
nand U7358 (N_7358,N_1980,N_1102);
nand U7359 (N_7359,N_947,N_787);
or U7360 (N_7360,N_4606,N_2897);
nand U7361 (N_7361,N_1487,N_1037);
nor U7362 (N_7362,N_4890,N_3062);
nor U7363 (N_7363,N_113,N_4103);
or U7364 (N_7364,N_1989,N_3430);
nand U7365 (N_7365,N_4385,N_4289);
or U7366 (N_7366,N_418,N_1613);
nand U7367 (N_7367,N_2814,N_3251);
nand U7368 (N_7368,N_4459,N_4875);
nand U7369 (N_7369,N_3469,N_4672);
or U7370 (N_7370,N_2017,N_323);
and U7371 (N_7371,N_4291,N_1303);
nor U7372 (N_7372,N_3228,N_1710);
nand U7373 (N_7373,N_1045,N_133);
or U7374 (N_7374,N_3383,N_1472);
nand U7375 (N_7375,N_4948,N_3933);
xor U7376 (N_7376,N_4695,N_248);
or U7377 (N_7377,N_1640,N_1312);
and U7378 (N_7378,N_278,N_264);
and U7379 (N_7379,N_1496,N_2891);
or U7380 (N_7380,N_1309,N_2364);
nor U7381 (N_7381,N_3401,N_558);
or U7382 (N_7382,N_1165,N_1409);
or U7383 (N_7383,N_1949,N_3058);
or U7384 (N_7384,N_2500,N_4494);
and U7385 (N_7385,N_609,N_4714);
nor U7386 (N_7386,N_878,N_1326);
nor U7387 (N_7387,N_2912,N_2846);
and U7388 (N_7388,N_2979,N_2637);
nand U7389 (N_7389,N_4181,N_3634);
nand U7390 (N_7390,N_2581,N_3413);
nor U7391 (N_7391,N_1580,N_2628);
nand U7392 (N_7392,N_3698,N_4647);
nor U7393 (N_7393,N_4344,N_4747);
and U7394 (N_7394,N_659,N_1366);
nand U7395 (N_7395,N_4280,N_838);
or U7396 (N_7396,N_3597,N_4069);
nand U7397 (N_7397,N_3571,N_3066);
nor U7398 (N_7398,N_2800,N_2344);
or U7399 (N_7399,N_2507,N_3619);
nand U7400 (N_7400,N_9,N_3737);
nor U7401 (N_7401,N_1113,N_4902);
nor U7402 (N_7402,N_782,N_2437);
and U7403 (N_7403,N_3372,N_3904);
and U7404 (N_7404,N_1521,N_4038);
or U7405 (N_7405,N_4585,N_487);
xnor U7406 (N_7406,N_2544,N_3872);
xnor U7407 (N_7407,N_1315,N_774);
nor U7408 (N_7408,N_1691,N_735);
and U7409 (N_7409,N_4901,N_3812);
xor U7410 (N_7410,N_2975,N_4116);
or U7411 (N_7411,N_4245,N_3475);
or U7412 (N_7412,N_288,N_3558);
nor U7413 (N_7413,N_4438,N_4777);
or U7414 (N_7414,N_4319,N_2771);
or U7415 (N_7415,N_1035,N_3009);
and U7416 (N_7416,N_1002,N_2263);
and U7417 (N_7417,N_3834,N_676);
xnor U7418 (N_7418,N_1438,N_4608);
and U7419 (N_7419,N_2367,N_303);
nor U7420 (N_7420,N_367,N_3656);
and U7421 (N_7421,N_3937,N_109);
or U7422 (N_7422,N_3916,N_1622);
xor U7423 (N_7423,N_3375,N_3532);
or U7424 (N_7424,N_4277,N_527);
nand U7425 (N_7425,N_1218,N_1147);
xor U7426 (N_7426,N_1292,N_2116);
or U7427 (N_7427,N_3910,N_3414);
nor U7428 (N_7428,N_2406,N_4373);
nor U7429 (N_7429,N_505,N_3601);
or U7430 (N_7430,N_3117,N_755);
or U7431 (N_7431,N_1781,N_3321);
and U7432 (N_7432,N_960,N_1674);
and U7433 (N_7433,N_1038,N_1382);
nand U7434 (N_7434,N_4179,N_684);
or U7435 (N_7435,N_3432,N_902);
xnor U7436 (N_7436,N_641,N_2390);
nand U7437 (N_7437,N_1752,N_2003);
nand U7438 (N_7438,N_339,N_564);
and U7439 (N_7439,N_3563,N_2750);
nor U7440 (N_7440,N_1658,N_3461);
or U7441 (N_7441,N_3787,N_2457);
and U7442 (N_7442,N_3057,N_472);
and U7443 (N_7443,N_1571,N_2219);
and U7444 (N_7444,N_3419,N_1705);
and U7445 (N_7445,N_4744,N_1846);
nand U7446 (N_7446,N_2018,N_217);
or U7447 (N_7447,N_205,N_2312);
xnor U7448 (N_7448,N_3278,N_3298);
and U7449 (N_7449,N_305,N_671);
and U7450 (N_7450,N_3448,N_338);
and U7451 (N_7451,N_4512,N_1328);
nor U7452 (N_7452,N_4465,N_2626);
xnor U7453 (N_7453,N_2490,N_157);
and U7454 (N_7454,N_984,N_4911);
nand U7455 (N_7455,N_1346,N_3995);
nor U7456 (N_7456,N_4275,N_238);
nor U7457 (N_7457,N_791,N_3090);
xnor U7458 (N_7458,N_3852,N_3498);
xor U7459 (N_7459,N_4708,N_1933);
nor U7460 (N_7460,N_2711,N_1914);
or U7461 (N_7461,N_4372,N_499);
nand U7462 (N_7462,N_357,N_3810);
or U7463 (N_7463,N_839,N_482);
nand U7464 (N_7464,N_3335,N_2050);
or U7465 (N_7465,N_1182,N_1738);
nand U7466 (N_7466,N_1108,N_1821);
xor U7467 (N_7467,N_2827,N_187);
or U7468 (N_7468,N_1958,N_3722);
or U7469 (N_7469,N_4294,N_2005);
nor U7470 (N_7470,N_4774,N_931);
or U7471 (N_7471,N_3653,N_522);
or U7472 (N_7472,N_2417,N_4376);
nand U7473 (N_7473,N_1796,N_4625);
nand U7474 (N_7474,N_965,N_3097);
and U7475 (N_7475,N_3198,N_828);
nor U7476 (N_7476,N_4942,N_3238);
nand U7477 (N_7477,N_4166,N_86);
nor U7478 (N_7478,N_1015,N_2656);
and U7479 (N_7479,N_3222,N_4760);
nor U7480 (N_7480,N_4183,N_1649);
nor U7481 (N_7481,N_4460,N_269);
nand U7482 (N_7482,N_4988,N_1365);
and U7483 (N_7483,N_1604,N_2440);
xnor U7484 (N_7484,N_437,N_763);
nand U7485 (N_7485,N_2670,N_2766);
nor U7486 (N_7486,N_4665,N_2962);
nand U7487 (N_7487,N_4928,N_2243);
and U7488 (N_7488,N_2497,N_796);
nor U7489 (N_7489,N_1718,N_2964);
nand U7490 (N_7490,N_3957,N_2158);
or U7491 (N_7491,N_1632,N_2657);
and U7492 (N_7492,N_2820,N_645);
nor U7493 (N_7493,N_876,N_4578);
and U7494 (N_7494,N_713,N_2321);
or U7495 (N_7495,N_2090,N_4127);
nor U7496 (N_7496,N_535,N_4107);
nand U7497 (N_7497,N_832,N_2184);
nor U7498 (N_7498,N_4035,N_4253);
xnor U7499 (N_7499,N_3479,N_545);
and U7500 (N_7500,N_1250,N_330);
nand U7501 (N_7501,N_738,N_4562);
xor U7502 (N_7502,N_2813,N_2061);
or U7503 (N_7503,N_4358,N_3579);
nand U7504 (N_7504,N_3354,N_3671);
or U7505 (N_7505,N_3018,N_281);
and U7506 (N_7506,N_1335,N_2818);
or U7507 (N_7507,N_1111,N_442);
xnor U7508 (N_7508,N_1714,N_3139);
and U7509 (N_7509,N_495,N_1641);
nand U7510 (N_7510,N_799,N_1026);
nor U7511 (N_7511,N_4673,N_4458);
nand U7512 (N_7512,N_4782,N_4895);
nand U7513 (N_7513,N_2910,N_224);
nor U7514 (N_7514,N_1952,N_1751);
and U7515 (N_7515,N_441,N_4411);
nand U7516 (N_7516,N_4657,N_2155);
and U7517 (N_7517,N_2109,N_3986);
nand U7518 (N_7518,N_3278,N_2423);
and U7519 (N_7519,N_2328,N_1619);
or U7520 (N_7520,N_1816,N_1402);
and U7521 (N_7521,N_650,N_1486);
nor U7522 (N_7522,N_4844,N_3082);
or U7523 (N_7523,N_4166,N_1398);
or U7524 (N_7524,N_1919,N_2451);
nand U7525 (N_7525,N_2362,N_1634);
nand U7526 (N_7526,N_4999,N_1774);
and U7527 (N_7527,N_778,N_4401);
xnor U7528 (N_7528,N_3284,N_2818);
and U7529 (N_7529,N_4828,N_3641);
nor U7530 (N_7530,N_2133,N_1496);
and U7531 (N_7531,N_2502,N_2966);
nand U7532 (N_7532,N_2786,N_4500);
nand U7533 (N_7533,N_4743,N_2280);
nand U7534 (N_7534,N_263,N_4945);
xnor U7535 (N_7535,N_1886,N_2367);
nand U7536 (N_7536,N_855,N_1805);
nand U7537 (N_7537,N_4263,N_1182);
or U7538 (N_7538,N_289,N_4614);
nand U7539 (N_7539,N_540,N_2896);
xor U7540 (N_7540,N_2729,N_1066);
nand U7541 (N_7541,N_4319,N_1382);
or U7542 (N_7542,N_2566,N_1181);
xnor U7543 (N_7543,N_4192,N_3708);
nor U7544 (N_7544,N_4005,N_1620);
and U7545 (N_7545,N_3871,N_1905);
and U7546 (N_7546,N_4810,N_2969);
or U7547 (N_7547,N_896,N_1031);
or U7548 (N_7548,N_4351,N_4735);
nor U7549 (N_7549,N_25,N_3644);
or U7550 (N_7550,N_4355,N_3639);
or U7551 (N_7551,N_2495,N_2931);
xor U7552 (N_7552,N_2934,N_241);
and U7553 (N_7553,N_3133,N_696);
nand U7554 (N_7554,N_1072,N_827);
nor U7555 (N_7555,N_1093,N_402);
nand U7556 (N_7556,N_1639,N_2940);
or U7557 (N_7557,N_2189,N_2863);
and U7558 (N_7558,N_1919,N_4902);
xor U7559 (N_7559,N_1516,N_3161);
or U7560 (N_7560,N_1184,N_1537);
nand U7561 (N_7561,N_1115,N_627);
and U7562 (N_7562,N_1393,N_4809);
nand U7563 (N_7563,N_1505,N_1286);
nor U7564 (N_7564,N_3706,N_3254);
or U7565 (N_7565,N_917,N_4111);
xor U7566 (N_7566,N_2333,N_870);
or U7567 (N_7567,N_4010,N_3793);
or U7568 (N_7568,N_871,N_664);
nor U7569 (N_7569,N_1059,N_4343);
nand U7570 (N_7570,N_133,N_3218);
or U7571 (N_7571,N_4738,N_4797);
and U7572 (N_7572,N_4940,N_4651);
nand U7573 (N_7573,N_494,N_4675);
or U7574 (N_7574,N_4525,N_3808);
nor U7575 (N_7575,N_4111,N_1628);
nor U7576 (N_7576,N_2779,N_4588);
nor U7577 (N_7577,N_2991,N_2219);
nand U7578 (N_7578,N_2166,N_71);
or U7579 (N_7579,N_2395,N_3478);
and U7580 (N_7580,N_3427,N_491);
nor U7581 (N_7581,N_4641,N_888);
nand U7582 (N_7582,N_3879,N_1133);
nor U7583 (N_7583,N_442,N_1289);
and U7584 (N_7584,N_2407,N_313);
or U7585 (N_7585,N_3627,N_903);
or U7586 (N_7586,N_1848,N_1508);
nand U7587 (N_7587,N_3389,N_4752);
nor U7588 (N_7588,N_397,N_3361);
nor U7589 (N_7589,N_1370,N_1369);
nor U7590 (N_7590,N_2607,N_57);
nand U7591 (N_7591,N_2512,N_1292);
nand U7592 (N_7592,N_4701,N_3936);
nand U7593 (N_7593,N_2408,N_2955);
nand U7594 (N_7594,N_3692,N_765);
nor U7595 (N_7595,N_3431,N_4670);
xnor U7596 (N_7596,N_3200,N_2543);
nor U7597 (N_7597,N_595,N_1217);
nor U7598 (N_7598,N_2080,N_4680);
or U7599 (N_7599,N_1635,N_3515);
nor U7600 (N_7600,N_2030,N_1659);
nand U7601 (N_7601,N_3903,N_0);
and U7602 (N_7602,N_2735,N_2617);
or U7603 (N_7603,N_3975,N_3424);
and U7604 (N_7604,N_557,N_1601);
nand U7605 (N_7605,N_3008,N_740);
or U7606 (N_7606,N_3402,N_4164);
xnor U7607 (N_7607,N_4013,N_3502);
nand U7608 (N_7608,N_801,N_1116);
nand U7609 (N_7609,N_1906,N_2331);
nand U7610 (N_7610,N_99,N_4395);
nor U7611 (N_7611,N_4975,N_956);
xor U7612 (N_7612,N_2946,N_3542);
and U7613 (N_7613,N_812,N_2129);
xnor U7614 (N_7614,N_601,N_4874);
or U7615 (N_7615,N_35,N_2534);
and U7616 (N_7616,N_2236,N_4887);
and U7617 (N_7617,N_2825,N_2160);
nand U7618 (N_7618,N_341,N_2404);
or U7619 (N_7619,N_2865,N_2423);
nand U7620 (N_7620,N_2437,N_337);
and U7621 (N_7621,N_431,N_2742);
xnor U7622 (N_7622,N_2927,N_54);
or U7623 (N_7623,N_364,N_2275);
nor U7624 (N_7624,N_4228,N_4550);
and U7625 (N_7625,N_4158,N_1580);
and U7626 (N_7626,N_1843,N_539);
or U7627 (N_7627,N_3305,N_2444);
or U7628 (N_7628,N_4814,N_1666);
nor U7629 (N_7629,N_3260,N_3018);
nand U7630 (N_7630,N_240,N_2396);
and U7631 (N_7631,N_328,N_3469);
and U7632 (N_7632,N_3607,N_3956);
and U7633 (N_7633,N_1971,N_2215);
and U7634 (N_7634,N_759,N_2224);
nand U7635 (N_7635,N_4158,N_1013);
nand U7636 (N_7636,N_3207,N_1957);
nand U7637 (N_7637,N_1133,N_2255);
and U7638 (N_7638,N_1497,N_3421);
nand U7639 (N_7639,N_509,N_2227);
nor U7640 (N_7640,N_579,N_3832);
nor U7641 (N_7641,N_4551,N_2325);
or U7642 (N_7642,N_4225,N_1490);
and U7643 (N_7643,N_3896,N_2485);
nor U7644 (N_7644,N_885,N_1360);
nand U7645 (N_7645,N_3150,N_3322);
and U7646 (N_7646,N_16,N_747);
nor U7647 (N_7647,N_3978,N_2646);
and U7648 (N_7648,N_3560,N_2164);
or U7649 (N_7649,N_3728,N_385);
or U7650 (N_7650,N_602,N_4694);
and U7651 (N_7651,N_779,N_901);
nand U7652 (N_7652,N_2933,N_3647);
or U7653 (N_7653,N_399,N_1015);
or U7654 (N_7654,N_3788,N_4915);
or U7655 (N_7655,N_4835,N_1380);
or U7656 (N_7656,N_4762,N_4997);
nor U7657 (N_7657,N_3036,N_4431);
xnor U7658 (N_7658,N_4527,N_1689);
nand U7659 (N_7659,N_3154,N_2325);
and U7660 (N_7660,N_2099,N_1313);
xor U7661 (N_7661,N_371,N_3597);
nor U7662 (N_7662,N_1171,N_376);
nor U7663 (N_7663,N_2411,N_3931);
nand U7664 (N_7664,N_4148,N_2527);
nor U7665 (N_7665,N_4230,N_3623);
or U7666 (N_7666,N_3951,N_3687);
xor U7667 (N_7667,N_3278,N_3710);
or U7668 (N_7668,N_2043,N_1512);
nand U7669 (N_7669,N_4883,N_2025);
or U7670 (N_7670,N_4591,N_3672);
and U7671 (N_7671,N_4658,N_605);
and U7672 (N_7672,N_2231,N_1367);
and U7673 (N_7673,N_2034,N_3468);
or U7674 (N_7674,N_2447,N_4235);
and U7675 (N_7675,N_3789,N_178);
and U7676 (N_7676,N_2460,N_2320);
nor U7677 (N_7677,N_1799,N_867);
or U7678 (N_7678,N_1736,N_4500);
and U7679 (N_7679,N_1445,N_1789);
and U7680 (N_7680,N_1105,N_2142);
or U7681 (N_7681,N_4881,N_681);
nand U7682 (N_7682,N_2525,N_1290);
nand U7683 (N_7683,N_3964,N_1809);
and U7684 (N_7684,N_3752,N_1340);
nand U7685 (N_7685,N_3577,N_1659);
nand U7686 (N_7686,N_702,N_1920);
or U7687 (N_7687,N_1186,N_4897);
nor U7688 (N_7688,N_4605,N_3695);
and U7689 (N_7689,N_2333,N_2388);
nor U7690 (N_7690,N_3285,N_3383);
nand U7691 (N_7691,N_4821,N_1388);
nand U7692 (N_7692,N_3972,N_4494);
and U7693 (N_7693,N_398,N_588);
nor U7694 (N_7694,N_1235,N_508);
or U7695 (N_7695,N_421,N_2556);
or U7696 (N_7696,N_2890,N_420);
and U7697 (N_7697,N_4782,N_1352);
nand U7698 (N_7698,N_4130,N_1637);
nor U7699 (N_7699,N_4637,N_4712);
xor U7700 (N_7700,N_613,N_4527);
nor U7701 (N_7701,N_4809,N_2959);
or U7702 (N_7702,N_4778,N_2091);
nand U7703 (N_7703,N_4763,N_4538);
nand U7704 (N_7704,N_2434,N_1063);
or U7705 (N_7705,N_1742,N_59);
nand U7706 (N_7706,N_2280,N_903);
and U7707 (N_7707,N_2182,N_4050);
and U7708 (N_7708,N_4630,N_2414);
nand U7709 (N_7709,N_2605,N_2938);
nor U7710 (N_7710,N_1356,N_4294);
nand U7711 (N_7711,N_740,N_4326);
nor U7712 (N_7712,N_2551,N_3148);
nand U7713 (N_7713,N_3069,N_2897);
nand U7714 (N_7714,N_352,N_3527);
nor U7715 (N_7715,N_712,N_3783);
xnor U7716 (N_7716,N_2923,N_3774);
nand U7717 (N_7717,N_1650,N_1211);
or U7718 (N_7718,N_42,N_1969);
xnor U7719 (N_7719,N_513,N_2833);
and U7720 (N_7720,N_4188,N_1207);
and U7721 (N_7721,N_4872,N_960);
or U7722 (N_7722,N_560,N_4762);
or U7723 (N_7723,N_334,N_4491);
nor U7724 (N_7724,N_1189,N_2513);
nor U7725 (N_7725,N_3771,N_63);
xnor U7726 (N_7726,N_3501,N_4600);
nor U7727 (N_7727,N_942,N_2339);
or U7728 (N_7728,N_2598,N_2835);
or U7729 (N_7729,N_1599,N_3666);
nand U7730 (N_7730,N_2024,N_4578);
nand U7731 (N_7731,N_2510,N_2574);
and U7732 (N_7732,N_4663,N_3282);
nand U7733 (N_7733,N_4884,N_2482);
nor U7734 (N_7734,N_1247,N_2820);
or U7735 (N_7735,N_450,N_2453);
or U7736 (N_7736,N_3163,N_2249);
and U7737 (N_7737,N_3999,N_2098);
or U7738 (N_7738,N_1470,N_4307);
and U7739 (N_7739,N_3205,N_545);
nor U7740 (N_7740,N_1781,N_3461);
or U7741 (N_7741,N_3559,N_4978);
or U7742 (N_7742,N_396,N_3461);
xnor U7743 (N_7743,N_392,N_2839);
or U7744 (N_7744,N_3555,N_2109);
and U7745 (N_7745,N_3348,N_4580);
nand U7746 (N_7746,N_2205,N_3442);
xnor U7747 (N_7747,N_932,N_1645);
or U7748 (N_7748,N_114,N_4217);
nand U7749 (N_7749,N_3975,N_4383);
or U7750 (N_7750,N_3507,N_4894);
or U7751 (N_7751,N_4977,N_1023);
and U7752 (N_7752,N_4744,N_2696);
xnor U7753 (N_7753,N_1029,N_3449);
xnor U7754 (N_7754,N_3281,N_2232);
or U7755 (N_7755,N_2405,N_1518);
nor U7756 (N_7756,N_1333,N_3534);
nand U7757 (N_7757,N_1243,N_3999);
nor U7758 (N_7758,N_649,N_762);
and U7759 (N_7759,N_1011,N_3458);
and U7760 (N_7760,N_940,N_1493);
nand U7761 (N_7761,N_3477,N_1830);
and U7762 (N_7762,N_2621,N_1740);
or U7763 (N_7763,N_2050,N_4231);
nor U7764 (N_7764,N_2068,N_1866);
or U7765 (N_7765,N_2775,N_2683);
nor U7766 (N_7766,N_1549,N_1922);
nor U7767 (N_7767,N_4262,N_3398);
nor U7768 (N_7768,N_802,N_3400);
or U7769 (N_7769,N_4415,N_3834);
and U7770 (N_7770,N_112,N_65);
or U7771 (N_7771,N_3172,N_2770);
or U7772 (N_7772,N_1289,N_3833);
and U7773 (N_7773,N_2099,N_126);
and U7774 (N_7774,N_2765,N_3313);
nor U7775 (N_7775,N_4564,N_4945);
or U7776 (N_7776,N_2934,N_4187);
and U7777 (N_7777,N_4139,N_3174);
and U7778 (N_7778,N_1979,N_4355);
and U7779 (N_7779,N_95,N_2813);
and U7780 (N_7780,N_2907,N_722);
or U7781 (N_7781,N_4442,N_2022);
nand U7782 (N_7782,N_2819,N_1950);
and U7783 (N_7783,N_3952,N_1319);
nand U7784 (N_7784,N_1585,N_2297);
nor U7785 (N_7785,N_4676,N_651);
nor U7786 (N_7786,N_435,N_1339);
xnor U7787 (N_7787,N_4201,N_2475);
nand U7788 (N_7788,N_883,N_473);
or U7789 (N_7789,N_1495,N_4855);
xnor U7790 (N_7790,N_1820,N_101);
and U7791 (N_7791,N_1248,N_1341);
nor U7792 (N_7792,N_2613,N_4161);
and U7793 (N_7793,N_4452,N_4280);
or U7794 (N_7794,N_4643,N_4945);
nand U7795 (N_7795,N_219,N_4053);
and U7796 (N_7796,N_1523,N_703);
nor U7797 (N_7797,N_3327,N_2924);
and U7798 (N_7798,N_3115,N_1224);
nor U7799 (N_7799,N_2556,N_136);
xor U7800 (N_7800,N_356,N_3756);
or U7801 (N_7801,N_1103,N_978);
or U7802 (N_7802,N_407,N_947);
or U7803 (N_7803,N_366,N_1820);
xnor U7804 (N_7804,N_849,N_4186);
or U7805 (N_7805,N_1708,N_3547);
nand U7806 (N_7806,N_2721,N_1464);
nor U7807 (N_7807,N_171,N_3579);
nand U7808 (N_7808,N_1275,N_3006);
nor U7809 (N_7809,N_2021,N_1547);
xnor U7810 (N_7810,N_4712,N_2819);
xor U7811 (N_7811,N_1797,N_2788);
xnor U7812 (N_7812,N_1911,N_3783);
nor U7813 (N_7813,N_4946,N_2056);
nand U7814 (N_7814,N_924,N_1969);
or U7815 (N_7815,N_4846,N_168);
xnor U7816 (N_7816,N_2080,N_45);
or U7817 (N_7817,N_4827,N_3830);
nand U7818 (N_7818,N_3505,N_3317);
nor U7819 (N_7819,N_302,N_1668);
or U7820 (N_7820,N_2683,N_4780);
nor U7821 (N_7821,N_1112,N_746);
or U7822 (N_7822,N_1664,N_1438);
xor U7823 (N_7823,N_3176,N_957);
or U7824 (N_7824,N_3412,N_4655);
xnor U7825 (N_7825,N_4675,N_2092);
or U7826 (N_7826,N_4213,N_380);
nor U7827 (N_7827,N_1644,N_3032);
nor U7828 (N_7828,N_3094,N_809);
and U7829 (N_7829,N_4122,N_1212);
nand U7830 (N_7830,N_4366,N_3205);
or U7831 (N_7831,N_1189,N_1827);
xnor U7832 (N_7832,N_2962,N_2845);
and U7833 (N_7833,N_3172,N_4842);
and U7834 (N_7834,N_3737,N_260);
or U7835 (N_7835,N_3508,N_3546);
nor U7836 (N_7836,N_3154,N_2534);
xnor U7837 (N_7837,N_2528,N_3785);
or U7838 (N_7838,N_3557,N_4407);
nand U7839 (N_7839,N_1035,N_4464);
or U7840 (N_7840,N_2275,N_2597);
xor U7841 (N_7841,N_3456,N_3362);
and U7842 (N_7842,N_1323,N_2536);
and U7843 (N_7843,N_1399,N_1907);
nor U7844 (N_7844,N_1631,N_4208);
xnor U7845 (N_7845,N_2357,N_987);
nor U7846 (N_7846,N_389,N_2049);
nand U7847 (N_7847,N_4484,N_517);
and U7848 (N_7848,N_4352,N_1066);
and U7849 (N_7849,N_245,N_4775);
nor U7850 (N_7850,N_2831,N_1552);
nand U7851 (N_7851,N_1694,N_2430);
nand U7852 (N_7852,N_4552,N_3674);
or U7853 (N_7853,N_3379,N_2310);
nand U7854 (N_7854,N_4219,N_2218);
or U7855 (N_7855,N_4603,N_1634);
or U7856 (N_7856,N_520,N_3974);
nand U7857 (N_7857,N_2046,N_1519);
xnor U7858 (N_7858,N_1383,N_1826);
nand U7859 (N_7859,N_3521,N_3300);
and U7860 (N_7860,N_3844,N_4996);
xnor U7861 (N_7861,N_3577,N_3475);
and U7862 (N_7862,N_4654,N_4402);
nand U7863 (N_7863,N_3905,N_4510);
nand U7864 (N_7864,N_1791,N_3372);
nand U7865 (N_7865,N_3276,N_2862);
nand U7866 (N_7866,N_4433,N_3889);
nor U7867 (N_7867,N_2075,N_4981);
nor U7868 (N_7868,N_2334,N_4783);
or U7869 (N_7869,N_3009,N_572);
nand U7870 (N_7870,N_969,N_3181);
xnor U7871 (N_7871,N_2896,N_3595);
nand U7872 (N_7872,N_2364,N_1881);
xor U7873 (N_7873,N_4201,N_3339);
nand U7874 (N_7874,N_2629,N_3008);
nor U7875 (N_7875,N_1469,N_817);
and U7876 (N_7876,N_665,N_2712);
nand U7877 (N_7877,N_4846,N_4606);
or U7878 (N_7878,N_3468,N_3016);
nand U7879 (N_7879,N_235,N_3296);
or U7880 (N_7880,N_4159,N_3379);
nor U7881 (N_7881,N_1573,N_1982);
nand U7882 (N_7882,N_2992,N_4359);
or U7883 (N_7883,N_903,N_2449);
nor U7884 (N_7884,N_4916,N_2465);
nor U7885 (N_7885,N_4224,N_2226);
nor U7886 (N_7886,N_1307,N_1266);
nor U7887 (N_7887,N_1300,N_282);
nor U7888 (N_7888,N_4054,N_700);
and U7889 (N_7889,N_1590,N_700);
or U7890 (N_7890,N_480,N_3617);
xor U7891 (N_7891,N_4046,N_1655);
xnor U7892 (N_7892,N_4731,N_2740);
or U7893 (N_7893,N_1828,N_4875);
or U7894 (N_7894,N_4846,N_1773);
or U7895 (N_7895,N_4156,N_3555);
nand U7896 (N_7896,N_1090,N_424);
nand U7897 (N_7897,N_3771,N_2042);
nor U7898 (N_7898,N_125,N_895);
nor U7899 (N_7899,N_1200,N_1391);
and U7900 (N_7900,N_3218,N_2674);
nand U7901 (N_7901,N_2346,N_1006);
nor U7902 (N_7902,N_3277,N_4280);
or U7903 (N_7903,N_3327,N_1104);
or U7904 (N_7904,N_3128,N_127);
nand U7905 (N_7905,N_2360,N_1723);
and U7906 (N_7906,N_4295,N_265);
and U7907 (N_7907,N_97,N_4774);
xor U7908 (N_7908,N_2800,N_3960);
nand U7909 (N_7909,N_4778,N_4406);
nor U7910 (N_7910,N_3556,N_1456);
or U7911 (N_7911,N_2860,N_1110);
nand U7912 (N_7912,N_4239,N_3604);
and U7913 (N_7913,N_4072,N_2219);
nor U7914 (N_7914,N_4769,N_764);
and U7915 (N_7915,N_410,N_1448);
nand U7916 (N_7916,N_223,N_834);
nor U7917 (N_7917,N_2528,N_4660);
and U7918 (N_7918,N_634,N_3740);
nand U7919 (N_7919,N_4509,N_3358);
and U7920 (N_7920,N_588,N_3619);
nand U7921 (N_7921,N_506,N_3856);
nand U7922 (N_7922,N_364,N_2263);
nor U7923 (N_7923,N_502,N_3358);
nand U7924 (N_7924,N_2726,N_3665);
xor U7925 (N_7925,N_3445,N_2577);
or U7926 (N_7926,N_4205,N_595);
or U7927 (N_7927,N_2364,N_3487);
nor U7928 (N_7928,N_1045,N_3974);
nor U7929 (N_7929,N_3589,N_4002);
nand U7930 (N_7930,N_2123,N_2568);
xor U7931 (N_7931,N_2200,N_4472);
nand U7932 (N_7932,N_3389,N_3150);
and U7933 (N_7933,N_376,N_2612);
and U7934 (N_7934,N_2766,N_1510);
xnor U7935 (N_7935,N_308,N_1812);
and U7936 (N_7936,N_1013,N_4357);
and U7937 (N_7937,N_4521,N_1100);
or U7938 (N_7938,N_2613,N_1473);
nand U7939 (N_7939,N_3887,N_4082);
and U7940 (N_7940,N_1701,N_3379);
or U7941 (N_7941,N_1786,N_4514);
or U7942 (N_7942,N_4179,N_191);
or U7943 (N_7943,N_486,N_6);
nand U7944 (N_7944,N_3513,N_284);
and U7945 (N_7945,N_2264,N_3048);
or U7946 (N_7946,N_811,N_1018);
nor U7947 (N_7947,N_1875,N_3435);
and U7948 (N_7948,N_1639,N_540);
or U7949 (N_7949,N_2485,N_2711);
and U7950 (N_7950,N_53,N_2410);
xor U7951 (N_7951,N_987,N_525);
nand U7952 (N_7952,N_3613,N_658);
nand U7953 (N_7953,N_1215,N_3723);
and U7954 (N_7954,N_1575,N_2488);
nor U7955 (N_7955,N_4087,N_2700);
nand U7956 (N_7956,N_427,N_4590);
and U7957 (N_7957,N_2897,N_2746);
or U7958 (N_7958,N_2634,N_1059);
or U7959 (N_7959,N_290,N_3007);
and U7960 (N_7960,N_4962,N_4616);
xor U7961 (N_7961,N_3020,N_2225);
nor U7962 (N_7962,N_1561,N_1180);
or U7963 (N_7963,N_4950,N_3980);
xor U7964 (N_7964,N_4225,N_3078);
nand U7965 (N_7965,N_3966,N_173);
or U7966 (N_7966,N_4683,N_1963);
and U7967 (N_7967,N_3225,N_1067);
or U7968 (N_7968,N_1100,N_4467);
nand U7969 (N_7969,N_1153,N_3591);
or U7970 (N_7970,N_1024,N_979);
nor U7971 (N_7971,N_2,N_221);
nor U7972 (N_7972,N_4311,N_4212);
or U7973 (N_7973,N_4993,N_243);
nor U7974 (N_7974,N_2200,N_4363);
xnor U7975 (N_7975,N_3685,N_4046);
and U7976 (N_7976,N_4011,N_2066);
or U7977 (N_7977,N_4497,N_2894);
nand U7978 (N_7978,N_4207,N_743);
nand U7979 (N_7979,N_2646,N_1002);
and U7980 (N_7980,N_2508,N_3629);
and U7981 (N_7981,N_2652,N_2265);
and U7982 (N_7982,N_317,N_682);
nor U7983 (N_7983,N_724,N_4118);
nand U7984 (N_7984,N_576,N_966);
nor U7985 (N_7985,N_324,N_1908);
and U7986 (N_7986,N_2774,N_462);
xor U7987 (N_7987,N_565,N_4571);
nand U7988 (N_7988,N_523,N_91);
nor U7989 (N_7989,N_1097,N_3814);
nor U7990 (N_7990,N_2026,N_3921);
nor U7991 (N_7991,N_1563,N_1994);
xor U7992 (N_7992,N_3795,N_4141);
nor U7993 (N_7993,N_4136,N_1536);
nor U7994 (N_7994,N_4312,N_2611);
nand U7995 (N_7995,N_2148,N_3666);
nand U7996 (N_7996,N_3121,N_4481);
or U7997 (N_7997,N_152,N_1662);
nor U7998 (N_7998,N_3304,N_4608);
and U7999 (N_7999,N_2512,N_2148);
and U8000 (N_8000,N_1003,N_1973);
xor U8001 (N_8001,N_3817,N_2117);
or U8002 (N_8002,N_4252,N_3324);
and U8003 (N_8003,N_1050,N_4240);
nand U8004 (N_8004,N_2894,N_3258);
xnor U8005 (N_8005,N_4277,N_4043);
or U8006 (N_8006,N_1907,N_3872);
nand U8007 (N_8007,N_861,N_3721);
nand U8008 (N_8008,N_3869,N_1157);
and U8009 (N_8009,N_4444,N_4775);
nor U8010 (N_8010,N_2221,N_2832);
nand U8011 (N_8011,N_3289,N_3070);
xor U8012 (N_8012,N_2945,N_1603);
and U8013 (N_8013,N_4022,N_4112);
nor U8014 (N_8014,N_449,N_1703);
nand U8015 (N_8015,N_1069,N_4284);
nor U8016 (N_8016,N_139,N_3560);
nor U8017 (N_8017,N_3753,N_2389);
nand U8018 (N_8018,N_1768,N_2709);
and U8019 (N_8019,N_3454,N_1669);
or U8020 (N_8020,N_1367,N_810);
and U8021 (N_8021,N_3596,N_4418);
nand U8022 (N_8022,N_4216,N_3714);
and U8023 (N_8023,N_225,N_1051);
or U8024 (N_8024,N_1778,N_713);
or U8025 (N_8025,N_2350,N_1167);
nor U8026 (N_8026,N_763,N_4553);
nor U8027 (N_8027,N_1549,N_2034);
nand U8028 (N_8028,N_2345,N_3255);
and U8029 (N_8029,N_1091,N_3004);
nor U8030 (N_8030,N_1856,N_3207);
nand U8031 (N_8031,N_2136,N_1530);
xor U8032 (N_8032,N_4991,N_4429);
or U8033 (N_8033,N_2836,N_1676);
and U8034 (N_8034,N_3670,N_4654);
nand U8035 (N_8035,N_4270,N_3194);
nor U8036 (N_8036,N_1535,N_4110);
and U8037 (N_8037,N_4340,N_4379);
nor U8038 (N_8038,N_1547,N_4069);
and U8039 (N_8039,N_2704,N_1306);
nor U8040 (N_8040,N_264,N_2974);
nor U8041 (N_8041,N_1086,N_4107);
nor U8042 (N_8042,N_3644,N_550);
or U8043 (N_8043,N_882,N_2333);
and U8044 (N_8044,N_4782,N_3496);
nor U8045 (N_8045,N_685,N_1774);
xnor U8046 (N_8046,N_1857,N_4507);
and U8047 (N_8047,N_3205,N_4298);
or U8048 (N_8048,N_3168,N_2317);
or U8049 (N_8049,N_3049,N_3465);
nand U8050 (N_8050,N_3966,N_3598);
xor U8051 (N_8051,N_71,N_1595);
nand U8052 (N_8052,N_2466,N_741);
xnor U8053 (N_8053,N_466,N_186);
and U8054 (N_8054,N_4686,N_2132);
and U8055 (N_8055,N_1321,N_2627);
nand U8056 (N_8056,N_4579,N_3467);
or U8057 (N_8057,N_4613,N_2580);
xor U8058 (N_8058,N_4959,N_4578);
nor U8059 (N_8059,N_2386,N_208);
nand U8060 (N_8060,N_2704,N_2813);
nand U8061 (N_8061,N_4886,N_2923);
xor U8062 (N_8062,N_2269,N_552);
nor U8063 (N_8063,N_2006,N_4352);
nor U8064 (N_8064,N_596,N_2035);
or U8065 (N_8065,N_4552,N_4875);
and U8066 (N_8066,N_3245,N_3640);
xnor U8067 (N_8067,N_143,N_2401);
and U8068 (N_8068,N_217,N_2914);
nand U8069 (N_8069,N_971,N_1413);
nand U8070 (N_8070,N_762,N_2428);
or U8071 (N_8071,N_421,N_4543);
nor U8072 (N_8072,N_3622,N_4289);
nor U8073 (N_8073,N_3835,N_4650);
nor U8074 (N_8074,N_1660,N_3882);
and U8075 (N_8075,N_1064,N_2790);
nand U8076 (N_8076,N_2763,N_2796);
and U8077 (N_8077,N_1884,N_3757);
xnor U8078 (N_8078,N_1116,N_4876);
or U8079 (N_8079,N_2349,N_3427);
and U8080 (N_8080,N_493,N_1455);
nor U8081 (N_8081,N_632,N_701);
nor U8082 (N_8082,N_2320,N_1857);
xor U8083 (N_8083,N_1875,N_17);
nand U8084 (N_8084,N_975,N_3323);
nor U8085 (N_8085,N_3559,N_3716);
nor U8086 (N_8086,N_4946,N_2640);
nand U8087 (N_8087,N_1935,N_2352);
nor U8088 (N_8088,N_4678,N_928);
or U8089 (N_8089,N_40,N_31);
nor U8090 (N_8090,N_791,N_2145);
nor U8091 (N_8091,N_3314,N_1397);
nand U8092 (N_8092,N_820,N_3603);
or U8093 (N_8093,N_1874,N_304);
or U8094 (N_8094,N_3238,N_1997);
or U8095 (N_8095,N_3711,N_2877);
nor U8096 (N_8096,N_1250,N_4598);
or U8097 (N_8097,N_28,N_506);
or U8098 (N_8098,N_409,N_2892);
or U8099 (N_8099,N_1911,N_2954);
or U8100 (N_8100,N_1250,N_1378);
nor U8101 (N_8101,N_67,N_330);
or U8102 (N_8102,N_3130,N_556);
nor U8103 (N_8103,N_4504,N_218);
xor U8104 (N_8104,N_3642,N_283);
and U8105 (N_8105,N_1663,N_320);
nand U8106 (N_8106,N_1301,N_3530);
and U8107 (N_8107,N_2003,N_1364);
nand U8108 (N_8108,N_2850,N_3238);
and U8109 (N_8109,N_3563,N_4422);
nor U8110 (N_8110,N_390,N_721);
nor U8111 (N_8111,N_551,N_285);
nand U8112 (N_8112,N_2726,N_4549);
nor U8113 (N_8113,N_805,N_3907);
nand U8114 (N_8114,N_1,N_4332);
and U8115 (N_8115,N_4730,N_724);
nor U8116 (N_8116,N_3198,N_1127);
nand U8117 (N_8117,N_1719,N_1176);
nand U8118 (N_8118,N_1078,N_290);
or U8119 (N_8119,N_4092,N_2908);
or U8120 (N_8120,N_4010,N_265);
nand U8121 (N_8121,N_1165,N_4349);
and U8122 (N_8122,N_2732,N_2399);
nand U8123 (N_8123,N_3909,N_1929);
and U8124 (N_8124,N_4574,N_376);
and U8125 (N_8125,N_766,N_248);
and U8126 (N_8126,N_2677,N_3573);
nand U8127 (N_8127,N_2434,N_1662);
or U8128 (N_8128,N_55,N_817);
nand U8129 (N_8129,N_1319,N_3498);
or U8130 (N_8130,N_3517,N_3401);
or U8131 (N_8131,N_3682,N_2294);
nor U8132 (N_8132,N_3980,N_3601);
and U8133 (N_8133,N_4823,N_1243);
nor U8134 (N_8134,N_4896,N_2202);
nand U8135 (N_8135,N_1842,N_1874);
nand U8136 (N_8136,N_4422,N_1752);
nor U8137 (N_8137,N_427,N_4213);
nand U8138 (N_8138,N_1299,N_3373);
and U8139 (N_8139,N_1438,N_2205);
or U8140 (N_8140,N_994,N_4947);
or U8141 (N_8141,N_3100,N_1817);
nor U8142 (N_8142,N_4849,N_4427);
or U8143 (N_8143,N_1459,N_2262);
nand U8144 (N_8144,N_2904,N_1559);
or U8145 (N_8145,N_2956,N_321);
nor U8146 (N_8146,N_3011,N_707);
nand U8147 (N_8147,N_2039,N_4165);
and U8148 (N_8148,N_3776,N_2506);
or U8149 (N_8149,N_4253,N_2213);
nand U8150 (N_8150,N_4697,N_463);
nor U8151 (N_8151,N_1222,N_3496);
nor U8152 (N_8152,N_2759,N_80);
and U8153 (N_8153,N_1083,N_1131);
nand U8154 (N_8154,N_296,N_1938);
nand U8155 (N_8155,N_1505,N_4371);
or U8156 (N_8156,N_4891,N_3265);
or U8157 (N_8157,N_1958,N_2039);
xnor U8158 (N_8158,N_3180,N_2310);
and U8159 (N_8159,N_4008,N_3095);
and U8160 (N_8160,N_3741,N_2737);
nor U8161 (N_8161,N_360,N_94);
nand U8162 (N_8162,N_3913,N_4570);
or U8163 (N_8163,N_4873,N_667);
xor U8164 (N_8164,N_2642,N_2429);
nor U8165 (N_8165,N_2519,N_4883);
nand U8166 (N_8166,N_2153,N_4647);
and U8167 (N_8167,N_1688,N_91);
or U8168 (N_8168,N_4090,N_1429);
nand U8169 (N_8169,N_1725,N_575);
and U8170 (N_8170,N_4095,N_2501);
and U8171 (N_8171,N_1560,N_1368);
xnor U8172 (N_8172,N_4447,N_4837);
or U8173 (N_8173,N_2313,N_261);
nor U8174 (N_8174,N_1259,N_2501);
nor U8175 (N_8175,N_217,N_2115);
nor U8176 (N_8176,N_1597,N_3889);
xnor U8177 (N_8177,N_2561,N_529);
nor U8178 (N_8178,N_2005,N_3955);
and U8179 (N_8179,N_3969,N_466);
xnor U8180 (N_8180,N_4240,N_130);
nor U8181 (N_8181,N_433,N_4403);
nand U8182 (N_8182,N_2959,N_2686);
nor U8183 (N_8183,N_37,N_3493);
or U8184 (N_8184,N_212,N_2723);
nand U8185 (N_8185,N_705,N_4332);
nor U8186 (N_8186,N_4126,N_2342);
or U8187 (N_8187,N_3184,N_3210);
or U8188 (N_8188,N_4148,N_2301);
nand U8189 (N_8189,N_145,N_1955);
nand U8190 (N_8190,N_46,N_2841);
xor U8191 (N_8191,N_1746,N_3674);
and U8192 (N_8192,N_1192,N_4226);
nor U8193 (N_8193,N_356,N_1201);
nand U8194 (N_8194,N_443,N_3331);
nand U8195 (N_8195,N_1036,N_2509);
nand U8196 (N_8196,N_3270,N_2844);
and U8197 (N_8197,N_3046,N_2174);
nand U8198 (N_8198,N_4537,N_3452);
xor U8199 (N_8199,N_2877,N_4573);
nand U8200 (N_8200,N_3223,N_2790);
or U8201 (N_8201,N_1733,N_778);
or U8202 (N_8202,N_3804,N_3367);
nor U8203 (N_8203,N_4622,N_2045);
or U8204 (N_8204,N_1484,N_2455);
or U8205 (N_8205,N_94,N_1806);
nor U8206 (N_8206,N_3948,N_812);
and U8207 (N_8207,N_1142,N_3557);
nor U8208 (N_8208,N_1067,N_4004);
nand U8209 (N_8209,N_831,N_357);
nor U8210 (N_8210,N_1325,N_1574);
nand U8211 (N_8211,N_3320,N_4872);
nor U8212 (N_8212,N_377,N_4847);
or U8213 (N_8213,N_224,N_4029);
or U8214 (N_8214,N_3266,N_2569);
xnor U8215 (N_8215,N_4634,N_1879);
or U8216 (N_8216,N_4836,N_3481);
nor U8217 (N_8217,N_3174,N_4825);
xnor U8218 (N_8218,N_4856,N_617);
and U8219 (N_8219,N_3980,N_460);
nand U8220 (N_8220,N_2336,N_4180);
nand U8221 (N_8221,N_4626,N_3935);
nand U8222 (N_8222,N_3042,N_4080);
nand U8223 (N_8223,N_3681,N_1478);
or U8224 (N_8224,N_1240,N_4553);
or U8225 (N_8225,N_3117,N_593);
nand U8226 (N_8226,N_1086,N_1215);
nand U8227 (N_8227,N_4976,N_2788);
and U8228 (N_8228,N_219,N_705);
xor U8229 (N_8229,N_364,N_3768);
nor U8230 (N_8230,N_629,N_1990);
and U8231 (N_8231,N_4293,N_3979);
or U8232 (N_8232,N_228,N_3036);
nand U8233 (N_8233,N_1572,N_3173);
nor U8234 (N_8234,N_3217,N_1327);
xor U8235 (N_8235,N_3817,N_3970);
nand U8236 (N_8236,N_1381,N_4594);
nand U8237 (N_8237,N_4622,N_3213);
and U8238 (N_8238,N_4575,N_2246);
nor U8239 (N_8239,N_2279,N_4186);
nand U8240 (N_8240,N_2446,N_2990);
and U8241 (N_8241,N_3100,N_3135);
or U8242 (N_8242,N_2557,N_1422);
nand U8243 (N_8243,N_4337,N_2167);
nor U8244 (N_8244,N_2313,N_1590);
nand U8245 (N_8245,N_2557,N_3231);
and U8246 (N_8246,N_1164,N_3210);
nand U8247 (N_8247,N_3925,N_4309);
and U8248 (N_8248,N_519,N_1960);
nor U8249 (N_8249,N_4924,N_2182);
or U8250 (N_8250,N_3546,N_1326);
nor U8251 (N_8251,N_2764,N_2072);
or U8252 (N_8252,N_4983,N_2640);
nor U8253 (N_8253,N_1709,N_2430);
xor U8254 (N_8254,N_2109,N_2502);
nor U8255 (N_8255,N_3314,N_3274);
or U8256 (N_8256,N_3106,N_210);
nor U8257 (N_8257,N_4386,N_2045);
nor U8258 (N_8258,N_2710,N_370);
and U8259 (N_8259,N_4237,N_2517);
and U8260 (N_8260,N_2158,N_4926);
nor U8261 (N_8261,N_2,N_3400);
or U8262 (N_8262,N_4609,N_3145);
or U8263 (N_8263,N_3585,N_227);
and U8264 (N_8264,N_3562,N_28);
and U8265 (N_8265,N_3294,N_256);
or U8266 (N_8266,N_3685,N_2808);
or U8267 (N_8267,N_1986,N_3844);
xnor U8268 (N_8268,N_721,N_4879);
and U8269 (N_8269,N_2549,N_1540);
and U8270 (N_8270,N_1014,N_982);
nor U8271 (N_8271,N_3350,N_470);
or U8272 (N_8272,N_3401,N_1720);
and U8273 (N_8273,N_4176,N_3633);
nand U8274 (N_8274,N_1174,N_1415);
and U8275 (N_8275,N_768,N_1728);
nand U8276 (N_8276,N_4301,N_3726);
nand U8277 (N_8277,N_2818,N_2397);
nand U8278 (N_8278,N_4155,N_1200);
nor U8279 (N_8279,N_769,N_4983);
and U8280 (N_8280,N_1760,N_4567);
and U8281 (N_8281,N_4981,N_1494);
and U8282 (N_8282,N_4116,N_2137);
and U8283 (N_8283,N_4967,N_3737);
or U8284 (N_8284,N_2599,N_4671);
or U8285 (N_8285,N_1310,N_2799);
or U8286 (N_8286,N_758,N_1620);
or U8287 (N_8287,N_402,N_4762);
or U8288 (N_8288,N_3628,N_3949);
nor U8289 (N_8289,N_3237,N_1483);
xor U8290 (N_8290,N_3367,N_311);
nor U8291 (N_8291,N_4396,N_4504);
and U8292 (N_8292,N_354,N_1299);
nor U8293 (N_8293,N_3678,N_3518);
or U8294 (N_8294,N_1035,N_3911);
or U8295 (N_8295,N_2395,N_802);
xnor U8296 (N_8296,N_3385,N_4582);
or U8297 (N_8297,N_1176,N_1269);
and U8298 (N_8298,N_424,N_1997);
nand U8299 (N_8299,N_1602,N_3144);
or U8300 (N_8300,N_2585,N_4616);
or U8301 (N_8301,N_3209,N_1521);
nand U8302 (N_8302,N_4055,N_3925);
nand U8303 (N_8303,N_2743,N_3881);
or U8304 (N_8304,N_1103,N_291);
nand U8305 (N_8305,N_2015,N_3166);
or U8306 (N_8306,N_4416,N_3562);
or U8307 (N_8307,N_2015,N_4654);
nand U8308 (N_8308,N_3927,N_2215);
and U8309 (N_8309,N_766,N_470);
nor U8310 (N_8310,N_3300,N_2569);
or U8311 (N_8311,N_2919,N_2428);
nor U8312 (N_8312,N_2900,N_485);
and U8313 (N_8313,N_1562,N_2262);
or U8314 (N_8314,N_1844,N_3762);
nand U8315 (N_8315,N_2913,N_3506);
or U8316 (N_8316,N_4681,N_2635);
xor U8317 (N_8317,N_2972,N_1564);
nor U8318 (N_8318,N_2806,N_4940);
or U8319 (N_8319,N_1106,N_4094);
nand U8320 (N_8320,N_3221,N_2043);
nor U8321 (N_8321,N_4028,N_1639);
and U8322 (N_8322,N_2085,N_4048);
or U8323 (N_8323,N_3548,N_1677);
and U8324 (N_8324,N_2727,N_78);
and U8325 (N_8325,N_25,N_4118);
and U8326 (N_8326,N_1269,N_2790);
nor U8327 (N_8327,N_2666,N_4618);
nand U8328 (N_8328,N_545,N_2744);
and U8329 (N_8329,N_625,N_3800);
nand U8330 (N_8330,N_4205,N_1782);
nor U8331 (N_8331,N_4154,N_205);
xor U8332 (N_8332,N_4398,N_4827);
and U8333 (N_8333,N_3255,N_1107);
and U8334 (N_8334,N_4814,N_3607);
nor U8335 (N_8335,N_2622,N_1494);
nor U8336 (N_8336,N_3522,N_1439);
or U8337 (N_8337,N_4750,N_3074);
nor U8338 (N_8338,N_2884,N_1788);
nand U8339 (N_8339,N_4657,N_3059);
xor U8340 (N_8340,N_1049,N_1526);
or U8341 (N_8341,N_2862,N_3245);
and U8342 (N_8342,N_4133,N_2796);
nand U8343 (N_8343,N_1136,N_3319);
xnor U8344 (N_8344,N_2415,N_494);
and U8345 (N_8345,N_1536,N_4812);
and U8346 (N_8346,N_191,N_253);
nor U8347 (N_8347,N_1204,N_192);
and U8348 (N_8348,N_2063,N_2575);
and U8349 (N_8349,N_122,N_833);
nand U8350 (N_8350,N_691,N_1062);
nand U8351 (N_8351,N_2249,N_1803);
nor U8352 (N_8352,N_2312,N_2152);
nor U8353 (N_8353,N_3800,N_399);
nand U8354 (N_8354,N_2748,N_624);
nor U8355 (N_8355,N_784,N_3280);
or U8356 (N_8356,N_374,N_1938);
nand U8357 (N_8357,N_4032,N_1904);
and U8358 (N_8358,N_430,N_4532);
or U8359 (N_8359,N_2688,N_2372);
or U8360 (N_8360,N_2852,N_3539);
nor U8361 (N_8361,N_938,N_4061);
or U8362 (N_8362,N_4075,N_1731);
nand U8363 (N_8363,N_2067,N_2608);
and U8364 (N_8364,N_4700,N_586);
and U8365 (N_8365,N_1804,N_876);
xnor U8366 (N_8366,N_190,N_3804);
or U8367 (N_8367,N_2057,N_1708);
xor U8368 (N_8368,N_1778,N_1981);
or U8369 (N_8369,N_2125,N_1793);
nor U8370 (N_8370,N_1934,N_723);
or U8371 (N_8371,N_2540,N_778);
nor U8372 (N_8372,N_2420,N_1213);
nand U8373 (N_8373,N_2310,N_3825);
nand U8374 (N_8374,N_1524,N_2754);
nor U8375 (N_8375,N_3077,N_1249);
nand U8376 (N_8376,N_4219,N_4013);
nand U8377 (N_8377,N_2637,N_2085);
and U8378 (N_8378,N_733,N_2789);
or U8379 (N_8379,N_4793,N_3014);
nand U8380 (N_8380,N_1512,N_2658);
xor U8381 (N_8381,N_1315,N_3424);
xnor U8382 (N_8382,N_761,N_2539);
nor U8383 (N_8383,N_2344,N_2779);
nand U8384 (N_8384,N_3779,N_4363);
or U8385 (N_8385,N_1202,N_1949);
nand U8386 (N_8386,N_182,N_3572);
or U8387 (N_8387,N_1501,N_20);
nand U8388 (N_8388,N_1417,N_691);
or U8389 (N_8389,N_3181,N_2918);
or U8390 (N_8390,N_2339,N_1412);
xnor U8391 (N_8391,N_3368,N_1825);
or U8392 (N_8392,N_2753,N_3847);
nand U8393 (N_8393,N_3580,N_2069);
or U8394 (N_8394,N_2934,N_2278);
nor U8395 (N_8395,N_4258,N_1891);
nor U8396 (N_8396,N_1172,N_4152);
nand U8397 (N_8397,N_1571,N_2512);
nand U8398 (N_8398,N_299,N_559);
and U8399 (N_8399,N_931,N_2411);
nand U8400 (N_8400,N_3922,N_4403);
nor U8401 (N_8401,N_3561,N_3691);
and U8402 (N_8402,N_3778,N_2747);
nand U8403 (N_8403,N_151,N_4014);
nand U8404 (N_8404,N_1797,N_3684);
nand U8405 (N_8405,N_1973,N_1868);
or U8406 (N_8406,N_4273,N_2231);
nor U8407 (N_8407,N_464,N_4072);
nand U8408 (N_8408,N_3198,N_2248);
nor U8409 (N_8409,N_3624,N_3087);
nand U8410 (N_8410,N_594,N_2846);
nand U8411 (N_8411,N_1174,N_3686);
nor U8412 (N_8412,N_256,N_725);
and U8413 (N_8413,N_357,N_1762);
or U8414 (N_8414,N_2622,N_2091);
and U8415 (N_8415,N_3415,N_1292);
and U8416 (N_8416,N_3839,N_4370);
or U8417 (N_8417,N_1866,N_2584);
and U8418 (N_8418,N_1037,N_4613);
nand U8419 (N_8419,N_3106,N_2498);
and U8420 (N_8420,N_2460,N_3343);
or U8421 (N_8421,N_67,N_4759);
or U8422 (N_8422,N_2651,N_3342);
and U8423 (N_8423,N_1958,N_3364);
nor U8424 (N_8424,N_1581,N_2966);
or U8425 (N_8425,N_4286,N_3005);
nor U8426 (N_8426,N_1734,N_3692);
and U8427 (N_8427,N_1260,N_1121);
and U8428 (N_8428,N_3531,N_4040);
and U8429 (N_8429,N_3129,N_1438);
nand U8430 (N_8430,N_1436,N_3828);
and U8431 (N_8431,N_3766,N_991);
nor U8432 (N_8432,N_290,N_945);
xor U8433 (N_8433,N_4476,N_300);
or U8434 (N_8434,N_4232,N_3177);
or U8435 (N_8435,N_3419,N_2259);
or U8436 (N_8436,N_2008,N_3834);
nand U8437 (N_8437,N_1955,N_3844);
and U8438 (N_8438,N_3102,N_1526);
nor U8439 (N_8439,N_1906,N_3321);
xor U8440 (N_8440,N_4548,N_3483);
or U8441 (N_8441,N_2348,N_1384);
nand U8442 (N_8442,N_4478,N_3103);
nand U8443 (N_8443,N_3768,N_4772);
or U8444 (N_8444,N_856,N_2799);
xnor U8445 (N_8445,N_4002,N_839);
or U8446 (N_8446,N_1523,N_1464);
or U8447 (N_8447,N_3826,N_4982);
or U8448 (N_8448,N_622,N_117);
nand U8449 (N_8449,N_4464,N_1370);
nand U8450 (N_8450,N_4985,N_3029);
and U8451 (N_8451,N_2357,N_594);
and U8452 (N_8452,N_4382,N_3063);
and U8453 (N_8453,N_3397,N_241);
nor U8454 (N_8454,N_4116,N_4090);
or U8455 (N_8455,N_99,N_3825);
nand U8456 (N_8456,N_2115,N_3072);
and U8457 (N_8457,N_122,N_1588);
and U8458 (N_8458,N_2890,N_4953);
and U8459 (N_8459,N_929,N_2116);
nand U8460 (N_8460,N_2004,N_1441);
nor U8461 (N_8461,N_4775,N_4209);
nand U8462 (N_8462,N_4833,N_3158);
nand U8463 (N_8463,N_4722,N_4555);
nor U8464 (N_8464,N_2886,N_3264);
or U8465 (N_8465,N_1125,N_2302);
nand U8466 (N_8466,N_953,N_227);
nand U8467 (N_8467,N_1520,N_3173);
and U8468 (N_8468,N_2580,N_4487);
xor U8469 (N_8469,N_3571,N_3862);
and U8470 (N_8470,N_3262,N_4862);
nor U8471 (N_8471,N_772,N_2397);
nor U8472 (N_8472,N_3919,N_473);
or U8473 (N_8473,N_1242,N_1449);
xor U8474 (N_8474,N_2441,N_3480);
nand U8475 (N_8475,N_227,N_3119);
and U8476 (N_8476,N_4143,N_79);
nand U8477 (N_8477,N_1951,N_2280);
or U8478 (N_8478,N_3741,N_3799);
and U8479 (N_8479,N_3700,N_3040);
and U8480 (N_8480,N_2317,N_275);
or U8481 (N_8481,N_3113,N_1758);
or U8482 (N_8482,N_3716,N_3954);
or U8483 (N_8483,N_3169,N_4329);
xnor U8484 (N_8484,N_3403,N_324);
nor U8485 (N_8485,N_3960,N_434);
nand U8486 (N_8486,N_440,N_2601);
and U8487 (N_8487,N_2713,N_203);
or U8488 (N_8488,N_3756,N_649);
or U8489 (N_8489,N_362,N_2353);
xnor U8490 (N_8490,N_959,N_4074);
and U8491 (N_8491,N_4711,N_4802);
and U8492 (N_8492,N_4290,N_1847);
and U8493 (N_8493,N_4646,N_4973);
and U8494 (N_8494,N_1362,N_3303);
and U8495 (N_8495,N_3315,N_1831);
and U8496 (N_8496,N_3198,N_2728);
and U8497 (N_8497,N_1481,N_4777);
and U8498 (N_8498,N_3935,N_1712);
nand U8499 (N_8499,N_2447,N_1655);
and U8500 (N_8500,N_2943,N_3743);
nor U8501 (N_8501,N_777,N_2077);
or U8502 (N_8502,N_1505,N_4737);
xor U8503 (N_8503,N_4327,N_3141);
nor U8504 (N_8504,N_4483,N_2116);
nand U8505 (N_8505,N_1143,N_2990);
nand U8506 (N_8506,N_3688,N_4624);
or U8507 (N_8507,N_2362,N_1024);
and U8508 (N_8508,N_887,N_685);
nand U8509 (N_8509,N_4217,N_1384);
and U8510 (N_8510,N_2345,N_1238);
nand U8511 (N_8511,N_1305,N_2812);
or U8512 (N_8512,N_2484,N_298);
nor U8513 (N_8513,N_308,N_1565);
nor U8514 (N_8514,N_642,N_12);
xnor U8515 (N_8515,N_1266,N_894);
nor U8516 (N_8516,N_4916,N_4640);
or U8517 (N_8517,N_3664,N_4772);
or U8518 (N_8518,N_1612,N_4958);
or U8519 (N_8519,N_1900,N_578);
or U8520 (N_8520,N_804,N_2601);
nand U8521 (N_8521,N_4773,N_4271);
nor U8522 (N_8522,N_1552,N_1744);
nand U8523 (N_8523,N_542,N_194);
or U8524 (N_8524,N_2325,N_1264);
nor U8525 (N_8525,N_2506,N_1300);
nor U8526 (N_8526,N_4368,N_3815);
nand U8527 (N_8527,N_2487,N_3327);
or U8528 (N_8528,N_3216,N_3300);
nand U8529 (N_8529,N_2683,N_648);
nor U8530 (N_8530,N_3826,N_3208);
or U8531 (N_8531,N_2353,N_2247);
nand U8532 (N_8532,N_2044,N_1215);
and U8533 (N_8533,N_2914,N_414);
xnor U8534 (N_8534,N_1024,N_397);
nor U8535 (N_8535,N_3011,N_2461);
nand U8536 (N_8536,N_2842,N_46);
and U8537 (N_8537,N_920,N_2324);
nor U8538 (N_8538,N_3841,N_4040);
or U8539 (N_8539,N_716,N_84);
nor U8540 (N_8540,N_3307,N_574);
nor U8541 (N_8541,N_2548,N_4506);
or U8542 (N_8542,N_1176,N_2756);
or U8543 (N_8543,N_2083,N_4791);
nand U8544 (N_8544,N_4982,N_4903);
or U8545 (N_8545,N_2054,N_3143);
and U8546 (N_8546,N_3300,N_2119);
or U8547 (N_8547,N_202,N_2924);
xnor U8548 (N_8548,N_4603,N_3592);
and U8549 (N_8549,N_3883,N_3674);
or U8550 (N_8550,N_37,N_2412);
or U8551 (N_8551,N_641,N_1490);
or U8552 (N_8552,N_334,N_2232);
or U8553 (N_8553,N_728,N_884);
or U8554 (N_8554,N_3679,N_4319);
or U8555 (N_8555,N_2729,N_87);
nand U8556 (N_8556,N_1044,N_345);
or U8557 (N_8557,N_2167,N_1342);
and U8558 (N_8558,N_2192,N_3090);
nor U8559 (N_8559,N_88,N_3093);
or U8560 (N_8560,N_1271,N_2816);
nand U8561 (N_8561,N_1414,N_695);
nor U8562 (N_8562,N_37,N_1070);
and U8563 (N_8563,N_4635,N_2775);
nand U8564 (N_8564,N_3321,N_3710);
nor U8565 (N_8565,N_1307,N_1990);
nor U8566 (N_8566,N_2702,N_3085);
nor U8567 (N_8567,N_129,N_3486);
or U8568 (N_8568,N_18,N_4082);
nor U8569 (N_8569,N_1376,N_773);
nor U8570 (N_8570,N_3704,N_2589);
xnor U8571 (N_8571,N_3748,N_2115);
or U8572 (N_8572,N_884,N_2738);
nand U8573 (N_8573,N_233,N_4506);
and U8574 (N_8574,N_2959,N_4248);
or U8575 (N_8575,N_2755,N_3257);
nand U8576 (N_8576,N_4750,N_3529);
nand U8577 (N_8577,N_3501,N_162);
nand U8578 (N_8578,N_3059,N_1436);
xor U8579 (N_8579,N_4684,N_2731);
nor U8580 (N_8580,N_3107,N_2758);
nor U8581 (N_8581,N_1438,N_442);
nor U8582 (N_8582,N_2127,N_3987);
and U8583 (N_8583,N_543,N_412);
and U8584 (N_8584,N_2573,N_3984);
nor U8585 (N_8585,N_4331,N_2657);
or U8586 (N_8586,N_2311,N_4423);
nor U8587 (N_8587,N_3012,N_3915);
nand U8588 (N_8588,N_3150,N_4670);
nand U8589 (N_8589,N_1499,N_1346);
or U8590 (N_8590,N_3859,N_46);
nor U8591 (N_8591,N_2963,N_4291);
and U8592 (N_8592,N_4147,N_348);
and U8593 (N_8593,N_4859,N_2174);
and U8594 (N_8594,N_3226,N_3006);
nand U8595 (N_8595,N_4633,N_2354);
nand U8596 (N_8596,N_679,N_1673);
nor U8597 (N_8597,N_3353,N_2557);
and U8598 (N_8598,N_4350,N_3086);
nand U8599 (N_8599,N_4419,N_2015);
nand U8600 (N_8600,N_2721,N_270);
and U8601 (N_8601,N_2314,N_4063);
nand U8602 (N_8602,N_3518,N_3049);
nor U8603 (N_8603,N_2003,N_3915);
nand U8604 (N_8604,N_1030,N_1512);
or U8605 (N_8605,N_2383,N_2903);
and U8606 (N_8606,N_1857,N_2329);
nand U8607 (N_8607,N_3953,N_1758);
or U8608 (N_8608,N_3024,N_3959);
nor U8609 (N_8609,N_2122,N_1835);
nor U8610 (N_8610,N_3648,N_2587);
nor U8611 (N_8611,N_4193,N_88);
xor U8612 (N_8612,N_1140,N_4079);
or U8613 (N_8613,N_4235,N_4285);
nand U8614 (N_8614,N_3052,N_2757);
nand U8615 (N_8615,N_1510,N_4098);
nor U8616 (N_8616,N_4906,N_4004);
nand U8617 (N_8617,N_1717,N_1913);
nand U8618 (N_8618,N_4771,N_1532);
nand U8619 (N_8619,N_4146,N_952);
nor U8620 (N_8620,N_4379,N_2883);
xor U8621 (N_8621,N_2340,N_3086);
nor U8622 (N_8622,N_2902,N_464);
nor U8623 (N_8623,N_830,N_2736);
or U8624 (N_8624,N_1817,N_53);
nor U8625 (N_8625,N_2,N_3463);
or U8626 (N_8626,N_1366,N_3266);
nor U8627 (N_8627,N_1487,N_4620);
and U8628 (N_8628,N_1540,N_2536);
nor U8629 (N_8629,N_138,N_3671);
and U8630 (N_8630,N_3888,N_2235);
nand U8631 (N_8631,N_2471,N_2165);
nor U8632 (N_8632,N_433,N_2121);
or U8633 (N_8633,N_621,N_4342);
nor U8634 (N_8634,N_1184,N_681);
or U8635 (N_8635,N_2106,N_4846);
nand U8636 (N_8636,N_2034,N_2707);
nand U8637 (N_8637,N_4874,N_580);
nand U8638 (N_8638,N_1867,N_3686);
or U8639 (N_8639,N_4898,N_4319);
nor U8640 (N_8640,N_4699,N_2034);
and U8641 (N_8641,N_1106,N_2614);
or U8642 (N_8642,N_1520,N_1509);
and U8643 (N_8643,N_4359,N_3317);
or U8644 (N_8644,N_3725,N_999);
and U8645 (N_8645,N_2482,N_2514);
nand U8646 (N_8646,N_1715,N_1740);
xnor U8647 (N_8647,N_4726,N_4079);
or U8648 (N_8648,N_675,N_4598);
and U8649 (N_8649,N_3219,N_3169);
nor U8650 (N_8650,N_2462,N_3276);
nor U8651 (N_8651,N_154,N_1122);
or U8652 (N_8652,N_3662,N_289);
or U8653 (N_8653,N_987,N_563);
or U8654 (N_8654,N_878,N_4451);
and U8655 (N_8655,N_4809,N_1715);
nor U8656 (N_8656,N_2068,N_94);
nor U8657 (N_8657,N_4419,N_1239);
nand U8658 (N_8658,N_3628,N_2932);
nor U8659 (N_8659,N_2573,N_4046);
nor U8660 (N_8660,N_2461,N_4622);
nand U8661 (N_8661,N_3179,N_336);
or U8662 (N_8662,N_4029,N_1739);
nand U8663 (N_8663,N_538,N_789);
or U8664 (N_8664,N_198,N_3458);
nor U8665 (N_8665,N_2674,N_1645);
or U8666 (N_8666,N_4638,N_2189);
and U8667 (N_8667,N_2159,N_3273);
nor U8668 (N_8668,N_3787,N_213);
or U8669 (N_8669,N_1594,N_1954);
and U8670 (N_8670,N_3558,N_4039);
nand U8671 (N_8671,N_2062,N_2449);
and U8672 (N_8672,N_446,N_1691);
nor U8673 (N_8673,N_1896,N_4275);
and U8674 (N_8674,N_4176,N_447);
or U8675 (N_8675,N_4651,N_4536);
or U8676 (N_8676,N_2161,N_1394);
or U8677 (N_8677,N_1137,N_1723);
and U8678 (N_8678,N_3702,N_1942);
nor U8679 (N_8679,N_1147,N_4197);
nor U8680 (N_8680,N_133,N_2978);
xnor U8681 (N_8681,N_3467,N_2850);
nor U8682 (N_8682,N_3136,N_1588);
and U8683 (N_8683,N_3370,N_4220);
and U8684 (N_8684,N_801,N_942);
and U8685 (N_8685,N_4884,N_695);
and U8686 (N_8686,N_1896,N_3947);
nor U8687 (N_8687,N_4409,N_4907);
nand U8688 (N_8688,N_4964,N_1985);
nor U8689 (N_8689,N_3327,N_3388);
nor U8690 (N_8690,N_3856,N_3719);
or U8691 (N_8691,N_3273,N_2173);
nand U8692 (N_8692,N_2103,N_129);
and U8693 (N_8693,N_1566,N_948);
or U8694 (N_8694,N_4672,N_1573);
xor U8695 (N_8695,N_2947,N_1550);
and U8696 (N_8696,N_2340,N_3637);
and U8697 (N_8697,N_206,N_1559);
xnor U8698 (N_8698,N_3151,N_1615);
nor U8699 (N_8699,N_686,N_542);
nand U8700 (N_8700,N_1148,N_978);
and U8701 (N_8701,N_4204,N_4732);
or U8702 (N_8702,N_3093,N_1139);
nand U8703 (N_8703,N_2374,N_4341);
nand U8704 (N_8704,N_3259,N_3181);
nor U8705 (N_8705,N_961,N_2986);
nor U8706 (N_8706,N_1510,N_268);
or U8707 (N_8707,N_2873,N_4635);
nand U8708 (N_8708,N_3332,N_4903);
xor U8709 (N_8709,N_2844,N_3561);
nor U8710 (N_8710,N_3288,N_389);
nor U8711 (N_8711,N_2153,N_4418);
nor U8712 (N_8712,N_1511,N_1853);
nor U8713 (N_8713,N_2391,N_3051);
nor U8714 (N_8714,N_2067,N_77);
and U8715 (N_8715,N_2797,N_1635);
or U8716 (N_8716,N_347,N_4387);
nand U8717 (N_8717,N_4591,N_1227);
or U8718 (N_8718,N_506,N_1921);
and U8719 (N_8719,N_2202,N_1079);
xor U8720 (N_8720,N_276,N_2055);
nor U8721 (N_8721,N_4688,N_1140);
nor U8722 (N_8722,N_4724,N_4089);
and U8723 (N_8723,N_634,N_1785);
and U8724 (N_8724,N_2921,N_4336);
nor U8725 (N_8725,N_4872,N_2855);
or U8726 (N_8726,N_3540,N_4696);
nor U8727 (N_8727,N_3221,N_4411);
or U8728 (N_8728,N_2424,N_3375);
and U8729 (N_8729,N_3260,N_176);
or U8730 (N_8730,N_733,N_2699);
nand U8731 (N_8731,N_510,N_2432);
nand U8732 (N_8732,N_3509,N_2747);
or U8733 (N_8733,N_4282,N_3409);
and U8734 (N_8734,N_837,N_2627);
xor U8735 (N_8735,N_3077,N_2141);
and U8736 (N_8736,N_3295,N_405);
and U8737 (N_8737,N_4404,N_3083);
or U8738 (N_8738,N_488,N_4849);
and U8739 (N_8739,N_1617,N_2932);
or U8740 (N_8740,N_2913,N_1374);
nand U8741 (N_8741,N_3401,N_1621);
nor U8742 (N_8742,N_9,N_60);
nor U8743 (N_8743,N_4241,N_4868);
nand U8744 (N_8744,N_4648,N_3622);
nand U8745 (N_8745,N_2215,N_362);
nand U8746 (N_8746,N_954,N_965);
nor U8747 (N_8747,N_1858,N_1549);
nor U8748 (N_8748,N_360,N_2521);
or U8749 (N_8749,N_3086,N_1359);
nand U8750 (N_8750,N_397,N_4408);
xor U8751 (N_8751,N_4164,N_4201);
or U8752 (N_8752,N_984,N_1900);
and U8753 (N_8753,N_3970,N_1982);
nand U8754 (N_8754,N_537,N_2655);
and U8755 (N_8755,N_282,N_3315);
nor U8756 (N_8756,N_3955,N_1262);
and U8757 (N_8757,N_650,N_3635);
or U8758 (N_8758,N_4618,N_4488);
nand U8759 (N_8759,N_2430,N_3900);
or U8760 (N_8760,N_2264,N_558);
and U8761 (N_8761,N_1091,N_478);
nor U8762 (N_8762,N_4939,N_3855);
nand U8763 (N_8763,N_501,N_1079);
nor U8764 (N_8764,N_1097,N_4043);
or U8765 (N_8765,N_187,N_4123);
nor U8766 (N_8766,N_2331,N_4527);
xnor U8767 (N_8767,N_4369,N_533);
nand U8768 (N_8768,N_2811,N_2688);
and U8769 (N_8769,N_4033,N_108);
nand U8770 (N_8770,N_4855,N_4849);
or U8771 (N_8771,N_3284,N_3037);
nor U8772 (N_8772,N_339,N_4830);
or U8773 (N_8773,N_1,N_2241);
and U8774 (N_8774,N_2164,N_330);
nor U8775 (N_8775,N_2234,N_1493);
nand U8776 (N_8776,N_2340,N_4858);
or U8777 (N_8777,N_1144,N_40);
nor U8778 (N_8778,N_3338,N_1376);
nand U8779 (N_8779,N_1879,N_1615);
xnor U8780 (N_8780,N_1340,N_3131);
nand U8781 (N_8781,N_2952,N_2582);
and U8782 (N_8782,N_725,N_1300);
xnor U8783 (N_8783,N_984,N_521);
and U8784 (N_8784,N_987,N_2456);
nor U8785 (N_8785,N_2862,N_4875);
or U8786 (N_8786,N_2825,N_2161);
xor U8787 (N_8787,N_1810,N_4376);
nand U8788 (N_8788,N_1973,N_3513);
xor U8789 (N_8789,N_269,N_1225);
and U8790 (N_8790,N_1195,N_4882);
nand U8791 (N_8791,N_278,N_4893);
nand U8792 (N_8792,N_3227,N_2275);
and U8793 (N_8793,N_922,N_1164);
and U8794 (N_8794,N_4845,N_2498);
and U8795 (N_8795,N_996,N_4364);
and U8796 (N_8796,N_92,N_2520);
xor U8797 (N_8797,N_2760,N_1819);
nor U8798 (N_8798,N_4078,N_2345);
and U8799 (N_8799,N_4329,N_2094);
nand U8800 (N_8800,N_3320,N_1752);
or U8801 (N_8801,N_2325,N_2527);
xor U8802 (N_8802,N_1785,N_26);
nor U8803 (N_8803,N_3239,N_4093);
nor U8804 (N_8804,N_2575,N_4320);
and U8805 (N_8805,N_4657,N_684);
nor U8806 (N_8806,N_227,N_1744);
or U8807 (N_8807,N_2887,N_722);
and U8808 (N_8808,N_1304,N_4209);
and U8809 (N_8809,N_2736,N_3237);
nor U8810 (N_8810,N_2249,N_2163);
or U8811 (N_8811,N_3128,N_3030);
nand U8812 (N_8812,N_3198,N_1474);
nor U8813 (N_8813,N_4872,N_1631);
xor U8814 (N_8814,N_1912,N_1166);
nand U8815 (N_8815,N_4294,N_3262);
xnor U8816 (N_8816,N_1894,N_1431);
and U8817 (N_8817,N_3928,N_4839);
or U8818 (N_8818,N_4086,N_1105);
or U8819 (N_8819,N_4550,N_3798);
xor U8820 (N_8820,N_3465,N_4176);
and U8821 (N_8821,N_2074,N_1632);
nand U8822 (N_8822,N_2223,N_4528);
nand U8823 (N_8823,N_4465,N_4381);
nor U8824 (N_8824,N_1827,N_2336);
nand U8825 (N_8825,N_4203,N_174);
or U8826 (N_8826,N_767,N_3857);
nor U8827 (N_8827,N_4710,N_806);
xnor U8828 (N_8828,N_3392,N_2953);
or U8829 (N_8829,N_1313,N_1338);
xor U8830 (N_8830,N_4361,N_2735);
nor U8831 (N_8831,N_3592,N_2069);
nand U8832 (N_8832,N_3115,N_513);
and U8833 (N_8833,N_2304,N_1293);
nor U8834 (N_8834,N_2948,N_3221);
nor U8835 (N_8835,N_3796,N_1225);
or U8836 (N_8836,N_2932,N_4110);
or U8837 (N_8837,N_2865,N_4506);
and U8838 (N_8838,N_1417,N_3548);
nor U8839 (N_8839,N_4102,N_252);
or U8840 (N_8840,N_3727,N_736);
or U8841 (N_8841,N_3285,N_4732);
and U8842 (N_8842,N_3704,N_4266);
nand U8843 (N_8843,N_3262,N_1180);
nor U8844 (N_8844,N_404,N_270);
or U8845 (N_8845,N_2037,N_3787);
nor U8846 (N_8846,N_2703,N_1315);
nor U8847 (N_8847,N_2460,N_2578);
or U8848 (N_8848,N_585,N_784);
nor U8849 (N_8849,N_4938,N_4394);
nand U8850 (N_8850,N_2811,N_1354);
nand U8851 (N_8851,N_3586,N_4384);
and U8852 (N_8852,N_942,N_2159);
and U8853 (N_8853,N_749,N_1417);
or U8854 (N_8854,N_519,N_1825);
nor U8855 (N_8855,N_4605,N_4867);
nand U8856 (N_8856,N_1217,N_984);
nor U8857 (N_8857,N_2510,N_2934);
nor U8858 (N_8858,N_86,N_911);
nor U8859 (N_8859,N_2660,N_3067);
or U8860 (N_8860,N_627,N_525);
or U8861 (N_8861,N_273,N_3478);
nand U8862 (N_8862,N_492,N_4522);
nor U8863 (N_8863,N_3864,N_4673);
or U8864 (N_8864,N_4179,N_3009);
nand U8865 (N_8865,N_1516,N_884);
and U8866 (N_8866,N_1043,N_1873);
and U8867 (N_8867,N_4628,N_2982);
nor U8868 (N_8868,N_3670,N_2335);
nor U8869 (N_8869,N_508,N_2017);
nand U8870 (N_8870,N_4244,N_488);
nand U8871 (N_8871,N_4127,N_1730);
nor U8872 (N_8872,N_4837,N_4509);
or U8873 (N_8873,N_255,N_4541);
and U8874 (N_8874,N_3966,N_4983);
nand U8875 (N_8875,N_1289,N_2219);
nand U8876 (N_8876,N_3911,N_2012);
nor U8877 (N_8877,N_4702,N_420);
and U8878 (N_8878,N_1544,N_1883);
nor U8879 (N_8879,N_4222,N_2604);
and U8880 (N_8880,N_1523,N_2663);
nand U8881 (N_8881,N_2829,N_2885);
or U8882 (N_8882,N_225,N_960);
xnor U8883 (N_8883,N_4950,N_3241);
nor U8884 (N_8884,N_1300,N_1625);
nor U8885 (N_8885,N_961,N_3152);
or U8886 (N_8886,N_3831,N_3931);
nand U8887 (N_8887,N_2407,N_2308);
or U8888 (N_8888,N_2195,N_2001);
and U8889 (N_8889,N_3853,N_3770);
nor U8890 (N_8890,N_3990,N_4785);
or U8891 (N_8891,N_3899,N_2917);
and U8892 (N_8892,N_491,N_1212);
nand U8893 (N_8893,N_1118,N_3810);
xnor U8894 (N_8894,N_4846,N_1674);
nor U8895 (N_8895,N_4946,N_1152);
nor U8896 (N_8896,N_935,N_1888);
or U8897 (N_8897,N_4846,N_1996);
nor U8898 (N_8898,N_921,N_2790);
nand U8899 (N_8899,N_3552,N_2749);
and U8900 (N_8900,N_1645,N_1775);
or U8901 (N_8901,N_1026,N_4460);
nor U8902 (N_8902,N_1449,N_2418);
or U8903 (N_8903,N_3285,N_3983);
nor U8904 (N_8904,N_2352,N_802);
and U8905 (N_8905,N_4565,N_1318);
or U8906 (N_8906,N_568,N_370);
and U8907 (N_8907,N_4728,N_51);
nand U8908 (N_8908,N_4939,N_360);
and U8909 (N_8909,N_1060,N_4755);
and U8910 (N_8910,N_684,N_527);
or U8911 (N_8911,N_1181,N_764);
nor U8912 (N_8912,N_2309,N_4830);
and U8913 (N_8913,N_2226,N_597);
nand U8914 (N_8914,N_4771,N_1997);
or U8915 (N_8915,N_4337,N_4964);
nand U8916 (N_8916,N_4760,N_2799);
xor U8917 (N_8917,N_2642,N_4033);
and U8918 (N_8918,N_3890,N_2856);
or U8919 (N_8919,N_3646,N_2860);
and U8920 (N_8920,N_1897,N_3831);
nor U8921 (N_8921,N_107,N_842);
or U8922 (N_8922,N_2684,N_294);
and U8923 (N_8923,N_319,N_3712);
nand U8924 (N_8924,N_4527,N_4197);
nand U8925 (N_8925,N_4978,N_201);
xor U8926 (N_8926,N_1542,N_585);
xor U8927 (N_8927,N_2462,N_2097);
nand U8928 (N_8928,N_105,N_1562);
nand U8929 (N_8929,N_4285,N_4839);
nor U8930 (N_8930,N_2636,N_2080);
nor U8931 (N_8931,N_1976,N_3415);
and U8932 (N_8932,N_1994,N_1322);
and U8933 (N_8933,N_3140,N_2579);
or U8934 (N_8934,N_4523,N_4988);
nand U8935 (N_8935,N_1967,N_2744);
or U8936 (N_8936,N_574,N_3420);
or U8937 (N_8937,N_2799,N_2355);
or U8938 (N_8938,N_2753,N_1332);
and U8939 (N_8939,N_3393,N_3136);
nand U8940 (N_8940,N_2538,N_3597);
or U8941 (N_8941,N_4096,N_502);
or U8942 (N_8942,N_800,N_1146);
nand U8943 (N_8943,N_3461,N_719);
and U8944 (N_8944,N_770,N_3499);
or U8945 (N_8945,N_117,N_1510);
xor U8946 (N_8946,N_3266,N_308);
nor U8947 (N_8947,N_1663,N_2411);
xnor U8948 (N_8948,N_2955,N_4925);
or U8949 (N_8949,N_698,N_1919);
and U8950 (N_8950,N_4392,N_2951);
nand U8951 (N_8951,N_4017,N_807);
and U8952 (N_8952,N_1943,N_4348);
and U8953 (N_8953,N_4341,N_2799);
nor U8954 (N_8954,N_4952,N_849);
and U8955 (N_8955,N_3269,N_2062);
nor U8956 (N_8956,N_3485,N_414);
nand U8957 (N_8957,N_1802,N_4353);
and U8958 (N_8958,N_4077,N_4964);
and U8959 (N_8959,N_4720,N_1246);
or U8960 (N_8960,N_2442,N_3109);
nor U8961 (N_8961,N_2572,N_1543);
nor U8962 (N_8962,N_3247,N_2820);
xor U8963 (N_8963,N_3614,N_349);
xor U8964 (N_8964,N_108,N_516);
nor U8965 (N_8965,N_3522,N_3342);
nand U8966 (N_8966,N_1129,N_4037);
xnor U8967 (N_8967,N_2476,N_2853);
or U8968 (N_8968,N_2552,N_361);
and U8969 (N_8969,N_2439,N_3015);
or U8970 (N_8970,N_4538,N_142);
nand U8971 (N_8971,N_1301,N_3422);
nand U8972 (N_8972,N_1033,N_3342);
nand U8973 (N_8973,N_1747,N_482);
xnor U8974 (N_8974,N_1560,N_2953);
nor U8975 (N_8975,N_151,N_626);
and U8976 (N_8976,N_3736,N_340);
or U8977 (N_8977,N_3433,N_3817);
nand U8978 (N_8978,N_1497,N_4697);
or U8979 (N_8979,N_814,N_3623);
nor U8980 (N_8980,N_4206,N_1948);
or U8981 (N_8981,N_3314,N_4104);
nand U8982 (N_8982,N_4536,N_3326);
and U8983 (N_8983,N_438,N_3232);
or U8984 (N_8984,N_2507,N_839);
nand U8985 (N_8985,N_3390,N_432);
or U8986 (N_8986,N_1377,N_3724);
or U8987 (N_8987,N_2809,N_4102);
nor U8988 (N_8988,N_4041,N_1431);
xnor U8989 (N_8989,N_1592,N_1702);
and U8990 (N_8990,N_1576,N_2789);
xnor U8991 (N_8991,N_1658,N_1733);
or U8992 (N_8992,N_378,N_4556);
or U8993 (N_8993,N_218,N_266);
and U8994 (N_8994,N_844,N_4336);
nor U8995 (N_8995,N_2802,N_3169);
and U8996 (N_8996,N_3029,N_3921);
nand U8997 (N_8997,N_4003,N_3624);
or U8998 (N_8998,N_4609,N_2362);
nor U8999 (N_8999,N_3943,N_2425);
or U9000 (N_9000,N_2629,N_4805);
and U9001 (N_9001,N_4938,N_2052);
and U9002 (N_9002,N_2421,N_2020);
or U9003 (N_9003,N_3944,N_4392);
nor U9004 (N_9004,N_1608,N_292);
nand U9005 (N_9005,N_3193,N_2644);
nor U9006 (N_9006,N_2329,N_2885);
nand U9007 (N_9007,N_2734,N_2861);
and U9008 (N_9008,N_1892,N_2851);
nand U9009 (N_9009,N_189,N_422);
or U9010 (N_9010,N_295,N_3185);
nor U9011 (N_9011,N_86,N_1521);
or U9012 (N_9012,N_4532,N_3432);
nand U9013 (N_9013,N_1582,N_902);
nand U9014 (N_9014,N_3412,N_3837);
nand U9015 (N_9015,N_3576,N_2076);
xnor U9016 (N_9016,N_1049,N_879);
nor U9017 (N_9017,N_4690,N_4168);
and U9018 (N_9018,N_4886,N_2622);
or U9019 (N_9019,N_4251,N_1928);
and U9020 (N_9020,N_1146,N_2749);
nor U9021 (N_9021,N_4187,N_3245);
and U9022 (N_9022,N_3154,N_1509);
nand U9023 (N_9023,N_4252,N_2389);
and U9024 (N_9024,N_3558,N_2744);
and U9025 (N_9025,N_1511,N_2493);
nand U9026 (N_9026,N_2820,N_3922);
or U9027 (N_9027,N_3102,N_1883);
nand U9028 (N_9028,N_2446,N_4346);
nor U9029 (N_9029,N_1614,N_1510);
xor U9030 (N_9030,N_4908,N_356);
nand U9031 (N_9031,N_4080,N_4258);
and U9032 (N_9032,N_4811,N_958);
xnor U9033 (N_9033,N_3174,N_1482);
nand U9034 (N_9034,N_4799,N_1757);
or U9035 (N_9035,N_4753,N_3233);
and U9036 (N_9036,N_420,N_2157);
and U9037 (N_9037,N_1282,N_3053);
nor U9038 (N_9038,N_249,N_3114);
nor U9039 (N_9039,N_555,N_884);
xor U9040 (N_9040,N_96,N_1202);
and U9041 (N_9041,N_1339,N_978);
nor U9042 (N_9042,N_1035,N_4728);
or U9043 (N_9043,N_4828,N_1377);
and U9044 (N_9044,N_274,N_3704);
and U9045 (N_9045,N_2139,N_2769);
xor U9046 (N_9046,N_2851,N_3999);
or U9047 (N_9047,N_3407,N_4989);
nor U9048 (N_9048,N_4064,N_4037);
nor U9049 (N_9049,N_1052,N_2330);
nand U9050 (N_9050,N_1781,N_1050);
nand U9051 (N_9051,N_1255,N_713);
nor U9052 (N_9052,N_3688,N_1753);
or U9053 (N_9053,N_1738,N_3227);
or U9054 (N_9054,N_567,N_4029);
nand U9055 (N_9055,N_1889,N_2996);
nor U9056 (N_9056,N_1062,N_411);
or U9057 (N_9057,N_1465,N_2105);
xnor U9058 (N_9058,N_3630,N_522);
xnor U9059 (N_9059,N_1273,N_113);
nand U9060 (N_9060,N_4468,N_4773);
nand U9061 (N_9061,N_4649,N_4854);
nand U9062 (N_9062,N_1119,N_150);
or U9063 (N_9063,N_127,N_346);
or U9064 (N_9064,N_1248,N_1344);
and U9065 (N_9065,N_2740,N_1892);
nor U9066 (N_9066,N_4295,N_2197);
nand U9067 (N_9067,N_4693,N_4133);
nand U9068 (N_9068,N_747,N_146);
nor U9069 (N_9069,N_4277,N_3639);
nor U9070 (N_9070,N_592,N_4586);
or U9071 (N_9071,N_2608,N_1526);
xnor U9072 (N_9072,N_65,N_4650);
nor U9073 (N_9073,N_4650,N_4164);
nand U9074 (N_9074,N_4367,N_1405);
nand U9075 (N_9075,N_1840,N_3849);
nand U9076 (N_9076,N_1845,N_271);
nor U9077 (N_9077,N_20,N_688);
or U9078 (N_9078,N_4826,N_2939);
or U9079 (N_9079,N_3885,N_1074);
nor U9080 (N_9080,N_3388,N_2443);
or U9081 (N_9081,N_1719,N_4558);
nor U9082 (N_9082,N_842,N_514);
and U9083 (N_9083,N_4818,N_877);
or U9084 (N_9084,N_4028,N_3881);
or U9085 (N_9085,N_358,N_91);
nor U9086 (N_9086,N_1533,N_1645);
xnor U9087 (N_9087,N_1451,N_425);
nor U9088 (N_9088,N_986,N_3040);
nor U9089 (N_9089,N_3504,N_2706);
nand U9090 (N_9090,N_2137,N_4819);
or U9091 (N_9091,N_125,N_906);
or U9092 (N_9092,N_1593,N_3172);
or U9093 (N_9093,N_2926,N_2947);
nand U9094 (N_9094,N_22,N_3346);
and U9095 (N_9095,N_2957,N_630);
and U9096 (N_9096,N_341,N_2400);
xor U9097 (N_9097,N_4741,N_2556);
nor U9098 (N_9098,N_1083,N_1549);
xnor U9099 (N_9099,N_3458,N_3834);
or U9100 (N_9100,N_1912,N_3128);
or U9101 (N_9101,N_2788,N_4554);
or U9102 (N_9102,N_1643,N_3978);
xor U9103 (N_9103,N_547,N_3424);
nor U9104 (N_9104,N_142,N_1145);
nor U9105 (N_9105,N_2050,N_2798);
or U9106 (N_9106,N_3983,N_3135);
and U9107 (N_9107,N_45,N_2324);
or U9108 (N_9108,N_2523,N_923);
nor U9109 (N_9109,N_4133,N_1750);
and U9110 (N_9110,N_2988,N_3262);
or U9111 (N_9111,N_3716,N_485);
nor U9112 (N_9112,N_2290,N_2765);
and U9113 (N_9113,N_3103,N_2668);
nor U9114 (N_9114,N_4906,N_3066);
nor U9115 (N_9115,N_328,N_1377);
nand U9116 (N_9116,N_3553,N_1093);
nor U9117 (N_9117,N_2203,N_3984);
nor U9118 (N_9118,N_543,N_1365);
or U9119 (N_9119,N_763,N_3508);
nand U9120 (N_9120,N_4638,N_4122);
nand U9121 (N_9121,N_2437,N_373);
and U9122 (N_9122,N_1203,N_3558);
nor U9123 (N_9123,N_519,N_2555);
or U9124 (N_9124,N_549,N_204);
nor U9125 (N_9125,N_3810,N_3933);
nand U9126 (N_9126,N_3573,N_2035);
or U9127 (N_9127,N_1942,N_2262);
nor U9128 (N_9128,N_1131,N_4766);
xor U9129 (N_9129,N_3287,N_3709);
nand U9130 (N_9130,N_3887,N_4568);
and U9131 (N_9131,N_2157,N_2723);
nand U9132 (N_9132,N_900,N_137);
and U9133 (N_9133,N_3891,N_2686);
nor U9134 (N_9134,N_2706,N_2161);
nor U9135 (N_9135,N_4166,N_920);
or U9136 (N_9136,N_457,N_2559);
nor U9137 (N_9137,N_628,N_2496);
nand U9138 (N_9138,N_2033,N_4558);
or U9139 (N_9139,N_4705,N_3885);
xor U9140 (N_9140,N_3560,N_450);
nor U9141 (N_9141,N_3299,N_4336);
or U9142 (N_9142,N_296,N_334);
nor U9143 (N_9143,N_689,N_1962);
and U9144 (N_9144,N_3484,N_383);
and U9145 (N_9145,N_1543,N_4137);
nor U9146 (N_9146,N_3692,N_2489);
xnor U9147 (N_9147,N_1050,N_2486);
and U9148 (N_9148,N_2999,N_4870);
or U9149 (N_9149,N_3583,N_3785);
nor U9150 (N_9150,N_3277,N_654);
and U9151 (N_9151,N_1813,N_2492);
and U9152 (N_9152,N_4454,N_4630);
or U9153 (N_9153,N_297,N_3845);
xor U9154 (N_9154,N_4390,N_107);
nand U9155 (N_9155,N_4870,N_4204);
nor U9156 (N_9156,N_3259,N_1872);
nand U9157 (N_9157,N_1987,N_552);
xor U9158 (N_9158,N_588,N_4649);
nand U9159 (N_9159,N_1344,N_2718);
and U9160 (N_9160,N_2510,N_3903);
or U9161 (N_9161,N_4157,N_4162);
xor U9162 (N_9162,N_2993,N_2634);
and U9163 (N_9163,N_833,N_1209);
nor U9164 (N_9164,N_4110,N_3248);
or U9165 (N_9165,N_3068,N_2441);
and U9166 (N_9166,N_2342,N_587);
nor U9167 (N_9167,N_1881,N_3971);
or U9168 (N_9168,N_2395,N_3388);
or U9169 (N_9169,N_4444,N_1035);
or U9170 (N_9170,N_1337,N_3415);
nor U9171 (N_9171,N_1269,N_966);
and U9172 (N_9172,N_3395,N_1975);
and U9173 (N_9173,N_1354,N_4606);
nand U9174 (N_9174,N_379,N_3341);
nand U9175 (N_9175,N_2099,N_7);
and U9176 (N_9176,N_820,N_3014);
and U9177 (N_9177,N_4821,N_165);
nor U9178 (N_9178,N_1027,N_1704);
nor U9179 (N_9179,N_1429,N_1995);
or U9180 (N_9180,N_2889,N_3699);
xor U9181 (N_9181,N_3058,N_3577);
xor U9182 (N_9182,N_632,N_1302);
or U9183 (N_9183,N_2224,N_1962);
nor U9184 (N_9184,N_3126,N_382);
nand U9185 (N_9185,N_277,N_883);
or U9186 (N_9186,N_4891,N_757);
and U9187 (N_9187,N_1394,N_4748);
and U9188 (N_9188,N_1019,N_192);
or U9189 (N_9189,N_4171,N_4356);
and U9190 (N_9190,N_263,N_2627);
xor U9191 (N_9191,N_652,N_3118);
or U9192 (N_9192,N_404,N_4683);
nor U9193 (N_9193,N_378,N_3127);
nand U9194 (N_9194,N_2601,N_3237);
nor U9195 (N_9195,N_1306,N_2766);
or U9196 (N_9196,N_679,N_1030);
or U9197 (N_9197,N_2749,N_2989);
nand U9198 (N_9198,N_4351,N_4601);
and U9199 (N_9199,N_282,N_4792);
nand U9200 (N_9200,N_495,N_2307);
or U9201 (N_9201,N_2481,N_3942);
nand U9202 (N_9202,N_2692,N_2096);
nand U9203 (N_9203,N_2910,N_345);
nor U9204 (N_9204,N_3827,N_3499);
or U9205 (N_9205,N_1196,N_4906);
nand U9206 (N_9206,N_1055,N_4812);
or U9207 (N_9207,N_3960,N_4217);
xor U9208 (N_9208,N_4900,N_1186);
and U9209 (N_9209,N_3074,N_2940);
nor U9210 (N_9210,N_862,N_1395);
nand U9211 (N_9211,N_1854,N_479);
xor U9212 (N_9212,N_1146,N_1410);
or U9213 (N_9213,N_4320,N_3346);
and U9214 (N_9214,N_2681,N_1561);
or U9215 (N_9215,N_3271,N_1927);
and U9216 (N_9216,N_4309,N_3904);
or U9217 (N_9217,N_4552,N_997);
nor U9218 (N_9218,N_1351,N_3244);
nand U9219 (N_9219,N_1952,N_4808);
and U9220 (N_9220,N_1713,N_4970);
and U9221 (N_9221,N_4,N_2938);
or U9222 (N_9222,N_2974,N_4869);
or U9223 (N_9223,N_4168,N_4576);
nand U9224 (N_9224,N_1800,N_4647);
or U9225 (N_9225,N_2235,N_2348);
nand U9226 (N_9226,N_2289,N_1971);
nor U9227 (N_9227,N_1763,N_874);
and U9228 (N_9228,N_675,N_2679);
nand U9229 (N_9229,N_1403,N_3646);
nor U9230 (N_9230,N_3299,N_3988);
or U9231 (N_9231,N_224,N_546);
and U9232 (N_9232,N_1060,N_4745);
or U9233 (N_9233,N_4893,N_1114);
nor U9234 (N_9234,N_3539,N_4990);
nor U9235 (N_9235,N_3014,N_2386);
or U9236 (N_9236,N_2823,N_874);
and U9237 (N_9237,N_517,N_4593);
nand U9238 (N_9238,N_3840,N_1299);
or U9239 (N_9239,N_1444,N_3148);
nor U9240 (N_9240,N_2824,N_2599);
nor U9241 (N_9241,N_3666,N_2132);
nor U9242 (N_9242,N_3115,N_3914);
nand U9243 (N_9243,N_3491,N_4218);
and U9244 (N_9244,N_2916,N_3514);
nor U9245 (N_9245,N_3266,N_1615);
and U9246 (N_9246,N_4105,N_1678);
or U9247 (N_9247,N_1480,N_4724);
nand U9248 (N_9248,N_2847,N_2328);
nor U9249 (N_9249,N_4894,N_637);
xor U9250 (N_9250,N_3727,N_2768);
or U9251 (N_9251,N_1096,N_2897);
or U9252 (N_9252,N_3545,N_3351);
or U9253 (N_9253,N_4947,N_1710);
xor U9254 (N_9254,N_2786,N_2444);
nand U9255 (N_9255,N_4382,N_2840);
and U9256 (N_9256,N_657,N_3999);
or U9257 (N_9257,N_4368,N_1187);
nor U9258 (N_9258,N_3842,N_540);
nor U9259 (N_9259,N_3691,N_4366);
nor U9260 (N_9260,N_864,N_2204);
nor U9261 (N_9261,N_1408,N_532);
nor U9262 (N_9262,N_1811,N_4917);
or U9263 (N_9263,N_506,N_909);
xor U9264 (N_9264,N_3899,N_4870);
or U9265 (N_9265,N_378,N_2423);
nand U9266 (N_9266,N_1991,N_3771);
or U9267 (N_9267,N_3261,N_4940);
or U9268 (N_9268,N_490,N_1958);
and U9269 (N_9269,N_558,N_4125);
and U9270 (N_9270,N_4595,N_3953);
nor U9271 (N_9271,N_56,N_1437);
xor U9272 (N_9272,N_2159,N_3408);
or U9273 (N_9273,N_4125,N_586);
or U9274 (N_9274,N_3406,N_4030);
nor U9275 (N_9275,N_3781,N_4507);
xnor U9276 (N_9276,N_2632,N_768);
nor U9277 (N_9277,N_4611,N_2409);
or U9278 (N_9278,N_2141,N_1649);
and U9279 (N_9279,N_3548,N_2183);
or U9280 (N_9280,N_3700,N_3748);
nor U9281 (N_9281,N_1193,N_1987);
xor U9282 (N_9282,N_796,N_1424);
or U9283 (N_9283,N_3657,N_1195);
or U9284 (N_9284,N_4650,N_1741);
nor U9285 (N_9285,N_3608,N_1429);
xnor U9286 (N_9286,N_4119,N_2028);
and U9287 (N_9287,N_1322,N_2900);
and U9288 (N_9288,N_3586,N_1624);
and U9289 (N_9289,N_4445,N_1213);
nand U9290 (N_9290,N_1787,N_1625);
nand U9291 (N_9291,N_4932,N_1563);
nor U9292 (N_9292,N_3110,N_3042);
nand U9293 (N_9293,N_3862,N_1235);
and U9294 (N_9294,N_3375,N_1217);
or U9295 (N_9295,N_3156,N_483);
and U9296 (N_9296,N_3602,N_3975);
or U9297 (N_9297,N_3747,N_4725);
and U9298 (N_9298,N_3625,N_4542);
xor U9299 (N_9299,N_1406,N_2585);
nand U9300 (N_9300,N_3781,N_912);
xor U9301 (N_9301,N_260,N_3230);
nor U9302 (N_9302,N_2274,N_581);
nor U9303 (N_9303,N_580,N_4304);
nand U9304 (N_9304,N_3044,N_2806);
nand U9305 (N_9305,N_2793,N_162);
or U9306 (N_9306,N_532,N_3821);
or U9307 (N_9307,N_3310,N_4221);
and U9308 (N_9308,N_4398,N_1985);
or U9309 (N_9309,N_2907,N_4878);
nor U9310 (N_9310,N_4774,N_4007);
xnor U9311 (N_9311,N_553,N_3263);
nor U9312 (N_9312,N_4767,N_1396);
or U9313 (N_9313,N_683,N_183);
nand U9314 (N_9314,N_2375,N_2212);
or U9315 (N_9315,N_3105,N_4441);
nand U9316 (N_9316,N_1166,N_3488);
or U9317 (N_9317,N_4908,N_1021);
nand U9318 (N_9318,N_1735,N_2463);
nand U9319 (N_9319,N_853,N_3017);
nor U9320 (N_9320,N_3688,N_1703);
and U9321 (N_9321,N_3996,N_2778);
nand U9322 (N_9322,N_670,N_1463);
nor U9323 (N_9323,N_3349,N_3531);
nor U9324 (N_9324,N_3762,N_3305);
or U9325 (N_9325,N_4492,N_2668);
and U9326 (N_9326,N_2268,N_2451);
or U9327 (N_9327,N_3173,N_4192);
nor U9328 (N_9328,N_4697,N_3636);
nand U9329 (N_9329,N_1252,N_3016);
nand U9330 (N_9330,N_2757,N_2942);
xnor U9331 (N_9331,N_810,N_1645);
nor U9332 (N_9332,N_4362,N_857);
nor U9333 (N_9333,N_4875,N_2126);
or U9334 (N_9334,N_3753,N_1438);
or U9335 (N_9335,N_3111,N_4003);
nor U9336 (N_9336,N_3657,N_1434);
nor U9337 (N_9337,N_2496,N_289);
xor U9338 (N_9338,N_69,N_2202);
nand U9339 (N_9339,N_599,N_3892);
nor U9340 (N_9340,N_3539,N_2048);
xor U9341 (N_9341,N_1818,N_3882);
nand U9342 (N_9342,N_2269,N_4119);
and U9343 (N_9343,N_201,N_2964);
and U9344 (N_9344,N_2316,N_1885);
and U9345 (N_9345,N_3025,N_2413);
or U9346 (N_9346,N_3570,N_1704);
xnor U9347 (N_9347,N_1904,N_2601);
nand U9348 (N_9348,N_2622,N_318);
and U9349 (N_9349,N_870,N_4526);
nor U9350 (N_9350,N_2676,N_2349);
and U9351 (N_9351,N_962,N_4228);
xor U9352 (N_9352,N_1004,N_538);
or U9353 (N_9353,N_4025,N_2342);
nor U9354 (N_9354,N_1535,N_3408);
and U9355 (N_9355,N_17,N_2117);
and U9356 (N_9356,N_504,N_1800);
nand U9357 (N_9357,N_4626,N_2039);
and U9358 (N_9358,N_433,N_4492);
and U9359 (N_9359,N_590,N_2718);
nand U9360 (N_9360,N_1227,N_1181);
or U9361 (N_9361,N_4186,N_3049);
and U9362 (N_9362,N_3705,N_4128);
or U9363 (N_9363,N_2691,N_2275);
nor U9364 (N_9364,N_3685,N_4769);
nor U9365 (N_9365,N_2559,N_3742);
xnor U9366 (N_9366,N_2736,N_979);
and U9367 (N_9367,N_2766,N_783);
or U9368 (N_9368,N_2235,N_3519);
or U9369 (N_9369,N_3006,N_3854);
nand U9370 (N_9370,N_4188,N_1088);
or U9371 (N_9371,N_1303,N_423);
and U9372 (N_9372,N_316,N_2022);
and U9373 (N_9373,N_1293,N_1852);
nor U9374 (N_9374,N_2191,N_1886);
nand U9375 (N_9375,N_4300,N_2654);
nor U9376 (N_9376,N_3893,N_3288);
or U9377 (N_9377,N_375,N_2496);
nand U9378 (N_9378,N_4171,N_3029);
nor U9379 (N_9379,N_708,N_1690);
and U9380 (N_9380,N_4036,N_985);
nand U9381 (N_9381,N_722,N_1092);
and U9382 (N_9382,N_4868,N_2365);
nand U9383 (N_9383,N_1989,N_913);
nor U9384 (N_9384,N_492,N_446);
or U9385 (N_9385,N_4716,N_1716);
nor U9386 (N_9386,N_4693,N_1238);
nor U9387 (N_9387,N_3886,N_849);
and U9388 (N_9388,N_19,N_1339);
or U9389 (N_9389,N_2301,N_633);
or U9390 (N_9390,N_3936,N_2615);
and U9391 (N_9391,N_1642,N_1580);
nor U9392 (N_9392,N_1360,N_384);
nand U9393 (N_9393,N_2009,N_998);
nor U9394 (N_9394,N_220,N_1937);
nor U9395 (N_9395,N_3759,N_4942);
nand U9396 (N_9396,N_765,N_4983);
nor U9397 (N_9397,N_1446,N_1100);
or U9398 (N_9398,N_1428,N_4793);
or U9399 (N_9399,N_625,N_4181);
or U9400 (N_9400,N_166,N_3547);
xnor U9401 (N_9401,N_804,N_220);
and U9402 (N_9402,N_3824,N_2944);
and U9403 (N_9403,N_4712,N_300);
and U9404 (N_9404,N_3063,N_1241);
nor U9405 (N_9405,N_3103,N_1411);
nand U9406 (N_9406,N_199,N_4583);
or U9407 (N_9407,N_37,N_2620);
nand U9408 (N_9408,N_2688,N_3838);
nand U9409 (N_9409,N_2124,N_4381);
and U9410 (N_9410,N_184,N_1609);
and U9411 (N_9411,N_4442,N_4748);
nor U9412 (N_9412,N_4827,N_1618);
and U9413 (N_9413,N_1065,N_3988);
and U9414 (N_9414,N_3142,N_1897);
or U9415 (N_9415,N_1054,N_1853);
and U9416 (N_9416,N_4829,N_2691);
nor U9417 (N_9417,N_2556,N_3662);
and U9418 (N_9418,N_2645,N_215);
and U9419 (N_9419,N_4651,N_3669);
xnor U9420 (N_9420,N_511,N_2245);
or U9421 (N_9421,N_2116,N_439);
nor U9422 (N_9422,N_1206,N_3573);
or U9423 (N_9423,N_3318,N_4493);
or U9424 (N_9424,N_4659,N_1769);
or U9425 (N_9425,N_58,N_2017);
and U9426 (N_9426,N_363,N_756);
and U9427 (N_9427,N_2168,N_3262);
or U9428 (N_9428,N_4539,N_3910);
or U9429 (N_9429,N_1839,N_256);
and U9430 (N_9430,N_3100,N_2597);
and U9431 (N_9431,N_284,N_431);
or U9432 (N_9432,N_274,N_1758);
or U9433 (N_9433,N_136,N_617);
nor U9434 (N_9434,N_4047,N_3127);
nor U9435 (N_9435,N_1598,N_793);
nor U9436 (N_9436,N_3698,N_2440);
nor U9437 (N_9437,N_1975,N_2497);
xnor U9438 (N_9438,N_4563,N_2039);
nor U9439 (N_9439,N_679,N_2643);
or U9440 (N_9440,N_4342,N_3145);
nand U9441 (N_9441,N_2772,N_4078);
and U9442 (N_9442,N_2608,N_3359);
and U9443 (N_9443,N_504,N_704);
nor U9444 (N_9444,N_1966,N_3751);
or U9445 (N_9445,N_1242,N_3221);
or U9446 (N_9446,N_749,N_385);
nand U9447 (N_9447,N_105,N_2518);
nor U9448 (N_9448,N_4770,N_2377);
nor U9449 (N_9449,N_2531,N_4075);
and U9450 (N_9450,N_1443,N_2629);
or U9451 (N_9451,N_4849,N_2078);
nand U9452 (N_9452,N_1650,N_4455);
nor U9453 (N_9453,N_2839,N_429);
or U9454 (N_9454,N_2752,N_345);
and U9455 (N_9455,N_3969,N_3745);
or U9456 (N_9456,N_3855,N_2495);
and U9457 (N_9457,N_439,N_1737);
xor U9458 (N_9458,N_1175,N_4234);
xor U9459 (N_9459,N_1791,N_1891);
nor U9460 (N_9460,N_3286,N_1989);
nor U9461 (N_9461,N_3284,N_1131);
and U9462 (N_9462,N_1395,N_2936);
and U9463 (N_9463,N_3808,N_1179);
nor U9464 (N_9464,N_617,N_3966);
nand U9465 (N_9465,N_2583,N_2341);
and U9466 (N_9466,N_2537,N_1136);
and U9467 (N_9467,N_3747,N_329);
nor U9468 (N_9468,N_1135,N_1133);
and U9469 (N_9469,N_2919,N_783);
nand U9470 (N_9470,N_4099,N_4947);
xor U9471 (N_9471,N_507,N_4343);
nand U9472 (N_9472,N_136,N_2287);
nand U9473 (N_9473,N_888,N_2830);
nor U9474 (N_9474,N_459,N_638);
nor U9475 (N_9475,N_3546,N_875);
nand U9476 (N_9476,N_3364,N_2722);
nand U9477 (N_9477,N_4472,N_2692);
nor U9478 (N_9478,N_4646,N_2361);
or U9479 (N_9479,N_4220,N_3103);
xor U9480 (N_9480,N_55,N_2917);
or U9481 (N_9481,N_2006,N_3564);
nor U9482 (N_9482,N_2781,N_4668);
nor U9483 (N_9483,N_3887,N_4225);
nand U9484 (N_9484,N_4052,N_2059);
nand U9485 (N_9485,N_2501,N_3383);
or U9486 (N_9486,N_487,N_3122);
or U9487 (N_9487,N_3316,N_4475);
nor U9488 (N_9488,N_4699,N_4705);
xor U9489 (N_9489,N_617,N_1308);
and U9490 (N_9490,N_4811,N_3699);
or U9491 (N_9491,N_4620,N_2363);
and U9492 (N_9492,N_1175,N_191);
nor U9493 (N_9493,N_2525,N_858);
nor U9494 (N_9494,N_3427,N_3373);
nor U9495 (N_9495,N_1703,N_1070);
xor U9496 (N_9496,N_1102,N_3055);
or U9497 (N_9497,N_4214,N_1881);
nor U9498 (N_9498,N_2460,N_2251);
nand U9499 (N_9499,N_481,N_3929);
or U9500 (N_9500,N_4145,N_4410);
xnor U9501 (N_9501,N_3682,N_2764);
or U9502 (N_9502,N_3091,N_1737);
and U9503 (N_9503,N_4525,N_584);
nand U9504 (N_9504,N_1027,N_2478);
xnor U9505 (N_9505,N_370,N_1990);
or U9506 (N_9506,N_2418,N_2569);
and U9507 (N_9507,N_1962,N_3331);
xnor U9508 (N_9508,N_2566,N_3172);
nor U9509 (N_9509,N_2609,N_4689);
nand U9510 (N_9510,N_1902,N_642);
nand U9511 (N_9511,N_954,N_616);
and U9512 (N_9512,N_970,N_1862);
or U9513 (N_9513,N_4944,N_1322);
nor U9514 (N_9514,N_2483,N_2520);
and U9515 (N_9515,N_4823,N_1887);
and U9516 (N_9516,N_3893,N_2612);
nor U9517 (N_9517,N_3770,N_1855);
or U9518 (N_9518,N_3787,N_3317);
nand U9519 (N_9519,N_832,N_719);
and U9520 (N_9520,N_1462,N_2081);
nand U9521 (N_9521,N_44,N_4470);
or U9522 (N_9522,N_4382,N_2686);
nor U9523 (N_9523,N_4177,N_4534);
or U9524 (N_9524,N_1040,N_966);
nand U9525 (N_9525,N_1845,N_2331);
or U9526 (N_9526,N_4323,N_3940);
xnor U9527 (N_9527,N_3680,N_1414);
and U9528 (N_9528,N_2293,N_1200);
and U9529 (N_9529,N_3395,N_2394);
nor U9530 (N_9530,N_3560,N_4398);
and U9531 (N_9531,N_299,N_3091);
nor U9532 (N_9532,N_1294,N_4484);
and U9533 (N_9533,N_2067,N_2948);
or U9534 (N_9534,N_4512,N_1209);
nand U9535 (N_9535,N_3108,N_2865);
or U9536 (N_9536,N_1412,N_132);
or U9537 (N_9537,N_3514,N_2190);
or U9538 (N_9538,N_4881,N_2343);
nand U9539 (N_9539,N_1805,N_3489);
nor U9540 (N_9540,N_3928,N_2591);
and U9541 (N_9541,N_1783,N_2148);
nor U9542 (N_9542,N_3555,N_4439);
or U9543 (N_9543,N_1614,N_1237);
nand U9544 (N_9544,N_998,N_4972);
or U9545 (N_9545,N_3936,N_172);
and U9546 (N_9546,N_3480,N_48);
or U9547 (N_9547,N_3804,N_1941);
or U9548 (N_9548,N_3831,N_1801);
nor U9549 (N_9549,N_3876,N_1908);
or U9550 (N_9550,N_4047,N_3582);
xor U9551 (N_9551,N_1631,N_518);
nor U9552 (N_9552,N_2421,N_19);
nor U9553 (N_9553,N_3419,N_3159);
or U9554 (N_9554,N_3137,N_4566);
or U9555 (N_9555,N_2413,N_891);
nor U9556 (N_9556,N_2993,N_2678);
nor U9557 (N_9557,N_1445,N_3603);
or U9558 (N_9558,N_687,N_3958);
nor U9559 (N_9559,N_979,N_4672);
nand U9560 (N_9560,N_1693,N_4661);
and U9561 (N_9561,N_4309,N_4692);
or U9562 (N_9562,N_1695,N_4367);
nand U9563 (N_9563,N_246,N_4339);
nand U9564 (N_9564,N_3438,N_881);
nor U9565 (N_9565,N_1398,N_3882);
xor U9566 (N_9566,N_4025,N_1748);
nand U9567 (N_9567,N_4159,N_83);
or U9568 (N_9568,N_2900,N_1965);
nand U9569 (N_9569,N_2342,N_2885);
or U9570 (N_9570,N_1036,N_1889);
and U9571 (N_9571,N_499,N_817);
or U9572 (N_9572,N_1644,N_4896);
and U9573 (N_9573,N_2159,N_3113);
nor U9574 (N_9574,N_4955,N_655);
nor U9575 (N_9575,N_1923,N_2491);
or U9576 (N_9576,N_3083,N_3616);
nor U9577 (N_9577,N_3482,N_495);
xnor U9578 (N_9578,N_1417,N_1147);
and U9579 (N_9579,N_1749,N_3462);
or U9580 (N_9580,N_4037,N_3120);
and U9581 (N_9581,N_4883,N_2549);
xnor U9582 (N_9582,N_73,N_4371);
or U9583 (N_9583,N_3848,N_3938);
nor U9584 (N_9584,N_8,N_3832);
and U9585 (N_9585,N_2702,N_2592);
nor U9586 (N_9586,N_1449,N_3771);
nor U9587 (N_9587,N_4358,N_3530);
and U9588 (N_9588,N_1951,N_637);
or U9589 (N_9589,N_3921,N_925);
and U9590 (N_9590,N_1969,N_4513);
and U9591 (N_9591,N_4224,N_2596);
and U9592 (N_9592,N_2217,N_2700);
and U9593 (N_9593,N_3272,N_456);
nor U9594 (N_9594,N_3937,N_3215);
or U9595 (N_9595,N_268,N_4645);
or U9596 (N_9596,N_1629,N_4393);
or U9597 (N_9597,N_1321,N_1430);
and U9598 (N_9598,N_874,N_1500);
nand U9599 (N_9599,N_4711,N_479);
xnor U9600 (N_9600,N_366,N_2298);
nand U9601 (N_9601,N_2260,N_4959);
and U9602 (N_9602,N_2658,N_930);
nor U9603 (N_9603,N_4768,N_2683);
xor U9604 (N_9604,N_3281,N_4903);
or U9605 (N_9605,N_3395,N_2783);
or U9606 (N_9606,N_3736,N_2022);
and U9607 (N_9607,N_329,N_2499);
and U9608 (N_9608,N_943,N_440);
nand U9609 (N_9609,N_511,N_143);
or U9610 (N_9610,N_4717,N_4470);
nor U9611 (N_9611,N_2068,N_2076);
or U9612 (N_9612,N_3299,N_1445);
or U9613 (N_9613,N_1560,N_2613);
or U9614 (N_9614,N_3480,N_4654);
xnor U9615 (N_9615,N_1440,N_2075);
or U9616 (N_9616,N_1067,N_2203);
xor U9617 (N_9617,N_2965,N_4708);
nand U9618 (N_9618,N_3726,N_4027);
and U9619 (N_9619,N_1389,N_1403);
and U9620 (N_9620,N_997,N_726);
or U9621 (N_9621,N_1824,N_3016);
or U9622 (N_9622,N_316,N_2572);
nor U9623 (N_9623,N_3729,N_4188);
and U9624 (N_9624,N_4500,N_2620);
xor U9625 (N_9625,N_2646,N_3285);
and U9626 (N_9626,N_4271,N_249);
and U9627 (N_9627,N_4649,N_4150);
xor U9628 (N_9628,N_716,N_3671);
xor U9629 (N_9629,N_4208,N_2681);
or U9630 (N_9630,N_1368,N_1063);
and U9631 (N_9631,N_4888,N_2434);
or U9632 (N_9632,N_2180,N_1039);
and U9633 (N_9633,N_2078,N_3927);
nand U9634 (N_9634,N_4057,N_3906);
or U9635 (N_9635,N_218,N_4100);
nor U9636 (N_9636,N_3006,N_37);
or U9637 (N_9637,N_3096,N_2432);
and U9638 (N_9638,N_32,N_3660);
or U9639 (N_9639,N_671,N_2320);
nand U9640 (N_9640,N_973,N_358);
and U9641 (N_9641,N_3040,N_4276);
xor U9642 (N_9642,N_718,N_2116);
nor U9643 (N_9643,N_2111,N_3221);
xor U9644 (N_9644,N_1845,N_3807);
and U9645 (N_9645,N_4687,N_2074);
and U9646 (N_9646,N_3844,N_4439);
nor U9647 (N_9647,N_2426,N_2675);
xor U9648 (N_9648,N_4132,N_4274);
and U9649 (N_9649,N_4390,N_477);
xor U9650 (N_9650,N_2873,N_3156);
nor U9651 (N_9651,N_4451,N_2890);
xor U9652 (N_9652,N_546,N_1354);
nand U9653 (N_9653,N_2522,N_4019);
nand U9654 (N_9654,N_80,N_1528);
nor U9655 (N_9655,N_4003,N_2311);
and U9656 (N_9656,N_434,N_3617);
nor U9657 (N_9657,N_358,N_1488);
and U9658 (N_9658,N_1351,N_3456);
xnor U9659 (N_9659,N_3188,N_1830);
nand U9660 (N_9660,N_2075,N_2638);
or U9661 (N_9661,N_694,N_3317);
and U9662 (N_9662,N_3206,N_2104);
and U9663 (N_9663,N_864,N_2629);
xor U9664 (N_9664,N_753,N_2847);
xor U9665 (N_9665,N_1054,N_3259);
nand U9666 (N_9666,N_4084,N_69);
or U9667 (N_9667,N_4899,N_2869);
and U9668 (N_9668,N_880,N_3063);
or U9669 (N_9669,N_4372,N_773);
nor U9670 (N_9670,N_4204,N_2366);
or U9671 (N_9671,N_725,N_4326);
and U9672 (N_9672,N_2464,N_378);
nand U9673 (N_9673,N_2879,N_2699);
nand U9674 (N_9674,N_532,N_3869);
nand U9675 (N_9675,N_4736,N_2018);
xor U9676 (N_9676,N_183,N_251);
nor U9677 (N_9677,N_1416,N_1072);
nand U9678 (N_9678,N_2570,N_4426);
or U9679 (N_9679,N_920,N_4622);
and U9680 (N_9680,N_2894,N_4890);
nor U9681 (N_9681,N_2282,N_1778);
nand U9682 (N_9682,N_3319,N_4044);
and U9683 (N_9683,N_3833,N_3047);
and U9684 (N_9684,N_1432,N_2496);
nor U9685 (N_9685,N_3080,N_177);
nor U9686 (N_9686,N_35,N_2717);
nor U9687 (N_9687,N_1827,N_1571);
nor U9688 (N_9688,N_3651,N_2394);
nand U9689 (N_9689,N_1412,N_2745);
xnor U9690 (N_9690,N_4650,N_2177);
nor U9691 (N_9691,N_1354,N_2145);
or U9692 (N_9692,N_344,N_87);
and U9693 (N_9693,N_697,N_1439);
nand U9694 (N_9694,N_4424,N_3199);
nand U9695 (N_9695,N_1063,N_3840);
nor U9696 (N_9696,N_1872,N_3740);
or U9697 (N_9697,N_1288,N_3824);
or U9698 (N_9698,N_1612,N_911);
and U9699 (N_9699,N_1968,N_3679);
xor U9700 (N_9700,N_1344,N_1512);
nand U9701 (N_9701,N_1585,N_4723);
or U9702 (N_9702,N_532,N_990);
or U9703 (N_9703,N_2248,N_2953);
nand U9704 (N_9704,N_3383,N_332);
and U9705 (N_9705,N_4854,N_2918);
and U9706 (N_9706,N_2230,N_3877);
and U9707 (N_9707,N_746,N_4444);
nor U9708 (N_9708,N_3941,N_2964);
xor U9709 (N_9709,N_1754,N_3296);
nor U9710 (N_9710,N_2975,N_2965);
nor U9711 (N_9711,N_2455,N_3679);
and U9712 (N_9712,N_3233,N_4233);
nor U9713 (N_9713,N_2306,N_492);
or U9714 (N_9714,N_2235,N_3065);
xor U9715 (N_9715,N_43,N_2862);
or U9716 (N_9716,N_4880,N_413);
nand U9717 (N_9717,N_3349,N_4012);
nand U9718 (N_9718,N_3152,N_2615);
nand U9719 (N_9719,N_3115,N_310);
or U9720 (N_9720,N_3044,N_4561);
or U9721 (N_9721,N_1691,N_2002);
or U9722 (N_9722,N_3816,N_770);
or U9723 (N_9723,N_975,N_835);
nor U9724 (N_9724,N_1503,N_487);
and U9725 (N_9725,N_671,N_1241);
nand U9726 (N_9726,N_2820,N_2019);
nor U9727 (N_9727,N_2494,N_4455);
or U9728 (N_9728,N_4183,N_2536);
or U9729 (N_9729,N_3902,N_3148);
and U9730 (N_9730,N_387,N_3080);
xor U9731 (N_9731,N_3043,N_1094);
and U9732 (N_9732,N_484,N_68);
nand U9733 (N_9733,N_2664,N_4426);
and U9734 (N_9734,N_743,N_3465);
nor U9735 (N_9735,N_1875,N_3378);
or U9736 (N_9736,N_3056,N_1253);
xnor U9737 (N_9737,N_217,N_1129);
nor U9738 (N_9738,N_4548,N_1618);
nor U9739 (N_9739,N_45,N_2051);
and U9740 (N_9740,N_1153,N_4532);
nor U9741 (N_9741,N_510,N_2707);
nor U9742 (N_9742,N_1747,N_791);
nand U9743 (N_9743,N_473,N_2096);
nand U9744 (N_9744,N_2596,N_4240);
nor U9745 (N_9745,N_1103,N_3611);
nand U9746 (N_9746,N_730,N_3276);
nor U9747 (N_9747,N_3611,N_1115);
nor U9748 (N_9748,N_3572,N_3996);
and U9749 (N_9749,N_3752,N_3948);
xor U9750 (N_9750,N_3854,N_1189);
nand U9751 (N_9751,N_1893,N_234);
and U9752 (N_9752,N_4156,N_4379);
nand U9753 (N_9753,N_401,N_2131);
or U9754 (N_9754,N_1587,N_1232);
nand U9755 (N_9755,N_1180,N_4609);
nand U9756 (N_9756,N_3497,N_4253);
nand U9757 (N_9757,N_918,N_3940);
nor U9758 (N_9758,N_4443,N_1195);
or U9759 (N_9759,N_4075,N_54);
nand U9760 (N_9760,N_714,N_1000);
xor U9761 (N_9761,N_577,N_4408);
or U9762 (N_9762,N_3376,N_1008);
and U9763 (N_9763,N_1616,N_2102);
and U9764 (N_9764,N_4129,N_4344);
nor U9765 (N_9765,N_4,N_844);
xor U9766 (N_9766,N_1945,N_3562);
nand U9767 (N_9767,N_1841,N_1497);
nand U9768 (N_9768,N_2123,N_3156);
or U9769 (N_9769,N_3648,N_4692);
or U9770 (N_9770,N_144,N_1243);
xnor U9771 (N_9771,N_196,N_832);
and U9772 (N_9772,N_1697,N_764);
or U9773 (N_9773,N_2310,N_3078);
and U9774 (N_9774,N_4600,N_4273);
nand U9775 (N_9775,N_316,N_3344);
nand U9776 (N_9776,N_2497,N_1121);
nor U9777 (N_9777,N_1035,N_3375);
nand U9778 (N_9778,N_4118,N_3796);
nand U9779 (N_9779,N_3065,N_848);
nand U9780 (N_9780,N_1433,N_2700);
or U9781 (N_9781,N_1701,N_456);
and U9782 (N_9782,N_944,N_1148);
nor U9783 (N_9783,N_3544,N_4410);
and U9784 (N_9784,N_4017,N_2056);
nor U9785 (N_9785,N_1274,N_4162);
and U9786 (N_9786,N_4656,N_2846);
nand U9787 (N_9787,N_38,N_3368);
nand U9788 (N_9788,N_4910,N_4841);
nand U9789 (N_9789,N_46,N_2464);
xnor U9790 (N_9790,N_1883,N_501);
or U9791 (N_9791,N_3877,N_4221);
nor U9792 (N_9792,N_1893,N_2765);
nor U9793 (N_9793,N_3910,N_3350);
nor U9794 (N_9794,N_4005,N_2513);
and U9795 (N_9795,N_4136,N_2804);
nor U9796 (N_9796,N_1891,N_849);
and U9797 (N_9797,N_1505,N_2896);
or U9798 (N_9798,N_2103,N_153);
or U9799 (N_9799,N_2180,N_1478);
and U9800 (N_9800,N_2177,N_283);
nor U9801 (N_9801,N_4698,N_2175);
or U9802 (N_9802,N_3933,N_128);
nand U9803 (N_9803,N_498,N_2281);
and U9804 (N_9804,N_4608,N_1546);
nor U9805 (N_9805,N_1903,N_2897);
xor U9806 (N_9806,N_4302,N_3982);
xnor U9807 (N_9807,N_2779,N_4948);
nand U9808 (N_9808,N_3189,N_4293);
or U9809 (N_9809,N_3821,N_2515);
and U9810 (N_9810,N_880,N_3618);
nand U9811 (N_9811,N_1620,N_2492);
nor U9812 (N_9812,N_4274,N_4702);
and U9813 (N_9813,N_960,N_336);
and U9814 (N_9814,N_1389,N_1043);
and U9815 (N_9815,N_3132,N_581);
xor U9816 (N_9816,N_1902,N_4918);
or U9817 (N_9817,N_4910,N_1484);
nor U9818 (N_9818,N_103,N_3870);
nor U9819 (N_9819,N_2219,N_3208);
and U9820 (N_9820,N_1395,N_3246);
or U9821 (N_9821,N_718,N_1565);
nor U9822 (N_9822,N_4825,N_2087);
xnor U9823 (N_9823,N_4976,N_375);
or U9824 (N_9824,N_59,N_4558);
or U9825 (N_9825,N_4785,N_2003);
nand U9826 (N_9826,N_116,N_4690);
nor U9827 (N_9827,N_1302,N_4678);
nor U9828 (N_9828,N_2315,N_4416);
nor U9829 (N_9829,N_1420,N_4727);
nor U9830 (N_9830,N_70,N_4918);
or U9831 (N_9831,N_3622,N_4539);
and U9832 (N_9832,N_719,N_3994);
nand U9833 (N_9833,N_3910,N_4265);
nand U9834 (N_9834,N_1096,N_1263);
nor U9835 (N_9835,N_992,N_4693);
nor U9836 (N_9836,N_460,N_1892);
nand U9837 (N_9837,N_4679,N_1584);
nand U9838 (N_9838,N_718,N_2341);
and U9839 (N_9839,N_1597,N_4045);
nor U9840 (N_9840,N_4077,N_2491);
xor U9841 (N_9841,N_1448,N_2791);
and U9842 (N_9842,N_1578,N_373);
nor U9843 (N_9843,N_3314,N_1094);
nand U9844 (N_9844,N_3202,N_1077);
or U9845 (N_9845,N_3716,N_1597);
nor U9846 (N_9846,N_4904,N_4297);
and U9847 (N_9847,N_2118,N_4104);
nand U9848 (N_9848,N_1087,N_1965);
xor U9849 (N_9849,N_2895,N_447);
or U9850 (N_9850,N_2493,N_1239);
or U9851 (N_9851,N_1908,N_1865);
xnor U9852 (N_9852,N_3784,N_3906);
nand U9853 (N_9853,N_4517,N_934);
and U9854 (N_9854,N_4152,N_4044);
and U9855 (N_9855,N_2302,N_2629);
nor U9856 (N_9856,N_2242,N_2308);
nor U9857 (N_9857,N_4933,N_2884);
or U9858 (N_9858,N_798,N_1460);
nand U9859 (N_9859,N_1673,N_2645);
nor U9860 (N_9860,N_1383,N_1916);
and U9861 (N_9861,N_3927,N_4367);
or U9862 (N_9862,N_1061,N_146);
or U9863 (N_9863,N_3549,N_2011);
nor U9864 (N_9864,N_1694,N_4540);
nor U9865 (N_9865,N_3214,N_434);
nor U9866 (N_9866,N_1165,N_818);
xnor U9867 (N_9867,N_1379,N_3164);
or U9868 (N_9868,N_4781,N_2926);
nand U9869 (N_9869,N_3986,N_1849);
nor U9870 (N_9870,N_451,N_4463);
and U9871 (N_9871,N_2982,N_2882);
nand U9872 (N_9872,N_4433,N_4214);
and U9873 (N_9873,N_346,N_3258);
or U9874 (N_9874,N_3010,N_146);
and U9875 (N_9875,N_1810,N_3669);
nand U9876 (N_9876,N_4814,N_4883);
and U9877 (N_9877,N_2746,N_1907);
nand U9878 (N_9878,N_3678,N_4293);
nand U9879 (N_9879,N_2062,N_1374);
nand U9880 (N_9880,N_3357,N_3101);
and U9881 (N_9881,N_1586,N_554);
nand U9882 (N_9882,N_4391,N_3214);
and U9883 (N_9883,N_613,N_4095);
nor U9884 (N_9884,N_4114,N_2084);
or U9885 (N_9885,N_3999,N_2718);
and U9886 (N_9886,N_3806,N_2032);
nand U9887 (N_9887,N_4938,N_2993);
nand U9888 (N_9888,N_2165,N_3235);
and U9889 (N_9889,N_245,N_1907);
nand U9890 (N_9890,N_3489,N_1215);
nor U9891 (N_9891,N_1698,N_1015);
or U9892 (N_9892,N_894,N_2057);
or U9893 (N_9893,N_3314,N_574);
or U9894 (N_9894,N_4651,N_939);
xnor U9895 (N_9895,N_3971,N_3542);
and U9896 (N_9896,N_401,N_1054);
nor U9897 (N_9897,N_202,N_2254);
nand U9898 (N_9898,N_4794,N_1080);
or U9899 (N_9899,N_3693,N_1144);
or U9900 (N_9900,N_2212,N_3940);
or U9901 (N_9901,N_261,N_3796);
and U9902 (N_9902,N_4120,N_661);
nand U9903 (N_9903,N_1415,N_976);
nor U9904 (N_9904,N_4598,N_321);
nand U9905 (N_9905,N_3641,N_343);
and U9906 (N_9906,N_13,N_3250);
nand U9907 (N_9907,N_4132,N_2468);
and U9908 (N_9908,N_4139,N_4520);
xnor U9909 (N_9909,N_1559,N_1468);
nand U9910 (N_9910,N_2077,N_4333);
nand U9911 (N_9911,N_4913,N_4466);
nor U9912 (N_9912,N_2190,N_2242);
and U9913 (N_9913,N_1858,N_19);
xnor U9914 (N_9914,N_1587,N_3079);
and U9915 (N_9915,N_3798,N_2915);
or U9916 (N_9916,N_4574,N_231);
nand U9917 (N_9917,N_3153,N_2468);
nor U9918 (N_9918,N_2467,N_1716);
nor U9919 (N_9919,N_1307,N_817);
nand U9920 (N_9920,N_2889,N_2345);
and U9921 (N_9921,N_4759,N_4703);
and U9922 (N_9922,N_4544,N_2843);
or U9923 (N_9923,N_1591,N_1525);
nor U9924 (N_9924,N_4405,N_653);
and U9925 (N_9925,N_3920,N_3277);
nand U9926 (N_9926,N_2835,N_1995);
or U9927 (N_9927,N_4867,N_1317);
and U9928 (N_9928,N_2669,N_1807);
nand U9929 (N_9929,N_4262,N_232);
nor U9930 (N_9930,N_381,N_473);
nor U9931 (N_9931,N_4445,N_4154);
and U9932 (N_9932,N_3626,N_3214);
xnor U9933 (N_9933,N_2549,N_4474);
nand U9934 (N_9934,N_2538,N_244);
nor U9935 (N_9935,N_1323,N_4800);
nor U9936 (N_9936,N_1227,N_2831);
nor U9937 (N_9937,N_1412,N_2730);
nand U9938 (N_9938,N_3311,N_3648);
and U9939 (N_9939,N_3311,N_268);
or U9940 (N_9940,N_2343,N_2146);
nand U9941 (N_9941,N_2194,N_2113);
or U9942 (N_9942,N_2992,N_3740);
nand U9943 (N_9943,N_592,N_3080);
nor U9944 (N_9944,N_1487,N_2921);
or U9945 (N_9945,N_582,N_4754);
and U9946 (N_9946,N_758,N_4754);
or U9947 (N_9947,N_4983,N_2221);
nor U9948 (N_9948,N_1846,N_3309);
and U9949 (N_9949,N_1141,N_1390);
or U9950 (N_9950,N_3175,N_2926);
and U9951 (N_9951,N_2039,N_2223);
nor U9952 (N_9952,N_1595,N_2854);
nand U9953 (N_9953,N_3898,N_1994);
and U9954 (N_9954,N_1311,N_614);
or U9955 (N_9955,N_2453,N_1876);
or U9956 (N_9956,N_381,N_3775);
nor U9957 (N_9957,N_3220,N_3263);
nor U9958 (N_9958,N_1351,N_3392);
nand U9959 (N_9959,N_954,N_3016);
or U9960 (N_9960,N_3212,N_814);
nor U9961 (N_9961,N_2507,N_462);
and U9962 (N_9962,N_3762,N_3237);
nand U9963 (N_9963,N_4638,N_2948);
and U9964 (N_9964,N_3910,N_4538);
nand U9965 (N_9965,N_3510,N_3639);
nand U9966 (N_9966,N_2415,N_256);
or U9967 (N_9967,N_4838,N_741);
nand U9968 (N_9968,N_3630,N_4808);
or U9969 (N_9969,N_2420,N_221);
nor U9970 (N_9970,N_3622,N_3982);
or U9971 (N_9971,N_1774,N_2884);
nand U9972 (N_9972,N_3963,N_2034);
nand U9973 (N_9973,N_1482,N_4155);
nand U9974 (N_9974,N_2038,N_566);
nor U9975 (N_9975,N_1752,N_1091);
nor U9976 (N_9976,N_3938,N_4920);
and U9977 (N_9977,N_4716,N_3864);
nand U9978 (N_9978,N_4233,N_3882);
nor U9979 (N_9979,N_4689,N_3128);
or U9980 (N_9980,N_3748,N_190);
nand U9981 (N_9981,N_2577,N_876);
xor U9982 (N_9982,N_2647,N_1228);
and U9983 (N_9983,N_4694,N_4030);
nand U9984 (N_9984,N_2040,N_2177);
nor U9985 (N_9985,N_4919,N_1913);
nor U9986 (N_9986,N_894,N_2873);
nand U9987 (N_9987,N_3272,N_3309);
and U9988 (N_9988,N_3261,N_2633);
or U9989 (N_9989,N_4822,N_3796);
and U9990 (N_9990,N_977,N_3274);
nor U9991 (N_9991,N_1710,N_4571);
or U9992 (N_9992,N_3520,N_1053);
nand U9993 (N_9993,N_21,N_4766);
nor U9994 (N_9994,N_760,N_1300);
nand U9995 (N_9995,N_2736,N_3692);
nand U9996 (N_9996,N_1353,N_4878);
or U9997 (N_9997,N_300,N_4298);
and U9998 (N_9998,N_783,N_4716);
or U9999 (N_9999,N_4241,N_2390);
nand U10000 (N_10000,N_9093,N_9092);
nand U10001 (N_10001,N_8447,N_5223);
nand U10002 (N_10002,N_5539,N_9268);
or U10003 (N_10003,N_8184,N_8116);
nand U10004 (N_10004,N_8412,N_8309);
nor U10005 (N_10005,N_6821,N_5900);
and U10006 (N_10006,N_8435,N_5073);
nand U10007 (N_10007,N_7246,N_7377);
nand U10008 (N_10008,N_5801,N_6098);
nor U10009 (N_10009,N_7337,N_6058);
nand U10010 (N_10010,N_9238,N_5427);
or U10011 (N_10011,N_5270,N_9713);
xor U10012 (N_10012,N_8034,N_7473);
nand U10013 (N_10013,N_8994,N_8598);
and U10014 (N_10014,N_7595,N_5786);
or U10015 (N_10015,N_8332,N_7422);
nor U10016 (N_10016,N_8455,N_7856);
or U10017 (N_10017,N_5982,N_7723);
nand U10018 (N_10018,N_8000,N_5522);
xor U10019 (N_10019,N_8298,N_5456);
nand U10020 (N_10020,N_9070,N_9976);
nor U10021 (N_10021,N_9365,N_5703);
and U10022 (N_10022,N_9729,N_9431);
nor U10023 (N_10023,N_9981,N_6219);
or U10024 (N_10024,N_8896,N_5015);
and U10025 (N_10025,N_7431,N_7387);
xor U10026 (N_10026,N_8381,N_6707);
and U10027 (N_10027,N_5261,N_7861);
and U10028 (N_10028,N_7730,N_7604);
nand U10029 (N_10029,N_6012,N_6889);
or U10030 (N_10030,N_7352,N_6141);
and U10031 (N_10031,N_5082,N_6005);
or U10032 (N_10032,N_6506,N_7032);
and U10033 (N_10033,N_9900,N_8263);
and U10034 (N_10034,N_8901,N_8392);
nand U10035 (N_10035,N_9791,N_9775);
and U10036 (N_10036,N_7225,N_9044);
or U10037 (N_10037,N_7612,N_9979);
nor U10038 (N_10038,N_5376,N_5318);
or U10039 (N_10039,N_5398,N_8758);
or U10040 (N_10040,N_7209,N_7119);
nor U10041 (N_10041,N_8395,N_5624);
or U10042 (N_10042,N_6958,N_8905);
nor U10043 (N_10043,N_6049,N_6309);
or U10044 (N_10044,N_7654,N_8433);
or U10045 (N_10045,N_8658,N_8421);
nand U10046 (N_10046,N_7641,N_9228);
nor U10047 (N_10047,N_6087,N_9800);
and U10048 (N_10048,N_5290,N_9127);
and U10049 (N_10049,N_8159,N_5650);
or U10050 (N_10050,N_6205,N_5319);
nor U10051 (N_10051,N_8834,N_5127);
nor U10052 (N_10052,N_9465,N_7076);
or U10053 (N_10053,N_7778,N_8594);
or U10054 (N_10054,N_6969,N_8883);
and U10055 (N_10055,N_5680,N_5674);
and U10056 (N_10056,N_5083,N_8868);
and U10057 (N_10057,N_8647,N_5894);
and U10058 (N_10058,N_5193,N_5600);
nor U10059 (N_10059,N_6231,N_8308);
and U10060 (N_10060,N_7287,N_5219);
nor U10061 (N_10061,N_8441,N_6366);
nor U10062 (N_10062,N_5930,N_7622);
or U10063 (N_10063,N_8700,N_5014);
nor U10064 (N_10064,N_7136,N_6149);
nand U10065 (N_10065,N_8838,N_8873);
and U10066 (N_10066,N_8058,N_9869);
xnor U10067 (N_10067,N_9962,N_6666);
and U10068 (N_10068,N_7981,N_9653);
and U10069 (N_10069,N_9523,N_6314);
xor U10070 (N_10070,N_5050,N_7598);
nor U10071 (N_10071,N_7333,N_7334);
nand U10072 (N_10072,N_8836,N_5716);
and U10073 (N_10073,N_9757,N_8393);
nor U10074 (N_10074,N_6796,N_8375);
xnor U10075 (N_10075,N_5599,N_6382);
or U10076 (N_10076,N_8856,N_5307);
or U10077 (N_10077,N_8108,N_6802);
nor U10078 (N_10078,N_6625,N_9320);
or U10079 (N_10079,N_7794,N_9084);
nand U10080 (N_10080,N_6723,N_6959);
and U10081 (N_10081,N_5120,N_7220);
and U10082 (N_10082,N_5285,N_7293);
and U10083 (N_10083,N_6510,N_6851);
and U10084 (N_10084,N_5134,N_9796);
nand U10085 (N_10085,N_9876,N_9016);
xor U10086 (N_10086,N_5559,N_9363);
nand U10087 (N_10087,N_5577,N_7573);
nand U10088 (N_10088,N_6761,N_5934);
or U10089 (N_10089,N_6494,N_9087);
or U10090 (N_10090,N_6072,N_6916);
nand U10091 (N_10091,N_9546,N_8404);
or U10092 (N_10092,N_6080,N_7505);
and U10093 (N_10093,N_6700,N_8489);
nand U10094 (N_10094,N_5243,N_8466);
nor U10095 (N_10095,N_7330,N_7481);
xnor U10096 (N_10096,N_8270,N_7608);
nor U10097 (N_10097,N_5336,N_8220);
and U10098 (N_10098,N_8287,N_7355);
or U10099 (N_10099,N_7004,N_6412);
nor U10100 (N_10100,N_5288,N_7365);
xnor U10101 (N_10101,N_8065,N_9417);
nor U10102 (N_10102,N_8078,N_9132);
or U10103 (N_10103,N_7177,N_7303);
or U10104 (N_10104,N_7736,N_9797);
xnor U10105 (N_10105,N_8444,N_6957);
or U10106 (N_10106,N_9277,N_8004);
or U10107 (N_10107,N_7945,N_6227);
nor U10108 (N_10108,N_5545,N_5173);
nand U10109 (N_10109,N_5423,N_8888);
xnor U10110 (N_10110,N_6552,N_5094);
nand U10111 (N_10111,N_7851,N_7675);
xnor U10112 (N_10112,N_7357,N_9231);
nand U10113 (N_10113,N_7876,N_5171);
nor U10114 (N_10114,N_7682,N_6538);
nor U10115 (N_10115,N_6099,N_7253);
nor U10116 (N_10116,N_8234,N_8294);
nor U10117 (N_10117,N_6863,N_8338);
nor U10118 (N_10118,N_8218,N_6277);
xnor U10119 (N_10119,N_8509,N_8469);
nor U10120 (N_10120,N_9836,N_7688);
nand U10121 (N_10121,N_9780,N_5037);
or U10122 (N_10122,N_8321,N_6777);
or U10123 (N_10123,N_9234,N_5080);
or U10124 (N_10124,N_6711,N_5925);
nor U10125 (N_10125,N_5414,N_9590);
and U10126 (N_10126,N_7019,N_8349);
or U10127 (N_10127,N_8724,N_6931);
nor U10128 (N_10128,N_9740,N_5021);
nor U10129 (N_10129,N_9772,N_8819);
or U10130 (N_10130,N_6606,N_8961);
nand U10131 (N_10131,N_8286,N_7163);
and U10132 (N_10132,N_6319,N_5633);
and U10133 (N_10133,N_7074,N_5868);
xor U10134 (N_10134,N_8808,N_5890);
nand U10135 (N_10135,N_9897,N_5670);
or U10136 (N_10136,N_9715,N_9115);
or U10137 (N_10137,N_8477,N_6101);
nor U10138 (N_10138,N_7782,N_9873);
nor U10139 (N_10139,N_8747,N_7035);
xnor U10140 (N_10140,N_5400,N_6850);
xnor U10141 (N_10141,N_8824,N_9269);
xor U10142 (N_10142,N_7575,N_5441);
and U10143 (N_10143,N_6767,N_6428);
nand U10144 (N_10144,N_7819,N_8992);
xnor U10145 (N_10145,N_7788,N_9583);
or U10146 (N_10146,N_8314,N_9705);
and U10147 (N_10147,N_9743,N_6394);
and U10148 (N_10148,N_9709,N_6993);
and U10149 (N_10149,N_5353,N_7460);
xor U10150 (N_10150,N_5753,N_7503);
or U10151 (N_10151,N_8809,N_5097);
or U10152 (N_10152,N_7686,N_6987);
nor U10153 (N_10153,N_9942,N_7541);
and U10154 (N_10154,N_8170,N_8219);
nand U10155 (N_10155,N_9823,N_9236);
xnor U10156 (N_10156,N_5118,N_7314);
nand U10157 (N_10157,N_7551,N_5865);
nor U10158 (N_10158,N_5513,N_9028);
nand U10159 (N_10159,N_7058,N_9654);
nor U10160 (N_10160,N_6264,N_6455);
and U10161 (N_10161,N_7214,N_5342);
and U10162 (N_10162,N_6295,N_8514);
nor U10163 (N_10163,N_8796,N_7423);
and U10164 (N_10164,N_6832,N_7366);
or U10165 (N_10165,N_7168,N_9659);
or U10166 (N_10166,N_9700,N_5540);
and U10167 (N_10167,N_6335,N_9901);
nand U10168 (N_10168,N_7192,N_8984);
nor U10169 (N_10169,N_5326,N_9062);
nand U10170 (N_10170,N_9924,N_6939);
nand U10171 (N_10171,N_9121,N_9241);
or U10172 (N_10172,N_5845,N_8621);
nand U10173 (N_10173,N_6259,N_9160);
and U10174 (N_10174,N_6252,N_8068);
and U10175 (N_10175,N_9510,N_7112);
or U10176 (N_10176,N_9537,N_7984);
nor U10177 (N_10177,N_5755,N_8127);
nor U10178 (N_10178,N_7661,N_7956);
and U10179 (N_10179,N_9059,N_7180);
nand U10180 (N_10180,N_5280,N_5210);
xor U10181 (N_10181,N_6617,N_5343);
nor U10182 (N_10182,N_5308,N_9822);
and U10183 (N_10183,N_6733,N_8527);
or U10184 (N_10184,N_5681,N_6285);
or U10185 (N_10185,N_8342,N_5259);
and U10186 (N_10186,N_8979,N_8148);
nor U10187 (N_10187,N_7797,N_8832);
or U10188 (N_10188,N_6131,N_7637);
or U10189 (N_10189,N_9799,N_7687);
nand U10190 (N_10190,N_5146,N_8546);
nand U10191 (N_10191,N_7920,N_7444);
or U10192 (N_10192,N_6191,N_7063);
nor U10193 (N_10193,N_6649,N_7605);
nand U10194 (N_10194,N_9538,N_8966);
or U10195 (N_10195,N_6357,N_5517);
and U10196 (N_10196,N_5084,N_9903);
nand U10197 (N_10197,N_6561,N_7972);
nor U10198 (N_10198,N_6006,N_7060);
nand U10199 (N_10199,N_9141,N_6002);
nor U10200 (N_10200,N_8794,N_5999);
nand U10201 (N_10201,N_5964,N_7765);
nand U10202 (N_10202,N_5036,N_8307);
or U10203 (N_10203,N_6694,N_5740);
nand U10204 (N_10204,N_8419,N_8829);
nor U10205 (N_10205,N_5920,N_7010);
xnor U10206 (N_10206,N_9221,N_9877);
or U10207 (N_10207,N_6864,N_8776);
nor U10208 (N_10208,N_6887,N_7174);
or U10209 (N_10209,N_9894,N_8153);
nor U10210 (N_10210,N_9484,N_5834);
xnor U10211 (N_10211,N_7036,N_9854);
nor U10212 (N_10212,N_7581,N_9592);
and U10213 (N_10213,N_6396,N_6135);
and U10214 (N_10214,N_6464,N_8132);
nand U10215 (N_10215,N_8595,N_5238);
or U10216 (N_10216,N_9932,N_6981);
or U10217 (N_10217,N_5415,N_9022);
xor U10218 (N_10218,N_5076,N_7184);
or U10219 (N_10219,N_8432,N_9525);
xnor U10220 (N_10220,N_9349,N_6047);
nand U10221 (N_10221,N_9071,N_6329);
nand U10222 (N_10222,N_8122,N_6435);
nor U10223 (N_10223,N_9145,N_9315);
nand U10224 (N_10224,N_6325,N_7190);
nand U10225 (N_10225,N_8316,N_9374);
nor U10226 (N_10226,N_6615,N_6917);
nand U10227 (N_10227,N_7140,N_5085);
nor U10228 (N_10228,N_8329,N_7540);
nor U10229 (N_10229,N_5142,N_5265);
and U10230 (N_10230,N_8361,N_5231);
or U10231 (N_10231,N_8891,N_7409);
xor U10232 (N_10232,N_5821,N_6500);
and U10233 (N_10233,N_8448,N_6346);
and U10234 (N_10234,N_9898,N_9761);
and U10235 (N_10235,N_6288,N_8784);
xnor U10236 (N_10236,N_5425,N_8827);
nor U10237 (N_10237,N_9051,N_5725);
nand U10238 (N_10238,N_9636,N_8135);
and U10239 (N_10239,N_5018,N_9156);
nand U10240 (N_10240,N_6239,N_7594);
nand U10241 (N_10241,N_5711,N_7202);
nor U10242 (N_10242,N_5241,N_6833);
xor U10243 (N_10243,N_5370,N_8145);
or U10244 (N_10244,N_5516,N_7960);
nand U10245 (N_10245,N_5862,N_5025);
nand U10246 (N_10246,N_9007,N_8865);
nand U10247 (N_10247,N_8565,N_9909);
nand U10248 (N_10248,N_6161,N_8011);
nor U10249 (N_10249,N_7370,N_7850);
nand U10250 (N_10250,N_7285,N_6766);
nor U10251 (N_10251,N_8430,N_7371);
nand U10252 (N_10252,N_5067,N_7544);
xor U10253 (N_10253,N_9576,N_5974);
or U10254 (N_10254,N_5424,N_6210);
nor U10255 (N_10255,N_7345,N_7590);
or U10256 (N_10256,N_9435,N_6271);
or U10257 (N_10257,N_9809,N_8652);
or U10258 (N_10258,N_6417,N_8463);
nand U10259 (N_10259,N_7924,N_6838);
and U10260 (N_10260,N_8745,N_5731);
nand U10261 (N_10261,N_8975,N_6626);
nand U10262 (N_10262,N_5225,N_9929);
and U10263 (N_10263,N_6203,N_6248);
or U10264 (N_10264,N_9362,N_7832);
and U10265 (N_10265,N_9855,N_6964);
and U10266 (N_10266,N_9168,N_5388);
nor U10267 (N_10267,N_7006,N_7212);
and U10268 (N_10268,N_9112,N_5092);
nand U10269 (N_10269,N_9124,N_5813);
nor U10270 (N_10270,N_6572,N_9596);
nand U10271 (N_10271,N_7891,N_5978);
and U10272 (N_10272,N_9728,N_9805);
nand U10273 (N_10273,N_8426,N_5258);
xor U10274 (N_10274,N_5131,N_7243);
nor U10275 (N_10275,N_5064,N_6770);
nor U10276 (N_10276,N_8360,N_8212);
nand U10277 (N_10277,N_6204,N_5734);
nor U10278 (N_10278,N_6608,N_9214);
nand U10279 (N_10279,N_6923,N_5751);
xor U10280 (N_10280,N_5929,N_5121);
and U10281 (N_10281,N_6845,N_8738);
nand U10282 (N_10282,N_6318,N_7497);
xor U10283 (N_10283,N_9066,N_8233);
nand U10284 (N_10284,N_5768,N_8547);
nand U10285 (N_10285,N_6393,N_5159);
nor U10286 (N_10286,N_8549,N_5389);
nand U10287 (N_10287,N_7955,N_5792);
xor U10288 (N_10288,N_7729,N_5569);
or U10289 (N_10289,N_7635,N_9722);
nand U10290 (N_10290,N_7383,N_9196);
or U10291 (N_10291,N_9328,N_9184);
nor U10292 (N_10292,N_9993,N_8920);
nand U10293 (N_10293,N_9842,N_5857);
nor U10294 (N_10294,N_9853,N_8356);
or U10295 (N_10295,N_7615,N_5320);
xor U10296 (N_10296,N_5510,N_8492);
nand U10297 (N_10297,N_9001,N_8578);
nor U10298 (N_10298,N_5613,N_9216);
nor U10299 (N_10299,N_5799,N_5724);
or U10300 (N_10300,N_8271,N_9532);
nand U10301 (N_10301,N_6092,N_8845);
nor U10302 (N_10302,N_7773,N_6377);
and U10303 (N_10303,N_8908,N_8622);
nand U10304 (N_10304,N_8519,N_8552);
and U10305 (N_10305,N_6493,N_9543);
and U10306 (N_10306,N_9208,N_9192);
or U10307 (N_10307,N_6487,N_9283);
and U10308 (N_10308,N_8810,N_6880);
nor U10309 (N_10309,N_6787,N_9025);
or U10310 (N_10310,N_6320,N_7821);
and U10311 (N_10311,N_5068,N_6356);
nor U10312 (N_10312,N_7017,N_5739);
nor U10313 (N_10313,N_6590,N_7089);
or U10314 (N_10314,N_7676,N_9663);
and U10315 (N_10315,N_8493,N_9479);
and U10316 (N_10316,N_7659,N_6575);
and U10317 (N_10317,N_8198,N_5268);
xor U10318 (N_10318,N_5662,N_6890);
nor U10319 (N_10319,N_7562,N_5292);
nand U10320 (N_10320,N_5413,N_6673);
xnor U10321 (N_10321,N_5497,N_8762);
or U10322 (N_10322,N_7309,N_8215);
and U10323 (N_10323,N_7249,N_7815);
nand U10324 (N_10324,N_8767,N_5515);
nor U10325 (N_10325,N_6088,N_8670);
and U10326 (N_10326,N_9173,N_5224);
xor U10327 (N_10327,N_6730,N_7304);
nor U10328 (N_10328,N_9442,N_8079);
nand U10329 (N_10329,N_9542,N_6717);
or U10330 (N_10330,N_8005,N_6280);
and U10331 (N_10331,N_9864,N_8335);
or U10332 (N_10332,N_9978,N_5150);
and U10333 (N_10333,N_6429,N_8373);
and U10334 (N_10334,N_5010,N_8663);
and U10335 (N_10335,N_6508,N_8534);
nand U10336 (N_10336,N_6643,N_7609);
or U10337 (N_10337,N_9021,N_5181);
and U10338 (N_10338,N_9194,N_9263);
nor U10339 (N_10339,N_6984,N_9138);
nand U10340 (N_10340,N_7959,N_8781);
and U10341 (N_10341,N_7786,N_7325);
nand U10342 (N_10342,N_8502,N_6308);
and U10343 (N_10343,N_9865,N_8878);
nand U10344 (N_10344,N_8551,N_8821);
or U10345 (N_10345,N_5311,N_8968);
and U10346 (N_10346,N_7436,N_9925);
or U10347 (N_10347,N_7923,N_6491);
or U10348 (N_10348,N_7138,N_5723);
nand U10349 (N_10349,N_8111,N_7098);
xor U10350 (N_10350,N_7651,N_9222);
and U10351 (N_10351,N_5876,N_6297);
nor U10352 (N_10352,N_5034,N_7708);
nor U10353 (N_10353,N_7440,N_6118);
nand U10354 (N_10354,N_9755,N_7082);
xnor U10355 (N_10355,N_7488,N_9860);
nor U10356 (N_10356,N_9834,N_6482);
nor U10357 (N_10357,N_8450,N_5331);
nor U10358 (N_10358,N_6083,N_9446);
nor U10359 (N_10359,N_8788,N_9650);
nand U10360 (N_10360,N_9660,N_9848);
nor U10361 (N_10361,N_8452,N_5765);
nand U10362 (N_10362,N_8563,N_9563);
nor U10363 (N_10363,N_8561,N_6342);
and U10364 (N_10364,N_6650,N_8474);
nand U10365 (N_10365,N_5718,N_6143);
nor U10366 (N_10366,N_9426,N_9614);
and U10367 (N_10367,N_7029,N_6839);
nor U10368 (N_10368,N_6907,N_5757);
nand U10369 (N_10369,N_9770,N_9610);
or U10370 (N_10370,N_6165,N_7545);
xnor U10371 (N_10371,N_9181,N_6028);
or U10372 (N_10372,N_8117,N_8339);
or U10373 (N_10373,N_5209,N_5450);
or U10374 (N_10374,N_5374,N_6877);
nand U10375 (N_10375,N_6004,N_9344);
nand U10376 (N_10376,N_7644,N_7648);
nand U10377 (N_10377,N_6378,N_7106);
xor U10378 (N_10378,N_5759,N_8280);
nor U10379 (N_10379,N_7110,N_7234);
nand U10380 (N_10380,N_9451,N_5598);
or U10381 (N_10381,N_8445,N_6104);
nand U10382 (N_10382,N_5295,N_7295);
and U10383 (N_10383,N_9551,N_6411);
nor U10384 (N_10384,N_5781,N_5602);
nand U10385 (N_10385,N_8933,N_6648);
or U10386 (N_10386,N_6175,N_8853);
and U10387 (N_10387,N_6898,N_6499);
nand U10388 (N_10388,N_5445,N_5140);
or U10389 (N_10389,N_5991,N_6944);
or U10390 (N_10390,N_5428,N_7454);
nor U10391 (N_10391,N_6486,N_9685);
or U10392 (N_10392,N_6604,N_8768);
and U10393 (N_10393,N_7576,N_9314);
and U10394 (N_10394,N_6578,N_7529);
nand U10395 (N_10395,N_7747,N_6076);
and U10396 (N_10396,N_8383,N_6952);
nand U10397 (N_10397,N_5483,N_9104);
and U10398 (N_10398,N_5587,N_6284);
and U10399 (N_10399,N_8697,N_6278);
xnor U10400 (N_10400,N_7227,N_8709);
nor U10401 (N_10401,N_8195,N_7327);
nand U10402 (N_10402,N_8147,N_6128);
nand U10403 (N_10403,N_5610,N_5944);
xnor U10404 (N_10404,N_9109,N_9767);
or U10405 (N_10405,N_6609,N_8366);
nor U10406 (N_10406,N_8268,N_6915);
nor U10407 (N_10407,N_5283,N_6612);
nor U10408 (N_10408,N_5529,N_7874);
or U10409 (N_10409,N_5090,N_9436);
and U10410 (N_10410,N_5299,N_5583);
nor U10411 (N_10411,N_9731,N_9085);
xor U10412 (N_10412,N_9422,N_8748);
and U10413 (N_10413,N_6731,N_6808);
and U10414 (N_10414,N_5957,N_7419);
nor U10415 (N_10415,N_7415,N_7274);
nor U10416 (N_10416,N_7780,N_9516);
and U10417 (N_10417,N_5931,N_7754);
and U10418 (N_10418,N_9689,N_7939);
or U10419 (N_10419,N_7313,N_9662);
or U10420 (N_10420,N_5047,N_8753);
and U10421 (N_10421,N_6448,N_6168);
nor U10422 (N_10422,N_9180,N_9564);
nor U10423 (N_10423,N_7777,N_8012);
nor U10424 (N_10424,N_5381,N_9339);
and U10425 (N_10425,N_7618,N_7349);
nand U10426 (N_10426,N_9101,N_9667);
nand U10427 (N_10427,N_9644,N_5485);
nand U10428 (N_10428,N_7187,N_5861);
or U10429 (N_10429,N_5315,N_8730);
and U10430 (N_10430,N_6742,N_5380);
nor U10431 (N_10431,N_6370,N_7047);
nand U10432 (N_10432,N_6044,N_7629);
xor U10433 (N_10433,N_9769,N_5668);
or U10434 (N_10434,N_7181,N_8222);
and U10435 (N_10435,N_9704,N_8562);
or U10436 (N_10436,N_5864,N_5158);
and U10437 (N_10437,N_8624,N_8424);
nand U10438 (N_10438,N_6550,N_6790);
or U10439 (N_10439,N_9506,N_8168);
or U10440 (N_10440,N_8128,N_6975);
and U10441 (N_10441,N_8711,N_8027);
nand U10442 (N_10442,N_7455,N_6199);
and U10443 (N_10443,N_9683,N_7869);
or U10444 (N_10444,N_5479,N_9242);
or U10445 (N_10445,N_5779,N_7845);
xor U10446 (N_10446,N_5756,N_9130);
nand U10447 (N_10447,N_7271,N_8941);
nand U10448 (N_10448,N_8998,N_9255);
nor U10449 (N_10449,N_9079,N_7809);
nand U10450 (N_10450,N_6746,N_6654);
nor U10451 (N_10451,N_6275,N_7178);
nor U10452 (N_10452,N_8974,N_5760);
nor U10453 (N_10453,N_9649,N_5558);
and U10454 (N_10454,N_8760,N_8144);
and U10455 (N_10455,N_9633,N_6904);
nor U10456 (N_10456,N_7524,N_6444);
or U10457 (N_10457,N_6922,N_7697);
nand U10458 (N_10458,N_9992,N_7430);
nand U10459 (N_10459,N_5986,N_6762);
or U10460 (N_10460,N_8086,N_7302);
and U10461 (N_10461,N_6925,N_6462);
or U10462 (N_10462,N_7568,N_9091);
xnor U10463 (N_10463,N_8440,N_8325);
xnor U10464 (N_10464,N_8725,N_7559);
nand U10465 (N_10465,N_5321,N_5357);
nor U10466 (N_10466,N_5547,N_6662);
nor U10467 (N_10467,N_9814,N_9163);
nand U10468 (N_10468,N_8623,N_6639);
nor U10469 (N_10469,N_8706,N_7395);
or U10470 (N_10470,N_8851,N_7698);
or U10471 (N_10471,N_6465,N_6769);
or U10472 (N_10472,N_6977,N_9285);
or U10473 (N_10473,N_5761,N_5069);
xor U10474 (N_10474,N_6226,N_7701);
or U10475 (N_10475,N_6849,N_8620);
nand U10476 (N_10476,N_6886,N_5111);
or U10477 (N_10477,N_5685,N_7465);
or U10478 (N_10478,N_5625,N_6690);
nand U10479 (N_10479,N_6286,N_8283);
or U10480 (N_10480,N_7479,N_5783);
nand U10481 (N_10481,N_7783,N_7114);
and U10482 (N_10482,N_9878,N_7018);
xor U10483 (N_10483,N_8459,N_5623);
xor U10484 (N_10484,N_6685,N_7854);
nand U10485 (N_10485,N_6071,N_5538);
or U10486 (N_10486,N_8376,N_7397);
xnor U10487 (N_10487,N_9802,N_6292);
nand U10488 (N_10488,N_9024,N_9574);
xor U10489 (N_10489,N_6313,N_7707);
or U10490 (N_10490,N_5910,N_8893);
nand U10491 (N_10491,N_6995,N_5155);
nor U10492 (N_10492,N_6830,N_5970);
xnor U10493 (N_10493,N_6339,N_6438);
nor U10494 (N_10494,N_7012,N_5690);
nor U10495 (N_10495,N_7170,N_5256);
nor U10496 (N_10496,N_8110,N_8109);
and U10497 (N_10497,N_7808,N_6139);
nand U10498 (N_10498,N_9500,N_7752);
xnor U10499 (N_10499,N_5228,N_9535);
and U10500 (N_10500,N_6816,N_8370);
xnor U10501 (N_10501,N_5678,N_9777);
nand U10502 (N_10502,N_7160,N_9812);
and U10503 (N_10503,N_9201,N_6729);
nand U10504 (N_10504,N_5628,N_7224);
nor U10505 (N_10505,N_9927,N_5593);
nand U10506 (N_10506,N_6440,N_9625);
xnor U10507 (N_10507,N_6712,N_8648);
and U10508 (N_10508,N_9259,N_8482);
nor U10509 (N_10509,N_6069,N_5462);
nand U10510 (N_10510,N_8465,N_6737);
or U10511 (N_10511,N_6601,N_8969);
nor U10512 (N_10512,N_8284,N_5274);
and U10513 (N_10513,N_7962,N_8290);
xor U10514 (N_10514,N_8397,N_6812);
nand U10515 (N_10515,N_7805,N_5272);
nor U10516 (N_10516,N_5169,N_5561);
and U10517 (N_10517,N_5310,N_5498);
nor U10518 (N_10518,N_6413,N_9707);
or U10519 (N_10519,N_8291,N_7796);
xor U10520 (N_10520,N_9881,N_6225);
or U10521 (N_10521,N_7367,N_5654);
and U10522 (N_10522,N_8101,N_9473);
nor U10523 (N_10523,N_7310,N_5636);
nor U10524 (N_10524,N_9033,N_8499);
or U10525 (N_10525,N_5975,N_8363);
and U10526 (N_10526,N_9494,N_5156);
nand U10527 (N_10527,N_6803,N_9959);
and U10528 (N_10528,N_8491,N_9064);
and U10529 (N_10529,N_9969,N_5844);
and U10530 (N_10530,N_8657,N_6537);
nor U10531 (N_10531,N_7478,N_6543);
nor U10532 (N_10532,N_9988,N_7528);
nor U10533 (N_10533,N_6794,N_7746);
xnor U10534 (N_10534,N_9961,N_6775);
nor U10535 (N_10535,N_6784,N_8543);
nand U10536 (N_10536,N_7802,N_9586);
nand U10537 (N_10537,N_5129,N_5108);
and U10538 (N_10538,N_5530,N_7237);
xor U10539 (N_10539,N_6369,N_6591);
nor U10540 (N_10540,N_8679,N_5719);
nor U10541 (N_10541,N_7953,N_5300);
nand U10542 (N_10542,N_7484,N_9264);
nand U10543 (N_10543,N_5896,N_9017);
nor U10544 (N_10544,N_6772,N_9664);
or U10545 (N_10545,N_6119,N_7070);
and U10546 (N_10546,N_6095,N_8367);
or U10547 (N_10547,N_5165,N_5895);
and U10548 (N_10548,N_7897,N_5672);
or U10549 (N_10549,N_9159,N_6198);
xnor U10550 (N_10550,N_7554,N_6041);
or U10551 (N_10551,N_8391,N_9459);
xor U10552 (N_10552,N_7695,N_6437);
and U10553 (N_10553,N_8371,N_8311);
or U10554 (N_10554,N_7188,N_5297);
or U10555 (N_10555,N_9569,N_6527);
and U10556 (N_10556,N_5289,N_5431);
nand U10557 (N_10557,N_5713,N_7405);
nor U10558 (N_10558,N_5867,N_6375);
or U10559 (N_10559,N_9623,N_7871);
nor U10560 (N_10560,N_7589,N_8564);
nand U10561 (N_10561,N_7870,N_5178);
xor U10562 (N_10562,N_7647,N_5254);
nand U10563 (N_10563,N_8061,N_5434);
nor U10564 (N_10564,N_9675,N_8130);
and U10565 (N_10565,N_9191,N_6368);
nand U10566 (N_10566,N_7428,N_5962);
nor U10567 (N_10567,N_7597,N_8256);
nand U10568 (N_10568,N_7685,N_5494);
and U10569 (N_10569,N_6459,N_8226);
and U10570 (N_10570,N_8991,N_8579);
nor U10571 (N_10571,N_7968,N_8605);
xnor U10572 (N_10572,N_8055,N_7335);
nor U10573 (N_10573,N_5035,N_5885);
or U10574 (N_10574,N_9960,N_7584);
nand U10575 (N_10575,N_9453,N_7011);
and U10576 (N_10576,N_6683,N_5989);
or U10577 (N_10577,N_5113,N_5206);
and U10578 (N_10578,N_5179,N_5448);
and U10579 (N_10579,N_9237,N_9373);
or U10580 (N_10580,N_8866,N_6680);
xnor U10581 (N_10581,N_9301,N_8507);
or U10582 (N_10582,N_5746,N_9845);
nor U10583 (N_10583,N_9134,N_8948);
xnor U10584 (N_10584,N_6439,N_8945);
or U10585 (N_10585,N_7677,N_6888);
and U10586 (N_10586,N_7683,N_7265);
xnor U10587 (N_10587,N_6531,N_8051);
nand U10588 (N_10588,N_7893,N_6970);
and U10589 (N_10589,N_9454,N_9378);
nor U10590 (N_10590,N_6569,N_6709);
xnor U10591 (N_10591,N_6903,N_7526);
nor U10592 (N_10592,N_6333,N_8182);
nand U10593 (N_10593,N_9348,N_7221);
and U10594 (N_10594,N_6799,N_6351);
nor U10595 (N_10595,N_6189,N_8406);
nor U10596 (N_10596,N_6820,N_8940);
and U10597 (N_10597,N_5688,N_5446);
or U10598 (N_10598,N_7046,N_6122);
nor U10599 (N_10599,N_9493,N_8114);
and U10600 (N_10600,N_6420,N_9973);
or U10601 (N_10601,N_8511,N_5536);
and U10602 (N_10602,N_8713,N_7305);
nor U10603 (N_10603,N_8584,N_6502);
xnor U10604 (N_10604,N_5123,N_6138);
or U10605 (N_10605,N_6345,N_9225);
nand U10606 (N_10606,N_9498,N_8685);
xor U10607 (N_10607,N_8982,N_8299);
and U10608 (N_10608,N_8177,N_6557);
or U10609 (N_10609,N_5754,N_5470);
nor U10610 (N_10610,N_7083,N_9577);
and U10611 (N_10611,N_9832,N_9316);
nand U10612 (N_10612,N_6051,N_9794);
nand U10613 (N_10613,N_8718,N_8989);
xor U10614 (N_10614,N_6310,N_8942);
nor U10615 (N_10615,N_8458,N_5733);
or U10616 (N_10616,N_9045,N_5891);
or U10617 (N_10617,N_5617,N_9447);
nand U10618 (N_10618,N_8680,N_5042);
and U10619 (N_10619,N_8726,N_5619);
xor U10620 (N_10620,N_8364,N_5840);
xor U10621 (N_10621,N_6895,N_7418);
or U10622 (N_10622,N_9545,N_6042);
or U10623 (N_10623,N_5809,N_7898);
and U10624 (N_10624,N_5226,N_5524);
or U10625 (N_10625,N_6267,N_5091);
nand U10626 (N_10626,N_5913,N_9308);
nor U10627 (N_10627,N_8241,N_7966);
or U10628 (N_10628,N_7030,N_5266);
and U10629 (N_10629,N_6103,N_9597);
and U10630 (N_10630,N_5742,N_9275);
or U10631 (N_10631,N_6187,N_7374);
or U10632 (N_10632,N_5005,N_8327);
and U10633 (N_10633,N_9721,N_5041);
nor U10634 (N_10634,N_7183,N_9239);
or U10635 (N_10635,N_7602,N_8684);
or U10636 (N_10636,N_8720,N_9967);
and U10637 (N_10637,N_8575,N_7291);
and U10638 (N_10638,N_8456,N_6720);
or U10639 (N_10639,N_6774,N_8134);
or U10640 (N_10640,N_9395,N_5597);
nand U10641 (N_10641,N_5147,N_6614);
xnor U10642 (N_10642,N_7734,N_8591);
nand U10643 (N_10643,N_7311,N_6137);
and U10644 (N_10644,N_7703,N_6544);
nand U10645 (N_10645,N_7748,N_9945);
nor U10646 (N_10646,N_7215,N_9670);
nand U10647 (N_10647,N_7343,N_5578);
nand U10648 (N_10648,N_9920,N_6726);
and U10649 (N_10649,N_8518,N_8510);
or U10650 (N_10650,N_5639,N_9738);
nand U10651 (N_10651,N_5887,N_6177);
xnor U10652 (N_10652,N_9509,N_7087);
nand U10653 (N_10653,N_9617,N_7525);
or U10654 (N_10654,N_6814,N_8276);
nor U10655 (N_10655,N_5984,N_9847);
xnor U10656 (N_10656,N_8274,N_6505);
nor U10657 (N_10657,N_9615,N_9331);
or U10658 (N_10658,N_5237,N_5963);
nor U10659 (N_10659,N_8097,N_9910);
and U10660 (N_10660,N_8142,N_8250);
nand U10661 (N_10661,N_9407,N_9274);
and U10662 (N_10662,N_7957,N_7996);
nand U10663 (N_10663,N_8446,N_7264);
nor U10664 (N_10664,N_7614,N_5588);
nand U10665 (N_10665,N_8272,N_9952);
nand U10666 (N_10666,N_6302,N_8632);
or U10667 (N_10667,N_9616,N_8615);
or U10668 (N_10668,N_5787,N_8503);
and U10669 (N_10669,N_9206,N_6855);
nor U10670 (N_10670,N_8353,N_5291);
xnor U10671 (N_10671,N_5007,N_5939);
nand U10672 (N_10672,N_7144,N_6659);
nor U10673 (N_10673,N_7952,N_7315);
or U10674 (N_10674,N_5788,N_9443);
nor U10675 (N_10675,N_7531,N_8818);
nor U10676 (N_10676,N_9984,N_5013);
or U10677 (N_10677,N_8739,N_8324);
or U10678 (N_10678,N_9094,N_7296);
nor U10679 (N_10679,N_9930,N_9751);
nand U10680 (N_10680,N_7363,N_9690);
and U10681 (N_10681,N_8695,N_7245);
or U10682 (N_10682,N_5914,N_9678);
nand U10683 (N_10683,N_5363,N_8255);
and U10684 (N_10684,N_9476,N_8264);
nand U10685 (N_10685,N_6235,N_8230);
and U10686 (N_10686,N_9725,N_9006);
and U10687 (N_10687,N_6408,N_5465);
nand U10688 (N_10688,N_8764,N_8885);
nor U10689 (N_10689,N_5531,N_5393);
or U10690 (N_10690,N_8691,N_9148);
or U10691 (N_10691,N_7259,N_7899);
nor U10692 (N_10692,N_9122,N_7466);
xor U10693 (N_10693,N_7825,N_6867);
or U10694 (N_10694,N_7535,N_7250);
or U10695 (N_10695,N_8536,N_9343);
nor U10696 (N_10696,N_8886,N_6196);
xor U10697 (N_10697,N_6074,N_7396);
nor U10698 (N_10698,N_9397,N_9039);
xnor U10699 (N_10699,N_7217,N_6935);
and U10700 (N_10700,N_8046,N_9783);
or U10701 (N_10701,N_7918,N_6107);
and U10702 (N_10702,N_9547,N_8898);
nor U10703 (N_10703,N_8642,N_9914);
and U10704 (N_10704,N_5382,N_8468);
or U10705 (N_10705,N_5222,N_9922);
nand U10706 (N_10706,N_6540,N_7537);
and U10707 (N_10707,N_7511,N_8422);
nor U10708 (N_10708,N_6283,N_8703);
or U10709 (N_10709,N_6595,N_5003);
or U10710 (N_10710,N_5573,N_5432);
and U10711 (N_10711,N_7741,N_6084);
and U10712 (N_10712,N_6125,N_6556);
or U10713 (N_10713,N_8861,N_8535);
nor U10714 (N_10714,N_6725,N_8839);
nand U10715 (N_10715,N_8009,N_5006);
or U10716 (N_10716,N_9687,N_9964);
nand U10717 (N_10717,N_9941,N_8904);
nor U10718 (N_10718,N_6593,N_6266);
nor U10719 (N_10719,N_5467,N_5971);
nand U10720 (N_10720,N_5563,N_8667);
nor U10721 (N_10721,N_9703,N_6133);
nor U10722 (N_10722,N_7970,N_9828);
nand U10723 (N_10723,N_7500,N_9188);
xnor U10724 (N_10724,N_9179,N_5646);
nand U10725 (N_10725,N_6167,N_6571);
and U10726 (N_10726,N_9736,N_8035);
and U10727 (N_10727,N_6542,N_5190);
and U10728 (N_10728,N_7742,N_5124);
and U10729 (N_10729,N_6819,N_7162);
or U10730 (N_10730,N_7443,N_9548);
nor U10731 (N_10731,N_6011,N_5107);
or U10732 (N_10732,N_9521,N_6255);
nand U10733 (N_10733,N_5248,N_9244);
and U10734 (N_10734,N_6140,N_9560);
nand U10735 (N_10735,N_9487,N_5263);
nand U10736 (N_10736,N_6714,N_5785);
or U10737 (N_10737,N_7906,N_7113);
nor U10738 (N_10738,N_8495,N_9502);
nor U10739 (N_10739,N_7692,N_8516);
nor U10740 (N_10740,N_7284,N_5058);
or U10741 (N_10741,N_9197,N_6710);
or U10742 (N_10742,N_5655,N_5056);
xor U10743 (N_10743,N_7001,N_9171);
xor U10744 (N_10744,N_9719,N_5808);
and U10745 (N_10745,N_5514,N_9334);
or U10746 (N_10746,N_6037,N_7995);
or U10747 (N_10747,N_8166,N_5686);
xnor U10748 (N_10748,N_7740,N_6548);
and U10749 (N_10749,N_5941,N_8612);
nand U10750 (N_10750,N_7756,N_9737);
nand U10751 (N_10751,N_8334,N_5605);
or U10752 (N_10752,N_6209,N_7381);
or U10753 (N_10753,N_7633,N_9752);
or U10754 (N_10754,N_8143,N_8180);
nand U10755 (N_10755,N_5992,N_9748);
nand U10756 (N_10756,N_6180,N_7901);
xnor U10757 (N_10757,N_6705,N_9298);
or U10758 (N_10758,N_9937,N_9496);
nor U10759 (N_10759,N_9060,N_5352);
nand U10760 (N_10760,N_8637,N_8646);
nand U10761 (N_10761,N_8413,N_7625);
and U10762 (N_10762,N_7964,N_8464);
and U10763 (N_10763,N_7317,N_6262);
or U10764 (N_10764,N_9380,N_6962);
nor U10765 (N_10765,N_7767,N_6024);
or U10766 (N_10766,N_5794,N_9074);
xor U10767 (N_10767,N_9075,N_8654);
and U10768 (N_10768,N_7882,N_9948);
and U10769 (N_10769,N_8418,N_9217);
or U10770 (N_10770,N_9119,N_6870);
and U10771 (N_10771,N_8428,N_7308);
and U10772 (N_10772,N_5273,N_7490);
nand U10773 (N_10773,N_5903,N_5884);
or U10774 (N_10774,N_7003,N_5454);
nand U10775 (N_10775,N_6019,N_7450);
and U10776 (N_10776,N_7057,N_6480);
or U10777 (N_10777,N_5373,N_5264);
xor U10778 (N_10778,N_9773,N_6093);
or U10779 (N_10779,N_9488,N_9357);
nor U10780 (N_10780,N_5411,N_7434);
and U10781 (N_10781,N_5552,N_9080);
nand U10782 (N_10782,N_7373,N_9050);
and U10783 (N_10783,N_8251,N_8774);
xor U10784 (N_10784,N_7101,N_5378);
nand U10785 (N_10785,N_7743,N_8090);
nand U10786 (N_10786,N_8515,N_9778);
xnor U10787 (N_10787,N_7561,N_7248);
nor U10788 (N_10788,N_8045,N_5904);
nor U10789 (N_10789,N_5656,N_8227);
nor U10790 (N_10790,N_9570,N_7849);
or U10791 (N_10791,N_7519,N_5694);
or U10792 (N_10792,N_9333,N_9841);
or U10793 (N_10793,N_8932,N_7858);
nand U10794 (N_10794,N_6885,N_5151);
nor U10795 (N_10795,N_7758,N_5882);
nor U10796 (N_10796,N_8531,N_9656);
nand U10797 (N_10797,N_6738,N_5476);
xor U10798 (N_10798,N_8599,N_9645);
nor U10799 (N_10799,N_5481,N_6282);
xor U10800 (N_10800,N_5584,N_5512);
and U10801 (N_10801,N_5762,N_8870);
nand U10802 (N_10802,N_5698,N_6498);
nor U10803 (N_10803,N_9727,N_9935);
or U10804 (N_10804,N_9399,N_5770);
xnor U10805 (N_10805,N_9987,N_5200);
nand U10806 (N_10806,N_6565,N_6813);
nor U10807 (N_10807,N_7318,N_8442);
or U10808 (N_10808,N_9105,N_9405);
or U10809 (N_10809,N_5826,N_6146);
or U10810 (N_10810,N_5251,N_9297);
nand U10811 (N_10811,N_6754,N_5747);
xnor U10812 (N_10812,N_6933,N_7760);
and U10813 (N_10813,N_8249,N_9588);
xor U10814 (N_10814,N_8372,N_6386);
xnor U10815 (N_10815,N_8486,N_7967);
nor U10816 (N_10816,N_8414,N_9330);
nand U10817 (N_10817,N_6588,N_7402);
nand U10818 (N_10818,N_7550,N_6365);
and U10819 (N_10819,N_6109,N_5194);
nand U10820 (N_10820,N_5106,N_9788);
nor U10821 (N_10821,N_5863,N_6678);
or U10822 (N_10822,N_9902,N_9456);
xor U10823 (N_10823,N_6645,N_6642);
or U10824 (N_10824,N_5983,N_7611);
or U10825 (N_10825,N_7329,N_8088);
and U10826 (N_10826,N_8977,N_5271);
xor U10827 (N_10827,N_9776,N_8560);
and U10828 (N_10828,N_7572,N_7810);
nor U10829 (N_10829,N_7865,N_9843);
and U10830 (N_10830,N_6748,N_5774);
nand U10831 (N_10831,N_7185,N_7231);
or U10832 (N_10832,N_5016,N_7842);
and U10833 (N_10833,N_9608,N_7242);
nor U10834 (N_10834,N_7015,N_6831);
and U10835 (N_10835,N_8141,N_6344);
and U10836 (N_10836,N_8826,N_8721);
or U10837 (N_10837,N_8728,N_7848);
and U10838 (N_10838,N_5825,N_5504);
or U10839 (N_10839,N_5848,N_6630);
and U10840 (N_10840,N_9826,N_5631);
nand U10841 (N_10841,N_9522,N_7713);
or U10842 (N_10842,N_8790,N_9042);
nor U10843 (N_10843,N_5812,N_6322);
nand U10844 (N_10844,N_5267,N_8028);
nand U10845 (N_10845,N_8848,N_8675);
nand U10846 (N_10846,N_8121,N_9889);
nor U10847 (N_10847,N_8952,N_6509);
nand U10848 (N_10848,N_5277,N_8415);
nand U10849 (N_10849,N_9041,N_6257);
and U10850 (N_10850,N_5528,N_9970);
nor U10851 (N_10851,N_9375,N_7596);
nand U10852 (N_10852,N_6974,N_7624);
nor U10853 (N_10853,N_8084,N_8344);
and U10854 (N_10854,N_8500,N_5255);
nand U10855 (N_10855,N_6127,N_6771);
nor U10856 (N_10856,N_8751,N_9342);
xor U10857 (N_10857,N_5052,N_6563);
or U10858 (N_10858,N_9223,N_8708);
xnor U10859 (N_10859,N_8326,N_6463);
nor U10860 (N_10860,N_6478,N_7260);
xor U10861 (N_10861,N_5022,N_5287);
and U10862 (N_10862,N_9390,N_7206);
or U10863 (N_10863,N_8659,N_5748);
and U10864 (N_10864,N_6334,N_7885);
nor U10865 (N_10865,N_7803,N_7902);
nor U10866 (N_10866,N_9097,N_7577);
and U10867 (N_10867,N_9991,N_8095);
and U10868 (N_10868,N_6834,N_8732);
nor U10869 (N_10869,N_9240,N_7844);
or U10870 (N_10870,N_5933,N_8601);
nand U10871 (N_10871,N_9120,N_5012);
or U10872 (N_10872,N_7548,N_5215);
and U10873 (N_10873,N_5927,N_5383);
or U10874 (N_10874,N_6009,N_8015);
nor U10875 (N_10875,N_9526,N_6433);
or U10876 (N_10876,N_7353,N_8577);
xor U10877 (N_10877,N_9098,N_5500);
nor U10878 (N_10878,N_5901,N_5804);
nor U10879 (N_10879,N_5923,N_8884);
or U10880 (N_10880,N_7745,N_5478);
nor U10881 (N_10881,N_9990,N_5918);
nor U10882 (N_10882,N_5491,N_5521);
nor U10883 (N_10883,N_5850,N_5912);
nand U10884 (N_10884,N_5772,N_5346);
or U10885 (N_10885,N_8611,N_6421);
and U10886 (N_10886,N_9972,N_7052);
nand U10887 (N_10887,N_5532,N_8385);
or U10888 (N_10888,N_8242,N_8588);
or U10889 (N_10889,N_9198,N_7833);
nand U10890 (N_10890,N_6077,N_6179);
nor U10891 (N_10891,N_5764,N_5189);
xor U10892 (N_10892,N_9470,N_8750);
nor U10893 (N_10893,N_7356,N_6477);
or U10894 (N_10894,N_9210,N_6954);
xnor U10895 (N_10895,N_8791,N_7759);
nand U10896 (N_10896,N_7426,N_8915);
nor U10897 (N_10897,N_6238,N_8496);
or U10898 (N_10898,N_8733,N_9215);
nor U10899 (N_10899,N_6163,N_8971);
nor U10900 (N_10900,N_8172,N_5253);
nor U10901 (N_10901,N_7024,N_9460);
nand U10902 (N_10902,N_5216,N_6635);
xnor U10903 (N_10903,N_7491,N_6398);
xnor U10904 (N_10904,N_7755,N_5811);
nor U10905 (N_10905,N_5827,N_8102);
nand U10906 (N_10906,N_6577,N_7149);
or U10907 (N_10907,N_6924,N_6014);
nand U10908 (N_10908,N_5658,N_8854);
and U10909 (N_10909,N_6489,N_6576);
or U10910 (N_10910,N_7982,N_9475);
nor U10911 (N_10911,N_6223,N_6702);
nand U10912 (N_10912,N_8523,N_6722);
nor U10913 (N_10913,N_7591,N_5119);
or U10914 (N_10914,N_7056,N_9164);
nor U10915 (N_10915,N_9058,N_8336);
and U10916 (N_10916,N_6534,N_6105);
or U10917 (N_10917,N_5871,N_5700);
or U10918 (N_10918,N_6782,N_5019);
nand U10919 (N_10919,N_9669,N_5328);
nand U10920 (N_10920,N_6669,N_7139);
and U10921 (N_10921,N_9648,N_7693);
nand U10922 (N_10922,N_7171,N_5609);
or U10923 (N_10923,N_5188,N_7361);
nor U10924 (N_10924,N_7931,N_8485);
nor U10925 (N_10925,N_9983,N_8175);
xor U10926 (N_10926,N_6656,N_7838);
and U10927 (N_10927,N_6545,N_6596);
or U10928 (N_10928,N_7339,N_6560);
nand U10929 (N_10929,N_9890,N_8083);
nor U10930 (N_10930,N_6020,N_7665);
and U10931 (N_10931,N_6585,N_7961);
nand U10932 (N_10932,N_6503,N_9896);
or U10933 (N_10933,N_6485,N_5657);
nor U10934 (N_10934,N_7050,N_5412);
nand U10935 (N_10935,N_9257,N_8662);
nor U10936 (N_10936,N_9377,N_6240);
and U10937 (N_10937,N_9556,N_9905);
or U10938 (N_10938,N_7427,N_7841);
nor U10939 (N_10939,N_9601,N_7715);
nand U10940 (N_10940,N_7517,N_5301);
nand U10941 (N_10941,N_8377,N_5626);
nand U10942 (N_10942,N_9611,N_9020);
and U10943 (N_10943,N_6340,N_9116);
nor U10944 (N_10944,N_5560,N_5161);
nand U10945 (N_10945,N_5033,N_5489);
xnor U10946 (N_10946,N_8799,N_9155);
nand U10947 (N_10947,N_8544,N_6946);
or U10948 (N_10948,N_7917,N_5397);
nor U10949 (N_10949,N_9409,N_7189);
nor U10950 (N_10950,N_6251,N_5511);
nand U10951 (N_10951,N_8741,N_9503);
or U10952 (N_10952,N_8773,N_8705);
nor U10953 (N_10953,N_5717,N_8661);
nor U10954 (N_10954,N_6392,N_5027);
nor U10955 (N_10955,N_9884,N_7565);
nand U10956 (N_10956,N_5784,N_6559);
or U10957 (N_10957,N_5176,N_5789);
or U10958 (N_10958,N_9507,N_9195);
or U10959 (N_10959,N_6268,N_6015);
and U10960 (N_10960,N_6265,N_5815);
nand U10961 (N_10961,N_9921,N_9520);
and U10962 (N_10962,N_8472,N_9501);
nor U10963 (N_10963,N_9514,N_9167);
xnor U10964 (N_10964,N_7547,N_9771);
or U10965 (N_10965,N_5304,N_6874);
nand U10966 (N_10966,N_9482,N_6136);
xor U10967 (N_10967,N_7607,N_8976);
nor U10968 (N_10968,N_7064,N_7042);
nor U10969 (N_10969,N_6202,N_6985);
and U10970 (N_10970,N_8618,N_7986);
and U10971 (N_10971,N_7501,N_5293);
and U10972 (N_10972,N_7630,N_7827);
nand U10973 (N_10973,N_8777,N_9643);
or U10974 (N_10974,N_6667,N_5071);
nor U10975 (N_10975,N_7621,N_9825);
and U10976 (N_10976,N_5351,N_5507);
nand U10977 (N_10977,N_5473,N_9550);
xor U10978 (N_10978,N_7670,N_9189);
nor U10979 (N_10979,N_9862,N_5408);
and U10980 (N_10980,N_8710,N_5355);
nand U10981 (N_10981,N_5911,N_8213);
nor U10982 (N_10982,N_7822,N_8018);
and U10983 (N_10983,N_8614,N_8047);
nand U10984 (N_10984,N_7061,N_8107);
and U10985 (N_10985,N_9953,N_5117);
or U10986 (N_10986,N_7770,N_8766);
nand U10987 (N_10987,N_8150,N_5706);
nand U10988 (N_10988,N_8919,N_5969);
nor U10989 (N_10989,N_9529,N_9536);
nor U10990 (N_10990,N_7784,N_5854);
or U10991 (N_10991,N_9177,N_9354);
or U10992 (N_10992,N_7509,N_6940);
and U10993 (N_10993,N_5936,N_7044);
and U10994 (N_10994,N_5361,N_5078);
or U10995 (N_10995,N_5477,N_7538);
nor U10996 (N_10996,N_5641,N_6123);
nor U10997 (N_10997,N_5098,N_7400);
or U10998 (N_10998,N_5749,N_7272);
nor U10999 (N_10999,N_9892,N_9966);
or U11000 (N_11000,N_8687,N_8749);
or U11001 (N_11001,N_6425,N_7238);
and U11002 (N_11002,N_6193,N_7088);
or U11003 (N_11003,N_5130,N_6797);
or U11004 (N_11004,N_9428,N_9439);
nand U11005 (N_11005,N_8775,N_6331);
and U11006 (N_11006,N_9306,N_5630);
and U11007 (N_11007,N_8899,N_6519);
and U11008 (N_11008,N_8306,N_7276);
nand U11009 (N_11009,N_5100,N_5775);
xnor U11010 (N_11010,N_9326,N_9370);
or U11011 (N_11011,N_5892,N_8387);
nand U11012 (N_11012,N_7792,N_8024);
nand U11013 (N_11013,N_5141,N_6882);
or U11014 (N_11014,N_7530,N_7229);
nand U11015 (N_11015,N_6961,N_7159);
xor U11016 (N_11016,N_6164,N_7988);
xor U11017 (N_11017,N_8158,N_9053);
nor U11018 (N_11018,N_5554,N_6792);
and U11019 (N_11019,N_9288,N_6884);
nor U11020 (N_11020,N_8434,N_8494);
nor U11021 (N_11021,N_7772,N_9054);
nand U11022 (N_11022,N_7930,N_9762);
or U11023 (N_11023,N_7889,N_9403);
nor U11024 (N_11024,N_6902,N_9887);
nand U11025 (N_11025,N_7282,N_8935);
xor U11026 (N_11026,N_7105,N_7442);
and U11027 (N_11027,N_6170,N_9289);
or U11028 (N_11028,N_6789,N_8934);
and U11029 (N_11029,N_6384,N_7100);
and U11030 (N_11030,N_6646,N_7508);
or U11031 (N_11031,N_7131,N_5484);
and U11032 (N_11032,N_8525,N_9637);
nor U11033 (N_11033,N_7718,N_5135);
xor U11034 (N_11034,N_5174,N_9440);
nand U11035 (N_11035,N_5199,N_7040);
and U11036 (N_11036,N_5144,N_7649);
or U11037 (N_11037,N_8454,N_9337);
or U11038 (N_11038,N_8582,N_7109);
nand U11039 (N_11039,N_6971,N_6272);
xnor U11040 (N_11040,N_7867,N_8460);
and U11041 (N_11041,N_9284,N_7639);
nor U11042 (N_11042,N_5506,N_6057);
or U11043 (N_11043,N_9445,N_8247);
nand U11044 (N_11044,N_8295,N_9938);
xor U11045 (N_11045,N_7804,N_8847);
or U11046 (N_11046,N_5640,N_7376);
or U11047 (N_11047,N_6324,N_5837);
nand U11048 (N_11048,N_5535,N_9712);
nor U11049 (N_11049,N_5534,N_9303);
nand U11050 (N_11050,N_7610,N_7592);
nand U11051 (N_11051,N_6460,N_5404);
and U11052 (N_11052,N_5252,N_6801);
and U11053 (N_11053,N_6279,N_8202);
nor U11054 (N_11054,N_5244,N_6706);
nor U11055 (N_11055,N_7210,N_9928);
nand U11056 (N_11056,N_9524,N_6504);
and U11057 (N_11057,N_7757,N_8840);
or U11058 (N_11058,N_5710,N_8822);
or U11059 (N_11059,N_8927,N_8913);
and U11060 (N_11060,N_6174,N_5525);
or U11061 (N_11061,N_5831,N_8300);
and U11062 (N_11062,N_8165,N_5667);
nor U11063 (N_11063,N_6875,N_5973);
xor U11064 (N_11064,N_8702,N_6793);
and U11065 (N_11065,N_6045,N_7791);
nand U11066 (N_11066,N_7182,N_5421);
and U11067 (N_11067,N_6220,N_9632);
or U11068 (N_11068,N_6976,N_6633);
and U11069 (N_11069,N_8410,N_6029);
or U11070 (N_11070,N_9885,N_5589);
or U11071 (N_11071,N_9313,N_6906);
nor U11072 (N_11072,N_7141,N_5523);
nor U11073 (N_11073,N_5548,N_6300);
nand U11074 (N_11074,N_9696,N_8803);
nand U11075 (N_11075,N_6718,N_8475);
nand U11076 (N_11076,N_5683,N_8129);
or U11077 (N_11077,N_9389,N_8881);
nor U11078 (N_11078,N_7468,N_9593);
nand U11079 (N_11079,N_6753,N_8909);
and U11080 (N_11080,N_7268,N_5482);
or U11081 (N_11081,N_9874,N_9213);
or U11082 (N_11082,N_6511,N_6134);
or U11083 (N_11083,N_7523,N_9247);
or U11084 (N_11084,N_9355,N_7691);
or U11085 (N_11085,N_6376,N_6173);
xor U11086 (N_11086,N_8765,N_5822);
nor U11087 (N_11087,N_5729,N_7807);
nor U11088 (N_11088,N_8754,N_8520);
nor U11089 (N_11089,N_5712,N_5339);
or U11090 (N_11090,N_6547,N_7855);
nor U11091 (N_11091,N_8900,N_6741);
and U11092 (N_11092,N_9176,N_5095);
nor U11093 (N_11093,N_5466,N_7439);
or U11094 (N_11094,N_8396,N_5394);
nand U11095 (N_11095,N_7204,N_6473);
nand U11096 (N_11096,N_7985,N_5607);
and U11097 (N_11097,N_5541,N_8644);
xor U11098 (N_11098,N_8597,N_7429);
and U11099 (N_11099,N_5737,N_9723);
xnor U11100 (N_11100,N_8154,N_6900);
xor U11101 (N_11101,N_6495,N_5475);
and U11102 (N_11102,N_9369,N_6117);
and U11103 (N_11103,N_6983,N_5898);
nand U11104 (N_11104,N_9418,N_5492);
nor U11105 (N_11105,N_6947,N_7067);
nand U11106 (N_11106,N_5359,N_5031);
nor U11107 (N_11107,N_8157,N_9803);
nand U11108 (N_11108,N_8488,N_8641);
or U11109 (N_11109,N_7175,N_5797);
and U11110 (N_11110,N_5878,N_8389);
or U11111 (N_11111,N_9974,N_7033);
nor U11112 (N_11112,N_8592,N_7814);
nand U11113 (N_11113,N_6636,N_6162);
nor U11114 (N_11114,N_6010,N_7619);
nor U11115 (N_11115,N_6941,N_5814);
nand U11116 (N_11116,N_7877,N_7720);
xnor U11117 (N_11117,N_8921,N_8963);
nand U11118 (N_11118,N_7393,N_8841);
nand U11119 (N_11119,N_8333,N_6151);
or U11120 (N_11120,N_6178,N_6873);
or U11121 (N_11121,N_9517,N_7912);
nand U11122 (N_11122,N_7579,N_6114);
xor U11123 (N_11123,N_5437,N_7301);
nor U11124 (N_11124,N_8050,N_8665);
or U11125 (N_11125,N_7007,N_6963);
nor U11126 (N_11126,N_6914,N_6195);
nand U11127 (N_11127,N_5773,N_7534);
nor U11128 (N_11128,N_5457,N_6708);
nor U11129 (N_11129,N_6750,N_5665);
nor U11130 (N_11130,N_8674,N_5126);
nor U11131 (N_11131,N_7196,N_8194);
nand U11132 (N_11132,N_9880,N_7129);
nor U11133 (N_11133,N_5839,N_5061);
or U11134 (N_11134,N_6603,N_5115);
or U11135 (N_11135,N_7998,N_9262);
and U11136 (N_11136,N_9891,N_9603);
nand U11137 (N_11137,N_8407,N_6619);
xnor U11138 (N_11138,N_9674,N_8416);
or U11139 (N_11139,N_6978,N_6899);
nand U11140 (N_11140,N_7776,N_5325);
nand U11141 (N_11141,N_7681,N_8497);
nand U11142 (N_11142,N_8253,N_9801);
nor U11143 (N_11143,N_9883,N_5358);
nor U11144 (N_11144,N_8453,N_9218);
or U11145 (N_11145,N_6663,N_8858);
and U11146 (N_11146,N_8990,N_9286);
or U11147 (N_11147,N_6943,N_8723);
nand U11148 (N_11148,N_7425,N_6397);
or U11149 (N_11149,N_5110,N_7881);
nor U11150 (N_11150,N_5961,N_8823);
and U11151 (N_11151,N_5218,N_9174);
nor U11152 (N_11152,N_8010,N_6383);
or U11153 (N_11153,N_5782,N_8929);
or U11154 (N_11154,N_7286,N_5537);
xnor U11155 (N_11155,N_9477,N_6541);
or U11156 (N_11156,N_9273,N_5557);
nand U11157 (N_11157,N_5185,N_8104);
and U11158 (N_11158,N_6795,N_8279);
or U11159 (N_11159,N_7837,N_8943);
xnor U11160 (N_11160,N_6573,N_9726);
xnor U11161 (N_11161,N_8188,N_8354);
nand U11162 (N_11162,N_7620,N_9906);
or U11163 (N_11163,N_5395,N_5433);
or U11164 (N_11164,N_5590,N_6715);
nor U11165 (N_11165,N_8694,N_8567);
or U11166 (N_11166,N_8022,N_6075);
or U11167 (N_11167,N_9412,N_7992);
nor U11168 (N_11168,N_8319,N_8960);
or U11169 (N_11169,N_6273,N_7585);
and U11170 (N_11170,N_8052,N_7650);
and U11171 (N_11171,N_6913,N_7907);
or U11172 (N_11172,N_5843,N_5763);
and U11173 (N_11173,N_9673,N_9899);
or U11174 (N_11174,N_8629,N_8471);
and U11175 (N_11175,N_8014,N_8091);
and U11176 (N_11176,N_8556,N_6461);
and U11177 (N_11177,N_8245,N_5419);
nand U11178 (N_11178,N_6858,N_9018);
nor U11179 (N_11179,N_5614,N_8717);
nor U11180 (N_11180,N_7895,N_8092);
and U11181 (N_11181,N_8722,N_7563);
xor U11182 (N_11182,N_7472,N_7150);
or U11183 (N_11183,N_7452,N_9338);
nor U11184 (N_11184,N_7761,N_6432);
nand U11185 (N_11185,N_6102,N_8320);
or U11186 (N_11186,N_5406,N_7459);
nand U11187 (N_11187,N_6215,N_7751);
nor U11188 (N_11188,N_7239,N_8040);
nand U11189 (N_11189,N_7513,N_9998);
nand U11190 (N_11190,N_5816,N_5204);
and U11191 (N_11191,N_9464,N_5728);
nor U11192 (N_11192,N_7915,N_6651);
nand U11193 (N_11193,N_5306,N_5870);
or U11194 (N_11194,N_9111,N_8163);
nor U11195 (N_11195,N_5780,N_9323);
nand U11196 (N_11196,N_9455,N_6594);
and U11197 (N_11197,N_6597,N_5940);
nand U11198 (N_11198,N_9912,N_5627);
nand U11199 (N_11199,N_6586,N_7090);
and U11200 (N_11200,N_5945,N_8678);
or U11201 (N_11201,N_5875,N_5055);
nand U11202 (N_11202,N_5329,N_9364);
nand U11203 (N_11203,N_7532,N_5709);
xor U11204 (N_11204,N_9019,N_6472);
or U11205 (N_11205,N_9733,N_8743);
xor U11206 (N_11206,N_7735,N_6307);
and U11207 (N_11207,N_5201,N_8789);
nor U11208 (N_11208,N_5823,N_9299);
xnor U11209 (N_11209,N_8716,N_6692);
nor U11210 (N_11210,N_8655,N_6234);
nand U11211 (N_11211,N_9359,N_7048);
nor U11212 (N_11212,N_8119,N_5572);
or U11213 (N_11213,N_6090,N_8949);
nand U11214 (N_11214,N_6030,N_7273);
xor U11215 (N_11215,N_7167,N_5608);
and U11216 (N_11216,N_8273,N_7020);
xnor U11217 (N_11217,N_5116,N_5191);
nand U11218 (N_11218,N_8409,N_7518);
and U11219 (N_11219,N_7258,N_9072);
nand U11220 (N_11220,N_5459,N_6610);
and U11221 (N_11221,N_9749,N_9867);
or U11222 (N_11222,N_8616,N_8467);
nor U11223 (N_11223,N_8690,N_7820);
xor U11224 (N_11224,N_7257,N_7172);
xnor U11225 (N_11225,N_6823,N_7256);
or U11226 (N_11226,N_6836,N_5576);
or U11227 (N_11227,N_9821,N_6516);
and U11228 (N_11228,N_8895,N_6431);
and U11229 (N_11229,N_5866,N_7471);
and U11230 (N_11230,N_8288,N_9253);
or U11231 (N_11231,N_5060,N_7684);
nand U11232 (N_11232,N_8501,N_8470);
nand U11233 (N_11233,N_5059,N_8664);
nor U11234 (N_11234,N_9486,N_9319);
nand U11235 (N_11235,N_9995,N_6956);
and U11236 (N_11236,N_7664,N_7469);
nand U11237 (N_11237,N_7072,N_9784);
or U11238 (N_11238,N_6321,N_8639);
or U11239 (N_11239,N_8879,N_8688);
nand U11240 (N_11240,N_6749,N_9471);
xor U11241 (N_11241,N_6144,N_6261);
nor U11242 (N_11242,N_8816,N_5985);
nor U11243 (N_11243,N_5726,N_7328);
or U11244 (N_11244,N_5407,N_7823);
xnor U11245 (N_11245,N_8423,N_7847);
and U11246 (N_11246,N_9697,N_6524);
nand U11247 (N_11247,N_5881,N_9584);
xor U11248 (N_11248,N_8345,N_7799);
xnor U11249 (N_11249,N_9954,N_8569);
xor U11250 (N_11250,N_8323,N_8634);
or U11251 (N_11251,N_9518,N_5543);
xnor U11252 (N_11252,N_8894,N_8056);
nor U11253 (N_11253,N_8115,N_9580);
or U11254 (N_11254,N_9076,N_7617);
nor U11255 (N_11255,N_5905,N_6860);
nand U11256 (N_11256,N_5948,N_7522);
xor U11257 (N_11257,N_7839,N_6304);
nor U11258 (N_11258,N_9527,N_8903);
nand U11259 (N_11259,N_9499,N_9859);
or U11260 (N_11260,N_7653,N_8737);
nor U11261 (N_11261,N_7447,N_6785);
nand U11262 (N_11262,N_6973,N_7195);
or U11263 (N_11263,N_8411,N_7476);
nand U11264 (N_11264,N_7492,N_9813);
or U11265 (N_11265,N_7474,N_9068);
and U11266 (N_11266,N_7482,N_8887);
nand U11267 (N_11267,N_9573,N_6467);
nor U11268 (N_11268,N_6097,N_7146);
nand U11269 (N_11269,N_8817,N_5795);
and U11270 (N_11270,N_8185,N_5879);
and U11271 (N_11271,N_5732,N_8530);
xor U11272 (N_11272,N_6079,N_8673);
nor U11273 (N_11273,N_5691,N_8033);
xor U11274 (N_11274,N_8872,N_6338);
and U11275 (N_11275,N_9067,N_6953);
nor U11276 (N_11276,N_9381,N_8164);
and U11277 (N_11277,N_9619,N_5460);
or U11278 (N_11278,N_6299,N_9671);
nand U11279 (N_11279,N_6763,N_7937);
xnor U11280 (N_11280,N_9278,N_6185);
and U11281 (N_11281,N_6153,N_8512);
xnor U11282 (N_11282,N_5937,N_7824);
or U11283 (N_11283,N_7448,N_6878);
nor U11284 (N_11284,N_5902,N_8793);
or U11285 (N_11285,N_6381,N_6631);
xnor U11286 (N_11286,N_7094,N_8235);
and U11287 (N_11287,N_5830,N_8063);
xor U11288 (N_11288,N_6517,N_7275);
or U11289 (N_11289,N_6159,N_7424);
or U11290 (N_11290,N_9073,N_6522);
and U11291 (N_11291,N_5832,N_9295);
or U11292 (N_11292,N_6696,N_7254);
or U11293 (N_11293,N_5164,N_8174);
or U11294 (N_11294,N_9133,N_9466);
and U11295 (N_11295,N_8576,N_8677);
and U11296 (N_11296,N_8315,N_7358);
and U11297 (N_11297,N_7817,N_9554);
nor U11298 (N_11298,N_9628,N_8451);
nand U11299 (N_11299,N_9647,N_6100);
and U11300 (N_11300,N_5396,N_8187);
nand U11301 (N_11301,N_6171,N_6081);
and U11302 (N_11302,N_8696,N_8953);
or U11303 (N_11303,N_5958,N_8504);
nand U11304 (N_11304,N_9043,N_8066);
or U11305 (N_11305,N_7456,N_9252);
nor U11306 (N_11306,N_8693,N_9483);
nor U11307 (N_11307,N_9606,N_9187);
or U11308 (N_11308,N_5736,N_8399);
nor U11309 (N_11309,N_6468,N_5663);
and U11310 (N_11310,N_6989,N_7663);
or U11311 (N_11311,N_9735,N_7798);
nor U11312 (N_11312,N_8439,N_6201);
and U11313 (N_11313,N_5038,N_6181);
or U11314 (N_11314,N_9281,N_7486);
xor U11315 (N_11315,N_6033,N_7569);
or U11316 (N_11316,N_5214,N_6183);
or U11317 (N_11317,N_6671,N_6551);
nand U11318 (N_11318,N_8533,N_5332);
nand U11319 (N_11319,N_7480,N_7115);
or U11320 (N_11320,N_6670,N_6207);
nand U11321 (N_11321,N_5132,N_8742);
nand U11322 (N_11322,N_9011,N_9806);
nand U11323 (N_11323,N_5386,N_8752);
and U11324 (N_11324,N_5405,N_5702);
xnor U11325 (N_11325,N_7991,N_9620);
nand U11326 (N_11326,N_7732,N_8481);
or U11327 (N_11327,N_8804,N_9701);
and U11328 (N_11328,N_5103,N_6343);
or U11329 (N_11329,N_6768,N_8007);
or U11330 (N_11330,N_5451,N_8837);
or U11331 (N_11331,N_5883,N_6244);
and U11332 (N_11332,N_6129,N_6270);
xnor U11333 (N_11333,N_7483,N_9004);
nor U11334 (N_11334,N_7211,N_5705);
and U11335 (N_11335,N_5349,N_5651);
nor U11336 (N_11336,N_6441,N_9368);
nand U11337 (N_11337,N_7290,N_8053);
nor U11338 (N_11338,N_7938,N_6106);
nor U11339 (N_11339,N_8124,N_8825);
xnor U11340 (N_11340,N_7811,N_9336);
or U11341 (N_11341,N_7616,N_7634);
and U11342 (N_11342,N_6399,N_7411);
or U11343 (N_11343,N_5909,N_5262);
nand U11344 (N_11344,N_8330,N_8585);
nor U11345 (N_11345,N_6025,N_6328);
nand U11346 (N_11346,N_8123,N_9061);
nand U11347 (N_11347,N_9706,N_6747);
nand U11348 (N_11348,N_8701,N_7126);
nor U11349 (N_11349,N_8003,N_7949);
nor U11350 (N_11350,N_7421,N_5148);
nand U11351 (N_11351,N_5233,N_7414);
nand U11352 (N_11352,N_6241,N_8683);
or U11353 (N_11353,N_9372,N_9512);
nor U11354 (N_11354,N_7348,N_8062);
or U11355 (N_11355,N_9739,N_9462);
nand U11356 (N_11356,N_9949,N_5908);
and U11357 (N_11357,N_9768,N_5368);
nor U11358 (N_11358,N_6046,N_5081);
and U11359 (N_11359,N_6526,N_7543);
nor U11360 (N_11360,N_7613,N_8201);
nand U11361 (N_11361,N_8210,N_9789);
and U11362 (N_11362,N_6385,N_7724);
or U11363 (N_11363,N_5125,N_5026);
and U11364 (N_11364,N_6085,N_7680);
nor U11365 (N_11365,N_8362,N_5249);
nand U11366 (N_11366,N_9581,N_5247);
or U11367 (N_11367,N_9077,N_9714);
nor U11368 (N_11368,N_9858,N_9207);
nor U11369 (N_11369,N_6740,N_8890);
nand U11370 (N_11370,N_9504,N_6326);
nor U11371 (N_11371,N_9819,N_7662);
nor U11372 (N_11372,N_6291,N_7236);
nand U11373 (N_11373,N_6921,N_6697);
or U11374 (N_11374,N_6579,N_8528);
nand U11375 (N_11375,N_8462,N_9258);
and U11376 (N_11376,N_9125,N_7417);
and U11377 (N_11377,N_9568,N_5585);
and U11378 (N_11378,N_6395,N_6188);
or U11379 (N_11379,N_7407,N_8609);
nand U11380 (N_11380,N_8358,N_7142);
and U11381 (N_11381,N_7043,N_5000);
or U11382 (N_11382,N_6807,N_6689);
or U11383 (N_11383,N_6992,N_9318);
and U11384 (N_11384,N_5679,N_9515);
or U11385 (N_11385,N_6021,N_6124);
nand U11386 (N_11386,N_8125,N_9746);
nor U11387 (N_11387,N_9312,N_5946);
and U11388 (N_11388,N_7812,N_9612);
nor U11389 (N_11389,N_6323,N_8425);
nor U11390 (N_11390,N_6154,N_6698);
nand U11391 (N_11391,N_7626,N_5842);
nand U11392 (N_11392,N_7344,N_9490);
and U11393 (N_11393,N_7934,N_6998);
nor U11394 (N_11394,N_6497,N_5136);
and U11395 (N_11395,N_8573,N_8828);
nand U11396 (N_11396,N_9144,N_6672);
and U11397 (N_11397,N_9203,N_8600);
nand U11398 (N_11398,N_6893,N_5965);
nand U11399 (N_11399,N_5139,N_9106);
or U11400 (N_11400,N_9327,N_8676);
and U11401 (N_11401,N_9250,N_8513);
and U11402 (N_11402,N_8814,N_6484);
or U11403 (N_11403,N_9681,N_9193);
or U11404 (N_11404,N_7909,N_5367);
nor U11405 (N_11405,N_7657,N_9351);
or U11406 (N_11406,N_5987,N_8744);
or U11407 (N_11407,N_8365,N_8031);
nor U11408 (N_11408,N_7244,N_9975);
or U11409 (N_11409,N_9082,N_5802);
or U11410 (N_11410,N_7826,N_8554);
xnor U11411 (N_11411,N_7672,N_7944);
or U11412 (N_11412,N_8603,N_8792);
xnor U11413 (N_11413,N_5420,N_9404);
nor U11414 (N_11414,N_7834,N_8224);
or U11415 (N_11415,N_8734,N_8833);
nand U11416 (N_11416,N_7710,N_9398);
xor U11417 (N_11417,N_9711,N_8266);
and U11418 (N_11418,N_7346,N_7919);
or U11419 (N_11419,N_8731,N_8863);
or U11420 (N_11420,N_8581,N_7753);
or U11421 (N_11421,N_6848,N_8815);
or U11422 (N_11422,N_5087,N_8133);
and U11423 (N_11423,N_6574,N_9630);
and U11424 (N_11424,N_5574,N_6237);
and U11425 (N_11425,N_9379,N_9202);
and U11426 (N_11426,N_6687,N_8876);
or U11427 (N_11427,N_5580,N_7107);
or U11428 (N_11428,N_6306,N_5449);
and U11429 (N_11429,N_6703,N_7997);
xnor U11430 (N_11430,N_6211,N_7940);
nand U11431 (N_11431,N_6113,N_9335);
nand U11432 (N_11432,N_6693,N_9587);
and U11433 (N_11433,N_9792,N_8437);
nand U11434 (N_11434,N_5501,N_8231);
and U11435 (N_11435,N_6507,N_9599);
nand U11436 (N_11436,N_5735,N_7843);
or U11437 (N_11437,N_5275,N_8002);
nor U11438 (N_11438,N_6250,N_6809);
xnor U11439 (N_11439,N_7280,N_7866);
nand U11440 (N_11440,N_6847,N_8193);
or U11441 (N_11441,N_5979,N_9276);
and U11442 (N_11442,N_9759,N_9481);
nor U11443 (N_11443,N_8369,N_8038);
xnor U11444 (N_11444,N_9916,N_8645);
nor U11445 (N_11445,N_5818,N_9154);
and U11446 (N_11446,N_9936,N_6824);
nand U11447 (N_11447,N_6228,N_9110);
and U11448 (N_11448,N_6126,N_7980);
nand U11449 (N_11449,N_8232,N_8707);
or U11450 (N_11450,N_6078,N_7872);
and U11451 (N_11451,N_8131,N_9744);
nand U11452 (N_11452,N_6414,N_6788);
and U11453 (N_11453,N_6032,N_9943);
or U11454 (N_11454,N_5417,N_7123);
or U11455 (N_11455,N_5820,N_9266);
nor U11456 (N_11456,N_7864,N_6054);
nor U11457 (N_11457,N_7059,N_7475);
nand U11458 (N_11458,N_5874,N_8643);
and U11459 (N_11459,N_8874,N_9152);
xnor U11460 (N_11460,N_7341,N_9956);
or U11461 (N_11461,N_5648,N_9682);
or U11462 (N_11462,N_7077,N_5956);
nand U11463 (N_11463,N_9212,N_8478);
or U11464 (N_11464,N_5928,N_9402);
or U11465 (N_11465,N_5496,N_9957);
nor U11466 (N_11466,N_8265,N_8583);
nor U11467 (N_11467,N_6242,N_6253);
or U11468 (N_11468,N_8699,N_9750);
nor U11469 (N_11469,N_6066,N_6355);
and U11470 (N_11470,N_5872,N_6424);
and U11471 (N_11471,N_9023,N_5330);
xor U11472 (N_11472,N_9423,N_5776);
and U11473 (N_11473,N_6349,N_5239);
nand U11474 (N_11474,N_9838,N_7135);
nor U11475 (N_11475,N_9047,N_8082);
nor U11476 (N_11476,N_6229,N_5917);
or U11477 (N_11477,N_9230,N_7292);
nand U11478 (N_11478,N_9391,N_9508);
nor U11479 (N_11479,N_9358,N_5851);
nand U11480 (N_11480,N_9808,N_9631);
nand U11481 (N_11481,N_9951,N_5162);
and U11482 (N_11482,N_7390,N_8069);
xnor U11483 (N_11483,N_9143,N_7051);
or U11484 (N_11484,N_9248,N_8113);
nand U11485 (N_11485,N_6317,N_7179);
nand U11486 (N_11486,N_8120,N_7073);
nor U11487 (N_11487,N_5860,N_6290);
and U11488 (N_11488,N_7078,N_9926);
and U11489 (N_11489,N_6407,N_8277);
nor U11490 (N_11490,N_6108,N_8457);
and U11491 (N_11491,N_9411,N_8786);
nor U11492 (N_11492,N_9175,N_6778);
nand U11493 (N_11493,N_7416,N_5553);
nand U11494 (N_11494,N_9999,N_9386);
or U11495 (N_11495,N_7207,N_8162);
and U11496 (N_11496,N_5172,N_7388);
or U11497 (N_11497,N_8590,N_6713);
nand U11498 (N_11498,N_5645,N_7152);
nand U11499 (N_11499,N_5020,N_9282);
xor U11500 (N_11500,N_5556,N_5435);
nor U11501 (N_11501,N_5829,N_9199);
nand U11502 (N_11502,N_6361,N_7096);
xnor U11503 (N_11503,N_6337,N_8303);
nor U11504 (N_11504,N_9366,N_5122);
or U11505 (N_11505,N_6865,N_5101);
or U11506 (N_11506,N_9850,N_6400);
xnor U11507 (N_11507,N_9469,N_8553);
and U11508 (N_11508,N_9589,N_9829);
nand U11509 (N_11509,N_8341,N_5075);
and U11510 (N_11510,N_9695,N_5350);
and U11511 (N_11511,N_6418,N_8926);
nand U11512 (N_11512,N_5416,N_7016);
nand U11513 (N_11513,N_8993,N_8139);
nand U11514 (N_11514,N_8715,N_7656);
and U11515 (N_11515,N_7721,N_8889);
nor U11516 (N_11516,N_8073,N_6852);
nand U11517 (N_11517,N_7462,N_7158);
nand U11518 (N_11518,N_7487,N_7336);
and U11519 (N_11519,N_6232,N_7574);
nand U11520 (N_11520,N_6247,N_5440);
nand U11521 (N_11521,N_7186,N_6405);
nor U11522 (N_11522,N_5695,N_6584);
nor U11523 (N_11523,N_8965,N_7558);
or U11524 (N_11524,N_7294,N_5152);
xnor U11525 (N_11525,N_8443,N_9150);
and U11526 (N_11526,N_8305,N_9243);
nand U11527 (N_11527,N_6695,N_5303);
nand U11528 (N_11528,N_6372,N_8181);
xnor U11529 (N_11529,N_8228,N_9626);
nand U11530 (N_11530,N_9394,N_9613);
nor U11531 (N_11531,N_6744,N_5967);
nor U11532 (N_11532,N_6479,N_9229);
and U11533 (N_11533,N_6818,N_7652);
nand U11534 (N_11534,N_8780,N_8076);
xnor U11535 (N_11535,N_5916,N_8521);
or U11536 (N_11536,N_7386,N_6938);
or U11537 (N_11537,N_6316,N_7398);
nor U11538 (N_11538,N_8736,N_7401);
nand U11539 (N_11539,N_5488,N_6379);
nand U11540 (N_11540,N_6064,N_6406);
nor U11541 (N_11541,N_8524,N_9866);
or U11542 (N_11542,N_8586,N_9427);
or U11543 (N_11543,N_8957,N_6488);
nor U11544 (N_11544,N_6622,N_7117);
nor U11545 (N_11545,N_9055,N_5778);
and U11546 (N_11546,N_6716,N_7350);
or U11547 (N_11547,N_7567,N_8239);
or U11548 (N_11548,N_5422,N_6668);
nand U11549 (N_11549,N_7993,N_7979);
and U11550 (N_11550,N_6416,N_6920);
nor U11551 (N_11551,N_8169,N_7080);
and U11552 (N_11552,N_5057,N_8761);
nor U11553 (N_11553,N_7323,N_7910);
and U11554 (N_11554,N_8907,N_5447);
nor U11555 (N_11555,N_5722,N_5338);
nor U11556 (N_11556,N_8043,N_6035);
nand U11557 (N_11557,N_8539,N_9785);
nand U11558 (N_11558,N_5951,N_6520);
and U11559 (N_11559,N_8289,N_5886);
nand U11560 (N_11560,N_9907,N_5949);
nor U11561 (N_11561,N_6130,N_9553);
nor U11562 (N_11562,N_8574,N_8558);
nand U11563 (N_11563,N_5137,N_6387);
nand U11564 (N_11564,N_7582,N_6760);
and U11565 (N_11565,N_9779,N_5791);
xnor U11566 (N_11566,N_5988,N_7380);
nand U11567 (N_11567,N_6815,N_6094);
or U11568 (N_11568,N_6827,N_9753);
nor U11569 (N_11569,N_9839,N_6256);
and U11570 (N_11570,N_5652,N_5953);
or U11571 (N_11571,N_9420,N_5980);
or U11572 (N_11572,N_7831,N_5313);
or U11573 (N_11573,N_9131,N_7933);
nand U11574 (N_11574,N_9272,N_6857);
nor U11575 (N_11575,N_5853,N_9720);
nand U11576 (N_11576,N_5752,N_8297);
nand U11577 (N_11577,N_6854,N_7240);
or U11578 (N_11578,N_5518,N_6230);
nor U11579 (N_11579,N_5687,N_5555);
xor U11580 (N_11580,N_5533,N_9030);
or U11581 (N_11581,N_8755,N_9040);
or U11582 (N_11582,N_7013,N_7983);
or U11583 (N_11583,N_7976,N_5684);
nor U11584 (N_11584,N_6554,N_7580);
and U11585 (N_11585,N_7116,N_7739);
and U11586 (N_11586,N_6876,N_5469);
xor U11587 (N_11587,N_9511,N_7764);
nand U11588 (N_11588,N_9324,N_8532);
nand U11589 (N_11589,N_9270,N_7728);
and U11590 (N_11590,N_8947,N_9260);
and U11591 (N_11591,N_7999,N_8386);
xnor U11592 (N_11592,N_8681,N_6979);
nand U11593 (N_11593,N_5461,N_5990);
nand U11594 (N_11594,N_5066,N_7208);
and U11595 (N_11595,N_8351,N_9424);
and U11596 (N_11596,N_8368,N_5947);
and U11597 (N_11597,N_9923,N_8862);
or U11598 (N_11598,N_6157,N_5236);
or U11599 (N_11599,N_5298,N_8855);
and U11600 (N_11600,N_6492,N_5305);
nor U11601 (N_11601,N_9140,N_7801);
xnor U11602 (N_11602,N_7354,N_8317);
nand U11603 (N_11603,N_5240,N_8098);
nand U11604 (N_11604,N_6452,N_6866);
or U11605 (N_11605,N_5968,N_8692);
and U11606 (N_11606,N_8911,N_7705);
or U11607 (N_11607,N_6846,N_7319);
nand U11608 (N_11608,N_6445,N_8048);
and U11609 (N_11609,N_6132,N_5568);
and U11610 (N_11610,N_8191,N_6719);
nor U11611 (N_11611,N_6674,N_7878);
xor U11612 (N_11612,N_7564,N_8044);
nor U11613 (N_11613,N_5212,N_7606);
or U11614 (N_11614,N_9211,N_8352);
and U11615 (N_11615,N_5177,N_9461);
and U11616 (N_11616,N_9688,N_9893);
or U11617 (N_11617,N_5869,N_8811);
xnor U11618 (N_11618,N_9982,N_8260);
nor U11619 (N_11619,N_6966,N_5333);
nor U11620 (N_11620,N_7298,N_6067);
and U11621 (N_11621,N_8735,N_9591);
nor U11622 (N_11622,N_8771,N_9763);
or U11623 (N_11623,N_8408,N_6389);
and U11624 (N_11624,N_7205,N_7994);
or U11625 (N_11625,N_5114,N_8206);
xor U11626 (N_11626,N_5138,N_9413);
nor U11627 (N_11627,N_8619,N_9558);
nand U11628 (N_11628,N_8041,N_8548);
xnor U11629 (N_11629,N_7914,N_7364);
and U11630 (N_11630,N_5954,N_8830);
nand U11631 (N_11631,N_8204,N_9083);
nand U11632 (N_11632,N_8649,N_5966);
and U11633 (N_11633,N_9065,N_9756);
and U11634 (N_11634,N_9758,N_9505);
nor U11635 (N_11635,N_8962,N_7332);
xor U11636 (N_11636,N_8805,N_6627);
nor U11637 (N_11637,N_7506,N_5803);
and U11638 (N_11638,N_8596,N_9717);
or U11639 (N_11639,N_9692,N_6453);
nand U11640 (N_11640,N_6022,N_6675);
xor U11641 (N_11641,N_5043,N_7702);
and U11642 (N_11642,N_7351,N_7495);
nor U11643 (N_11643,N_7896,N_7603);
or U11644 (N_11644,N_6909,N_5546);
nor U11645 (N_11645,N_6218,N_5314);
and U11646 (N_11646,N_5847,N_5581);
nor U11647 (N_11647,N_7671,N_7646);
or U11648 (N_11648,N_7588,N_7095);
nor U11649 (N_11649,N_8508,N_7892);
and U11650 (N_11650,N_6929,N_7570);
nand U11651 (N_11651,N_9787,N_6200);
nor U11652 (N_11652,N_9716,N_7066);
nand U11653 (N_11653,N_6628,N_8906);
nor U11654 (N_11654,N_9086,N_7763);
and U11655 (N_11655,N_6456,N_7251);
nor U11656 (N_11656,N_9672,N_5697);
nor U11657 (N_11657,N_7025,N_6048);
or U11658 (N_11658,N_8846,N_7571);
or U11659 (N_11659,N_6991,N_6745);
and U11660 (N_11660,N_5468,N_7880);
nor U11661 (N_11661,N_8328,N_7408);
nor U11662 (N_11662,N_6217,N_8983);
nor U11663 (N_11663,N_6786,N_9003);
nor U11664 (N_11664,N_9137,N_9579);
or U11665 (N_11665,N_6216,N_5838);
and U11666 (N_11666,N_9539,N_8236);
and U11667 (N_11667,N_7875,N_8787);
nor U11668 (N_11668,N_7133,N_7404);
and U11669 (N_11669,N_5505,N_9904);
nor U11670 (N_11670,N_7840,N_9385);
nor U11671 (N_11671,N_5208,N_8074);
or U11672 (N_11672,N_6562,N_9699);
or U11673 (N_11673,N_7041,N_6287);
nand U11674 (N_11674,N_6972,N_5362);
nand U11675 (N_11675,N_6221,N_9646);
or U11676 (N_11676,N_6391,N_9474);
nor U11677 (N_11677,N_9882,N_5888);
nor U11678 (N_11678,N_9302,N_8186);
nand U11679 (N_11679,N_8719,N_9513);
nand U11680 (N_11680,N_6613,N_7081);
xnor U11681 (N_11681,N_6471,N_6070);
and U11682 (N_11682,N_5317,N_5771);
nand U11683 (N_11683,N_8656,N_8633);
nor U11684 (N_11684,N_6600,N_7147);
and U11685 (N_11685,N_8772,N_7627);
nor U11686 (N_11686,N_9827,N_8660);
and U11687 (N_11687,N_9305,N_8401);
nor U11688 (N_11688,N_9096,N_6607);
nor U11689 (N_11689,N_6918,N_5282);
nand U11690 (N_11690,N_6728,N_5286);
and U11691 (N_11691,N_5480,N_5364);
nor U11692 (N_11692,N_6599,N_8151);
and U11693 (N_11693,N_6166,N_6781);
or U11694 (N_11694,N_9742,N_5604);
and U11695 (N_11695,N_8800,N_9347);
and U11696 (N_11696,N_9724,N_7954);
xnor U11697 (N_11697,N_6111,N_9624);
nand U11698 (N_11698,N_5671,N_6872);
nand U11699 (N_11699,N_8917,N_7005);
xnor U11700 (N_11700,N_6305,N_5347);
or U11701 (N_11701,N_9457,N_7766);
nand U11702 (N_11702,N_5029,N_6926);
and U11703 (N_11703,N_6908,N_6949);
xor U11704 (N_11704,N_6176,N_5245);
xor U11705 (N_11705,N_9986,N_7666);
or U11706 (N_11706,N_9565,N_7974);
and U11707 (N_11707,N_7498,N_5766);
and U11708 (N_11708,N_6736,N_5096);
and U11709 (N_11709,N_5232,N_7375);
nand U11710 (N_11710,N_6841,N_8461);
nor U11711 (N_11711,N_6332,N_9345);
nor U11712 (N_11712,N_6644,N_9444);
and U11713 (N_11713,N_8668,N_9561);
nand U11714 (N_11714,N_8617,N_9032);
and U11715 (N_11715,N_7546,N_5198);
and U11716 (N_11716,N_6423,N_8666);
nand U11717 (N_11717,N_8844,N_6091);
xnor U11718 (N_11718,N_9950,N_9205);
nor U11719 (N_11719,N_6861,N_6910);
or U11720 (N_11720,N_5741,N_6073);
nand U11721 (N_11721,N_7278,N_7368);
or U11722 (N_11722,N_9300,N_6980);
nor U11723 (N_11723,N_6616,N_5526);
xnor U11724 (N_11724,N_5453,N_6404);
and U11725 (N_11725,N_7586,N_9356);
nor U11726 (N_11726,N_5592,N_9108);
and U11727 (N_11727,N_5509,N_5938);
nand U11728 (N_11728,N_8882,N_7926);
nor U11729 (N_11729,N_5487,N_5575);
nor U11730 (N_11730,N_6688,N_9126);
nor U11731 (N_11731,N_7441,N_8189);
and U11732 (N_11732,N_9519,N_6632);
or U11733 (N_11733,N_5993,N_6052);
or U11734 (N_11734,N_8106,N_7445);
or U11735 (N_11735,N_7725,N_9309);
xnor U11736 (N_11736,N_5180,N_9367);
nand U11737 (N_11737,N_7863,N_6263);
or U11738 (N_11738,N_9600,N_9005);
and U11739 (N_11739,N_7512,N_7950);
or U11740 (N_11740,N_7859,N_6825);
nor U11741 (N_11741,N_9977,N_8714);
or U11742 (N_11742,N_6348,N_9985);
xor U11743 (N_11743,N_5402,N_9530);
and U11744 (N_11744,N_7118,N_5542);
or U11745 (N_11745,N_8964,N_6967);
nand U11746 (N_11746,N_8635,N_8016);
or U11747 (N_11747,N_5024,N_9271);
and U11748 (N_11748,N_6990,N_5205);
nor U11749 (N_11749,N_7793,N_7111);
nand U11750 (N_11750,N_8944,N_5186);
nor U11751 (N_11751,N_7055,N_7674);
nor U11752 (N_11752,N_7173,N_6620);
and U11753 (N_11753,N_6208,N_7795);
nor U11754 (N_11754,N_7928,N_8813);
nor U11755 (N_11755,N_7642,N_9492);
and U11756 (N_11756,N_5981,N_7022);
and U11757 (N_11757,N_7154,N_7539);
and U11758 (N_11758,N_7560,N_8017);
nand U11759 (N_11759,N_9123,N_7394);
and U11760 (N_11760,N_6298,N_9489);
nand U11761 (N_11761,N_6096,N_7516);
nor U11762 (N_11762,N_5356,N_5070);
nor U11763 (N_11763,N_7726,N_9408);
nand U11764 (N_11764,N_8246,N_5666);
nand U11765 (N_11765,N_5458,N_8479);
nand U11766 (N_11766,N_8698,N_9480);
xnor U11767 (N_11767,N_7477,N_5769);
nor U11768 (N_11768,N_8096,N_5932);
nand U11769 (N_11769,N_9294,N_6783);
nand U11770 (N_11770,N_6474,N_6948);
and U11771 (N_11771,N_8978,N_5418);
and U11772 (N_11772,N_6752,N_5279);
and U11773 (N_11773,N_9811,N_9595);
nor U11774 (N_11774,N_7722,N_5644);
nor U11775 (N_11775,N_5183,N_7936);
and U11776 (N_11776,N_5996,N_7062);
nand U11777 (N_11777,N_5669,N_8864);
nor U11778 (N_11778,N_7921,N_9261);
nor U11779 (N_11779,N_7316,N_9185);
nor U11780 (N_11780,N_7164,N_9256);
or U11781 (N_11781,N_9280,N_6592);
nand U11782 (N_11782,N_9057,N_7835);
or U11783 (N_11783,N_5758,N_6062);
nor U11784 (N_11784,N_6828,N_7201);
nor U11785 (N_11785,N_7161,N_9090);
xor U11786 (N_11786,N_5998,N_9816);
and U11787 (N_11787,N_6222,N_8388);
or U11788 (N_11788,N_8473,N_9818);
nor U11789 (N_11789,N_6000,N_5426);
or U11790 (N_11790,N_7420,N_9946);
or U11791 (N_11791,N_6142,N_9151);
or U11792 (N_11792,N_5369,N_8857);
nor U11793 (N_11793,N_9360,N_5777);
nand U11794 (N_11794,N_6236,N_9393);
and U11795 (N_11795,N_6862,N_6791);
and U11796 (N_11796,N_9913,N_6555);
nor U11797 (N_11797,N_6112,N_6003);
and U11798 (N_11798,N_5493,N_5430);
or U11799 (N_11799,N_7775,N_5379);
or U11800 (N_11800,N_5841,N_5472);
nor U11801 (N_11801,N_9026,N_7514);
and U11802 (N_11802,N_7121,N_8146);
nor U11803 (N_11803,N_7935,N_6036);
xnor U11804 (N_11804,N_9182,N_9793);
and U11805 (N_11805,N_7338,N_5730);
xor U11806 (N_11806,N_9170,N_5112);
or U11807 (N_11807,N_5221,N_7134);
nor U11808 (N_11808,N_8072,N_7947);
and U11809 (N_11809,N_8262,N_6994);
and U11810 (N_11810,N_9807,N_7946);
or U11811 (N_11811,N_9293,N_7638);
nor U11812 (N_11812,N_7699,N_9421);
and U11813 (N_11813,N_5074,N_5133);
and U11814 (N_11814,N_8727,N_5921);
nand U11815 (N_11815,N_5994,N_7668);
xnor U11816 (N_11816,N_5955,N_9149);
and U11817 (N_11817,N_7883,N_7219);
or U11818 (N_11818,N_7852,N_9857);
or U11819 (N_11819,N_6367,N_8867);
and U11820 (N_11820,N_9437,N_6454);
nor U11821 (N_11821,N_9765,N_6598);
xor U11822 (N_11822,N_5281,N_7958);
and U11823 (N_11823,N_6426,N_9410);
or U11824 (N_11824,N_8835,N_6982);
and U11825 (N_11825,N_7470,N_6186);
xor U11826 (N_11826,N_7277,N_9396);
or U11827 (N_11827,N_7927,N_6686);
and U11828 (N_11828,N_6293,N_5595);
nor U11829 (N_11829,N_9528,N_9046);
xnor U11830 (N_11830,N_8269,N_8566);
or U11831 (N_11831,N_7200,N_5354);
xor U11832 (N_11832,N_9609,N_6274);
nand U11833 (N_11833,N_8651,N_9341);
xor U11834 (N_11834,N_6341,N_5893);
nand U11835 (N_11835,N_7502,N_9038);
and U11836 (N_11836,N_6986,N_6665);
xnor U11837 (N_11837,N_6214,N_9232);
and U11838 (N_11838,N_7711,N_6549);
nand U11839 (N_11839,N_7086,N_7053);
nand U11840 (N_11840,N_6469,N_5596);
nand U11841 (N_11841,N_6525,N_8013);
and U11842 (N_11842,N_6514,N_9638);
and U11843 (N_11843,N_7038,N_9401);
nand U11844 (N_11844,N_8192,N_5011);
or U11845 (N_11845,N_5184,N_5390);
nand U11846 (N_11846,N_5664,N_5246);
nor U11847 (N_11847,N_7169,N_9968);
and U11848 (N_11848,N_9429,N_9049);
and U11849 (N_11849,N_8778,N_6158);
xnor U11850 (N_11850,N_7071,N_8259);
nand U11851 (N_11851,N_7322,N_7326);
nor U11852 (N_11852,N_7860,N_6089);
xnor U11853 (N_11853,N_5959,N_6063);
and U11854 (N_11854,N_6806,N_5586);
and U11855 (N_11855,N_5276,N_6892);
xnor U11856 (N_11856,N_6430,N_7873);
and U11857 (N_11857,N_9939,N_9376);
nor U11858 (N_11858,N_9142,N_9557);
nand U11859 (N_11859,N_5855,N_9012);
xnor U11860 (N_11860,N_5260,N_7694);
nor U11861 (N_11861,N_5677,N_7137);
and U11862 (N_11862,N_7252,N_8875);
nand U11863 (N_11863,N_8379,N_7925);
or U11864 (N_11864,N_9585,N_5089);
nor U11865 (N_11865,N_5708,N_6354);
and U11866 (N_11866,N_6732,N_9540);
and U11867 (N_11867,N_8190,N_6942);
or U11868 (N_11868,N_6739,N_5387);
nor U11869 (N_11869,N_5154,N_9008);
and U11870 (N_11870,N_6289,N_5692);
nand U11871 (N_11871,N_5229,N_6704);
and U11872 (N_11872,N_9254,N_6086);
and U11873 (N_11873,N_9764,N_7846);
or U11874 (N_11874,N_5880,N_6618);
nor U11875 (N_11875,N_5045,N_8229);
or U11876 (N_11876,N_8067,N_8357);
xor U11877 (N_11877,N_9947,N_6120);
or U11878 (N_11878,N_9760,N_5202);
and U11879 (N_11879,N_6043,N_9441);
and U11880 (N_11880,N_5618,N_7818);
nor U11881 (N_11881,N_7360,N_8640);
nor U11882 (N_11882,N_5873,N_7218);
nand U11883 (N_11883,N_9989,N_5455);
or U11884 (N_11884,N_9081,N_5693);
or U11885 (N_11885,N_9698,N_9541);
nor U11886 (N_11886,N_5743,N_5196);
xnor U11887 (N_11887,N_8039,N_8997);
nand U11888 (N_11888,N_6691,N_6960);
or U11889 (N_11889,N_7990,N_9562);
nand U11890 (N_11890,N_8006,N_7145);
nand U11891 (N_11891,N_8770,N_9350);
and U11892 (N_11892,N_7359,N_7894);
and U11893 (N_11893,N_8207,N_6566);
or U11894 (N_11894,N_8089,N_9063);
or U11895 (N_11895,N_6621,N_6891);
or U11896 (N_11896,N_6363,N_6853);
or U11897 (N_11897,N_8950,N_7267);
or U11898 (N_11898,N_9798,N_7021);
or U11899 (N_11899,N_9035,N_7299);
nor U11900 (N_11900,N_8985,N_6312);
nand U11901 (N_11901,N_7464,N_7122);
and U11902 (N_11902,N_9745,N_9290);
or U11903 (N_11903,N_7342,N_9406);
nor U11904 (N_11904,N_6868,N_9414);
nor U11905 (N_11905,N_6581,N_7262);
or U11906 (N_11906,N_8712,N_7093);
or U11907 (N_11907,N_8860,N_5567);
and U11908 (N_11908,N_7520,N_6016);
or U11909 (N_11909,N_9618,N_7507);
or U11910 (N_11910,N_5836,N_9037);
or U11911 (N_11911,N_9052,N_5217);
or U11912 (N_11912,N_6822,N_6155);
and U11913 (N_11913,N_8400,N_7193);
or U11914 (N_11914,N_6359,N_9095);
or U11915 (N_11915,N_8394,N_8054);
nor U11916 (N_11916,N_8483,N_8431);
nand U11917 (N_11917,N_8023,N_9157);
nand U11918 (N_11918,N_9863,N_7324);
or U11919 (N_11919,N_9153,N_8746);
nor U11920 (N_11920,N_8398,N_6443);
nor U11921 (N_11921,N_6039,N_8094);
nand U11922 (N_11922,N_7951,N_7714);
xnor U11923 (N_11923,N_7191,N_5579);
or U11924 (N_11924,N_5527,N_9100);
and U11925 (N_11925,N_6258,N_7542);
xor U11926 (N_11926,N_6800,N_9676);
nand U11927 (N_11927,N_5128,N_5877);
nor U11928 (N_11928,N_9113,N_5611);
or U11929 (N_11929,N_6249,N_6533);
xnor U11930 (N_11930,N_5182,N_9014);
xor U11931 (N_11931,N_6558,N_9786);
nor U11932 (N_11932,N_5341,N_6804);
xnor U11933 (N_11933,N_8517,N_9227);
and U11934 (N_11934,N_5044,N_7853);
xnor U11935 (N_11935,N_8795,N_8238);
nor U11936 (N_11936,N_6192,N_8602);
or U11937 (N_11937,N_7039,N_6449);
or U11938 (N_11938,N_6624,N_6843);
xor U11939 (N_11939,N_6532,N_8211);
nand U11940 (N_11940,N_8126,N_5079);
or U11941 (N_11941,N_8568,N_7499);
and U11942 (N_11942,N_8589,N_8972);
or U11943 (N_11943,N_8438,N_7716);
nand U11944 (N_11944,N_7203,N_9691);
and U11945 (N_11945,N_5474,N_9467);
nor U11946 (N_11946,N_8240,N_5566);
xnor U11947 (N_11947,N_8359,N_5028);
and U11948 (N_11948,N_6919,N_5257);
nand U11949 (N_11949,N_7978,N_6145);
and U11950 (N_11950,N_9934,N_8346);
or U11951 (N_11951,N_7413,N_7643);
xor U11952 (N_11952,N_7904,N_5105);
and U11953 (N_11953,N_7601,N_8653);
nor U11954 (N_11954,N_5952,N_6476);
nand U11955 (N_11955,N_9332,N_6660);
nand U11956 (N_11956,N_9955,N_9029);
nand U11957 (N_11957,N_7989,N_8923);
nor U11958 (N_11958,N_7515,N_8820);
xor U11959 (N_11959,N_6446,N_6027);
nand U11960 (N_11960,N_7658,N_5001);
nor U11961 (N_11961,N_7045,N_8156);
or U11962 (N_11962,N_7779,N_7230);
and U11963 (N_11963,N_5344,N_9226);
xor U11964 (N_11964,N_8278,N_8337);
xnor U11965 (N_11965,N_8312,N_6681);
and U11966 (N_11966,N_9607,N_8910);
nand U11967 (N_11967,N_5643,N_8740);
nand U11968 (N_11968,N_8348,N_8071);
xor U11969 (N_11969,N_5889,N_7689);
or U11970 (N_11970,N_9190,N_9392);
nor U11971 (N_11971,N_8542,N_5002);
or U11972 (N_11972,N_8225,N_5950);
nor U11973 (N_11973,N_9129,N_9015);
or U11974 (N_11974,N_5835,N_6184);
nand U11975 (N_11975,N_7451,N_7738);
or U11976 (N_11976,N_9114,N_5401);
or U11977 (N_11977,N_5606,N_8801);
and U11978 (N_11978,N_8429,N_9088);
and U11979 (N_11979,N_7306,N_5727);
nor U11980 (N_11980,N_5149,N_8155);
or U11981 (N_11981,N_9449,N_8138);
nor U11982 (N_11982,N_8350,N_9317);
and U11983 (N_11983,N_9997,N_5738);
nor U11984 (N_11984,N_5562,N_6434);
nand U11985 (N_11985,N_5220,N_5302);
and U11986 (N_11986,N_5675,N_8682);
and U11987 (N_11987,N_9629,N_5464);
nand U11988 (N_11988,N_8087,N_8081);
nand U11989 (N_11989,N_9747,N_6589);
or U11990 (N_11990,N_8812,N_8343);
xnor U11991 (N_11991,N_5499,N_9310);
nand U11992 (N_11992,N_9835,N_9710);
nand U11993 (N_11993,N_9694,N_9438);
or U11994 (N_11994,N_9400,N_9908);
and U11995 (N_11995,N_7002,N_9099);
nor U11996 (N_11996,N_5805,N_7521);
nor U11997 (N_11997,N_7774,N_8318);
and U11998 (N_11998,N_5942,N_5676);
and U11999 (N_11999,N_8613,N_9658);
nor U12000 (N_12000,N_9549,N_9103);
or U12001 (N_12001,N_7263,N_9146);
nor U12002 (N_12002,N_6951,N_9322);
nand U12003 (N_12003,N_8480,N_8686);
or U12004 (N_12004,N_7049,N_8636);
nand U12005 (N_12005,N_6829,N_5849);
nor U12006 (N_12006,N_8209,N_9870);
nor U12007 (N_12007,N_7199,N_7297);
and U12008 (N_12008,N_7737,N_6436);
or U12009 (N_12009,N_5443,N_9824);
nor U12010 (N_12010,N_5065,N_6647);
or U12011 (N_12011,N_8449,N_7911);
nand U12012 (N_12012,N_9571,N_6001);
xor U12013 (N_12013,N_6276,N_9552);
or U12014 (N_12014,N_6945,N_8892);
and U12015 (N_12015,N_5439,N_6038);
or U12016 (N_12016,N_6955,N_8897);
and U12017 (N_12017,N_5638,N_8037);
nand U12018 (N_12018,N_5508,N_7886);
nor U12019 (N_12019,N_9267,N_5972);
nand U12020 (N_12020,N_7165,N_5906);
nand U12021 (N_12021,N_7527,N_7241);
nand U12022 (N_12022,N_8557,N_6623);
or U12023 (N_12023,N_9652,N_9010);
and U12024 (N_12024,N_7884,N_9321);
and U12025 (N_12025,N_8606,N_9642);
or U12026 (N_12026,N_5327,N_7566);
nor U12027 (N_12027,N_8103,N_9622);
nand U12028 (N_12028,N_6150,N_6758);
nor U12029 (N_12029,N_6583,N_5767);
xor U12030 (N_12030,N_9996,N_6358);
nor U12031 (N_12031,N_5846,N_6402);
nand U12032 (N_12032,N_9219,N_6856);
nor U12033 (N_12033,N_5242,N_9432);
xor U12034 (N_12034,N_6466,N_8999);
or U12035 (N_12035,N_7913,N_5213);
nor U12036 (N_12036,N_6773,N_6523);
nor U12037 (N_12037,N_7378,N_9730);
and U12038 (N_12038,N_5721,N_7813);
or U12039 (N_12039,N_8020,N_5828);
nand U12040 (N_12040,N_6518,N_7552);
xor U12041 (N_12041,N_7235,N_6172);
and U12042 (N_12042,N_5163,N_7391);
and U12043 (N_12043,N_9598,N_7097);
xnor U12044 (N_12044,N_5166,N_8476);
nor U12045 (N_12045,N_9774,N_6727);
and U12046 (N_12046,N_8570,N_7130);
xnor U12047 (N_12047,N_7372,N_6528);
or U12048 (N_12048,N_9810,N_5635);
nand U12049 (N_12049,N_8042,N_5312);
nand U12050 (N_12050,N_6881,N_5235);
nor U12051 (N_12051,N_9209,N_7879);
nand U12052 (N_12052,N_8267,N_5187);
and U12053 (N_12053,N_5995,N_9846);
nand U12054 (N_12054,N_8008,N_8604);
or U12055 (N_12055,N_5620,N_8374);
and U12056 (N_12056,N_9139,N_8161);
and U12057 (N_12057,N_9463,N_8417);
nor U12058 (N_12058,N_9458,N_5399);
nor U12059 (N_12059,N_8257,N_6896);
or U12060 (N_12060,N_8580,N_9621);
nor U12061 (N_12061,N_9680,N_8526);
nand U12062 (N_12062,N_5919,N_6213);
and U12063 (N_12063,N_5040,N_8672);
or U12064 (N_12064,N_9118,N_7075);
or U12065 (N_12065,N_6190,N_6260);
nand U12066 (N_12066,N_6055,N_8032);
xor U12067 (N_12067,N_7969,N_6871);
xnor U12068 (N_12068,N_8914,N_7600);
nor U12069 (N_12069,N_9013,N_7198);
or U12070 (N_12070,N_7226,N_6269);
and U12071 (N_12071,N_9578,N_7593);
and U12072 (N_12072,N_7916,N_8946);
xor U12073 (N_12073,N_7987,N_7269);
and U12074 (N_12074,N_9031,N_7678);
nor U12075 (N_12075,N_9249,N_6844);
nor U12076 (N_12076,N_8959,N_6224);
or U12077 (N_12077,N_6965,N_9566);
and U12078 (N_12078,N_7153,N_7712);
or U12079 (N_12079,N_9292,N_8105);
or U12080 (N_12080,N_9000,N_6018);
or U12081 (N_12081,N_7312,N_8152);
nor U12082 (N_12082,N_6842,N_7127);
nand U12083 (N_12083,N_8304,N_5824);
nor U12084 (N_12084,N_7079,N_8085);
nand U12085 (N_12085,N_8030,N_6388);
nor U12086 (N_12086,N_9651,N_8571);
and U12087 (N_12087,N_5392,N_7771);
or U12088 (N_12088,N_8292,N_8331);
or U12089 (N_12089,N_8293,N_8427);
xnor U12090 (N_12090,N_6364,N_9235);
nor U12091 (N_12091,N_5051,N_6999);
nand U12092 (N_12092,N_7435,N_7092);
nor U12093 (N_12093,N_7536,N_8075);
or U12094 (N_12094,N_9533,N_8384);
or U12095 (N_12095,N_7948,N_6564);
nand U12096 (N_12096,N_7977,N_7787);
nand U12097 (N_12097,N_9434,N_8254);
and U12098 (N_12098,N_9602,N_8281);
nand U12099 (N_12099,N_7496,N_6751);
and U12100 (N_12100,N_7623,N_6347);
and U12101 (N_12101,N_5924,N_6410);
and U12102 (N_12102,N_6353,N_5551);
nor U12103 (N_12103,N_6930,N_5519);
and U12104 (N_12104,N_9635,N_8149);
and U12105 (N_12105,N_5660,N_7412);
xnor U12106 (N_12106,N_9732,N_8704);
nand U12107 (N_12107,N_9102,N_5365);
nand U12108 (N_12108,N_8001,N_6826);
or U12109 (N_12109,N_9605,N_8099);
nand U12110 (N_12110,N_8669,N_8996);
nor U12111 (N_12111,N_9852,N_5502);
and U12112 (N_12112,N_9868,N_7124);
xnor U12113 (N_12113,N_9820,N_7830);
and U12114 (N_12114,N_5197,N_8842);
xor U12115 (N_12115,N_5642,N_6724);
nand U12116 (N_12116,N_8021,N_5377);
nand U12117 (N_12117,N_7223,N_8610);
xor U12118 (N_12118,N_8981,N_9766);
and U12119 (N_12119,N_8877,N_7583);
nand U12120 (N_12120,N_9915,N_7027);
nor U12121 (N_12121,N_5385,N_5410);
or U12122 (N_12122,N_8540,N_7261);
nand U12123 (N_12123,N_6869,N_5366);
nand U12124 (N_12124,N_7862,N_5316);
xor U12125 (N_12125,N_6513,N_8176);
xor U12126 (N_12126,N_6521,N_8179);
nand U12127 (N_12127,N_5629,N_7166);
nor U12128 (N_12128,N_8285,N_9895);
and U12129 (N_12129,N_8559,N_9128);
or U12130 (N_12130,N_9718,N_5634);
xor U12131 (N_12131,N_5296,N_7806);
or U12132 (N_12132,N_6934,N_7281);
xor U12133 (N_12133,N_7908,N_5160);
or U12134 (N_12134,N_9980,N_9450);
nor U12135 (N_12135,N_5495,N_9911);
nand U12136 (N_12136,N_5175,N_7673);
or U12137 (N_12137,N_7640,N_7709);
or U12138 (N_12138,N_7023,N_8221);
and U12139 (N_12139,N_5093,N_9204);
or U12140 (N_12140,N_5926,N_5915);
nand U12141 (N_12141,N_6148,N_7028);
nor U12142 (N_12142,N_5063,N_8785);
nor U12143 (N_12143,N_9604,N_7504);
or U12144 (N_12144,N_5503,N_6390);
xnor U12145 (N_12145,N_6115,N_7463);
and U12146 (N_12146,N_6638,N_6676);
or U12147 (N_12147,N_7151,N_6212);
nor U12148 (N_12148,N_8136,N_9965);
or U12149 (N_12149,N_7009,N_5309);
or U12150 (N_12150,N_7768,N_7000);
or U12151 (N_12151,N_7489,N_8625);
nor U12152 (N_12152,N_6637,N_7255);
or U12153 (N_12153,N_6427,N_8490);
or U12154 (N_12154,N_5612,N_7438);
nor U12155 (N_12155,N_7667,N_8487);
xor U12156 (N_12156,N_9166,N_9036);
and U12157 (N_12157,N_6301,N_8689);
nand U12158 (N_12158,N_8980,N_8382);
and U12159 (N_12159,N_9172,N_6458);
nand U12160 (N_12160,N_8203,N_5899);
nor U12161 (N_12161,N_7587,N_7289);
nor U12162 (N_12162,N_7132,N_5622);
nor U12163 (N_12163,N_5707,N_9224);
nor U12164 (N_12164,N_6050,N_7631);
nand U12165 (N_12165,N_5673,N_5143);
or U12166 (N_12166,N_8402,N_6764);
xnor U12167 (N_12167,N_6059,N_5520);
nand U12168 (N_12168,N_9817,N_8340);
nor U12169 (N_12169,N_5324,N_8380);
and U12170 (N_12170,N_5211,N_5429);
and U12171 (N_12171,N_7553,N_6116);
and U12172 (N_12172,N_6336,N_8347);
or U12173 (N_12173,N_9183,N_6451);
nand U12174 (N_12174,N_9640,N_8275);
or U12175 (N_12175,N_5997,N_5463);
and U12176 (N_12176,N_6536,N_6611);
xor U12177 (N_12177,N_8850,N_6997);
and U12178 (N_12178,N_7690,N_6928);
nand U12179 (N_12179,N_9544,N_9468);
xor U12180 (N_12180,N_6937,N_8631);
and U12181 (N_12181,N_7054,N_8628);
or U12182 (N_12182,N_6805,N_5745);
and U12183 (N_12183,N_6677,N_7157);
and U12184 (N_12184,N_8880,N_8955);
and U12185 (N_12185,N_7099,N_8550);
nand U12186 (N_12186,N_7069,N_8956);
or U12187 (N_12187,N_7632,N_5168);
nand U12188 (N_12188,N_7037,N_7790);
nand U12189 (N_12189,N_8925,N_7494);
and U12190 (N_12190,N_7065,N_7800);
or U12191 (N_12191,N_9433,N_6380);
nor U12192 (N_12192,N_8995,N_7727);
nand U12193 (N_12193,N_9279,N_9531);
nand U12194 (N_12194,N_6664,N_9840);
nand U12195 (N_12195,N_5009,N_6743);
nor U12196 (N_12196,N_6901,N_5054);
or U12197 (N_12197,N_9246,N_6629);
xnor U12198 (N_12198,N_6490,N_6060);
nand U12199 (N_12199,N_7379,N_5696);
nor U12200 (N_12200,N_7660,N_7973);
and U12201 (N_12201,N_9497,N_7789);
nor U12202 (N_12202,N_9641,N_5858);
and U12203 (N_12203,N_8077,N_7197);
nor U12204 (N_12204,N_7385,N_8205);
xnor U12205 (N_12205,N_7900,N_7533);
and U12206 (N_12206,N_8859,N_8954);
and U12207 (N_12207,N_6546,N_9329);
or U12208 (N_12208,N_9856,N_9888);
nor U12209 (N_12209,N_8080,N_8798);
and U12210 (N_12210,N_6735,N_8807);
nand U12211 (N_12211,N_8100,N_5452);
xor U12212 (N_12212,N_5403,N_9078);
nor U12213 (N_12213,N_8137,N_7148);
xor U12214 (N_12214,N_5810,N_9919);
or U12215 (N_12215,N_6352,N_8973);
nand U12216 (N_12216,N_9963,N_8869);
and U12217 (N_12217,N_5203,N_6988);
nand U12218 (N_12218,N_6835,N_7155);
and U12219 (N_12219,N_9871,N_7369);
nor U12220 (N_12220,N_8938,N_8036);
nor U12221 (N_12221,N_8769,N_6023);
nand U12222 (N_12222,N_8243,N_9009);
and U12223 (N_12223,N_8797,N_5714);
nand U12224 (N_12224,N_6776,N_9686);
and U12225 (N_12225,N_5601,N_9027);
xnor U12226 (N_12226,N_6655,N_8420);
nand U12227 (N_12227,N_8650,N_9383);
nor U12228 (N_12228,N_9056,N_5549);
and U12229 (N_12229,N_8537,N_9200);
and U12230 (N_12230,N_6779,N_6447);
nor U12231 (N_12231,N_9782,N_8541);
nor U12232 (N_12232,N_5852,N_9325);
nor U12233 (N_12233,N_8924,N_6759);
nor U12234 (N_12234,N_9340,N_5935);
and U12235 (N_12235,N_6470,N_9790);
nand U12236 (N_12236,N_7432,N_9804);
and U12237 (N_12237,N_7731,N_8064);
and U12238 (N_12238,N_9815,N_6034);
nand U12239 (N_12239,N_7449,N_9415);
and U12240 (N_12240,N_5284,N_9944);
nor U12241 (N_12241,N_6194,N_8310);
nand U12242 (N_12242,N_8436,N_5032);
nor U12243 (N_12243,N_8967,N_5603);
and U12244 (N_12244,N_7362,N_9559);
xnor U12245 (N_12245,N_7213,N_6810);
nand U12246 (N_12246,N_9382,N_8607);
or U12247 (N_12247,N_5335,N_5104);
or U12248 (N_12248,N_5544,N_7331);
nand U12249 (N_12249,N_6121,N_6206);
and U12250 (N_12250,N_8671,N_9861);
and U12251 (N_12251,N_9594,N_6653);
xnor U12252 (N_12252,N_8173,N_8355);
and U12253 (N_12253,N_8049,N_8070);
nor U12254 (N_12254,N_9708,N_9162);
nand U12255 (N_12255,N_8849,N_8178);
nand U12256 (N_12256,N_6996,N_9165);
nand U12257 (N_12257,N_6912,N_7857);
and U12258 (N_12258,N_8936,N_9452);
nand U12259 (N_12259,N_5269,N_5030);
and U12260 (N_12260,N_7453,N_6008);
nor U12261 (N_12261,N_5637,N_8608);
xnor U12262 (N_12262,N_8626,N_5088);
or U12263 (N_12263,N_7216,N_6897);
nand U12264 (N_12264,N_6640,N_8783);
or U12265 (N_12265,N_8302,N_5391);
nor U12266 (N_12266,N_9872,N_6859);
nor U12267 (N_12267,N_6879,N_7410);
nor U12268 (N_12268,N_7700,N_9567);
or U12269 (N_12269,N_9419,N_9352);
nor U12270 (N_12270,N_6535,N_5444);
nor U12271 (N_12271,N_9702,N_6160);
and U12272 (N_12272,N_9781,N_8572);
nor U12273 (N_12273,N_5819,N_9186);
nand U12274 (N_12274,N_5649,N_8505);
nor U12275 (N_12275,N_7437,N_9287);
and U12276 (N_12276,N_6450,N_6798);
nand U12277 (N_12277,N_8160,N_7406);
xnor U12278 (N_12278,N_5564,N_9117);
nor U12279 (N_12279,N_6684,N_6246);
or U12280 (N_12280,N_7929,N_6894);
or U12281 (N_12281,N_6065,N_8529);
nand U12282 (N_12282,N_9448,N_8498);
or U12283 (N_12283,N_6496,N_6515);
nand U12284 (N_12284,N_9657,N_8390);
or U12285 (N_12285,N_9684,N_6580);
and U12286 (N_12286,N_9233,N_6233);
or U12287 (N_12287,N_8843,N_8248);
xnor U12288 (N_12288,N_9693,N_9555);
nand U12289 (N_12289,N_7128,N_8059);
nand U12290 (N_12290,N_7232,N_6932);
nor U12291 (N_12291,N_5744,N_5227);
and U12292 (N_12292,N_6360,N_7458);
xnor U12293 (N_12293,N_6422,N_7971);
xor U12294 (N_12294,N_6658,N_7868);
or U12295 (N_12295,N_8118,N_5442);
nor U12296 (N_12296,N_8296,N_7283);
or U12297 (N_12297,N_5360,N_6056);
nand U12298 (N_12298,N_8902,N_7467);
nand U12299 (N_12299,N_7578,N_6169);
nor U12300 (N_12300,N_5976,N_5790);
nand U12301 (N_12301,N_9831,N_8244);
and U12302 (N_12302,N_5099,N_6013);
nand U12303 (N_12303,N_9734,N_7704);
xnor U12304 (N_12304,N_8593,N_5384);
nor U12305 (N_12305,N_8918,N_5072);
or U12306 (N_12306,N_5334,N_8988);
nor U12307 (N_12307,N_8029,N_8216);
or U12308 (N_12308,N_7555,N_7288);
or U12309 (N_12309,N_8986,N_6530);
or U12310 (N_12310,N_5960,N_6147);
or U12311 (N_12311,N_5234,N_6529);
nor U12312 (N_12312,N_8167,N_9875);
and U12313 (N_12313,N_6197,N_7108);
nor U12314 (N_12314,N_9668,N_7836);
or U12315 (N_12315,N_7233,N_8378);
and U12316 (N_12316,N_7556,N_8301);
and U12317 (N_12317,N_5715,N_6936);
nor U12318 (N_12318,N_6701,N_8545);
nand U12319 (N_12319,N_5720,N_7669);
and U12320 (N_12320,N_9851,N_9931);
and U12321 (N_12321,N_5109,N_7829);
or U12322 (N_12322,N_9666,N_8199);
nor U12323 (N_12323,N_6570,N_5348);
nor U12324 (N_12324,N_6837,N_9844);
and U12325 (N_12325,N_7034,N_6755);
or U12326 (N_12326,N_5615,N_9371);
or U12327 (N_12327,N_9107,N_5859);
nand U12328 (N_12328,N_5371,N_8322);
nand U12329 (N_12329,N_5943,N_7717);
nand U12330 (N_12330,N_7457,N_8484);
nor U12331 (N_12331,N_6082,N_6634);
or U12332 (N_12332,N_8171,N_9485);
or U12333 (N_12333,N_5798,N_8759);
and U12334 (N_12334,N_5471,N_9879);
or U12335 (N_12335,N_6602,N_6457);
nand U12336 (N_12336,N_9169,N_9245);
or U12337 (N_12337,N_8802,N_9830);
and U12338 (N_12338,N_6026,N_7965);
and U12339 (N_12339,N_8555,N_5004);
nand U12340 (N_12340,N_7493,N_8252);
or U12341 (N_12341,N_9220,N_8026);
nand U12342 (N_12342,N_6587,N_6780);
and U12343 (N_12343,N_7389,N_6567);
and U12344 (N_12344,N_8970,N_5230);
xnor U12345 (N_12345,N_6765,N_7485);
and U12346 (N_12346,N_8912,N_7384);
and U12347 (N_12347,N_9918,N_6061);
and U12348 (N_12348,N_6373,N_9353);
xnor U12349 (N_12349,N_5659,N_7628);
nor U12350 (N_12350,N_9849,N_6327);
nand U12351 (N_12351,N_6481,N_6699);
or U12352 (N_12352,N_7120,N_9940);
nand U12353 (N_12353,N_6442,N_5647);
and U12354 (N_12354,N_7599,N_9627);
or U12355 (N_12355,N_7905,N_5486);
or U12356 (N_12356,N_7270,N_6315);
nor U12357 (N_12357,N_6968,N_6415);
nor U12358 (N_12358,N_5565,N_5077);
nand U12359 (N_12359,N_7300,N_9311);
nand U12360 (N_12360,N_6243,N_9425);
or U12361 (N_12361,N_7785,N_5102);
or U12362 (N_12362,N_5621,N_5322);
nor U12363 (N_12363,N_8282,N_7446);
nand U12364 (N_12364,N_5571,N_7461);
or U12365 (N_12365,N_8057,N_5689);
or U12366 (N_12366,N_8763,N_6110);
nor U12367 (N_12367,N_9387,N_5409);
and U12368 (N_12368,N_7008,N_7156);
nand U12369 (N_12369,N_5682,N_6652);
or U12370 (N_12370,N_5049,N_7084);
nand U12371 (N_12371,N_7557,N_9677);
xor U12372 (N_12372,N_6927,N_7943);
nand U12373 (N_12373,N_6296,N_5796);
and U12374 (N_12374,N_9933,N_6757);
nand U12375 (N_12375,N_9416,N_9795);
and U12376 (N_12376,N_9582,N_9251);
and U12377 (N_12377,N_6254,N_9741);
nor U12378 (N_12378,N_5616,N_9069);
and U12379 (N_12379,N_9384,N_5591);
nor U12380 (N_12380,N_8261,N_8782);
or U12381 (N_12381,N_8922,N_8060);
or U12382 (N_12382,N_5294,N_5661);
nor U12383 (N_12383,N_5582,N_7125);
xor U12384 (N_12384,N_8196,N_9837);
xor U12385 (N_12385,N_5046,N_6419);
nor U12386 (N_12386,N_9430,N_9048);
and U12387 (N_12387,N_6245,N_6303);
and U12388 (N_12388,N_8958,N_6017);
or U12389 (N_12389,N_5170,N_9346);
nand U12390 (N_12390,N_9291,N_7433);
and U12391 (N_12391,N_7176,N_6053);
nand U12392 (N_12392,N_6371,N_7392);
xnor U12393 (N_12393,N_7762,N_8729);
and U12394 (N_12394,N_5039,N_6582);
and U12395 (N_12395,N_8237,N_8217);
or U12396 (N_12396,N_7696,N_5806);
nor U12397 (N_12397,N_7014,N_8214);
and U12398 (N_12398,N_6553,N_5632);
and U12399 (N_12399,N_6512,N_8405);
nor U12400 (N_12400,N_7750,N_7247);
nor U12401 (N_12401,N_8025,N_6905);
nand U12402 (N_12402,N_6401,N_8140);
or U12403 (N_12403,N_5250,N_6605);
or U12404 (N_12404,N_5345,N_8831);
xor U12405 (N_12405,N_9634,N_6641);
or U12406 (N_12406,N_7031,N_9388);
nand U12407 (N_12407,N_5701,N_8403);
or U12408 (N_12408,N_7510,N_7963);
nor U12409 (N_12409,N_5704,N_6501);
xor U12410 (N_12410,N_5922,N_8208);
nand U12411 (N_12411,N_7382,N_9661);
nor U12412 (N_12412,N_5153,N_9886);
nand U12413 (N_12413,N_9491,N_7719);
and U12414 (N_12414,N_9002,N_7085);
and U12415 (N_12415,N_7816,N_9655);
nor U12416 (N_12416,N_5699,N_9089);
nand U12417 (N_12417,N_9178,N_9495);
or U12418 (N_12418,N_6911,N_8930);
nor U12419 (N_12419,N_7307,N_8630);
nor U12420 (N_12420,N_7706,N_6682);
or U12421 (N_12421,N_7321,N_9958);
or U12422 (N_12422,N_5833,N_5807);
nor U12423 (N_12423,N_6182,N_6350);
and U12424 (N_12424,N_6362,N_9304);
and U12425 (N_12425,N_7890,N_8538);
and U12426 (N_12426,N_8852,N_8019);
nor U12427 (N_12427,N_7744,N_5340);
nand U12428 (N_12428,N_9917,N_9833);
xnor U12429 (N_12429,N_5008,N_9639);
or U12430 (N_12430,N_8951,N_6657);
nor U12431 (N_12431,N_9478,N_9147);
nand U12432 (N_12432,N_6311,N_7679);
xor U12433 (N_12433,N_6409,N_6840);
or U12434 (N_12434,N_5372,N_5337);
nand U12435 (N_12435,N_7749,N_7279);
and U12436 (N_12436,N_6330,N_9665);
xnor U12437 (N_12437,N_8806,N_5856);
or U12438 (N_12438,N_5145,N_5490);
nor U12439 (N_12439,N_5800,N_9679);
nor U12440 (N_12440,N_7091,N_5375);
xnor U12441 (N_12441,N_7549,N_8757);
and U12442 (N_12442,N_8258,N_8183);
or U12443 (N_12443,N_9971,N_6068);
nor U12444 (N_12444,N_9575,N_8871);
xor U12445 (N_12445,N_7320,N_5323);
xnor U12446 (N_12446,N_8931,N_6950);
and U12447 (N_12447,N_6152,N_5062);
nand U12448 (N_12448,N_5192,N_8522);
nand U12449 (N_12449,N_6817,N_6156);
and U12450 (N_12450,N_9307,N_7903);
and U12451 (N_12451,N_9034,N_7103);
or U12452 (N_12452,N_6281,N_5594);
nor U12453 (N_12453,N_9754,N_7655);
or U12454 (N_12454,N_5438,N_6475);
and U12455 (N_12455,N_5167,N_5086);
nor U12456 (N_12456,N_8587,N_8627);
and U12457 (N_12457,N_6483,N_6294);
or U12458 (N_12458,N_8093,N_6374);
and U12459 (N_12459,N_7026,N_9572);
or U12460 (N_12460,N_8506,N_6661);
nand U12461 (N_12461,N_6756,N_9158);
and U12462 (N_12462,N_7102,N_8756);
and U12463 (N_12463,N_6539,N_7068);
or U12464 (N_12464,N_5195,N_9136);
nor U12465 (N_12465,N_7975,N_9135);
and U12466 (N_12466,N_8916,N_7941);
and U12467 (N_12467,N_7733,N_6403);
nor U12468 (N_12468,N_7143,N_6721);
or U12469 (N_12469,N_5907,N_5023);
xnor U12470 (N_12470,N_7769,N_6734);
nand U12471 (N_12471,N_7636,N_7888);
nor U12472 (N_12472,N_6040,N_6883);
nand U12473 (N_12473,N_5207,N_7828);
and U12474 (N_12474,N_5570,N_8112);
nor U12475 (N_12475,N_5550,N_8987);
nand U12476 (N_12476,N_6811,N_7922);
and U12477 (N_12477,N_7194,N_6031);
xor U12478 (N_12478,N_7403,N_5897);
xnor U12479 (N_12479,N_7104,N_5793);
and U12480 (N_12480,N_5157,N_7228);
and U12481 (N_12481,N_9265,N_9994);
nor U12482 (N_12482,N_7340,N_8313);
and U12483 (N_12483,N_9534,N_8638);
and U12484 (N_12484,N_5977,N_5048);
nor U12485 (N_12485,N_7781,N_9161);
or U12486 (N_12486,N_8937,N_6679);
and U12487 (N_12487,N_8200,N_7266);
and U12488 (N_12488,N_7932,N_8939);
nor U12489 (N_12489,N_5278,N_9361);
nand U12490 (N_12490,N_7887,N_5750);
nor U12491 (N_12491,N_5653,N_7399);
nand U12492 (N_12492,N_8223,N_5053);
or U12493 (N_12493,N_7222,N_5436);
nor U12494 (N_12494,N_9472,N_6568);
nor U12495 (N_12495,N_8928,N_5817);
or U12496 (N_12496,N_7942,N_9296);
nor U12497 (N_12497,N_8197,N_6007);
nand U12498 (N_12498,N_7645,N_8779);
nor U12499 (N_12499,N_5017,N_7347);
and U12500 (N_12500,N_6141,N_9114);
or U12501 (N_12501,N_9200,N_7748);
nand U12502 (N_12502,N_7331,N_8975);
and U12503 (N_12503,N_8731,N_9271);
or U12504 (N_12504,N_5705,N_5490);
or U12505 (N_12505,N_7553,N_9683);
xnor U12506 (N_12506,N_5207,N_5754);
nand U12507 (N_12507,N_8896,N_9652);
xnor U12508 (N_12508,N_8457,N_8925);
or U12509 (N_12509,N_7698,N_6674);
nor U12510 (N_12510,N_8026,N_9052);
xor U12511 (N_12511,N_7601,N_5781);
xor U12512 (N_12512,N_7594,N_6042);
nand U12513 (N_12513,N_8846,N_7157);
nor U12514 (N_12514,N_6884,N_7214);
or U12515 (N_12515,N_8658,N_6634);
and U12516 (N_12516,N_6215,N_5967);
nand U12517 (N_12517,N_5381,N_9830);
and U12518 (N_12518,N_6152,N_7805);
or U12519 (N_12519,N_9214,N_5008);
and U12520 (N_12520,N_8566,N_9591);
or U12521 (N_12521,N_9103,N_9372);
and U12522 (N_12522,N_6595,N_8484);
nand U12523 (N_12523,N_6349,N_9502);
and U12524 (N_12524,N_7787,N_7095);
or U12525 (N_12525,N_8403,N_8937);
xnor U12526 (N_12526,N_5456,N_8854);
nor U12527 (N_12527,N_8190,N_7104);
or U12528 (N_12528,N_6083,N_9566);
or U12529 (N_12529,N_8571,N_9632);
nand U12530 (N_12530,N_7036,N_7985);
or U12531 (N_12531,N_6774,N_7436);
xor U12532 (N_12532,N_8385,N_7178);
and U12533 (N_12533,N_7920,N_5264);
nor U12534 (N_12534,N_6797,N_9966);
and U12535 (N_12535,N_5546,N_6797);
and U12536 (N_12536,N_6210,N_7347);
xor U12537 (N_12537,N_6873,N_7222);
and U12538 (N_12538,N_7843,N_9914);
or U12539 (N_12539,N_6378,N_9926);
or U12540 (N_12540,N_7089,N_6207);
nor U12541 (N_12541,N_5739,N_8940);
or U12542 (N_12542,N_5017,N_6392);
nor U12543 (N_12543,N_5160,N_5581);
nor U12544 (N_12544,N_7086,N_6093);
nor U12545 (N_12545,N_9036,N_5216);
nand U12546 (N_12546,N_6062,N_7475);
and U12547 (N_12547,N_7056,N_8714);
xnor U12548 (N_12548,N_8955,N_7800);
or U12549 (N_12549,N_7367,N_7885);
nor U12550 (N_12550,N_8540,N_6920);
nor U12551 (N_12551,N_5151,N_6838);
and U12552 (N_12552,N_5700,N_6131);
nand U12553 (N_12553,N_8668,N_6818);
and U12554 (N_12554,N_8812,N_5046);
xor U12555 (N_12555,N_6263,N_9910);
and U12556 (N_12556,N_5995,N_7883);
and U12557 (N_12557,N_6390,N_5332);
nor U12558 (N_12558,N_5475,N_6072);
or U12559 (N_12559,N_7783,N_7957);
and U12560 (N_12560,N_9875,N_7622);
and U12561 (N_12561,N_5859,N_9754);
nor U12562 (N_12562,N_6540,N_6824);
or U12563 (N_12563,N_9709,N_7925);
and U12564 (N_12564,N_6881,N_7733);
xnor U12565 (N_12565,N_6706,N_8955);
nor U12566 (N_12566,N_8880,N_6683);
or U12567 (N_12567,N_9884,N_5475);
or U12568 (N_12568,N_5970,N_7084);
nand U12569 (N_12569,N_5285,N_7858);
or U12570 (N_12570,N_8108,N_6438);
xor U12571 (N_12571,N_5178,N_9300);
and U12572 (N_12572,N_6970,N_5203);
or U12573 (N_12573,N_7067,N_5870);
nand U12574 (N_12574,N_9111,N_6670);
and U12575 (N_12575,N_7528,N_7320);
nand U12576 (N_12576,N_8494,N_7998);
nand U12577 (N_12577,N_6696,N_6160);
nand U12578 (N_12578,N_9906,N_7643);
nand U12579 (N_12579,N_5522,N_9617);
nor U12580 (N_12580,N_9724,N_5577);
and U12581 (N_12581,N_5653,N_9658);
nor U12582 (N_12582,N_6793,N_8123);
or U12583 (N_12583,N_5208,N_7156);
or U12584 (N_12584,N_7396,N_8341);
nand U12585 (N_12585,N_8271,N_7281);
nor U12586 (N_12586,N_8776,N_8911);
xnor U12587 (N_12587,N_5017,N_6514);
or U12588 (N_12588,N_6126,N_7891);
and U12589 (N_12589,N_5422,N_8941);
xor U12590 (N_12590,N_5848,N_6383);
nor U12591 (N_12591,N_8295,N_7126);
nor U12592 (N_12592,N_8221,N_5542);
and U12593 (N_12593,N_7513,N_7029);
or U12594 (N_12594,N_8934,N_9098);
and U12595 (N_12595,N_7615,N_5278);
nand U12596 (N_12596,N_8567,N_9250);
and U12597 (N_12597,N_7626,N_7863);
or U12598 (N_12598,N_8084,N_7141);
nor U12599 (N_12599,N_5489,N_8177);
or U12600 (N_12600,N_9134,N_7030);
or U12601 (N_12601,N_5209,N_7209);
or U12602 (N_12602,N_8882,N_6754);
nor U12603 (N_12603,N_9298,N_7574);
nand U12604 (N_12604,N_9209,N_8511);
nand U12605 (N_12605,N_7268,N_9998);
nor U12606 (N_12606,N_7468,N_5944);
nor U12607 (N_12607,N_6775,N_6418);
or U12608 (N_12608,N_8251,N_9610);
xor U12609 (N_12609,N_6976,N_8121);
nand U12610 (N_12610,N_8476,N_9826);
nor U12611 (N_12611,N_8994,N_9444);
or U12612 (N_12612,N_9994,N_5913);
nand U12613 (N_12613,N_8637,N_7048);
nand U12614 (N_12614,N_5602,N_9298);
and U12615 (N_12615,N_9844,N_7781);
nand U12616 (N_12616,N_7478,N_5035);
and U12617 (N_12617,N_8475,N_6579);
and U12618 (N_12618,N_7995,N_7900);
xor U12619 (N_12619,N_9410,N_7490);
or U12620 (N_12620,N_6706,N_7118);
xnor U12621 (N_12621,N_7226,N_9534);
or U12622 (N_12622,N_7244,N_8754);
nor U12623 (N_12623,N_6433,N_5187);
and U12624 (N_12624,N_9277,N_7737);
xor U12625 (N_12625,N_5864,N_7589);
or U12626 (N_12626,N_9353,N_8222);
nand U12627 (N_12627,N_7659,N_6178);
or U12628 (N_12628,N_5595,N_6681);
and U12629 (N_12629,N_8540,N_5897);
xor U12630 (N_12630,N_8014,N_9603);
or U12631 (N_12631,N_9575,N_8047);
or U12632 (N_12632,N_7024,N_8202);
nand U12633 (N_12633,N_6305,N_9272);
nand U12634 (N_12634,N_6046,N_6760);
or U12635 (N_12635,N_8719,N_6064);
or U12636 (N_12636,N_5088,N_9575);
xnor U12637 (N_12637,N_9636,N_6071);
and U12638 (N_12638,N_6599,N_9758);
nand U12639 (N_12639,N_9150,N_9238);
nor U12640 (N_12640,N_7758,N_6551);
nor U12641 (N_12641,N_6353,N_6857);
xor U12642 (N_12642,N_5722,N_9204);
xnor U12643 (N_12643,N_5726,N_7863);
or U12644 (N_12644,N_6426,N_5670);
or U12645 (N_12645,N_8343,N_8101);
nor U12646 (N_12646,N_7661,N_8859);
and U12647 (N_12647,N_8438,N_7046);
and U12648 (N_12648,N_6343,N_6787);
nand U12649 (N_12649,N_7501,N_5758);
nor U12650 (N_12650,N_9211,N_7824);
nand U12651 (N_12651,N_9857,N_9738);
nand U12652 (N_12652,N_6844,N_8997);
nor U12653 (N_12653,N_9619,N_7094);
or U12654 (N_12654,N_7911,N_6926);
nand U12655 (N_12655,N_7645,N_6644);
and U12656 (N_12656,N_5165,N_9730);
and U12657 (N_12657,N_6658,N_7204);
nor U12658 (N_12658,N_6755,N_6974);
or U12659 (N_12659,N_5958,N_5561);
nand U12660 (N_12660,N_8320,N_5787);
nand U12661 (N_12661,N_7024,N_6239);
xnor U12662 (N_12662,N_5827,N_6952);
nand U12663 (N_12663,N_6559,N_8953);
xor U12664 (N_12664,N_9390,N_7362);
and U12665 (N_12665,N_7920,N_8330);
nand U12666 (N_12666,N_7630,N_5017);
and U12667 (N_12667,N_6403,N_6537);
and U12668 (N_12668,N_7006,N_9039);
nand U12669 (N_12669,N_6183,N_7294);
and U12670 (N_12670,N_5818,N_9838);
or U12671 (N_12671,N_6638,N_8643);
nand U12672 (N_12672,N_7468,N_9057);
nand U12673 (N_12673,N_8740,N_5395);
and U12674 (N_12674,N_8031,N_6206);
nand U12675 (N_12675,N_9432,N_9531);
or U12676 (N_12676,N_8436,N_9500);
nor U12677 (N_12677,N_7669,N_5107);
and U12678 (N_12678,N_6296,N_8148);
or U12679 (N_12679,N_7159,N_8219);
nor U12680 (N_12680,N_9794,N_9117);
xnor U12681 (N_12681,N_7149,N_7448);
nor U12682 (N_12682,N_8204,N_9449);
or U12683 (N_12683,N_8450,N_5973);
nand U12684 (N_12684,N_5113,N_6508);
nand U12685 (N_12685,N_8104,N_6612);
nor U12686 (N_12686,N_7203,N_6645);
and U12687 (N_12687,N_8028,N_8188);
nor U12688 (N_12688,N_5197,N_6167);
and U12689 (N_12689,N_6404,N_8003);
and U12690 (N_12690,N_6182,N_6577);
nor U12691 (N_12691,N_6892,N_9348);
or U12692 (N_12692,N_9080,N_9588);
nor U12693 (N_12693,N_5793,N_8593);
nand U12694 (N_12694,N_8553,N_9942);
nand U12695 (N_12695,N_6354,N_8307);
or U12696 (N_12696,N_7536,N_5187);
nor U12697 (N_12697,N_7089,N_6659);
or U12698 (N_12698,N_8612,N_5922);
or U12699 (N_12699,N_7564,N_6180);
and U12700 (N_12700,N_7743,N_5786);
nand U12701 (N_12701,N_9448,N_7806);
and U12702 (N_12702,N_6155,N_8062);
and U12703 (N_12703,N_5374,N_5672);
or U12704 (N_12704,N_6830,N_7868);
or U12705 (N_12705,N_8412,N_6491);
or U12706 (N_12706,N_6935,N_7722);
or U12707 (N_12707,N_6204,N_9970);
or U12708 (N_12708,N_6725,N_9358);
nand U12709 (N_12709,N_7190,N_8808);
nand U12710 (N_12710,N_6279,N_7961);
xor U12711 (N_12711,N_5878,N_9298);
or U12712 (N_12712,N_8052,N_7516);
nor U12713 (N_12713,N_9528,N_6695);
or U12714 (N_12714,N_6652,N_5768);
xor U12715 (N_12715,N_6166,N_5572);
or U12716 (N_12716,N_9093,N_8636);
nor U12717 (N_12717,N_5937,N_7943);
and U12718 (N_12718,N_8397,N_6467);
and U12719 (N_12719,N_5974,N_9039);
or U12720 (N_12720,N_9777,N_6441);
and U12721 (N_12721,N_9726,N_6506);
nor U12722 (N_12722,N_6953,N_6276);
nor U12723 (N_12723,N_7705,N_6519);
or U12724 (N_12724,N_5700,N_9051);
or U12725 (N_12725,N_5649,N_8254);
nor U12726 (N_12726,N_7114,N_9864);
xor U12727 (N_12727,N_5578,N_7059);
and U12728 (N_12728,N_6571,N_7171);
or U12729 (N_12729,N_5894,N_8025);
or U12730 (N_12730,N_8337,N_8913);
nor U12731 (N_12731,N_6378,N_7110);
nor U12732 (N_12732,N_9870,N_8963);
nor U12733 (N_12733,N_5863,N_7246);
and U12734 (N_12734,N_6705,N_7587);
and U12735 (N_12735,N_6068,N_8832);
nand U12736 (N_12736,N_7182,N_7593);
nand U12737 (N_12737,N_8172,N_5026);
nand U12738 (N_12738,N_9625,N_6580);
or U12739 (N_12739,N_6649,N_9340);
nor U12740 (N_12740,N_6443,N_7591);
nor U12741 (N_12741,N_9332,N_7608);
and U12742 (N_12742,N_7076,N_8638);
nand U12743 (N_12743,N_5230,N_5774);
and U12744 (N_12744,N_8392,N_5683);
and U12745 (N_12745,N_5754,N_9563);
or U12746 (N_12746,N_7908,N_6500);
or U12747 (N_12747,N_6184,N_8871);
and U12748 (N_12748,N_6890,N_8846);
and U12749 (N_12749,N_7803,N_5614);
xnor U12750 (N_12750,N_9600,N_8999);
nand U12751 (N_12751,N_9454,N_7974);
nand U12752 (N_12752,N_9468,N_9721);
nor U12753 (N_12753,N_5685,N_7766);
or U12754 (N_12754,N_9422,N_5797);
nor U12755 (N_12755,N_9300,N_6292);
and U12756 (N_12756,N_5256,N_5364);
and U12757 (N_12757,N_6682,N_6054);
and U12758 (N_12758,N_8256,N_8000);
nor U12759 (N_12759,N_5084,N_5231);
and U12760 (N_12760,N_5547,N_8251);
nand U12761 (N_12761,N_6362,N_9201);
xnor U12762 (N_12762,N_9650,N_8179);
and U12763 (N_12763,N_5061,N_6907);
or U12764 (N_12764,N_5250,N_8679);
or U12765 (N_12765,N_6166,N_9844);
nor U12766 (N_12766,N_8916,N_5157);
xnor U12767 (N_12767,N_8005,N_8057);
or U12768 (N_12768,N_6958,N_5243);
or U12769 (N_12769,N_5057,N_6923);
nor U12770 (N_12770,N_7488,N_9359);
or U12771 (N_12771,N_9439,N_9004);
nand U12772 (N_12772,N_8484,N_5473);
xnor U12773 (N_12773,N_7941,N_7048);
nor U12774 (N_12774,N_7169,N_9583);
and U12775 (N_12775,N_6158,N_5375);
nor U12776 (N_12776,N_8625,N_8757);
nor U12777 (N_12777,N_6917,N_7677);
or U12778 (N_12778,N_5039,N_8407);
and U12779 (N_12779,N_8049,N_7168);
and U12780 (N_12780,N_9539,N_8562);
nand U12781 (N_12781,N_9987,N_8874);
xnor U12782 (N_12782,N_6656,N_9832);
and U12783 (N_12783,N_8465,N_8737);
xnor U12784 (N_12784,N_8151,N_9846);
xnor U12785 (N_12785,N_9535,N_5216);
or U12786 (N_12786,N_7501,N_8397);
or U12787 (N_12787,N_9407,N_7472);
nor U12788 (N_12788,N_5349,N_6964);
nor U12789 (N_12789,N_8318,N_6425);
or U12790 (N_12790,N_8211,N_6389);
and U12791 (N_12791,N_7889,N_9743);
nor U12792 (N_12792,N_6224,N_6206);
and U12793 (N_12793,N_8524,N_7124);
xor U12794 (N_12794,N_6827,N_8713);
or U12795 (N_12795,N_9192,N_9391);
nand U12796 (N_12796,N_7412,N_5697);
or U12797 (N_12797,N_7802,N_8758);
nand U12798 (N_12798,N_7957,N_5465);
nand U12799 (N_12799,N_7034,N_6539);
or U12800 (N_12800,N_7956,N_9997);
and U12801 (N_12801,N_8978,N_7207);
nand U12802 (N_12802,N_9507,N_5687);
nor U12803 (N_12803,N_7261,N_7457);
and U12804 (N_12804,N_9049,N_8930);
or U12805 (N_12805,N_7285,N_9673);
nand U12806 (N_12806,N_9065,N_6385);
nand U12807 (N_12807,N_6313,N_9244);
or U12808 (N_12808,N_5268,N_5738);
or U12809 (N_12809,N_7800,N_5370);
and U12810 (N_12810,N_7235,N_9606);
and U12811 (N_12811,N_6775,N_7862);
nand U12812 (N_12812,N_6316,N_7248);
and U12813 (N_12813,N_7172,N_7173);
or U12814 (N_12814,N_6797,N_6233);
nand U12815 (N_12815,N_5505,N_6156);
nand U12816 (N_12816,N_7840,N_8577);
nor U12817 (N_12817,N_6025,N_7251);
nor U12818 (N_12818,N_6907,N_7551);
and U12819 (N_12819,N_8301,N_8095);
or U12820 (N_12820,N_7461,N_6970);
xor U12821 (N_12821,N_6551,N_9393);
nor U12822 (N_12822,N_7543,N_5415);
and U12823 (N_12823,N_6753,N_9189);
nor U12824 (N_12824,N_7251,N_5764);
or U12825 (N_12825,N_5483,N_5436);
nand U12826 (N_12826,N_8663,N_6338);
or U12827 (N_12827,N_7450,N_8457);
and U12828 (N_12828,N_8029,N_5185);
nand U12829 (N_12829,N_5203,N_6721);
nor U12830 (N_12830,N_8175,N_8282);
and U12831 (N_12831,N_9035,N_6115);
xnor U12832 (N_12832,N_9204,N_9175);
nand U12833 (N_12833,N_5864,N_7819);
xnor U12834 (N_12834,N_8337,N_7578);
and U12835 (N_12835,N_8172,N_6520);
xor U12836 (N_12836,N_9537,N_9117);
and U12837 (N_12837,N_7028,N_6862);
or U12838 (N_12838,N_6898,N_5276);
nor U12839 (N_12839,N_9044,N_7727);
nand U12840 (N_12840,N_7340,N_6698);
nor U12841 (N_12841,N_8467,N_5238);
nand U12842 (N_12842,N_7246,N_8254);
and U12843 (N_12843,N_5777,N_7351);
nand U12844 (N_12844,N_6259,N_9764);
nor U12845 (N_12845,N_8231,N_8136);
or U12846 (N_12846,N_7621,N_7111);
or U12847 (N_12847,N_7441,N_7645);
or U12848 (N_12848,N_9594,N_6111);
nand U12849 (N_12849,N_5696,N_8898);
nor U12850 (N_12850,N_8173,N_7235);
or U12851 (N_12851,N_9271,N_5093);
and U12852 (N_12852,N_8263,N_9291);
nand U12853 (N_12853,N_5204,N_9430);
nand U12854 (N_12854,N_7402,N_6367);
xnor U12855 (N_12855,N_7721,N_5605);
nand U12856 (N_12856,N_6510,N_8608);
nand U12857 (N_12857,N_8542,N_7713);
nor U12858 (N_12858,N_5181,N_5123);
nand U12859 (N_12859,N_6498,N_5725);
nand U12860 (N_12860,N_5696,N_7600);
nor U12861 (N_12861,N_6280,N_8219);
or U12862 (N_12862,N_5082,N_7349);
and U12863 (N_12863,N_6035,N_7672);
nand U12864 (N_12864,N_9266,N_6136);
xor U12865 (N_12865,N_8320,N_9455);
or U12866 (N_12866,N_5116,N_6307);
nand U12867 (N_12867,N_7157,N_5017);
nor U12868 (N_12868,N_8067,N_6055);
nor U12869 (N_12869,N_8085,N_9235);
xnor U12870 (N_12870,N_5055,N_9610);
nor U12871 (N_12871,N_6971,N_7052);
or U12872 (N_12872,N_8216,N_7877);
and U12873 (N_12873,N_7303,N_7614);
nor U12874 (N_12874,N_6266,N_8802);
nor U12875 (N_12875,N_5156,N_8606);
nand U12876 (N_12876,N_6299,N_5853);
nand U12877 (N_12877,N_9943,N_5381);
and U12878 (N_12878,N_8606,N_9343);
and U12879 (N_12879,N_9572,N_6417);
nor U12880 (N_12880,N_8400,N_5157);
or U12881 (N_12881,N_9460,N_8028);
nand U12882 (N_12882,N_8378,N_6183);
or U12883 (N_12883,N_8643,N_8036);
nor U12884 (N_12884,N_7220,N_5056);
nor U12885 (N_12885,N_7985,N_6195);
nor U12886 (N_12886,N_7423,N_9558);
and U12887 (N_12887,N_9308,N_5736);
nor U12888 (N_12888,N_8023,N_9817);
or U12889 (N_12889,N_5650,N_7419);
nor U12890 (N_12890,N_5282,N_7144);
nor U12891 (N_12891,N_9029,N_5973);
and U12892 (N_12892,N_8732,N_5048);
and U12893 (N_12893,N_7421,N_8565);
nand U12894 (N_12894,N_8779,N_7709);
or U12895 (N_12895,N_9135,N_8546);
and U12896 (N_12896,N_5021,N_8039);
and U12897 (N_12897,N_6734,N_8182);
xnor U12898 (N_12898,N_5559,N_6791);
nand U12899 (N_12899,N_8244,N_6786);
and U12900 (N_12900,N_7995,N_5846);
or U12901 (N_12901,N_8513,N_6548);
nand U12902 (N_12902,N_7280,N_5728);
and U12903 (N_12903,N_9408,N_6555);
and U12904 (N_12904,N_8914,N_7655);
nor U12905 (N_12905,N_8399,N_7769);
or U12906 (N_12906,N_9007,N_5495);
and U12907 (N_12907,N_9238,N_6415);
nand U12908 (N_12908,N_8825,N_8786);
or U12909 (N_12909,N_8764,N_8468);
nand U12910 (N_12910,N_5296,N_6585);
xnor U12911 (N_12911,N_8721,N_8907);
nor U12912 (N_12912,N_5403,N_7363);
nand U12913 (N_12913,N_9792,N_5439);
nor U12914 (N_12914,N_7285,N_7326);
nand U12915 (N_12915,N_7647,N_8908);
or U12916 (N_12916,N_5748,N_8631);
or U12917 (N_12917,N_5121,N_6419);
nand U12918 (N_12918,N_6891,N_9994);
and U12919 (N_12919,N_6274,N_6639);
or U12920 (N_12920,N_8352,N_7194);
nand U12921 (N_12921,N_7108,N_8049);
nand U12922 (N_12922,N_6131,N_6558);
xor U12923 (N_12923,N_5684,N_5512);
nor U12924 (N_12924,N_8792,N_6570);
and U12925 (N_12925,N_7385,N_7811);
nand U12926 (N_12926,N_5644,N_7939);
nor U12927 (N_12927,N_7451,N_6341);
or U12928 (N_12928,N_7885,N_7125);
nand U12929 (N_12929,N_7620,N_7327);
nor U12930 (N_12930,N_8264,N_6154);
and U12931 (N_12931,N_7706,N_5633);
nor U12932 (N_12932,N_5274,N_7760);
nor U12933 (N_12933,N_6291,N_6702);
nand U12934 (N_12934,N_6572,N_7841);
xor U12935 (N_12935,N_5260,N_8098);
and U12936 (N_12936,N_8124,N_6183);
and U12937 (N_12937,N_5252,N_9813);
nor U12938 (N_12938,N_9592,N_5634);
or U12939 (N_12939,N_7237,N_6537);
and U12940 (N_12940,N_9207,N_8248);
and U12941 (N_12941,N_5210,N_5782);
and U12942 (N_12942,N_8210,N_7567);
nor U12943 (N_12943,N_7367,N_9260);
xor U12944 (N_12944,N_7636,N_6553);
or U12945 (N_12945,N_8159,N_8977);
or U12946 (N_12946,N_6904,N_5472);
or U12947 (N_12947,N_9065,N_9347);
or U12948 (N_12948,N_5939,N_6780);
nor U12949 (N_12949,N_7669,N_7735);
nor U12950 (N_12950,N_7910,N_8502);
xnor U12951 (N_12951,N_5826,N_6509);
nand U12952 (N_12952,N_6976,N_5788);
xor U12953 (N_12953,N_5766,N_9584);
and U12954 (N_12954,N_9649,N_9644);
and U12955 (N_12955,N_9683,N_9177);
and U12956 (N_12956,N_6028,N_5842);
nor U12957 (N_12957,N_8831,N_7388);
nand U12958 (N_12958,N_7028,N_5051);
nor U12959 (N_12959,N_9734,N_6024);
and U12960 (N_12960,N_7145,N_7531);
or U12961 (N_12961,N_7466,N_9996);
nor U12962 (N_12962,N_8133,N_7814);
nand U12963 (N_12963,N_7985,N_8696);
and U12964 (N_12964,N_5487,N_6102);
nor U12965 (N_12965,N_9430,N_6632);
nand U12966 (N_12966,N_8585,N_5558);
nor U12967 (N_12967,N_9060,N_6174);
nand U12968 (N_12968,N_6128,N_6966);
and U12969 (N_12969,N_5139,N_5744);
nand U12970 (N_12970,N_6082,N_7175);
nand U12971 (N_12971,N_8037,N_7879);
nor U12972 (N_12972,N_6550,N_8406);
and U12973 (N_12973,N_5879,N_9060);
nand U12974 (N_12974,N_8562,N_5668);
nand U12975 (N_12975,N_7189,N_7104);
xor U12976 (N_12976,N_9286,N_5976);
nand U12977 (N_12977,N_7320,N_7584);
nor U12978 (N_12978,N_8855,N_6291);
nor U12979 (N_12979,N_8641,N_9080);
and U12980 (N_12980,N_5796,N_8692);
or U12981 (N_12981,N_9713,N_7892);
and U12982 (N_12982,N_7212,N_7962);
xnor U12983 (N_12983,N_6237,N_7264);
nand U12984 (N_12984,N_5206,N_7195);
nor U12985 (N_12985,N_5602,N_8466);
nor U12986 (N_12986,N_6395,N_7719);
or U12987 (N_12987,N_9665,N_6430);
nand U12988 (N_12988,N_8789,N_8515);
nor U12989 (N_12989,N_6017,N_8208);
nor U12990 (N_12990,N_8340,N_9445);
nor U12991 (N_12991,N_9132,N_7440);
or U12992 (N_12992,N_7924,N_8521);
nor U12993 (N_12993,N_5082,N_6326);
or U12994 (N_12994,N_7252,N_5015);
and U12995 (N_12995,N_7858,N_7227);
or U12996 (N_12996,N_6566,N_6257);
xor U12997 (N_12997,N_8568,N_7924);
nor U12998 (N_12998,N_8984,N_8643);
nand U12999 (N_12999,N_9038,N_8527);
or U13000 (N_13000,N_6835,N_6784);
nand U13001 (N_13001,N_5118,N_7620);
nand U13002 (N_13002,N_9785,N_9750);
nand U13003 (N_13003,N_5052,N_7455);
nand U13004 (N_13004,N_5061,N_5100);
and U13005 (N_13005,N_5132,N_6778);
nand U13006 (N_13006,N_7228,N_7644);
or U13007 (N_13007,N_5355,N_6747);
xnor U13008 (N_13008,N_9545,N_9277);
nand U13009 (N_13009,N_6630,N_9829);
and U13010 (N_13010,N_9547,N_9985);
xor U13011 (N_13011,N_9367,N_6293);
nand U13012 (N_13012,N_7695,N_6467);
and U13013 (N_13013,N_6533,N_5179);
xor U13014 (N_13014,N_5787,N_7684);
nor U13015 (N_13015,N_5165,N_8047);
or U13016 (N_13016,N_5117,N_6723);
or U13017 (N_13017,N_9539,N_9841);
or U13018 (N_13018,N_8498,N_5551);
xnor U13019 (N_13019,N_7032,N_6235);
and U13020 (N_13020,N_9821,N_5979);
xnor U13021 (N_13021,N_7930,N_5068);
nand U13022 (N_13022,N_5479,N_7231);
and U13023 (N_13023,N_7161,N_7748);
and U13024 (N_13024,N_8116,N_9782);
nor U13025 (N_13025,N_9746,N_6803);
and U13026 (N_13026,N_5592,N_8688);
and U13027 (N_13027,N_9526,N_7401);
nor U13028 (N_13028,N_6438,N_9696);
nand U13029 (N_13029,N_7440,N_7845);
nand U13030 (N_13030,N_8892,N_8358);
or U13031 (N_13031,N_7282,N_5337);
and U13032 (N_13032,N_5253,N_7484);
and U13033 (N_13033,N_6581,N_7358);
nor U13034 (N_13034,N_5652,N_8882);
xnor U13035 (N_13035,N_7391,N_9537);
and U13036 (N_13036,N_9304,N_9268);
nand U13037 (N_13037,N_8270,N_7879);
or U13038 (N_13038,N_6959,N_8368);
nor U13039 (N_13039,N_5914,N_8489);
nor U13040 (N_13040,N_5979,N_7098);
nor U13041 (N_13041,N_5197,N_6899);
xnor U13042 (N_13042,N_9010,N_9626);
and U13043 (N_13043,N_6511,N_5457);
nand U13044 (N_13044,N_5252,N_5066);
and U13045 (N_13045,N_6952,N_6413);
or U13046 (N_13046,N_7864,N_9330);
and U13047 (N_13047,N_9332,N_8270);
nand U13048 (N_13048,N_6489,N_6870);
nor U13049 (N_13049,N_6912,N_5510);
nand U13050 (N_13050,N_6247,N_8105);
or U13051 (N_13051,N_9847,N_7882);
xor U13052 (N_13052,N_6179,N_6502);
xnor U13053 (N_13053,N_5691,N_5801);
xnor U13054 (N_13054,N_9837,N_8335);
or U13055 (N_13055,N_6669,N_7169);
and U13056 (N_13056,N_8402,N_6180);
xnor U13057 (N_13057,N_8307,N_8451);
nand U13058 (N_13058,N_5303,N_7101);
or U13059 (N_13059,N_6671,N_7030);
xnor U13060 (N_13060,N_5992,N_6308);
xnor U13061 (N_13061,N_5582,N_9516);
and U13062 (N_13062,N_6608,N_6151);
nand U13063 (N_13063,N_9042,N_8405);
xor U13064 (N_13064,N_6001,N_9001);
or U13065 (N_13065,N_7659,N_5199);
xnor U13066 (N_13066,N_9193,N_9677);
or U13067 (N_13067,N_5802,N_5123);
nor U13068 (N_13068,N_5435,N_6422);
xor U13069 (N_13069,N_7342,N_8348);
or U13070 (N_13070,N_5803,N_6401);
nand U13071 (N_13071,N_5321,N_6046);
or U13072 (N_13072,N_7733,N_5083);
nor U13073 (N_13073,N_9814,N_8819);
nor U13074 (N_13074,N_8361,N_6957);
nand U13075 (N_13075,N_5476,N_7764);
and U13076 (N_13076,N_9150,N_6879);
and U13077 (N_13077,N_5320,N_7707);
or U13078 (N_13078,N_9703,N_5393);
nor U13079 (N_13079,N_7286,N_9532);
nor U13080 (N_13080,N_6568,N_6622);
or U13081 (N_13081,N_7188,N_5790);
nor U13082 (N_13082,N_9456,N_7764);
nand U13083 (N_13083,N_6415,N_7148);
and U13084 (N_13084,N_7429,N_8642);
nor U13085 (N_13085,N_7333,N_5496);
nor U13086 (N_13086,N_5202,N_9606);
or U13087 (N_13087,N_8345,N_6855);
and U13088 (N_13088,N_8453,N_5452);
nand U13089 (N_13089,N_6633,N_7801);
nor U13090 (N_13090,N_6386,N_9513);
xnor U13091 (N_13091,N_9757,N_8690);
and U13092 (N_13092,N_8457,N_6344);
or U13093 (N_13093,N_9296,N_6381);
or U13094 (N_13094,N_9879,N_9549);
or U13095 (N_13095,N_9700,N_7841);
or U13096 (N_13096,N_5708,N_8516);
and U13097 (N_13097,N_9266,N_5046);
xnor U13098 (N_13098,N_6014,N_6293);
or U13099 (N_13099,N_7406,N_7600);
and U13100 (N_13100,N_8103,N_8180);
or U13101 (N_13101,N_8029,N_9130);
and U13102 (N_13102,N_9932,N_5065);
nor U13103 (N_13103,N_6979,N_9700);
and U13104 (N_13104,N_8697,N_6159);
nand U13105 (N_13105,N_7314,N_8513);
nor U13106 (N_13106,N_9528,N_8207);
nand U13107 (N_13107,N_6064,N_6571);
and U13108 (N_13108,N_7461,N_7933);
nand U13109 (N_13109,N_8270,N_6068);
nand U13110 (N_13110,N_8621,N_6733);
or U13111 (N_13111,N_8614,N_8858);
nand U13112 (N_13112,N_8365,N_6168);
nand U13113 (N_13113,N_9372,N_6647);
nand U13114 (N_13114,N_9914,N_9962);
nand U13115 (N_13115,N_9701,N_8297);
nor U13116 (N_13116,N_8898,N_5586);
xnor U13117 (N_13117,N_9738,N_7015);
or U13118 (N_13118,N_7132,N_8410);
and U13119 (N_13119,N_7863,N_7909);
and U13120 (N_13120,N_8576,N_6045);
or U13121 (N_13121,N_6670,N_6162);
nand U13122 (N_13122,N_7034,N_9331);
and U13123 (N_13123,N_5878,N_5125);
xor U13124 (N_13124,N_5771,N_9893);
nor U13125 (N_13125,N_7503,N_8714);
nor U13126 (N_13126,N_6340,N_5429);
or U13127 (N_13127,N_8932,N_8457);
or U13128 (N_13128,N_6424,N_6467);
or U13129 (N_13129,N_9545,N_9604);
nor U13130 (N_13130,N_8718,N_7863);
or U13131 (N_13131,N_8477,N_7756);
and U13132 (N_13132,N_9226,N_6996);
and U13133 (N_13133,N_6316,N_5016);
nor U13134 (N_13134,N_5049,N_7999);
nor U13135 (N_13135,N_9691,N_9883);
and U13136 (N_13136,N_5656,N_7164);
or U13137 (N_13137,N_7445,N_7146);
and U13138 (N_13138,N_8456,N_5384);
nand U13139 (N_13139,N_9541,N_5762);
and U13140 (N_13140,N_5666,N_5345);
or U13141 (N_13141,N_5030,N_7891);
nand U13142 (N_13142,N_7615,N_9647);
nand U13143 (N_13143,N_6025,N_9198);
nor U13144 (N_13144,N_7629,N_6665);
nand U13145 (N_13145,N_8683,N_9270);
nand U13146 (N_13146,N_7649,N_6149);
nand U13147 (N_13147,N_5616,N_7402);
or U13148 (N_13148,N_7711,N_7581);
and U13149 (N_13149,N_9023,N_6737);
or U13150 (N_13150,N_5685,N_5281);
nand U13151 (N_13151,N_9133,N_5640);
and U13152 (N_13152,N_9928,N_6493);
nand U13153 (N_13153,N_5856,N_5569);
or U13154 (N_13154,N_6745,N_5830);
xor U13155 (N_13155,N_6896,N_9375);
nor U13156 (N_13156,N_8401,N_5483);
or U13157 (N_13157,N_9204,N_7213);
and U13158 (N_13158,N_7850,N_9267);
xor U13159 (N_13159,N_7911,N_8091);
nand U13160 (N_13160,N_7288,N_9895);
xor U13161 (N_13161,N_7718,N_9210);
and U13162 (N_13162,N_7978,N_9120);
and U13163 (N_13163,N_6359,N_7560);
nand U13164 (N_13164,N_5123,N_9449);
and U13165 (N_13165,N_6530,N_9035);
or U13166 (N_13166,N_8262,N_7482);
and U13167 (N_13167,N_9016,N_8426);
and U13168 (N_13168,N_9613,N_9633);
nor U13169 (N_13169,N_7204,N_8375);
nor U13170 (N_13170,N_9981,N_8480);
or U13171 (N_13171,N_5814,N_6523);
or U13172 (N_13172,N_6493,N_7151);
and U13173 (N_13173,N_7980,N_5410);
and U13174 (N_13174,N_9614,N_6056);
and U13175 (N_13175,N_7382,N_5557);
or U13176 (N_13176,N_5397,N_7759);
or U13177 (N_13177,N_7188,N_5371);
nor U13178 (N_13178,N_5490,N_6711);
nand U13179 (N_13179,N_7263,N_8187);
nor U13180 (N_13180,N_6980,N_7127);
or U13181 (N_13181,N_6541,N_9663);
nand U13182 (N_13182,N_8403,N_6417);
nor U13183 (N_13183,N_5485,N_6272);
and U13184 (N_13184,N_7309,N_8107);
and U13185 (N_13185,N_7481,N_7233);
or U13186 (N_13186,N_8548,N_8463);
nand U13187 (N_13187,N_7615,N_9573);
or U13188 (N_13188,N_7247,N_9776);
nor U13189 (N_13189,N_9703,N_5908);
and U13190 (N_13190,N_9176,N_8116);
nand U13191 (N_13191,N_9141,N_9042);
nand U13192 (N_13192,N_8010,N_8137);
nor U13193 (N_13193,N_9790,N_9895);
or U13194 (N_13194,N_6897,N_7263);
nand U13195 (N_13195,N_5757,N_6393);
nor U13196 (N_13196,N_8990,N_5720);
nand U13197 (N_13197,N_9827,N_6476);
and U13198 (N_13198,N_5337,N_9284);
nand U13199 (N_13199,N_5151,N_6424);
nand U13200 (N_13200,N_8827,N_7855);
nand U13201 (N_13201,N_7594,N_7616);
and U13202 (N_13202,N_8320,N_8540);
or U13203 (N_13203,N_5859,N_6529);
and U13204 (N_13204,N_7786,N_9855);
or U13205 (N_13205,N_8434,N_5323);
xor U13206 (N_13206,N_9319,N_5762);
nand U13207 (N_13207,N_9138,N_7123);
nor U13208 (N_13208,N_9781,N_7135);
nand U13209 (N_13209,N_8127,N_5085);
nand U13210 (N_13210,N_6776,N_5123);
xor U13211 (N_13211,N_5794,N_7320);
nor U13212 (N_13212,N_9778,N_5939);
or U13213 (N_13213,N_8144,N_5027);
and U13214 (N_13214,N_6723,N_9248);
nand U13215 (N_13215,N_8035,N_9167);
or U13216 (N_13216,N_9624,N_9918);
nand U13217 (N_13217,N_8371,N_7261);
and U13218 (N_13218,N_7053,N_6138);
and U13219 (N_13219,N_7652,N_6756);
nor U13220 (N_13220,N_6091,N_6081);
nor U13221 (N_13221,N_6790,N_5951);
nand U13222 (N_13222,N_5140,N_7667);
nor U13223 (N_13223,N_8437,N_5813);
nor U13224 (N_13224,N_8899,N_8303);
and U13225 (N_13225,N_6287,N_5108);
or U13226 (N_13226,N_9249,N_9598);
nor U13227 (N_13227,N_8931,N_9952);
or U13228 (N_13228,N_7146,N_7744);
nand U13229 (N_13229,N_7578,N_8560);
and U13230 (N_13230,N_6397,N_6615);
xor U13231 (N_13231,N_6530,N_8529);
and U13232 (N_13232,N_8261,N_7214);
nand U13233 (N_13233,N_6834,N_8772);
or U13234 (N_13234,N_5805,N_8258);
xnor U13235 (N_13235,N_7349,N_5671);
nand U13236 (N_13236,N_9820,N_5333);
and U13237 (N_13237,N_5125,N_7267);
nand U13238 (N_13238,N_5604,N_7596);
or U13239 (N_13239,N_9516,N_8644);
or U13240 (N_13240,N_8685,N_8167);
and U13241 (N_13241,N_6150,N_7170);
nand U13242 (N_13242,N_5846,N_7719);
or U13243 (N_13243,N_9735,N_7701);
nor U13244 (N_13244,N_7413,N_5790);
and U13245 (N_13245,N_9204,N_8938);
nor U13246 (N_13246,N_9460,N_6875);
nor U13247 (N_13247,N_6245,N_8261);
nand U13248 (N_13248,N_8815,N_8406);
and U13249 (N_13249,N_9810,N_5115);
or U13250 (N_13250,N_9717,N_7287);
and U13251 (N_13251,N_7117,N_7493);
xnor U13252 (N_13252,N_8824,N_8375);
nor U13253 (N_13253,N_5461,N_9823);
nor U13254 (N_13254,N_6221,N_9307);
or U13255 (N_13255,N_8080,N_6023);
nand U13256 (N_13256,N_6468,N_7431);
and U13257 (N_13257,N_6873,N_5921);
xnor U13258 (N_13258,N_5114,N_8764);
nand U13259 (N_13259,N_7144,N_8284);
nand U13260 (N_13260,N_7382,N_8744);
nand U13261 (N_13261,N_5215,N_8572);
and U13262 (N_13262,N_6865,N_6715);
nor U13263 (N_13263,N_8078,N_5301);
nor U13264 (N_13264,N_6215,N_6698);
xor U13265 (N_13265,N_9649,N_6804);
nor U13266 (N_13266,N_6393,N_6525);
and U13267 (N_13267,N_9791,N_5783);
or U13268 (N_13268,N_9422,N_6468);
and U13269 (N_13269,N_7039,N_6077);
or U13270 (N_13270,N_8851,N_5653);
nor U13271 (N_13271,N_5476,N_7772);
nand U13272 (N_13272,N_6396,N_6268);
or U13273 (N_13273,N_8586,N_7251);
nor U13274 (N_13274,N_5448,N_9835);
xnor U13275 (N_13275,N_5706,N_7166);
and U13276 (N_13276,N_9042,N_5393);
and U13277 (N_13277,N_5731,N_8425);
or U13278 (N_13278,N_8304,N_5683);
nor U13279 (N_13279,N_8483,N_6993);
or U13280 (N_13280,N_9726,N_7946);
nand U13281 (N_13281,N_5743,N_7814);
xnor U13282 (N_13282,N_7134,N_8445);
or U13283 (N_13283,N_5966,N_8502);
or U13284 (N_13284,N_7974,N_8933);
nand U13285 (N_13285,N_9092,N_5540);
and U13286 (N_13286,N_5909,N_6807);
nand U13287 (N_13287,N_6799,N_6286);
nand U13288 (N_13288,N_7043,N_8953);
and U13289 (N_13289,N_5343,N_9563);
and U13290 (N_13290,N_7266,N_8942);
and U13291 (N_13291,N_8243,N_9174);
xnor U13292 (N_13292,N_5168,N_7001);
nor U13293 (N_13293,N_5948,N_8340);
nand U13294 (N_13294,N_5708,N_9731);
or U13295 (N_13295,N_5127,N_9111);
nand U13296 (N_13296,N_8456,N_5732);
nor U13297 (N_13297,N_6858,N_8302);
nor U13298 (N_13298,N_8338,N_6781);
and U13299 (N_13299,N_9528,N_5771);
nor U13300 (N_13300,N_5287,N_5586);
nor U13301 (N_13301,N_8577,N_5412);
nor U13302 (N_13302,N_9825,N_9586);
or U13303 (N_13303,N_5529,N_9228);
nand U13304 (N_13304,N_6103,N_5882);
nand U13305 (N_13305,N_9521,N_8135);
and U13306 (N_13306,N_5354,N_7442);
and U13307 (N_13307,N_8147,N_8813);
and U13308 (N_13308,N_7987,N_6782);
or U13309 (N_13309,N_6860,N_5271);
and U13310 (N_13310,N_9585,N_6999);
and U13311 (N_13311,N_5048,N_6294);
or U13312 (N_13312,N_6615,N_9175);
nand U13313 (N_13313,N_6510,N_5504);
nand U13314 (N_13314,N_8286,N_5685);
nand U13315 (N_13315,N_6220,N_9026);
and U13316 (N_13316,N_9216,N_7563);
xor U13317 (N_13317,N_8998,N_8624);
nor U13318 (N_13318,N_7384,N_6067);
nand U13319 (N_13319,N_8075,N_6478);
xnor U13320 (N_13320,N_8354,N_5926);
and U13321 (N_13321,N_6078,N_7929);
xor U13322 (N_13322,N_5189,N_8971);
or U13323 (N_13323,N_9455,N_6200);
and U13324 (N_13324,N_7437,N_8339);
or U13325 (N_13325,N_7018,N_5373);
nor U13326 (N_13326,N_7589,N_7644);
and U13327 (N_13327,N_6498,N_5860);
nor U13328 (N_13328,N_8061,N_8492);
or U13329 (N_13329,N_9313,N_9871);
nor U13330 (N_13330,N_6857,N_8674);
or U13331 (N_13331,N_8890,N_5040);
and U13332 (N_13332,N_6168,N_6042);
and U13333 (N_13333,N_7545,N_8633);
xnor U13334 (N_13334,N_8415,N_6594);
xnor U13335 (N_13335,N_5566,N_6184);
or U13336 (N_13336,N_7499,N_6832);
xnor U13337 (N_13337,N_6637,N_9792);
nor U13338 (N_13338,N_6106,N_6162);
nand U13339 (N_13339,N_7666,N_5100);
nand U13340 (N_13340,N_7052,N_7226);
xor U13341 (N_13341,N_6537,N_7896);
nand U13342 (N_13342,N_8151,N_7843);
nand U13343 (N_13343,N_5398,N_7697);
xnor U13344 (N_13344,N_7305,N_8603);
or U13345 (N_13345,N_7658,N_6568);
xnor U13346 (N_13346,N_8066,N_6082);
nand U13347 (N_13347,N_8023,N_5919);
and U13348 (N_13348,N_8692,N_6905);
nor U13349 (N_13349,N_9496,N_5664);
or U13350 (N_13350,N_8021,N_8529);
and U13351 (N_13351,N_8482,N_5257);
or U13352 (N_13352,N_7367,N_6373);
or U13353 (N_13353,N_9229,N_8216);
nor U13354 (N_13354,N_6974,N_5574);
nand U13355 (N_13355,N_5386,N_6511);
nor U13356 (N_13356,N_5965,N_9526);
nor U13357 (N_13357,N_5475,N_9594);
and U13358 (N_13358,N_8787,N_6949);
and U13359 (N_13359,N_8549,N_8299);
or U13360 (N_13360,N_9830,N_8627);
nand U13361 (N_13361,N_7432,N_9894);
nor U13362 (N_13362,N_9500,N_5505);
xnor U13363 (N_13363,N_8831,N_8270);
nor U13364 (N_13364,N_7168,N_5880);
nor U13365 (N_13365,N_5125,N_7976);
or U13366 (N_13366,N_9635,N_6719);
nand U13367 (N_13367,N_5317,N_5044);
nor U13368 (N_13368,N_9526,N_5589);
nand U13369 (N_13369,N_6086,N_8894);
nand U13370 (N_13370,N_8081,N_7424);
or U13371 (N_13371,N_8195,N_6071);
and U13372 (N_13372,N_7251,N_7230);
or U13373 (N_13373,N_6752,N_5767);
nor U13374 (N_13374,N_9484,N_9903);
nor U13375 (N_13375,N_7860,N_6847);
and U13376 (N_13376,N_7978,N_8796);
and U13377 (N_13377,N_5841,N_8749);
or U13378 (N_13378,N_8891,N_6280);
and U13379 (N_13379,N_7798,N_9069);
nor U13380 (N_13380,N_5921,N_8393);
xor U13381 (N_13381,N_8468,N_6763);
nor U13382 (N_13382,N_5859,N_9766);
nand U13383 (N_13383,N_7347,N_6240);
xnor U13384 (N_13384,N_6225,N_6231);
xnor U13385 (N_13385,N_9458,N_8890);
nor U13386 (N_13386,N_8771,N_8853);
or U13387 (N_13387,N_8963,N_6589);
nand U13388 (N_13388,N_8167,N_6545);
or U13389 (N_13389,N_6902,N_8234);
nor U13390 (N_13390,N_8370,N_7357);
nor U13391 (N_13391,N_9248,N_6793);
nand U13392 (N_13392,N_9535,N_8417);
and U13393 (N_13393,N_5754,N_9224);
nor U13394 (N_13394,N_7252,N_7914);
nor U13395 (N_13395,N_6647,N_8073);
or U13396 (N_13396,N_5761,N_6860);
nor U13397 (N_13397,N_5898,N_8554);
xnor U13398 (N_13398,N_9094,N_9498);
xnor U13399 (N_13399,N_8243,N_8241);
or U13400 (N_13400,N_5263,N_8286);
and U13401 (N_13401,N_7848,N_7421);
nor U13402 (N_13402,N_7059,N_5512);
nand U13403 (N_13403,N_7827,N_8869);
nor U13404 (N_13404,N_8250,N_5037);
or U13405 (N_13405,N_6048,N_5607);
nand U13406 (N_13406,N_9874,N_9532);
xnor U13407 (N_13407,N_5700,N_6536);
and U13408 (N_13408,N_5547,N_9591);
and U13409 (N_13409,N_9142,N_9190);
nand U13410 (N_13410,N_6498,N_8787);
nand U13411 (N_13411,N_7370,N_5711);
nand U13412 (N_13412,N_9971,N_5845);
nand U13413 (N_13413,N_8535,N_6942);
nor U13414 (N_13414,N_8745,N_8650);
and U13415 (N_13415,N_9087,N_9283);
nand U13416 (N_13416,N_5354,N_9268);
and U13417 (N_13417,N_5170,N_7065);
and U13418 (N_13418,N_8859,N_7658);
xnor U13419 (N_13419,N_8610,N_9531);
and U13420 (N_13420,N_5839,N_6844);
and U13421 (N_13421,N_9396,N_6376);
xor U13422 (N_13422,N_8425,N_8349);
nand U13423 (N_13423,N_9847,N_8150);
and U13424 (N_13424,N_9636,N_8343);
nand U13425 (N_13425,N_7258,N_8644);
or U13426 (N_13426,N_5961,N_6555);
and U13427 (N_13427,N_7838,N_5973);
nor U13428 (N_13428,N_8115,N_5414);
and U13429 (N_13429,N_9712,N_6233);
nand U13430 (N_13430,N_6298,N_5261);
and U13431 (N_13431,N_9256,N_8087);
xor U13432 (N_13432,N_5489,N_5472);
and U13433 (N_13433,N_9076,N_8023);
nor U13434 (N_13434,N_7849,N_9475);
nor U13435 (N_13435,N_7463,N_9339);
nand U13436 (N_13436,N_7659,N_6689);
and U13437 (N_13437,N_6710,N_6507);
and U13438 (N_13438,N_8504,N_9091);
nand U13439 (N_13439,N_5558,N_7633);
or U13440 (N_13440,N_5410,N_5973);
and U13441 (N_13441,N_7731,N_6897);
nor U13442 (N_13442,N_9708,N_9520);
nand U13443 (N_13443,N_7537,N_6023);
or U13444 (N_13444,N_6859,N_6022);
and U13445 (N_13445,N_5932,N_9116);
xor U13446 (N_13446,N_8325,N_5470);
nand U13447 (N_13447,N_7731,N_6652);
nor U13448 (N_13448,N_7565,N_6360);
nor U13449 (N_13449,N_6852,N_8163);
and U13450 (N_13450,N_8734,N_7465);
and U13451 (N_13451,N_7026,N_5882);
or U13452 (N_13452,N_7511,N_9236);
or U13453 (N_13453,N_6866,N_9739);
or U13454 (N_13454,N_8260,N_9329);
nor U13455 (N_13455,N_6710,N_5270);
nand U13456 (N_13456,N_5770,N_7572);
or U13457 (N_13457,N_5100,N_5393);
or U13458 (N_13458,N_6078,N_9194);
or U13459 (N_13459,N_8487,N_6333);
nor U13460 (N_13460,N_5804,N_5728);
and U13461 (N_13461,N_8589,N_7891);
nand U13462 (N_13462,N_9584,N_5743);
nor U13463 (N_13463,N_8568,N_9544);
xnor U13464 (N_13464,N_5993,N_7516);
nor U13465 (N_13465,N_8402,N_6614);
and U13466 (N_13466,N_5943,N_9448);
nand U13467 (N_13467,N_6476,N_7677);
and U13468 (N_13468,N_9145,N_6294);
and U13469 (N_13469,N_5431,N_7364);
nand U13470 (N_13470,N_6044,N_7537);
or U13471 (N_13471,N_9902,N_6436);
nand U13472 (N_13472,N_6131,N_8708);
nor U13473 (N_13473,N_7839,N_8721);
and U13474 (N_13474,N_6510,N_7353);
and U13475 (N_13475,N_9853,N_8248);
nor U13476 (N_13476,N_5981,N_7089);
nor U13477 (N_13477,N_7340,N_6124);
or U13478 (N_13478,N_7192,N_9813);
and U13479 (N_13479,N_9770,N_7523);
or U13480 (N_13480,N_9166,N_5566);
nor U13481 (N_13481,N_8505,N_9738);
or U13482 (N_13482,N_9725,N_6229);
nor U13483 (N_13483,N_6028,N_6068);
and U13484 (N_13484,N_7024,N_6762);
or U13485 (N_13485,N_8214,N_5057);
nand U13486 (N_13486,N_8743,N_6676);
nor U13487 (N_13487,N_7254,N_8123);
nor U13488 (N_13488,N_9776,N_6984);
and U13489 (N_13489,N_6808,N_5530);
and U13490 (N_13490,N_9025,N_6841);
or U13491 (N_13491,N_5549,N_9034);
or U13492 (N_13492,N_5254,N_7526);
nand U13493 (N_13493,N_6097,N_6139);
xor U13494 (N_13494,N_5250,N_9988);
nand U13495 (N_13495,N_8123,N_9579);
and U13496 (N_13496,N_5847,N_8344);
and U13497 (N_13497,N_9668,N_7097);
xor U13498 (N_13498,N_8253,N_9025);
nand U13499 (N_13499,N_5772,N_8675);
nand U13500 (N_13500,N_9183,N_7528);
nor U13501 (N_13501,N_8150,N_6117);
nor U13502 (N_13502,N_7677,N_8099);
xnor U13503 (N_13503,N_7252,N_5115);
nand U13504 (N_13504,N_7703,N_8750);
nand U13505 (N_13505,N_8571,N_9716);
or U13506 (N_13506,N_5638,N_5183);
or U13507 (N_13507,N_9700,N_9806);
nor U13508 (N_13508,N_8293,N_7710);
or U13509 (N_13509,N_7915,N_7114);
and U13510 (N_13510,N_7750,N_7934);
xor U13511 (N_13511,N_9806,N_9155);
xnor U13512 (N_13512,N_6664,N_8825);
and U13513 (N_13513,N_7282,N_7074);
nand U13514 (N_13514,N_5997,N_6552);
nand U13515 (N_13515,N_6478,N_7773);
and U13516 (N_13516,N_8163,N_9353);
xor U13517 (N_13517,N_9385,N_9012);
nand U13518 (N_13518,N_9081,N_7085);
and U13519 (N_13519,N_6235,N_6797);
and U13520 (N_13520,N_5569,N_6355);
and U13521 (N_13521,N_8074,N_5252);
or U13522 (N_13522,N_6572,N_7409);
nor U13523 (N_13523,N_9666,N_5660);
and U13524 (N_13524,N_5859,N_6933);
or U13525 (N_13525,N_9507,N_7193);
nand U13526 (N_13526,N_5949,N_7145);
and U13527 (N_13527,N_8123,N_8127);
nor U13528 (N_13528,N_5952,N_6600);
xor U13529 (N_13529,N_6957,N_8260);
nor U13530 (N_13530,N_7547,N_6953);
and U13531 (N_13531,N_5310,N_9936);
nand U13532 (N_13532,N_6287,N_8434);
and U13533 (N_13533,N_5750,N_7035);
nor U13534 (N_13534,N_6814,N_7505);
nor U13535 (N_13535,N_8792,N_7530);
nand U13536 (N_13536,N_5409,N_5538);
nand U13537 (N_13537,N_8147,N_9693);
nor U13538 (N_13538,N_6491,N_6810);
or U13539 (N_13539,N_9048,N_5900);
xor U13540 (N_13540,N_5833,N_5460);
or U13541 (N_13541,N_9279,N_6987);
nand U13542 (N_13542,N_9701,N_5312);
nand U13543 (N_13543,N_8526,N_5133);
or U13544 (N_13544,N_5305,N_6918);
nor U13545 (N_13545,N_6810,N_6742);
xnor U13546 (N_13546,N_8372,N_6895);
nand U13547 (N_13547,N_7062,N_5936);
and U13548 (N_13548,N_7297,N_8893);
or U13549 (N_13549,N_5233,N_8876);
nor U13550 (N_13550,N_5037,N_6712);
xor U13551 (N_13551,N_9669,N_9426);
and U13552 (N_13552,N_5260,N_6385);
nor U13553 (N_13553,N_8980,N_6401);
nor U13554 (N_13554,N_7673,N_9035);
or U13555 (N_13555,N_8528,N_8987);
xor U13556 (N_13556,N_8567,N_9721);
or U13557 (N_13557,N_6451,N_5431);
nand U13558 (N_13558,N_5459,N_9107);
and U13559 (N_13559,N_5622,N_9896);
and U13560 (N_13560,N_8897,N_6662);
or U13561 (N_13561,N_9947,N_8663);
and U13562 (N_13562,N_9576,N_5877);
nor U13563 (N_13563,N_5196,N_7612);
or U13564 (N_13564,N_5638,N_8255);
or U13565 (N_13565,N_5031,N_8233);
nor U13566 (N_13566,N_8636,N_5405);
or U13567 (N_13567,N_7771,N_7597);
nand U13568 (N_13568,N_5134,N_6770);
xor U13569 (N_13569,N_8875,N_7948);
nor U13570 (N_13570,N_9462,N_6961);
nand U13571 (N_13571,N_6706,N_7978);
and U13572 (N_13572,N_6455,N_9236);
nand U13573 (N_13573,N_7056,N_7723);
and U13574 (N_13574,N_7094,N_9153);
nor U13575 (N_13575,N_9954,N_6401);
and U13576 (N_13576,N_8332,N_6207);
nand U13577 (N_13577,N_7432,N_7988);
or U13578 (N_13578,N_8825,N_9208);
or U13579 (N_13579,N_5891,N_5324);
and U13580 (N_13580,N_7801,N_7814);
and U13581 (N_13581,N_9381,N_6119);
xor U13582 (N_13582,N_7581,N_5225);
and U13583 (N_13583,N_8225,N_8091);
and U13584 (N_13584,N_7479,N_9260);
nand U13585 (N_13585,N_5246,N_9159);
or U13586 (N_13586,N_5133,N_6470);
nor U13587 (N_13587,N_5051,N_8404);
and U13588 (N_13588,N_7620,N_8900);
xor U13589 (N_13589,N_8988,N_9551);
nor U13590 (N_13590,N_6443,N_8164);
or U13591 (N_13591,N_6066,N_7202);
nor U13592 (N_13592,N_6166,N_6349);
nand U13593 (N_13593,N_8370,N_6448);
and U13594 (N_13594,N_9977,N_9204);
nor U13595 (N_13595,N_6591,N_8673);
nor U13596 (N_13596,N_6258,N_7581);
and U13597 (N_13597,N_7577,N_7795);
nand U13598 (N_13598,N_7906,N_5646);
or U13599 (N_13599,N_9317,N_9405);
nor U13600 (N_13600,N_6002,N_8282);
or U13601 (N_13601,N_8140,N_5097);
nand U13602 (N_13602,N_6464,N_9893);
and U13603 (N_13603,N_8508,N_8087);
nand U13604 (N_13604,N_9313,N_9502);
or U13605 (N_13605,N_9743,N_9697);
and U13606 (N_13606,N_5745,N_5735);
and U13607 (N_13607,N_8317,N_8650);
nand U13608 (N_13608,N_6355,N_5111);
nor U13609 (N_13609,N_8027,N_9812);
xor U13610 (N_13610,N_9635,N_6643);
nand U13611 (N_13611,N_8251,N_8383);
nor U13612 (N_13612,N_6001,N_5680);
nand U13613 (N_13613,N_8334,N_9308);
nand U13614 (N_13614,N_9697,N_9216);
or U13615 (N_13615,N_6602,N_5314);
nor U13616 (N_13616,N_7801,N_9660);
xor U13617 (N_13617,N_9565,N_6428);
nand U13618 (N_13618,N_5140,N_8705);
xnor U13619 (N_13619,N_7463,N_8183);
and U13620 (N_13620,N_6986,N_7462);
nand U13621 (N_13621,N_8160,N_9582);
and U13622 (N_13622,N_8130,N_8924);
or U13623 (N_13623,N_6012,N_7426);
or U13624 (N_13624,N_5159,N_8145);
nor U13625 (N_13625,N_6109,N_9052);
xnor U13626 (N_13626,N_8255,N_5052);
nor U13627 (N_13627,N_5521,N_8787);
nand U13628 (N_13628,N_9039,N_6924);
and U13629 (N_13629,N_5765,N_9869);
nor U13630 (N_13630,N_6680,N_8114);
or U13631 (N_13631,N_7462,N_6636);
nand U13632 (N_13632,N_7045,N_9812);
and U13633 (N_13633,N_8812,N_5894);
nand U13634 (N_13634,N_5717,N_7229);
nand U13635 (N_13635,N_7144,N_6967);
or U13636 (N_13636,N_6571,N_7181);
nand U13637 (N_13637,N_7188,N_6502);
nand U13638 (N_13638,N_5508,N_6786);
nand U13639 (N_13639,N_7269,N_5401);
and U13640 (N_13640,N_7121,N_7521);
xor U13641 (N_13641,N_7529,N_5824);
and U13642 (N_13642,N_8597,N_5486);
nor U13643 (N_13643,N_9750,N_6199);
or U13644 (N_13644,N_6216,N_9992);
xor U13645 (N_13645,N_7628,N_7209);
and U13646 (N_13646,N_6336,N_8363);
nand U13647 (N_13647,N_7058,N_8673);
nor U13648 (N_13648,N_8841,N_8715);
or U13649 (N_13649,N_5846,N_7815);
and U13650 (N_13650,N_5442,N_8753);
and U13651 (N_13651,N_5821,N_5419);
nand U13652 (N_13652,N_8975,N_6557);
nor U13653 (N_13653,N_8836,N_7573);
nand U13654 (N_13654,N_8926,N_5124);
nand U13655 (N_13655,N_8423,N_7300);
nor U13656 (N_13656,N_9157,N_5184);
nand U13657 (N_13657,N_5030,N_9575);
or U13658 (N_13658,N_7754,N_8077);
or U13659 (N_13659,N_9033,N_5085);
nand U13660 (N_13660,N_5731,N_7921);
nor U13661 (N_13661,N_9891,N_8949);
or U13662 (N_13662,N_9235,N_6826);
nand U13663 (N_13663,N_5654,N_9929);
nor U13664 (N_13664,N_9690,N_5054);
and U13665 (N_13665,N_7750,N_5840);
nand U13666 (N_13666,N_5503,N_9225);
nor U13667 (N_13667,N_9018,N_9105);
nor U13668 (N_13668,N_6845,N_9880);
or U13669 (N_13669,N_9709,N_8363);
nor U13670 (N_13670,N_9262,N_5234);
or U13671 (N_13671,N_6397,N_5230);
and U13672 (N_13672,N_9474,N_8266);
nand U13673 (N_13673,N_6375,N_7978);
and U13674 (N_13674,N_5719,N_7814);
or U13675 (N_13675,N_6567,N_7736);
xor U13676 (N_13676,N_7464,N_9884);
xor U13677 (N_13677,N_7168,N_8109);
nand U13678 (N_13678,N_5135,N_8514);
nor U13679 (N_13679,N_6074,N_9575);
nor U13680 (N_13680,N_6437,N_9564);
nand U13681 (N_13681,N_5542,N_8329);
nand U13682 (N_13682,N_8622,N_8026);
nor U13683 (N_13683,N_9168,N_8390);
nor U13684 (N_13684,N_9904,N_5244);
nor U13685 (N_13685,N_9445,N_9476);
nor U13686 (N_13686,N_5809,N_6426);
nand U13687 (N_13687,N_9070,N_9901);
and U13688 (N_13688,N_9790,N_6712);
and U13689 (N_13689,N_9228,N_9251);
and U13690 (N_13690,N_5243,N_6814);
or U13691 (N_13691,N_8377,N_5204);
nand U13692 (N_13692,N_8051,N_9943);
and U13693 (N_13693,N_8580,N_7521);
nor U13694 (N_13694,N_7817,N_9067);
or U13695 (N_13695,N_6088,N_9281);
nor U13696 (N_13696,N_5571,N_8243);
and U13697 (N_13697,N_9642,N_7598);
nand U13698 (N_13698,N_5731,N_9214);
nand U13699 (N_13699,N_8881,N_5369);
and U13700 (N_13700,N_7111,N_8140);
and U13701 (N_13701,N_7201,N_8256);
xnor U13702 (N_13702,N_9468,N_6773);
or U13703 (N_13703,N_9362,N_6916);
nand U13704 (N_13704,N_7635,N_6754);
xor U13705 (N_13705,N_7750,N_9728);
or U13706 (N_13706,N_9011,N_5446);
and U13707 (N_13707,N_7496,N_5660);
and U13708 (N_13708,N_9640,N_7639);
or U13709 (N_13709,N_9732,N_9916);
nand U13710 (N_13710,N_7110,N_6950);
nor U13711 (N_13711,N_7069,N_8169);
or U13712 (N_13712,N_8230,N_7756);
or U13713 (N_13713,N_5827,N_6444);
nand U13714 (N_13714,N_8973,N_8607);
and U13715 (N_13715,N_9505,N_8662);
and U13716 (N_13716,N_9582,N_6136);
or U13717 (N_13717,N_6468,N_8161);
nand U13718 (N_13718,N_8495,N_8754);
nand U13719 (N_13719,N_9005,N_9490);
nor U13720 (N_13720,N_8131,N_5592);
nand U13721 (N_13721,N_5473,N_7828);
xnor U13722 (N_13722,N_7867,N_6183);
and U13723 (N_13723,N_8888,N_8360);
nor U13724 (N_13724,N_8006,N_6907);
nor U13725 (N_13725,N_7708,N_5505);
or U13726 (N_13726,N_8801,N_7404);
or U13727 (N_13727,N_9209,N_7362);
and U13728 (N_13728,N_8162,N_6707);
nor U13729 (N_13729,N_5211,N_7030);
xnor U13730 (N_13730,N_5273,N_8276);
and U13731 (N_13731,N_5713,N_7479);
and U13732 (N_13732,N_6001,N_9094);
or U13733 (N_13733,N_5008,N_9449);
nor U13734 (N_13734,N_7974,N_5123);
nor U13735 (N_13735,N_9872,N_6038);
xnor U13736 (N_13736,N_8203,N_8896);
nand U13737 (N_13737,N_7580,N_5687);
or U13738 (N_13738,N_9728,N_6435);
nor U13739 (N_13739,N_9513,N_8864);
nand U13740 (N_13740,N_7731,N_8766);
or U13741 (N_13741,N_5671,N_8666);
nand U13742 (N_13742,N_5553,N_5384);
or U13743 (N_13743,N_8130,N_8942);
or U13744 (N_13744,N_7007,N_8828);
nor U13745 (N_13745,N_8746,N_6471);
nand U13746 (N_13746,N_8217,N_5563);
nand U13747 (N_13747,N_7151,N_9645);
or U13748 (N_13748,N_9196,N_8314);
nand U13749 (N_13749,N_9144,N_7889);
nand U13750 (N_13750,N_5132,N_9069);
or U13751 (N_13751,N_6910,N_6283);
or U13752 (N_13752,N_6271,N_7503);
and U13753 (N_13753,N_9820,N_6304);
nand U13754 (N_13754,N_6508,N_9765);
xor U13755 (N_13755,N_6974,N_8615);
nand U13756 (N_13756,N_6324,N_9986);
nor U13757 (N_13757,N_8089,N_6682);
nor U13758 (N_13758,N_6536,N_9954);
nor U13759 (N_13759,N_5579,N_7691);
and U13760 (N_13760,N_6572,N_8505);
nor U13761 (N_13761,N_6258,N_9671);
nand U13762 (N_13762,N_6767,N_6853);
and U13763 (N_13763,N_7698,N_8041);
nand U13764 (N_13764,N_7852,N_8866);
nor U13765 (N_13765,N_5931,N_9613);
nor U13766 (N_13766,N_5985,N_6650);
xnor U13767 (N_13767,N_8634,N_9271);
nand U13768 (N_13768,N_8407,N_5854);
nor U13769 (N_13769,N_9487,N_7261);
or U13770 (N_13770,N_6057,N_6817);
or U13771 (N_13771,N_5671,N_7465);
or U13772 (N_13772,N_7287,N_8831);
and U13773 (N_13773,N_7355,N_9761);
nand U13774 (N_13774,N_8029,N_9287);
and U13775 (N_13775,N_8188,N_9880);
and U13776 (N_13776,N_9732,N_6594);
xor U13777 (N_13777,N_5028,N_8267);
nor U13778 (N_13778,N_9641,N_7634);
nand U13779 (N_13779,N_6128,N_9835);
nand U13780 (N_13780,N_8467,N_7953);
nand U13781 (N_13781,N_5596,N_8579);
nor U13782 (N_13782,N_7910,N_9929);
xnor U13783 (N_13783,N_9478,N_9974);
and U13784 (N_13784,N_7190,N_6997);
or U13785 (N_13785,N_6136,N_5084);
and U13786 (N_13786,N_9885,N_7206);
and U13787 (N_13787,N_6220,N_7997);
nand U13788 (N_13788,N_5770,N_8595);
xor U13789 (N_13789,N_9634,N_6826);
and U13790 (N_13790,N_8800,N_9860);
xnor U13791 (N_13791,N_7470,N_7127);
nand U13792 (N_13792,N_9588,N_7516);
or U13793 (N_13793,N_9515,N_5099);
nor U13794 (N_13794,N_9260,N_9815);
and U13795 (N_13795,N_9004,N_5097);
nand U13796 (N_13796,N_5836,N_7639);
or U13797 (N_13797,N_8070,N_5766);
nor U13798 (N_13798,N_5225,N_5064);
nand U13799 (N_13799,N_8482,N_6467);
nand U13800 (N_13800,N_6314,N_8462);
or U13801 (N_13801,N_7636,N_7192);
nand U13802 (N_13802,N_8330,N_5417);
or U13803 (N_13803,N_9272,N_5019);
and U13804 (N_13804,N_8074,N_7014);
and U13805 (N_13805,N_8393,N_9891);
nand U13806 (N_13806,N_6920,N_5011);
or U13807 (N_13807,N_6970,N_6407);
and U13808 (N_13808,N_9743,N_9910);
nor U13809 (N_13809,N_8709,N_7094);
or U13810 (N_13810,N_9492,N_9313);
nand U13811 (N_13811,N_9888,N_5040);
or U13812 (N_13812,N_9955,N_6570);
or U13813 (N_13813,N_8275,N_7517);
nor U13814 (N_13814,N_7925,N_7409);
nand U13815 (N_13815,N_9501,N_5317);
or U13816 (N_13816,N_5054,N_6430);
or U13817 (N_13817,N_6721,N_8632);
nor U13818 (N_13818,N_8830,N_7116);
nand U13819 (N_13819,N_8390,N_5644);
and U13820 (N_13820,N_7447,N_7749);
or U13821 (N_13821,N_8174,N_6629);
or U13822 (N_13822,N_9132,N_8491);
or U13823 (N_13823,N_7187,N_9941);
or U13824 (N_13824,N_6231,N_6007);
nand U13825 (N_13825,N_7201,N_8721);
or U13826 (N_13826,N_7255,N_8629);
xor U13827 (N_13827,N_7785,N_5232);
nand U13828 (N_13828,N_8818,N_7737);
nand U13829 (N_13829,N_5213,N_7810);
nor U13830 (N_13830,N_6787,N_5673);
or U13831 (N_13831,N_6806,N_9689);
and U13832 (N_13832,N_9103,N_5932);
and U13833 (N_13833,N_9535,N_6204);
and U13834 (N_13834,N_5561,N_7792);
and U13835 (N_13835,N_9166,N_6063);
nor U13836 (N_13836,N_5126,N_5197);
or U13837 (N_13837,N_7152,N_8270);
nand U13838 (N_13838,N_8345,N_6189);
or U13839 (N_13839,N_7369,N_9753);
nand U13840 (N_13840,N_6862,N_5799);
and U13841 (N_13841,N_8775,N_8865);
nand U13842 (N_13842,N_6944,N_9266);
xor U13843 (N_13843,N_8264,N_5035);
nand U13844 (N_13844,N_9853,N_5409);
nor U13845 (N_13845,N_6007,N_9769);
or U13846 (N_13846,N_8676,N_7160);
nor U13847 (N_13847,N_9724,N_7080);
nand U13848 (N_13848,N_8806,N_6216);
nor U13849 (N_13849,N_8557,N_5418);
nor U13850 (N_13850,N_7974,N_6286);
nor U13851 (N_13851,N_6779,N_8014);
xor U13852 (N_13852,N_8838,N_5862);
nand U13853 (N_13853,N_9370,N_7751);
and U13854 (N_13854,N_5082,N_7231);
nor U13855 (N_13855,N_5512,N_7687);
nor U13856 (N_13856,N_6670,N_7448);
nand U13857 (N_13857,N_7614,N_6778);
nand U13858 (N_13858,N_6446,N_6468);
nor U13859 (N_13859,N_8604,N_8361);
nor U13860 (N_13860,N_6832,N_5330);
and U13861 (N_13861,N_9022,N_5878);
or U13862 (N_13862,N_8501,N_5979);
and U13863 (N_13863,N_5465,N_5932);
nor U13864 (N_13864,N_8207,N_6236);
nor U13865 (N_13865,N_6073,N_5840);
and U13866 (N_13866,N_7463,N_5857);
nand U13867 (N_13867,N_6822,N_6395);
or U13868 (N_13868,N_6680,N_9184);
nor U13869 (N_13869,N_8724,N_5036);
and U13870 (N_13870,N_6272,N_6408);
and U13871 (N_13871,N_9737,N_5760);
nor U13872 (N_13872,N_9912,N_7300);
and U13873 (N_13873,N_7819,N_5739);
nor U13874 (N_13874,N_8272,N_6887);
nor U13875 (N_13875,N_9023,N_6914);
and U13876 (N_13876,N_6098,N_9243);
or U13877 (N_13877,N_7674,N_6194);
nor U13878 (N_13878,N_8786,N_7600);
and U13879 (N_13879,N_5144,N_5193);
nor U13880 (N_13880,N_6725,N_5725);
or U13881 (N_13881,N_8447,N_5944);
nand U13882 (N_13882,N_8133,N_5924);
nor U13883 (N_13883,N_8595,N_7689);
nand U13884 (N_13884,N_9100,N_9802);
nor U13885 (N_13885,N_9916,N_7018);
xor U13886 (N_13886,N_8174,N_9395);
or U13887 (N_13887,N_9642,N_5542);
nor U13888 (N_13888,N_9416,N_8270);
and U13889 (N_13889,N_6403,N_8816);
and U13890 (N_13890,N_9379,N_8568);
nand U13891 (N_13891,N_7630,N_9365);
nor U13892 (N_13892,N_8787,N_7500);
and U13893 (N_13893,N_6643,N_8307);
nor U13894 (N_13894,N_9820,N_7703);
nor U13895 (N_13895,N_9502,N_9243);
nor U13896 (N_13896,N_9016,N_8712);
nand U13897 (N_13897,N_9254,N_8137);
and U13898 (N_13898,N_9244,N_8535);
or U13899 (N_13899,N_5017,N_6833);
or U13900 (N_13900,N_6091,N_7480);
nor U13901 (N_13901,N_7814,N_8212);
and U13902 (N_13902,N_9408,N_7832);
or U13903 (N_13903,N_5926,N_9204);
and U13904 (N_13904,N_5363,N_9962);
or U13905 (N_13905,N_6031,N_5855);
or U13906 (N_13906,N_9057,N_9924);
nand U13907 (N_13907,N_6862,N_5016);
nor U13908 (N_13908,N_5110,N_5862);
or U13909 (N_13909,N_7640,N_7512);
nor U13910 (N_13910,N_9839,N_7399);
or U13911 (N_13911,N_6536,N_9225);
nand U13912 (N_13912,N_7616,N_9720);
or U13913 (N_13913,N_6017,N_7556);
xor U13914 (N_13914,N_8676,N_5323);
or U13915 (N_13915,N_8843,N_8716);
and U13916 (N_13916,N_6891,N_8447);
and U13917 (N_13917,N_8655,N_7642);
xnor U13918 (N_13918,N_7504,N_5128);
and U13919 (N_13919,N_7330,N_7476);
and U13920 (N_13920,N_6334,N_6754);
and U13921 (N_13921,N_6323,N_6359);
and U13922 (N_13922,N_9675,N_6992);
or U13923 (N_13923,N_8598,N_9955);
xnor U13924 (N_13924,N_5830,N_6165);
xor U13925 (N_13925,N_5904,N_8851);
nand U13926 (N_13926,N_8346,N_9762);
nor U13927 (N_13927,N_7663,N_5804);
and U13928 (N_13928,N_8592,N_6549);
or U13929 (N_13929,N_6611,N_5003);
nor U13930 (N_13930,N_8613,N_6417);
nor U13931 (N_13931,N_7134,N_9922);
nand U13932 (N_13932,N_9858,N_5731);
and U13933 (N_13933,N_8718,N_8290);
and U13934 (N_13934,N_6004,N_5591);
nand U13935 (N_13935,N_7194,N_5276);
or U13936 (N_13936,N_9471,N_6564);
and U13937 (N_13937,N_5176,N_8716);
nand U13938 (N_13938,N_6517,N_8724);
and U13939 (N_13939,N_9612,N_9493);
nand U13940 (N_13940,N_9810,N_6071);
or U13941 (N_13941,N_7266,N_7610);
nor U13942 (N_13942,N_9755,N_8519);
and U13943 (N_13943,N_9491,N_7554);
nand U13944 (N_13944,N_9578,N_9883);
and U13945 (N_13945,N_5831,N_5095);
and U13946 (N_13946,N_5892,N_5109);
or U13947 (N_13947,N_6038,N_5763);
nor U13948 (N_13948,N_6713,N_7932);
nand U13949 (N_13949,N_5645,N_5613);
or U13950 (N_13950,N_7125,N_7916);
nand U13951 (N_13951,N_5563,N_6762);
and U13952 (N_13952,N_7531,N_8722);
nor U13953 (N_13953,N_9853,N_8986);
nor U13954 (N_13954,N_7092,N_8665);
or U13955 (N_13955,N_7349,N_6222);
xor U13956 (N_13956,N_9039,N_7825);
nor U13957 (N_13957,N_7557,N_8613);
and U13958 (N_13958,N_6007,N_8181);
nor U13959 (N_13959,N_6457,N_8612);
and U13960 (N_13960,N_5317,N_8442);
or U13961 (N_13961,N_8858,N_7847);
or U13962 (N_13962,N_9990,N_6443);
nand U13963 (N_13963,N_6118,N_6961);
and U13964 (N_13964,N_7181,N_6822);
and U13965 (N_13965,N_7561,N_5546);
or U13966 (N_13966,N_6010,N_9751);
or U13967 (N_13967,N_5482,N_6358);
and U13968 (N_13968,N_5595,N_7726);
nand U13969 (N_13969,N_6598,N_6070);
and U13970 (N_13970,N_9239,N_8739);
nor U13971 (N_13971,N_9014,N_7433);
nor U13972 (N_13972,N_7471,N_6682);
and U13973 (N_13973,N_8695,N_6355);
nand U13974 (N_13974,N_5778,N_6863);
nand U13975 (N_13975,N_5508,N_6734);
or U13976 (N_13976,N_7377,N_7158);
nand U13977 (N_13977,N_8886,N_6022);
nor U13978 (N_13978,N_6058,N_8716);
or U13979 (N_13979,N_6576,N_5752);
nand U13980 (N_13980,N_9129,N_8754);
or U13981 (N_13981,N_6308,N_8417);
or U13982 (N_13982,N_5060,N_6587);
nand U13983 (N_13983,N_7927,N_6843);
nand U13984 (N_13984,N_9357,N_7342);
xor U13985 (N_13985,N_5333,N_5737);
nand U13986 (N_13986,N_9077,N_7594);
xor U13987 (N_13987,N_5610,N_5584);
nor U13988 (N_13988,N_8976,N_7647);
or U13989 (N_13989,N_5277,N_9630);
or U13990 (N_13990,N_9272,N_9542);
and U13991 (N_13991,N_9995,N_7718);
or U13992 (N_13992,N_9447,N_6413);
xor U13993 (N_13993,N_6699,N_9270);
or U13994 (N_13994,N_9294,N_7169);
nand U13995 (N_13995,N_9385,N_5126);
or U13996 (N_13996,N_6454,N_9706);
nor U13997 (N_13997,N_6419,N_8459);
and U13998 (N_13998,N_9687,N_8203);
nor U13999 (N_13999,N_6609,N_6477);
or U14000 (N_14000,N_7335,N_8474);
nand U14001 (N_14001,N_9549,N_9020);
nand U14002 (N_14002,N_5352,N_5502);
nand U14003 (N_14003,N_9061,N_5803);
and U14004 (N_14004,N_8218,N_9499);
nor U14005 (N_14005,N_6224,N_9923);
nor U14006 (N_14006,N_9926,N_9456);
or U14007 (N_14007,N_6617,N_5700);
and U14008 (N_14008,N_9408,N_7158);
nand U14009 (N_14009,N_9002,N_5578);
and U14010 (N_14010,N_6554,N_9378);
nand U14011 (N_14011,N_5250,N_7573);
nand U14012 (N_14012,N_6327,N_6497);
nor U14013 (N_14013,N_8984,N_6312);
xnor U14014 (N_14014,N_8233,N_9556);
and U14015 (N_14015,N_6051,N_7146);
xnor U14016 (N_14016,N_5541,N_9520);
and U14017 (N_14017,N_7589,N_9290);
and U14018 (N_14018,N_6035,N_9118);
and U14019 (N_14019,N_8273,N_7927);
nand U14020 (N_14020,N_5375,N_7836);
and U14021 (N_14021,N_8427,N_9132);
or U14022 (N_14022,N_9080,N_9397);
or U14023 (N_14023,N_8850,N_9932);
nand U14024 (N_14024,N_9463,N_6167);
xor U14025 (N_14025,N_6852,N_6736);
nand U14026 (N_14026,N_5287,N_6774);
or U14027 (N_14027,N_8316,N_9809);
and U14028 (N_14028,N_6883,N_9802);
or U14029 (N_14029,N_9775,N_9383);
nand U14030 (N_14030,N_6607,N_7991);
xor U14031 (N_14031,N_5717,N_5175);
or U14032 (N_14032,N_7334,N_7124);
nor U14033 (N_14033,N_8098,N_7260);
or U14034 (N_14034,N_8933,N_5824);
xor U14035 (N_14035,N_6197,N_6501);
and U14036 (N_14036,N_8176,N_9013);
xnor U14037 (N_14037,N_6732,N_5857);
nand U14038 (N_14038,N_6194,N_6719);
nand U14039 (N_14039,N_9121,N_7171);
nand U14040 (N_14040,N_7279,N_6373);
nor U14041 (N_14041,N_5677,N_6044);
nor U14042 (N_14042,N_9516,N_6969);
nand U14043 (N_14043,N_7663,N_6537);
or U14044 (N_14044,N_7829,N_6659);
and U14045 (N_14045,N_7347,N_8784);
nor U14046 (N_14046,N_8049,N_5543);
nor U14047 (N_14047,N_5254,N_5282);
nand U14048 (N_14048,N_5530,N_5030);
or U14049 (N_14049,N_6257,N_7544);
or U14050 (N_14050,N_8207,N_9279);
nand U14051 (N_14051,N_9273,N_9501);
and U14052 (N_14052,N_6327,N_7796);
nand U14053 (N_14053,N_9936,N_7640);
or U14054 (N_14054,N_9467,N_6642);
nor U14055 (N_14055,N_5311,N_5543);
and U14056 (N_14056,N_6587,N_7767);
or U14057 (N_14057,N_5022,N_7495);
nand U14058 (N_14058,N_6000,N_7003);
xnor U14059 (N_14059,N_6373,N_9546);
and U14060 (N_14060,N_7029,N_8890);
nand U14061 (N_14061,N_6240,N_5441);
nor U14062 (N_14062,N_6923,N_8180);
nand U14063 (N_14063,N_5823,N_8272);
or U14064 (N_14064,N_6054,N_5960);
xor U14065 (N_14065,N_5710,N_8689);
xor U14066 (N_14066,N_7691,N_7584);
or U14067 (N_14067,N_9267,N_8149);
nor U14068 (N_14068,N_5427,N_5377);
or U14069 (N_14069,N_9945,N_9236);
or U14070 (N_14070,N_5816,N_7734);
and U14071 (N_14071,N_7279,N_5681);
xor U14072 (N_14072,N_7397,N_6121);
xnor U14073 (N_14073,N_8439,N_8150);
nor U14074 (N_14074,N_7618,N_5402);
or U14075 (N_14075,N_8708,N_8251);
nor U14076 (N_14076,N_5702,N_9989);
xor U14077 (N_14077,N_6694,N_6615);
xor U14078 (N_14078,N_7341,N_8300);
or U14079 (N_14079,N_5004,N_7575);
nor U14080 (N_14080,N_8434,N_6153);
and U14081 (N_14081,N_5470,N_5423);
xnor U14082 (N_14082,N_9747,N_8071);
or U14083 (N_14083,N_7731,N_5368);
or U14084 (N_14084,N_5949,N_9626);
xnor U14085 (N_14085,N_7280,N_8660);
nor U14086 (N_14086,N_7638,N_9065);
nor U14087 (N_14087,N_9183,N_8241);
or U14088 (N_14088,N_7790,N_6475);
nand U14089 (N_14089,N_8433,N_7677);
nor U14090 (N_14090,N_5822,N_8518);
or U14091 (N_14091,N_8129,N_7328);
or U14092 (N_14092,N_6613,N_9029);
nor U14093 (N_14093,N_5037,N_7103);
nand U14094 (N_14094,N_5235,N_8629);
xnor U14095 (N_14095,N_6325,N_9590);
or U14096 (N_14096,N_8960,N_9920);
or U14097 (N_14097,N_8644,N_5075);
nor U14098 (N_14098,N_6749,N_6261);
or U14099 (N_14099,N_8990,N_6534);
xor U14100 (N_14100,N_8215,N_8457);
nor U14101 (N_14101,N_7656,N_8721);
or U14102 (N_14102,N_6815,N_8370);
and U14103 (N_14103,N_6781,N_6189);
or U14104 (N_14104,N_5891,N_7008);
nand U14105 (N_14105,N_9752,N_8410);
nand U14106 (N_14106,N_5469,N_5339);
or U14107 (N_14107,N_7453,N_7071);
or U14108 (N_14108,N_8256,N_9140);
nand U14109 (N_14109,N_8391,N_5253);
nor U14110 (N_14110,N_7960,N_5489);
nor U14111 (N_14111,N_8180,N_8082);
nand U14112 (N_14112,N_7017,N_6902);
or U14113 (N_14113,N_9070,N_9755);
xor U14114 (N_14114,N_7446,N_8789);
nor U14115 (N_14115,N_5033,N_6300);
and U14116 (N_14116,N_9580,N_9102);
nand U14117 (N_14117,N_8533,N_8196);
nand U14118 (N_14118,N_8177,N_5161);
and U14119 (N_14119,N_6617,N_9442);
and U14120 (N_14120,N_9094,N_6527);
nand U14121 (N_14121,N_9147,N_9906);
xor U14122 (N_14122,N_9233,N_7817);
nand U14123 (N_14123,N_9054,N_9334);
xor U14124 (N_14124,N_6283,N_6098);
nor U14125 (N_14125,N_8097,N_5530);
nor U14126 (N_14126,N_9364,N_5546);
nand U14127 (N_14127,N_9870,N_7953);
nor U14128 (N_14128,N_5994,N_7079);
or U14129 (N_14129,N_9353,N_6328);
or U14130 (N_14130,N_8013,N_7158);
nor U14131 (N_14131,N_6737,N_5505);
xor U14132 (N_14132,N_5652,N_8275);
nand U14133 (N_14133,N_6209,N_6736);
xor U14134 (N_14134,N_5039,N_7015);
and U14135 (N_14135,N_6649,N_9726);
nor U14136 (N_14136,N_5982,N_9351);
or U14137 (N_14137,N_8624,N_5261);
or U14138 (N_14138,N_5409,N_6525);
and U14139 (N_14139,N_6534,N_7092);
nor U14140 (N_14140,N_7440,N_8391);
nand U14141 (N_14141,N_7132,N_9824);
or U14142 (N_14142,N_5951,N_5744);
xor U14143 (N_14143,N_5638,N_6033);
and U14144 (N_14144,N_8416,N_7994);
and U14145 (N_14145,N_6521,N_5042);
or U14146 (N_14146,N_7424,N_7591);
or U14147 (N_14147,N_5553,N_7942);
or U14148 (N_14148,N_5999,N_9669);
nor U14149 (N_14149,N_6065,N_8834);
nand U14150 (N_14150,N_5300,N_7437);
nand U14151 (N_14151,N_6087,N_7320);
nand U14152 (N_14152,N_7252,N_9938);
nor U14153 (N_14153,N_9209,N_8343);
nor U14154 (N_14154,N_8879,N_6202);
nor U14155 (N_14155,N_5719,N_6990);
or U14156 (N_14156,N_9023,N_8980);
and U14157 (N_14157,N_8174,N_8095);
nand U14158 (N_14158,N_6334,N_6478);
nand U14159 (N_14159,N_6651,N_8772);
nand U14160 (N_14160,N_5073,N_7178);
nand U14161 (N_14161,N_9917,N_5568);
nand U14162 (N_14162,N_7854,N_8597);
xor U14163 (N_14163,N_6654,N_9001);
nand U14164 (N_14164,N_5648,N_9294);
and U14165 (N_14165,N_8451,N_9928);
nor U14166 (N_14166,N_6871,N_9021);
nor U14167 (N_14167,N_9030,N_6759);
and U14168 (N_14168,N_8429,N_8972);
and U14169 (N_14169,N_9228,N_7238);
and U14170 (N_14170,N_9674,N_6918);
or U14171 (N_14171,N_8916,N_8997);
and U14172 (N_14172,N_8540,N_5849);
nand U14173 (N_14173,N_5850,N_9031);
nor U14174 (N_14174,N_7629,N_5641);
nor U14175 (N_14175,N_5444,N_8543);
or U14176 (N_14176,N_5382,N_7701);
and U14177 (N_14177,N_7770,N_9832);
or U14178 (N_14178,N_5744,N_9784);
or U14179 (N_14179,N_8924,N_9745);
and U14180 (N_14180,N_7761,N_9711);
xnor U14181 (N_14181,N_5670,N_7210);
and U14182 (N_14182,N_9603,N_9577);
xnor U14183 (N_14183,N_6365,N_6226);
or U14184 (N_14184,N_7065,N_8179);
and U14185 (N_14185,N_7364,N_7771);
or U14186 (N_14186,N_6945,N_6333);
nand U14187 (N_14187,N_6527,N_5932);
and U14188 (N_14188,N_5819,N_9098);
nand U14189 (N_14189,N_5846,N_5222);
or U14190 (N_14190,N_6938,N_9772);
and U14191 (N_14191,N_8865,N_9084);
nand U14192 (N_14192,N_7628,N_5943);
and U14193 (N_14193,N_8503,N_7318);
or U14194 (N_14194,N_6974,N_6363);
or U14195 (N_14195,N_6356,N_9382);
nor U14196 (N_14196,N_6294,N_8071);
nor U14197 (N_14197,N_7076,N_9061);
and U14198 (N_14198,N_8548,N_9740);
nor U14199 (N_14199,N_5108,N_7638);
and U14200 (N_14200,N_5389,N_8436);
nor U14201 (N_14201,N_5546,N_6374);
xor U14202 (N_14202,N_5658,N_5845);
nor U14203 (N_14203,N_5350,N_9254);
and U14204 (N_14204,N_6694,N_8942);
or U14205 (N_14205,N_8409,N_6782);
and U14206 (N_14206,N_7681,N_8765);
nor U14207 (N_14207,N_7062,N_8389);
xor U14208 (N_14208,N_6543,N_8873);
nor U14209 (N_14209,N_5723,N_8757);
and U14210 (N_14210,N_8655,N_5561);
and U14211 (N_14211,N_9021,N_9640);
and U14212 (N_14212,N_5619,N_8590);
and U14213 (N_14213,N_9212,N_6541);
and U14214 (N_14214,N_6788,N_5943);
nand U14215 (N_14215,N_8245,N_6387);
and U14216 (N_14216,N_6510,N_6420);
nand U14217 (N_14217,N_5962,N_7121);
and U14218 (N_14218,N_8517,N_6179);
nor U14219 (N_14219,N_5956,N_5768);
and U14220 (N_14220,N_5952,N_6347);
and U14221 (N_14221,N_5776,N_6921);
and U14222 (N_14222,N_7629,N_7983);
nand U14223 (N_14223,N_5247,N_5454);
and U14224 (N_14224,N_7835,N_9201);
nand U14225 (N_14225,N_7893,N_8130);
or U14226 (N_14226,N_7652,N_6794);
nor U14227 (N_14227,N_6749,N_7742);
xnor U14228 (N_14228,N_9291,N_9491);
nor U14229 (N_14229,N_5951,N_9824);
nand U14230 (N_14230,N_5138,N_7205);
and U14231 (N_14231,N_6307,N_5309);
or U14232 (N_14232,N_9440,N_6219);
nand U14233 (N_14233,N_7205,N_5975);
nor U14234 (N_14234,N_7885,N_9659);
and U14235 (N_14235,N_9283,N_6024);
nand U14236 (N_14236,N_9005,N_5791);
nand U14237 (N_14237,N_7269,N_6490);
and U14238 (N_14238,N_5078,N_6049);
nor U14239 (N_14239,N_8384,N_9187);
nand U14240 (N_14240,N_6376,N_5548);
nor U14241 (N_14241,N_8050,N_5097);
or U14242 (N_14242,N_5489,N_5969);
or U14243 (N_14243,N_7570,N_5313);
nand U14244 (N_14244,N_5264,N_8003);
or U14245 (N_14245,N_9367,N_5808);
and U14246 (N_14246,N_9464,N_8497);
or U14247 (N_14247,N_6851,N_6323);
or U14248 (N_14248,N_9225,N_5484);
or U14249 (N_14249,N_8015,N_7570);
nor U14250 (N_14250,N_8075,N_8973);
nor U14251 (N_14251,N_6022,N_8414);
nand U14252 (N_14252,N_7331,N_5479);
nor U14253 (N_14253,N_7486,N_5380);
or U14254 (N_14254,N_6234,N_5330);
nand U14255 (N_14255,N_6790,N_8589);
nor U14256 (N_14256,N_6178,N_9723);
or U14257 (N_14257,N_6756,N_5373);
and U14258 (N_14258,N_5121,N_8512);
nor U14259 (N_14259,N_7564,N_5537);
nand U14260 (N_14260,N_8416,N_5746);
nor U14261 (N_14261,N_7251,N_7789);
or U14262 (N_14262,N_8109,N_7063);
xnor U14263 (N_14263,N_6110,N_7638);
nand U14264 (N_14264,N_7827,N_8278);
nand U14265 (N_14265,N_8945,N_5568);
and U14266 (N_14266,N_5458,N_9814);
nor U14267 (N_14267,N_6326,N_8139);
or U14268 (N_14268,N_5019,N_6883);
or U14269 (N_14269,N_6356,N_6553);
or U14270 (N_14270,N_5538,N_9527);
nand U14271 (N_14271,N_9509,N_7368);
nand U14272 (N_14272,N_9548,N_5518);
nand U14273 (N_14273,N_5984,N_5748);
and U14274 (N_14274,N_5012,N_8918);
or U14275 (N_14275,N_9070,N_5948);
nor U14276 (N_14276,N_7843,N_5275);
nor U14277 (N_14277,N_9743,N_8413);
nor U14278 (N_14278,N_5910,N_5210);
and U14279 (N_14279,N_8196,N_7766);
and U14280 (N_14280,N_8927,N_6774);
xor U14281 (N_14281,N_6677,N_6810);
and U14282 (N_14282,N_9736,N_7873);
or U14283 (N_14283,N_6652,N_8345);
nand U14284 (N_14284,N_5758,N_7787);
and U14285 (N_14285,N_6973,N_8269);
or U14286 (N_14286,N_5116,N_5677);
xnor U14287 (N_14287,N_8688,N_7443);
or U14288 (N_14288,N_7205,N_6148);
nor U14289 (N_14289,N_5963,N_9122);
or U14290 (N_14290,N_7376,N_8636);
xor U14291 (N_14291,N_9583,N_8916);
and U14292 (N_14292,N_8159,N_7071);
xor U14293 (N_14293,N_8108,N_6772);
nand U14294 (N_14294,N_9757,N_9157);
xor U14295 (N_14295,N_8351,N_8808);
or U14296 (N_14296,N_9372,N_9343);
and U14297 (N_14297,N_8426,N_9285);
and U14298 (N_14298,N_7145,N_7056);
nor U14299 (N_14299,N_8556,N_5004);
or U14300 (N_14300,N_9046,N_5636);
or U14301 (N_14301,N_7321,N_5700);
xnor U14302 (N_14302,N_5266,N_9265);
and U14303 (N_14303,N_8318,N_8163);
nand U14304 (N_14304,N_8180,N_9190);
or U14305 (N_14305,N_9812,N_7549);
nand U14306 (N_14306,N_7480,N_5051);
nor U14307 (N_14307,N_6821,N_6063);
or U14308 (N_14308,N_8515,N_5992);
or U14309 (N_14309,N_6467,N_5507);
nand U14310 (N_14310,N_6149,N_6808);
and U14311 (N_14311,N_8841,N_5157);
and U14312 (N_14312,N_7936,N_8145);
and U14313 (N_14313,N_5918,N_6869);
nand U14314 (N_14314,N_7914,N_9275);
nor U14315 (N_14315,N_7031,N_5100);
or U14316 (N_14316,N_5666,N_7511);
or U14317 (N_14317,N_6325,N_9893);
and U14318 (N_14318,N_7471,N_9468);
or U14319 (N_14319,N_7042,N_5885);
xnor U14320 (N_14320,N_8137,N_5790);
or U14321 (N_14321,N_6057,N_7635);
nor U14322 (N_14322,N_5379,N_8641);
or U14323 (N_14323,N_6625,N_6339);
and U14324 (N_14324,N_6242,N_5322);
or U14325 (N_14325,N_8526,N_6999);
and U14326 (N_14326,N_5747,N_9444);
xor U14327 (N_14327,N_8773,N_5199);
nor U14328 (N_14328,N_9181,N_9570);
or U14329 (N_14329,N_8899,N_5488);
nand U14330 (N_14330,N_9335,N_7113);
nand U14331 (N_14331,N_8065,N_7561);
xnor U14332 (N_14332,N_9900,N_9322);
xor U14333 (N_14333,N_9643,N_5788);
and U14334 (N_14334,N_8272,N_9698);
and U14335 (N_14335,N_7381,N_6978);
or U14336 (N_14336,N_9671,N_7370);
or U14337 (N_14337,N_5425,N_9144);
or U14338 (N_14338,N_7968,N_9508);
or U14339 (N_14339,N_7497,N_6641);
and U14340 (N_14340,N_8848,N_6411);
nand U14341 (N_14341,N_5057,N_6780);
xnor U14342 (N_14342,N_8686,N_8885);
nor U14343 (N_14343,N_8207,N_7041);
and U14344 (N_14344,N_8231,N_5958);
or U14345 (N_14345,N_8199,N_7842);
xor U14346 (N_14346,N_6280,N_9188);
or U14347 (N_14347,N_5168,N_8342);
or U14348 (N_14348,N_8556,N_7851);
and U14349 (N_14349,N_9270,N_9637);
xor U14350 (N_14350,N_6309,N_5903);
nor U14351 (N_14351,N_6794,N_6581);
nand U14352 (N_14352,N_6311,N_6776);
nand U14353 (N_14353,N_9501,N_6081);
nand U14354 (N_14354,N_5091,N_5065);
and U14355 (N_14355,N_8199,N_8474);
nand U14356 (N_14356,N_9024,N_5202);
or U14357 (N_14357,N_6217,N_9464);
xor U14358 (N_14358,N_5688,N_7559);
and U14359 (N_14359,N_6701,N_7391);
and U14360 (N_14360,N_6401,N_7087);
nand U14361 (N_14361,N_9649,N_6665);
nor U14362 (N_14362,N_5134,N_6364);
nand U14363 (N_14363,N_6412,N_5522);
nand U14364 (N_14364,N_5424,N_7874);
and U14365 (N_14365,N_5047,N_7086);
or U14366 (N_14366,N_5366,N_6204);
and U14367 (N_14367,N_9292,N_5011);
xor U14368 (N_14368,N_7609,N_8557);
xor U14369 (N_14369,N_9268,N_6510);
nor U14370 (N_14370,N_9245,N_9437);
nor U14371 (N_14371,N_6931,N_9010);
and U14372 (N_14372,N_5588,N_6466);
or U14373 (N_14373,N_5459,N_6961);
xnor U14374 (N_14374,N_5737,N_6739);
nand U14375 (N_14375,N_8345,N_8810);
nor U14376 (N_14376,N_6894,N_5399);
and U14377 (N_14377,N_9341,N_5363);
xnor U14378 (N_14378,N_5267,N_6376);
and U14379 (N_14379,N_7352,N_5269);
xor U14380 (N_14380,N_8481,N_9780);
or U14381 (N_14381,N_8653,N_7899);
nand U14382 (N_14382,N_6457,N_5931);
or U14383 (N_14383,N_9837,N_5780);
nor U14384 (N_14384,N_5453,N_7322);
nor U14385 (N_14385,N_6452,N_5451);
or U14386 (N_14386,N_5166,N_7131);
or U14387 (N_14387,N_7053,N_9689);
nor U14388 (N_14388,N_9825,N_5238);
nor U14389 (N_14389,N_5704,N_8942);
and U14390 (N_14390,N_7596,N_9190);
or U14391 (N_14391,N_7022,N_6057);
nand U14392 (N_14392,N_9002,N_5408);
or U14393 (N_14393,N_7039,N_6996);
and U14394 (N_14394,N_5910,N_5823);
or U14395 (N_14395,N_6619,N_6134);
or U14396 (N_14396,N_6348,N_9799);
or U14397 (N_14397,N_9633,N_6814);
nor U14398 (N_14398,N_9411,N_5951);
nor U14399 (N_14399,N_6748,N_9076);
nand U14400 (N_14400,N_8865,N_6698);
nand U14401 (N_14401,N_9385,N_7173);
and U14402 (N_14402,N_9786,N_9950);
and U14403 (N_14403,N_9578,N_5918);
or U14404 (N_14404,N_5616,N_5428);
nor U14405 (N_14405,N_9233,N_9250);
xor U14406 (N_14406,N_9792,N_7910);
or U14407 (N_14407,N_6968,N_7924);
nor U14408 (N_14408,N_6737,N_6795);
nand U14409 (N_14409,N_8559,N_6285);
and U14410 (N_14410,N_7441,N_5705);
nor U14411 (N_14411,N_9505,N_7498);
nor U14412 (N_14412,N_8662,N_9603);
and U14413 (N_14413,N_7651,N_6097);
and U14414 (N_14414,N_8346,N_8084);
xnor U14415 (N_14415,N_5270,N_6658);
nor U14416 (N_14416,N_5769,N_6335);
and U14417 (N_14417,N_8835,N_7102);
and U14418 (N_14418,N_7082,N_5835);
nand U14419 (N_14419,N_5941,N_9856);
nand U14420 (N_14420,N_9333,N_7224);
nor U14421 (N_14421,N_6715,N_5273);
xnor U14422 (N_14422,N_7641,N_6545);
or U14423 (N_14423,N_8195,N_8327);
nor U14424 (N_14424,N_5540,N_8507);
nor U14425 (N_14425,N_9195,N_9032);
xor U14426 (N_14426,N_8649,N_6706);
or U14427 (N_14427,N_8710,N_9894);
or U14428 (N_14428,N_5944,N_7167);
or U14429 (N_14429,N_8101,N_5368);
and U14430 (N_14430,N_9231,N_5887);
or U14431 (N_14431,N_5320,N_9105);
and U14432 (N_14432,N_8736,N_8729);
nor U14433 (N_14433,N_6782,N_9715);
xnor U14434 (N_14434,N_9593,N_9130);
nand U14435 (N_14435,N_9388,N_7776);
nand U14436 (N_14436,N_9091,N_7512);
or U14437 (N_14437,N_5850,N_6681);
and U14438 (N_14438,N_8917,N_7520);
nand U14439 (N_14439,N_5004,N_6385);
nor U14440 (N_14440,N_9152,N_9675);
nor U14441 (N_14441,N_7627,N_6177);
nor U14442 (N_14442,N_7482,N_8651);
nand U14443 (N_14443,N_7523,N_9668);
and U14444 (N_14444,N_7917,N_7956);
nand U14445 (N_14445,N_5693,N_5898);
nor U14446 (N_14446,N_5277,N_5619);
and U14447 (N_14447,N_6513,N_8458);
and U14448 (N_14448,N_7215,N_7512);
xnor U14449 (N_14449,N_5945,N_5224);
or U14450 (N_14450,N_5857,N_7514);
or U14451 (N_14451,N_9987,N_5827);
and U14452 (N_14452,N_9436,N_9848);
or U14453 (N_14453,N_9978,N_7672);
nand U14454 (N_14454,N_7506,N_5039);
nor U14455 (N_14455,N_5671,N_9751);
nand U14456 (N_14456,N_8777,N_7648);
or U14457 (N_14457,N_8553,N_9652);
or U14458 (N_14458,N_9342,N_7317);
nand U14459 (N_14459,N_6410,N_8128);
or U14460 (N_14460,N_8995,N_9007);
nor U14461 (N_14461,N_6586,N_7184);
xor U14462 (N_14462,N_6578,N_8769);
nand U14463 (N_14463,N_7101,N_6848);
nand U14464 (N_14464,N_6563,N_5555);
xor U14465 (N_14465,N_5052,N_6391);
nand U14466 (N_14466,N_7539,N_6195);
and U14467 (N_14467,N_6848,N_8143);
nor U14468 (N_14468,N_5168,N_5774);
nor U14469 (N_14469,N_7413,N_7374);
nand U14470 (N_14470,N_6802,N_7663);
nor U14471 (N_14471,N_8388,N_5676);
nand U14472 (N_14472,N_6761,N_7734);
nand U14473 (N_14473,N_8604,N_6966);
nor U14474 (N_14474,N_9458,N_9819);
or U14475 (N_14475,N_6157,N_8755);
nor U14476 (N_14476,N_5647,N_5358);
or U14477 (N_14477,N_5912,N_7157);
nor U14478 (N_14478,N_9935,N_8044);
nor U14479 (N_14479,N_5164,N_6671);
and U14480 (N_14480,N_8099,N_9079);
nand U14481 (N_14481,N_7889,N_7211);
nand U14482 (N_14482,N_5526,N_8473);
xnor U14483 (N_14483,N_7832,N_9637);
nor U14484 (N_14484,N_9458,N_6698);
and U14485 (N_14485,N_9063,N_9303);
or U14486 (N_14486,N_7801,N_5829);
and U14487 (N_14487,N_6374,N_6787);
or U14488 (N_14488,N_7995,N_8406);
and U14489 (N_14489,N_5712,N_7454);
nor U14490 (N_14490,N_7625,N_8385);
or U14491 (N_14491,N_7694,N_9750);
or U14492 (N_14492,N_7567,N_7931);
or U14493 (N_14493,N_6178,N_5013);
or U14494 (N_14494,N_7862,N_9807);
nor U14495 (N_14495,N_8505,N_5983);
nor U14496 (N_14496,N_5749,N_9967);
and U14497 (N_14497,N_7358,N_8333);
nand U14498 (N_14498,N_5153,N_7329);
nand U14499 (N_14499,N_8305,N_5852);
and U14500 (N_14500,N_7231,N_9410);
or U14501 (N_14501,N_6649,N_6772);
and U14502 (N_14502,N_9693,N_7031);
nor U14503 (N_14503,N_7697,N_6949);
nand U14504 (N_14504,N_5467,N_5968);
or U14505 (N_14505,N_8299,N_6756);
or U14506 (N_14506,N_9778,N_9743);
xnor U14507 (N_14507,N_9646,N_5660);
and U14508 (N_14508,N_7098,N_8682);
or U14509 (N_14509,N_5296,N_9194);
and U14510 (N_14510,N_5724,N_7384);
xnor U14511 (N_14511,N_6786,N_7798);
and U14512 (N_14512,N_5864,N_9735);
and U14513 (N_14513,N_5223,N_8981);
xnor U14514 (N_14514,N_5867,N_9059);
nand U14515 (N_14515,N_7229,N_5887);
or U14516 (N_14516,N_6558,N_9315);
or U14517 (N_14517,N_5969,N_9846);
nor U14518 (N_14518,N_8089,N_5442);
nor U14519 (N_14519,N_5392,N_5939);
and U14520 (N_14520,N_9585,N_5014);
nor U14521 (N_14521,N_8060,N_6602);
and U14522 (N_14522,N_9210,N_6636);
or U14523 (N_14523,N_8836,N_6893);
or U14524 (N_14524,N_7783,N_9162);
nand U14525 (N_14525,N_8447,N_6979);
nand U14526 (N_14526,N_6993,N_6418);
nor U14527 (N_14527,N_7749,N_7978);
or U14528 (N_14528,N_5203,N_5879);
nand U14529 (N_14529,N_6231,N_7965);
xnor U14530 (N_14530,N_7375,N_9472);
xnor U14531 (N_14531,N_5776,N_6670);
and U14532 (N_14532,N_9158,N_9862);
or U14533 (N_14533,N_8621,N_5018);
and U14534 (N_14534,N_7175,N_7820);
or U14535 (N_14535,N_7938,N_9688);
or U14536 (N_14536,N_8575,N_8185);
and U14537 (N_14537,N_5321,N_6288);
or U14538 (N_14538,N_9734,N_6890);
or U14539 (N_14539,N_5718,N_5123);
and U14540 (N_14540,N_9726,N_8716);
or U14541 (N_14541,N_5818,N_9191);
xnor U14542 (N_14542,N_5134,N_9543);
or U14543 (N_14543,N_5863,N_8803);
nand U14544 (N_14544,N_8261,N_9133);
and U14545 (N_14545,N_5432,N_7216);
and U14546 (N_14546,N_6671,N_7357);
or U14547 (N_14547,N_7354,N_5213);
nor U14548 (N_14548,N_7340,N_6826);
xnor U14549 (N_14549,N_9565,N_5002);
and U14550 (N_14550,N_6078,N_7374);
or U14551 (N_14551,N_5160,N_6480);
nand U14552 (N_14552,N_5702,N_8903);
nand U14553 (N_14553,N_7230,N_8486);
or U14554 (N_14554,N_7674,N_7086);
nor U14555 (N_14555,N_5221,N_7080);
nor U14556 (N_14556,N_8142,N_5897);
nand U14557 (N_14557,N_7547,N_7118);
nor U14558 (N_14558,N_6121,N_8167);
or U14559 (N_14559,N_5454,N_9916);
and U14560 (N_14560,N_5760,N_8316);
nand U14561 (N_14561,N_6578,N_8827);
nand U14562 (N_14562,N_5560,N_7258);
or U14563 (N_14563,N_5738,N_5537);
nand U14564 (N_14564,N_9586,N_8367);
xor U14565 (N_14565,N_7753,N_9501);
and U14566 (N_14566,N_6869,N_9061);
nor U14567 (N_14567,N_6256,N_5372);
nor U14568 (N_14568,N_5865,N_8643);
nand U14569 (N_14569,N_5157,N_6204);
or U14570 (N_14570,N_5440,N_8253);
nor U14571 (N_14571,N_6769,N_9179);
and U14572 (N_14572,N_5797,N_6953);
xnor U14573 (N_14573,N_7656,N_6444);
nand U14574 (N_14574,N_5250,N_6359);
nor U14575 (N_14575,N_9021,N_5201);
and U14576 (N_14576,N_8377,N_6086);
nor U14577 (N_14577,N_5272,N_6864);
and U14578 (N_14578,N_8539,N_7902);
nor U14579 (N_14579,N_8975,N_9773);
nor U14580 (N_14580,N_6655,N_7572);
nor U14581 (N_14581,N_7594,N_9745);
and U14582 (N_14582,N_7031,N_8870);
nand U14583 (N_14583,N_7075,N_9468);
or U14584 (N_14584,N_5677,N_6435);
or U14585 (N_14585,N_7130,N_7490);
nand U14586 (N_14586,N_8250,N_6426);
and U14587 (N_14587,N_5034,N_8020);
and U14588 (N_14588,N_7868,N_6044);
or U14589 (N_14589,N_5926,N_9418);
or U14590 (N_14590,N_7398,N_9245);
nand U14591 (N_14591,N_6057,N_5492);
and U14592 (N_14592,N_5053,N_5753);
and U14593 (N_14593,N_5906,N_8043);
nand U14594 (N_14594,N_9176,N_5630);
nor U14595 (N_14595,N_8165,N_7252);
and U14596 (N_14596,N_8051,N_7811);
nand U14597 (N_14597,N_8661,N_6099);
and U14598 (N_14598,N_9572,N_5107);
or U14599 (N_14599,N_7131,N_7467);
or U14600 (N_14600,N_6953,N_8191);
xnor U14601 (N_14601,N_7360,N_9673);
nand U14602 (N_14602,N_9401,N_5619);
or U14603 (N_14603,N_6771,N_9190);
or U14604 (N_14604,N_9433,N_7191);
nand U14605 (N_14605,N_6396,N_8306);
and U14606 (N_14606,N_6218,N_8806);
xor U14607 (N_14607,N_6674,N_8196);
xor U14608 (N_14608,N_9662,N_8169);
xor U14609 (N_14609,N_5861,N_7522);
and U14610 (N_14610,N_6420,N_9232);
and U14611 (N_14611,N_7055,N_8787);
nand U14612 (N_14612,N_5431,N_8863);
or U14613 (N_14613,N_5271,N_6033);
xor U14614 (N_14614,N_7816,N_6032);
xor U14615 (N_14615,N_8925,N_8999);
and U14616 (N_14616,N_9789,N_8159);
or U14617 (N_14617,N_9918,N_9014);
nand U14618 (N_14618,N_7059,N_7530);
and U14619 (N_14619,N_8189,N_6594);
or U14620 (N_14620,N_5405,N_9446);
nor U14621 (N_14621,N_6351,N_7842);
xnor U14622 (N_14622,N_6654,N_5709);
or U14623 (N_14623,N_5232,N_6450);
nor U14624 (N_14624,N_7588,N_7096);
and U14625 (N_14625,N_6839,N_8550);
or U14626 (N_14626,N_9856,N_8469);
and U14627 (N_14627,N_7215,N_9064);
nand U14628 (N_14628,N_6044,N_9086);
nor U14629 (N_14629,N_6210,N_9237);
or U14630 (N_14630,N_5156,N_9587);
nor U14631 (N_14631,N_6723,N_9257);
and U14632 (N_14632,N_6284,N_8444);
nand U14633 (N_14633,N_6141,N_9704);
and U14634 (N_14634,N_5496,N_6813);
xor U14635 (N_14635,N_6176,N_8399);
or U14636 (N_14636,N_9821,N_8416);
nand U14637 (N_14637,N_8179,N_9226);
or U14638 (N_14638,N_6935,N_9884);
nor U14639 (N_14639,N_8162,N_5587);
nand U14640 (N_14640,N_9388,N_7618);
nand U14641 (N_14641,N_6907,N_8439);
or U14642 (N_14642,N_7524,N_8974);
or U14643 (N_14643,N_5941,N_9248);
and U14644 (N_14644,N_7251,N_5819);
and U14645 (N_14645,N_9435,N_7078);
and U14646 (N_14646,N_5450,N_7193);
nand U14647 (N_14647,N_6936,N_7803);
nand U14648 (N_14648,N_5637,N_8725);
or U14649 (N_14649,N_9883,N_7358);
xor U14650 (N_14650,N_8037,N_5373);
or U14651 (N_14651,N_6806,N_6781);
or U14652 (N_14652,N_9504,N_5407);
nor U14653 (N_14653,N_5636,N_8816);
or U14654 (N_14654,N_6410,N_5509);
and U14655 (N_14655,N_7835,N_8683);
or U14656 (N_14656,N_9482,N_8984);
or U14657 (N_14657,N_6940,N_8961);
nand U14658 (N_14658,N_7018,N_9501);
nand U14659 (N_14659,N_6558,N_8420);
or U14660 (N_14660,N_8914,N_7729);
nand U14661 (N_14661,N_6918,N_6323);
nor U14662 (N_14662,N_5906,N_5573);
nand U14663 (N_14663,N_6459,N_7918);
nor U14664 (N_14664,N_9326,N_5172);
xor U14665 (N_14665,N_7543,N_7300);
nand U14666 (N_14666,N_7755,N_7992);
and U14667 (N_14667,N_8055,N_5157);
nand U14668 (N_14668,N_9355,N_8010);
xnor U14669 (N_14669,N_9432,N_5657);
or U14670 (N_14670,N_6128,N_8209);
nand U14671 (N_14671,N_9570,N_7910);
nand U14672 (N_14672,N_9028,N_8390);
nor U14673 (N_14673,N_6174,N_8168);
or U14674 (N_14674,N_6699,N_5703);
and U14675 (N_14675,N_6834,N_9400);
and U14676 (N_14676,N_5305,N_9199);
nor U14677 (N_14677,N_8929,N_5061);
or U14678 (N_14678,N_8146,N_9619);
nor U14679 (N_14679,N_8855,N_7014);
nand U14680 (N_14680,N_6673,N_8178);
and U14681 (N_14681,N_6395,N_5397);
xnor U14682 (N_14682,N_6740,N_8366);
or U14683 (N_14683,N_6288,N_6316);
or U14684 (N_14684,N_5505,N_5724);
and U14685 (N_14685,N_6843,N_5215);
and U14686 (N_14686,N_7842,N_6653);
nor U14687 (N_14687,N_6851,N_8389);
nand U14688 (N_14688,N_8934,N_6103);
and U14689 (N_14689,N_9318,N_8913);
or U14690 (N_14690,N_5870,N_9459);
nand U14691 (N_14691,N_6945,N_8767);
and U14692 (N_14692,N_9074,N_8785);
or U14693 (N_14693,N_8446,N_8281);
xor U14694 (N_14694,N_5664,N_8741);
and U14695 (N_14695,N_8819,N_8760);
nand U14696 (N_14696,N_6577,N_5031);
nand U14697 (N_14697,N_5588,N_9905);
or U14698 (N_14698,N_5577,N_9713);
or U14699 (N_14699,N_7986,N_7463);
or U14700 (N_14700,N_6230,N_7615);
or U14701 (N_14701,N_8916,N_5178);
nor U14702 (N_14702,N_5276,N_6444);
nor U14703 (N_14703,N_5205,N_9389);
or U14704 (N_14704,N_5138,N_8379);
xor U14705 (N_14705,N_5860,N_6348);
nand U14706 (N_14706,N_5112,N_7191);
and U14707 (N_14707,N_5128,N_5492);
nand U14708 (N_14708,N_6008,N_8371);
nand U14709 (N_14709,N_9444,N_7686);
nand U14710 (N_14710,N_7205,N_9480);
and U14711 (N_14711,N_9428,N_8892);
xor U14712 (N_14712,N_8178,N_8272);
or U14713 (N_14713,N_5709,N_5330);
xor U14714 (N_14714,N_9617,N_8378);
and U14715 (N_14715,N_6790,N_7272);
nand U14716 (N_14716,N_9659,N_5810);
nor U14717 (N_14717,N_9822,N_9501);
and U14718 (N_14718,N_9605,N_9731);
and U14719 (N_14719,N_8092,N_7581);
or U14720 (N_14720,N_7227,N_8031);
nor U14721 (N_14721,N_5380,N_5946);
and U14722 (N_14722,N_8766,N_8010);
nand U14723 (N_14723,N_8692,N_9111);
or U14724 (N_14724,N_6949,N_6504);
nor U14725 (N_14725,N_9514,N_9980);
or U14726 (N_14726,N_7909,N_5349);
nor U14727 (N_14727,N_8935,N_6056);
xor U14728 (N_14728,N_9477,N_8614);
nor U14729 (N_14729,N_9882,N_8450);
nor U14730 (N_14730,N_8647,N_5398);
xnor U14731 (N_14731,N_7278,N_5211);
nor U14732 (N_14732,N_6118,N_8295);
nor U14733 (N_14733,N_5056,N_8209);
or U14734 (N_14734,N_9216,N_8112);
nor U14735 (N_14735,N_8664,N_8554);
and U14736 (N_14736,N_7018,N_7946);
nor U14737 (N_14737,N_5699,N_7829);
and U14738 (N_14738,N_5172,N_8107);
or U14739 (N_14739,N_7905,N_8544);
and U14740 (N_14740,N_9336,N_7718);
nand U14741 (N_14741,N_8336,N_7090);
nor U14742 (N_14742,N_7090,N_8193);
nand U14743 (N_14743,N_9749,N_5409);
and U14744 (N_14744,N_6363,N_8118);
and U14745 (N_14745,N_6754,N_5401);
nand U14746 (N_14746,N_9501,N_6402);
or U14747 (N_14747,N_5921,N_9006);
or U14748 (N_14748,N_6510,N_8454);
nor U14749 (N_14749,N_7779,N_6666);
and U14750 (N_14750,N_8020,N_9470);
xnor U14751 (N_14751,N_5934,N_9706);
nand U14752 (N_14752,N_5135,N_9758);
and U14753 (N_14753,N_6129,N_6437);
and U14754 (N_14754,N_5546,N_6694);
xor U14755 (N_14755,N_6669,N_8679);
nor U14756 (N_14756,N_9031,N_5405);
nand U14757 (N_14757,N_8703,N_8479);
and U14758 (N_14758,N_6266,N_6747);
and U14759 (N_14759,N_6647,N_5042);
or U14760 (N_14760,N_8484,N_9634);
nand U14761 (N_14761,N_5920,N_6664);
or U14762 (N_14762,N_5612,N_5691);
or U14763 (N_14763,N_7865,N_8137);
nand U14764 (N_14764,N_7555,N_8863);
or U14765 (N_14765,N_6318,N_8001);
and U14766 (N_14766,N_9914,N_7887);
nor U14767 (N_14767,N_8124,N_5099);
or U14768 (N_14768,N_6177,N_6162);
xor U14769 (N_14769,N_6889,N_7337);
or U14770 (N_14770,N_8342,N_9719);
and U14771 (N_14771,N_8694,N_9752);
nand U14772 (N_14772,N_8420,N_5099);
and U14773 (N_14773,N_6420,N_6740);
or U14774 (N_14774,N_7557,N_8824);
and U14775 (N_14775,N_8171,N_9336);
and U14776 (N_14776,N_8538,N_6515);
nor U14777 (N_14777,N_8295,N_9262);
nand U14778 (N_14778,N_8953,N_6445);
or U14779 (N_14779,N_6177,N_7770);
and U14780 (N_14780,N_5436,N_7033);
nand U14781 (N_14781,N_5966,N_5426);
and U14782 (N_14782,N_5554,N_7363);
and U14783 (N_14783,N_5048,N_9685);
or U14784 (N_14784,N_6723,N_5979);
nand U14785 (N_14785,N_6819,N_6426);
or U14786 (N_14786,N_5796,N_7931);
and U14787 (N_14787,N_7483,N_5244);
and U14788 (N_14788,N_9194,N_5238);
or U14789 (N_14789,N_5052,N_8196);
and U14790 (N_14790,N_9554,N_5740);
xor U14791 (N_14791,N_8922,N_5551);
nand U14792 (N_14792,N_8012,N_5949);
xnor U14793 (N_14793,N_5092,N_5287);
or U14794 (N_14794,N_7842,N_5500);
and U14795 (N_14795,N_6048,N_7129);
and U14796 (N_14796,N_7248,N_8010);
nand U14797 (N_14797,N_8053,N_8080);
nor U14798 (N_14798,N_6035,N_7120);
nand U14799 (N_14799,N_7826,N_5705);
and U14800 (N_14800,N_6824,N_5334);
nand U14801 (N_14801,N_5098,N_8759);
and U14802 (N_14802,N_5529,N_8739);
or U14803 (N_14803,N_5303,N_7035);
nand U14804 (N_14804,N_9917,N_6060);
nor U14805 (N_14805,N_8244,N_6348);
or U14806 (N_14806,N_5335,N_7687);
or U14807 (N_14807,N_9795,N_7781);
and U14808 (N_14808,N_8986,N_7645);
or U14809 (N_14809,N_6766,N_9468);
and U14810 (N_14810,N_7335,N_5853);
nor U14811 (N_14811,N_9254,N_9169);
nor U14812 (N_14812,N_6006,N_8268);
or U14813 (N_14813,N_5864,N_8600);
or U14814 (N_14814,N_6928,N_8187);
xnor U14815 (N_14815,N_8006,N_8973);
nand U14816 (N_14816,N_9319,N_6191);
nor U14817 (N_14817,N_5471,N_7977);
or U14818 (N_14818,N_8496,N_8930);
xnor U14819 (N_14819,N_6724,N_8668);
nor U14820 (N_14820,N_7609,N_6668);
or U14821 (N_14821,N_6840,N_8909);
and U14822 (N_14822,N_7739,N_6368);
nor U14823 (N_14823,N_8833,N_7688);
nor U14824 (N_14824,N_5019,N_6104);
or U14825 (N_14825,N_5714,N_9755);
and U14826 (N_14826,N_8877,N_6889);
nor U14827 (N_14827,N_6697,N_6206);
nand U14828 (N_14828,N_6702,N_8358);
or U14829 (N_14829,N_7125,N_7980);
nand U14830 (N_14830,N_6024,N_7367);
or U14831 (N_14831,N_6725,N_9082);
nor U14832 (N_14832,N_9740,N_8194);
and U14833 (N_14833,N_6739,N_5187);
nor U14834 (N_14834,N_8487,N_6508);
nand U14835 (N_14835,N_9785,N_6390);
or U14836 (N_14836,N_9966,N_8767);
nand U14837 (N_14837,N_7376,N_7613);
nor U14838 (N_14838,N_5075,N_6452);
and U14839 (N_14839,N_9157,N_7791);
or U14840 (N_14840,N_9016,N_8969);
and U14841 (N_14841,N_6202,N_5233);
or U14842 (N_14842,N_5726,N_5847);
and U14843 (N_14843,N_8855,N_7843);
and U14844 (N_14844,N_5886,N_7995);
or U14845 (N_14845,N_8484,N_7137);
nand U14846 (N_14846,N_5691,N_7990);
nor U14847 (N_14847,N_6268,N_6717);
xor U14848 (N_14848,N_5376,N_9530);
and U14849 (N_14849,N_9568,N_9654);
or U14850 (N_14850,N_6463,N_5060);
nand U14851 (N_14851,N_9526,N_6272);
or U14852 (N_14852,N_7109,N_6490);
and U14853 (N_14853,N_5405,N_9940);
and U14854 (N_14854,N_5384,N_5535);
and U14855 (N_14855,N_9080,N_8332);
and U14856 (N_14856,N_9993,N_5997);
or U14857 (N_14857,N_6389,N_9948);
and U14858 (N_14858,N_8167,N_8682);
nor U14859 (N_14859,N_9218,N_6154);
nor U14860 (N_14860,N_6035,N_6244);
nand U14861 (N_14861,N_5383,N_5672);
or U14862 (N_14862,N_8303,N_7199);
xnor U14863 (N_14863,N_8699,N_9085);
nor U14864 (N_14864,N_5863,N_8371);
nor U14865 (N_14865,N_5393,N_8566);
or U14866 (N_14866,N_9378,N_8637);
and U14867 (N_14867,N_5695,N_8296);
or U14868 (N_14868,N_8566,N_5958);
nor U14869 (N_14869,N_9336,N_6331);
or U14870 (N_14870,N_5916,N_9391);
or U14871 (N_14871,N_8906,N_9029);
nand U14872 (N_14872,N_8494,N_6391);
and U14873 (N_14873,N_6237,N_8109);
nor U14874 (N_14874,N_9039,N_7978);
nand U14875 (N_14875,N_5955,N_9107);
or U14876 (N_14876,N_5489,N_9636);
nor U14877 (N_14877,N_9607,N_9939);
xnor U14878 (N_14878,N_5590,N_8225);
xnor U14879 (N_14879,N_8552,N_6126);
and U14880 (N_14880,N_9743,N_5922);
nor U14881 (N_14881,N_8649,N_8421);
or U14882 (N_14882,N_6880,N_5621);
or U14883 (N_14883,N_5408,N_9867);
or U14884 (N_14884,N_7694,N_8035);
xor U14885 (N_14885,N_9053,N_6937);
nand U14886 (N_14886,N_6726,N_9374);
nor U14887 (N_14887,N_8540,N_6697);
xnor U14888 (N_14888,N_7385,N_9435);
and U14889 (N_14889,N_7659,N_6036);
nor U14890 (N_14890,N_9643,N_6751);
or U14891 (N_14891,N_5039,N_9948);
xor U14892 (N_14892,N_6332,N_5813);
nand U14893 (N_14893,N_5434,N_7588);
nor U14894 (N_14894,N_9393,N_5282);
or U14895 (N_14895,N_5757,N_8624);
and U14896 (N_14896,N_7495,N_7325);
nor U14897 (N_14897,N_9512,N_5325);
or U14898 (N_14898,N_7423,N_6618);
or U14899 (N_14899,N_8571,N_5405);
or U14900 (N_14900,N_7217,N_6222);
nor U14901 (N_14901,N_6072,N_8069);
nor U14902 (N_14902,N_7082,N_9436);
or U14903 (N_14903,N_6895,N_6907);
nor U14904 (N_14904,N_9902,N_7143);
and U14905 (N_14905,N_6224,N_6601);
nand U14906 (N_14906,N_6622,N_8622);
or U14907 (N_14907,N_6243,N_9168);
or U14908 (N_14908,N_8010,N_6673);
xor U14909 (N_14909,N_6334,N_8606);
or U14910 (N_14910,N_8178,N_7133);
nor U14911 (N_14911,N_7363,N_5891);
and U14912 (N_14912,N_5930,N_5821);
or U14913 (N_14913,N_7889,N_5699);
nor U14914 (N_14914,N_6288,N_7492);
xor U14915 (N_14915,N_6553,N_9249);
nor U14916 (N_14916,N_8267,N_5693);
or U14917 (N_14917,N_7762,N_7283);
xor U14918 (N_14918,N_6744,N_5567);
and U14919 (N_14919,N_8548,N_6054);
and U14920 (N_14920,N_6228,N_5120);
nor U14921 (N_14921,N_5046,N_8644);
or U14922 (N_14922,N_7656,N_7493);
nand U14923 (N_14923,N_8602,N_7967);
and U14924 (N_14924,N_8169,N_5871);
nor U14925 (N_14925,N_8196,N_5502);
or U14926 (N_14926,N_9596,N_8418);
nor U14927 (N_14927,N_9113,N_6265);
xor U14928 (N_14928,N_6408,N_7816);
xnor U14929 (N_14929,N_7762,N_5270);
nor U14930 (N_14930,N_5113,N_5107);
or U14931 (N_14931,N_5059,N_6114);
and U14932 (N_14932,N_7800,N_9929);
xnor U14933 (N_14933,N_7584,N_9165);
or U14934 (N_14934,N_6762,N_7416);
nor U14935 (N_14935,N_7148,N_9326);
nand U14936 (N_14936,N_9162,N_8085);
nor U14937 (N_14937,N_9166,N_6619);
nor U14938 (N_14938,N_6837,N_8870);
xor U14939 (N_14939,N_6249,N_6465);
nor U14940 (N_14940,N_8080,N_7400);
nand U14941 (N_14941,N_5228,N_5110);
or U14942 (N_14942,N_6130,N_6557);
nand U14943 (N_14943,N_9514,N_5944);
nor U14944 (N_14944,N_9496,N_6696);
nor U14945 (N_14945,N_9226,N_9639);
nand U14946 (N_14946,N_8484,N_8599);
xor U14947 (N_14947,N_5623,N_6576);
nand U14948 (N_14948,N_7152,N_8748);
or U14949 (N_14949,N_9124,N_8634);
nor U14950 (N_14950,N_8898,N_9016);
and U14951 (N_14951,N_6112,N_7390);
xnor U14952 (N_14952,N_5812,N_6685);
and U14953 (N_14953,N_8848,N_5956);
nand U14954 (N_14954,N_5002,N_9986);
xor U14955 (N_14955,N_7524,N_6645);
or U14956 (N_14956,N_6069,N_8888);
or U14957 (N_14957,N_6728,N_7514);
nor U14958 (N_14958,N_7431,N_8028);
nand U14959 (N_14959,N_8826,N_6374);
or U14960 (N_14960,N_8391,N_6739);
nor U14961 (N_14961,N_9329,N_6067);
xnor U14962 (N_14962,N_8161,N_7929);
xnor U14963 (N_14963,N_5873,N_7505);
or U14964 (N_14964,N_9331,N_5953);
nor U14965 (N_14965,N_6220,N_8093);
or U14966 (N_14966,N_6875,N_7498);
xnor U14967 (N_14967,N_5236,N_9754);
and U14968 (N_14968,N_6381,N_5430);
nand U14969 (N_14969,N_6500,N_9935);
nand U14970 (N_14970,N_6953,N_5447);
or U14971 (N_14971,N_5060,N_8640);
nor U14972 (N_14972,N_6721,N_8290);
nor U14973 (N_14973,N_5170,N_8556);
xnor U14974 (N_14974,N_7365,N_8045);
or U14975 (N_14975,N_7018,N_9198);
nand U14976 (N_14976,N_7891,N_8725);
nand U14977 (N_14977,N_9215,N_9100);
and U14978 (N_14978,N_8413,N_5839);
and U14979 (N_14979,N_9898,N_8058);
xnor U14980 (N_14980,N_5071,N_8762);
nor U14981 (N_14981,N_8872,N_9771);
and U14982 (N_14982,N_9913,N_7040);
nand U14983 (N_14983,N_9719,N_9765);
nand U14984 (N_14984,N_7322,N_5473);
nor U14985 (N_14985,N_6992,N_6273);
and U14986 (N_14986,N_9146,N_5015);
and U14987 (N_14987,N_5671,N_9550);
nor U14988 (N_14988,N_6706,N_6468);
or U14989 (N_14989,N_5570,N_6451);
xor U14990 (N_14990,N_7465,N_6411);
xnor U14991 (N_14991,N_8316,N_6051);
or U14992 (N_14992,N_5971,N_9107);
xor U14993 (N_14993,N_6275,N_8334);
nor U14994 (N_14994,N_6674,N_8801);
and U14995 (N_14995,N_6066,N_5132);
or U14996 (N_14996,N_8211,N_7109);
and U14997 (N_14997,N_8015,N_7352);
and U14998 (N_14998,N_9071,N_8393);
or U14999 (N_14999,N_5580,N_6033);
nand UO_0 (O_0,N_10023,N_14888);
nor UO_1 (O_1,N_13824,N_12574);
nand UO_2 (O_2,N_10921,N_12590);
or UO_3 (O_3,N_13290,N_11687);
and UO_4 (O_4,N_14180,N_11479);
nor UO_5 (O_5,N_10999,N_13461);
nand UO_6 (O_6,N_14796,N_12551);
nor UO_7 (O_7,N_11347,N_11926);
and UO_8 (O_8,N_12595,N_12358);
nand UO_9 (O_9,N_12132,N_13894);
or UO_10 (O_10,N_11706,N_14355);
nand UO_11 (O_11,N_10404,N_11741);
nor UO_12 (O_12,N_12429,N_11048);
and UO_13 (O_13,N_14605,N_14498);
or UO_14 (O_14,N_10277,N_11950);
nand UO_15 (O_15,N_10082,N_12219);
or UO_16 (O_16,N_11498,N_14816);
or UO_17 (O_17,N_12710,N_11744);
and UO_18 (O_18,N_12143,N_14442);
nor UO_19 (O_19,N_13495,N_11276);
xor UO_20 (O_20,N_13336,N_10775);
or UO_21 (O_21,N_13718,N_12999);
and UO_22 (O_22,N_12950,N_13086);
or UO_23 (O_23,N_12077,N_10294);
nor UO_24 (O_24,N_11110,N_12631);
or UO_25 (O_25,N_14099,N_14366);
or UO_26 (O_26,N_11337,N_14273);
or UO_27 (O_27,N_13273,N_12474);
or UO_28 (O_28,N_13269,N_12044);
or UO_29 (O_29,N_12071,N_12180);
and UO_30 (O_30,N_12096,N_10722);
nand UO_31 (O_31,N_12571,N_13164);
and UO_32 (O_32,N_14214,N_13808);
nor UO_33 (O_33,N_11222,N_11211);
and UO_34 (O_34,N_12689,N_13554);
xor UO_35 (O_35,N_11683,N_11619);
or UO_36 (O_36,N_11157,N_10201);
nor UO_37 (O_37,N_14669,N_13312);
nand UO_38 (O_38,N_11753,N_14074);
and UO_39 (O_39,N_12681,N_13660);
xor UO_40 (O_40,N_10191,N_14729);
nor UO_41 (O_41,N_12786,N_12570);
nor UO_42 (O_42,N_11848,N_12258);
or UO_43 (O_43,N_11327,N_14028);
or UO_44 (O_44,N_10944,N_11053);
nor UO_45 (O_45,N_13570,N_11981);
xor UO_46 (O_46,N_12482,N_12741);
or UO_47 (O_47,N_11174,N_11465);
nand UO_48 (O_48,N_14218,N_12194);
or UO_49 (O_49,N_14087,N_13748);
or UO_50 (O_50,N_12680,N_12790);
nor UO_51 (O_51,N_14489,N_10701);
and UO_52 (O_52,N_10276,N_11705);
or UO_53 (O_53,N_11778,N_11729);
and UO_54 (O_54,N_10186,N_10432);
nand UO_55 (O_55,N_11226,N_12218);
and UO_56 (O_56,N_14385,N_13036);
nor UO_57 (O_57,N_10427,N_14915);
xor UO_58 (O_58,N_11014,N_11641);
xnor UO_59 (O_59,N_12127,N_10766);
xor UO_60 (O_60,N_14504,N_12199);
and UO_61 (O_61,N_14001,N_10199);
nand UO_62 (O_62,N_11032,N_14072);
nand UO_63 (O_63,N_10688,N_13536);
or UO_64 (O_64,N_13756,N_13484);
nor UO_65 (O_65,N_12022,N_12300);
nand UO_66 (O_66,N_12820,N_10095);
nor UO_67 (O_67,N_14270,N_13120);
nor UO_68 (O_68,N_13629,N_13735);
and UO_69 (O_69,N_13278,N_13933);
and UO_70 (O_70,N_13754,N_13724);
nor UO_71 (O_71,N_11727,N_14511);
nand UO_72 (O_72,N_10721,N_14726);
nand UO_73 (O_73,N_12424,N_14964);
nor UO_74 (O_74,N_13927,N_14762);
nor UO_75 (O_75,N_10417,N_10763);
or UO_76 (O_76,N_13931,N_13821);
and UO_77 (O_77,N_11350,N_10174);
xor UO_78 (O_78,N_10675,N_12328);
xor UO_79 (O_79,N_12940,N_12533);
or UO_80 (O_80,N_13863,N_11849);
and UO_81 (O_81,N_12014,N_10636);
nor UO_82 (O_82,N_11771,N_13643);
nor UO_83 (O_83,N_11566,N_12417);
or UO_84 (O_84,N_10853,N_14575);
or UO_85 (O_85,N_10937,N_12515);
nor UO_86 (O_86,N_14369,N_14759);
nand UO_87 (O_87,N_12109,N_12283);
nand UO_88 (O_88,N_14421,N_11446);
and UO_89 (O_89,N_11628,N_11224);
and UO_90 (O_90,N_14121,N_13326);
nor UO_91 (O_91,N_11120,N_12379);
or UO_92 (O_92,N_13242,N_11766);
and UO_93 (O_93,N_12523,N_13609);
xor UO_94 (O_94,N_12364,N_14226);
nand UO_95 (O_95,N_12384,N_10153);
nor UO_96 (O_96,N_11976,N_12753);
nor UO_97 (O_97,N_10181,N_12341);
nor UO_98 (O_98,N_11671,N_11349);
nor UO_99 (O_99,N_14512,N_13227);
and UO_100 (O_100,N_14215,N_13076);
nor UO_101 (O_101,N_13910,N_11166);
and UO_102 (O_102,N_12536,N_13248);
and UO_103 (O_103,N_11360,N_13407);
nand UO_104 (O_104,N_14004,N_10112);
and UO_105 (O_105,N_11597,N_13587);
nor UO_106 (O_106,N_14325,N_14526);
nand UO_107 (O_107,N_13328,N_12240);
nand UO_108 (O_108,N_13752,N_13982);
nand UO_109 (O_109,N_10274,N_13552);
or UO_110 (O_110,N_14140,N_13625);
and UO_111 (O_111,N_12971,N_13794);
or UO_112 (O_112,N_12373,N_11554);
xor UO_113 (O_113,N_13930,N_13160);
and UO_114 (O_114,N_10617,N_10829);
nor UO_115 (O_115,N_11750,N_13736);
and UO_116 (O_116,N_12177,N_14296);
nand UO_117 (O_117,N_13404,N_14297);
nor UO_118 (O_118,N_12943,N_10660);
nor UO_119 (O_119,N_14918,N_12110);
or UO_120 (O_120,N_11861,N_11912);
nand UO_121 (O_121,N_14225,N_13985);
nand UO_122 (O_122,N_12618,N_14542);
or UO_123 (O_123,N_14606,N_13459);
nand UO_124 (O_124,N_13283,N_12727);
and UO_125 (O_125,N_12716,N_13132);
and UO_126 (O_126,N_12748,N_14491);
nor UO_127 (O_127,N_10791,N_10542);
nand UO_128 (O_128,N_12131,N_11815);
nor UO_129 (O_129,N_14801,N_11290);
nand UO_130 (O_130,N_14707,N_10416);
nand UO_131 (O_131,N_11837,N_11036);
and UO_132 (O_132,N_13241,N_10588);
nand UO_133 (O_133,N_12253,N_11204);
xor UO_134 (O_134,N_11150,N_13934);
nor UO_135 (O_135,N_14375,N_14785);
and UO_136 (O_136,N_14795,N_11225);
nor UO_137 (O_137,N_10391,N_13551);
or UO_138 (O_138,N_11335,N_14673);
or UO_139 (O_139,N_10342,N_11678);
or UO_140 (O_140,N_11408,N_10590);
xnor UO_141 (O_141,N_12732,N_12828);
or UO_142 (O_142,N_12863,N_10407);
or UO_143 (O_143,N_13127,N_12900);
and UO_144 (O_144,N_12150,N_12207);
and UO_145 (O_145,N_14363,N_10692);
nand UO_146 (O_146,N_14557,N_14129);
nor UO_147 (O_147,N_12566,N_11844);
xor UO_148 (O_148,N_14714,N_14591);
or UO_149 (O_149,N_11432,N_13006);
nor UO_150 (O_150,N_10121,N_10892);
or UO_151 (O_151,N_11605,N_11203);
or UO_152 (O_152,N_13712,N_10682);
nor UO_153 (O_153,N_14681,N_11700);
or UO_154 (O_154,N_12170,N_13214);
nor UO_155 (O_155,N_12182,N_13973);
or UO_156 (O_156,N_11832,N_11828);
nand UO_157 (O_157,N_13650,N_11154);
nand UO_158 (O_158,N_13354,N_12204);
nand UO_159 (O_159,N_11199,N_12511);
and UO_160 (O_160,N_12498,N_10240);
and UO_161 (O_161,N_10378,N_11076);
nor UO_162 (O_162,N_10658,N_12643);
or UO_163 (O_163,N_11910,N_14108);
nand UO_164 (O_164,N_13993,N_13038);
nand UO_165 (O_165,N_13568,N_14400);
or UO_166 (O_166,N_13637,N_10699);
nand UO_167 (O_167,N_10200,N_11924);
nor UO_168 (O_168,N_12966,N_13122);
nor UO_169 (O_169,N_11846,N_12298);
or UO_170 (O_170,N_11853,N_14638);
nand UO_171 (O_171,N_10243,N_11739);
nor UO_172 (O_172,N_11717,N_14590);
nor UO_173 (O_173,N_12137,N_10321);
nor UO_174 (O_174,N_13817,N_11546);
nand UO_175 (O_175,N_10235,N_14402);
and UO_176 (O_176,N_14247,N_13003);
and UO_177 (O_177,N_10176,N_10712);
and UO_178 (O_178,N_14329,N_10832);
nand UO_179 (O_179,N_11428,N_11718);
or UO_180 (O_180,N_14328,N_10093);
nand UO_181 (O_181,N_11988,N_11643);
xor UO_182 (O_182,N_12469,N_10324);
and UO_183 (O_183,N_12366,N_11599);
or UO_184 (O_184,N_14688,N_14833);
or UO_185 (O_185,N_14172,N_12147);
and UO_186 (O_186,N_13196,N_14520);
nand UO_187 (O_187,N_11132,N_11669);
and UO_188 (O_188,N_14177,N_12227);
nand UO_189 (O_189,N_10630,N_13085);
and UO_190 (O_190,N_13117,N_12015);
xnor UO_191 (O_191,N_11538,N_12405);
or UO_192 (O_192,N_12836,N_13009);
and UO_193 (O_193,N_14570,N_14268);
and UO_194 (O_194,N_13295,N_11770);
or UO_195 (O_195,N_13473,N_12393);
and UO_196 (O_196,N_10696,N_11136);
nor UO_197 (O_197,N_13381,N_13679);
or UO_198 (O_198,N_14710,N_13088);
or UO_199 (O_199,N_11920,N_10461);
nor UO_200 (O_200,N_12237,N_13593);
or UO_201 (O_201,N_12333,N_10025);
or UO_202 (O_202,N_12020,N_14784);
or UO_203 (O_203,N_14308,N_11959);
nand UO_204 (O_204,N_14317,N_10164);
or UO_205 (O_205,N_14536,N_11441);
and UO_206 (O_206,N_14102,N_10189);
or UO_207 (O_207,N_10469,N_12839);
and UO_208 (O_208,N_10054,N_10884);
xor UO_209 (O_209,N_12981,N_11756);
nor UO_210 (O_210,N_13791,N_13775);
xor UO_211 (O_211,N_14101,N_11351);
nand UO_212 (O_212,N_13298,N_10325);
xnor UO_213 (O_213,N_11625,N_12290);
or UO_214 (O_214,N_12857,N_11536);
nand UO_215 (O_215,N_13800,N_13440);
nand UO_216 (O_216,N_14486,N_10949);
or UO_217 (O_217,N_12687,N_14163);
nand UO_218 (O_218,N_14885,N_12104);
nor UO_219 (O_219,N_13705,N_11201);
and UO_220 (O_220,N_12598,N_13246);
or UO_221 (O_221,N_12270,N_13016);
or UO_222 (O_222,N_13492,N_10552);
or UO_223 (O_223,N_12905,N_11230);
and UO_224 (O_224,N_11042,N_11210);
xor UO_225 (O_225,N_13345,N_10604);
or UO_226 (O_226,N_14272,N_11922);
nand UO_227 (O_227,N_12221,N_11758);
and UO_228 (O_228,N_14462,N_13681);
or UO_229 (O_229,N_11077,N_11421);
nand UO_230 (O_230,N_14517,N_11831);
or UO_231 (O_231,N_14998,N_13600);
xor UO_232 (O_232,N_10083,N_11906);
and UO_233 (O_233,N_11930,N_10206);
or UO_234 (O_234,N_13193,N_14629);
and UO_235 (O_235,N_10908,N_10380);
and UO_236 (O_236,N_14005,N_11659);
nand UO_237 (O_237,N_12963,N_13654);
and UO_238 (O_238,N_10345,N_11262);
and UO_239 (O_239,N_12446,N_10741);
and UO_240 (O_240,N_11790,N_11638);
nor UO_241 (O_241,N_13900,N_14053);
or UO_242 (O_242,N_14126,N_11997);
or UO_243 (O_243,N_11244,N_10700);
or UO_244 (O_244,N_14783,N_12667);
nand UO_245 (O_245,N_11152,N_13682);
nand UO_246 (O_246,N_12370,N_14020);
and UO_247 (O_247,N_11447,N_10942);
nand UO_248 (O_248,N_11374,N_12367);
nor UO_249 (O_249,N_14139,N_13953);
xor UO_250 (O_250,N_11819,N_14967);
nor UO_251 (O_251,N_11962,N_14950);
or UO_252 (O_252,N_14691,N_12359);
and UO_253 (O_253,N_13939,N_11061);
nand UO_254 (O_254,N_12045,N_11975);
and UO_255 (O_255,N_12733,N_13444);
and UO_256 (O_256,N_14025,N_13453);
nand UO_257 (O_257,N_14948,N_14877);
nor UO_258 (O_258,N_14834,N_10671);
or UO_259 (O_259,N_10151,N_14713);
and UO_260 (O_260,N_13481,N_12233);
nand UO_261 (O_261,N_10585,N_13413);
nand UO_262 (O_262,N_12171,N_12747);
or UO_263 (O_263,N_13441,N_10177);
and UO_264 (O_264,N_10953,N_12396);
or UO_265 (O_265,N_13247,N_10845);
and UO_266 (O_266,N_14789,N_11401);
nor UO_267 (O_267,N_12398,N_14709);
or UO_268 (O_268,N_14157,N_12146);
xor UO_269 (O_269,N_12202,N_11562);
and UO_270 (O_270,N_10070,N_10792);
and UO_271 (O_271,N_12785,N_12038);
nor UO_272 (O_272,N_10381,N_10064);
and UO_273 (O_273,N_13222,N_11213);
nand UO_274 (O_274,N_12974,N_11109);
nor UO_275 (O_275,N_13675,N_10724);
nor UO_276 (O_276,N_10410,N_13667);
and UO_277 (O_277,N_12872,N_12156);
xnor UO_278 (O_278,N_11434,N_12457);
and UO_279 (O_279,N_11573,N_11851);
or UO_280 (O_280,N_12535,N_13129);
nor UO_281 (O_281,N_10074,N_14650);
nand UO_282 (O_282,N_12419,N_12580);
or UO_283 (O_283,N_11874,N_14130);
nand UO_284 (O_284,N_14541,N_10735);
nand UO_285 (O_285,N_12627,N_13400);
xnor UO_286 (O_286,N_13813,N_10827);
nor UO_287 (O_287,N_12195,N_13175);
or UO_288 (O_288,N_14427,N_12018);
nand UO_289 (O_289,N_11168,N_14151);
nand UO_290 (O_290,N_14501,N_13566);
nand UO_291 (O_291,N_11913,N_11563);
and UO_292 (O_292,N_11326,N_13251);
nor UO_293 (O_293,N_12501,N_12175);
and UO_294 (O_294,N_12039,N_11747);
and UO_295 (O_295,N_13201,N_14937);
nor UO_296 (O_296,N_11875,N_12059);
and UO_297 (O_297,N_12811,N_12010);
and UO_298 (O_298,N_11696,N_13811);
nand UO_299 (O_299,N_11068,N_13877);
and UO_300 (O_300,N_10184,N_14093);
or UO_301 (O_301,N_12877,N_12174);
or UO_302 (O_302,N_12234,N_14391);
or UO_303 (O_303,N_14131,N_11570);
or UO_304 (O_304,N_14029,N_13915);
nand UO_305 (O_305,N_13659,N_13389);
or UO_306 (O_306,N_13823,N_10613);
nor UO_307 (O_307,N_11453,N_14479);
nand UO_308 (O_308,N_10029,N_13778);
nor UO_309 (O_309,N_10223,N_12115);
nor UO_310 (O_310,N_11888,N_14746);
nand UO_311 (O_311,N_12691,N_11319);
xnor UO_312 (O_312,N_12885,N_13186);
nand UO_313 (O_313,N_12578,N_12738);
nor UO_314 (O_314,N_11508,N_14209);
xor UO_315 (O_315,N_12463,N_13968);
or UO_316 (O_316,N_10799,N_12639);
xnor UO_317 (O_317,N_12389,N_11013);
or UO_318 (O_318,N_14313,N_13083);
and UO_319 (O_319,N_12422,N_12685);
nand UO_320 (O_320,N_12599,N_11794);
or UO_321 (O_321,N_13102,N_12767);
nor UO_322 (O_322,N_11274,N_14412);
nor UO_323 (O_323,N_12899,N_12649);
nor UO_324 (O_324,N_13014,N_12678);
or UO_325 (O_325,N_11496,N_12168);
or UO_326 (O_326,N_11062,N_14892);
and UO_327 (O_327,N_10595,N_14627);
nand UO_328 (O_328,N_11125,N_10089);
and UO_329 (O_329,N_10894,N_10218);
or UO_330 (O_330,N_14070,N_13482);
xnor UO_331 (O_331,N_12470,N_14264);
xor UO_332 (O_332,N_10049,N_10533);
nor UO_333 (O_333,N_11209,N_12061);
or UO_334 (O_334,N_13366,N_12878);
and UO_335 (O_335,N_10042,N_11929);
xor UO_336 (O_336,N_10879,N_14105);
nor UO_337 (O_337,N_10111,N_12778);
and UO_338 (O_338,N_10303,N_11801);
nand UO_339 (O_339,N_10088,N_12140);
or UO_340 (O_340,N_12461,N_13063);
nand UO_341 (O_341,N_10150,N_11364);
nand UO_342 (O_342,N_14815,N_13279);
nor UO_343 (O_343,N_13284,N_11473);
or UO_344 (O_344,N_13046,N_14411);
xnor UO_345 (O_345,N_10652,N_13789);
xor UO_346 (O_346,N_14342,N_14406);
nand UO_347 (O_347,N_14263,N_13433);
and UO_348 (O_348,N_11942,N_14899);
nand UO_349 (O_349,N_11431,N_12453);
xor UO_350 (O_350,N_12997,N_14481);
or UO_351 (O_351,N_13128,N_13673);
or UO_352 (O_352,N_10914,N_14257);
nand UO_353 (O_353,N_13402,N_14869);
and UO_354 (O_354,N_11300,N_14698);
xnor UO_355 (O_355,N_11019,N_12225);
and UO_356 (O_356,N_12998,N_11995);
nand UO_357 (O_357,N_13626,N_13642);
nor UO_358 (O_358,N_11951,N_10057);
nand UO_359 (O_359,N_14128,N_12697);
or UO_360 (O_360,N_12694,N_14267);
and UO_361 (O_361,N_14019,N_10233);
nor UO_362 (O_362,N_11070,N_12534);
nand UO_363 (O_363,N_14534,N_11207);
and UO_364 (O_364,N_14780,N_10073);
and UO_365 (O_365,N_10183,N_10965);
and UO_366 (O_366,N_13337,N_10771);
or UO_367 (O_367,N_11504,N_14751);
xnor UO_368 (O_368,N_11067,N_12274);
nor UO_369 (O_369,N_13344,N_13097);
nor UO_370 (O_370,N_12336,N_13511);
or UO_371 (O_371,N_14805,N_13467);
or UO_372 (O_372,N_13049,N_14572);
and UO_373 (O_373,N_10536,N_10230);
nor UO_374 (O_374,N_13819,N_12852);
nor UO_375 (O_375,N_13253,N_14357);
nand UO_376 (O_376,N_12855,N_14024);
nor UO_377 (O_377,N_12945,N_12079);
or UO_378 (O_378,N_10840,N_14771);
or UO_379 (O_379,N_12583,N_14907);
nand UO_380 (O_380,N_12901,N_10185);
nand UO_381 (O_381,N_10566,N_13176);
nand UO_382 (O_382,N_12325,N_14881);
and UO_383 (O_383,N_13890,N_10897);
xor UO_384 (O_384,N_13445,N_11193);
or UO_385 (O_385,N_14659,N_11020);
and UO_386 (O_386,N_11507,N_12692);
and UO_387 (O_387,N_10528,N_12822);
or UO_388 (O_388,N_13213,N_13207);
nand UO_389 (O_389,N_14050,N_11463);
and UO_390 (O_390,N_11609,N_13320);
nor UO_391 (O_391,N_10104,N_12390);
nand UO_392 (O_392,N_12564,N_12016);
and UO_393 (O_393,N_14419,N_12939);
and UO_394 (O_394,N_13442,N_14772);
or UO_395 (O_395,N_11186,N_12527);
and UO_396 (O_396,N_10197,N_11390);
and UO_397 (O_397,N_10866,N_13498);
nand UO_398 (O_398,N_14678,N_11155);
xnor UO_399 (O_399,N_10021,N_10118);
nand UO_400 (O_400,N_10020,N_12883);
and UO_401 (O_401,N_14721,N_10920);
nor UO_402 (O_402,N_10260,N_14192);
and UO_403 (O_403,N_11572,N_13699);
nor UO_404 (O_404,N_10951,N_13469);
nor UO_405 (O_405,N_14201,N_13762);
nor UO_406 (O_406,N_10117,N_13121);
and UO_407 (O_407,N_10835,N_11212);
nand UO_408 (O_408,N_14240,N_13543);
nand UO_409 (O_409,N_10705,N_10710);
and UO_410 (O_410,N_12540,N_11579);
and UO_411 (O_411,N_14530,N_14345);
nand UO_412 (O_412,N_10108,N_10273);
or UO_413 (O_413,N_11899,N_12669);
nor UO_414 (O_414,N_10368,N_14873);
nor UO_415 (O_415,N_13403,N_14879);
and UO_416 (O_416,N_12604,N_14608);
nand UO_417 (O_417,N_11194,N_14010);
or UO_418 (O_418,N_10437,N_13258);
and UO_419 (O_419,N_14523,N_14125);
or UO_420 (O_420,N_13861,N_12572);
and UO_421 (O_421,N_14528,N_11632);
nor UO_422 (O_422,N_12661,N_12126);
and UO_423 (O_423,N_10603,N_13218);
and UO_424 (O_424,N_14809,N_11118);
xor UO_425 (O_425,N_13056,N_12647);
nor UO_426 (O_426,N_14543,N_11363);
xor UO_427 (O_427,N_12655,N_14495);
and UO_428 (O_428,N_13598,N_12445);
nor UO_429 (O_429,N_13395,N_11901);
or UO_430 (O_430,N_13617,N_11075);
xor UO_431 (O_431,N_12737,N_12295);
xor UO_432 (O_432,N_13100,N_10779);
nor UO_433 (O_433,N_12774,N_10402);
or UO_434 (O_434,N_10062,N_14935);
nand UO_435 (O_435,N_14734,N_11397);
and UO_436 (O_436,N_10995,N_10823);
nand UO_437 (O_437,N_11568,N_14114);
xnor UO_438 (O_438,N_13450,N_12522);
xnor UO_439 (O_439,N_14316,N_10134);
or UO_440 (O_440,N_14231,N_13026);
and UO_441 (O_441,N_13239,N_11862);
or UO_442 (O_442,N_14995,N_11416);
nor UO_443 (O_443,N_13019,N_10389);
xor UO_444 (O_444,N_13562,N_12214);
or UO_445 (O_445,N_10561,N_10475);
and UO_446 (O_446,N_11603,N_12795);
and UO_447 (O_447,N_13886,N_13177);
or UO_448 (O_448,N_14248,N_12965);
and UO_449 (O_449,N_13304,N_12443);
or UO_450 (O_450,N_12832,N_13540);
or UO_451 (O_451,N_14826,N_12635);
and UO_452 (O_452,N_12791,N_11044);
nand UO_453 (O_453,N_13959,N_11514);
xnor UO_454 (O_454,N_10903,N_11492);
and UO_455 (O_455,N_12755,N_12846);
nor UO_456 (O_456,N_13181,N_12141);
nand UO_457 (O_457,N_10606,N_14052);
nand UO_458 (O_458,N_14259,N_11805);
and UO_459 (O_459,N_11820,N_10996);
nand UO_460 (O_460,N_11633,N_13115);
nand UO_461 (O_461,N_12276,N_10399);
and UO_462 (O_462,N_11620,N_12824);
and UO_463 (O_463,N_10238,N_13301);
nor UO_464 (O_464,N_12212,N_12941);
or UO_465 (O_465,N_11802,N_13062);
nand UO_466 (O_466,N_13869,N_14104);
or UO_467 (O_467,N_10030,N_12190);
nand UO_468 (O_468,N_13928,N_11500);
or UO_469 (O_469,N_14037,N_10401);
or UO_470 (O_470,N_13670,N_13452);
xor UO_471 (O_471,N_10553,N_10060);
or UO_472 (O_472,N_13691,N_14884);
and UO_473 (O_473,N_12596,N_14813);
or UO_474 (O_474,N_10154,N_13040);
nand UO_475 (O_475,N_14914,N_11331);
nand UO_476 (O_476,N_13401,N_13348);
and UO_477 (O_477,N_13760,N_10281);
xnor UO_478 (O_478,N_14786,N_12722);
nand UO_479 (O_479,N_12705,N_13647);
nand UO_480 (O_480,N_11153,N_12348);
and UO_481 (O_481,N_11486,N_11163);
nand UO_482 (O_482,N_14444,N_14832);
and UO_483 (O_483,N_14574,N_12056);
nand UO_484 (O_484,N_10305,N_11518);
nand UO_485 (O_485,N_12259,N_12456);
nor UO_486 (O_486,N_13285,N_14360);
xor UO_487 (O_487,N_13096,N_10599);
xnor UO_488 (O_488,N_10750,N_13472);
nor UO_489 (O_489,N_13588,N_14141);
or UO_490 (O_490,N_10616,N_11792);
nor UO_491 (O_491,N_10669,N_11824);
xnor UO_492 (O_492,N_12118,N_11501);
and UO_493 (O_493,N_11050,N_10952);
and UO_494 (O_494,N_11784,N_12271);
xor UO_495 (O_495,N_13583,N_10194);
and UO_496 (O_496,N_11969,N_12884);
or UO_497 (O_497,N_14588,N_14671);
nor UO_498 (O_498,N_13761,N_14212);
nor UO_499 (O_499,N_13112,N_10644);
nor UO_500 (O_500,N_14338,N_10365);
nor UO_501 (O_501,N_10090,N_12082);
nand UO_502 (O_502,N_13464,N_11281);
and UO_503 (O_503,N_14794,N_13657);
nand UO_504 (O_504,N_10301,N_11285);
nor UO_505 (O_505,N_12693,N_14073);
and UO_506 (O_506,N_10472,N_11935);
nor UO_507 (O_507,N_10159,N_12651);
nor UO_508 (O_508,N_10486,N_13135);
and UO_509 (O_509,N_13665,N_13544);
nor UO_510 (O_510,N_12450,N_11393);
or UO_511 (O_511,N_12784,N_12838);
xor UO_512 (O_512,N_12376,N_11631);
or UO_513 (O_513,N_12833,N_14625);
and UO_514 (O_514,N_13359,N_11371);
nand UO_515 (O_515,N_11847,N_13281);
and UO_516 (O_516,N_11245,N_11232);
nor UO_517 (O_517,N_13002,N_12394);
nor UO_518 (O_518,N_14975,N_12413);
xnor UO_519 (O_519,N_13728,N_14535);
nor UO_520 (O_520,N_11022,N_10812);
and UO_521 (O_521,N_11105,N_12876);
and UO_522 (O_522,N_10422,N_13205);
nand UO_523 (O_523,N_13105,N_12781);
nand UO_524 (O_524,N_10678,N_13870);
and UO_525 (O_525,N_11111,N_12011);
and UO_526 (O_526,N_12871,N_10384);
and UO_527 (O_527,N_11046,N_11797);
nor UO_528 (O_528,N_13184,N_11133);
nor UO_529 (O_529,N_14562,N_10205);
and UO_530 (O_530,N_10997,N_12349);
nand UO_531 (O_531,N_13338,N_14558);
nor UO_532 (O_532,N_11923,N_12829);
and UO_533 (O_533,N_14559,N_10795);
nor UO_534 (O_534,N_14470,N_12892);
or UO_535 (O_535,N_10442,N_14033);
or UO_536 (O_536,N_12881,N_12414);
nor UO_537 (O_537,N_10072,N_12510);
nor UO_538 (O_538,N_13828,N_11558);
nand UO_539 (O_539,N_10846,N_10481);
or UO_540 (O_540,N_10822,N_14017);
and UO_541 (O_541,N_10405,N_11978);
nor UO_542 (O_542,N_14705,N_11656);
or UO_543 (O_543,N_13827,N_14333);
or UO_544 (O_544,N_10058,N_12645);
and UO_545 (O_545,N_12497,N_10786);
nor UO_546 (O_546,N_14343,N_11873);
nand UO_547 (O_547,N_11143,N_10430);
nor UO_548 (O_548,N_14755,N_10237);
and UO_549 (O_549,N_11868,N_13524);
nor UO_550 (O_550,N_14494,N_11429);
xnor UO_551 (O_551,N_14990,N_12906);
and UO_552 (O_552,N_10115,N_14368);
xnor UO_553 (O_553,N_14438,N_10283);
nand UO_554 (O_554,N_10693,N_11968);
or UO_555 (O_555,N_14891,N_14509);
xor UO_556 (O_556,N_10703,N_11540);
nor UO_557 (O_557,N_10014,N_12568);
or UO_558 (O_558,N_11535,N_14991);
or UO_559 (O_559,N_11722,N_14525);
and UO_560 (O_560,N_10452,N_12186);
and UO_561 (O_561,N_14931,N_11782);
or UO_562 (O_562,N_12615,N_13169);
nor UO_563 (O_563,N_11925,N_11989);
nand UO_564 (O_564,N_10152,N_12592);
and UO_565 (O_565,N_10719,N_10387);
or UO_566 (O_566,N_13265,N_10105);
nor UO_567 (O_567,N_13964,N_12070);
or UO_568 (O_568,N_10814,N_10813);
nor UO_569 (O_569,N_13872,N_10143);
and UO_570 (O_570,N_13232,N_11016);
xnor UO_571 (O_571,N_13156,N_10412);
nor UO_572 (O_572,N_14763,N_14977);
xnor UO_573 (O_573,N_10131,N_12552);
or UO_574 (O_574,N_12848,N_14448);
and UO_575 (O_575,N_13731,N_12993);
or UO_576 (O_576,N_10984,N_14490);
nand UO_577 (O_577,N_12264,N_13310);
or UO_578 (O_578,N_11481,N_12054);
nor UO_579 (O_579,N_12920,N_11693);
and UO_580 (O_580,N_14655,N_13216);
nand UO_581 (O_581,N_11804,N_13010);
and UO_582 (O_582,N_12211,N_12267);
and UO_583 (O_583,N_12814,N_12287);
and UO_584 (O_584,N_10026,N_10320);
and UO_585 (O_585,N_10262,N_10519);
or UO_586 (O_586,N_14457,N_10992);
and UO_587 (O_587,N_13980,N_13209);
nor UO_588 (O_588,N_10508,N_10061);
nor UO_589 (O_589,N_13475,N_12628);
or UO_590 (O_590,N_13580,N_14009);
nand UO_591 (O_591,N_14704,N_10284);
and UO_592 (O_592,N_11183,N_14577);
or UO_593 (O_593,N_13510,N_14521);
nand UO_594 (O_594,N_13797,N_13614);
nor UO_595 (O_595,N_10936,N_10296);
or UO_596 (O_596,N_14842,N_13393);
nor UO_597 (O_597,N_10683,N_14938);
or UO_598 (O_598,N_14835,N_11099);
nand UO_599 (O_599,N_11840,N_14825);
nor UO_600 (O_600,N_10211,N_13891);
xor UO_601 (O_601,N_14600,N_11459);
nand UO_602 (O_602,N_12129,N_11780);
nor UO_603 (O_603,N_10883,N_10156);
xnor UO_604 (O_604,N_11320,N_10868);
nor UO_605 (O_605,N_13892,N_11505);
or UO_606 (O_606,N_10720,N_10376);
nand UO_607 (O_607,N_11857,N_14202);
nor UO_608 (O_608,N_12757,N_12425);
nor UO_609 (O_609,N_12908,N_13742);
or UO_610 (O_610,N_11776,N_13740);
nand UO_611 (O_611,N_10970,N_11217);
nand UO_612 (O_612,N_11591,N_12380);
and UO_613 (O_613,N_10446,N_13415);
nor UO_614 (O_614,N_11970,N_12381);
and UO_615 (O_615,N_12777,N_14466);
nand UO_616 (O_616,N_11476,N_11682);
and UO_617 (O_617,N_13053,N_11661);
and UO_618 (O_618,N_12034,N_14170);
nor UO_619 (O_619,N_13592,N_10697);
nor UO_620 (O_620,N_13843,N_10040);
nor UO_621 (O_621,N_11614,N_13028);
nor UO_622 (O_622,N_12229,N_10525);
nand UO_623 (O_623,N_14184,N_10594);
and UO_624 (O_624,N_11556,N_12477);
xnor UO_625 (O_625,N_12193,N_10232);
and UO_626 (O_626,N_11716,N_14597);
and UO_627 (O_627,N_13126,N_14876);
nor UO_628 (O_628,N_11324,N_11686);
nor UO_629 (O_629,N_13680,N_11256);
and UO_630 (O_630,N_14724,N_10484);
nand UO_631 (O_631,N_14191,N_12739);
xor UO_632 (O_632,N_12594,N_11093);
xor UO_633 (O_633,N_14337,N_12656);
xnor UO_634 (O_634,N_13233,N_12718);
or UO_635 (O_635,N_11724,N_12342);
or UO_636 (O_636,N_12874,N_11676);
or UO_637 (O_637,N_11420,N_11600);
and UO_638 (O_638,N_13250,N_11991);
and UO_639 (O_639,N_12119,N_13549);
nand UO_640 (O_640,N_11662,N_14295);
and UO_641 (O_641,N_13686,N_13436);
or UO_642 (O_642,N_13483,N_12427);
or UO_643 (O_643,N_12975,N_14144);
and UO_644 (O_644,N_13888,N_14903);
and UO_645 (O_645,N_13074,N_14468);
and UO_646 (O_646,N_10160,N_14428);
nor UO_647 (O_647,N_12024,N_10887);
and UO_648 (O_648,N_12236,N_12520);
and UO_649 (O_649,N_12983,N_10650);
nor UO_650 (O_650,N_11037,N_10207);
or UO_651 (O_651,N_11356,N_14800);
and UO_652 (O_652,N_13229,N_12302);
and UO_653 (O_653,N_13282,N_11394);
xor UO_654 (O_654,N_10267,N_14162);
and UO_655 (O_655,N_12793,N_10520);
nor UO_656 (O_656,N_14963,N_10581);
nor UO_657 (O_657,N_14423,N_12531);
nand UO_658 (O_658,N_14403,N_14136);
nor UO_659 (O_659,N_13148,N_12013);
nor UO_660 (O_660,N_13961,N_11996);
nor UO_661 (O_661,N_14571,N_10038);
xnor UO_662 (O_662,N_10573,N_12640);
or UO_663 (O_663,N_12107,N_11523);
nand UO_664 (O_664,N_12653,N_12033);
nor UO_665 (O_665,N_10044,N_11858);
nand UO_666 (O_666,N_13094,N_11301);
xnor UO_667 (O_667,N_13606,N_14068);
nand UO_668 (O_668,N_11228,N_11798);
nand UO_669 (O_669,N_11474,N_14221);
nand UO_670 (O_670,N_13385,N_12799);
or UO_671 (O_671,N_10809,N_11581);
nand UO_672 (O_672,N_14186,N_11220);
and UO_673 (O_673,N_13143,N_12938);
or UO_674 (O_674,N_10931,N_11261);
nand UO_675 (O_675,N_10247,N_12027);
and UO_676 (O_676,N_11180,N_14962);
nand UO_677 (O_677,N_13256,N_10767);
or UO_678 (O_678,N_13145,N_11078);
nor UO_679 (O_679,N_14651,N_13596);
nand UO_680 (O_680,N_12094,N_13124);
nor UO_681 (O_681,N_13849,N_12666);
xnor UO_682 (O_682,N_13411,N_10986);
nor UO_683 (O_683,N_10745,N_13685);
or UO_684 (O_684,N_14808,N_13648);
and UO_685 (O_685,N_10423,N_13390);
xor UO_686 (O_686,N_11196,N_13683);
nor UO_687 (O_687,N_14863,N_13874);
or UO_688 (O_688,N_12665,N_10085);
or UO_689 (O_689,N_11497,N_10390);
and UO_690 (O_690,N_13198,N_12503);
xnor UO_691 (O_691,N_12437,N_11490);
nor UO_692 (O_692,N_13909,N_10339);
nand UO_693 (O_693,N_14095,N_12148);
nor UO_694 (O_694,N_14348,N_14002);
nand UO_695 (O_695,N_14804,N_14843);
or UO_696 (O_696,N_13702,N_10801);
nand UO_697 (O_697,N_12254,N_11470);
nor UO_698 (O_698,N_13349,N_14547);
and UO_699 (O_699,N_12324,N_10572);
xor UO_700 (O_700,N_11783,N_12198);
nand UO_701 (O_701,N_14431,N_12982);
or UO_702 (O_702,N_12262,N_14513);
or UO_703 (O_703,N_13101,N_14997);
and UO_704 (O_704,N_12291,N_12922);
nand UO_705 (O_705,N_12304,N_11362);
nand UO_706 (O_706,N_12151,N_13287);
or UO_707 (O_707,N_12363,N_13418);
and UO_708 (O_708,N_14817,N_13497);
nor UO_709 (O_709,N_12930,N_12454);
or UO_710 (O_710,N_13512,N_10919);
nand UO_711 (O_711,N_13369,N_10464);
xor UO_712 (O_712,N_10834,N_12978);
nor UO_713 (O_713,N_12375,N_13687);
nor UO_714 (O_714,N_10760,N_12842);
nor UO_715 (O_715,N_10962,N_14702);
nand UO_716 (O_716,N_13770,N_13162);
nand UO_717 (O_717,N_10500,N_14586);
and UO_718 (O_718,N_13638,N_14730);
and UO_719 (O_719,N_14265,N_13845);
nor UO_720 (O_720,N_13912,N_12060);
nor UO_721 (O_721,N_11977,N_11084);
or UO_722 (O_722,N_14051,N_14239);
or UO_723 (O_723,N_11344,N_10001);
and UO_724 (O_724,N_11402,N_12928);
or UO_725 (O_725,N_12752,N_14880);
or UO_726 (O_726,N_14619,N_12936);
and UO_727 (O_727,N_10742,N_10366);
nand UO_728 (O_728,N_10526,N_10713);
nand UO_729 (O_729,N_11626,N_14810);
or UO_730 (O_730,N_13478,N_10583);
nand UO_731 (O_731,N_13197,N_12606);
nand UO_732 (O_732,N_11892,N_13548);
nand UO_733 (O_733,N_10797,N_10438);
or UO_734 (O_734,N_10302,N_12548);
or UO_735 (O_735,N_11905,N_11731);
nand UO_736 (O_736,N_10686,N_13044);
or UO_737 (O_737,N_10811,N_12452);
and UO_738 (O_738,N_12835,N_12117);
xor UO_739 (O_739,N_14372,N_14341);
and UO_740 (O_740,N_11530,N_14420);
nand UO_741 (O_741,N_11707,N_14731);
nor UO_742 (O_742,N_14615,N_14648);
or UO_743 (O_743,N_12305,N_14485);
and UO_744 (O_744,N_12035,N_13272);
or UO_745 (O_745,N_10768,N_13260);
xnor UO_746 (O_746,N_12557,N_12989);
nor UO_747 (O_747,N_14388,N_13509);
and UO_748 (O_748,N_13391,N_10256);
or UO_749 (O_749,N_11485,N_14694);
and UO_750 (O_750,N_13889,N_13815);
nand UO_751 (O_751,N_10097,N_13814);
and UO_752 (O_752,N_10972,N_13779);
nor UO_753 (O_753,N_10878,N_14576);
nor UO_754 (O_754,N_13489,N_11184);
and UO_755 (O_755,N_10035,N_10010);
nor UO_756 (O_756,N_10147,N_11367);
and UO_757 (O_757,N_10102,N_10103);
nor UO_758 (O_758,N_13384,N_14837);
or UO_759 (O_759,N_13895,N_11308);
nor UO_760 (O_760,N_12674,N_12213);
nor UO_761 (O_761,N_10755,N_14340);
nor UO_762 (O_762,N_11006,N_13111);
and UO_763 (O_763,N_13692,N_10698);
nor UO_764 (O_764,N_14471,N_11116);
nand UO_765 (O_765,N_11864,N_10842);
nand UO_766 (O_766,N_12354,N_12708);
nand UO_767 (O_767,N_12958,N_13332);
or UO_768 (O_768,N_10331,N_10297);
and UO_769 (O_769,N_11258,N_11838);
or UO_770 (O_770,N_12844,N_14906);
and UO_771 (O_771,N_10448,N_14015);
xor UO_772 (O_772,N_11963,N_14745);
nor UO_773 (O_773,N_10677,N_14189);
nand UO_774 (O_774,N_11938,N_10790);
nor UO_775 (O_775,N_10824,N_13963);
and UO_776 (O_776,N_13023,N_13624);
or UO_777 (O_777,N_12787,N_11219);
and UO_778 (O_778,N_11456,N_14618);
nand UO_779 (O_779,N_11004,N_13938);
nand UO_780 (O_780,N_11811,N_10728);
nor UO_781 (O_781,N_14007,N_13628);
or UO_782 (O_782,N_12924,N_14459);
nor UO_783 (O_783,N_13106,N_10165);
nand UO_784 (O_784,N_11098,N_13057);
nor UO_785 (O_785,N_12279,N_14416);
nor UO_786 (O_786,N_12217,N_10086);
or UO_787 (O_787,N_14469,N_12575);
xnor UO_788 (O_788,N_10825,N_11665);
or UO_789 (O_789,N_11085,N_14284);
and UO_790 (O_790,N_10732,N_11512);
nor UO_791 (O_791,N_11477,N_13611);
and UO_792 (O_792,N_10420,N_10431);
nand UO_793 (O_793,N_13942,N_10122);
nand UO_794 (O_794,N_10855,N_14851);
nand UO_795 (O_795,N_14549,N_13717);
nor UO_796 (O_796,N_14875,N_12659);
nand UO_797 (O_797,N_12915,N_14038);
and UO_798 (O_798,N_13674,N_13358);
xor UO_799 (O_799,N_12409,N_13954);
or UO_800 (O_800,N_13634,N_12455);
and UO_801 (O_801,N_11482,N_14410);
nand UO_802 (O_802,N_13553,N_13329);
nand UO_803 (O_803,N_14253,N_11613);
xnor UO_804 (O_804,N_10280,N_14208);
nor UO_805 (O_805,N_11982,N_11594);
nor UO_806 (O_806,N_10748,N_12486);
and UO_807 (O_807,N_14982,N_12095);
and UO_808 (O_808,N_11164,N_11928);
or UO_809 (O_809,N_10544,N_14934);
and UO_810 (O_810,N_13972,N_11332);
or UO_811 (O_811,N_11947,N_10538);
nand UO_812 (O_812,N_13480,N_10602);
nor UO_813 (O_813,N_12121,N_14841);
and UO_814 (O_814,N_11328,N_13427);
nand UO_815 (O_815,N_14846,N_12909);
nor UO_816 (O_816,N_13425,N_13847);
and UO_817 (O_817,N_14452,N_14440);
or UO_818 (O_818,N_14195,N_10123);
or UO_819 (O_819,N_11762,N_13695);
and UO_820 (O_820,N_13142,N_14617);
and UO_821 (O_821,N_14079,N_11438);
or UO_822 (O_822,N_10917,N_13990);
and UO_823 (O_823,N_12644,N_12128);
and UO_824 (O_824,N_14656,N_10880);
nor UO_825 (O_825,N_12088,N_12902);
and UO_826 (O_826,N_11971,N_10328);
or UO_827 (O_827,N_14291,N_13590);
and UO_828 (O_828,N_10462,N_11713);
nand UO_829 (O_829,N_14000,N_14628);
nor UO_830 (O_830,N_10990,N_10598);
nor UO_831 (O_831,N_12139,N_14374);
and UO_832 (O_832,N_12030,N_13898);
and UO_833 (O_833,N_13753,N_10261);
nor UO_834 (O_834,N_13677,N_10408);
nand UO_835 (O_835,N_12581,N_10621);
nand UO_836 (O_836,N_11461,N_14390);
nand UO_837 (O_837,N_12192,N_11894);
and UO_838 (O_838,N_12507,N_11484);
nand UO_839 (O_839,N_12356,N_11243);
nand UO_840 (O_840,N_11515,N_10947);
or UO_841 (O_841,N_13557,N_12837);
nand UO_842 (O_842,N_14370,N_14581);
or UO_843 (O_843,N_10190,N_13785);
and UO_844 (O_844,N_14732,N_12352);
xnor UO_845 (O_845,N_13133,N_10173);
nand UO_846 (O_846,N_14276,N_13603);
and UO_847 (O_847,N_14910,N_13346);
or UO_848 (O_848,N_14478,N_11435);
nor UO_849 (O_849,N_14871,N_14080);
nand UO_850 (O_850,N_11513,N_13630);
or UO_851 (O_851,N_13039,N_14505);
or UO_852 (O_852,N_11958,N_12853);
and UO_853 (O_853,N_14301,N_13263);
and UO_854 (O_854,N_11720,N_13706);
nor UO_855 (O_855,N_13131,N_14598);
xnor UO_856 (O_856,N_13621,N_12897);
nand UO_857 (O_857,N_13965,N_11664);
xor UO_858 (O_858,N_11878,N_11531);
nor UO_859 (O_859,N_13726,N_12440);
and UO_860 (O_860,N_14774,N_14039);
nand UO_861 (O_861,N_11681,N_12197);
nand UO_862 (O_862,N_11859,N_11200);
nor UO_863 (O_863,N_14269,N_11941);
nand UO_864 (O_864,N_14078,N_13270);
nand UO_865 (O_865,N_12610,N_12357);
nand UO_866 (O_866,N_14919,N_13392);
and UO_867 (O_867,N_14133,N_10132);
or UO_868 (O_868,N_12475,N_10839);
and UO_869 (O_869,N_14992,N_11649);
or UO_870 (O_870,N_11503,N_11795);
and UO_871 (O_871,N_10856,N_10415);
and UO_872 (O_872,N_10769,N_10439);
xnor UO_873 (O_873,N_11684,N_10291);
nand UO_874 (O_874,N_13179,N_13844);
nor UO_875 (O_875,N_11175,N_10640);
nor UO_876 (O_876,N_11791,N_11081);
or UO_877 (O_877,N_14480,N_10547);
nand UO_878 (O_878,N_12383,N_11897);
nand UO_879 (O_879,N_10645,N_11437);
nand UO_880 (O_880,N_10066,N_12933);
nand UO_881 (O_881,N_14076,N_12889);
xnor UO_882 (O_882,N_14047,N_12990);
xnor UO_883 (O_883,N_10004,N_12249);
nor UO_884 (O_884,N_13901,N_13975);
nand UO_885 (O_885,N_13662,N_14533);
and UO_886 (O_886,N_14048,N_14578);
nand UO_887 (O_887,N_14096,N_14929);
and UO_888 (O_888,N_14298,N_10032);
nor UO_889 (O_889,N_13838,N_10974);
and UO_890 (O_890,N_10290,N_14059);
xor UO_891 (O_891,N_10388,N_12743);
nand UO_892 (O_892,N_14687,N_14958);
or UO_893 (O_893,N_10045,N_11478);
nor UO_894 (O_894,N_12312,N_10632);
or UO_895 (O_895,N_14266,N_13261);
nand UO_896 (O_896,N_14217,N_10137);
xnor UO_897 (O_897,N_11586,N_10398);
or UO_898 (O_898,N_12796,N_12111);
nand UO_899 (O_899,N_12307,N_13107);
and UO_900 (O_900,N_13866,N_14312);
nand UO_901 (O_901,N_11772,N_11112);
nand UO_902 (O_902,N_13316,N_11674);
and UO_903 (O_903,N_10400,N_10482);
nor UO_904 (O_904,N_11691,N_10709);
nor UO_905 (O_905,N_13906,N_11557);
or UO_906 (O_906,N_13958,N_12431);
and UO_907 (O_907,N_12715,N_12979);
xnor UO_908 (O_908,N_13199,N_12744);
nor UO_909 (O_909,N_11198,N_11158);
and UO_910 (O_910,N_11549,N_14632);
nand UO_911 (O_911,N_10157,N_12947);
nor UO_912 (O_912,N_14176,N_13688);
or UO_913 (O_913,N_14213,N_11333);
or UO_914 (O_914,N_11457,N_13394);
and UO_915 (O_915,N_11714,N_13503);
or UO_916 (O_916,N_10907,N_13042);
nand UO_917 (O_917,N_13627,N_12320);
or UO_918 (O_918,N_10571,N_10477);
and UO_919 (O_919,N_12544,N_14647);
and UO_920 (O_920,N_14747,N_10627);
nor UO_921 (O_921,N_11449,N_14309);
or UO_922 (O_922,N_12954,N_10752);
nor UO_923 (O_923,N_12812,N_11823);
nor UO_924 (O_924,N_13725,N_10094);
or UO_925 (O_925,N_11103,N_11652);
and UO_926 (O_926,N_13055,N_13296);
nand UO_927 (O_927,N_10875,N_10651);
nor UO_928 (O_928,N_13771,N_14287);
or UO_929 (O_929,N_13021,N_12091);
nor UO_930 (O_930,N_11966,N_11012);
nor UO_931 (O_931,N_14321,N_10485);
or UO_932 (O_932,N_11064,N_11786);
xor UO_933 (O_933,N_13428,N_12361);
nor UO_934 (O_934,N_10382,N_10579);
nand UO_935 (O_935,N_14961,N_11025);
nand UO_936 (O_936,N_10352,N_11239);
nand UO_937 (O_937,N_11379,N_13388);
or UO_938 (O_938,N_13171,N_14091);
or UO_939 (O_939,N_13504,N_11961);
xnor UO_940 (O_940,N_10424,N_14680);
and UO_941 (O_941,N_10219,N_14754);
or UO_942 (O_942,N_11151,N_13419);
nand UO_943 (O_943,N_11268,N_13945);
or UO_944 (O_944,N_13999,N_13215);
nand UO_945 (O_945,N_13743,N_14787);
or UO_946 (O_946,N_13422,N_13781);
nor UO_947 (O_947,N_10928,N_12711);
nor UO_948 (O_948,N_11761,N_10546);
and UO_949 (O_949,N_10964,N_13676);
and UO_950 (O_950,N_14132,N_13514);
or UO_951 (O_951,N_11825,N_11192);
nor UO_952 (O_952,N_12084,N_14838);
nand UO_953 (O_953,N_10299,N_12779);
nand UO_954 (O_954,N_13608,N_13077);
nand UO_955 (O_955,N_10135,N_10443);
nor UO_956 (O_956,N_13357,N_13182);
nor UO_957 (O_957,N_12771,N_11960);
nand UO_958 (O_958,N_12248,N_13881);
nand UO_959 (O_959,N_11080,N_13073);
nand UO_960 (O_960,N_12764,N_10815);
or UO_961 (O_961,N_11191,N_12273);
and UO_962 (O_962,N_11793,N_13166);
nor UO_963 (O_963,N_12724,N_11908);
nand UO_964 (O_964,N_11162,N_14246);
xnor UO_965 (O_965,N_12102,N_11576);
or UO_966 (O_966,N_12547,N_12289);
and UO_967 (O_967,N_12000,N_10758);
and UO_968 (O_968,N_11399,N_11915);
nand UO_969 (O_969,N_11252,N_14941);
nor UO_970 (O_970,N_12408,N_12006);
nor UO_971 (O_971,N_12232,N_13949);
and UO_972 (O_972,N_13064,N_10053);
and UO_973 (O_973,N_14035,N_14864);
nand UO_974 (O_974,N_14782,N_10478);
or UO_975 (O_975,N_14496,N_10110);
nand UO_976 (O_976,N_13880,N_12601);
or UO_977 (O_977,N_11760,N_13173);
or UO_978 (O_978,N_14181,N_10455);
nor UO_979 (O_979,N_10955,N_12113);
nand UO_980 (O_980,N_13319,N_11233);
nand UO_981 (O_981,N_14966,N_14251);
nand UO_982 (O_982,N_11525,N_11945);
or UO_983 (O_983,N_12907,N_10371);
and UO_984 (O_984,N_14717,N_12481);
nor UO_985 (O_985,N_11265,N_13065);
or UO_986 (O_986,N_10893,N_13694);
and UO_987 (O_987,N_11635,N_10994);
xor UO_988 (O_988,N_10681,N_11933);
nor UO_989 (O_989,N_14026,N_10851);
nand UO_990 (O_990,N_13533,N_13271);
or UO_991 (O_991,N_11043,N_14696);
and UO_992 (O_992,N_10343,N_13139);
nand UO_993 (O_993,N_13977,N_11448);
and UO_994 (O_994,N_11346,N_14364);
and UO_995 (O_995,N_11267,N_14652);
xor UO_996 (O_996,N_13238,N_11389);
nand UO_997 (O_997,N_10783,N_11104);
nand UO_998 (O_998,N_12040,N_12611);
and UO_999 (O_999,N_12554,N_11710);
nand UO_1000 (O_1000,N_10954,N_11368);
and UO_1001 (O_1001,N_12657,N_10216);
and UO_1002 (O_1002,N_13138,N_12934);
or UO_1003 (O_1003,N_13921,N_14757);
or UO_1004 (O_1004,N_10322,N_14446);
nor UO_1005 (O_1005,N_10624,N_12582);
nor UO_1006 (O_1006,N_14224,N_12345);
or UO_1007 (O_1007,N_13496,N_11666);
xnor UO_1008 (O_1008,N_12619,N_10867);
nor UO_1009 (O_1009,N_12891,N_13641);
nor UO_1010 (O_1010,N_14944,N_12215);
and UO_1011 (O_1011,N_11774,N_11114);
or UO_1012 (O_1012,N_13114,N_13334);
and UO_1013 (O_1013,N_11667,N_12031);
nand UO_1014 (O_1014,N_11653,N_13266);
nand UO_1015 (O_1015,N_11886,N_14450);
nand UO_1016 (O_1016,N_13799,N_11826);
nor UO_1017 (O_1017,N_10287,N_10221);
and UO_1018 (O_1018,N_12662,N_12542);
and UO_1019 (O_1019,N_10619,N_14928);
nand UO_1020 (O_1020,N_12823,N_13837);
or UO_1021 (O_1021,N_10545,N_13605);
and UO_1022 (O_1022,N_13075,N_13195);
or UO_1023 (O_1023,N_14620,N_11141);
and UO_1024 (O_1024,N_10307,N_11703);
nand UO_1025 (O_1025,N_13458,N_10171);
nand UO_1026 (O_1026,N_12663,N_11071);
xnor UO_1027 (O_1027,N_10327,N_13067);
and UO_1028 (O_1028,N_12746,N_13439);
nand UO_1029 (O_1029,N_14443,N_13719);
xor UO_1030 (O_1030,N_11146,N_11051);
nor UO_1031 (O_1031,N_14371,N_11596);
and UO_1032 (O_1032,N_10024,N_12050);
nand UO_1033 (O_1033,N_10622,N_10476);
xor UO_1034 (O_1034,N_13520,N_12562);
or UO_1035 (O_1035,N_12154,N_11927);
or UO_1036 (O_1036,N_10531,N_12343);
nand UO_1037 (O_1037,N_13237,N_12310);
nor UO_1038 (O_1038,N_10309,N_13851);
nand UO_1039 (O_1039,N_13421,N_10245);
or UO_1040 (O_1040,N_10496,N_10756);
nor UO_1041 (O_1041,N_11197,N_11867);
xor UO_1042 (O_1042,N_14737,N_14083);
nand UO_1043 (O_1043,N_14684,N_11916);
nand UO_1044 (O_1044,N_13351,N_10099);
or UO_1045 (O_1045,N_11509,N_11773);
and UO_1046 (O_1046,N_14492,N_14324);
nand UO_1047 (O_1047,N_14145,N_12630);
or UO_1048 (O_1048,N_10559,N_13672);
xor UO_1049 (O_1049,N_13830,N_11655);
xnor UO_1050 (O_1050,N_12347,N_13905);
or UO_1051 (O_1051,N_11238,N_13275);
or UO_1052 (O_1052,N_13212,N_14280);
nand UO_1053 (O_1053,N_11964,N_12849);
xnor UO_1054 (O_1054,N_11569,N_11165);
nand UO_1055 (O_1055,N_10254,N_12712);
and UO_1056 (O_1056,N_13741,N_14718);
nor UO_1057 (O_1057,N_13829,N_13610);
or UO_1058 (O_1058,N_14207,N_13228);
xnor UO_1059 (O_1059,N_14556,N_13873);
and UO_1060 (O_1060,N_13922,N_14954);
nor UO_1061 (O_1061,N_11914,N_11499);
or UO_1062 (O_1062,N_14042,N_14616);
nor UO_1063 (O_1063,N_12485,N_14286);
nor UO_1064 (O_1064,N_11442,N_11675);
xor UO_1065 (O_1065,N_10370,N_12001);
nor UO_1066 (O_1066,N_13738,N_14138);
xor UO_1067 (O_1067,N_14315,N_11240);
or UO_1068 (O_1068,N_10796,N_10222);
or UO_1069 (O_1069,N_10557,N_10810);
or UO_1070 (O_1070,N_10098,N_12116);
and UO_1071 (O_1071,N_12123,N_10800);
or UO_1072 (O_1072,N_12851,N_11047);
nand UO_1073 (O_1073,N_13978,N_11100);
xnor UO_1074 (O_1074,N_14852,N_12759);
xor UO_1075 (O_1075,N_13875,N_13764);
nor UO_1076 (O_1076,N_12831,N_10490);
nor UO_1077 (O_1077,N_14583,N_10966);
nor UO_1078 (O_1078,N_12436,N_10973);
and UO_1079 (O_1079,N_14318,N_10596);
nand UO_1080 (O_1080,N_10991,N_13206);
or UO_1081 (O_1081,N_10844,N_14089);
nor UO_1082 (O_1082,N_12493,N_10133);
and UO_1083 (O_1083,N_14609,N_12311);
and UO_1084 (O_1084,N_10252,N_12277);
xnor UO_1085 (O_1085,N_11121,N_13399);
nand UO_1086 (O_1086,N_11502,N_10306);
or UO_1087 (O_1087,N_11816,N_12402);
nand UO_1088 (O_1088,N_11763,N_13678);
and UO_1089 (O_1089,N_14500,N_12783);
and UO_1090 (O_1090,N_10242,N_10600);
nand UO_1091 (O_1091,N_12269,N_14299);
or UO_1092 (O_1092,N_13856,N_14952);
and UO_1093 (O_1093,N_13941,N_13987);
nor UO_1094 (O_1094,N_11690,N_12176);
or UO_1095 (O_1095,N_10360,N_13952);
and UO_1096 (O_1096,N_14260,N_13618);
nand UO_1097 (O_1097,N_13792,N_10830);
and UO_1098 (O_1098,N_11604,N_13589);
and UO_1099 (O_1099,N_13768,N_10653);
or UO_1100 (O_1100,N_11571,N_12051);
or UO_1101 (O_1101,N_13308,N_12887);
nand UO_1102 (O_1102,N_14733,N_11699);
and UO_1103 (O_1103,N_12489,N_11711);
nor UO_1104 (O_1104,N_12286,N_10647);
or UO_1105 (O_1105,N_11169,N_11353);
and UO_1106 (O_1106,N_11471,N_10100);
nand UO_1107 (O_1107,N_14021,N_12532);
nor UO_1108 (O_1108,N_11740,N_10821);
or UO_1109 (O_1109,N_12576,N_13305);
or UO_1110 (O_1110,N_14824,N_14434);
and UO_1111 (O_1111,N_11733,N_12586);
nand UO_1112 (O_1112,N_14996,N_13858);
nor UO_1113 (O_1113,N_14289,N_10694);
nand UO_1114 (O_1114,N_10332,N_13225);
nor UO_1115 (O_1115,N_12528,N_12636);
nor UO_1116 (O_1116,N_14836,N_14773);
and UO_1117 (O_1117,N_12043,N_12391);
nand UO_1118 (O_1118,N_13061,N_11737);
nand UO_1119 (O_1119,N_10357,N_11932);
nor UO_1120 (O_1120,N_14897,N_14766);
and UO_1121 (O_1121,N_10802,N_10672);
and UO_1122 (O_1122,N_13720,N_13236);
nand UO_1123 (O_1123,N_14584,N_14460);
nor UO_1124 (O_1124,N_10817,N_14679);
or UO_1125 (O_1125,N_12120,N_13698);
nor UO_1126 (O_1126,N_11688,N_13550);
nand UO_1127 (O_1127,N_13579,N_12466);
nand UO_1128 (O_1128,N_11584,N_13556);
or UO_1129 (O_1129,N_10764,N_12995);
xnor UO_1130 (O_1130,N_10784,N_11698);
nor UO_1131 (O_1131,N_14933,N_12491);
nor UO_1132 (O_1132,N_12509,N_14335);
nor UO_1133 (O_1133,N_14653,N_12404);
nand UO_1134 (O_1134,N_10084,N_12299);
nand UO_1135 (O_1135,N_12326,N_11391);
nor UO_1136 (O_1136,N_10865,N_14723);
nor UO_1137 (O_1137,N_11973,N_13860);
and UO_1138 (O_1138,N_10580,N_12646);
nand UO_1139 (O_1139,N_14862,N_13137);
nand UO_1140 (O_1140,N_11601,N_14553);
or UO_1141 (O_1141,N_12257,N_10737);
or UO_1142 (O_1142,N_13095,N_11382);
or UO_1143 (O_1143,N_13437,N_10912);
nand UO_1144 (O_1144,N_13146,N_10926);
and UO_1145 (O_1145,N_13163,N_11028);
xor UO_1146 (O_1146,N_12546,N_12898);
or UO_1147 (O_1147,N_13029,N_12967);
nand UO_1148 (O_1148,N_10975,N_12242);
nand UO_1149 (O_1149,N_12494,N_14292);
xnor UO_1150 (O_1150,N_10354,N_14014);
and UO_1151 (O_1151,N_13696,N_12403);
and UO_1152 (O_1152,N_14041,N_12047);
or UO_1153 (O_1153,N_10248,N_13595);
nand UO_1154 (O_1154,N_13937,N_11865);
and UO_1155 (O_1155,N_13318,N_13578);
nand UO_1156 (O_1156,N_13424,N_11339);
nor UO_1157 (O_1157,N_13159,N_11704);
and UO_1158 (O_1158,N_10348,N_10913);
or UO_1159 (O_1159,N_10819,N_14398);
nand UO_1160 (O_1160,N_14088,N_10803);
or UO_1161 (O_1161,N_10397,N_10130);
nor UO_1162 (O_1162,N_11288,N_11822);
and UO_1163 (O_1163,N_12108,N_10459);
and UO_1164 (O_1164,N_13559,N_14861);
nor UO_1165 (O_1165,N_14758,N_14243);
nor UO_1166 (O_1166,N_10516,N_14883);
and UO_1167 (O_1167,N_14119,N_10806);
and UO_1168 (O_1168,N_10861,N_13187);
or UO_1169 (O_1169,N_10548,N_14676);
or UO_1170 (O_1170,N_10114,N_13572);
or UO_1171 (O_1171,N_13616,N_10013);
or UO_1172 (O_1172,N_11008,N_14890);
nand UO_1173 (O_1173,N_11615,N_12210);
and UO_1174 (O_1174,N_14960,N_11248);
nor UO_1175 (O_1175,N_13862,N_14613);
nor UO_1176 (O_1176,N_13645,N_13935);
nor UO_1177 (O_1177,N_12613,N_11522);
nor UO_1178 (O_1178,N_10224,N_10445);
nor UO_1179 (O_1179,N_13986,N_13715);
or UO_1180 (O_1180,N_11721,N_10782);
and UO_1181 (O_1181,N_11956,N_11181);
nor UO_1182 (O_1182,N_10956,N_14927);
nand UO_1183 (O_1183,N_10447,N_13528);
or UO_1184 (O_1184,N_14433,N_13822);
nor UO_1185 (O_1185,N_14339,N_11039);
nor UO_1186 (O_1186,N_11426,N_10967);
nor UO_1187 (O_1187,N_12263,N_11297);
or UO_1188 (O_1188,N_12919,N_10691);
nor UO_1189 (O_1189,N_14200,N_11066);
nor UO_1190 (O_1190,N_10337,N_14985);
nor UO_1191 (O_1191,N_13079,N_13379);
nor UO_1192 (O_1192,N_12886,N_11602);
nor UO_1193 (O_1193,N_13154,N_14404);
or UO_1194 (O_1194,N_11672,N_12092);
and UO_1195 (O_1195,N_10805,N_10031);
nor UO_1196 (O_1196,N_10007,N_14596);
or UO_1197 (O_1197,N_10541,N_10518);
nand UO_1198 (O_1198,N_12350,N_11618);
nor UO_1199 (O_1199,N_14546,N_14106);
and UO_1200 (O_1200,N_10501,N_11126);
or UO_1201 (O_1201,N_10979,N_12654);
nor UO_1202 (O_1202,N_14675,N_12632);
and UO_1203 (O_1203,N_12706,N_13563);
nand UO_1204 (O_1204,N_13362,N_13991);
or UO_1205 (O_1205,N_14334,N_11657);
nor UO_1206 (O_1206,N_13267,N_12369);
and UO_1207 (O_1207,N_14649,N_12714);
or UO_1208 (O_1208,N_10170,N_14858);
and UO_1209 (O_1209,N_11247,N_14814);
nand UO_1210 (O_1210,N_10124,N_13244);
nand UO_1211 (O_1211,N_14164,N_13663);
nor UO_1212 (O_1212,N_10708,N_11469);
nand UO_1213 (O_1213,N_12770,N_11058);
nor UO_1214 (O_1214,N_12399,N_13396);
nand UO_1215 (O_1215,N_14971,N_14633);
nor UO_1216 (O_1216,N_14283,N_14663);
nor UO_1217 (O_1217,N_12003,N_10069);
nor UO_1218 (O_1218,N_14045,N_12937);
xnor UO_1219 (O_1219,N_12076,N_12322);
nor UO_1220 (O_1220,N_12602,N_13835);
nand UO_1221 (O_1221,N_12623,N_12953);
or UO_1222 (O_1222,N_13380,N_13098);
and UO_1223 (O_1223,N_11003,N_13919);
nor UO_1224 (O_1224,N_11537,N_14699);
nand UO_1225 (O_1225,N_10852,N_14587);
nor UO_1226 (O_1226,N_10456,N_11937);
and UO_1227 (O_1227,N_13313,N_12049);
nor UO_1228 (O_1228,N_14503,N_14351);
or UO_1229 (O_1229,N_11303,N_14274);
nor UO_1230 (O_1230,N_14331,N_12278);
nor UO_1231 (O_1231,N_10757,N_12053);
and UO_1232 (O_1232,N_12723,N_10192);
and UO_1233 (O_1233,N_12067,N_14765);
or UO_1234 (O_1234,N_14367,N_11187);
and UO_1235 (O_1235,N_11018,N_12329);
nand UO_1236 (O_1236,N_11065,N_14595);
or UO_1237 (O_1237,N_14564,N_12768);
or UO_1238 (O_1238,N_11419,N_11095);
nand UO_1239 (O_1239,N_13651,N_13853);
nor UO_1240 (O_1240,N_12172,N_12241);
or UO_1241 (O_1241,N_11338,N_13331);
and UO_1242 (O_1242,N_13303,N_11173);
and UO_1243 (O_1243,N_13291,N_10109);
nor UO_1244 (O_1244,N_12448,N_11974);
nand UO_1245 (O_1245,N_10440,N_13547);
or UO_1246 (O_1246,N_11130,N_11170);
or UO_1247 (O_1247,N_14193,N_14507);
and UO_1248 (O_1248,N_13420,N_14467);
or UO_1249 (O_1249,N_12245,N_11876);
and UO_1250 (O_1250,N_11887,N_12415);
and UO_1251 (O_1251,N_14573,N_13537);
and UO_1252 (O_1252,N_13567,N_12530);
nor UO_1253 (O_1253,N_10993,N_13926);
or UO_1254 (O_1254,N_11269,N_12675);
nand UO_1255 (O_1255,N_10804,N_13235);
and UO_1256 (O_1256,N_13531,N_11660);
nand UO_1257 (O_1257,N_11185,N_11548);
or UO_1258 (O_1258,N_10649,N_13335);
and UO_1259 (O_1259,N_10664,N_14848);
nand UO_1260 (O_1260,N_12761,N_13701);
or UO_1261 (O_1261,N_14409,N_10329);
and UO_1262 (O_1262,N_14386,N_12888);
nand UO_1263 (O_1263,N_10275,N_14389);
or UO_1264 (O_1264,N_14821,N_14373);
nand UO_1265 (O_1265,N_10587,N_13024);
nor UO_1266 (O_1266,N_13535,N_14418);
nand UO_1267 (O_1267,N_10612,N_13974);
nor UO_1268 (O_1268,N_10940,N_11292);
and UO_1269 (O_1269,N_12447,N_12495);
nor UO_1270 (O_1270,N_13585,N_12921);
or UO_1271 (O_1271,N_10326,N_12987);
or UO_1272 (O_1272,N_11595,N_12707);
nand UO_1273 (O_1273,N_11949,N_14611);
xnor UO_1274 (O_1274,N_10738,N_13777);
nand UO_1275 (O_1275,N_10695,N_14667);
or UO_1276 (O_1276,N_10540,N_12858);
nand UO_1277 (O_1277,N_11400,N_12609);
nor UO_1278 (O_1278,N_13311,N_13729);
or UO_1279 (O_1279,N_10434,N_13970);
nand UO_1280 (O_1280,N_11216,N_11882);
xor UO_1281 (O_1281,N_11278,N_12124);
nor UO_1282 (O_1282,N_11918,N_13405);
xor UO_1283 (O_1283,N_11765,N_13355);
nand UO_1284 (O_1284,N_12964,N_11409);
xor UO_1285 (O_1285,N_14454,N_10019);
or UO_1286 (O_1286,N_10065,N_14739);
or UO_1287 (O_1287,N_13315,N_12181);
nor UO_1288 (O_1288,N_10080,N_13377);
xor UO_1289 (O_1289,N_13555,N_13226);
nor UO_1290 (O_1290,N_13776,N_14708);
nor UO_1291 (O_1291,N_14100,N_11642);
or UO_1292 (O_1292,N_13723,N_10436);
nand UO_1293 (O_1293,N_13297,N_10946);
nand UO_1294 (O_1294,N_10515,N_11980);
nor UO_1295 (O_1295,N_11145,N_12183);
and UO_1296 (O_1296,N_12224,N_11091);
and UO_1297 (O_1297,N_14336,N_13782);
xnor UO_1298 (O_1298,N_11271,N_10162);
and UO_1299 (O_1299,N_12247,N_12074);
or UO_1300 (O_1300,N_14603,N_13745);
xor UO_1301 (O_1301,N_13155,N_12340);
nand UO_1302 (O_1302,N_11325,N_14711);
xnor UO_1303 (O_1303,N_10716,N_11636);
nor UO_1304 (O_1304,N_12231,N_13904);
nor UO_1305 (O_1305,N_10558,N_10393);
or UO_1306 (O_1306,N_14555,N_12317);
nor UO_1307 (O_1307,N_12395,N_10425);
and UO_1308 (O_1308,N_12519,N_13468);
or UO_1309 (O_1309,N_10146,N_10507);
nor UO_1310 (O_1310,N_14077,N_14098);
nand UO_1311 (O_1311,N_11767,N_13721);
or UO_1312 (O_1312,N_10068,N_11955);
or UO_1313 (O_1313,N_10910,N_13521);
or UO_1314 (O_1314,N_13170,N_11015);
xnor UO_1315 (O_1315,N_12002,N_10589);
nor UO_1316 (O_1316,N_13923,N_11528);
and UO_1317 (O_1317,N_11979,N_10759);
nor UO_1318 (O_1318,N_13294,N_13810);
or UO_1319 (O_1319,N_11296,N_12800);
nand UO_1320 (O_1320,N_14898,N_14911);
nor UO_1321 (O_1321,N_12164,N_12196);
nor UO_1322 (O_1322,N_10517,N_13918);
or UO_1323 (O_1323,N_11952,N_11745);
and UO_1324 (O_1324,N_13507,N_10498);
nor UO_1325 (O_1325,N_13542,N_10597);
nand UO_1326 (O_1326,N_14953,N_10902);
nor UO_1327 (O_1327,N_10998,N_14662);
nor UO_1328 (O_1328,N_12802,N_11236);
nand UO_1329 (O_1329,N_13668,N_10905);
xnor UO_1330 (O_1330,N_12896,N_11315);
xnor UO_1331 (O_1331,N_12293,N_12972);
or UO_1332 (O_1332,N_14252,N_13365);
nand UO_1333 (O_1333,N_10727,N_11757);
and UO_1334 (O_1334,N_12926,N_11992);
and UO_1335 (O_1335,N_11629,N_13426);
nor UO_1336 (O_1336,N_12797,N_11639);
and UO_1337 (O_1337,N_10523,N_10560);
nor UO_1338 (O_1338,N_14769,N_14970);
nand UO_1339 (O_1339,N_11545,N_11658);
nand UO_1340 (O_1340,N_11373,N_10863);
or UO_1341 (O_1341,N_10575,N_11835);
nand UO_1342 (O_1342,N_11383,N_11454);
nand UO_1343 (O_1343,N_10373,N_10334);
and UO_1344 (O_1344,N_13574,N_13809);
and UO_1345 (O_1345,N_11302,N_12923);
and UO_1346 (O_1346,N_12360,N_13084);
and UO_1347 (O_1347,N_14167,N_12538);
xor UO_1348 (O_1348,N_10120,N_12625);
and UO_1349 (O_1349,N_12773,N_11555);
xnor UO_1350 (O_1350,N_10654,N_11418);
nor UO_1351 (O_1351,N_14346,N_14839);
xor UO_1352 (O_1352,N_14188,N_10987);
xnor UO_1353 (O_1353,N_13615,N_14046);
nand UO_1354 (O_1354,N_11723,N_11117);
nand UO_1355 (O_1355,N_13150,N_10961);
nand UO_1356 (O_1356,N_13612,N_13255);
xor UO_1357 (O_1357,N_10733,N_14537);
nor UO_1358 (O_1358,N_10577,N_14356);
nand UO_1359 (O_1359,N_10444,N_12558);
or UO_1360 (O_1360,N_13158,N_10626);
and UO_1361 (O_1361,N_13183,N_13652);
nor UO_1362 (O_1362,N_14670,N_11451);
nand UO_1363 (O_1363,N_13417,N_14569);
and UO_1364 (O_1364,N_11781,N_11939);
nand UO_1365 (O_1365,N_11967,N_14194);
and UO_1366 (O_1366,N_14432,N_14307);
nor UO_1367 (O_1367,N_10203,N_14896);
or UO_1368 (O_1368,N_12251,N_14631);
and UO_1369 (O_1369,N_11171,N_11427);
nand UO_1370 (O_1370,N_10119,N_13012);
and UO_1371 (O_1371,N_13353,N_14027);
nor UO_1372 (O_1372,N_11138,N_10492);
or UO_1373 (O_1373,N_14955,N_14165);
xnor UO_1374 (O_1374,N_13623,N_13224);
nand UO_1375 (O_1375,N_13842,N_13041);
nor UO_1376 (O_1376,N_11587,N_13737);
nand UO_1377 (O_1377,N_12086,N_14262);
nand UO_1378 (O_1378,N_11263,N_14792);
or UO_1379 (O_1379,N_11830,N_12133);
nand UO_1380 (O_1380,N_10253,N_13981);
or UO_1381 (O_1381,N_13410,N_14552);
nor UO_1382 (O_1382,N_11283,N_11161);
and UO_1383 (O_1383,N_11128,N_14439);
nor UO_1384 (O_1384,N_12226,N_14514);
nor UO_1385 (O_1385,N_14199,N_12388);
nand UO_1386 (O_1386,N_13113,N_10314);
or UO_1387 (O_1387,N_12894,N_14261);
nor UO_1388 (O_1388,N_11627,N_11560);
or UO_1389 (O_1389,N_10457,N_13018);
or UO_1390 (O_1390,N_12337,N_10182);
nand UO_1391 (O_1391,N_11789,N_10668);
xnor UO_1392 (O_1392,N_14793,N_13025);
nor UO_1393 (O_1393,N_12944,N_13370);
nand UO_1394 (O_1394,N_13151,N_13635);
or UO_1395 (O_1395,N_12955,N_11341);
and UO_1396 (O_1396,N_10960,N_10319);
and UO_1397 (O_1397,N_11972,N_10101);
and UO_1398 (O_1398,N_13575,N_10743);
nor UO_1399 (O_1399,N_12702,N_13147);
nor UO_1400 (O_1400,N_14330,N_11188);
or UO_1401 (O_1401,N_13099,N_11553);
or UO_1402 (O_1402,N_13457,N_10113);
and UO_1403 (O_1403,N_14529,N_13462);
nand UO_1404 (O_1404,N_10142,N_12929);
and UO_1405 (O_1405,N_14012,N_12228);
nand UO_1406 (O_1406,N_14854,N_12873);
and UO_1407 (O_1407,N_13871,N_10854);
nor UO_1408 (O_1408,N_14912,N_10747);
nor UO_1409 (O_1409,N_14303,N_14081);
and UO_1410 (O_1410,N_14567,N_10925);
or UO_1411 (O_1411,N_12893,N_10139);
or UO_1412 (O_1412,N_14484,N_10924);
nand UO_1413 (O_1413,N_10841,N_13368);
and UO_1414 (O_1414,N_12488,N_14781);
and UO_1415 (O_1415,N_11277,N_11376);
nor UO_1416 (O_1416,N_11190,N_12808);
or UO_1417 (O_1417,N_11384,N_14236);
or UO_1418 (O_1418,N_14032,N_14901);
nand UO_1419 (O_1419,N_13833,N_11948);
and UO_1420 (O_1420,N_10008,N_10629);
nor UO_1421 (O_1421,N_13831,N_13989);
or UO_1422 (O_1422,N_10208,N_12960);
nor UO_1423 (O_1423,N_10266,N_10862);
nand UO_1424 (O_1424,N_12243,N_10145);
nand UO_1425 (O_1425,N_13950,N_10285);
or UO_1426 (O_1426,N_10138,N_11806);
nand UO_1427 (O_1427,N_12912,N_14111);
and UO_1428 (O_1428,N_11855,N_14644);
or UO_1429 (O_1429,N_14493,N_12332);
and UO_1430 (O_1430,N_13449,N_10574);
xor UO_1431 (O_1431,N_10009,N_13565);
and UO_1432 (O_1432,N_12956,N_12867);
xor UO_1433 (O_1433,N_10751,N_12265);
or UO_1434 (O_1434,N_12879,N_10772);
nor UO_1435 (O_1435,N_13324,N_10971);
or UO_1436 (O_1436,N_11206,N_12728);
nor UO_1437 (O_1437,N_12418,N_10214);
nor UO_1438 (O_1438,N_11654,N_10395);
nor UO_1439 (O_1439,N_12303,N_11000);
or UO_1440 (O_1440,N_14322,N_10667);
and UO_1441 (O_1441,N_12250,N_14358);
nor UO_1442 (O_1442,N_13001,N_10957);
or UO_1443 (O_1443,N_13289,N_13321);
or UO_1444 (O_1444,N_13571,N_14893);
nand UO_1445 (O_1445,N_13373,N_10362);
nor UO_1446 (O_1446,N_14926,N_10315);
and UO_1447 (O_1447,N_11074,N_14451);
and UO_1448 (O_1448,N_12840,N_11310);
and UO_1449 (O_1449,N_11282,N_10514);
or UO_1450 (O_1450,N_11083,N_11343);
nor UO_1451 (O_1451,N_12573,N_10411);
and UO_1452 (O_1452,N_10922,N_13947);
nor UO_1453 (O_1453,N_14791,N_10136);
or UO_1454 (O_1454,N_12068,N_13322);
and UO_1455 (O_1455,N_10375,N_13408);
nand UO_1456 (O_1456,N_10317,N_14134);
nor UO_1457 (O_1457,N_13903,N_12994);
and UO_1458 (O_1458,N_14728,N_11358);
or UO_1459 (O_1459,N_11673,N_10615);
and UO_1460 (O_1460,N_14743,N_11779);
and UO_1461 (O_1461,N_14807,N_13576);
xor UO_1462 (O_1462,N_13767,N_10158);
nor UO_1463 (O_1463,N_10831,N_11575);
and UO_1464 (O_1464,N_14968,N_12735);
and UO_1465 (O_1465,N_13846,N_10983);
or UO_1466 (O_1466,N_11034,N_11229);
nor UO_1467 (O_1467,N_14502,N_14233);
or UO_1468 (O_1468,N_12025,N_13818);
nand UO_1469 (O_1469,N_14277,N_11234);
xnor UO_1470 (O_1470,N_13341,N_14222);
nor UO_1471 (O_1471,N_10295,N_13091);
or UO_1472 (O_1472,N_12433,N_14582);
nor UO_1473 (O_1473,N_11495,N_11871);
nor UO_1474 (O_1474,N_10419,N_12007);
or UO_1475 (O_1475,N_11702,N_10453);
and UO_1476 (O_1476,N_11884,N_11775);
nand UO_1477 (O_1477,N_12670,N_14692);
and UO_1478 (O_1478,N_12323,N_10250);
nand UO_1479 (O_1479,N_12673,N_12794);
or UO_1480 (O_1480,N_14161,N_10129);
or UO_1481 (O_1481,N_14579,N_10872);
or UO_1482 (O_1482,N_11564,N_11624);
and UO_1483 (O_1483,N_13573,N_12315);
xor UO_1484 (O_1484,N_12734,N_11023);
nand UO_1485 (O_1485,N_11921,N_14323);
nand UO_1486 (O_1486,N_11359,N_11534);
nand UO_1487 (O_1487,N_10228,N_13352);
nor UO_1488 (O_1488,N_13203,N_11694);
nor UO_1489 (O_1489,N_12073,N_10264);
nor UO_1490 (O_1490,N_14086,N_14872);
nand UO_1491 (O_1491,N_14799,N_11547);
or UO_1492 (O_1492,N_13538,N_10633);
nor UO_1493 (O_1493,N_10340,N_13759);
nor UO_1494 (O_1494,N_12335,N_11377);
nand UO_1495 (O_1495,N_10318,N_12362);
nand UO_1496 (O_1496,N_14630,N_14361);
and UO_1497 (O_1497,N_13259,N_13693);
or UO_1498 (O_1498,N_14319,N_13604);
and UO_1499 (O_1499,N_12191,N_10435);
nor UO_1500 (O_1500,N_13020,N_14085);
xor UO_1501 (O_1501,N_10499,N_11799);
xnor UO_1502 (O_1502,N_13979,N_11987);
and UO_1503 (O_1503,N_11904,N_14857);
nor UO_1504 (O_1504,N_13398,N_12850);
and UO_1505 (O_1505,N_11316,N_11651);
nor UO_1506 (O_1506,N_11423,N_10673);
nor UO_1507 (O_1507,N_10428,N_10506);
or UO_1508 (O_1508,N_14326,N_10107);
and UO_1509 (O_1509,N_10637,N_14986);
nand UO_1510 (O_1510,N_12860,N_10787);
nor UO_1511 (O_1511,N_10620,N_10383);
nor UO_1512 (O_1512,N_10985,N_10933);
nor UO_1513 (O_1513,N_11214,N_14205);
or UO_1514 (O_1514,N_14959,N_11189);
nor UO_1515 (O_1515,N_12641,N_14637);
nor UO_1516 (O_1516,N_14332,N_11680);
or UO_1517 (O_1517,N_12932,N_13855);
and UO_1518 (O_1518,N_11663,N_10717);
nand UO_1519 (O_1519,N_12803,N_11291);
nor UO_1520 (O_1520,N_10175,N_10210);
nand UO_1521 (O_1521,N_12699,N_14819);
nand UO_1522 (O_1522,N_11593,N_14185);
and UO_1523 (O_1523,N_13465,N_13932);
nand UO_1524 (O_1524,N_10789,N_11539);
nor UO_1525 (O_1525,N_12961,N_10168);
xnor UO_1526 (O_1526,N_14822,N_14011);
and UO_1527 (O_1527,N_11129,N_13584);
nand UO_1528 (O_1528,N_12517,N_10258);
nand UO_1529 (O_1529,N_10346,N_14994);
nor UO_1530 (O_1530,N_10539,N_14285);
nand UO_1531 (O_1531,N_11640,N_12854);
nand UO_1532 (O_1532,N_14256,N_12826);
nand UO_1533 (O_1533,N_10704,N_14797);
and UO_1534 (O_1534,N_14055,N_11590);
and UO_1535 (O_1535,N_11458,N_14123);
or UO_1536 (O_1536,N_13653,N_13911);
xnor UO_1537 (O_1537,N_12935,N_12062);
nor UO_1538 (O_1538,N_12019,N_12063);
nor UO_1539 (O_1539,N_14279,N_14271);
and UO_1540 (O_1540,N_14472,N_13649);
and UO_1541 (O_1541,N_14749,N_11366);
nand UO_1542 (O_1542,N_13859,N_10563);
or UO_1543 (O_1543,N_12426,N_12513);
and UO_1544 (O_1544,N_14160,N_11856);
and UO_1545 (O_1545,N_10052,N_14461);
and UO_1546 (O_1546,N_13908,N_14946);
or UO_1547 (O_1547,N_11424,N_12080);
and UO_1548 (O_1548,N_12057,N_12173);
or UO_1549 (O_1549,N_11139,N_10551);
or UO_1550 (O_1550,N_14449,N_12959);
or UO_1551 (O_1551,N_12428,N_13302);
nor UO_1552 (O_1552,N_13217,N_14137);
and UO_1553 (O_1553,N_11182,N_10406);
and UO_1554 (O_1554,N_12847,N_12672);
or UO_1555 (O_1555,N_14258,N_14987);
xnor UO_1556 (O_1556,N_11880,N_11235);
nand UO_1557 (O_1557,N_12970,N_14887);
nand UO_1558 (O_1558,N_14422,N_13240);
or UO_1559 (O_1559,N_10605,N_13646);
nand UO_1560 (O_1560,N_13317,N_11038);
nand UO_1561 (O_1561,N_10948,N_12112);
or UO_1562 (O_1562,N_14593,N_12208);
nand UO_1563 (O_1563,N_11415,N_13801);
nand UO_1564 (O_1564,N_10489,N_13333);
nor UO_1565 (O_1565,N_11430,N_12816);
nand UO_1566 (O_1566,N_11583,N_14701);
or UO_1567 (O_1567,N_13751,N_11818);
xnor UO_1568 (O_1568,N_10833,N_14117);
nor UO_1569 (O_1569,N_12460,N_12875);
and UO_1570 (O_1570,N_10941,N_13807);
nand UO_1571 (O_1571,N_14359,N_13772);
xnor UO_1572 (O_1572,N_12209,N_14853);
nor UO_1573 (O_1573,N_14146,N_11708);
or UO_1574 (O_1574,N_10379,N_10483);
nand UO_1575 (O_1575,N_14886,N_13110);
nor UO_1576 (O_1576,N_12462,N_11223);
nor UO_1577 (O_1577,N_14381,N_12046);
nor UO_1578 (O_1578,N_11054,N_10308);
nand UO_1579 (O_1579,N_13223,N_11370);
nor UO_1580 (O_1580,N_14580,N_13523);
nand UO_1581 (O_1581,N_10012,N_14377);
nor UO_1582 (O_1582,N_10655,N_12321);
and UO_1583 (O_1583,N_12105,N_11748);
or UO_1584 (O_1584,N_14742,N_10220);
nand UO_1585 (O_1585,N_11746,N_14905);
or UO_1586 (O_1586,N_14844,N_13755);
and UO_1587 (O_1587,N_12624,N_13090);
nand UO_1588 (O_1588,N_14043,N_13262);
nand UO_1589 (O_1589,N_12652,N_14700);
xor UO_1590 (O_1590,N_12505,N_11944);
nor UO_1591 (O_1591,N_14090,N_14806);
or UO_1592 (O_1592,N_10976,N_10746);
nand UO_1593 (O_1593,N_14984,N_14847);
xor UO_1594 (O_1594,N_11097,N_10226);
or UO_1595 (O_1595,N_12252,N_13230);
or UO_1596 (O_1596,N_10323,N_11231);
xor UO_1597 (O_1597,N_13168,N_13916);
xnor UO_1598 (O_1598,N_10911,N_12946);
and UO_1599 (O_1599,N_12629,N_14894);
nor UO_1600 (O_1600,N_10511,N_14767);
and UO_1601 (O_1601,N_13432,N_12144);
nor UO_1602 (O_1602,N_14599,N_12660);
nand UO_1603 (O_1603,N_14175,N_12720);
and UO_1604 (O_1604,N_12895,N_11957);
or UO_1605 (O_1605,N_13984,N_11526);
or UO_1606 (O_1606,N_13988,N_13619);
nand UO_1607 (O_1607,N_13971,N_11334);
nor UO_1608 (O_1608,N_13431,N_10369);
nand UO_1609 (O_1609,N_11460,N_11317);
nand UO_1610 (O_1610,N_10684,N_10006);
and UO_1611 (O_1611,N_13078,N_14166);
nand UO_1612 (O_1612,N_11852,N_11289);
or UO_1613 (O_1613,N_11298,N_10491);
and UO_1614 (O_1614,N_14453,N_10470);
nor UO_1615 (O_1615,N_14232,N_12638);
nor UO_1616 (O_1616,N_10349,N_14347);
nand UO_1617 (O_1617,N_13330,N_11810);
and UO_1618 (O_1618,N_14865,N_12205);
nor UO_1619 (O_1619,N_13564,N_13887);
nand UO_1620 (O_1620,N_10958,N_11578);
and UO_1621 (O_1621,N_14384,N_14155);
and UO_1622 (O_1622,N_14683,N_14666);
nor UO_1623 (O_1623,N_10535,N_10562);
nand UO_1624 (O_1624,N_13035,N_10059);
nand UO_1625 (O_1625,N_12134,N_14352);
and UO_1626 (O_1626,N_10988,N_13108);
nand UO_1627 (O_1627,N_10744,N_12430);
or UO_1628 (O_1628,N_11266,N_11072);
nand UO_1629 (O_1629,N_11551,N_10272);
nor UO_1630 (O_1630,N_11800,N_11357);
xnor UO_1631 (O_1631,N_10631,N_11254);
nand UO_1632 (O_1632,N_13599,N_14516);
nor UO_1633 (O_1633,N_14978,N_14828);
or UO_1634 (O_1634,N_14016,N_10310);
nand UO_1635 (O_1635,N_11896,N_12167);
and UO_1636 (O_1636,N_13383,N_12988);
or UO_1637 (O_1637,N_13447,N_11087);
and UO_1638 (O_1638,N_11052,N_12508);
or UO_1639 (O_1639,N_14756,N_11101);
and UO_1640 (O_1640,N_12476,N_12187);
nand UO_1641 (O_1641,N_12543,N_13848);
nand UO_1642 (O_1642,N_12821,N_12704);
or UO_1643 (O_1643,N_12306,N_11751);
xor UO_1644 (O_1644,N_10169,N_14643);
nand UO_1645 (O_1645,N_12758,N_10898);
and UO_1646 (O_1646,N_11902,N_12904);
nand UO_1647 (O_1647,N_11940,N_10043);
or UO_1648 (O_1648,N_13716,N_14441);
and UO_1649 (O_1649,N_12159,N_14640);
or UO_1650 (O_1650,N_10213,N_13594);
nor UO_1651 (O_1651,N_12319,N_14254);
or UO_1652 (O_1652,N_13210,N_12529);
xnor UO_1653 (O_1653,N_14657,N_12355);
or UO_1654 (O_1654,N_14720,N_14725);
xor UO_1655 (O_1655,N_13868,N_12081);
and UO_1656 (O_1656,N_10899,N_10047);
and UO_1657 (O_1657,N_14855,N_10774);
nor UO_1658 (O_1658,N_13423,N_12614);
xnor UO_1659 (O_1659,N_14551,N_13655);
nand UO_1660 (O_1660,N_14143,N_12751);
nand UO_1661 (O_1661,N_10554,N_10316);
xnor UO_1662 (O_1662,N_14238,N_13864);
and UO_1663 (O_1663,N_11787,N_11622);
and UO_1664 (O_1664,N_10225,N_11202);
nand UO_1665 (O_1665,N_10092,N_14174);
nand UO_1666 (O_1666,N_14148,N_14677);
or UO_1667 (O_1667,N_12149,N_12160);
nand UO_1668 (O_1668,N_11903,N_11839);
nand UO_1669 (O_1669,N_13374,N_12696);
or UO_1670 (O_1670,N_11668,N_11069);
and UO_1671 (O_1671,N_10895,N_10359);
nand UO_1672 (O_1672,N_13515,N_14084);
or UO_1673 (O_1673,N_12138,N_12996);
xor UO_1674 (O_1674,N_10204,N_13092);
or UO_1675 (O_1675,N_13951,N_13689);
or UO_1676 (O_1676,N_11712,N_12135);
nor UO_1677 (O_1677,N_10657,N_13069);
or UO_1678 (O_1678,N_10549,N_10711);
nand UO_1679 (O_1679,N_10828,N_11106);
and UO_1680 (O_1680,N_13081,N_14658);
and UO_1681 (O_1681,N_10480,N_11293);
nand UO_1682 (O_1682,N_10509,N_10363);
nor UO_1683 (O_1683,N_14506,N_11715);
nand UO_1684 (O_1684,N_12246,N_10479);
or UO_1685 (O_1685,N_13976,N_13116);
nand UO_1686 (O_1686,N_10055,N_14744);
nor UO_1687 (O_1687,N_12682,N_11645);
and UO_1688 (O_1688,N_13327,N_12165);
nand UO_1689 (O_1689,N_11348,N_14936);
nand UO_1690 (O_1690,N_13517,N_11608);
nor UO_1691 (O_1691,N_10300,N_10289);
nand UO_1692 (O_1692,N_14940,N_12272);
xor UO_1693 (O_1693,N_11403,N_11648);
or UO_1694 (O_1694,N_12504,N_10016);
and UO_1695 (O_1695,N_12977,N_13254);
nor UO_1696 (O_1696,N_11102,N_13640);
or UO_1697 (O_1697,N_12695,N_10543);
xor UO_1698 (O_1698,N_14642,N_12561);
and UO_1699 (O_1699,N_13059,N_13532);
nor UO_1700 (O_1700,N_10471,N_11527);
nor UO_1701 (O_1701,N_14135,N_11821);
nand UO_1702 (O_1702,N_12760,N_14956);
nor UO_1703 (O_1703,N_12512,N_12166);
or UO_1704 (O_1704,N_12861,N_10873);
nand UO_1705 (O_1705,N_11280,N_10959);
nand UO_1706 (O_1706,N_13948,N_14752);
nand UO_1707 (O_1707,N_13243,N_12483);
xnor UO_1708 (O_1708,N_13034,N_12280);
or UO_1709 (O_1709,N_13839,N_11679);
nor UO_1710 (O_1710,N_13995,N_14951);
nor UO_1711 (O_1711,N_14216,N_11392);
and UO_1712 (O_1712,N_13708,N_13832);
nor UO_1713 (O_1713,N_14018,N_13983);
and UO_1714 (O_1714,N_13907,N_14294);
nand UO_1715 (O_1715,N_13031,N_11845);
and UO_1716 (O_1716,N_10188,N_12037);
nand UO_1717 (O_1717,N_11160,N_10037);
nor UO_1718 (O_1718,N_13812,N_12297);
nor UO_1719 (O_1719,N_14006,N_12809);
or UO_1720 (O_1720,N_10643,N_12230);
nor UO_1721 (O_1721,N_14237,N_12472);
and UO_1722 (O_1722,N_10702,N_13430);
and UO_1723 (O_1723,N_10212,N_11817);
or UO_1724 (O_1724,N_10773,N_14245);
and UO_1725 (O_1725,N_10263,N_14602);
nand UO_1726 (O_1726,N_14275,N_10257);
and UO_1727 (O_1727,N_14482,N_11253);
nand UO_1728 (O_1728,N_14895,N_10848);
and UO_1729 (O_1729,N_14607,N_13397);
or UO_1730 (O_1730,N_14860,N_10017);
and UO_1731 (O_1731,N_13477,N_14654);
xor UO_1732 (O_1732,N_13917,N_10679);
nand UO_1733 (O_1733,N_11769,N_14003);
and UO_1734 (O_1734,N_10978,N_14818);
or UO_1735 (O_1735,N_12622,N_14979);
and UO_1736 (O_1736,N_11144,N_13119);
and UO_1737 (O_1737,N_14314,N_11877);
nand UO_1738 (O_1738,N_13929,N_10901);
or UO_1739 (O_1739,N_14685,N_14183);
nor UO_1740 (O_1740,N_13722,N_11866);
or UO_1741 (O_1741,N_11142,N_13867);
nand UO_1742 (O_1742,N_10126,N_12664);
or UO_1743 (O_1743,N_10278,N_10689);
xor UO_1744 (O_1744,N_14519,N_14779);
and UO_1745 (O_1745,N_11082,N_11644);
or UO_1746 (O_1746,N_10251,N_10259);
and UO_1747 (O_1747,N_10623,N_11985);
nand UO_1748 (O_1748,N_11294,N_12500);
nor UO_1749 (O_1749,N_11270,N_14753);
or UO_1750 (O_1750,N_10015,N_11788);
nor UO_1751 (O_1751,N_10607,N_10847);
nor UO_1752 (O_1752,N_11984,N_10078);
or UO_1753 (O_1753,N_13490,N_12465);
nand UO_1754 (O_1754,N_10570,N_13474);
and UO_1755 (O_1755,N_10808,N_14350);
nand UO_1756 (O_1756,N_11148,N_10635);
or UO_1757 (O_1757,N_14976,N_12078);
and UO_1758 (O_1758,N_12841,N_14674);
or UO_1759 (O_1759,N_14230,N_10896);
nor UO_1760 (O_1760,N_12650,N_14798);
nand UO_1761 (O_1761,N_14518,N_11898);
nand UO_1762 (O_1762,N_11241,N_14932);
and UO_1763 (O_1763,N_10468,N_10377);
nand UO_1764 (O_1764,N_13007,N_14693);
nand UO_1765 (O_1765,N_14768,N_11208);
or UO_1766 (O_1766,N_11520,N_10969);
and UO_1767 (O_1767,N_12285,N_13149);
and UO_1768 (O_1768,N_12957,N_14544);
xnor UO_1769 (O_1769,N_10209,N_11611);
nand UO_1770 (O_1770,N_12658,N_12819);
nor UO_1771 (O_1771,N_13414,N_10663);
nand UO_1772 (O_1772,N_11307,N_10077);
and UO_1773 (O_1773,N_11946,N_12524);
and UO_1774 (O_1774,N_14425,N_10890);
nand UO_1775 (O_1775,N_11728,N_14197);
nand UO_1776 (O_1776,N_11719,N_11024);
nand UO_1777 (O_1777,N_10555,N_13446);
nor UO_1778 (O_1778,N_11585,N_13508);
or UO_1779 (O_1779,N_12017,N_11010);
and UO_1780 (O_1780,N_11565,N_11318);
or UO_1781 (O_1781,N_12387,N_10241);
nand UO_1782 (O_1782,N_12189,N_10187);
nand UO_1783 (O_1783,N_13703,N_14531);
xnor UO_1784 (O_1784,N_13470,N_10860);
or UO_1785 (O_1785,N_12179,N_13276);
nor UO_1786 (O_1786,N_13434,N_12444);
or UO_1787 (O_1787,N_13443,N_10144);
nand UO_1788 (O_1788,N_12780,N_13429);
or UO_1789 (O_1789,N_14878,N_12344);
or UO_1790 (O_1790,N_14497,N_12754);
xor UO_1791 (O_1791,N_12973,N_14945);
and UO_1792 (O_1792,N_11040,N_13601);
nand UO_1793 (O_1793,N_14424,N_10943);
nand UO_1794 (O_1794,N_10510,N_13093);
or UO_1795 (O_1795,N_12585,N_12152);
and UO_1796 (O_1796,N_13455,N_10780);
or UO_1797 (O_1797,N_11011,N_10676);
xor UO_1798 (O_1798,N_10355,N_14722);
nor UO_1799 (O_1799,N_12677,N_11953);
and UO_1800 (O_1800,N_10502,N_14250);
nor UO_1801 (O_1801,N_11322,N_10871);
nand UO_1802 (O_1802,N_13913,N_12792);
or UO_1803 (O_1803,N_11994,N_12976);
and UO_1804 (O_1804,N_12726,N_11264);
nand UO_1805 (O_1805,N_10268,N_14062);
nand UO_1806 (O_1806,N_14527,N_11221);
and UO_1807 (O_1807,N_14827,N_14049);
or UO_1808 (O_1808,N_14697,N_10067);
xnor UO_1809 (O_1809,N_12185,N_11701);
and UO_1810 (O_1810,N_14376,N_12587);
or UO_1811 (O_1811,N_11749,N_13476);
nand UO_1812 (O_1812,N_12075,N_14634);
nand UO_1813 (O_1813,N_14770,N_13485);
or UO_1814 (O_1814,N_11730,N_14646);
nand UO_1815 (O_1815,N_13671,N_11450);
or UO_1816 (O_1816,N_12565,N_12178);
nand UO_1817 (O_1817,N_11516,N_13000);
nor UO_1818 (O_1818,N_12294,N_14972);
and UO_1819 (O_1819,N_10793,N_10503);
and UO_1820 (O_1820,N_12309,N_14823);
xor UO_1821 (O_1821,N_11273,N_10537);
and UO_1822 (O_1822,N_12368,N_14305);
xor UO_1823 (O_1823,N_12385,N_13734);
nor UO_1824 (O_1824,N_11284,N_14223);
nand UO_1825 (O_1825,N_13620,N_14203);
and UO_1826 (O_1826,N_14464,N_14196);
nand UO_1827 (O_1827,N_10870,N_11122);
or UO_1828 (O_1828,N_12467,N_14601);
nand UO_1829 (O_1829,N_12145,N_12818);
or UO_1830 (O_1830,N_13486,N_14060);
or UO_1831 (O_1831,N_10271,N_10196);
nand UO_1832 (O_1832,N_11854,N_11580);
and UO_1833 (O_1833,N_13194,N_11026);
nand UO_1834 (O_1834,N_13141,N_12392);
nand UO_1835 (O_1835,N_13416,N_10513);
nand UO_1836 (O_1836,N_11060,N_11306);
and UO_1837 (O_1837,N_14508,N_13920);
nand UO_1838 (O_1838,N_14660,N_12742);
or UO_1839 (O_1839,N_10195,N_14554);
xor UO_1840 (O_1840,N_14829,N_14594);
nor UO_1841 (O_1841,N_13082,N_14859);
or UO_1842 (O_1842,N_12559,N_10488);
or UO_1843 (O_1843,N_14499,N_11732);
or UO_1844 (O_1844,N_14811,N_10450);
and UO_1845 (O_1845,N_12130,N_14344);
or UO_1846 (O_1846,N_11936,N_11738);
or UO_1847 (O_1847,N_11309,N_13220);
or UO_1848 (O_1848,N_12518,N_11242);
nor UO_1849 (O_1849,N_14788,N_14290);
and UO_1850 (O_1850,N_13286,N_12577);
nand UO_1851 (O_1851,N_11907,N_10022);
nor UO_1852 (O_1852,N_12261,N_13518);
nand UO_1853 (O_1853,N_10364,N_14110);
or UO_1854 (O_1854,N_11031,N_14538);
nand UO_1855 (O_1855,N_12825,N_11803);
and UO_1856 (O_1856,N_13529,N_12282);
xnor UO_1857 (O_1857,N_13161,N_11881);
or UO_1858 (O_1858,N_12161,N_14840);
nand UO_1859 (O_1859,N_11361,N_13769);
and UO_1860 (O_1860,N_10467,N_11178);
nand UO_1861 (O_1861,N_12334,N_13435);
and UO_1862 (O_1862,N_10140,N_12066);
nor UO_1863 (O_1863,N_13805,N_14624);
xnor UO_1864 (O_1864,N_14568,N_12591);
nor UO_1865 (O_1865,N_13639,N_14158);
or UO_1866 (O_1866,N_11483,N_10723);
and UO_1867 (O_1867,N_13896,N_13841);
or UO_1868 (O_1868,N_14415,N_13850);
nand UO_1869 (O_1869,N_12008,N_14456);
nand UO_1870 (O_1870,N_10982,N_12012);
and UO_1871 (O_1871,N_14560,N_11119);
nand UO_1872 (O_1872,N_10661,N_14909);
xor UO_1873 (O_1873,N_12725,N_10906);
nand UO_1874 (O_1874,N_12962,N_13749);
and UO_1875 (O_1875,N_14300,N_10521);
xnor UO_1876 (O_1876,N_10236,N_12980);
and UO_1877 (O_1877,N_13746,N_10441);
nand UO_1878 (O_1878,N_11414,N_11891);
or UO_1879 (O_1879,N_10313,N_11742);
nor UO_1880 (O_1880,N_13299,N_13300);
or UO_1881 (O_1881,N_13766,N_12968);
xnor UO_1882 (O_1882,N_13577,N_10286);
nand UO_1883 (O_1883,N_11063,N_12948);
nor UO_1884 (O_1884,N_10418,N_12683);
nor UO_1885 (O_1885,N_13730,N_13249);
nand UO_1886 (O_1886,N_12756,N_11279);
or UO_1887 (O_1887,N_13957,N_12798);
xor UO_1888 (O_1888,N_10350,N_13264);
nand UO_1889 (O_1889,N_14690,N_10642);
nor UO_1890 (O_1890,N_13879,N_13448);
nor UO_1891 (O_1891,N_13707,N_13560);
and UO_1892 (O_1892,N_12365,N_10386);
and UO_1893 (O_1893,N_13306,N_14320);
xnor UO_1894 (O_1894,N_12772,N_11809);
or UO_1895 (O_1895,N_10244,N_11543);
or UO_1896 (O_1896,N_11149,N_13966);
and UO_1897 (O_1897,N_10659,N_14293);
and UO_1898 (O_1898,N_10977,N_14515);
or UO_1899 (O_1899,N_14228,N_14868);
xor UO_1900 (O_1900,N_12407,N_12690);
and UO_1901 (O_1901,N_13709,N_10857);
nand UO_1902 (O_1902,N_14071,N_11455);
xnor UO_1903 (O_1903,N_12005,N_12351);
nor UO_1904 (O_1904,N_14116,N_10076);
xor UO_1905 (O_1905,N_11237,N_11759);
nand UO_1906 (O_1906,N_11697,N_13967);
nor UO_1907 (O_1907,N_11027,N_12136);
nand UO_1908 (O_1908,N_10149,N_13787);
and UO_1909 (O_1909,N_10229,N_11218);
and UO_1910 (O_1910,N_12313,N_11425);
nand UO_1911 (O_1911,N_11215,N_14916);
and UO_1912 (O_1912,N_14635,N_10311);
nor UO_1913 (O_1913,N_10487,N_11544);
nor UO_1914 (O_1914,N_12162,N_11796);
or UO_1915 (O_1915,N_10586,N_12560);
or UO_1916 (O_1916,N_14173,N_11001);
nor UO_1917 (O_1917,N_10935,N_13406);
nand UO_1918 (O_1918,N_14983,N_13956);
or UO_1919 (O_1919,N_12353,N_11412);
nor UO_1920 (O_1920,N_10217,N_12567);
nand UO_1921 (O_1921,N_12789,N_13733);
nor UO_1922 (O_1922,N_10715,N_10056);
nor UO_1923 (O_1923,N_12255,N_12103);
nor UO_1924 (O_1924,N_13342,N_12913);
and UO_1925 (O_1925,N_14387,N_12284);
nor UO_1926 (O_1926,N_12158,N_11365);
and UO_1927 (O_1927,N_14107,N_11227);
xor UO_1928 (O_1928,N_10079,N_11398);
or UO_1929 (O_1929,N_13104,N_11260);
nor UO_1930 (O_1930,N_12807,N_14623);
nor UO_1931 (O_1931,N_13361,N_11610);
xnor UO_1932 (O_1932,N_14115,N_10269);
or UO_1933 (O_1933,N_12400,N_12788);
and UO_1934 (O_1934,N_13180,N_13793);
and UO_1935 (O_1935,N_14522,N_10794);
or UO_1936 (O_1936,N_10859,N_10063);
nor UO_1937 (O_1937,N_13527,N_11506);
nand UO_1938 (O_1938,N_11954,N_11314);
nand UO_1939 (O_1939,N_12065,N_13174);
and UO_1940 (O_1940,N_10749,N_12620);
and UO_1941 (O_1941,N_14405,N_12330);
and UO_1942 (O_1942,N_14150,N_10128);
or UO_1943 (O_1943,N_12089,N_14706);
and UO_1944 (O_1944,N_11056,N_13208);
nor UO_1945 (O_1945,N_10989,N_14830);
and UO_1946 (O_1946,N_13914,N_14790);
xor UO_1947 (O_1947,N_12671,N_10215);
or UO_1948 (O_1948,N_12411,N_13519);
and UO_1949 (O_1949,N_11375,N_13463);
nand UO_1950 (O_1950,N_12026,N_13636);
nor UO_1951 (O_1951,N_11736,N_11589);
nand UO_1952 (O_1952,N_11096,N_13364);
nand UO_1953 (O_1953,N_11147,N_11167);
or UO_1954 (O_1954,N_12200,N_10610);
nand UO_1955 (O_1955,N_11354,N_12382);
or UO_1956 (O_1956,N_11321,N_11582);
or UO_1957 (O_1957,N_10048,N_11588);
nand UO_1958 (O_1958,N_12377,N_12862);
nor UO_1959 (O_1959,N_10473,N_10609);
xnor UO_1960 (O_1960,N_11468,N_11405);
nor UO_1961 (O_1961,N_11035,N_13471);
xnor UO_1962 (O_1962,N_14008,N_11445);
nor UO_1963 (O_1963,N_14458,N_11355);
or UO_1964 (O_1964,N_12617,N_12281);
nor UO_1965 (O_1965,N_13591,N_13700);
nor UO_1966 (O_1966,N_13774,N_14178);
or UO_1967 (O_1967,N_10888,N_10249);
and UO_1968 (O_1968,N_12700,N_13878);
nand UO_1969 (O_1969,N_12521,N_13051);
or UO_1970 (O_1970,N_11413,N_14023);
or UO_1971 (O_1971,N_11092,N_12917);
nor UO_1972 (O_1972,N_11552,N_11108);
nand UO_1973 (O_1973,N_14354,N_14510);
nand UO_1974 (O_1974,N_10816,N_10934);
nor UO_1975 (O_1975,N_12506,N_11983);
xnor UO_1976 (O_1976,N_10358,N_10304);
or UO_1977 (O_1977,N_12386,N_14235);
or UO_1978 (O_1978,N_12776,N_12266);
nor UO_1979 (O_1979,N_13125,N_13293);
nor UO_1980 (O_1980,N_12055,N_13252);
nand UO_1981 (O_1981,N_10000,N_12478);
nor UO_1982 (O_1982,N_13033,N_12442);
and UO_1983 (O_1983,N_12372,N_10950);
xnor UO_1984 (O_1984,N_10265,N_14682);
nor UO_1985 (O_1985,N_12815,N_12169);
nand UO_1986 (O_1986,N_13008,N_12459);
nand UO_1987 (O_1987,N_12331,N_11049);
or UO_1988 (O_1988,N_13387,N_12701);
xnor UO_1989 (O_1989,N_12869,N_12449);
and UO_1990 (O_1990,N_11323,N_13711);
xor UO_1991 (O_1991,N_10433,N_13602);
or UO_1992 (O_1992,N_10889,N_11567);
nand UO_1993 (O_1993,N_14153,N_12087);
nor UO_1994 (O_1994,N_13152,N_10753);
or UO_1995 (O_1995,N_10161,N_13962);
and UO_1996 (O_1996,N_14408,N_13454);
xnor UO_1997 (O_1997,N_12406,N_10885);
nand UO_1998 (O_1998,N_11045,N_10385);
and UO_1999 (O_1999,N_10625,N_10584);
endmodule