module basic_2000_20000_2500_100_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
nor U0 (N_0,In_1654,In_116);
xor U1 (N_1,In_1063,In_372);
and U2 (N_2,In_484,In_925);
xor U3 (N_3,In_710,In_1016);
nor U4 (N_4,In_232,In_1446);
nand U5 (N_5,In_949,In_1352);
or U6 (N_6,In_1754,In_1583);
nor U7 (N_7,In_1637,In_934);
nand U8 (N_8,In_721,In_1800);
nor U9 (N_9,In_162,In_986);
nand U10 (N_10,In_1031,In_1171);
nand U11 (N_11,In_709,In_1460);
xor U12 (N_12,In_494,In_1557);
nor U13 (N_13,In_1051,In_502);
nand U14 (N_14,In_327,In_1799);
nor U15 (N_15,In_430,In_115);
nand U16 (N_16,In_1407,In_1209);
or U17 (N_17,In_237,In_633);
or U18 (N_18,In_1372,In_577);
nand U19 (N_19,In_888,In_666);
nor U20 (N_20,In_50,In_195);
or U21 (N_21,In_1683,In_747);
nand U22 (N_22,In_617,In_530);
nand U23 (N_23,In_1138,In_632);
xor U24 (N_24,In_91,In_1285);
nand U25 (N_25,In_1392,In_1199);
nand U26 (N_26,In_156,In_875);
xor U27 (N_27,In_388,In_450);
nor U28 (N_28,In_1593,In_319);
xnor U29 (N_29,In_624,In_396);
or U30 (N_30,In_680,In_314);
xor U31 (N_31,In_687,In_762);
nand U32 (N_32,In_256,In_532);
nand U33 (N_33,In_1228,In_1995);
nand U34 (N_34,In_220,In_235);
xnor U35 (N_35,In_1316,In_1625);
or U36 (N_36,In_379,In_1510);
xor U37 (N_37,In_1920,In_773);
nand U38 (N_38,In_198,In_1350);
nand U39 (N_39,In_616,In_917);
xnor U40 (N_40,In_700,In_1850);
and U41 (N_41,In_1572,In_1853);
xnor U42 (N_42,In_161,In_600);
nand U43 (N_43,In_1948,In_144);
xnor U44 (N_44,In_1010,In_950);
xnor U45 (N_45,In_705,In_1685);
and U46 (N_46,In_1284,In_1842);
nand U47 (N_47,In_610,In_1576);
nand U48 (N_48,In_1459,In_1355);
and U49 (N_49,In_1789,In_1487);
and U50 (N_50,In_1207,In_1613);
or U51 (N_51,In_1471,In_1830);
xor U52 (N_52,In_692,In_1709);
xor U53 (N_53,In_879,In_631);
and U54 (N_54,In_273,In_104);
or U55 (N_55,In_127,In_1560);
or U56 (N_56,In_1480,In_734);
xor U57 (N_57,In_1473,In_973);
and U58 (N_58,In_92,In_1766);
and U59 (N_59,In_1634,In_320);
nor U60 (N_60,In_158,In_89);
nor U61 (N_61,In_301,In_318);
and U62 (N_62,In_575,In_258);
nand U63 (N_63,In_1246,In_1542);
xnor U64 (N_64,In_1906,In_1931);
nand U65 (N_65,In_1732,In_1564);
and U66 (N_66,In_339,In_1202);
nor U67 (N_67,In_248,In_1890);
nor U68 (N_68,In_1369,In_1304);
xnor U69 (N_69,In_15,In_583);
nand U70 (N_70,In_1580,In_30);
or U71 (N_71,In_1029,In_839);
or U72 (N_72,In_668,In_41);
nor U73 (N_73,In_1598,In_128);
and U74 (N_74,In_1532,In_1096);
nor U75 (N_75,In_1255,In_1200);
and U76 (N_76,In_1731,In_20);
or U77 (N_77,In_310,In_1933);
or U78 (N_78,In_1729,In_465);
nor U79 (N_79,In_1341,In_1782);
xor U80 (N_80,In_8,In_1054);
xnor U81 (N_81,In_1911,In_880);
or U82 (N_82,In_1693,In_612);
nand U83 (N_83,In_462,In_1896);
nor U84 (N_84,In_1677,In_1043);
nor U85 (N_85,In_19,In_11);
nand U86 (N_86,In_1705,In_179);
or U87 (N_87,In_820,In_1032);
and U88 (N_88,In_1891,In_857);
and U89 (N_89,In_1434,In_253);
and U90 (N_90,In_227,In_814);
nand U91 (N_91,In_935,In_1380);
and U92 (N_92,In_120,In_1433);
and U93 (N_93,In_1702,In_803);
nand U94 (N_94,In_1025,In_1047);
xor U95 (N_95,In_1111,In_619);
and U96 (N_96,In_216,In_1189);
nor U97 (N_97,In_404,In_169);
nor U98 (N_98,In_982,In_654);
and U99 (N_99,In_1816,In_563);
nand U100 (N_100,In_1741,In_259);
nand U101 (N_101,In_675,In_594);
and U102 (N_102,In_1907,In_1104);
and U103 (N_103,In_1805,In_1205);
and U104 (N_104,In_546,In_1413);
and U105 (N_105,In_1971,In_1235);
nand U106 (N_106,In_1902,In_1397);
nor U107 (N_107,In_154,In_1052);
xnor U108 (N_108,In_1555,In_966);
xnor U109 (N_109,In_365,In_317);
and U110 (N_110,In_1354,In_1240);
or U111 (N_111,In_432,In_843);
or U112 (N_112,In_781,In_603);
and U113 (N_113,In_541,In_268);
nand U114 (N_114,In_171,In_1855);
or U115 (N_115,In_1894,In_138);
xor U116 (N_116,In_1497,In_326);
and U117 (N_117,In_1607,In_164);
nor U118 (N_118,In_1900,In_1441);
xnor U119 (N_119,In_27,In_1651);
xnor U120 (N_120,In_946,In_177);
and U121 (N_121,In_1857,In_533);
nand U122 (N_122,In_1156,In_1073);
xnor U123 (N_123,In_1961,In_470);
and U124 (N_124,In_688,In_1280);
xnor U125 (N_125,In_472,In_1938);
nand U126 (N_126,In_664,In_516);
nor U127 (N_127,In_1586,In_886);
nor U128 (N_128,In_608,In_1250);
and U129 (N_129,In_598,In_124);
nor U130 (N_130,In_1603,In_1829);
xor U131 (N_131,In_1681,In_1874);
or U132 (N_132,In_1868,In_1690);
xor U133 (N_133,In_436,In_1464);
and U134 (N_134,In_1884,In_1626);
xnor U135 (N_135,In_140,In_345);
xnor U136 (N_136,In_1468,In_1516);
nand U137 (N_137,In_485,In_410);
nand U138 (N_138,In_990,In_322);
xnor U139 (N_139,In_1489,In_1062);
nor U140 (N_140,In_1882,In_1181);
or U141 (N_141,In_419,In_1108);
nor U142 (N_142,In_125,In_627);
and U143 (N_143,In_393,In_553);
nand U144 (N_144,In_733,In_1292);
nand U145 (N_145,In_1180,In_76);
or U146 (N_146,In_228,In_1960);
nor U147 (N_147,In_330,In_1554);
xnor U148 (N_148,In_95,In_921);
xor U149 (N_149,In_1405,In_751);
nor U150 (N_150,In_337,In_163);
nor U151 (N_151,In_400,In_887);
nand U152 (N_152,In_1973,In_291);
nor U153 (N_153,In_1442,In_257);
or U154 (N_154,In_959,In_1887);
nand U155 (N_155,In_1262,In_55);
nor U156 (N_156,In_752,In_830);
or U157 (N_157,In_543,In_1779);
and U158 (N_158,In_1954,In_778);
and U159 (N_159,In_685,In_1035);
xnor U160 (N_160,In_867,In_1217);
nor U161 (N_161,In_1194,In_299);
or U162 (N_162,In_1265,In_359);
or U163 (N_163,In_791,In_962);
and U164 (N_164,In_1084,In_1358);
or U165 (N_165,In_335,In_1317);
or U166 (N_166,In_1764,In_518);
nand U167 (N_167,In_1475,In_1076);
xor U168 (N_168,In_449,In_1221);
or U169 (N_169,In_1389,In_423);
xor U170 (N_170,In_1849,In_565);
nand U171 (N_171,In_1937,In_1037);
or U172 (N_172,In_1421,In_1402);
xnor U173 (N_173,In_1122,In_1154);
nand U174 (N_174,In_1708,In_1295);
xnor U175 (N_175,In_1655,In_1865);
nor U176 (N_176,In_996,In_1);
and U177 (N_177,In_838,In_1190);
and U178 (N_178,In_1206,In_1747);
nand U179 (N_179,In_1120,In_605);
xnor U180 (N_180,In_1985,In_836);
nand U181 (N_181,In_560,In_333);
xnor U182 (N_182,In_1270,In_1467);
or U183 (N_183,In_409,In_1962);
nor U184 (N_184,In_440,In_295);
and U185 (N_185,In_550,In_1058);
and U186 (N_186,In_913,In_1535);
xor U187 (N_187,In_1912,In_1632);
nand U188 (N_188,In_1130,In_985);
nor U189 (N_189,In_1835,In_902);
xor U190 (N_190,In_1077,In_1325);
or U191 (N_191,In_841,In_1771);
or U192 (N_192,In_1337,In_729);
and U193 (N_193,In_146,In_898);
nor U194 (N_194,In_662,In_606);
xor U195 (N_195,In_1290,In_939);
xnor U196 (N_196,In_191,In_453);
or U197 (N_197,In_1328,In_1211);
or U198 (N_198,In_1780,In_1293);
and U199 (N_199,In_389,In_1831);
and U200 (N_200,In_1386,In_368);
xor U201 (N_201,In_1457,In_35);
nor U202 (N_202,In_1496,In_1377);
xor U203 (N_203,In_1339,In_1932);
xor U204 (N_204,In_626,In_831);
and U205 (N_205,In_813,In_1977);
and U206 (N_206,In_527,In_278);
nand U207 (N_207,In_424,In_170);
nor U208 (N_208,N_171,In_101);
or U209 (N_209,In_1161,In_1485);
nand U210 (N_210,In_945,In_1989);
or U211 (N_211,In_1314,In_1256);
nor U212 (N_212,In_1346,In_306);
or U213 (N_213,In_402,In_1880);
and U214 (N_214,In_890,In_1301);
nor U215 (N_215,In_1231,In_1570);
nand U216 (N_216,In_1752,In_794);
xnor U217 (N_217,In_1746,In_1469);
and U218 (N_218,In_285,In_1042);
nor U219 (N_219,In_715,In_218);
or U220 (N_220,In_923,N_63);
nor U221 (N_221,In_1701,In_539);
and U222 (N_222,In_84,In_1373);
nand U223 (N_223,In_1118,In_1113);
and U224 (N_224,In_1309,In_375);
xnor U225 (N_225,In_599,In_1137);
xnor U226 (N_226,In_239,In_1670);
nand U227 (N_227,In_713,In_1079);
nand U228 (N_228,In_1975,In_1336);
or U229 (N_229,In_566,In_628);
nand U230 (N_230,In_1689,In_1501);
nor U231 (N_231,In_730,In_576);
and U232 (N_232,In_1187,In_1119);
or U233 (N_233,In_1023,In_593);
or U234 (N_234,In_1443,In_829);
or U235 (N_235,In_1768,In_1000);
and U236 (N_236,In_384,In_1125);
and U237 (N_237,In_215,In_1869);
nand U238 (N_238,In_37,In_549);
and U239 (N_239,In_315,In_455);
xor U240 (N_240,In_224,In_325);
or U241 (N_241,In_1198,In_1713);
nor U242 (N_242,In_1578,In_567);
nor U243 (N_243,In_611,In_102);
xnor U244 (N_244,In_815,In_995);
or U245 (N_245,In_821,In_614);
and U246 (N_246,In_1785,In_1984);
nand U247 (N_247,In_772,In_1514);
nor U248 (N_248,In_1784,In_1716);
nor U249 (N_249,In_477,In_444);
or U250 (N_250,In_1772,In_242);
or U251 (N_251,In_1979,In_718);
xor U252 (N_252,In_1676,In_1537);
or U253 (N_253,In_1271,In_60);
xor U254 (N_254,N_174,N_85);
and U255 (N_255,In_1222,In_183);
and U256 (N_256,In_323,In_361);
or U257 (N_257,In_134,In_172);
xnor U258 (N_258,In_1342,N_77);
nand U259 (N_259,In_1184,In_1002);
nor U260 (N_260,N_62,In_1717);
nand U261 (N_261,In_1820,In_765);
xor U262 (N_262,In_1349,In_1046);
or U263 (N_263,In_745,In_1275);
nor U264 (N_264,In_439,In_963);
xnor U265 (N_265,In_1627,In_1186);
nor U266 (N_266,In_1871,In_1993);
nand U267 (N_267,In_701,In_653);
nand U268 (N_268,N_162,In_105);
nor U269 (N_269,In_703,In_1415);
and U270 (N_270,In_87,In_415);
xnor U271 (N_271,In_407,In_1399);
nor U272 (N_272,In_214,In_834);
nand U273 (N_273,N_173,In_690);
and U274 (N_274,N_89,N_72);
xnor U275 (N_275,In_940,In_1671);
xor U276 (N_276,In_428,In_1463);
and U277 (N_277,In_999,In_1300);
nor U278 (N_278,In_1854,In_1233);
or U279 (N_279,N_61,In_647);
or U280 (N_280,In_1305,N_145);
xor U281 (N_281,In_1067,In_1692);
or U282 (N_282,In_1419,In_1218);
or U283 (N_283,N_27,In_133);
nor U284 (N_284,N_57,In_557);
xnor U285 (N_285,In_660,N_166);
nor U286 (N_286,In_1822,In_1263);
nand U287 (N_287,In_579,In_17);
or U288 (N_288,In_1318,In_304);
xnor U289 (N_289,N_81,In_1362);
nand U290 (N_290,In_1287,In_1517);
nor U291 (N_291,In_262,In_504);
nand U292 (N_292,N_65,In_1159);
nor U293 (N_293,N_191,N_20);
nand U294 (N_294,In_243,In_1841);
or U295 (N_295,In_302,In_1996);
xnor U296 (N_296,In_771,N_17);
nor U297 (N_297,In_1893,N_181);
or U298 (N_298,N_122,In_394);
and U299 (N_299,In_726,In_1101);
xor U300 (N_300,In_435,In_802);
or U301 (N_301,In_1174,In_1091);
nand U302 (N_302,In_1432,In_1639);
and U303 (N_303,In_665,In_294);
nand U304 (N_304,In_1718,In_569);
nor U305 (N_305,In_1359,In_1686);
nor U306 (N_306,In_1730,In_1635);
or U307 (N_307,In_1740,In_460);
nor U308 (N_308,In_537,In_1565);
or U309 (N_309,In_1698,In_1134);
or U310 (N_310,N_25,N_121);
nand U311 (N_311,In_872,In_1146);
and U312 (N_312,In_1321,In_1343);
or U313 (N_313,In_1930,In_1494);
xnor U314 (N_314,In_766,In_903);
nor U315 (N_315,In_88,In_1403);
or U316 (N_316,In_1599,In_1060);
nand U317 (N_317,In_1589,In_1112);
or U318 (N_318,In_947,In_641);
nand U319 (N_319,In_1951,N_147);
or U320 (N_320,N_73,In_1585);
and U321 (N_321,In_746,In_46);
nor U322 (N_322,In_1707,In_987);
nand U323 (N_323,In_942,In_1881);
or U324 (N_324,N_1,In_1541);
xnor U325 (N_325,In_1297,In_1162);
xor U326 (N_326,In_707,In_28);
nor U327 (N_327,In_868,In_279);
nand U328 (N_328,In_225,In_1584);
and U329 (N_329,N_139,In_1672);
or U330 (N_330,In_1382,In_817);
nor U331 (N_331,In_66,N_9);
and U332 (N_332,In_346,N_45);
nand U333 (N_333,In_932,In_334);
and U334 (N_334,In_558,In_490);
and U335 (N_335,In_1007,N_52);
xnor U336 (N_336,In_1085,In_205);
nand U337 (N_337,In_674,In_1109);
and U338 (N_338,In_1424,In_1965);
nand U339 (N_339,In_1472,In_274);
or U340 (N_340,In_184,In_1834);
or U341 (N_341,In_1796,In_63);
or U342 (N_342,N_68,In_406);
or U343 (N_343,In_1974,In_1858);
xor U344 (N_344,In_1330,In_130);
or U345 (N_345,In_1640,In_1664);
xor U346 (N_346,In_1748,In_152);
and U347 (N_347,In_336,In_1922);
or U348 (N_348,In_1970,In_1877);
xor U349 (N_349,In_551,In_209);
or U350 (N_350,In_731,In_374);
nor U351 (N_351,In_1567,In_1094);
nand U352 (N_352,In_178,In_39);
and U353 (N_353,In_1745,In_1688);
nand U354 (N_354,In_1963,In_1033);
and U355 (N_355,In_870,In_860);
xor U356 (N_356,In_1916,In_483);
nand U357 (N_357,In_906,In_1624);
or U358 (N_358,In_331,In_1164);
or U359 (N_359,N_14,In_1824);
or U360 (N_360,In_45,In_716);
nor U361 (N_361,In_1553,N_59);
and U362 (N_362,In_842,N_134);
or U363 (N_363,In_1212,In_1294);
nor U364 (N_364,N_197,In_1374);
or U365 (N_365,N_126,In_1600);
nand U366 (N_366,In_1024,In_1506);
nand U367 (N_367,In_623,In_905);
xor U368 (N_368,In_1398,In_1203);
nand U369 (N_369,In_1320,In_764);
nand U370 (N_370,In_637,In_5);
and U371 (N_371,In_1591,In_998);
nand U372 (N_372,In_1955,In_371);
or U373 (N_373,In_307,In_1710);
nand U374 (N_374,In_458,In_850);
and U375 (N_375,In_529,In_260);
and U376 (N_376,In_1158,In_1763);
xnor U377 (N_377,In_618,In_584);
or U378 (N_378,In_1420,In_33);
or U379 (N_379,In_1999,In_649);
and U380 (N_380,In_422,In_952);
and U381 (N_381,In_1451,In_572);
nor U382 (N_382,In_1022,N_107);
nor U383 (N_383,N_152,In_1719);
and U384 (N_384,In_193,In_1038);
nor U385 (N_385,In_1518,In_799);
xor U386 (N_386,In_426,In_1711);
nand U387 (N_387,In_1425,In_1185);
nor U388 (N_388,In_1777,N_185);
nor U389 (N_389,In_282,N_155);
xnor U390 (N_390,In_132,In_1596);
and U391 (N_391,In_1507,In_213);
xnor U392 (N_392,In_1550,In_1310);
xnor U393 (N_393,In_1527,In_1268);
and U394 (N_394,N_186,N_10);
nand U395 (N_395,In_240,In_1141);
nand U396 (N_396,In_1790,N_165);
nor U397 (N_397,In_1412,In_1525);
or U398 (N_398,In_1107,In_630);
nand U399 (N_399,In_1204,In_1662);
and U400 (N_400,In_1252,N_330);
nor U401 (N_401,In_1026,In_265);
nor U402 (N_402,In_702,In_974);
nand U403 (N_403,In_656,In_474);
and U404 (N_404,In_1491,In_1495);
nand U405 (N_405,N_178,In_1592);
or U406 (N_406,N_265,In_862);
nor U407 (N_407,N_199,In_1302);
or U408 (N_408,In_929,In_503);
xnor U409 (N_409,In_1006,N_373);
or U410 (N_410,In_1944,In_1311);
xnor U411 (N_411,In_1045,N_87);
and U412 (N_412,In_412,In_812);
nand U413 (N_413,N_26,In_1099);
nor U414 (N_414,N_15,In_1028);
nor U415 (N_415,In_80,In_420);
nor U416 (N_416,N_378,In_1547);
or U417 (N_417,In_1941,In_896);
nor U418 (N_418,In_809,In_827);
nor U419 (N_419,In_408,In_522);
nand U420 (N_420,N_84,In_943);
and U421 (N_421,In_369,In_1602);
xor U422 (N_422,In_1499,In_689);
xnor U423 (N_423,In_1697,In_1249);
and U424 (N_424,In_810,In_514);
or U425 (N_425,In_1604,In_1208);
or U426 (N_426,N_136,In_230);
xnor U427 (N_427,N_209,In_914);
nand U428 (N_428,N_95,In_431);
xnor U429 (N_429,N_109,In_145);
nand U430 (N_430,In_106,In_413);
xnor U431 (N_431,In_204,In_1658);
nand U432 (N_432,In_381,In_176);
xor U433 (N_433,In_524,In_1981);
nand U434 (N_434,In_1848,In_1148);
and U435 (N_435,In_1540,In_1106);
nor U436 (N_436,N_249,In_1213);
or U437 (N_437,In_936,N_350);
xor U438 (N_438,In_139,In_847);
xnor U439 (N_439,In_884,In_1642);
and U440 (N_440,In_1652,N_393);
nor U441 (N_441,N_398,In_51);
xor U442 (N_442,In_933,In_103);
xnor U443 (N_443,In_1673,In_1360);
nor U444 (N_444,In_182,In_385);
or U445 (N_445,In_679,N_53);
and U446 (N_446,In_779,In_293);
nand U447 (N_447,N_375,N_268);
nand U448 (N_448,N_138,In_1888);
nor U449 (N_449,In_1406,In_1781);
xor U450 (N_450,N_202,N_337);
and U451 (N_451,N_302,In_756);
xnor U452 (N_452,In_891,In_466);
xor U453 (N_453,In_376,In_481);
and U454 (N_454,In_1629,N_200);
nand U455 (N_455,N_341,N_238);
xor U456 (N_456,In_16,In_226);
and U457 (N_457,N_291,In_698);
or U458 (N_458,In_1843,In_964);
xnor U459 (N_459,In_693,N_314);
or U460 (N_460,In_24,In_108);
xor U461 (N_461,In_1605,In_283);
nor U462 (N_462,In_1126,In_750);
xor U463 (N_463,In_1068,N_359);
nor U464 (N_464,In_1562,In_1017);
and U465 (N_465,In_83,In_920);
or U466 (N_466,In_1381,In_1551);
and U467 (N_467,In_1261,N_243);
xnor U468 (N_468,In_1176,N_344);
and U469 (N_469,N_252,In_433);
xnor U470 (N_470,In_796,In_1003);
xor U471 (N_471,N_211,In_1327);
xor U472 (N_472,In_44,In_856);
or U473 (N_473,In_1219,In_1364);
nand U474 (N_474,In_221,In_10);
nand U475 (N_475,N_176,N_153);
or U476 (N_476,N_206,N_311);
or U477 (N_477,In_1744,In_924);
nand U478 (N_478,N_80,In_300);
xor U479 (N_479,In_31,In_1053);
xnor U480 (N_480,In_1066,In_793);
xor U481 (N_481,N_168,In_1075);
and U482 (N_482,N_343,In_960);
xor U483 (N_483,In_1755,In_1899);
nand U484 (N_484,In_1657,In_201);
or U485 (N_485,N_56,In_706);
nand U486 (N_486,In_1721,In_464);
nand U487 (N_487,N_320,In_1623);
nand U488 (N_488,In_927,In_34);
nor U489 (N_489,In_1956,In_1332);
and U490 (N_490,N_24,In_1170);
or U491 (N_491,N_217,In_267);
xor U492 (N_492,In_822,In_1964);
or U493 (N_493,In_1892,In_1823);
and U494 (N_494,N_34,In_673);
nor U495 (N_495,N_90,In_1682);
or U496 (N_496,In_129,In_954);
nor U497 (N_497,In_251,N_288);
xor U498 (N_498,N_362,In_1734);
or U499 (N_499,In_1409,In_732);
xnor U500 (N_500,N_105,N_167);
or U501 (N_501,In_1196,In_919);
nor U502 (N_502,In_364,In_3);
or U503 (N_503,In_536,In_727);
xor U504 (N_504,N_372,In_1175);
nand U505 (N_505,In_1315,In_96);
or U506 (N_506,In_1760,In_1254);
xor U507 (N_507,In_622,In_442);
or U508 (N_508,In_1753,In_1348);
and U509 (N_509,In_521,N_66);
and U510 (N_510,In_1172,In_437);
nand U511 (N_511,N_156,In_677);
or U512 (N_512,In_1408,In_1633);
nor U513 (N_513,In_186,N_111);
nand U514 (N_514,In_1787,In_1643);
xnor U515 (N_515,In_1152,In_1098);
nor U516 (N_516,In_362,In_1861);
nor U517 (N_517,In_1238,In_979);
nor U518 (N_518,In_510,In_271);
nand U519 (N_519,In_795,In_1323);
nor U520 (N_520,In_1917,In_534);
nand U521 (N_521,In_1601,In_1819);
nand U522 (N_522,In_4,In_509);
xnor U523 (N_523,In_378,In_545);
nand U524 (N_524,In_1059,In_1357);
or U525 (N_525,In_427,In_1012);
nor U526 (N_526,In_1462,N_380);
xor U527 (N_527,In_531,In_308);
nor U528 (N_528,N_264,In_784);
xnor U529 (N_529,In_1511,In_1793);
xor U530 (N_530,In_757,N_12);
nor U531 (N_531,In_1548,N_303);
or U532 (N_532,In_249,In_844);
or U533 (N_533,In_387,In_1559);
and U534 (N_534,In_869,In_972);
nand U535 (N_535,In_1935,In_219);
nand U536 (N_536,In_1361,In_1041);
and U537 (N_537,In_1197,In_479);
xor U538 (N_538,N_333,In_587);
nor U539 (N_539,N_371,In_487);
and U540 (N_540,In_661,In_1288);
nor U541 (N_541,In_136,In_1039);
xnor U542 (N_542,In_1724,N_0);
nor U543 (N_543,In_1173,In_1257);
or U544 (N_544,In_493,In_392);
and U545 (N_545,In_1385,N_389);
xnor U546 (N_546,In_446,In_1102);
nand U547 (N_547,In_1436,N_22);
nor U548 (N_548,In_159,In_1815);
xor U549 (N_549,In_1575,In_1864);
nand U550 (N_550,In_40,In_1476);
nor U551 (N_551,In_585,In_292);
or U552 (N_552,In_508,In_601);
nand U553 (N_553,In_672,In_864);
or U554 (N_554,In_1283,In_1505);
and U555 (N_555,In_118,In_1610);
or U556 (N_556,In_1241,N_31);
and U557 (N_557,In_1620,N_263);
nand U558 (N_558,In_1667,In_816);
nand U559 (N_559,In_1757,In_189);
or U560 (N_560,In_1946,In_1048);
nor U561 (N_561,In_1538,In_1492);
nor U562 (N_562,In_861,In_296);
nand U563 (N_563,In_1188,N_237);
nand U564 (N_564,In_429,In_528);
or U565 (N_565,In_753,In_650);
xnor U566 (N_566,In_1395,In_6);
nor U567 (N_567,In_1980,In_32);
nand U568 (N_568,In_1324,N_137);
nor U569 (N_569,N_51,In_748);
nor U570 (N_570,In_1247,In_1998);
and U571 (N_571,In_1286,In_596);
nand U572 (N_572,In_1387,In_754);
nor U573 (N_573,In_356,In_1738);
and U574 (N_574,N_83,In_109);
or U575 (N_575,In_863,N_347);
or U576 (N_576,In_941,In_909);
and U577 (N_577,In_1994,In_1020);
or U578 (N_578,In_491,N_112);
nand U579 (N_579,In_1939,In_1809);
xor U580 (N_580,In_1453,In_61);
nand U581 (N_581,In_1371,In_1437);
or U582 (N_582,In_131,In_699);
xnor U583 (N_583,In_1064,N_127);
and U584 (N_584,In_499,In_1544);
or U585 (N_585,In_775,In_241);
or U586 (N_586,In_849,In_1526);
xor U587 (N_587,In_266,In_1034);
nand U588 (N_588,In_958,N_269);
nor U589 (N_589,In_1226,In_1070);
nand U590 (N_590,In_1736,N_98);
and U591 (N_591,In_1366,In_497);
nor U592 (N_592,In_1840,N_37);
xnor U593 (N_593,In_895,In_681);
xnor U594 (N_594,In_1727,In_1267);
or U595 (N_595,In_648,N_386);
nand U596 (N_596,In_1791,In_1423);
nor U597 (N_597,N_193,N_149);
xnor U598 (N_598,In_1082,N_184);
or U599 (N_599,N_292,N_315);
xnor U600 (N_600,In_1802,In_682);
xor U601 (N_601,In_1619,N_187);
xnor U602 (N_602,In_1110,In_303);
and U603 (N_603,In_383,In_760);
or U604 (N_604,N_286,In_2);
or U605 (N_605,N_148,N_222);
nand U606 (N_606,In_1145,In_1743);
or U607 (N_607,In_930,In_1438);
nand U608 (N_608,In_1021,In_969);
xnor U609 (N_609,In_1873,In_948);
nand U610 (N_610,In_338,N_425);
xnor U611 (N_611,In_615,In_1333);
nand U612 (N_612,In_1934,N_283);
xnor U613 (N_613,In_956,In_1838);
nor U614 (N_614,In_1504,N_348);
xnor U615 (N_615,In_807,In_1050);
nor U616 (N_616,N_64,N_169);
nand U617 (N_617,In_85,N_198);
nor U618 (N_618,N_160,In_312);
xnor U619 (N_619,In_1281,In_840);
and U620 (N_620,In_1100,In_447);
or U621 (N_621,N_374,In_1243);
nor U622 (N_622,In_1244,N_313);
nand U623 (N_623,N_194,In_1879);
or U624 (N_624,In_1090,N_585);
or U625 (N_625,In_202,N_236);
or U626 (N_626,In_562,N_539);
nand U627 (N_627,N_196,In_486);
nor U628 (N_628,In_1832,In_1594);
and U629 (N_629,N_480,In_911);
nor U630 (N_630,In_349,N_5);
and U631 (N_631,In_658,In_1646);
nor U632 (N_632,N_579,In_1103);
xor U633 (N_633,N_13,In_1223);
nand U634 (N_634,N_154,In_1248);
xor U635 (N_635,In_357,N_228);
and U636 (N_636,N_290,N_210);
nand U637 (N_637,N_516,N_407);
xnor U638 (N_638,In_1528,In_1852);
nand U639 (N_639,In_1298,In_1151);
nand U640 (N_640,In_1513,N_207);
or U641 (N_641,In_559,N_491);
and U642 (N_642,In_1139,N_304);
and U643 (N_643,In_1401,In_953);
nand U644 (N_644,In_1160,N_253);
xnor U645 (N_645,In_1149,In_1011);
or U646 (N_646,In_1923,N_401);
or U647 (N_647,In_399,In_157);
or U648 (N_648,In_1872,In_284);
or U649 (N_649,In_403,N_232);
or U650 (N_650,In_1083,In_492);
nand U651 (N_651,In_643,N_47);
and U652 (N_652,N_535,In_75);
xor U653 (N_653,N_245,In_210);
nor U654 (N_654,In_1279,N_358);
nor U655 (N_655,N_266,In_1886);
or U656 (N_656,In_1778,In_498);
or U657 (N_657,N_392,In_469);
and U658 (N_658,In_739,In_967);
xor U659 (N_659,N_44,In_1430);
nand U660 (N_660,N_258,N_454);
or U661 (N_661,In_1679,N_125);
nor U662 (N_662,In_1282,In_425);
and U663 (N_663,N_352,In_607);
and U664 (N_664,N_574,N_301);
xnor U665 (N_665,N_460,N_188);
xor U666 (N_666,In_1237,N_349);
and U667 (N_667,In_873,In_1061);
nor U668 (N_668,In_1303,In_1523);
and U669 (N_669,In_329,In_1615);
and U670 (N_670,In_828,In_401);
nand U671 (N_671,N_30,In_1345);
nor U672 (N_672,In_1253,N_394);
nor U673 (N_673,In_704,In_590);
nor U674 (N_674,In_395,In_341);
or U675 (N_675,In_1929,N_39);
nor U676 (N_676,In_1384,N_470);
or U677 (N_677,N_221,N_270);
nor U678 (N_678,In_652,In_758);
nand U679 (N_679,In_1005,N_458);
xnor U680 (N_680,In_1648,In_725);
and U681 (N_681,N_218,N_327);
or U682 (N_682,In_1363,In_1897);
xnor U683 (N_683,In_1326,In_1936);
or U684 (N_684,N_332,In_275);
and U685 (N_685,In_1704,In_568);
xor U686 (N_686,In_1410,N_143);
xnor U687 (N_687,In_1515,N_369);
and U688 (N_688,In_1566,In_634);
and U689 (N_689,In_1329,In_1622);
nor U690 (N_690,In_366,In_411);
nand U691 (N_691,In_1379,N_23);
or U692 (N_692,In_74,In_1018);
xnor U693 (N_693,In_642,In_1128);
nand U694 (N_694,N_142,N_587);
xor U695 (N_695,N_443,N_205);
nand U696 (N_696,In_1153,N_248);
and U697 (N_697,In_686,In_352);
nand U698 (N_698,In_1694,In_208);
or U699 (N_699,In_854,In_1905);
and U700 (N_700,In_1618,N_317);
nand U701 (N_701,In_1488,In_1123);
xnor U702 (N_702,N_555,In_342);
xnor U703 (N_703,In_53,In_1910);
or U704 (N_704,N_88,In_1470);
and U705 (N_705,In_110,In_26);
xor U706 (N_706,In_1735,In_1774);
nor U707 (N_707,In_1131,In_1631);
and U708 (N_708,In_525,N_319);
nor U709 (N_709,N_54,In_554);
and U710 (N_710,N_489,In_386);
nor U711 (N_711,In_980,N_567);
nand U712 (N_712,In_1650,In_678);
or U713 (N_713,In_826,In_774);
nand U714 (N_714,In_663,In_1168);
or U715 (N_715,In_1983,In_683);
and U716 (N_716,In_1165,In_1019);
xnor U717 (N_717,In_7,N_259);
nor U718 (N_718,In_77,In_1909);
nand U719 (N_719,In_1479,In_473);
nand U720 (N_720,In_1474,N_216);
and U721 (N_721,In_255,In_107);
and U722 (N_722,N_547,In_1836);
xor U723 (N_723,In_1915,N_381);
and U724 (N_724,In_309,In_937);
and U725 (N_725,In_1178,In_1490);
xor U726 (N_726,N_468,In_1478);
nor U727 (N_727,In_165,In_1245);
and U728 (N_728,In_977,In_1621);
and U729 (N_729,In_344,In_1569);
nand U730 (N_730,In_1232,N_465);
xor U731 (N_731,In_1088,In_1444);
nor U732 (N_732,In_897,In_552);
nand U733 (N_733,N_411,In_1536);
nand U734 (N_734,In_1582,In_1508);
nor U735 (N_735,N_306,In_1477);
nor U736 (N_736,In_1455,In_719);
and U737 (N_737,In_370,In_276);
nor U738 (N_738,In_1870,In_931);
nor U739 (N_739,In_160,In_1552);
nor U740 (N_740,In_548,N_33);
xor U741 (N_741,In_69,N_563);
nor U742 (N_742,In_150,In_1057);
nor U743 (N_743,In_65,In_1015);
nor U744 (N_744,In_1638,N_158);
nand U745 (N_745,In_846,In_535);
or U746 (N_746,In_877,In_776);
or U747 (N_747,N_502,In_808);
nor U748 (N_748,N_434,In_1860);
or U749 (N_749,In_507,In_1368);
or U750 (N_750,In_1383,N_8);
nor U751 (N_751,In_1678,In_1684);
xnor U752 (N_752,N_519,In_989);
or U753 (N_753,N_213,In_175);
or U754 (N_754,N_430,N_130);
and U755 (N_755,In_382,In_1210);
and U756 (N_756,In_983,N_472);
xor U757 (N_757,In_777,In_993);
nand U758 (N_758,In_482,N_28);
or U759 (N_759,In_1224,N_231);
xor U760 (N_760,In_561,In_272);
nand U761 (N_761,In_955,N_104);
or U762 (N_762,In_523,N_335);
xnor U763 (N_763,In_1105,In_1659);
and U764 (N_764,In_244,In_667);
and U765 (N_765,N_583,N_7);
xor U766 (N_766,N_588,N_339);
nor U767 (N_767,In_461,N_223);
nor U768 (N_768,N_241,N_382);
or U769 (N_769,In_542,In_625);
and U770 (N_770,In_785,In_1696);
or U771 (N_771,N_580,In_443);
xor U772 (N_772,In_1143,In_111);
or U773 (N_773,In_1695,In_901);
and U774 (N_774,N_408,N_485);
and U775 (N_775,N_564,N_445);
nor U776 (N_776,In_1391,In_1502);
nor U777 (N_777,In_742,In_1273);
xor U778 (N_778,In_1259,N_49);
or U779 (N_779,N_402,N_536);
or U780 (N_780,In_1114,In_651);
nor U781 (N_781,In_866,In_1814);
and U782 (N_782,In_1806,N_599);
or U783 (N_783,N_510,N_477);
nand U784 (N_784,N_505,In_1065);
and U785 (N_785,In_744,In_1133);
nor U786 (N_786,N_42,N_11);
or U787 (N_787,In_112,In_944);
nor U788 (N_788,In_1876,In_78);
or U789 (N_789,N_363,N_474);
nor U790 (N_790,N_385,N_409);
nand U791 (N_791,In_1533,In_1396);
xor U792 (N_792,N_38,In_1878);
nor U793 (N_793,N_325,In_405);
nor U794 (N_794,In_59,N_546);
xnor U795 (N_795,N_183,N_255);
and U796 (N_796,N_551,N_391);
and U797 (N_797,N_541,N_569);
xnor U798 (N_798,In_360,In_367);
and U799 (N_799,In_1454,In_723);
or U800 (N_800,N_520,In_1759);
xnor U801 (N_801,In_289,N_100);
xor U802 (N_802,In_1097,N_761);
nand U803 (N_803,In_1895,In_1561);
nand U804 (N_804,In_380,In_1418);
nor U805 (N_805,In_916,In_1798);
nand U806 (N_806,In_1992,N_626);
or U807 (N_807,In_467,In_1988);
xnor U808 (N_808,N_791,In_1095);
nor U809 (N_809,In_582,In_991);
xnor U810 (N_810,N_779,N_117);
nor U811 (N_811,In_119,In_1908);
nor U812 (N_812,In_1086,In_254);
xor U813 (N_813,In_250,In_173);
or U814 (N_814,In_735,N_189);
nor U815 (N_815,In_1191,In_229);
nand U816 (N_816,N_2,N_414);
or U817 (N_817,N_782,In_1866);
xor U818 (N_818,In_1997,In_1390);
or U819 (N_819,N_351,N_298);
nor U820 (N_820,N_689,In_305);
nand U821 (N_821,N_4,In_783);
and U822 (N_822,In_1539,In_1597);
xnor U823 (N_823,In_1239,In_853);
xnor U824 (N_824,In_43,In_574);
xor U825 (N_825,In_855,In_1797);
nand U826 (N_826,In_513,In_22);
and U827 (N_827,In_155,In_231);
and U828 (N_828,N_608,N_702);
and U829 (N_829,N_778,In_199);
or U830 (N_830,N_478,In_899);
nor U831 (N_831,In_604,In_1767);
and U832 (N_832,In_1335,In_1666);
or U833 (N_833,N_496,N_598);
or U834 (N_834,In_117,N_312);
nor U835 (N_835,N_771,In_277);
nor U836 (N_836,In_573,In_1786);
and U837 (N_837,In_313,In_1773);
nand U838 (N_838,N_552,In_1440);
or U839 (N_839,In_644,N_638);
and U840 (N_840,In_501,N_735);
and U841 (N_841,In_1251,N_715);
and U842 (N_842,In_1577,In_72);
and U843 (N_843,In_1959,In_1647);
or U844 (N_844,N_544,N_287);
nor U845 (N_845,N_224,In_200);
nor U846 (N_846,In_804,N_32);
xnor U847 (N_847,N_669,In_36);
nand U848 (N_848,In_143,N_307);
nand U849 (N_849,In_1949,N_361);
nand U850 (N_850,N_441,N_300);
xnor U851 (N_851,N_482,In_1739);
nor U852 (N_852,N_501,In_938);
and U853 (N_853,In_246,In_1482);
xnor U854 (N_854,In_1338,N_762);
xor U855 (N_855,N_379,In_1529);
nor U856 (N_856,In_805,N_644);
or U857 (N_857,In_347,In_1737);
or U858 (N_858,In_166,In_1299);
nand U859 (N_859,In_280,In_976);
xor U860 (N_860,In_1968,N_651);
nor U861 (N_861,N_229,In_970);
nor U862 (N_862,N_758,In_555);
nor U863 (N_863,N_568,In_1521);
and U864 (N_864,N_717,N_582);
and U865 (N_865,N_749,In_741);
nand U866 (N_866,In_1435,N_540);
nand U867 (N_867,In_1157,In_1072);
nand U868 (N_868,N_367,N_672);
and U869 (N_869,N_612,In_1089);
xor U870 (N_870,N_120,N_360);
nand U871 (N_871,In_883,In_714);
xnor U872 (N_872,In_695,In_769);
nor U873 (N_873,In_167,In_1117);
xnor U874 (N_874,In_1914,In_708);
nand U875 (N_875,N_753,In_1483);
or U876 (N_876,N_455,In_1668);
or U877 (N_877,In_1942,In_1450);
xnor U878 (N_878,In_1982,N_278);
xor U879 (N_879,N_561,In_506);
xnor U880 (N_880,N_75,In_1214);
or U881 (N_881,In_1991,In_391);
and U882 (N_882,N_190,N_495);
and U883 (N_883,N_543,In_1150);
and U884 (N_884,In_770,N_356);
and U885 (N_885,N_416,N_93);
xor U886 (N_886,In_1712,N_647);
and U887 (N_887,N_667,N_719);
xor U888 (N_888,N_220,In_1611);
and U889 (N_889,N_645,In_12);
nor U890 (N_890,N_565,In_1856);
nand U891 (N_891,N_435,N_742);
and U892 (N_892,N_754,In_212);
xnor U893 (N_893,In_1044,N_701);
or U894 (N_894,In_1093,N_99);
or U895 (N_895,N_43,In_1278);
nor U896 (N_896,N_388,In_1078);
xor U897 (N_897,N_785,In_264);
or U898 (N_898,In_1236,N_512);
and U899 (N_899,In_994,In_196);
or U900 (N_900,In_328,N_663);
and U901 (N_901,In_992,In_350);
nand U902 (N_902,In_1568,N_711);
or U903 (N_903,N_357,N_631);
nor U904 (N_904,In_1573,In_1867);
nor U905 (N_905,N_438,In_500);
or U906 (N_906,In_609,In_595);
or U907 (N_907,N_310,N_494);
or U908 (N_908,N_586,In_1274);
nand U909 (N_909,In_358,N_466);
or U910 (N_910,In_1918,N_428);
and U911 (N_911,In_1807,N_366);
or U912 (N_912,N_60,In_457);
xnor U913 (N_913,N_695,N_793);
nand U914 (N_914,In_1201,N_297);
xor U915 (N_915,In_1166,In_755);
nand U916 (N_916,In_981,N_204);
or U917 (N_917,In_459,N_439);
or U918 (N_918,N_242,In_786);
or U919 (N_919,In_1136,In_538);
nor U920 (N_920,In_1049,In_1723);
and U921 (N_921,In_1733,In_1116);
or U922 (N_922,In_1449,N_614);
nand U923 (N_923,N_346,In_1266);
and U924 (N_924,In_1927,In_121);
nand U925 (N_925,N_497,In_1898);
and U926 (N_926,In_1630,In_471);
and U927 (N_927,N_618,In_882);
nand U928 (N_928,In_984,N_119);
or U929 (N_929,In_398,N_271);
xnor U930 (N_930,N_457,In_1312);
xor U931 (N_931,N_78,In_1127);
nand U932 (N_932,N_426,In_1486);
xor U933 (N_933,N_698,N_572);
nand U934 (N_934,N_581,N_538);
nor U935 (N_935,N_118,In_892);
and U936 (N_936,N_646,In_1788);
xor U937 (N_937,N_70,N_354);
or U938 (N_938,N_163,N_475);
nand U939 (N_939,N_687,N_177);
or U940 (N_940,In_712,N_71);
or U941 (N_941,N_710,In_1260);
nor U942 (N_942,N_257,N_450);
and U943 (N_943,In_373,N_161);
nand U944 (N_944,N_720,In_126);
nor U945 (N_945,In_297,In_556);
or U946 (N_946,In_1512,In_859);
and U947 (N_947,In_1144,N_650);
xnor U948 (N_948,N_694,In_1036);
and U949 (N_949,N_452,In_1628);
xor U950 (N_950,In_975,In_763);
nor U951 (N_951,In_222,In_188);
and U952 (N_952,N_150,N_246);
nor U953 (N_953,In_1649,In_269);
nand U954 (N_954,N_601,In_1817);
xnor U955 (N_955,In_73,N_624);
xnor U956 (N_956,N_128,In_181);
nor U957 (N_957,In_1913,N_140);
xor U958 (N_958,In_655,In_192);
xor U959 (N_959,N_96,N_21);
nor U960 (N_960,In_1447,In_743);
or U961 (N_961,N_513,In_912);
and U962 (N_962,N_649,N_692);
xor U963 (N_963,In_340,N_469);
nor U964 (N_964,In_1308,In_1163);
or U965 (N_965,N_370,N_449);
nand U966 (N_966,In_1925,In_1129);
or U967 (N_967,N_697,N_570);
nand U968 (N_968,In_1177,In_1056);
nor U969 (N_969,In_1990,In_1846);
xor U970 (N_970,N_442,In_211);
nand U971 (N_971,In_1092,In_1758);
nor U972 (N_972,In_915,In_1331);
xnor U973 (N_973,In_1195,In_1987);
and U974 (N_974,N_338,N_609);
xnor U975 (N_975,N_446,In_168);
xnor U976 (N_976,In_736,N_383);
xnor U977 (N_977,N_418,N_657);
and U978 (N_978,N_235,In_881);
nor U979 (N_979,In_149,In_1121);
xnor U980 (N_980,N_610,N_744);
nand U981 (N_981,In_180,N_102);
or U982 (N_982,N_741,In_1388);
nand U983 (N_983,N_578,In_1675);
nand U984 (N_984,N_106,In_1452);
xnor U985 (N_985,In_1115,In_1289);
and U986 (N_986,In_1531,N_240);
or U987 (N_987,N_170,N_417);
and U988 (N_988,N_693,N_267);
nand U989 (N_989,In_1656,In_1825);
nor U990 (N_990,In_520,N_308);
nand U991 (N_991,In_1714,In_1001);
and U992 (N_992,N_558,N_180);
nand U993 (N_993,N_730,N_691);
or U994 (N_994,N_284,N_620);
and U995 (N_995,In_889,In_592);
nand U996 (N_996,In_1940,In_1608);
and U997 (N_997,In_639,N_227);
or U998 (N_998,N_399,In_58);
or U999 (N_999,In_1722,N_737);
nand U1000 (N_1000,N_727,N_662);
nand U1001 (N_1001,In_1762,N_917);
nand U1002 (N_1002,N_929,In_1234);
xnor U1003 (N_1003,N_826,N_770);
nor U1004 (N_1004,N_830,In_1875);
or U1005 (N_1005,In_928,In_818);
xor U1006 (N_1006,N_935,In_893);
and U1007 (N_1007,In_1375,In_988);
xnor U1008 (N_1008,N_557,In_495);
or U1009 (N_1009,In_1367,N_958);
and U1010 (N_1010,In_1571,N_841);
or U1011 (N_1011,N_874,N_94);
or U1012 (N_1012,In_1503,In_64);
nor U1013 (N_1013,In_197,In_1069);
or U1014 (N_1014,N_521,N_760);
or U1015 (N_1015,N_824,In_997);
nand U1016 (N_1016,N_116,N_556);
nand U1017 (N_1017,N_973,N_808);
nor U1018 (N_1018,N_977,N_607);
nand U1019 (N_1019,N_6,In_696);
and U1020 (N_1020,In_1813,N_872);
and U1021 (N_1021,In_638,N_890);
or U1022 (N_1022,In_1416,N_964);
nand U1023 (N_1023,N_272,In_1417);
nand U1024 (N_1024,In_29,In_1795);
xnor U1025 (N_1025,In_1919,In_581);
and U1026 (N_1026,N_722,In_99);
nand U1027 (N_1027,N_704,In_353);
and U1028 (N_1028,N_406,N_619);
xor U1029 (N_1029,N_486,N_816);
nand U1030 (N_1030,In_141,In_1466);
nand U1031 (N_1031,In_722,N_410);
nor U1032 (N_1032,N_132,N_914);
or U1033 (N_1033,In_1921,N_675);
nor U1034 (N_1034,N_992,N_493);
and U1035 (N_1035,N_671,N_323);
nand U1036 (N_1036,N_767,N_769);
and U1037 (N_1037,In_1530,N_403);
or U1038 (N_1038,In_1242,N_273);
nor U1039 (N_1039,In_123,N_664);
nand U1040 (N_1040,N_340,N_861);
nor U1041 (N_1041,N_560,In_1182);
nand U1042 (N_1042,In_519,N_755);
nand U1043 (N_1043,N_792,N_837);
or U1044 (N_1044,N_36,In_1644);
xor U1045 (N_1045,In_1765,In_1703);
and U1046 (N_1046,N_508,In_961);
and U1047 (N_1047,In_14,N_46);
nor U1048 (N_1048,N_983,N_988);
nor U1049 (N_1049,In_417,In_1700);
and U1050 (N_1050,In_671,N_940);
or U1051 (N_1051,N_334,In_233);
xor U1052 (N_1052,In_1340,N_440);
or U1053 (N_1053,In_571,N_212);
and U1054 (N_1054,In_151,N_484);
nor U1055 (N_1055,In_194,N_621);
xnor U1056 (N_1056,N_699,N_528);
nand U1057 (N_1057,N_783,N_846);
nor U1058 (N_1058,N_797,In_907);
nand U1059 (N_1059,In_1587,N_812);
and U1060 (N_1060,In_1726,In_1641);
and U1061 (N_1061,In_1725,N_908);
nor U1062 (N_1062,N_627,In_659);
nand U1063 (N_1063,In_1400,N_774);
or U1064 (N_1064,In_287,N_483);
and U1065 (N_1065,N_941,N_275);
xor U1066 (N_1066,N_424,In_363);
and U1067 (N_1067,N_533,In_670);
nor U1068 (N_1068,In_1969,N_274);
or U1069 (N_1069,In_918,In_1590);
xor U1070 (N_1070,N_880,N_633);
and U1071 (N_1071,N_943,In_1804);
nor U1072 (N_1072,In_1009,N_129);
xnor U1073 (N_1073,In_238,In_1269);
and U1074 (N_1074,In_288,N_945);
or U1075 (N_1075,N_930,N_775);
nor U1076 (N_1076,N_776,In_1751);
xnor U1077 (N_1077,N_833,In_1404);
nand U1078 (N_1078,In_806,In_1458);
and U1079 (N_1079,N_534,N_464);
xor U1080 (N_1080,N_40,N_499);
nand U1081 (N_1081,N_642,N_787);
nand U1082 (N_1082,N_784,N_19);
or U1083 (N_1083,N_590,N_436);
nand U1084 (N_1084,In_18,N_653);
and U1085 (N_1085,In_1429,N_721);
xnor U1086 (N_1086,N_566,N_233);
and U1087 (N_1087,N_858,N_680);
xnor U1088 (N_1088,N_576,N_387);
or U1089 (N_1089,In_1926,N_928);
nor U1090 (N_1090,N_994,In_1353);
nor U1091 (N_1091,In_885,N_884);
nand U1092 (N_1092,In_1818,In_761);
xor U1093 (N_1093,N_766,N_835);
and U1094 (N_1094,In_1775,In_768);
and U1095 (N_1095,In_1614,In_824);
nand U1096 (N_1096,In_1344,In_1588);
or U1097 (N_1097,N_29,N_987);
nand U1098 (N_1098,N_309,In_1636);
xnor U1099 (N_1099,N_665,N_113);
nor U1100 (N_1100,In_720,In_1307);
and U1101 (N_1101,N_321,N_504);
nand U1102 (N_1102,N_571,N_688);
or U1103 (N_1103,N_74,N_971);
or U1104 (N_1104,N_423,In_1498);
nor U1105 (N_1105,In_21,In_478);
nand U1106 (N_1106,N_873,N_849);
and U1107 (N_1107,N_901,N_549);
xnor U1108 (N_1108,N_966,N_244);
nor U1109 (N_1109,In_25,N_529);
or U1110 (N_1110,N_41,In_1862);
xnor U1111 (N_1111,In_148,N_479);
nand U1112 (N_1112,In_782,In_965);
and U1113 (N_1113,N_606,N_724);
xor U1114 (N_1114,N_867,N_3);
nor U1115 (N_1115,In_515,N_965);
nor U1116 (N_1116,N_739,N_937);
and U1117 (N_1117,N_993,In_512);
or U1118 (N_1118,In_1833,In_1950);
xor U1119 (N_1119,In_135,N_811);
and U1120 (N_1120,In_1749,N_592);
nor U1121 (N_1121,N_962,N_836);
nand U1122 (N_1122,N_828,In_488);
and U1123 (N_1123,N_324,N_798);
nand U1124 (N_1124,N_822,N_634);
xor U1125 (N_1125,N_790,In_635);
nor U1126 (N_1126,In_832,N_921);
nor U1127 (N_1127,In_811,N_716);
xnor U1128 (N_1128,N_952,In_1839);
xor U1129 (N_1129,In_1966,N_876);
nand U1130 (N_1130,N_690,N_810);
xor U1131 (N_1131,N_604,N_492);
nor U1132 (N_1132,In_137,In_798);
nand U1133 (N_1133,In_1258,N_696);
nand U1134 (N_1134,In_1972,N_461);
nor U1135 (N_1135,N_451,In_1215);
and U1136 (N_1136,N_124,In_684);
nand U1137 (N_1137,N_840,N_751);
nand U1138 (N_1138,In_1522,In_1574);
nand U1139 (N_1139,N_823,In_1351);
and U1140 (N_1140,N_511,In_837);
and U1141 (N_1141,In_1296,In_57);
or U1142 (N_1142,N_639,N_577);
or U1143 (N_1143,N_718,In_865);
nor U1144 (N_1144,In_496,N_682);
or U1145 (N_1145,N_133,In_1378);
and U1146 (N_1146,N_655,N_55);
nor U1147 (N_1147,In_207,N_902);
nor U1148 (N_1148,N_419,In_1883);
xor U1149 (N_1149,N_815,N_738);
nand U1150 (N_1150,N_900,N_918);
xnor U1151 (N_1151,In_1810,In_1004);
nor U1152 (N_1152,N_507,N_613);
nand U1153 (N_1153,In_434,N_817);
or U1154 (N_1154,In_724,N_676);
xor U1155 (N_1155,In_351,N_405);
nand U1156 (N_1156,N_668,N_949);
and U1157 (N_1157,N_114,In_657);
or U1158 (N_1158,In_321,In_511);
and U1159 (N_1159,In_800,N_115);
nand U1160 (N_1160,N_842,N_584);
and U1161 (N_1161,N_462,In_526);
xnor U1162 (N_1162,N_530,N_262);
or U1163 (N_1163,In_728,In_833);
nor U1164 (N_1164,N_686,N_230);
or U1165 (N_1165,N_878,N_550);
nand U1166 (N_1166,N_654,In_261);
nand U1167 (N_1167,In_578,N_919);
xnor U1168 (N_1168,In_114,N_804);
nand U1169 (N_1169,In_1924,N_942);
nor U1170 (N_1170,N_247,N_376);
or U1171 (N_1171,N_215,In_789);
nand U1172 (N_1172,In_1953,In_348);
or U1173 (N_1173,In_591,In_1645);
nor U1174 (N_1174,N_827,N_907);
or U1175 (N_1175,N_305,N_905);
nand U1176 (N_1176,N_219,N_870);
nor U1177 (N_1177,N_487,In_343);
xor U1178 (N_1178,In_1500,In_697);
xor U1179 (N_1179,N_871,N_803);
xnor U1180 (N_1180,N_293,N_413);
nand U1181 (N_1181,N_794,N_909);
xnor U1182 (N_1182,N_648,N_195);
and U1183 (N_1183,N_747,In_418);
and U1184 (N_1184,N_851,N_875);
nor U1185 (N_1185,N_893,N_957);
nand U1186 (N_1186,In_1958,In_290);
xnor U1187 (N_1187,In_1947,N_277);
nand U1188 (N_1188,In_1481,N_972);
nand U1189 (N_1189,In_1792,N_801);
and U1190 (N_1190,N_159,In_1616);
nand U1191 (N_1191,In_245,In_1543);
or U1192 (N_1192,In_252,In_1687);
nand U1193 (N_1193,N_396,N_637);
nand U1194 (N_1194,N_674,N_526);
nand U1195 (N_1195,In_97,N_254);
or U1196 (N_1196,N_537,N_975);
nand U1197 (N_1197,In_1013,In_390);
and U1198 (N_1198,N_997,N_97);
or U1199 (N_1199,N_832,In_1728);
nor U1200 (N_1200,N_954,N_589);
and U1201 (N_1201,In_738,N_814);
and U1202 (N_1202,N_524,In_1556);
xor U1203 (N_1203,In_904,N_894);
and U1204 (N_1204,N_998,N_903);
nand U1205 (N_1205,N_1012,In_355);
nor U1206 (N_1206,N_1082,N_18);
nor U1207 (N_1207,N_179,N_628);
xnor U1208 (N_1208,N_927,N_1188);
and U1209 (N_1209,N_920,In_324);
nand U1210 (N_1210,N_700,In_588);
nor U1211 (N_1211,N_1016,N_889);
xor U1212 (N_1212,N_397,N_1144);
nand U1213 (N_1213,N_146,In_1606);
nor U1214 (N_1214,In_1803,N_756);
nand U1215 (N_1215,N_961,In_1365);
and U1216 (N_1216,N_108,In_142);
and U1217 (N_1217,In_1903,N_1070);
and U1218 (N_1218,N_1001,In_1699);
xnor U1219 (N_1219,In_1445,In_1534);
xnor U1220 (N_1220,In_1524,N_1186);
and U1221 (N_1221,N_605,N_103);
nor U1222 (N_1222,N_295,N_35);
or U1223 (N_1223,N_1004,N_473);
and U1224 (N_1224,In_1851,N_979);
xor U1225 (N_1225,N_1044,N_1150);
and U1226 (N_1226,N_882,In_629);
xor U1227 (N_1227,N_1112,In_669);
and U1228 (N_1228,N_1100,N_453);
nand U1229 (N_1229,In_1132,N_899);
or U1230 (N_1230,N_809,In_1183);
or U1231 (N_1231,In_823,In_926);
or U1232 (N_1232,N_1141,N_892);
xor U1233 (N_1233,N_1184,In_835);
nor U1234 (N_1234,N_1108,In_1706);
nand U1235 (N_1235,In_1216,In_876);
nand U1236 (N_1236,In_1414,N_384);
nand U1237 (N_1237,N_476,N_860);
nor U1238 (N_1238,N_172,N_444);
or U1239 (N_1239,N_1197,In_1812);
or U1240 (N_1240,In_0,In_38);
and U1241 (N_1241,N_422,N_447);
or U1242 (N_1242,N_970,N_895);
and U1243 (N_1243,N_853,N_891);
xor U1244 (N_1244,In_1808,N_101);
or U1245 (N_1245,N_1024,N_1088);
and U1246 (N_1246,N_1095,In_1147);
nor U1247 (N_1247,In_620,In_845);
or U1248 (N_1248,N_1071,In_1691);
xor U1249 (N_1249,In_1863,In_9);
nand U1250 (N_1250,N_1077,N_630);
and U1251 (N_1251,N_926,N_251);
or U1252 (N_1252,N_679,N_632);
or U1253 (N_1253,N_1157,N_1025);
nand U1254 (N_1254,N_881,N_331);
or U1255 (N_1255,N_915,N_1028);
or U1256 (N_1256,N_839,N_1042);
and U1257 (N_1257,N_1168,N_764);
and U1258 (N_1258,In_438,N_825);
nand U1259 (N_1259,N_463,N_1159);
or U1260 (N_1260,In_586,N_996);
and U1261 (N_1261,N_151,In_1769);
xnor U1262 (N_1262,N_947,N_1039);
and U1263 (N_1263,N_593,N_594);
nand U1264 (N_1264,N_1174,In_851);
nand U1265 (N_1265,N_879,N_316);
xor U1266 (N_1266,N_896,N_855);
nand U1267 (N_1267,In_640,N_1134);
xor U1268 (N_1268,N_805,N_1191);
nand U1269 (N_1269,In_819,N_913);
or U1270 (N_1270,In_691,In_1142);
and U1271 (N_1271,In_441,N_1137);
or U1272 (N_1272,N_1047,N_1121);
nand U1273 (N_1273,N_933,N_296);
or U1274 (N_1274,In_1276,In_1558);
and U1275 (N_1275,N_877,N_1033);
nand U1276 (N_1276,N_1161,N_532);
nand U1277 (N_1277,N_110,In_1074);
or U1278 (N_1278,N_1034,N_656);
nand U1279 (N_1279,N_597,In_1952);
nor U1280 (N_1280,N_1175,N_1138);
and U1281 (N_1281,In_281,N_723);
nand U1282 (N_1282,N_981,In_153);
or U1283 (N_1283,N_1139,N_427);
or U1284 (N_1284,N_1005,N_67);
nor U1285 (N_1285,In_1030,N_706);
nand U1286 (N_1286,In_636,N_58);
xnor U1287 (N_1287,N_883,In_780);
nor U1288 (N_1288,In_1674,In_1230);
or U1289 (N_1289,In_621,In_1431);
nor U1290 (N_1290,N_509,N_1199);
xnor U1291 (N_1291,In_1027,In_1967);
and U1292 (N_1292,In_1291,In_1663);
xnor U1293 (N_1293,N_1131,In_1665);
xor U1294 (N_1294,In_454,N_595);
or U1295 (N_1295,In_1376,N_773);
or U1296 (N_1296,N_364,N_395);
and U1297 (N_1297,N_745,N_910);
xnor U1298 (N_1298,N_1167,N_1050);
nor U1299 (N_1299,N_640,N_1045);
or U1300 (N_1300,N_898,N_951);
and U1301 (N_1301,N_788,In_1976);
nand U1302 (N_1302,In_1493,N_175);
xor U1303 (N_1303,In_1837,In_311);
or U1304 (N_1304,In_147,N_616);
nand U1305 (N_1305,In_1826,N_1015);
nor U1306 (N_1306,In_505,N_412);
nor U1307 (N_1307,N_862,N_732);
nor U1308 (N_1308,N_944,N_740);
nor U1309 (N_1309,N_1114,N_938);
or U1310 (N_1310,N_1026,N_684);
and U1311 (N_1311,N_729,In_468);
nor U1312 (N_1312,N_1059,N_931);
nor U1313 (N_1313,N_1193,In_878);
nand U1314 (N_1314,N_968,In_1229);
or U1315 (N_1315,N_1125,N_750);
and U1316 (N_1316,N_600,N_1073);
and U1317 (N_1317,N_1007,N_777);
and U1318 (N_1318,N_1118,N_1180);
xor U1319 (N_1319,N_932,N_1146);
nor U1320 (N_1320,N_336,N_559);
nor U1321 (N_1321,N_1123,In_787);
and U1322 (N_1322,In_1456,N_673);
nor U1323 (N_1323,In_871,N_1115);
nand U1324 (N_1324,N_1182,In_206);
xor U1325 (N_1325,N_1110,N_635);
and U1326 (N_1326,N_1195,N_1013);
or U1327 (N_1327,In_547,In_1313);
nor U1328 (N_1328,N_1080,In_1319);
nor U1329 (N_1329,In_968,N_1148);
or U1330 (N_1330,N_1084,N_1096);
or U1331 (N_1331,N_575,In_1393);
xnor U1332 (N_1332,In_1461,N_432);
nor U1333 (N_1333,N_602,N_906);
nand U1334 (N_1334,In_1167,N_1153);
nor U1335 (N_1335,N_1048,In_1563);
nor U1336 (N_1336,N_554,In_445);
xor U1337 (N_1337,N_847,N_897);
nor U1338 (N_1338,In_1901,In_1612);
nor U1339 (N_1339,In_1520,In_1579);
nor U1340 (N_1340,N_866,In_90);
and U1341 (N_1341,In_922,N_1020);
xor U1342 (N_1342,N_759,N_282);
or U1343 (N_1343,N_1064,In_476);
xor U1344 (N_1344,N_525,N_1171);
xnor U1345 (N_1345,In_316,N_806);
or U1346 (N_1346,In_1071,N_1156);
or U1347 (N_1347,N_144,N_1017);
nand U1348 (N_1348,N_829,In_42);
or U1349 (N_1349,N_1002,In_421);
xor U1350 (N_1350,N_518,N_641);
nor U1351 (N_1351,N_553,N_82);
xor U1352 (N_1352,In_790,N_925);
nor U1353 (N_1353,In_711,N_500);
nand U1354 (N_1354,N_1163,In_1448);
xnor U1355 (N_1355,N_1122,N_1068);
or U1356 (N_1356,In_788,N_1091);
nor U1357 (N_1357,N_904,In_236);
or U1358 (N_1358,N_522,N_956);
nand U1359 (N_1359,N_1128,N_780);
or U1360 (N_1360,N_1014,N_329);
or U1361 (N_1361,N_617,N_527);
and U1362 (N_1362,In_82,N_1066);
nand U1363 (N_1363,N_141,N_636);
nor U1364 (N_1364,N_850,N_1061);
or U1365 (N_1365,N_1187,N_1000);
nand U1366 (N_1366,N_1140,N_1097);
nor U1367 (N_1367,N_807,In_122);
xor U1368 (N_1368,In_67,N_748);
or U1369 (N_1369,N_318,N_888);
xnor U1370 (N_1370,N_1145,N_802);
nor U1371 (N_1371,N_1151,N_623);
and U1372 (N_1372,In_298,N_1190);
nand U1373 (N_1373,N_819,N_1189);
nor U1374 (N_1374,N_76,N_967);
or U1375 (N_1375,N_959,N_924);
and U1376 (N_1376,N_1119,In_1720);
or U1377 (N_1377,N_800,In_1411);
or U1378 (N_1378,N_562,In_694);
and U1379 (N_1379,N_934,N_1173);
nand U1380 (N_1380,In_1080,In_1546);
and U1381 (N_1381,N_1027,In_1986);
nand U1382 (N_1382,N_677,N_92);
nor U1383 (N_1383,In_1014,N_299);
nand U1384 (N_1384,In_1135,N_818);
xor U1385 (N_1385,In_223,N_1099);
or U1386 (N_1386,N_1063,N_1116);
nor U1387 (N_1387,In_263,N_545);
xnor U1388 (N_1388,In_1179,N_345);
or U1389 (N_1389,In_1124,In_1272);
xnor U1390 (N_1390,N_471,N_733);
xor U1391 (N_1391,In_1885,In_1220);
nor U1392 (N_1392,N_1036,N_573);
nor U1393 (N_1393,N_999,N_201);
nor U1394 (N_1394,N_1093,In_489);
or U1395 (N_1395,N_429,N_234);
xor U1396 (N_1396,N_652,In_1394);
or U1397 (N_1397,In_1821,N_629);
and U1398 (N_1398,N_353,N_1006);
and U1399 (N_1399,In_1087,In_1322);
xnor U1400 (N_1400,N_276,N_1065);
nor U1401 (N_1401,N_1333,N_1233);
nor U1402 (N_1402,In_1957,N_517);
nor U1403 (N_1403,In_740,N_1292);
nand U1404 (N_1404,In_217,In_1827);
nor U1405 (N_1405,N_531,N_420);
and U1406 (N_1406,N_821,N_1373);
and U1407 (N_1407,N_1294,N_1194);
or U1408 (N_1408,In_70,N_208);
nor U1409 (N_1409,N_1041,N_1391);
xnor U1410 (N_1410,In_900,N_1397);
and U1411 (N_1411,N_752,N_1213);
nand U1412 (N_1412,N_781,N_1354);
nor U1413 (N_1413,N_503,N_1087);
nand U1414 (N_1414,N_1057,In_737);
or U1415 (N_1415,N_1075,In_1347);
nor U1416 (N_1416,In_1945,N_1120);
xor U1417 (N_1417,N_1357,N_1244);
nand U1418 (N_1418,In_759,In_1761);
or U1419 (N_1419,N_1330,N_1386);
or U1420 (N_1420,N_795,In_13);
xor U1421 (N_1421,In_908,N_1086);
xor U1422 (N_1422,N_1222,In_1609);
or U1423 (N_1423,N_712,N_1388);
nand U1424 (N_1424,In_589,N_1287);
xor U1425 (N_1425,In_52,N_448);
xor U1426 (N_1426,N_1051,N_1142);
and U1427 (N_1427,N_659,N_1378);
nor U1428 (N_1428,N_1379,N_1255);
and U1429 (N_1429,N_845,N_864);
and U1430 (N_1430,N_986,In_1653);
and U1431 (N_1431,In_1595,N_1266);
or U1432 (N_1432,N_285,N_355);
xnor U1433 (N_1433,In_416,N_1253);
nand U1434 (N_1434,In_475,In_1426);
nand U1435 (N_1435,N_1268,N_1018);
xnor U1436 (N_1436,N_1105,In_749);
nand U1437 (N_1437,N_1343,In_825);
nor U1438 (N_1438,N_48,In_54);
nand U1439 (N_1439,N_923,N_1179);
nand U1440 (N_1440,N_886,N_400);
nand U1441 (N_1441,N_1226,N_1261);
xor U1442 (N_1442,N_1098,N_1126);
xnor U1443 (N_1443,N_1392,In_1859);
and U1444 (N_1444,N_1076,N_1106);
and U1445 (N_1445,N_685,N_705);
nand U1446 (N_1446,N_488,N_946);
or U1447 (N_1447,N_912,N_328);
nand U1448 (N_1448,N_1382,N_1009);
and U1449 (N_1449,N_1365,N_1327);
or U1450 (N_1450,N_1183,N_1085);
nor U1451 (N_1451,In_1484,N_1239);
xor U1452 (N_1452,N_1228,N_746);
nor U1453 (N_1453,N_1214,In_971);
xor U1454 (N_1454,N_281,N_1285);
and U1455 (N_1455,N_91,N_1201);
nand U1456 (N_1456,N_421,N_1277);
nand U1457 (N_1457,In_1040,N_433);
xor U1458 (N_1458,N_1362,N_1053);
nand U1459 (N_1459,N_615,N_1217);
nor U1460 (N_1460,N_1216,N_226);
xor U1461 (N_1461,In_848,In_86);
and U1462 (N_1462,In_570,In_792);
and U1463 (N_1463,N_955,N_731);
nor U1464 (N_1464,N_1055,In_1519);
xor U1465 (N_1465,N_969,N_734);
xnor U1466 (N_1466,N_1306,N_1074);
and U1467 (N_1467,N_1166,N_1282);
or U1468 (N_1468,N_1218,N_854);
xnor U1469 (N_1469,N_1160,N_1072);
nor U1470 (N_1470,In_1439,N_625);
and U1471 (N_1471,N_50,N_1318);
nor U1472 (N_1472,N_1103,N_948);
nand U1473 (N_1473,In_100,N_1181);
nor U1474 (N_1474,N_728,N_922);
nor U1475 (N_1475,N_1270,In_270);
xnor U1476 (N_1476,N_1321,In_448);
nor U1477 (N_1477,In_79,N_1236);
and U1478 (N_1478,N_1249,N_1364);
or U1479 (N_1479,In_894,N_848);
nand U1480 (N_1480,N_885,N_1288);
xor U1481 (N_1481,N_1247,N_1221);
and U1482 (N_1482,In_1715,N_736);
xor U1483 (N_1483,N_294,N_1035);
nand U1484 (N_1484,N_1062,N_768);
nor U1485 (N_1485,In_1801,N_838);
or U1486 (N_1486,N_1069,In_1742);
nor U1487 (N_1487,In_613,N_995);
nor U1488 (N_1488,In_1169,N_1308);
nand U1489 (N_1489,N_1325,N_865);
nand U1490 (N_1490,N_1052,N_1154);
xnor U1491 (N_1491,N_514,N_1374);
or U1492 (N_1492,N_1310,N_1368);
nand U1493 (N_1493,N_591,In_1549);
nor U1494 (N_1494,N_643,N_1324);
nor U1495 (N_1495,N_1037,N_1019);
and U1496 (N_1496,N_390,N_1229);
xor U1497 (N_1497,In_113,N_1272);
or U1498 (N_1498,In_978,In_676);
and U1499 (N_1499,In_48,N_953);
or U1500 (N_1500,N_1211,N_1049);
and U1501 (N_1501,N_1078,In_580);
nand U1502 (N_1502,N_1383,N_991);
nand U1503 (N_1503,N_1212,N_1328);
and U1504 (N_1504,N_1284,N_1370);
nor U1505 (N_1505,In_1756,N_1242);
xnor U1506 (N_1506,N_135,In_203);
nand U1507 (N_1507,N_1147,N_1300);
or U1508 (N_1508,N_1162,N_1235);
and U1509 (N_1509,In_1978,N_1207);
nor U1510 (N_1510,N_1319,In_1783);
or U1511 (N_1511,In_717,N_1023);
or U1512 (N_1512,N_1317,N_1203);
nand U1513 (N_1513,N_1279,N_1254);
and U1514 (N_1514,N_225,N_79);
nor U1515 (N_1515,N_1298,N_1101);
or U1516 (N_1516,N_1309,In_1844);
nor U1517 (N_1517,N_1381,N_661);
or U1518 (N_1518,N_1130,N_1297);
and U1519 (N_1519,N_1102,N_1315);
and U1520 (N_1520,N_869,In_1545);
and U1521 (N_1521,N_1352,N_976);
and U1522 (N_1522,N_1312,N_1079);
nand U1523 (N_1523,In_957,N_1132);
nand U1524 (N_1524,N_1267,N_1305);
or U1525 (N_1525,N_1081,In_540);
xnor U1526 (N_1526,In_93,N_985);
nand U1527 (N_1527,In_234,N_1043);
or U1528 (N_1528,N_820,N_523);
or U1529 (N_1529,N_404,N_1092);
and U1530 (N_1530,In_1193,N_1010);
nor U1531 (N_1531,In_1581,N_1329);
xor U1532 (N_1532,N_1399,In_247);
xnor U1533 (N_1533,In_1680,N_157);
and U1534 (N_1534,N_1363,N_1264);
or U1535 (N_1535,N_1143,In_1904);
nor U1536 (N_1536,In_1227,In_801);
and U1537 (N_1537,In_767,In_1428);
or U1538 (N_1538,In_174,In_1928);
xor U1539 (N_1539,N_725,N_1240);
nor U1540 (N_1540,N_763,N_1104);
xor U1541 (N_1541,In_852,N_1202);
nand U1542 (N_1542,N_1124,N_765);
and U1543 (N_1543,In_1509,N_1273);
or U1544 (N_1544,N_1347,N_481);
or U1545 (N_1545,N_456,N_856);
or U1546 (N_1546,N_707,N_1271);
and U1547 (N_1547,N_289,In_1669);
and U1548 (N_1548,N_713,N_1262);
nor U1549 (N_1549,N_1155,N_1278);
xor U1550 (N_1550,N_1387,In_1306);
xnor U1551 (N_1551,N_990,N_1299);
and U1552 (N_1552,N_342,N_1355);
nand U1553 (N_1553,N_868,N_1196);
or U1554 (N_1554,N_1313,In_187);
and U1555 (N_1555,In_1750,N_1296);
nand U1556 (N_1556,In_910,N_950);
or U1557 (N_1557,N_796,In_451);
or U1558 (N_1558,N_1339,N_1257);
xnor U1559 (N_1559,N_498,N_1136);
xor U1560 (N_1560,N_1170,N_1058);
or U1561 (N_1561,N_799,N_1275);
nor U1562 (N_1562,In_98,N_256);
or U1563 (N_1563,N_1209,N_1353);
nor U1564 (N_1564,N_1204,N_1366);
or U1565 (N_1565,N_1344,N_1276);
or U1566 (N_1566,N_670,N_757);
or U1567 (N_1567,In_1140,N_1398);
nand U1568 (N_1568,N_1263,N_1316);
xor U1569 (N_1569,N_1377,N_1056);
nand U1570 (N_1570,N_1224,In_1617);
or U1571 (N_1571,N_459,N_368);
nor U1572 (N_1572,N_1367,N_1248);
and U1573 (N_1573,N_960,In_377);
and U1574 (N_1574,N_1129,In_1055);
or U1575 (N_1575,N_1265,In_602);
xor U1576 (N_1576,N_131,N_467);
nand U1577 (N_1577,N_542,N_936);
nor U1578 (N_1578,N_1384,N_1295);
or U1579 (N_1579,In_1422,In_414);
xnor U1580 (N_1580,N_1380,N_279);
xnor U1581 (N_1581,N_1220,N_1011);
or U1582 (N_1582,N_1250,N_1107);
or U1583 (N_1583,N_1291,N_1260);
nand U1584 (N_1584,N_1237,N_1113);
or U1585 (N_1585,N_678,In_463);
nor U1586 (N_1586,N_1176,N_611);
nor U1587 (N_1587,N_1338,N_1165);
nand U1588 (N_1588,N_1178,In_23);
or U1589 (N_1589,N_1345,N_1054);
and U1590 (N_1590,N_1337,N_681);
nand U1591 (N_1591,In_1889,N_1293);
nand U1592 (N_1592,N_1031,N_911);
nor U1593 (N_1593,N_1234,N_1280);
nor U1594 (N_1594,In_1845,N_1395);
nor U1595 (N_1595,N_1246,N_1185);
and U1596 (N_1596,N_1256,N_1269);
and U1597 (N_1597,N_1205,In_1356);
nor U1598 (N_1598,N_1361,N_982);
xnor U1599 (N_1599,In_286,N_989);
and U1600 (N_1600,N_1400,N_1481);
and U1601 (N_1601,N_1589,N_1425);
or U1602 (N_1602,N_1543,N_1164);
nand U1603 (N_1603,N_1545,N_1434);
or U1604 (N_1604,N_1371,In_56);
xnor U1605 (N_1605,N_214,N_1536);
or U1606 (N_1606,N_1436,N_1417);
or U1607 (N_1607,N_1304,In_1847);
or U1608 (N_1608,N_1489,N_857);
or U1609 (N_1609,In_1370,N_844);
and U1610 (N_1610,N_1506,In_1828);
or U1611 (N_1611,N_714,N_1549);
xnor U1612 (N_1612,N_1480,N_1432);
nand U1613 (N_1613,N_1556,N_1408);
and U1614 (N_1614,N_1227,N_1564);
and U1615 (N_1615,N_1407,N_1430);
nor U1616 (N_1616,N_963,N_1349);
nor U1617 (N_1617,N_1200,N_1498);
nor U1618 (N_1618,N_1421,N_1029);
xor U1619 (N_1619,N_1431,N_1067);
and U1620 (N_1620,N_1369,N_1320);
and U1621 (N_1621,N_1516,N_1460);
xor U1622 (N_1622,In_1661,N_863);
xnor U1623 (N_1623,N_1356,N_1443);
xor U1624 (N_1624,In_354,N_1530);
nand U1625 (N_1625,N_1410,N_660);
or U1626 (N_1626,N_1094,N_1494);
and U1627 (N_1627,N_1538,N_250);
nand U1628 (N_1628,N_1360,N_1472);
nor U1629 (N_1629,N_261,N_1340);
xor U1630 (N_1630,N_1462,N_666);
nand U1631 (N_1631,N_1450,N_182);
or U1632 (N_1632,N_1418,N_1429);
nor U1633 (N_1633,N_1563,N_1350);
xnor U1634 (N_1634,In_397,In_81);
and U1635 (N_1635,In_452,N_1572);
nand U1636 (N_1636,N_1562,N_1520);
nor U1637 (N_1637,N_326,N_1133);
nand U1638 (N_1638,N_1326,N_1457);
nand U1639 (N_1639,N_786,N_1554);
and U1640 (N_1640,N_1442,N_887);
xnor U1641 (N_1641,N_1445,N_1437);
xnor U1642 (N_1642,N_1453,N_1485);
and U1643 (N_1643,N_1464,N_1289);
or U1644 (N_1644,N_1302,N_1060);
and U1645 (N_1645,N_1459,N_1493);
nor U1646 (N_1646,N_1559,N_1461);
xnor U1647 (N_1647,In_1155,N_1473);
xnor U1648 (N_1648,N_834,N_1567);
xnor U1649 (N_1649,N_1534,N_1513);
nand U1650 (N_1650,N_1358,In_1264);
or U1651 (N_1651,In_874,N_1465);
and U1652 (N_1652,N_1348,In_1770);
xnor U1653 (N_1653,N_703,N_1238);
or U1654 (N_1654,N_1008,N_1420);
or U1655 (N_1655,N_280,N_1507);
nand U1656 (N_1656,N_1149,N_978);
xor U1657 (N_1657,N_1585,N_1415);
nand U1658 (N_1658,In_94,In_47);
nor U1659 (N_1659,N_1413,N_1510);
and U1660 (N_1660,N_1514,N_1479);
nor U1661 (N_1661,N_1258,N_1484);
xor U1662 (N_1662,N_1511,N_1575);
nand U1663 (N_1663,N_1411,N_1083);
or U1664 (N_1664,N_1500,N_1535);
nor U1665 (N_1665,N_1566,N_1422);
and U1666 (N_1666,N_515,N_1581);
nor U1667 (N_1667,In_1776,N_1286);
nand U1668 (N_1668,N_1223,N_1283);
or U1669 (N_1669,N_1111,N_1515);
or U1670 (N_1670,N_843,In_597);
and U1671 (N_1671,N_1597,In_544);
nand U1672 (N_1672,N_1152,N_1331);
and U1673 (N_1673,N_1230,N_596);
and U1674 (N_1674,N_1522,N_1243);
nor U1675 (N_1675,N_1389,N_984);
nor U1676 (N_1676,N_1558,N_1586);
and U1677 (N_1677,N_164,N_1490);
nand U1678 (N_1678,N_1496,N_1590);
nor U1679 (N_1679,N_1588,N_1405);
and U1680 (N_1680,N_1341,N_1503);
or U1681 (N_1681,N_1548,N_1351);
nor U1682 (N_1682,N_1419,N_939);
nand U1683 (N_1683,N_1449,N_1529);
nand U1684 (N_1684,N_1525,N_1441);
xnor U1685 (N_1685,N_1206,N_1458);
or U1686 (N_1686,N_1332,N_1252);
and U1687 (N_1687,N_1426,N_1231);
xor U1688 (N_1688,N_1446,N_1497);
nor U1689 (N_1689,N_1463,N_1022);
or U1690 (N_1690,N_743,In_1334);
and U1691 (N_1691,N_1040,N_1523);
and U1692 (N_1692,N_1478,N_16);
xor U1693 (N_1693,N_1435,N_1215);
xnor U1694 (N_1694,N_1090,N_1396);
and U1695 (N_1695,N_1576,N_1281);
nand U1696 (N_1696,N_1471,N_506);
nand U1697 (N_1697,N_1482,N_1438);
nand U1698 (N_1698,N_1487,In_71);
or U1699 (N_1699,N_1393,N_1427);
xor U1700 (N_1700,N_772,N_1583);
or U1701 (N_1701,N_709,In_858);
and U1702 (N_1702,N_1467,In_190);
nor U1703 (N_1703,In_49,N_1375);
and U1704 (N_1704,N_1135,N_1251);
nor U1705 (N_1705,In_1008,N_192);
nor U1706 (N_1706,In_480,N_1158);
nand U1707 (N_1707,In_1943,N_726);
xnor U1708 (N_1708,N_1342,N_1533);
nand U1709 (N_1709,N_708,N_1447);
nor U1710 (N_1710,In_797,N_603);
and U1711 (N_1711,N_1501,N_1322);
and U1712 (N_1712,N_1172,N_1577);
nor U1713 (N_1713,N_1127,N_1492);
xor U1714 (N_1714,N_1596,N_1169);
and U1715 (N_1715,N_1495,N_813);
nand U1716 (N_1716,N_1046,N_1518);
or U1717 (N_1717,N_1334,N_260);
and U1718 (N_1718,N_1394,N_1030);
nand U1719 (N_1719,N_1521,N_1499);
and U1720 (N_1720,In_1811,N_1359);
nor U1721 (N_1721,N_1390,N_1504);
nand U1722 (N_1722,In_645,N_1470);
or U1723 (N_1723,In_1427,N_974);
or U1724 (N_1724,N_239,In_1277);
and U1725 (N_1725,N_1423,N_1477);
nand U1726 (N_1726,N_1451,N_1593);
or U1727 (N_1727,N_852,N_365);
nor U1728 (N_1728,N_1428,N_1561);
nand U1729 (N_1729,In_332,N_1376);
nor U1730 (N_1730,N_1038,N_1476);
and U1731 (N_1731,N_1444,N_1551);
xor U1732 (N_1732,N_1385,N_431);
nor U1733 (N_1733,In_1794,N_1565);
nand U1734 (N_1734,In_68,N_1526);
nor U1735 (N_1735,N_1486,N_622);
and U1736 (N_1736,N_1599,N_1594);
xnor U1737 (N_1737,N_1474,N_1311);
nor U1738 (N_1738,N_1595,N_831);
and U1739 (N_1739,N_1560,In_951);
nor U1740 (N_1740,N_1557,N_1323);
or U1741 (N_1741,N_1527,N_1483);
or U1742 (N_1742,N_1546,N_1210);
nor U1743 (N_1743,N_1177,N_1469);
or U1744 (N_1744,N_1274,N_1401);
or U1745 (N_1745,N_1468,N_1109);
nor U1746 (N_1746,N_1574,In_1465);
nand U1747 (N_1747,In_564,N_1488);
nand U1748 (N_1748,N_1532,N_1592);
nor U1749 (N_1749,N_1580,N_1303);
xnor U1750 (N_1750,In_1192,N_1117);
nor U1751 (N_1751,N_1584,N_1225);
and U1752 (N_1752,N_1512,N_1505);
xnor U1753 (N_1753,N_1089,N_1571);
nand U1754 (N_1754,In_62,N_1466);
nand U1755 (N_1755,N_1454,N_1569);
nor U1756 (N_1756,N_1573,N_1439);
nand U1757 (N_1757,N_1003,N_548);
xnor U1758 (N_1758,N_1259,In_456);
and U1759 (N_1759,N_658,N_1335);
or U1760 (N_1760,N_1208,N_490);
xnor U1761 (N_1761,N_1570,N_1502);
and U1762 (N_1762,N_1579,N_1032);
xnor U1763 (N_1763,N_1508,N_1412);
xor U1764 (N_1764,N_1568,N_1528);
and U1765 (N_1765,N_1416,N_86);
or U1766 (N_1766,N_1531,N_437);
nor U1767 (N_1767,N_1509,N_1307);
xor U1768 (N_1768,N_1245,N_1192);
xnor U1769 (N_1769,N_1414,N_1424);
nor U1770 (N_1770,N_1301,N_1519);
nand U1771 (N_1771,In_1081,N_1409);
and U1772 (N_1772,N_1198,N_1550);
nor U1773 (N_1773,N_203,In_517);
nor U1774 (N_1774,In_185,N_415);
xnor U1775 (N_1775,N_1448,N_1403);
and U1776 (N_1776,N_1578,N_1517);
xnor U1777 (N_1777,N_1021,N_1440);
nor U1778 (N_1778,N_1314,N_1372);
and U1779 (N_1779,N_1524,N_1433);
nand U1780 (N_1780,N_322,N_1537);
or U1781 (N_1781,N_69,N_1336);
nand U1782 (N_1782,N_789,N_1491);
xor U1783 (N_1783,N_1539,N_859);
xor U1784 (N_1784,N_1555,N_683);
and U1785 (N_1785,In_646,N_1475);
or U1786 (N_1786,N_1547,N_1587);
nor U1787 (N_1787,N_1552,N_916);
nor U1788 (N_1788,In_1660,N_1346);
and U1789 (N_1789,N_1232,N_1541);
and U1790 (N_1790,N_1219,N_1455);
nand U1791 (N_1791,N_123,N_1591);
nand U1792 (N_1792,N_1542,N_1598);
and U1793 (N_1793,N_980,N_1540);
nand U1794 (N_1794,N_1452,N_1404);
xnor U1795 (N_1795,N_1241,N_1456);
nand U1796 (N_1796,N_377,N_1544);
or U1797 (N_1797,N_1406,In_1225);
and U1798 (N_1798,N_1582,N_1402);
nand U1799 (N_1799,N_1290,N_1553);
xor U1800 (N_1800,N_1683,N_1791);
nor U1801 (N_1801,N_1706,N_1645);
and U1802 (N_1802,N_1705,N_1750);
xor U1803 (N_1803,N_1611,N_1735);
and U1804 (N_1804,N_1764,N_1771);
xnor U1805 (N_1805,N_1660,N_1752);
and U1806 (N_1806,N_1708,N_1635);
nor U1807 (N_1807,N_1648,N_1658);
and U1808 (N_1808,N_1676,N_1702);
or U1809 (N_1809,N_1642,N_1753);
and U1810 (N_1810,N_1798,N_1632);
nand U1811 (N_1811,N_1624,N_1736);
or U1812 (N_1812,N_1758,N_1696);
or U1813 (N_1813,N_1647,N_1685);
xor U1814 (N_1814,N_1672,N_1712);
nand U1815 (N_1815,N_1603,N_1691);
xor U1816 (N_1816,N_1761,N_1649);
nor U1817 (N_1817,N_1626,N_1693);
or U1818 (N_1818,N_1600,N_1663);
and U1819 (N_1819,N_1675,N_1612);
or U1820 (N_1820,N_1748,N_1602);
and U1821 (N_1821,N_1668,N_1733);
xnor U1822 (N_1822,N_1650,N_1621);
and U1823 (N_1823,N_1795,N_1796);
xnor U1824 (N_1824,N_1730,N_1757);
nand U1825 (N_1825,N_1615,N_1629);
nand U1826 (N_1826,N_1667,N_1792);
xor U1827 (N_1827,N_1732,N_1728);
nor U1828 (N_1828,N_1694,N_1794);
or U1829 (N_1829,N_1749,N_1745);
nand U1830 (N_1830,N_1727,N_1608);
nand U1831 (N_1831,N_1627,N_1695);
or U1832 (N_1832,N_1786,N_1759);
and U1833 (N_1833,N_1719,N_1697);
nand U1834 (N_1834,N_1605,N_1690);
nor U1835 (N_1835,N_1716,N_1657);
and U1836 (N_1836,N_1778,N_1737);
nand U1837 (N_1837,N_1684,N_1755);
nand U1838 (N_1838,N_1606,N_1744);
or U1839 (N_1839,N_1709,N_1613);
or U1840 (N_1840,N_1760,N_1666);
nor U1841 (N_1841,N_1742,N_1630);
nand U1842 (N_1842,N_1711,N_1780);
and U1843 (N_1843,N_1622,N_1789);
xor U1844 (N_1844,N_1639,N_1739);
or U1845 (N_1845,N_1665,N_1641);
nand U1846 (N_1846,N_1774,N_1765);
nor U1847 (N_1847,N_1769,N_1715);
or U1848 (N_1848,N_1721,N_1729);
xnor U1849 (N_1849,N_1781,N_1614);
or U1850 (N_1850,N_1674,N_1681);
nor U1851 (N_1851,N_1610,N_1671);
nor U1852 (N_1852,N_1664,N_1618);
and U1853 (N_1853,N_1646,N_1767);
nand U1854 (N_1854,N_1756,N_1625);
nand U1855 (N_1855,N_1634,N_1607);
or U1856 (N_1856,N_1740,N_1723);
or U1857 (N_1857,N_1689,N_1701);
nand U1858 (N_1858,N_1644,N_1718);
nor U1859 (N_1859,N_1777,N_1638);
nand U1860 (N_1860,N_1776,N_1656);
and U1861 (N_1861,N_1604,N_1643);
or U1862 (N_1862,N_1775,N_1637);
nand U1863 (N_1863,N_1703,N_1704);
nand U1864 (N_1864,N_1687,N_1653);
nor U1865 (N_1865,N_1787,N_1640);
nor U1866 (N_1866,N_1710,N_1680);
nand U1867 (N_1867,N_1746,N_1609);
xor U1868 (N_1868,N_1763,N_1636);
or U1869 (N_1869,N_1770,N_1785);
or U1870 (N_1870,N_1747,N_1726);
or U1871 (N_1871,N_1762,N_1790);
and U1872 (N_1872,N_1779,N_1682);
or U1873 (N_1873,N_1633,N_1751);
nor U1874 (N_1874,N_1720,N_1699);
or U1875 (N_1875,N_1722,N_1734);
and U1876 (N_1876,N_1686,N_1713);
xor U1877 (N_1877,N_1698,N_1788);
nand U1878 (N_1878,N_1766,N_1617);
and U1879 (N_1879,N_1724,N_1799);
nor U1880 (N_1880,N_1669,N_1784);
nand U1881 (N_1881,N_1717,N_1700);
nand U1882 (N_1882,N_1768,N_1679);
xor U1883 (N_1883,N_1782,N_1743);
or U1884 (N_1884,N_1731,N_1659);
xor U1885 (N_1885,N_1673,N_1652);
xor U1886 (N_1886,N_1654,N_1616);
xor U1887 (N_1887,N_1670,N_1754);
nor U1888 (N_1888,N_1714,N_1688);
or U1889 (N_1889,N_1772,N_1797);
or U1890 (N_1890,N_1661,N_1773);
xor U1891 (N_1891,N_1692,N_1677);
xor U1892 (N_1892,N_1631,N_1601);
nor U1893 (N_1893,N_1678,N_1619);
or U1894 (N_1894,N_1741,N_1707);
and U1895 (N_1895,N_1738,N_1655);
nand U1896 (N_1896,N_1620,N_1662);
and U1897 (N_1897,N_1783,N_1793);
and U1898 (N_1898,N_1628,N_1651);
nor U1899 (N_1899,N_1623,N_1725);
xor U1900 (N_1900,N_1716,N_1773);
nor U1901 (N_1901,N_1792,N_1719);
xor U1902 (N_1902,N_1656,N_1715);
xor U1903 (N_1903,N_1710,N_1749);
nor U1904 (N_1904,N_1680,N_1738);
or U1905 (N_1905,N_1714,N_1668);
and U1906 (N_1906,N_1677,N_1632);
xnor U1907 (N_1907,N_1740,N_1722);
or U1908 (N_1908,N_1670,N_1706);
xor U1909 (N_1909,N_1701,N_1777);
nor U1910 (N_1910,N_1739,N_1625);
nand U1911 (N_1911,N_1770,N_1613);
and U1912 (N_1912,N_1779,N_1766);
and U1913 (N_1913,N_1742,N_1607);
xnor U1914 (N_1914,N_1727,N_1764);
or U1915 (N_1915,N_1778,N_1671);
xor U1916 (N_1916,N_1641,N_1617);
xnor U1917 (N_1917,N_1757,N_1654);
and U1918 (N_1918,N_1759,N_1620);
nor U1919 (N_1919,N_1675,N_1693);
and U1920 (N_1920,N_1740,N_1625);
nand U1921 (N_1921,N_1733,N_1778);
and U1922 (N_1922,N_1672,N_1718);
nor U1923 (N_1923,N_1707,N_1619);
or U1924 (N_1924,N_1772,N_1799);
nor U1925 (N_1925,N_1784,N_1790);
and U1926 (N_1926,N_1717,N_1630);
or U1927 (N_1927,N_1751,N_1780);
nand U1928 (N_1928,N_1692,N_1661);
xnor U1929 (N_1929,N_1605,N_1764);
or U1930 (N_1930,N_1776,N_1603);
or U1931 (N_1931,N_1636,N_1701);
or U1932 (N_1932,N_1760,N_1626);
and U1933 (N_1933,N_1786,N_1615);
nor U1934 (N_1934,N_1762,N_1751);
and U1935 (N_1935,N_1634,N_1767);
and U1936 (N_1936,N_1767,N_1780);
and U1937 (N_1937,N_1632,N_1705);
nor U1938 (N_1938,N_1696,N_1629);
xor U1939 (N_1939,N_1606,N_1798);
and U1940 (N_1940,N_1760,N_1624);
nor U1941 (N_1941,N_1745,N_1777);
nor U1942 (N_1942,N_1727,N_1772);
xnor U1943 (N_1943,N_1626,N_1600);
xor U1944 (N_1944,N_1610,N_1678);
xor U1945 (N_1945,N_1784,N_1613);
or U1946 (N_1946,N_1662,N_1652);
or U1947 (N_1947,N_1673,N_1670);
and U1948 (N_1948,N_1669,N_1762);
or U1949 (N_1949,N_1739,N_1706);
xor U1950 (N_1950,N_1648,N_1641);
nor U1951 (N_1951,N_1678,N_1750);
nor U1952 (N_1952,N_1627,N_1683);
nor U1953 (N_1953,N_1623,N_1775);
nand U1954 (N_1954,N_1781,N_1669);
nand U1955 (N_1955,N_1653,N_1685);
and U1956 (N_1956,N_1658,N_1781);
nand U1957 (N_1957,N_1781,N_1635);
nor U1958 (N_1958,N_1618,N_1736);
xor U1959 (N_1959,N_1699,N_1696);
nand U1960 (N_1960,N_1750,N_1645);
nor U1961 (N_1961,N_1721,N_1607);
nand U1962 (N_1962,N_1780,N_1688);
nand U1963 (N_1963,N_1744,N_1712);
nand U1964 (N_1964,N_1784,N_1665);
nand U1965 (N_1965,N_1688,N_1788);
nor U1966 (N_1966,N_1758,N_1679);
nand U1967 (N_1967,N_1722,N_1697);
nor U1968 (N_1968,N_1660,N_1637);
nor U1969 (N_1969,N_1691,N_1703);
or U1970 (N_1970,N_1616,N_1714);
nand U1971 (N_1971,N_1629,N_1687);
xor U1972 (N_1972,N_1785,N_1717);
and U1973 (N_1973,N_1728,N_1739);
nor U1974 (N_1974,N_1735,N_1673);
or U1975 (N_1975,N_1669,N_1699);
xor U1976 (N_1976,N_1643,N_1732);
or U1977 (N_1977,N_1762,N_1772);
nor U1978 (N_1978,N_1670,N_1622);
nor U1979 (N_1979,N_1627,N_1650);
xnor U1980 (N_1980,N_1620,N_1790);
nand U1981 (N_1981,N_1737,N_1661);
xor U1982 (N_1982,N_1694,N_1642);
and U1983 (N_1983,N_1683,N_1796);
nand U1984 (N_1984,N_1793,N_1771);
or U1985 (N_1985,N_1731,N_1687);
or U1986 (N_1986,N_1655,N_1727);
and U1987 (N_1987,N_1687,N_1722);
or U1988 (N_1988,N_1759,N_1621);
or U1989 (N_1989,N_1792,N_1677);
and U1990 (N_1990,N_1734,N_1724);
xnor U1991 (N_1991,N_1640,N_1777);
nand U1992 (N_1992,N_1635,N_1796);
and U1993 (N_1993,N_1792,N_1631);
or U1994 (N_1994,N_1673,N_1719);
or U1995 (N_1995,N_1725,N_1765);
nor U1996 (N_1996,N_1793,N_1679);
or U1997 (N_1997,N_1633,N_1613);
xor U1998 (N_1998,N_1769,N_1701);
and U1999 (N_1999,N_1759,N_1779);
xnor U2000 (N_2000,N_1966,N_1898);
xor U2001 (N_2001,N_1955,N_1837);
nor U2002 (N_2002,N_1801,N_1877);
nand U2003 (N_2003,N_1927,N_1817);
and U2004 (N_2004,N_1942,N_1983);
and U2005 (N_2005,N_1826,N_1916);
nor U2006 (N_2006,N_1890,N_1883);
xnor U2007 (N_2007,N_1959,N_1870);
xor U2008 (N_2008,N_1882,N_1943);
nor U2009 (N_2009,N_1881,N_1841);
nor U2010 (N_2010,N_1824,N_1972);
nand U2011 (N_2011,N_1819,N_1969);
or U2012 (N_2012,N_1807,N_1874);
nor U2013 (N_2013,N_1957,N_1923);
xor U2014 (N_2014,N_1976,N_1834);
nand U2015 (N_2015,N_1995,N_1932);
or U2016 (N_2016,N_1853,N_1956);
and U2017 (N_2017,N_1864,N_1922);
or U2018 (N_2018,N_1852,N_1888);
or U2019 (N_2019,N_1988,N_1831);
nor U2020 (N_2020,N_1871,N_1989);
xnor U2021 (N_2021,N_1945,N_1896);
xor U2022 (N_2022,N_1921,N_1810);
xor U2023 (N_2023,N_1893,N_1805);
or U2024 (N_2024,N_1996,N_1986);
and U2025 (N_2025,N_1891,N_1939);
nand U2026 (N_2026,N_1878,N_1948);
nand U2027 (N_2027,N_1961,N_1894);
or U2028 (N_2028,N_1900,N_1967);
or U2029 (N_2029,N_1830,N_1999);
nand U2030 (N_2030,N_1971,N_1901);
nand U2031 (N_2031,N_1938,N_1910);
or U2032 (N_2032,N_1854,N_1886);
and U2033 (N_2033,N_1968,N_1985);
nand U2034 (N_2034,N_1859,N_1998);
xor U2035 (N_2035,N_1994,N_1940);
xor U2036 (N_2036,N_1931,N_1880);
xor U2037 (N_2037,N_1827,N_1873);
or U2038 (N_2038,N_1918,N_1821);
xor U2039 (N_2039,N_1876,N_1885);
nand U2040 (N_2040,N_1860,N_1964);
nor U2041 (N_2041,N_1899,N_1815);
or U2042 (N_2042,N_1872,N_1867);
nor U2043 (N_2043,N_1944,N_1935);
and U2044 (N_2044,N_1869,N_1808);
xnor U2045 (N_2045,N_1908,N_1823);
xnor U2046 (N_2046,N_1802,N_1952);
and U2047 (N_2047,N_1844,N_1920);
or U2048 (N_2048,N_1915,N_1855);
xor U2049 (N_2049,N_1958,N_1829);
nand U2050 (N_2050,N_1811,N_1847);
and U2051 (N_2051,N_1982,N_1946);
and U2052 (N_2052,N_1937,N_1849);
xnor U2053 (N_2053,N_1993,N_1947);
nand U2054 (N_2054,N_1858,N_1840);
and U2055 (N_2055,N_1909,N_1991);
and U2056 (N_2056,N_1990,N_1806);
and U2057 (N_2057,N_1965,N_1984);
xor U2058 (N_2058,N_1816,N_1933);
xor U2059 (N_2059,N_1820,N_1832);
nand U2060 (N_2060,N_1875,N_1842);
xnor U2061 (N_2061,N_1892,N_1809);
nand U2062 (N_2062,N_1925,N_1828);
or U2063 (N_2063,N_1917,N_1904);
and U2064 (N_2064,N_1838,N_1907);
nor U2065 (N_2065,N_1897,N_1836);
nor U2066 (N_2066,N_1903,N_1953);
xor U2067 (N_2067,N_1936,N_1863);
nand U2068 (N_2068,N_1887,N_1963);
and U2069 (N_2069,N_1919,N_1868);
or U2070 (N_2070,N_1914,N_1997);
or U2071 (N_2071,N_1839,N_1911);
nor U2072 (N_2072,N_1889,N_1848);
and U2073 (N_2073,N_1979,N_1913);
nor U2074 (N_2074,N_1950,N_1818);
nor U2075 (N_2075,N_1866,N_1962);
nand U2076 (N_2076,N_1906,N_1929);
and U2077 (N_2077,N_1865,N_1974);
and U2078 (N_2078,N_1924,N_1930);
and U2079 (N_2079,N_1845,N_1992);
or U2080 (N_2080,N_1949,N_1813);
and U2081 (N_2081,N_1934,N_1912);
or U2082 (N_2082,N_1835,N_1987);
and U2083 (N_2083,N_1941,N_1825);
or U2084 (N_2084,N_1977,N_1861);
or U2085 (N_2085,N_1926,N_1954);
or U2086 (N_2086,N_1975,N_1857);
nand U2087 (N_2087,N_1851,N_1856);
or U2088 (N_2088,N_1928,N_1804);
or U2089 (N_2089,N_1951,N_1905);
or U2090 (N_2090,N_1973,N_1862);
xor U2091 (N_2091,N_1850,N_1814);
xnor U2092 (N_2092,N_1833,N_1803);
nor U2093 (N_2093,N_1846,N_1902);
xor U2094 (N_2094,N_1822,N_1800);
nor U2095 (N_2095,N_1981,N_1884);
xor U2096 (N_2096,N_1978,N_1895);
nor U2097 (N_2097,N_1970,N_1879);
or U2098 (N_2098,N_1812,N_1960);
nor U2099 (N_2099,N_1843,N_1980);
xor U2100 (N_2100,N_1889,N_1815);
nor U2101 (N_2101,N_1843,N_1887);
nor U2102 (N_2102,N_1924,N_1980);
and U2103 (N_2103,N_1918,N_1872);
and U2104 (N_2104,N_1914,N_1934);
nor U2105 (N_2105,N_1973,N_1879);
and U2106 (N_2106,N_1826,N_1928);
or U2107 (N_2107,N_1856,N_1824);
or U2108 (N_2108,N_1971,N_1899);
or U2109 (N_2109,N_1997,N_1985);
or U2110 (N_2110,N_1913,N_1877);
and U2111 (N_2111,N_1884,N_1831);
nor U2112 (N_2112,N_1812,N_1808);
nor U2113 (N_2113,N_1863,N_1861);
and U2114 (N_2114,N_1940,N_1866);
and U2115 (N_2115,N_1991,N_1949);
nor U2116 (N_2116,N_1872,N_1943);
or U2117 (N_2117,N_1807,N_1868);
xor U2118 (N_2118,N_1912,N_1873);
and U2119 (N_2119,N_1975,N_1881);
nor U2120 (N_2120,N_1893,N_1867);
nand U2121 (N_2121,N_1838,N_1911);
nor U2122 (N_2122,N_1996,N_1943);
or U2123 (N_2123,N_1971,N_1879);
and U2124 (N_2124,N_1942,N_1949);
or U2125 (N_2125,N_1940,N_1843);
nand U2126 (N_2126,N_1886,N_1925);
nor U2127 (N_2127,N_1856,N_1933);
and U2128 (N_2128,N_1930,N_1904);
nand U2129 (N_2129,N_1936,N_1966);
nor U2130 (N_2130,N_1868,N_1929);
and U2131 (N_2131,N_1997,N_1890);
nor U2132 (N_2132,N_1845,N_1977);
nand U2133 (N_2133,N_1928,N_1817);
nand U2134 (N_2134,N_1957,N_1839);
or U2135 (N_2135,N_1803,N_1955);
and U2136 (N_2136,N_1987,N_1817);
xor U2137 (N_2137,N_1925,N_1834);
and U2138 (N_2138,N_1968,N_1961);
xor U2139 (N_2139,N_1814,N_1832);
nor U2140 (N_2140,N_1984,N_1843);
and U2141 (N_2141,N_1995,N_1800);
or U2142 (N_2142,N_1963,N_1894);
nor U2143 (N_2143,N_1898,N_1959);
nand U2144 (N_2144,N_1839,N_1858);
xnor U2145 (N_2145,N_1917,N_1994);
nor U2146 (N_2146,N_1927,N_1995);
xnor U2147 (N_2147,N_1865,N_1816);
nand U2148 (N_2148,N_1909,N_1895);
nor U2149 (N_2149,N_1866,N_1972);
nor U2150 (N_2150,N_1942,N_1961);
or U2151 (N_2151,N_1873,N_1869);
xnor U2152 (N_2152,N_1825,N_1893);
xnor U2153 (N_2153,N_1983,N_1809);
nand U2154 (N_2154,N_1927,N_1804);
and U2155 (N_2155,N_1937,N_1978);
nor U2156 (N_2156,N_1950,N_1899);
nand U2157 (N_2157,N_1941,N_1986);
nor U2158 (N_2158,N_1951,N_1898);
nand U2159 (N_2159,N_1962,N_1842);
nor U2160 (N_2160,N_1880,N_1866);
xnor U2161 (N_2161,N_1909,N_1815);
nor U2162 (N_2162,N_1912,N_1981);
or U2163 (N_2163,N_1913,N_1885);
or U2164 (N_2164,N_1888,N_1960);
xor U2165 (N_2165,N_1840,N_1968);
nand U2166 (N_2166,N_1958,N_1811);
or U2167 (N_2167,N_1840,N_1833);
nand U2168 (N_2168,N_1894,N_1863);
and U2169 (N_2169,N_1973,N_1920);
and U2170 (N_2170,N_1912,N_1922);
or U2171 (N_2171,N_1809,N_1844);
or U2172 (N_2172,N_1801,N_1906);
nand U2173 (N_2173,N_1820,N_1851);
xnor U2174 (N_2174,N_1902,N_1933);
nor U2175 (N_2175,N_1987,N_1869);
nand U2176 (N_2176,N_1935,N_1968);
xnor U2177 (N_2177,N_1901,N_1801);
xnor U2178 (N_2178,N_1972,N_1956);
xor U2179 (N_2179,N_1983,N_1893);
and U2180 (N_2180,N_1804,N_1831);
and U2181 (N_2181,N_1979,N_1834);
xnor U2182 (N_2182,N_1804,N_1955);
nor U2183 (N_2183,N_1971,N_1832);
and U2184 (N_2184,N_1918,N_1804);
or U2185 (N_2185,N_1893,N_1883);
and U2186 (N_2186,N_1900,N_1809);
and U2187 (N_2187,N_1950,N_1892);
nand U2188 (N_2188,N_1946,N_1898);
xor U2189 (N_2189,N_1912,N_1853);
xor U2190 (N_2190,N_1830,N_1955);
xor U2191 (N_2191,N_1902,N_1897);
nor U2192 (N_2192,N_1857,N_1996);
nor U2193 (N_2193,N_1974,N_1940);
nand U2194 (N_2194,N_1940,N_1833);
and U2195 (N_2195,N_1900,N_1810);
nand U2196 (N_2196,N_1970,N_1962);
xnor U2197 (N_2197,N_1897,N_1888);
or U2198 (N_2198,N_1853,N_1967);
nor U2199 (N_2199,N_1816,N_1959);
nand U2200 (N_2200,N_2142,N_2084);
nor U2201 (N_2201,N_2125,N_2199);
xor U2202 (N_2202,N_2088,N_2175);
or U2203 (N_2203,N_2153,N_2192);
nand U2204 (N_2204,N_2182,N_2021);
or U2205 (N_2205,N_2118,N_2188);
or U2206 (N_2206,N_2092,N_2059);
xnor U2207 (N_2207,N_2096,N_2179);
nor U2208 (N_2208,N_2020,N_2141);
xor U2209 (N_2209,N_2019,N_2060);
nor U2210 (N_2210,N_2053,N_2002);
and U2211 (N_2211,N_2154,N_2195);
nor U2212 (N_2212,N_2176,N_2052);
and U2213 (N_2213,N_2189,N_2036);
nor U2214 (N_2214,N_2187,N_2127);
nand U2215 (N_2215,N_2039,N_2105);
nand U2216 (N_2216,N_2093,N_2177);
nand U2217 (N_2217,N_2198,N_2013);
nor U2218 (N_2218,N_2112,N_2110);
xnor U2219 (N_2219,N_2076,N_2196);
and U2220 (N_2220,N_2180,N_2178);
or U2221 (N_2221,N_2169,N_2184);
and U2222 (N_2222,N_2094,N_2151);
xnor U2223 (N_2223,N_2121,N_2126);
nand U2224 (N_2224,N_2145,N_2140);
or U2225 (N_2225,N_2161,N_2097);
and U2226 (N_2226,N_2069,N_2029);
nor U2227 (N_2227,N_2087,N_2086);
nand U2228 (N_2228,N_2120,N_2091);
nand U2229 (N_2229,N_2168,N_2030);
and U2230 (N_2230,N_2155,N_2048);
nor U2231 (N_2231,N_2071,N_2134);
nand U2232 (N_2232,N_2018,N_2009);
nand U2233 (N_2233,N_2162,N_2133);
nand U2234 (N_2234,N_2051,N_2016);
nor U2235 (N_2235,N_2173,N_2164);
or U2236 (N_2236,N_2003,N_2080);
nor U2237 (N_2237,N_2111,N_2124);
nand U2238 (N_2238,N_2077,N_2174);
or U2239 (N_2239,N_2171,N_2011);
xnor U2240 (N_2240,N_2165,N_2072);
nor U2241 (N_2241,N_2146,N_2131);
and U2242 (N_2242,N_2108,N_2063);
nand U2243 (N_2243,N_2099,N_2159);
or U2244 (N_2244,N_2135,N_2115);
or U2245 (N_2245,N_2117,N_2104);
or U2246 (N_2246,N_2148,N_2101);
and U2247 (N_2247,N_2033,N_2103);
nor U2248 (N_2248,N_2089,N_2050);
or U2249 (N_2249,N_2194,N_2172);
xnor U2250 (N_2250,N_2058,N_2000);
and U2251 (N_2251,N_2037,N_2090);
and U2252 (N_2252,N_2047,N_2098);
and U2253 (N_2253,N_2191,N_2081);
or U2254 (N_2254,N_2137,N_2042);
nand U2255 (N_2255,N_2001,N_2054);
or U2256 (N_2256,N_2008,N_2005);
or U2257 (N_2257,N_2139,N_2044);
nor U2258 (N_2258,N_2181,N_2073);
nor U2259 (N_2259,N_2034,N_2113);
nand U2260 (N_2260,N_2065,N_2147);
or U2261 (N_2261,N_2022,N_2074);
nor U2262 (N_2262,N_2095,N_2043);
xnor U2263 (N_2263,N_2106,N_2109);
xnor U2264 (N_2264,N_2157,N_2079);
and U2265 (N_2265,N_2032,N_2057);
nand U2266 (N_2266,N_2055,N_2129);
nor U2267 (N_2267,N_2144,N_2170);
nor U2268 (N_2268,N_2028,N_2025);
and U2269 (N_2269,N_2152,N_2010);
nand U2270 (N_2270,N_2130,N_2017);
nor U2271 (N_2271,N_2070,N_2035);
xor U2272 (N_2272,N_2007,N_2041);
and U2273 (N_2273,N_2061,N_2160);
nand U2274 (N_2274,N_2085,N_2128);
nand U2275 (N_2275,N_2186,N_2049);
nand U2276 (N_2276,N_2012,N_2083);
nor U2277 (N_2277,N_2067,N_2107);
nand U2278 (N_2278,N_2102,N_2167);
nand U2279 (N_2279,N_2014,N_2190);
nor U2280 (N_2280,N_2143,N_2062);
nand U2281 (N_2281,N_2064,N_2166);
nor U2282 (N_2282,N_2075,N_2056);
xnor U2283 (N_2283,N_2046,N_2119);
nand U2284 (N_2284,N_2027,N_2138);
xnor U2285 (N_2285,N_2132,N_2163);
nor U2286 (N_2286,N_2100,N_2038);
nand U2287 (N_2287,N_2122,N_2183);
and U2288 (N_2288,N_2031,N_2004);
or U2289 (N_2289,N_2082,N_2078);
or U2290 (N_2290,N_2068,N_2040);
nor U2291 (N_2291,N_2193,N_2149);
and U2292 (N_2292,N_2136,N_2023);
nand U2293 (N_2293,N_2024,N_2114);
or U2294 (N_2294,N_2156,N_2015);
nor U2295 (N_2295,N_2006,N_2158);
xor U2296 (N_2296,N_2116,N_2123);
nand U2297 (N_2297,N_2045,N_2150);
nand U2298 (N_2298,N_2066,N_2197);
and U2299 (N_2299,N_2185,N_2026);
nor U2300 (N_2300,N_2043,N_2197);
or U2301 (N_2301,N_2051,N_2118);
nand U2302 (N_2302,N_2025,N_2062);
nand U2303 (N_2303,N_2199,N_2084);
and U2304 (N_2304,N_2146,N_2014);
and U2305 (N_2305,N_2037,N_2074);
and U2306 (N_2306,N_2039,N_2025);
nand U2307 (N_2307,N_2077,N_2090);
and U2308 (N_2308,N_2128,N_2019);
or U2309 (N_2309,N_2125,N_2107);
or U2310 (N_2310,N_2053,N_2178);
xor U2311 (N_2311,N_2010,N_2029);
nand U2312 (N_2312,N_2160,N_2065);
nor U2313 (N_2313,N_2134,N_2124);
xor U2314 (N_2314,N_2101,N_2120);
nand U2315 (N_2315,N_2093,N_2001);
xnor U2316 (N_2316,N_2138,N_2131);
nor U2317 (N_2317,N_2088,N_2014);
xnor U2318 (N_2318,N_2031,N_2043);
or U2319 (N_2319,N_2065,N_2078);
nand U2320 (N_2320,N_2149,N_2195);
and U2321 (N_2321,N_2122,N_2046);
nand U2322 (N_2322,N_2157,N_2127);
nand U2323 (N_2323,N_2130,N_2054);
nand U2324 (N_2324,N_2055,N_2095);
nand U2325 (N_2325,N_2049,N_2040);
and U2326 (N_2326,N_2026,N_2094);
nand U2327 (N_2327,N_2181,N_2131);
xnor U2328 (N_2328,N_2033,N_2026);
nor U2329 (N_2329,N_2010,N_2047);
xor U2330 (N_2330,N_2038,N_2173);
nand U2331 (N_2331,N_2062,N_2133);
or U2332 (N_2332,N_2010,N_2040);
nor U2333 (N_2333,N_2073,N_2018);
nor U2334 (N_2334,N_2014,N_2041);
nand U2335 (N_2335,N_2035,N_2031);
nand U2336 (N_2336,N_2097,N_2098);
xor U2337 (N_2337,N_2166,N_2164);
xor U2338 (N_2338,N_2053,N_2145);
and U2339 (N_2339,N_2047,N_2151);
and U2340 (N_2340,N_2110,N_2188);
nor U2341 (N_2341,N_2056,N_2135);
nor U2342 (N_2342,N_2056,N_2039);
xnor U2343 (N_2343,N_2159,N_2050);
nand U2344 (N_2344,N_2005,N_2186);
nor U2345 (N_2345,N_2009,N_2080);
nor U2346 (N_2346,N_2066,N_2102);
nand U2347 (N_2347,N_2181,N_2090);
and U2348 (N_2348,N_2051,N_2093);
or U2349 (N_2349,N_2193,N_2185);
and U2350 (N_2350,N_2007,N_2144);
or U2351 (N_2351,N_2051,N_2019);
nor U2352 (N_2352,N_2110,N_2063);
and U2353 (N_2353,N_2048,N_2077);
and U2354 (N_2354,N_2035,N_2186);
or U2355 (N_2355,N_2160,N_2018);
or U2356 (N_2356,N_2047,N_2196);
xor U2357 (N_2357,N_2058,N_2137);
and U2358 (N_2358,N_2061,N_2198);
or U2359 (N_2359,N_2003,N_2016);
xor U2360 (N_2360,N_2166,N_2102);
nor U2361 (N_2361,N_2018,N_2196);
nand U2362 (N_2362,N_2113,N_2187);
nor U2363 (N_2363,N_2116,N_2128);
nor U2364 (N_2364,N_2062,N_2049);
xor U2365 (N_2365,N_2139,N_2023);
or U2366 (N_2366,N_2003,N_2151);
and U2367 (N_2367,N_2021,N_2018);
nand U2368 (N_2368,N_2099,N_2145);
and U2369 (N_2369,N_2115,N_2143);
nor U2370 (N_2370,N_2016,N_2001);
nand U2371 (N_2371,N_2171,N_2105);
and U2372 (N_2372,N_2068,N_2039);
xor U2373 (N_2373,N_2061,N_2105);
and U2374 (N_2374,N_2192,N_2068);
nor U2375 (N_2375,N_2031,N_2166);
nand U2376 (N_2376,N_2036,N_2169);
or U2377 (N_2377,N_2076,N_2030);
nor U2378 (N_2378,N_2094,N_2010);
nand U2379 (N_2379,N_2009,N_2116);
or U2380 (N_2380,N_2171,N_2119);
nor U2381 (N_2381,N_2075,N_2008);
xnor U2382 (N_2382,N_2004,N_2198);
nand U2383 (N_2383,N_2173,N_2069);
or U2384 (N_2384,N_2162,N_2032);
and U2385 (N_2385,N_2000,N_2022);
nand U2386 (N_2386,N_2009,N_2193);
nor U2387 (N_2387,N_2193,N_2097);
and U2388 (N_2388,N_2187,N_2142);
nand U2389 (N_2389,N_2019,N_2132);
xor U2390 (N_2390,N_2108,N_2189);
nor U2391 (N_2391,N_2060,N_2166);
xor U2392 (N_2392,N_2143,N_2155);
nand U2393 (N_2393,N_2126,N_2034);
xor U2394 (N_2394,N_2020,N_2114);
nor U2395 (N_2395,N_2026,N_2123);
or U2396 (N_2396,N_2197,N_2048);
or U2397 (N_2397,N_2053,N_2194);
nor U2398 (N_2398,N_2058,N_2024);
xor U2399 (N_2399,N_2132,N_2117);
and U2400 (N_2400,N_2372,N_2283);
nand U2401 (N_2401,N_2257,N_2232);
or U2402 (N_2402,N_2324,N_2218);
nand U2403 (N_2403,N_2304,N_2291);
nor U2404 (N_2404,N_2332,N_2252);
nand U2405 (N_2405,N_2245,N_2254);
nor U2406 (N_2406,N_2351,N_2345);
xor U2407 (N_2407,N_2303,N_2357);
or U2408 (N_2408,N_2287,N_2322);
xor U2409 (N_2409,N_2361,N_2217);
or U2410 (N_2410,N_2233,N_2374);
xor U2411 (N_2411,N_2383,N_2275);
xor U2412 (N_2412,N_2373,N_2337);
nor U2413 (N_2413,N_2328,N_2201);
or U2414 (N_2414,N_2312,N_2350);
nor U2415 (N_2415,N_2323,N_2240);
xor U2416 (N_2416,N_2215,N_2264);
nand U2417 (N_2417,N_2256,N_2247);
xor U2418 (N_2418,N_2359,N_2307);
xnor U2419 (N_2419,N_2296,N_2284);
nand U2420 (N_2420,N_2259,N_2338);
and U2421 (N_2421,N_2297,N_2318);
xnor U2422 (N_2422,N_2321,N_2330);
or U2423 (N_2423,N_2334,N_2368);
or U2424 (N_2424,N_2279,N_2238);
xnor U2425 (N_2425,N_2389,N_2265);
nor U2426 (N_2426,N_2269,N_2305);
or U2427 (N_2427,N_2392,N_2298);
xnor U2428 (N_2428,N_2280,N_2276);
or U2429 (N_2429,N_2335,N_2277);
xor U2430 (N_2430,N_2382,N_2289);
xor U2431 (N_2431,N_2258,N_2213);
nand U2432 (N_2432,N_2248,N_2320);
nor U2433 (N_2433,N_2266,N_2356);
nor U2434 (N_2434,N_2250,N_2358);
or U2435 (N_2435,N_2292,N_2390);
xor U2436 (N_2436,N_2365,N_2377);
nand U2437 (N_2437,N_2237,N_2319);
xor U2438 (N_2438,N_2347,N_2263);
and U2439 (N_2439,N_2231,N_2262);
nand U2440 (N_2440,N_2226,N_2288);
or U2441 (N_2441,N_2253,N_2200);
nor U2442 (N_2442,N_2222,N_2267);
and U2443 (N_2443,N_2209,N_2230);
and U2444 (N_2444,N_2384,N_2235);
xor U2445 (N_2445,N_2327,N_2386);
nand U2446 (N_2446,N_2281,N_2329);
xor U2447 (N_2447,N_2221,N_2299);
nor U2448 (N_2448,N_2220,N_2225);
or U2449 (N_2449,N_2336,N_2313);
xnor U2450 (N_2450,N_2348,N_2204);
or U2451 (N_2451,N_2355,N_2344);
and U2452 (N_2452,N_2380,N_2360);
xor U2453 (N_2453,N_2272,N_2239);
or U2454 (N_2454,N_2223,N_2371);
nor U2455 (N_2455,N_2286,N_2273);
and U2456 (N_2456,N_2210,N_2228);
and U2457 (N_2457,N_2227,N_2364);
nor U2458 (N_2458,N_2376,N_2243);
and U2459 (N_2459,N_2278,N_2354);
or U2460 (N_2460,N_2310,N_2308);
and U2461 (N_2461,N_2293,N_2362);
xnor U2462 (N_2462,N_2268,N_2388);
and U2463 (N_2463,N_2366,N_2378);
xnor U2464 (N_2464,N_2370,N_2341);
xor U2465 (N_2465,N_2326,N_2241);
and U2466 (N_2466,N_2381,N_2219);
nand U2467 (N_2467,N_2260,N_2346);
xor U2468 (N_2468,N_2314,N_2242);
or U2469 (N_2469,N_2340,N_2391);
nor U2470 (N_2470,N_2317,N_2397);
and U2471 (N_2471,N_2385,N_2309);
nor U2472 (N_2472,N_2271,N_2244);
or U2473 (N_2473,N_2290,N_2379);
or U2474 (N_2474,N_2349,N_2207);
and U2475 (N_2475,N_2369,N_2301);
xor U2476 (N_2476,N_2203,N_2224);
or U2477 (N_2477,N_2333,N_2343);
or U2478 (N_2478,N_2270,N_2261);
xor U2479 (N_2479,N_2315,N_2229);
or U2480 (N_2480,N_2387,N_2367);
or U2481 (N_2481,N_2234,N_2285);
nand U2482 (N_2482,N_2255,N_2208);
nor U2483 (N_2483,N_2294,N_2339);
and U2484 (N_2484,N_2325,N_2306);
or U2485 (N_2485,N_2398,N_2399);
nand U2486 (N_2486,N_2300,N_2311);
and U2487 (N_2487,N_2214,N_2251);
and U2488 (N_2488,N_2202,N_2212);
and U2489 (N_2489,N_2274,N_2375);
xor U2490 (N_2490,N_2302,N_2394);
nand U2491 (N_2491,N_2205,N_2246);
or U2492 (N_2492,N_2206,N_2216);
xor U2493 (N_2493,N_2393,N_2352);
xnor U2494 (N_2494,N_2316,N_2396);
nor U2495 (N_2495,N_2211,N_2249);
or U2496 (N_2496,N_2236,N_2295);
xor U2497 (N_2497,N_2331,N_2282);
and U2498 (N_2498,N_2353,N_2342);
and U2499 (N_2499,N_2395,N_2363);
xor U2500 (N_2500,N_2361,N_2290);
or U2501 (N_2501,N_2376,N_2251);
and U2502 (N_2502,N_2203,N_2286);
xor U2503 (N_2503,N_2332,N_2202);
or U2504 (N_2504,N_2340,N_2250);
nand U2505 (N_2505,N_2339,N_2340);
nand U2506 (N_2506,N_2272,N_2385);
nor U2507 (N_2507,N_2371,N_2369);
xor U2508 (N_2508,N_2383,N_2273);
nand U2509 (N_2509,N_2240,N_2330);
or U2510 (N_2510,N_2392,N_2398);
and U2511 (N_2511,N_2336,N_2398);
nand U2512 (N_2512,N_2327,N_2270);
nand U2513 (N_2513,N_2380,N_2285);
nand U2514 (N_2514,N_2307,N_2218);
xor U2515 (N_2515,N_2332,N_2327);
nor U2516 (N_2516,N_2335,N_2302);
xor U2517 (N_2517,N_2346,N_2216);
and U2518 (N_2518,N_2310,N_2275);
nor U2519 (N_2519,N_2279,N_2340);
and U2520 (N_2520,N_2289,N_2237);
or U2521 (N_2521,N_2277,N_2258);
nor U2522 (N_2522,N_2212,N_2316);
xor U2523 (N_2523,N_2208,N_2215);
or U2524 (N_2524,N_2284,N_2323);
and U2525 (N_2525,N_2281,N_2261);
nand U2526 (N_2526,N_2376,N_2255);
xnor U2527 (N_2527,N_2312,N_2217);
nand U2528 (N_2528,N_2235,N_2336);
or U2529 (N_2529,N_2373,N_2361);
nor U2530 (N_2530,N_2234,N_2395);
nand U2531 (N_2531,N_2390,N_2231);
and U2532 (N_2532,N_2254,N_2232);
nand U2533 (N_2533,N_2221,N_2219);
and U2534 (N_2534,N_2383,N_2336);
and U2535 (N_2535,N_2340,N_2294);
nor U2536 (N_2536,N_2366,N_2357);
xor U2537 (N_2537,N_2332,N_2296);
and U2538 (N_2538,N_2274,N_2337);
xor U2539 (N_2539,N_2263,N_2310);
nor U2540 (N_2540,N_2269,N_2322);
and U2541 (N_2541,N_2276,N_2343);
nor U2542 (N_2542,N_2317,N_2324);
or U2543 (N_2543,N_2319,N_2245);
nand U2544 (N_2544,N_2294,N_2259);
nor U2545 (N_2545,N_2261,N_2311);
or U2546 (N_2546,N_2280,N_2318);
xnor U2547 (N_2547,N_2304,N_2228);
and U2548 (N_2548,N_2380,N_2231);
or U2549 (N_2549,N_2276,N_2275);
nand U2550 (N_2550,N_2381,N_2352);
nand U2551 (N_2551,N_2315,N_2305);
xor U2552 (N_2552,N_2328,N_2309);
or U2553 (N_2553,N_2269,N_2318);
or U2554 (N_2554,N_2218,N_2211);
nand U2555 (N_2555,N_2255,N_2284);
xor U2556 (N_2556,N_2226,N_2308);
or U2557 (N_2557,N_2336,N_2244);
and U2558 (N_2558,N_2388,N_2395);
and U2559 (N_2559,N_2287,N_2221);
nand U2560 (N_2560,N_2326,N_2316);
nor U2561 (N_2561,N_2278,N_2216);
and U2562 (N_2562,N_2367,N_2285);
nand U2563 (N_2563,N_2202,N_2284);
and U2564 (N_2564,N_2365,N_2280);
nand U2565 (N_2565,N_2231,N_2289);
and U2566 (N_2566,N_2255,N_2270);
or U2567 (N_2567,N_2315,N_2216);
or U2568 (N_2568,N_2226,N_2266);
nand U2569 (N_2569,N_2316,N_2204);
nand U2570 (N_2570,N_2361,N_2332);
or U2571 (N_2571,N_2279,N_2312);
nand U2572 (N_2572,N_2381,N_2241);
or U2573 (N_2573,N_2348,N_2279);
nand U2574 (N_2574,N_2264,N_2383);
nor U2575 (N_2575,N_2346,N_2337);
or U2576 (N_2576,N_2218,N_2317);
nor U2577 (N_2577,N_2367,N_2360);
nand U2578 (N_2578,N_2374,N_2280);
or U2579 (N_2579,N_2389,N_2379);
and U2580 (N_2580,N_2368,N_2312);
nor U2581 (N_2581,N_2303,N_2332);
and U2582 (N_2582,N_2391,N_2275);
nor U2583 (N_2583,N_2341,N_2358);
and U2584 (N_2584,N_2219,N_2276);
and U2585 (N_2585,N_2385,N_2297);
nor U2586 (N_2586,N_2263,N_2241);
xor U2587 (N_2587,N_2259,N_2237);
xnor U2588 (N_2588,N_2246,N_2376);
and U2589 (N_2589,N_2377,N_2242);
nand U2590 (N_2590,N_2261,N_2374);
nor U2591 (N_2591,N_2396,N_2326);
nor U2592 (N_2592,N_2268,N_2314);
xnor U2593 (N_2593,N_2231,N_2265);
or U2594 (N_2594,N_2345,N_2260);
nor U2595 (N_2595,N_2357,N_2311);
nor U2596 (N_2596,N_2343,N_2271);
or U2597 (N_2597,N_2322,N_2271);
or U2598 (N_2598,N_2396,N_2240);
nor U2599 (N_2599,N_2282,N_2233);
or U2600 (N_2600,N_2404,N_2556);
nand U2601 (N_2601,N_2591,N_2417);
xor U2602 (N_2602,N_2592,N_2427);
xor U2603 (N_2603,N_2434,N_2489);
xor U2604 (N_2604,N_2523,N_2543);
nand U2605 (N_2605,N_2576,N_2415);
or U2606 (N_2606,N_2590,N_2581);
nand U2607 (N_2607,N_2534,N_2428);
or U2608 (N_2608,N_2446,N_2533);
and U2609 (N_2609,N_2472,N_2536);
xor U2610 (N_2610,N_2578,N_2517);
and U2611 (N_2611,N_2450,N_2488);
and U2612 (N_2612,N_2430,N_2412);
and U2613 (N_2613,N_2483,N_2587);
or U2614 (N_2614,N_2492,N_2570);
and U2615 (N_2615,N_2572,N_2518);
nor U2616 (N_2616,N_2573,N_2432);
and U2617 (N_2617,N_2422,N_2526);
nand U2618 (N_2618,N_2530,N_2553);
xnor U2619 (N_2619,N_2445,N_2456);
or U2620 (N_2620,N_2495,N_2452);
nor U2621 (N_2621,N_2504,N_2481);
nor U2622 (N_2622,N_2583,N_2527);
nand U2623 (N_2623,N_2574,N_2540);
nor U2624 (N_2624,N_2549,N_2569);
xnor U2625 (N_2625,N_2515,N_2568);
or U2626 (N_2626,N_2555,N_2490);
nand U2627 (N_2627,N_2496,N_2405);
or U2628 (N_2628,N_2463,N_2544);
nor U2629 (N_2629,N_2541,N_2494);
and U2630 (N_2630,N_2577,N_2409);
nor U2631 (N_2631,N_2594,N_2493);
nand U2632 (N_2632,N_2589,N_2411);
or U2633 (N_2633,N_2438,N_2532);
nand U2634 (N_2634,N_2431,N_2444);
or U2635 (N_2635,N_2459,N_2598);
and U2636 (N_2636,N_2552,N_2559);
or U2637 (N_2637,N_2485,N_2538);
nor U2638 (N_2638,N_2406,N_2439);
nand U2639 (N_2639,N_2479,N_2449);
nand U2640 (N_2640,N_2524,N_2462);
and U2641 (N_2641,N_2595,N_2521);
or U2642 (N_2642,N_2471,N_2451);
and U2643 (N_2643,N_2546,N_2447);
and U2644 (N_2644,N_2407,N_2565);
nor U2645 (N_2645,N_2586,N_2505);
nand U2646 (N_2646,N_2453,N_2441);
and U2647 (N_2647,N_2484,N_2539);
xor U2648 (N_2648,N_2564,N_2465);
or U2649 (N_2649,N_2502,N_2503);
nand U2650 (N_2650,N_2477,N_2535);
and U2651 (N_2651,N_2480,N_2514);
and U2652 (N_2652,N_2507,N_2542);
or U2653 (N_2653,N_2478,N_2562);
xnor U2654 (N_2654,N_2413,N_2470);
or U2655 (N_2655,N_2597,N_2424);
nand U2656 (N_2656,N_2443,N_2403);
nor U2657 (N_2657,N_2571,N_2436);
xor U2658 (N_2658,N_2473,N_2425);
xnor U2659 (N_2659,N_2554,N_2548);
xor U2660 (N_2660,N_2516,N_2464);
nand U2661 (N_2661,N_2593,N_2575);
or U2662 (N_2662,N_2545,N_2561);
nand U2663 (N_2663,N_2402,N_2497);
nor U2664 (N_2664,N_2501,N_2566);
xnor U2665 (N_2665,N_2525,N_2580);
xor U2666 (N_2666,N_2537,N_2423);
nand U2667 (N_2667,N_2418,N_2557);
and U2668 (N_2668,N_2420,N_2508);
or U2669 (N_2669,N_2476,N_2512);
and U2670 (N_2670,N_2466,N_2558);
nand U2671 (N_2671,N_2588,N_2500);
xnor U2672 (N_2672,N_2454,N_2416);
nand U2673 (N_2673,N_2421,N_2522);
nand U2674 (N_2674,N_2551,N_2408);
nand U2675 (N_2675,N_2457,N_2509);
xnor U2676 (N_2676,N_2458,N_2531);
or U2677 (N_2677,N_2429,N_2519);
xnor U2678 (N_2678,N_2499,N_2582);
xnor U2679 (N_2679,N_2414,N_2474);
or U2680 (N_2680,N_2491,N_2529);
nand U2681 (N_2681,N_2596,N_2498);
nor U2682 (N_2682,N_2560,N_2510);
nand U2683 (N_2683,N_2455,N_2460);
nor U2684 (N_2684,N_2435,N_2426);
xnor U2685 (N_2685,N_2442,N_2400);
or U2686 (N_2686,N_2482,N_2599);
xnor U2687 (N_2687,N_2528,N_2579);
nand U2688 (N_2688,N_2448,N_2401);
nor U2689 (N_2689,N_2475,N_2520);
nor U2690 (N_2690,N_2567,N_2467);
nor U2691 (N_2691,N_2468,N_2440);
and U2692 (N_2692,N_2513,N_2419);
and U2693 (N_2693,N_2511,N_2584);
or U2694 (N_2694,N_2437,N_2410);
nand U2695 (N_2695,N_2487,N_2461);
nand U2696 (N_2696,N_2585,N_2506);
nor U2697 (N_2697,N_2550,N_2469);
nand U2698 (N_2698,N_2433,N_2486);
and U2699 (N_2699,N_2547,N_2563);
and U2700 (N_2700,N_2479,N_2574);
and U2701 (N_2701,N_2507,N_2592);
and U2702 (N_2702,N_2575,N_2578);
or U2703 (N_2703,N_2451,N_2417);
xnor U2704 (N_2704,N_2462,N_2454);
nor U2705 (N_2705,N_2522,N_2544);
or U2706 (N_2706,N_2401,N_2582);
xnor U2707 (N_2707,N_2400,N_2464);
or U2708 (N_2708,N_2564,N_2405);
and U2709 (N_2709,N_2513,N_2541);
nor U2710 (N_2710,N_2406,N_2404);
and U2711 (N_2711,N_2532,N_2452);
and U2712 (N_2712,N_2417,N_2572);
or U2713 (N_2713,N_2507,N_2531);
xor U2714 (N_2714,N_2578,N_2456);
or U2715 (N_2715,N_2509,N_2513);
nand U2716 (N_2716,N_2487,N_2495);
or U2717 (N_2717,N_2471,N_2586);
and U2718 (N_2718,N_2557,N_2422);
xor U2719 (N_2719,N_2594,N_2510);
or U2720 (N_2720,N_2515,N_2487);
or U2721 (N_2721,N_2547,N_2594);
nor U2722 (N_2722,N_2444,N_2497);
xor U2723 (N_2723,N_2506,N_2467);
and U2724 (N_2724,N_2470,N_2458);
xnor U2725 (N_2725,N_2430,N_2556);
and U2726 (N_2726,N_2476,N_2556);
nand U2727 (N_2727,N_2583,N_2417);
nand U2728 (N_2728,N_2594,N_2436);
nand U2729 (N_2729,N_2413,N_2593);
or U2730 (N_2730,N_2416,N_2571);
nand U2731 (N_2731,N_2590,N_2550);
nor U2732 (N_2732,N_2465,N_2591);
and U2733 (N_2733,N_2409,N_2418);
nor U2734 (N_2734,N_2459,N_2405);
nand U2735 (N_2735,N_2409,N_2448);
and U2736 (N_2736,N_2421,N_2537);
nor U2737 (N_2737,N_2433,N_2461);
or U2738 (N_2738,N_2445,N_2585);
nand U2739 (N_2739,N_2409,N_2506);
xor U2740 (N_2740,N_2409,N_2530);
nand U2741 (N_2741,N_2537,N_2592);
xor U2742 (N_2742,N_2469,N_2473);
nor U2743 (N_2743,N_2447,N_2418);
or U2744 (N_2744,N_2575,N_2508);
xor U2745 (N_2745,N_2503,N_2532);
nor U2746 (N_2746,N_2439,N_2433);
and U2747 (N_2747,N_2554,N_2427);
xor U2748 (N_2748,N_2445,N_2407);
xnor U2749 (N_2749,N_2459,N_2506);
nor U2750 (N_2750,N_2595,N_2490);
nand U2751 (N_2751,N_2430,N_2433);
and U2752 (N_2752,N_2489,N_2450);
or U2753 (N_2753,N_2511,N_2428);
xor U2754 (N_2754,N_2482,N_2506);
and U2755 (N_2755,N_2583,N_2462);
and U2756 (N_2756,N_2449,N_2551);
and U2757 (N_2757,N_2547,N_2517);
and U2758 (N_2758,N_2455,N_2433);
nor U2759 (N_2759,N_2573,N_2587);
and U2760 (N_2760,N_2593,N_2584);
or U2761 (N_2761,N_2416,N_2536);
nor U2762 (N_2762,N_2464,N_2413);
nand U2763 (N_2763,N_2402,N_2447);
nor U2764 (N_2764,N_2474,N_2464);
nand U2765 (N_2765,N_2531,N_2461);
and U2766 (N_2766,N_2453,N_2508);
nand U2767 (N_2767,N_2572,N_2567);
or U2768 (N_2768,N_2480,N_2512);
nor U2769 (N_2769,N_2554,N_2529);
xnor U2770 (N_2770,N_2475,N_2494);
or U2771 (N_2771,N_2589,N_2459);
and U2772 (N_2772,N_2578,N_2589);
nor U2773 (N_2773,N_2535,N_2595);
nor U2774 (N_2774,N_2542,N_2460);
nand U2775 (N_2775,N_2422,N_2561);
and U2776 (N_2776,N_2414,N_2543);
or U2777 (N_2777,N_2418,N_2450);
nor U2778 (N_2778,N_2553,N_2565);
xnor U2779 (N_2779,N_2400,N_2507);
nand U2780 (N_2780,N_2405,N_2522);
nor U2781 (N_2781,N_2533,N_2409);
nand U2782 (N_2782,N_2471,N_2412);
or U2783 (N_2783,N_2465,N_2507);
nor U2784 (N_2784,N_2522,N_2448);
nand U2785 (N_2785,N_2543,N_2458);
and U2786 (N_2786,N_2421,N_2597);
xor U2787 (N_2787,N_2535,N_2429);
or U2788 (N_2788,N_2500,N_2505);
nand U2789 (N_2789,N_2502,N_2587);
nand U2790 (N_2790,N_2452,N_2580);
nor U2791 (N_2791,N_2428,N_2455);
xnor U2792 (N_2792,N_2487,N_2542);
and U2793 (N_2793,N_2530,N_2404);
or U2794 (N_2794,N_2502,N_2441);
nand U2795 (N_2795,N_2457,N_2476);
xnor U2796 (N_2796,N_2545,N_2495);
and U2797 (N_2797,N_2477,N_2416);
or U2798 (N_2798,N_2556,N_2589);
and U2799 (N_2799,N_2557,N_2443);
or U2800 (N_2800,N_2696,N_2662);
or U2801 (N_2801,N_2652,N_2786);
xnor U2802 (N_2802,N_2691,N_2726);
nand U2803 (N_2803,N_2641,N_2714);
nor U2804 (N_2804,N_2703,N_2695);
and U2805 (N_2805,N_2797,N_2724);
xor U2806 (N_2806,N_2747,N_2710);
xor U2807 (N_2807,N_2784,N_2799);
and U2808 (N_2808,N_2748,N_2674);
nand U2809 (N_2809,N_2795,N_2625);
xor U2810 (N_2810,N_2755,N_2690);
nor U2811 (N_2811,N_2689,N_2779);
or U2812 (N_2812,N_2733,N_2774);
and U2813 (N_2813,N_2717,N_2741);
xor U2814 (N_2814,N_2738,N_2789);
or U2815 (N_2815,N_2701,N_2721);
nand U2816 (N_2816,N_2658,N_2629);
nand U2817 (N_2817,N_2688,N_2783);
nand U2818 (N_2818,N_2780,N_2788);
nand U2819 (N_2819,N_2796,N_2671);
and U2820 (N_2820,N_2608,N_2742);
xor U2821 (N_2821,N_2762,N_2634);
and U2822 (N_2822,N_2633,N_2759);
xnor U2823 (N_2823,N_2764,N_2749);
nand U2824 (N_2824,N_2772,N_2668);
nand U2825 (N_2825,N_2607,N_2723);
nor U2826 (N_2826,N_2720,N_2675);
nor U2827 (N_2827,N_2639,N_2781);
nand U2828 (N_2828,N_2771,N_2626);
nor U2829 (N_2829,N_2600,N_2640);
nand U2830 (N_2830,N_2654,N_2676);
xor U2831 (N_2831,N_2612,N_2790);
nor U2832 (N_2832,N_2643,N_2702);
or U2833 (N_2833,N_2673,N_2621);
nand U2834 (N_2834,N_2754,N_2740);
nand U2835 (N_2835,N_2642,N_2681);
or U2836 (N_2836,N_2704,N_2631);
nor U2837 (N_2837,N_2613,N_2773);
nand U2838 (N_2838,N_2650,N_2632);
or U2839 (N_2839,N_2678,N_2638);
xor U2840 (N_2840,N_2706,N_2793);
xor U2841 (N_2841,N_2619,N_2782);
nand U2842 (N_2842,N_2692,N_2627);
nor U2843 (N_2843,N_2653,N_2778);
or U2844 (N_2844,N_2656,N_2787);
nor U2845 (N_2845,N_2715,N_2649);
nand U2846 (N_2846,N_2729,N_2623);
or U2847 (N_2847,N_2635,N_2680);
or U2848 (N_2848,N_2611,N_2645);
nor U2849 (N_2849,N_2709,N_2760);
xnor U2850 (N_2850,N_2722,N_2769);
nor U2851 (N_2851,N_2616,N_2763);
and U2852 (N_2852,N_2767,N_2610);
nor U2853 (N_2853,N_2731,N_2604);
nor U2854 (N_2854,N_2756,N_2666);
nor U2855 (N_2855,N_2651,N_2734);
or U2856 (N_2856,N_2682,N_2670);
or U2857 (N_2857,N_2683,N_2669);
or U2858 (N_2858,N_2655,N_2730);
and U2859 (N_2859,N_2617,N_2694);
nand U2860 (N_2860,N_2644,N_2758);
nor U2861 (N_2861,N_2687,N_2685);
and U2862 (N_2862,N_2761,N_2737);
or U2863 (N_2863,N_2727,N_2744);
xnor U2864 (N_2864,N_2665,N_2770);
xnor U2865 (N_2865,N_2719,N_2746);
nor U2866 (N_2866,N_2708,N_2697);
or U2867 (N_2867,N_2765,N_2757);
nor U2868 (N_2868,N_2725,N_2750);
and U2869 (N_2869,N_2698,N_2766);
or U2870 (N_2870,N_2776,N_2728);
nor U2871 (N_2871,N_2699,N_2605);
nand U2872 (N_2872,N_2664,N_2603);
nand U2873 (N_2873,N_2768,N_2775);
and U2874 (N_2874,N_2646,N_2606);
nor U2875 (N_2875,N_2601,N_2777);
nor U2876 (N_2876,N_2667,N_2615);
nand U2877 (N_2877,N_2751,N_2679);
nand U2878 (N_2878,N_2677,N_2636);
xor U2879 (N_2879,N_2660,N_2745);
nor U2880 (N_2880,N_2657,N_2716);
xnor U2881 (N_2881,N_2628,N_2794);
or U2882 (N_2882,N_2618,N_2693);
or U2883 (N_2883,N_2718,N_2624);
xnor U2884 (N_2884,N_2735,N_2712);
and U2885 (N_2885,N_2732,N_2659);
nand U2886 (N_2886,N_2672,N_2791);
xnor U2887 (N_2887,N_2752,N_2648);
nor U2888 (N_2888,N_2739,N_2743);
or U2889 (N_2889,N_2647,N_2736);
nor U2890 (N_2890,N_2713,N_2785);
and U2891 (N_2891,N_2602,N_2661);
and U2892 (N_2892,N_2663,N_2630);
or U2893 (N_2893,N_2620,N_2705);
nor U2894 (N_2894,N_2798,N_2753);
nand U2895 (N_2895,N_2684,N_2637);
nor U2896 (N_2896,N_2622,N_2686);
xnor U2897 (N_2897,N_2609,N_2707);
nand U2898 (N_2898,N_2614,N_2700);
or U2899 (N_2899,N_2711,N_2792);
nand U2900 (N_2900,N_2702,N_2782);
nand U2901 (N_2901,N_2754,N_2703);
nor U2902 (N_2902,N_2687,N_2719);
xor U2903 (N_2903,N_2720,N_2749);
nand U2904 (N_2904,N_2721,N_2648);
xnor U2905 (N_2905,N_2663,N_2718);
and U2906 (N_2906,N_2678,N_2617);
and U2907 (N_2907,N_2748,N_2636);
or U2908 (N_2908,N_2647,N_2710);
nor U2909 (N_2909,N_2629,N_2652);
and U2910 (N_2910,N_2723,N_2637);
nor U2911 (N_2911,N_2608,N_2607);
nor U2912 (N_2912,N_2790,N_2741);
nor U2913 (N_2913,N_2787,N_2731);
or U2914 (N_2914,N_2779,N_2675);
and U2915 (N_2915,N_2756,N_2643);
xor U2916 (N_2916,N_2673,N_2644);
xor U2917 (N_2917,N_2632,N_2625);
or U2918 (N_2918,N_2770,N_2606);
nor U2919 (N_2919,N_2681,N_2688);
nand U2920 (N_2920,N_2626,N_2751);
and U2921 (N_2921,N_2743,N_2702);
and U2922 (N_2922,N_2681,N_2655);
nor U2923 (N_2923,N_2796,N_2784);
xnor U2924 (N_2924,N_2648,N_2683);
xor U2925 (N_2925,N_2638,N_2737);
nor U2926 (N_2926,N_2642,N_2614);
nand U2927 (N_2927,N_2710,N_2759);
and U2928 (N_2928,N_2652,N_2700);
xnor U2929 (N_2929,N_2658,N_2750);
and U2930 (N_2930,N_2778,N_2684);
nand U2931 (N_2931,N_2677,N_2694);
or U2932 (N_2932,N_2653,N_2622);
xnor U2933 (N_2933,N_2722,N_2720);
or U2934 (N_2934,N_2713,N_2733);
xor U2935 (N_2935,N_2776,N_2663);
nand U2936 (N_2936,N_2757,N_2715);
nor U2937 (N_2937,N_2707,N_2775);
and U2938 (N_2938,N_2756,N_2775);
nand U2939 (N_2939,N_2645,N_2746);
nand U2940 (N_2940,N_2728,N_2739);
or U2941 (N_2941,N_2770,N_2777);
and U2942 (N_2942,N_2777,N_2625);
or U2943 (N_2943,N_2604,N_2616);
nand U2944 (N_2944,N_2632,N_2687);
or U2945 (N_2945,N_2726,N_2714);
xnor U2946 (N_2946,N_2742,N_2715);
nand U2947 (N_2947,N_2696,N_2604);
nand U2948 (N_2948,N_2656,N_2707);
xnor U2949 (N_2949,N_2723,N_2703);
nand U2950 (N_2950,N_2651,N_2605);
nand U2951 (N_2951,N_2625,N_2780);
or U2952 (N_2952,N_2735,N_2650);
or U2953 (N_2953,N_2664,N_2727);
xor U2954 (N_2954,N_2737,N_2782);
xnor U2955 (N_2955,N_2757,N_2721);
and U2956 (N_2956,N_2639,N_2654);
xor U2957 (N_2957,N_2797,N_2759);
xnor U2958 (N_2958,N_2708,N_2720);
xnor U2959 (N_2959,N_2740,N_2636);
xor U2960 (N_2960,N_2635,N_2662);
and U2961 (N_2961,N_2788,N_2603);
and U2962 (N_2962,N_2663,N_2757);
and U2963 (N_2963,N_2724,N_2795);
or U2964 (N_2964,N_2618,N_2633);
xor U2965 (N_2965,N_2735,N_2760);
and U2966 (N_2966,N_2781,N_2753);
and U2967 (N_2967,N_2607,N_2772);
xor U2968 (N_2968,N_2662,N_2677);
and U2969 (N_2969,N_2733,N_2601);
nand U2970 (N_2970,N_2670,N_2771);
nand U2971 (N_2971,N_2766,N_2795);
nor U2972 (N_2972,N_2760,N_2648);
nor U2973 (N_2973,N_2652,N_2673);
nand U2974 (N_2974,N_2689,N_2616);
nor U2975 (N_2975,N_2664,N_2611);
xnor U2976 (N_2976,N_2677,N_2643);
nand U2977 (N_2977,N_2642,N_2602);
nand U2978 (N_2978,N_2799,N_2716);
and U2979 (N_2979,N_2654,N_2784);
xor U2980 (N_2980,N_2606,N_2741);
nand U2981 (N_2981,N_2758,N_2723);
xor U2982 (N_2982,N_2660,N_2727);
nand U2983 (N_2983,N_2774,N_2604);
and U2984 (N_2984,N_2767,N_2719);
xnor U2985 (N_2985,N_2683,N_2771);
and U2986 (N_2986,N_2696,N_2650);
xor U2987 (N_2987,N_2691,N_2710);
and U2988 (N_2988,N_2690,N_2704);
xnor U2989 (N_2989,N_2638,N_2608);
or U2990 (N_2990,N_2714,N_2774);
xor U2991 (N_2991,N_2619,N_2741);
nor U2992 (N_2992,N_2737,N_2774);
nand U2993 (N_2993,N_2729,N_2743);
and U2994 (N_2994,N_2763,N_2757);
nor U2995 (N_2995,N_2776,N_2712);
or U2996 (N_2996,N_2635,N_2760);
nor U2997 (N_2997,N_2652,N_2747);
nand U2998 (N_2998,N_2714,N_2649);
nor U2999 (N_2999,N_2602,N_2659);
nand U3000 (N_3000,N_2971,N_2802);
xor U3001 (N_3001,N_2968,N_2881);
and U3002 (N_3002,N_2957,N_2827);
and U3003 (N_3003,N_2973,N_2993);
or U3004 (N_3004,N_2811,N_2980);
nand U3005 (N_3005,N_2871,N_2847);
or U3006 (N_3006,N_2899,N_2874);
or U3007 (N_3007,N_2801,N_2922);
or U3008 (N_3008,N_2918,N_2844);
xnor U3009 (N_3009,N_2848,N_2815);
or U3010 (N_3010,N_2999,N_2877);
or U3011 (N_3011,N_2951,N_2806);
nor U3012 (N_3012,N_2902,N_2946);
nand U3013 (N_3013,N_2903,N_2897);
nor U3014 (N_3014,N_2875,N_2990);
or U3015 (N_3015,N_2850,N_2995);
or U3016 (N_3016,N_2914,N_2958);
nor U3017 (N_3017,N_2945,N_2950);
and U3018 (N_3018,N_2896,N_2808);
nand U3019 (N_3019,N_2885,N_2954);
nor U3020 (N_3020,N_2886,N_2864);
or U3021 (N_3021,N_2913,N_2837);
nor U3022 (N_3022,N_2934,N_2842);
nor U3023 (N_3023,N_2854,N_2887);
xnor U3024 (N_3024,N_2857,N_2805);
nor U3025 (N_3025,N_2966,N_2992);
and U3026 (N_3026,N_2972,N_2952);
and U3027 (N_3027,N_2942,N_2810);
and U3028 (N_3028,N_2927,N_2868);
nor U3029 (N_3029,N_2825,N_2838);
or U3030 (N_3030,N_2959,N_2943);
or U3031 (N_3031,N_2861,N_2843);
nor U3032 (N_3032,N_2823,N_2863);
xnor U3033 (N_3033,N_2814,N_2858);
nor U3034 (N_3034,N_2828,N_2878);
and U3035 (N_3035,N_2949,N_2905);
nand U3036 (N_3036,N_2818,N_2994);
nand U3037 (N_3037,N_2845,N_2860);
nand U3038 (N_3038,N_2944,N_2884);
nor U3039 (N_3039,N_2981,N_2901);
and U3040 (N_3040,N_2900,N_2925);
xnor U3041 (N_3041,N_2831,N_2872);
xor U3042 (N_3042,N_2907,N_2832);
nand U3043 (N_3043,N_2979,N_2933);
xor U3044 (N_3044,N_2867,N_2813);
or U3045 (N_3045,N_2879,N_2987);
or U3046 (N_3046,N_2873,N_2910);
nor U3047 (N_3047,N_2839,N_2841);
nor U3048 (N_3048,N_2812,N_2835);
or U3049 (N_3049,N_2865,N_2965);
xor U3050 (N_3050,N_2932,N_2894);
and U3051 (N_3051,N_2890,N_2807);
and U3052 (N_3052,N_2856,N_2975);
nand U3053 (N_3053,N_2817,N_2928);
xor U3054 (N_3054,N_2880,N_2988);
xnor U3055 (N_3055,N_2866,N_2820);
nand U3056 (N_3056,N_2803,N_2935);
xor U3057 (N_3057,N_2974,N_2908);
nor U3058 (N_3058,N_2969,N_2986);
nand U3059 (N_3059,N_2809,N_2826);
nand U3060 (N_3060,N_2898,N_2853);
nand U3061 (N_3061,N_2998,N_2930);
and U3062 (N_3062,N_2940,N_2924);
xnor U3063 (N_3063,N_2917,N_2985);
or U3064 (N_3064,N_2834,N_2893);
or U3065 (N_3065,N_2947,N_2983);
xor U3066 (N_3066,N_2816,N_2955);
or U3067 (N_3067,N_2984,N_2889);
and U3068 (N_3068,N_2859,N_2855);
or U3069 (N_3069,N_2911,N_2846);
and U3070 (N_3070,N_2840,N_2829);
and U3071 (N_3071,N_2851,N_2800);
nand U3072 (N_3072,N_2982,N_2912);
or U3073 (N_3073,N_2970,N_2937);
nor U3074 (N_3074,N_2916,N_2967);
nand U3075 (N_3075,N_2906,N_2956);
nor U3076 (N_3076,N_2962,N_2929);
xnor U3077 (N_3077,N_2804,N_2964);
xnor U3078 (N_3078,N_2991,N_2920);
or U3079 (N_3079,N_2976,N_2833);
nor U3080 (N_3080,N_2931,N_2939);
nand U3081 (N_3081,N_2936,N_2953);
nand U3082 (N_3082,N_2997,N_2869);
xor U3083 (N_3083,N_2862,N_2977);
nand U3084 (N_3084,N_2915,N_2824);
nor U3085 (N_3085,N_2888,N_2819);
or U3086 (N_3086,N_2919,N_2849);
xor U3087 (N_3087,N_2926,N_2960);
or U3088 (N_3088,N_2941,N_2978);
xor U3089 (N_3089,N_2852,N_2836);
nor U3090 (N_3090,N_2821,N_2996);
nor U3091 (N_3091,N_2882,N_2895);
nor U3092 (N_3092,N_2830,N_2870);
nand U3093 (N_3093,N_2989,N_2822);
xnor U3094 (N_3094,N_2923,N_2948);
nand U3095 (N_3095,N_2963,N_2904);
nand U3096 (N_3096,N_2909,N_2938);
nor U3097 (N_3097,N_2892,N_2883);
and U3098 (N_3098,N_2876,N_2961);
xnor U3099 (N_3099,N_2891,N_2921);
xor U3100 (N_3100,N_2960,N_2952);
nand U3101 (N_3101,N_2848,N_2936);
nor U3102 (N_3102,N_2954,N_2837);
nor U3103 (N_3103,N_2872,N_2833);
and U3104 (N_3104,N_2990,N_2948);
xor U3105 (N_3105,N_2839,N_2921);
nor U3106 (N_3106,N_2884,N_2997);
xor U3107 (N_3107,N_2939,N_2905);
xor U3108 (N_3108,N_2927,N_2914);
nor U3109 (N_3109,N_2866,N_2833);
nand U3110 (N_3110,N_2868,N_2976);
nor U3111 (N_3111,N_2848,N_2977);
nor U3112 (N_3112,N_2883,N_2933);
nor U3113 (N_3113,N_2892,N_2821);
nor U3114 (N_3114,N_2851,N_2884);
or U3115 (N_3115,N_2828,N_2810);
nand U3116 (N_3116,N_2863,N_2936);
and U3117 (N_3117,N_2967,N_2805);
xnor U3118 (N_3118,N_2981,N_2801);
nor U3119 (N_3119,N_2896,N_2832);
or U3120 (N_3120,N_2981,N_2954);
and U3121 (N_3121,N_2931,N_2854);
and U3122 (N_3122,N_2918,N_2838);
or U3123 (N_3123,N_2945,N_2931);
and U3124 (N_3124,N_2980,N_2927);
nor U3125 (N_3125,N_2910,N_2975);
and U3126 (N_3126,N_2858,N_2925);
nand U3127 (N_3127,N_2993,N_2843);
nand U3128 (N_3128,N_2963,N_2983);
or U3129 (N_3129,N_2881,N_2845);
and U3130 (N_3130,N_2834,N_2999);
and U3131 (N_3131,N_2958,N_2803);
xnor U3132 (N_3132,N_2844,N_2810);
or U3133 (N_3133,N_2943,N_2977);
nand U3134 (N_3134,N_2826,N_2924);
and U3135 (N_3135,N_2875,N_2817);
nand U3136 (N_3136,N_2912,N_2955);
nand U3137 (N_3137,N_2935,N_2893);
nor U3138 (N_3138,N_2984,N_2950);
or U3139 (N_3139,N_2995,N_2803);
nand U3140 (N_3140,N_2965,N_2939);
nand U3141 (N_3141,N_2937,N_2880);
or U3142 (N_3142,N_2962,N_2937);
and U3143 (N_3143,N_2910,N_2920);
nor U3144 (N_3144,N_2997,N_2852);
nand U3145 (N_3145,N_2928,N_2874);
or U3146 (N_3146,N_2874,N_2872);
nor U3147 (N_3147,N_2805,N_2868);
xor U3148 (N_3148,N_2834,N_2966);
or U3149 (N_3149,N_2966,N_2839);
xnor U3150 (N_3150,N_2897,N_2883);
or U3151 (N_3151,N_2915,N_2809);
and U3152 (N_3152,N_2975,N_2847);
or U3153 (N_3153,N_2953,N_2901);
or U3154 (N_3154,N_2830,N_2943);
nand U3155 (N_3155,N_2859,N_2825);
or U3156 (N_3156,N_2910,N_2953);
and U3157 (N_3157,N_2951,N_2903);
xnor U3158 (N_3158,N_2883,N_2867);
and U3159 (N_3159,N_2838,N_2833);
xor U3160 (N_3160,N_2807,N_2990);
nor U3161 (N_3161,N_2943,N_2885);
nor U3162 (N_3162,N_2840,N_2948);
nor U3163 (N_3163,N_2901,N_2929);
xnor U3164 (N_3164,N_2903,N_2914);
nand U3165 (N_3165,N_2831,N_2953);
or U3166 (N_3166,N_2829,N_2809);
or U3167 (N_3167,N_2987,N_2822);
and U3168 (N_3168,N_2922,N_2838);
xnor U3169 (N_3169,N_2841,N_2877);
and U3170 (N_3170,N_2882,N_2859);
and U3171 (N_3171,N_2833,N_2909);
nor U3172 (N_3172,N_2831,N_2862);
xnor U3173 (N_3173,N_2872,N_2929);
or U3174 (N_3174,N_2951,N_2843);
nor U3175 (N_3175,N_2978,N_2843);
or U3176 (N_3176,N_2892,N_2946);
xnor U3177 (N_3177,N_2842,N_2945);
nor U3178 (N_3178,N_2917,N_2833);
nor U3179 (N_3179,N_2940,N_2805);
nand U3180 (N_3180,N_2890,N_2953);
and U3181 (N_3181,N_2838,N_2990);
nor U3182 (N_3182,N_2941,N_2945);
or U3183 (N_3183,N_2834,N_2948);
xnor U3184 (N_3184,N_2854,N_2910);
or U3185 (N_3185,N_2985,N_2886);
nand U3186 (N_3186,N_2803,N_2900);
or U3187 (N_3187,N_2806,N_2899);
or U3188 (N_3188,N_2985,N_2817);
or U3189 (N_3189,N_2845,N_2853);
or U3190 (N_3190,N_2951,N_2889);
or U3191 (N_3191,N_2885,N_2974);
or U3192 (N_3192,N_2906,N_2932);
and U3193 (N_3193,N_2952,N_2994);
nand U3194 (N_3194,N_2856,N_2949);
xnor U3195 (N_3195,N_2907,N_2844);
and U3196 (N_3196,N_2962,N_2903);
and U3197 (N_3197,N_2800,N_2900);
or U3198 (N_3198,N_2862,N_2863);
nor U3199 (N_3199,N_2962,N_2812);
xnor U3200 (N_3200,N_3108,N_3053);
xor U3201 (N_3201,N_3071,N_3094);
xnor U3202 (N_3202,N_3164,N_3158);
nor U3203 (N_3203,N_3023,N_3013);
nor U3204 (N_3204,N_3119,N_3122);
xor U3205 (N_3205,N_3174,N_3155);
nor U3206 (N_3206,N_3171,N_3156);
xnor U3207 (N_3207,N_3188,N_3033);
nand U3208 (N_3208,N_3190,N_3031);
nor U3209 (N_3209,N_3168,N_3159);
xor U3210 (N_3210,N_3086,N_3145);
and U3211 (N_3211,N_3185,N_3152);
nor U3212 (N_3212,N_3007,N_3125);
xor U3213 (N_3213,N_3070,N_3181);
xor U3214 (N_3214,N_3110,N_3080);
and U3215 (N_3215,N_3061,N_3090);
nand U3216 (N_3216,N_3008,N_3045);
or U3217 (N_3217,N_3089,N_3097);
or U3218 (N_3218,N_3021,N_3054);
or U3219 (N_3219,N_3170,N_3016);
xor U3220 (N_3220,N_3076,N_3077);
xor U3221 (N_3221,N_3127,N_3025);
xor U3222 (N_3222,N_3088,N_3036);
nor U3223 (N_3223,N_3015,N_3177);
and U3224 (N_3224,N_3041,N_3121);
and U3225 (N_3225,N_3172,N_3098);
nand U3226 (N_3226,N_3091,N_3028);
or U3227 (N_3227,N_3129,N_3111);
xor U3228 (N_3228,N_3176,N_3116);
or U3229 (N_3229,N_3187,N_3065);
xnor U3230 (N_3230,N_3100,N_3131);
or U3231 (N_3231,N_3020,N_3047);
and U3232 (N_3232,N_3169,N_3140);
or U3233 (N_3233,N_3027,N_3042);
or U3234 (N_3234,N_3012,N_3058);
xnor U3235 (N_3235,N_3194,N_3124);
or U3236 (N_3236,N_3186,N_3082);
nand U3237 (N_3237,N_3019,N_3114);
and U3238 (N_3238,N_3150,N_3010);
or U3239 (N_3239,N_3128,N_3143);
or U3240 (N_3240,N_3104,N_3029);
or U3241 (N_3241,N_3189,N_3115);
or U3242 (N_3242,N_3030,N_3196);
xnor U3243 (N_3243,N_3151,N_3199);
or U3244 (N_3244,N_3101,N_3092);
nor U3245 (N_3245,N_3107,N_3160);
xor U3246 (N_3246,N_3146,N_3014);
and U3247 (N_3247,N_3120,N_3141);
xnor U3248 (N_3248,N_3022,N_3099);
nor U3249 (N_3249,N_3161,N_3001);
and U3250 (N_3250,N_3103,N_3118);
xnor U3251 (N_3251,N_3044,N_3073);
and U3252 (N_3252,N_3066,N_3050);
nand U3253 (N_3253,N_3018,N_3165);
nor U3254 (N_3254,N_3034,N_3195);
and U3255 (N_3255,N_3173,N_3087);
and U3256 (N_3256,N_3138,N_3005);
xnor U3257 (N_3257,N_3198,N_3084);
nand U3258 (N_3258,N_3137,N_3144);
nand U3259 (N_3259,N_3048,N_3072);
or U3260 (N_3260,N_3166,N_3024);
xor U3261 (N_3261,N_3037,N_3004);
or U3262 (N_3262,N_3043,N_3109);
nor U3263 (N_3263,N_3049,N_3069);
xnor U3264 (N_3264,N_3130,N_3126);
or U3265 (N_3265,N_3162,N_3074);
or U3266 (N_3266,N_3135,N_3052);
or U3267 (N_3267,N_3117,N_3179);
xnor U3268 (N_3268,N_3112,N_3148);
nand U3269 (N_3269,N_3095,N_3063);
nand U3270 (N_3270,N_3039,N_3184);
or U3271 (N_3271,N_3133,N_3134);
and U3272 (N_3272,N_3035,N_3093);
and U3273 (N_3273,N_3192,N_3003);
xor U3274 (N_3274,N_3157,N_3059);
and U3275 (N_3275,N_3085,N_3147);
nor U3276 (N_3276,N_3060,N_3132);
and U3277 (N_3277,N_3011,N_3081);
xnor U3278 (N_3278,N_3017,N_3032);
nor U3279 (N_3279,N_3079,N_3163);
and U3280 (N_3280,N_3006,N_3056);
nor U3281 (N_3281,N_3153,N_3040);
xnor U3282 (N_3282,N_3113,N_3167);
nand U3283 (N_3283,N_3154,N_3136);
and U3284 (N_3284,N_3096,N_3000);
nor U3285 (N_3285,N_3062,N_3175);
or U3286 (N_3286,N_3197,N_3002);
xor U3287 (N_3287,N_3182,N_3067);
xnor U3288 (N_3288,N_3083,N_3106);
or U3289 (N_3289,N_3105,N_3191);
nor U3290 (N_3290,N_3038,N_3180);
nor U3291 (N_3291,N_3178,N_3057);
xnor U3292 (N_3292,N_3102,N_3064);
nand U3293 (N_3293,N_3055,N_3139);
xor U3294 (N_3294,N_3046,N_3149);
nand U3295 (N_3295,N_3078,N_3026);
or U3296 (N_3296,N_3183,N_3009);
or U3297 (N_3297,N_3142,N_3075);
nand U3298 (N_3298,N_3123,N_3193);
xor U3299 (N_3299,N_3068,N_3051);
and U3300 (N_3300,N_3033,N_3128);
xnor U3301 (N_3301,N_3195,N_3100);
xnor U3302 (N_3302,N_3090,N_3175);
nor U3303 (N_3303,N_3099,N_3069);
and U3304 (N_3304,N_3059,N_3190);
nor U3305 (N_3305,N_3066,N_3087);
xor U3306 (N_3306,N_3105,N_3076);
nand U3307 (N_3307,N_3014,N_3089);
nand U3308 (N_3308,N_3110,N_3191);
or U3309 (N_3309,N_3082,N_3071);
xor U3310 (N_3310,N_3179,N_3052);
or U3311 (N_3311,N_3008,N_3194);
nand U3312 (N_3312,N_3155,N_3022);
and U3313 (N_3313,N_3108,N_3131);
nand U3314 (N_3314,N_3003,N_3012);
xor U3315 (N_3315,N_3146,N_3101);
nand U3316 (N_3316,N_3180,N_3024);
xnor U3317 (N_3317,N_3192,N_3113);
xor U3318 (N_3318,N_3143,N_3037);
nand U3319 (N_3319,N_3135,N_3197);
nand U3320 (N_3320,N_3190,N_3189);
or U3321 (N_3321,N_3085,N_3021);
nand U3322 (N_3322,N_3052,N_3140);
or U3323 (N_3323,N_3093,N_3063);
and U3324 (N_3324,N_3138,N_3120);
nand U3325 (N_3325,N_3011,N_3134);
and U3326 (N_3326,N_3042,N_3019);
nor U3327 (N_3327,N_3079,N_3170);
or U3328 (N_3328,N_3088,N_3146);
nand U3329 (N_3329,N_3074,N_3100);
xnor U3330 (N_3330,N_3009,N_3176);
and U3331 (N_3331,N_3041,N_3088);
nand U3332 (N_3332,N_3091,N_3140);
nor U3333 (N_3333,N_3169,N_3115);
nor U3334 (N_3334,N_3134,N_3189);
and U3335 (N_3335,N_3113,N_3027);
nand U3336 (N_3336,N_3023,N_3095);
and U3337 (N_3337,N_3189,N_3107);
nand U3338 (N_3338,N_3194,N_3159);
xnor U3339 (N_3339,N_3009,N_3067);
nor U3340 (N_3340,N_3189,N_3083);
or U3341 (N_3341,N_3166,N_3116);
nand U3342 (N_3342,N_3081,N_3124);
and U3343 (N_3343,N_3115,N_3167);
nand U3344 (N_3344,N_3058,N_3018);
xor U3345 (N_3345,N_3140,N_3156);
and U3346 (N_3346,N_3059,N_3173);
nor U3347 (N_3347,N_3028,N_3022);
xor U3348 (N_3348,N_3102,N_3190);
or U3349 (N_3349,N_3118,N_3186);
nand U3350 (N_3350,N_3086,N_3164);
nor U3351 (N_3351,N_3146,N_3078);
and U3352 (N_3352,N_3019,N_3040);
or U3353 (N_3353,N_3056,N_3191);
xnor U3354 (N_3354,N_3035,N_3110);
or U3355 (N_3355,N_3079,N_3109);
or U3356 (N_3356,N_3054,N_3159);
and U3357 (N_3357,N_3188,N_3097);
xnor U3358 (N_3358,N_3095,N_3079);
xor U3359 (N_3359,N_3099,N_3030);
nor U3360 (N_3360,N_3035,N_3057);
nor U3361 (N_3361,N_3197,N_3116);
nor U3362 (N_3362,N_3037,N_3166);
or U3363 (N_3363,N_3083,N_3186);
nand U3364 (N_3364,N_3058,N_3140);
nand U3365 (N_3365,N_3144,N_3066);
nand U3366 (N_3366,N_3033,N_3160);
and U3367 (N_3367,N_3012,N_3095);
or U3368 (N_3368,N_3084,N_3132);
xnor U3369 (N_3369,N_3190,N_3188);
nor U3370 (N_3370,N_3166,N_3197);
xor U3371 (N_3371,N_3032,N_3070);
nand U3372 (N_3372,N_3003,N_3081);
nor U3373 (N_3373,N_3011,N_3045);
or U3374 (N_3374,N_3034,N_3144);
or U3375 (N_3375,N_3170,N_3048);
nor U3376 (N_3376,N_3149,N_3163);
and U3377 (N_3377,N_3009,N_3062);
xnor U3378 (N_3378,N_3138,N_3176);
xnor U3379 (N_3379,N_3152,N_3193);
nand U3380 (N_3380,N_3089,N_3168);
and U3381 (N_3381,N_3081,N_3085);
and U3382 (N_3382,N_3083,N_3020);
nand U3383 (N_3383,N_3053,N_3102);
or U3384 (N_3384,N_3008,N_3107);
or U3385 (N_3385,N_3195,N_3095);
and U3386 (N_3386,N_3051,N_3059);
nand U3387 (N_3387,N_3124,N_3075);
or U3388 (N_3388,N_3126,N_3166);
or U3389 (N_3389,N_3196,N_3076);
nor U3390 (N_3390,N_3170,N_3169);
and U3391 (N_3391,N_3194,N_3127);
xor U3392 (N_3392,N_3097,N_3154);
or U3393 (N_3393,N_3129,N_3083);
xor U3394 (N_3394,N_3014,N_3139);
or U3395 (N_3395,N_3059,N_3023);
and U3396 (N_3396,N_3167,N_3026);
xor U3397 (N_3397,N_3158,N_3072);
or U3398 (N_3398,N_3094,N_3196);
nand U3399 (N_3399,N_3182,N_3176);
nor U3400 (N_3400,N_3255,N_3369);
and U3401 (N_3401,N_3276,N_3318);
xnor U3402 (N_3402,N_3265,N_3293);
nand U3403 (N_3403,N_3216,N_3379);
xor U3404 (N_3404,N_3262,N_3370);
xor U3405 (N_3405,N_3323,N_3337);
nand U3406 (N_3406,N_3210,N_3294);
and U3407 (N_3407,N_3260,N_3274);
nor U3408 (N_3408,N_3253,N_3214);
nand U3409 (N_3409,N_3233,N_3336);
xnor U3410 (N_3410,N_3392,N_3303);
nor U3411 (N_3411,N_3321,N_3236);
or U3412 (N_3412,N_3368,N_3249);
xnor U3413 (N_3413,N_3281,N_3334);
xor U3414 (N_3414,N_3315,N_3302);
or U3415 (N_3415,N_3374,N_3254);
and U3416 (N_3416,N_3247,N_3277);
or U3417 (N_3417,N_3311,N_3366);
nor U3418 (N_3418,N_3299,N_3341);
nand U3419 (N_3419,N_3385,N_3378);
or U3420 (N_3420,N_3215,N_3301);
nor U3421 (N_3421,N_3373,N_3328);
xor U3422 (N_3422,N_3342,N_3237);
xnor U3423 (N_3423,N_3339,N_3376);
or U3424 (N_3424,N_3324,N_3353);
nand U3425 (N_3425,N_3267,N_3396);
nor U3426 (N_3426,N_3352,N_3355);
or U3427 (N_3427,N_3242,N_3224);
nand U3428 (N_3428,N_3398,N_3359);
and U3429 (N_3429,N_3212,N_3211);
or U3430 (N_3430,N_3351,N_3218);
nor U3431 (N_3431,N_3291,N_3346);
or U3432 (N_3432,N_3363,N_3234);
nor U3433 (N_3433,N_3223,N_3387);
or U3434 (N_3434,N_3304,N_3270);
and U3435 (N_3435,N_3329,N_3313);
or U3436 (N_3436,N_3308,N_3297);
or U3437 (N_3437,N_3203,N_3382);
or U3438 (N_3438,N_3217,N_3258);
nand U3439 (N_3439,N_3225,N_3252);
and U3440 (N_3440,N_3213,N_3283);
and U3441 (N_3441,N_3381,N_3386);
and U3442 (N_3442,N_3280,N_3333);
or U3443 (N_3443,N_3331,N_3222);
nand U3444 (N_3444,N_3309,N_3298);
and U3445 (N_3445,N_3257,N_3372);
xor U3446 (N_3446,N_3231,N_3243);
nand U3447 (N_3447,N_3312,N_3350);
nor U3448 (N_3448,N_3221,N_3202);
xor U3449 (N_3449,N_3235,N_3228);
or U3450 (N_3450,N_3360,N_3390);
nand U3451 (N_3451,N_3284,N_3383);
and U3452 (N_3452,N_3232,N_3354);
or U3453 (N_3453,N_3357,N_3227);
or U3454 (N_3454,N_3380,N_3310);
or U3455 (N_3455,N_3200,N_3306);
xor U3456 (N_3456,N_3275,N_3250);
or U3457 (N_3457,N_3362,N_3229);
xnor U3458 (N_3458,N_3201,N_3305);
nor U3459 (N_3459,N_3316,N_3261);
or U3460 (N_3460,N_3240,N_3356);
nand U3461 (N_3461,N_3367,N_3246);
nand U3462 (N_3462,N_3327,N_3361);
or U3463 (N_3463,N_3271,N_3259);
or U3464 (N_3464,N_3371,N_3399);
or U3465 (N_3465,N_3285,N_3279);
and U3466 (N_3466,N_3348,N_3395);
nor U3467 (N_3467,N_3287,N_3375);
nor U3468 (N_3468,N_3300,N_3206);
nor U3469 (N_3469,N_3244,N_3343);
or U3470 (N_3470,N_3295,N_3209);
and U3471 (N_3471,N_3289,N_3322);
nor U3472 (N_3472,N_3317,N_3226);
nand U3473 (N_3473,N_3273,N_3364);
or U3474 (N_3474,N_3344,N_3347);
xnor U3475 (N_3475,N_3286,N_3264);
xor U3476 (N_3476,N_3245,N_3397);
nor U3477 (N_3477,N_3269,N_3296);
nand U3478 (N_3478,N_3340,N_3314);
and U3479 (N_3479,N_3389,N_3263);
and U3480 (N_3480,N_3338,N_3325);
or U3481 (N_3481,N_3365,N_3251);
or U3482 (N_3482,N_3384,N_3248);
nand U3483 (N_3483,N_3330,N_3241);
or U3484 (N_3484,N_3349,N_3358);
and U3485 (N_3485,N_3345,N_3220);
or U3486 (N_3486,N_3272,N_3268);
or U3487 (N_3487,N_3319,N_3278);
nand U3488 (N_3488,N_3335,N_3391);
and U3489 (N_3489,N_3377,N_3219);
or U3490 (N_3490,N_3393,N_3256);
nor U3491 (N_3491,N_3207,N_3282);
nor U3492 (N_3492,N_3208,N_3307);
or U3493 (N_3493,N_3204,N_3326);
nand U3494 (N_3494,N_3388,N_3239);
and U3495 (N_3495,N_3266,N_3292);
and U3496 (N_3496,N_3320,N_3238);
nor U3497 (N_3497,N_3394,N_3288);
or U3498 (N_3498,N_3230,N_3290);
and U3499 (N_3499,N_3332,N_3205);
or U3500 (N_3500,N_3313,N_3331);
xnor U3501 (N_3501,N_3307,N_3226);
xnor U3502 (N_3502,N_3211,N_3322);
or U3503 (N_3503,N_3324,N_3394);
or U3504 (N_3504,N_3298,N_3238);
and U3505 (N_3505,N_3254,N_3253);
xnor U3506 (N_3506,N_3378,N_3322);
nand U3507 (N_3507,N_3232,N_3222);
nor U3508 (N_3508,N_3373,N_3338);
nor U3509 (N_3509,N_3236,N_3249);
nand U3510 (N_3510,N_3363,N_3246);
nor U3511 (N_3511,N_3395,N_3341);
xor U3512 (N_3512,N_3344,N_3233);
nor U3513 (N_3513,N_3271,N_3236);
or U3514 (N_3514,N_3233,N_3350);
nand U3515 (N_3515,N_3392,N_3263);
nand U3516 (N_3516,N_3298,N_3352);
nor U3517 (N_3517,N_3306,N_3321);
nor U3518 (N_3518,N_3223,N_3363);
and U3519 (N_3519,N_3355,N_3381);
and U3520 (N_3520,N_3248,N_3268);
nor U3521 (N_3521,N_3302,N_3320);
nor U3522 (N_3522,N_3228,N_3295);
nand U3523 (N_3523,N_3375,N_3366);
nand U3524 (N_3524,N_3382,N_3249);
xor U3525 (N_3525,N_3245,N_3253);
and U3526 (N_3526,N_3317,N_3391);
nand U3527 (N_3527,N_3259,N_3216);
and U3528 (N_3528,N_3297,N_3307);
xor U3529 (N_3529,N_3295,N_3342);
nor U3530 (N_3530,N_3306,N_3371);
xnor U3531 (N_3531,N_3370,N_3261);
and U3532 (N_3532,N_3233,N_3259);
and U3533 (N_3533,N_3324,N_3304);
nand U3534 (N_3534,N_3358,N_3221);
nand U3535 (N_3535,N_3327,N_3252);
and U3536 (N_3536,N_3229,N_3221);
nor U3537 (N_3537,N_3202,N_3293);
nor U3538 (N_3538,N_3390,N_3285);
or U3539 (N_3539,N_3375,N_3258);
and U3540 (N_3540,N_3397,N_3341);
and U3541 (N_3541,N_3215,N_3344);
nor U3542 (N_3542,N_3380,N_3268);
and U3543 (N_3543,N_3278,N_3276);
or U3544 (N_3544,N_3322,N_3352);
nand U3545 (N_3545,N_3289,N_3259);
and U3546 (N_3546,N_3318,N_3344);
and U3547 (N_3547,N_3310,N_3215);
and U3548 (N_3548,N_3297,N_3344);
xor U3549 (N_3549,N_3323,N_3381);
and U3550 (N_3550,N_3255,N_3323);
nor U3551 (N_3551,N_3294,N_3296);
or U3552 (N_3552,N_3331,N_3268);
or U3553 (N_3553,N_3278,N_3247);
or U3554 (N_3554,N_3214,N_3385);
or U3555 (N_3555,N_3257,N_3349);
and U3556 (N_3556,N_3374,N_3380);
xnor U3557 (N_3557,N_3249,N_3379);
or U3558 (N_3558,N_3380,N_3217);
or U3559 (N_3559,N_3358,N_3373);
nand U3560 (N_3560,N_3217,N_3264);
and U3561 (N_3561,N_3267,N_3203);
or U3562 (N_3562,N_3214,N_3248);
nand U3563 (N_3563,N_3376,N_3206);
and U3564 (N_3564,N_3211,N_3288);
nand U3565 (N_3565,N_3274,N_3349);
and U3566 (N_3566,N_3300,N_3323);
xnor U3567 (N_3567,N_3211,N_3287);
and U3568 (N_3568,N_3303,N_3377);
xor U3569 (N_3569,N_3347,N_3349);
nand U3570 (N_3570,N_3252,N_3344);
and U3571 (N_3571,N_3216,N_3385);
or U3572 (N_3572,N_3347,N_3355);
and U3573 (N_3573,N_3331,N_3281);
nor U3574 (N_3574,N_3322,N_3279);
or U3575 (N_3575,N_3262,N_3256);
and U3576 (N_3576,N_3206,N_3379);
and U3577 (N_3577,N_3362,N_3219);
or U3578 (N_3578,N_3258,N_3334);
and U3579 (N_3579,N_3295,N_3213);
nor U3580 (N_3580,N_3303,N_3291);
nor U3581 (N_3581,N_3249,N_3302);
nor U3582 (N_3582,N_3232,N_3387);
and U3583 (N_3583,N_3322,N_3302);
xnor U3584 (N_3584,N_3253,N_3365);
or U3585 (N_3585,N_3378,N_3364);
nor U3586 (N_3586,N_3352,N_3241);
or U3587 (N_3587,N_3332,N_3377);
and U3588 (N_3588,N_3307,N_3210);
and U3589 (N_3589,N_3203,N_3264);
nand U3590 (N_3590,N_3346,N_3373);
nor U3591 (N_3591,N_3219,N_3202);
nor U3592 (N_3592,N_3293,N_3213);
nand U3593 (N_3593,N_3297,N_3272);
nand U3594 (N_3594,N_3223,N_3305);
or U3595 (N_3595,N_3353,N_3379);
xnor U3596 (N_3596,N_3393,N_3395);
xor U3597 (N_3597,N_3338,N_3358);
and U3598 (N_3598,N_3361,N_3211);
xor U3599 (N_3599,N_3290,N_3367);
or U3600 (N_3600,N_3517,N_3572);
xor U3601 (N_3601,N_3582,N_3563);
nor U3602 (N_3602,N_3495,N_3491);
nor U3603 (N_3603,N_3569,N_3512);
xor U3604 (N_3604,N_3550,N_3448);
nor U3605 (N_3605,N_3423,N_3535);
or U3606 (N_3606,N_3466,N_3591);
nor U3607 (N_3607,N_3509,N_3496);
xnor U3608 (N_3608,N_3475,N_3426);
nor U3609 (N_3609,N_3439,N_3493);
or U3610 (N_3610,N_3531,N_3523);
or U3611 (N_3611,N_3554,N_3457);
nand U3612 (N_3612,N_3539,N_3485);
xor U3613 (N_3613,N_3417,N_3469);
and U3614 (N_3614,N_3583,N_3590);
nand U3615 (N_3615,N_3589,N_3558);
nor U3616 (N_3616,N_3415,N_3463);
or U3617 (N_3617,N_3562,N_3593);
and U3618 (N_3618,N_3408,N_3413);
nand U3619 (N_3619,N_3406,N_3443);
nand U3620 (N_3620,N_3497,N_3503);
and U3621 (N_3621,N_3471,N_3551);
and U3622 (N_3622,N_3546,N_3479);
or U3623 (N_3623,N_3559,N_3483);
nand U3624 (N_3624,N_3409,N_3412);
or U3625 (N_3625,N_3459,N_3498);
nand U3626 (N_3626,N_3545,N_3599);
xor U3627 (N_3627,N_3587,N_3514);
nand U3628 (N_3628,N_3534,N_3460);
nor U3629 (N_3629,N_3574,N_3462);
or U3630 (N_3630,N_3541,N_3596);
nand U3631 (N_3631,N_3537,N_3424);
nor U3632 (N_3632,N_3547,N_3518);
or U3633 (N_3633,N_3404,N_3484);
nand U3634 (N_3634,N_3422,N_3414);
nor U3635 (N_3635,N_3428,N_3511);
nand U3636 (N_3636,N_3425,N_3568);
xnor U3637 (N_3637,N_3499,N_3510);
or U3638 (N_3638,N_3515,N_3480);
xor U3639 (N_3639,N_3565,N_3595);
or U3640 (N_3640,N_3433,N_3598);
or U3641 (N_3641,N_3437,N_3553);
nor U3642 (N_3642,N_3490,N_3580);
nand U3643 (N_3643,N_3405,N_3427);
nor U3644 (N_3644,N_3402,N_3488);
nand U3645 (N_3645,N_3419,N_3432);
and U3646 (N_3646,N_3473,N_3555);
xor U3647 (N_3647,N_3520,N_3489);
nand U3648 (N_3648,N_3504,N_3449);
xor U3649 (N_3649,N_3500,N_3430);
xnor U3650 (N_3650,N_3564,N_3465);
and U3651 (N_3651,N_3578,N_3516);
or U3652 (N_3652,N_3573,N_3476);
nand U3653 (N_3653,N_3416,N_3456);
or U3654 (N_3654,N_3442,N_3411);
or U3655 (N_3655,N_3431,N_3435);
and U3656 (N_3656,N_3577,N_3470);
and U3657 (N_3657,N_3410,N_3527);
xor U3658 (N_3658,N_3451,N_3401);
xnor U3659 (N_3659,N_3403,N_3513);
nor U3660 (N_3660,N_3561,N_3458);
xor U3661 (N_3661,N_3530,N_3481);
or U3662 (N_3662,N_3529,N_3447);
and U3663 (N_3663,N_3521,N_3532);
nor U3664 (N_3664,N_3592,N_3571);
nor U3665 (N_3665,N_3507,N_3557);
and U3666 (N_3666,N_3434,N_3474);
and U3667 (N_3667,N_3542,N_3570);
xnor U3668 (N_3668,N_3440,N_3536);
xor U3669 (N_3669,N_3524,N_3508);
nor U3670 (N_3670,N_3552,N_3444);
nor U3671 (N_3671,N_3581,N_3533);
or U3672 (N_3672,N_3455,N_3468);
xnor U3673 (N_3673,N_3494,N_3478);
and U3674 (N_3674,N_3454,N_3528);
and U3675 (N_3675,N_3438,N_3556);
nand U3676 (N_3676,N_3467,N_3586);
and U3677 (N_3677,N_3566,N_3453);
xor U3678 (N_3678,N_3487,N_3525);
or U3679 (N_3679,N_3588,N_3567);
or U3680 (N_3680,N_3421,N_3461);
nor U3681 (N_3681,N_3579,N_3501);
nand U3682 (N_3682,N_3429,N_3544);
xnor U3683 (N_3683,N_3505,N_3482);
and U3684 (N_3684,N_3450,N_3464);
and U3685 (N_3685,N_3472,N_3519);
and U3686 (N_3686,N_3441,N_3492);
xor U3687 (N_3687,N_3486,N_3560);
or U3688 (N_3688,N_3543,N_3540);
nand U3689 (N_3689,N_3506,N_3576);
nand U3690 (N_3690,N_3538,N_3400);
nor U3691 (N_3691,N_3597,N_3526);
nor U3692 (N_3692,N_3407,N_3446);
nand U3693 (N_3693,N_3477,N_3594);
and U3694 (N_3694,N_3452,N_3522);
or U3695 (N_3695,N_3548,N_3436);
or U3696 (N_3696,N_3420,N_3445);
nor U3697 (N_3697,N_3585,N_3575);
and U3698 (N_3698,N_3584,N_3502);
nor U3699 (N_3699,N_3418,N_3549);
xnor U3700 (N_3700,N_3473,N_3484);
xnor U3701 (N_3701,N_3477,N_3526);
nand U3702 (N_3702,N_3493,N_3574);
xnor U3703 (N_3703,N_3584,N_3452);
nor U3704 (N_3704,N_3521,N_3594);
and U3705 (N_3705,N_3468,N_3566);
and U3706 (N_3706,N_3488,N_3549);
nor U3707 (N_3707,N_3515,N_3483);
and U3708 (N_3708,N_3539,N_3445);
or U3709 (N_3709,N_3547,N_3440);
nor U3710 (N_3710,N_3567,N_3483);
or U3711 (N_3711,N_3487,N_3514);
and U3712 (N_3712,N_3583,N_3448);
or U3713 (N_3713,N_3476,N_3595);
or U3714 (N_3714,N_3592,N_3505);
nor U3715 (N_3715,N_3584,N_3580);
or U3716 (N_3716,N_3438,N_3484);
xor U3717 (N_3717,N_3535,N_3506);
or U3718 (N_3718,N_3496,N_3503);
nor U3719 (N_3719,N_3493,N_3566);
nor U3720 (N_3720,N_3516,N_3474);
nor U3721 (N_3721,N_3474,N_3512);
or U3722 (N_3722,N_3508,N_3526);
xor U3723 (N_3723,N_3565,N_3412);
or U3724 (N_3724,N_3459,N_3472);
or U3725 (N_3725,N_3409,N_3592);
xor U3726 (N_3726,N_3514,N_3406);
nor U3727 (N_3727,N_3520,N_3545);
nand U3728 (N_3728,N_3531,N_3489);
or U3729 (N_3729,N_3444,N_3592);
nor U3730 (N_3730,N_3440,N_3555);
or U3731 (N_3731,N_3541,N_3597);
or U3732 (N_3732,N_3442,N_3405);
or U3733 (N_3733,N_3483,N_3556);
nor U3734 (N_3734,N_3454,N_3483);
and U3735 (N_3735,N_3582,N_3420);
or U3736 (N_3736,N_3539,N_3595);
nor U3737 (N_3737,N_3520,N_3421);
nand U3738 (N_3738,N_3450,N_3482);
and U3739 (N_3739,N_3597,N_3522);
xnor U3740 (N_3740,N_3553,N_3406);
xor U3741 (N_3741,N_3434,N_3506);
or U3742 (N_3742,N_3502,N_3585);
nor U3743 (N_3743,N_3420,N_3528);
and U3744 (N_3744,N_3589,N_3403);
and U3745 (N_3745,N_3405,N_3495);
or U3746 (N_3746,N_3410,N_3419);
or U3747 (N_3747,N_3463,N_3502);
or U3748 (N_3748,N_3451,N_3568);
nor U3749 (N_3749,N_3423,N_3550);
nand U3750 (N_3750,N_3469,N_3563);
and U3751 (N_3751,N_3457,N_3444);
and U3752 (N_3752,N_3551,N_3515);
nor U3753 (N_3753,N_3542,N_3474);
and U3754 (N_3754,N_3571,N_3405);
or U3755 (N_3755,N_3476,N_3415);
or U3756 (N_3756,N_3492,N_3464);
nor U3757 (N_3757,N_3439,N_3406);
nand U3758 (N_3758,N_3546,N_3574);
nor U3759 (N_3759,N_3532,N_3450);
xnor U3760 (N_3760,N_3565,N_3466);
xnor U3761 (N_3761,N_3565,N_3411);
nor U3762 (N_3762,N_3419,N_3540);
and U3763 (N_3763,N_3447,N_3474);
or U3764 (N_3764,N_3458,N_3427);
xnor U3765 (N_3765,N_3513,N_3454);
and U3766 (N_3766,N_3464,N_3415);
nand U3767 (N_3767,N_3548,N_3577);
xnor U3768 (N_3768,N_3543,N_3419);
xor U3769 (N_3769,N_3521,N_3584);
nand U3770 (N_3770,N_3415,N_3400);
xor U3771 (N_3771,N_3426,N_3569);
and U3772 (N_3772,N_3474,N_3566);
nor U3773 (N_3773,N_3434,N_3579);
xor U3774 (N_3774,N_3440,N_3476);
or U3775 (N_3775,N_3562,N_3457);
nand U3776 (N_3776,N_3429,N_3443);
or U3777 (N_3777,N_3488,N_3524);
xnor U3778 (N_3778,N_3462,N_3483);
and U3779 (N_3779,N_3430,N_3434);
nand U3780 (N_3780,N_3448,N_3535);
and U3781 (N_3781,N_3424,N_3510);
nand U3782 (N_3782,N_3484,N_3429);
xor U3783 (N_3783,N_3456,N_3597);
and U3784 (N_3784,N_3542,N_3589);
nand U3785 (N_3785,N_3543,N_3429);
nand U3786 (N_3786,N_3447,N_3449);
xnor U3787 (N_3787,N_3500,N_3404);
or U3788 (N_3788,N_3437,N_3410);
xnor U3789 (N_3789,N_3550,N_3528);
nand U3790 (N_3790,N_3525,N_3511);
nand U3791 (N_3791,N_3525,N_3583);
xor U3792 (N_3792,N_3576,N_3436);
nor U3793 (N_3793,N_3491,N_3510);
xor U3794 (N_3794,N_3565,N_3450);
nand U3795 (N_3795,N_3538,N_3489);
or U3796 (N_3796,N_3430,N_3409);
or U3797 (N_3797,N_3555,N_3467);
nor U3798 (N_3798,N_3528,N_3536);
or U3799 (N_3799,N_3571,N_3547);
or U3800 (N_3800,N_3783,N_3794);
and U3801 (N_3801,N_3716,N_3753);
and U3802 (N_3802,N_3664,N_3767);
xor U3803 (N_3803,N_3708,N_3650);
nor U3804 (N_3804,N_3704,N_3639);
xor U3805 (N_3805,N_3606,N_3693);
and U3806 (N_3806,N_3775,N_3763);
and U3807 (N_3807,N_3697,N_3667);
nand U3808 (N_3808,N_3727,N_3799);
and U3809 (N_3809,N_3719,N_3654);
nand U3810 (N_3810,N_3698,N_3608);
xnor U3811 (N_3811,N_3702,N_3792);
and U3812 (N_3812,N_3750,N_3793);
or U3813 (N_3813,N_3648,N_3625);
or U3814 (N_3814,N_3661,N_3757);
nand U3815 (N_3815,N_3637,N_3721);
nand U3816 (N_3816,N_3689,N_3769);
nor U3817 (N_3817,N_3718,N_3680);
or U3818 (N_3818,N_3630,N_3610);
nand U3819 (N_3819,N_3772,N_3619);
and U3820 (N_3820,N_3600,N_3602);
or U3821 (N_3821,N_3642,N_3732);
xnor U3822 (N_3822,N_3634,N_3762);
nand U3823 (N_3823,N_3657,N_3731);
or U3824 (N_3824,N_3715,N_3622);
and U3825 (N_3825,N_3605,N_3751);
nor U3826 (N_3826,N_3707,N_3612);
xnor U3827 (N_3827,N_3623,N_3786);
xnor U3828 (N_3828,N_3699,N_3668);
nor U3829 (N_3829,N_3724,N_3649);
or U3830 (N_3830,N_3764,N_3720);
or U3831 (N_3831,N_3706,N_3616);
xnor U3832 (N_3832,N_3797,N_3709);
nor U3833 (N_3833,N_3692,N_3659);
or U3834 (N_3834,N_3736,N_3603);
nand U3835 (N_3835,N_3641,N_3628);
nand U3836 (N_3836,N_3643,N_3694);
xnor U3837 (N_3837,N_3695,N_3656);
or U3838 (N_3838,N_3743,N_3655);
nand U3839 (N_3839,N_3760,N_3636);
xor U3840 (N_3840,N_3742,N_3759);
nand U3841 (N_3841,N_3703,N_3611);
nand U3842 (N_3842,N_3678,N_3669);
and U3843 (N_3843,N_3761,N_3621);
and U3844 (N_3844,N_3677,N_3739);
nand U3845 (N_3845,N_3789,N_3725);
and U3846 (N_3846,N_3632,N_3631);
xor U3847 (N_3847,N_3766,N_3713);
nand U3848 (N_3848,N_3784,N_3674);
xor U3849 (N_3849,N_3754,N_3741);
nand U3850 (N_3850,N_3723,N_3635);
or U3851 (N_3851,N_3755,N_3613);
and U3852 (N_3852,N_3685,N_3690);
nor U3853 (N_3853,N_3712,N_3618);
or U3854 (N_3854,N_3691,N_3777);
nor U3855 (N_3855,N_3679,N_3737);
nand U3856 (N_3856,N_3620,N_3744);
nand U3857 (N_3857,N_3790,N_3666);
nor U3858 (N_3858,N_3627,N_3658);
nor U3859 (N_3859,N_3673,N_3758);
nand U3860 (N_3860,N_3660,N_3671);
nor U3861 (N_3861,N_3785,N_3729);
or U3862 (N_3862,N_3684,N_3774);
or U3863 (N_3863,N_3651,N_3711);
and U3864 (N_3864,N_3609,N_3682);
and U3865 (N_3865,N_3791,N_3752);
nor U3866 (N_3866,N_3734,N_3652);
xnor U3867 (N_3867,N_3787,N_3670);
nand U3868 (N_3868,N_3735,N_3738);
nand U3869 (N_3869,N_3747,N_3701);
or U3870 (N_3870,N_3645,N_3683);
nor U3871 (N_3871,N_3781,N_3617);
xnor U3872 (N_3872,N_3644,N_3624);
nor U3873 (N_3873,N_3795,N_3717);
xor U3874 (N_3874,N_3662,N_3629);
and U3875 (N_3875,N_3638,N_3733);
or U3876 (N_3876,N_3686,N_3676);
nor U3877 (N_3877,N_3756,N_3746);
xnor U3878 (N_3878,N_3771,N_3776);
and U3879 (N_3879,N_3798,N_3696);
and U3880 (N_3880,N_3663,N_3782);
xor U3881 (N_3881,N_3687,N_3626);
nand U3882 (N_3882,N_3615,N_3779);
or U3883 (N_3883,N_3646,N_3788);
and U3884 (N_3884,N_3607,N_3633);
xor U3885 (N_3885,N_3728,N_3796);
xor U3886 (N_3886,N_3778,N_3640);
or U3887 (N_3887,N_3748,N_3681);
nand U3888 (N_3888,N_3665,N_3604);
and U3889 (N_3889,N_3722,N_3647);
xor U3890 (N_3890,N_3688,N_3765);
xnor U3891 (N_3891,N_3780,N_3730);
xnor U3892 (N_3892,N_3768,N_3714);
and U3893 (N_3893,N_3601,N_3745);
or U3894 (N_3894,N_3749,N_3770);
and U3895 (N_3895,N_3740,N_3726);
or U3896 (N_3896,N_3705,N_3672);
or U3897 (N_3897,N_3700,N_3614);
and U3898 (N_3898,N_3773,N_3653);
or U3899 (N_3899,N_3675,N_3710);
or U3900 (N_3900,N_3624,N_3603);
xnor U3901 (N_3901,N_3647,N_3617);
and U3902 (N_3902,N_3708,N_3697);
and U3903 (N_3903,N_3700,N_3752);
nor U3904 (N_3904,N_3775,N_3628);
or U3905 (N_3905,N_3600,N_3722);
or U3906 (N_3906,N_3703,N_3637);
nor U3907 (N_3907,N_3720,N_3737);
xnor U3908 (N_3908,N_3640,N_3740);
nand U3909 (N_3909,N_3688,N_3698);
or U3910 (N_3910,N_3689,N_3715);
nand U3911 (N_3911,N_3639,N_3758);
nand U3912 (N_3912,N_3690,N_3770);
or U3913 (N_3913,N_3702,N_3750);
or U3914 (N_3914,N_3748,N_3649);
and U3915 (N_3915,N_3731,N_3680);
xnor U3916 (N_3916,N_3646,N_3601);
nand U3917 (N_3917,N_3744,N_3601);
and U3918 (N_3918,N_3665,N_3731);
xor U3919 (N_3919,N_3757,N_3647);
and U3920 (N_3920,N_3601,N_3798);
nand U3921 (N_3921,N_3757,N_3666);
nor U3922 (N_3922,N_3705,N_3719);
nand U3923 (N_3923,N_3733,N_3756);
or U3924 (N_3924,N_3646,N_3614);
xor U3925 (N_3925,N_3694,N_3726);
nand U3926 (N_3926,N_3646,N_3661);
and U3927 (N_3927,N_3629,N_3711);
nor U3928 (N_3928,N_3785,N_3633);
xnor U3929 (N_3929,N_3782,N_3656);
and U3930 (N_3930,N_3725,N_3619);
nor U3931 (N_3931,N_3796,N_3634);
and U3932 (N_3932,N_3646,N_3666);
xnor U3933 (N_3933,N_3763,N_3609);
or U3934 (N_3934,N_3723,N_3622);
xnor U3935 (N_3935,N_3763,N_3795);
nand U3936 (N_3936,N_3616,N_3699);
nand U3937 (N_3937,N_3747,N_3742);
nor U3938 (N_3938,N_3612,N_3683);
or U3939 (N_3939,N_3653,N_3728);
nor U3940 (N_3940,N_3615,N_3677);
and U3941 (N_3941,N_3788,N_3780);
xnor U3942 (N_3942,N_3780,N_3726);
xor U3943 (N_3943,N_3641,N_3610);
nand U3944 (N_3944,N_3723,N_3710);
or U3945 (N_3945,N_3709,N_3777);
xnor U3946 (N_3946,N_3639,N_3675);
and U3947 (N_3947,N_3792,N_3741);
and U3948 (N_3948,N_3780,N_3709);
and U3949 (N_3949,N_3728,N_3646);
xor U3950 (N_3950,N_3706,N_3675);
nor U3951 (N_3951,N_3770,N_3629);
nand U3952 (N_3952,N_3654,N_3678);
and U3953 (N_3953,N_3723,N_3777);
nand U3954 (N_3954,N_3635,N_3642);
or U3955 (N_3955,N_3763,N_3794);
or U3956 (N_3956,N_3680,N_3794);
or U3957 (N_3957,N_3639,N_3730);
xnor U3958 (N_3958,N_3634,N_3702);
nor U3959 (N_3959,N_3771,N_3694);
xor U3960 (N_3960,N_3611,N_3626);
and U3961 (N_3961,N_3769,N_3604);
nand U3962 (N_3962,N_3722,N_3698);
nand U3963 (N_3963,N_3653,N_3770);
or U3964 (N_3964,N_3766,N_3655);
nand U3965 (N_3965,N_3654,N_3721);
or U3966 (N_3966,N_3725,N_3652);
xnor U3967 (N_3967,N_3719,N_3754);
and U3968 (N_3968,N_3794,N_3744);
nand U3969 (N_3969,N_3673,N_3677);
nand U3970 (N_3970,N_3677,N_3786);
xor U3971 (N_3971,N_3727,N_3666);
xor U3972 (N_3972,N_3644,N_3739);
nor U3973 (N_3973,N_3607,N_3626);
nor U3974 (N_3974,N_3609,N_3621);
nand U3975 (N_3975,N_3623,N_3612);
nor U3976 (N_3976,N_3690,N_3679);
and U3977 (N_3977,N_3754,N_3779);
or U3978 (N_3978,N_3600,N_3608);
or U3979 (N_3979,N_3702,N_3799);
and U3980 (N_3980,N_3799,N_3629);
xor U3981 (N_3981,N_3784,N_3752);
or U3982 (N_3982,N_3688,N_3714);
nor U3983 (N_3983,N_3615,N_3735);
xor U3984 (N_3984,N_3723,N_3771);
xnor U3985 (N_3985,N_3768,N_3601);
xor U3986 (N_3986,N_3730,N_3638);
or U3987 (N_3987,N_3692,N_3688);
xor U3988 (N_3988,N_3609,N_3655);
nand U3989 (N_3989,N_3694,N_3655);
or U3990 (N_3990,N_3761,N_3714);
nor U3991 (N_3991,N_3795,N_3664);
nor U3992 (N_3992,N_3731,N_3605);
nor U3993 (N_3993,N_3756,N_3677);
nand U3994 (N_3994,N_3735,N_3792);
nor U3995 (N_3995,N_3605,N_3690);
nand U3996 (N_3996,N_3654,N_3731);
nand U3997 (N_3997,N_3746,N_3634);
and U3998 (N_3998,N_3773,N_3645);
nand U3999 (N_3999,N_3726,N_3737);
or U4000 (N_4000,N_3830,N_3896);
and U4001 (N_4001,N_3997,N_3960);
or U4002 (N_4002,N_3996,N_3843);
or U4003 (N_4003,N_3875,N_3818);
nor U4004 (N_4004,N_3994,N_3814);
nand U4005 (N_4005,N_3863,N_3976);
or U4006 (N_4006,N_3801,N_3924);
or U4007 (N_4007,N_3870,N_3858);
nor U4008 (N_4008,N_3805,N_3820);
xnor U4009 (N_4009,N_3901,N_3918);
nand U4010 (N_4010,N_3911,N_3826);
or U4011 (N_4011,N_3894,N_3926);
or U4012 (N_4012,N_3936,N_3902);
nor U4013 (N_4013,N_3981,N_3899);
nand U4014 (N_4014,N_3846,N_3861);
or U4015 (N_4015,N_3969,N_3889);
nor U4016 (N_4016,N_3922,N_3851);
nand U4017 (N_4017,N_3937,N_3874);
nor U4018 (N_4018,N_3945,N_3944);
nand U4019 (N_4019,N_3884,N_3856);
or U4020 (N_4020,N_3844,N_3860);
or U4021 (N_4021,N_3992,N_3970);
and U4022 (N_4022,N_3932,N_3838);
or U4023 (N_4023,N_3869,N_3935);
and U4024 (N_4024,N_3862,N_3954);
nor U4025 (N_4025,N_3809,N_3842);
nor U4026 (N_4026,N_3923,N_3892);
xor U4027 (N_4027,N_3957,N_3819);
or U4028 (N_4028,N_3912,N_3890);
and U4029 (N_4029,N_3947,N_3821);
and U4030 (N_4030,N_3950,N_3998);
or U4031 (N_4031,N_3823,N_3905);
nand U4032 (N_4032,N_3864,N_3828);
nor U4033 (N_4033,N_3930,N_3943);
nor U4034 (N_4034,N_3961,N_3877);
and U4035 (N_4035,N_3865,N_3964);
and U4036 (N_4036,N_3834,N_3979);
xnor U4037 (N_4037,N_3855,N_3891);
and U4038 (N_4038,N_3829,N_3816);
nor U4039 (N_4039,N_3822,N_3880);
and U4040 (N_4040,N_3853,N_3841);
nand U4041 (N_4041,N_3847,N_3803);
or U4042 (N_4042,N_3975,N_3854);
xnor U4043 (N_4043,N_3872,N_3968);
and U4044 (N_4044,N_3831,N_3906);
nor U4045 (N_4045,N_3807,N_3948);
nor U4046 (N_4046,N_3983,N_3832);
nand U4047 (N_4047,N_3852,N_3991);
and U4048 (N_4048,N_3993,N_3833);
and U4049 (N_4049,N_3859,N_3928);
xnor U4050 (N_4050,N_3910,N_3953);
and U4051 (N_4051,N_3956,N_3980);
xnor U4052 (N_4052,N_3929,N_3988);
xnor U4053 (N_4053,N_3837,N_3967);
nor U4054 (N_4054,N_3958,N_3972);
or U4055 (N_4055,N_3949,N_3882);
nor U4056 (N_4056,N_3914,N_3893);
nand U4057 (N_4057,N_3931,N_3873);
or U4058 (N_4058,N_3898,N_3920);
nand U4059 (N_4059,N_3999,N_3989);
or U4060 (N_4060,N_3987,N_3955);
nor U4061 (N_4061,N_3825,N_3900);
and U4062 (N_4062,N_3963,N_3804);
nor U4063 (N_4063,N_3977,N_3925);
or U4064 (N_4064,N_3995,N_3933);
or U4065 (N_4065,N_3857,N_3836);
nand U4066 (N_4066,N_3913,N_3840);
nor U4067 (N_4067,N_3962,N_3849);
nor U4068 (N_4068,N_3986,N_3941);
xor U4069 (N_4069,N_3966,N_3904);
nor U4070 (N_4070,N_3815,N_3878);
and U4071 (N_4071,N_3982,N_3824);
nor U4072 (N_4072,N_3984,N_3897);
xnor U4073 (N_4073,N_3802,N_3938);
and U4074 (N_4074,N_3908,N_3876);
and U4075 (N_4075,N_3903,N_3940);
or U4076 (N_4076,N_3919,N_3839);
and U4077 (N_4077,N_3800,N_3985);
nand U4078 (N_4078,N_3850,N_3871);
and U4079 (N_4079,N_3973,N_3952);
nor U4080 (N_4080,N_3845,N_3881);
or U4081 (N_4081,N_3946,N_3965);
or U4082 (N_4082,N_3868,N_3990);
xnor U4083 (N_4083,N_3812,N_3971);
nor U4084 (N_4084,N_3808,N_3886);
nand U4085 (N_4085,N_3927,N_3848);
and U4086 (N_4086,N_3888,N_3883);
nor U4087 (N_4087,N_3939,N_3879);
nor U4088 (N_4088,N_3810,N_3942);
and U4089 (N_4089,N_3835,N_3978);
xnor U4090 (N_4090,N_3951,N_3867);
nand U4091 (N_4091,N_3887,N_3885);
xnor U4092 (N_4092,N_3895,N_3959);
and U4093 (N_4093,N_3909,N_3827);
or U4094 (N_4094,N_3917,N_3813);
and U4095 (N_4095,N_3866,N_3974);
or U4096 (N_4096,N_3817,N_3806);
or U4097 (N_4097,N_3811,N_3921);
and U4098 (N_4098,N_3907,N_3916);
or U4099 (N_4099,N_3915,N_3934);
nand U4100 (N_4100,N_3966,N_3980);
nand U4101 (N_4101,N_3853,N_3889);
nand U4102 (N_4102,N_3946,N_3971);
and U4103 (N_4103,N_3861,N_3954);
xnor U4104 (N_4104,N_3894,N_3889);
nand U4105 (N_4105,N_3826,N_3837);
or U4106 (N_4106,N_3978,N_3801);
xnor U4107 (N_4107,N_3812,N_3977);
or U4108 (N_4108,N_3943,N_3802);
xor U4109 (N_4109,N_3938,N_3877);
and U4110 (N_4110,N_3962,N_3891);
xnor U4111 (N_4111,N_3925,N_3876);
xnor U4112 (N_4112,N_3897,N_3961);
and U4113 (N_4113,N_3802,N_3832);
or U4114 (N_4114,N_3936,N_3885);
xor U4115 (N_4115,N_3922,N_3942);
nor U4116 (N_4116,N_3969,N_3852);
nor U4117 (N_4117,N_3805,N_3914);
or U4118 (N_4118,N_3943,N_3801);
and U4119 (N_4119,N_3882,N_3802);
and U4120 (N_4120,N_3921,N_3924);
nand U4121 (N_4121,N_3863,N_3807);
and U4122 (N_4122,N_3970,N_3814);
nand U4123 (N_4123,N_3988,N_3898);
xnor U4124 (N_4124,N_3912,N_3905);
nor U4125 (N_4125,N_3802,N_3876);
and U4126 (N_4126,N_3836,N_3925);
and U4127 (N_4127,N_3887,N_3986);
xor U4128 (N_4128,N_3980,N_3960);
xor U4129 (N_4129,N_3817,N_3940);
or U4130 (N_4130,N_3935,N_3852);
and U4131 (N_4131,N_3856,N_3974);
nand U4132 (N_4132,N_3803,N_3862);
nor U4133 (N_4133,N_3813,N_3900);
nand U4134 (N_4134,N_3808,N_3819);
nor U4135 (N_4135,N_3868,N_3837);
and U4136 (N_4136,N_3860,N_3921);
and U4137 (N_4137,N_3810,N_3814);
nor U4138 (N_4138,N_3972,N_3959);
and U4139 (N_4139,N_3819,N_3870);
nor U4140 (N_4140,N_3804,N_3941);
and U4141 (N_4141,N_3847,N_3823);
nor U4142 (N_4142,N_3818,N_3978);
nor U4143 (N_4143,N_3940,N_3936);
xnor U4144 (N_4144,N_3905,N_3875);
xnor U4145 (N_4145,N_3861,N_3919);
nand U4146 (N_4146,N_3810,N_3978);
xnor U4147 (N_4147,N_3972,N_3811);
or U4148 (N_4148,N_3920,N_3986);
or U4149 (N_4149,N_3877,N_3872);
nand U4150 (N_4150,N_3861,N_3866);
xor U4151 (N_4151,N_3919,N_3806);
nand U4152 (N_4152,N_3954,N_3896);
nor U4153 (N_4153,N_3896,N_3938);
xnor U4154 (N_4154,N_3969,N_3858);
and U4155 (N_4155,N_3942,N_3881);
and U4156 (N_4156,N_3932,N_3827);
or U4157 (N_4157,N_3964,N_3889);
nand U4158 (N_4158,N_3960,N_3868);
nor U4159 (N_4159,N_3944,N_3803);
xor U4160 (N_4160,N_3854,N_3881);
or U4161 (N_4161,N_3885,N_3862);
and U4162 (N_4162,N_3809,N_3958);
and U4163 (N_4163,N_3904,N_3936);
nand U4164 (N_4164,N_3980,N_3833);
nand U4165 (N_4165,N_3848,N_3959);
and U4166 (N_4166,N_3922,N_3848);
xor U4167 (N_4167,N_3943,N_3811);
nand U4168 (N_4168,N_3998,N_3810);
or U4169 (N_4169,N_3979,N_3936);
and U4170 (N_4170,N_3982,N_3985);
xor U4171 (N_4171,N_3822,N_3988);
nor U4172 (N_4172,N_3821,N_3960);
or U4173 (N_4173,N_3863,N_3890);
nand U4174 (N_4174,N_3857,N_3807);
xnor U4175 (N_4175,N_3836,N_3914);
nand U4176 (N_4176,N_3948,N_3868);
xor U4177 (N_4177,N_3987,N_3887);
and U4178 (N_4178,N_3836,N_3899);
nor U4179 (N_4179,N_3908,N_3991);
nand U4180 (N_4180,N_3803,N_3917);
xor U4181 (N_4181,N_3925,N_3871);
and U4182 (N_4182,N_3966,N_3982);
xnor U4183 (N_4183,N_3846,N_3961);
nor U4184 (N_4184,N_3813,N_3885);
xor U4185 (N_4185,N_3980,N_3800);
nor U4186 (N_4186,N_3983,N_3831);
and U4187 (N_4187,N_3856,N_3889);
nand U4188 (N_4188,N_3833,N_3830);
nor U4189 (N_4189,N_3921,N_3856);
xnor U4190 (N_4190,N_3997,N_3897);
xor U4191 (N_4191,N_3956,N_3954);
nand U4192 (N_4192,N_3996,N_3992);
xor U4193 (N_4193,N_3872,N_3901);
or U4194 (N_4194,N_3952,N_3995);
xnor U4195 (N_4195,N_3962,N_3847);
nand U4196 (N_4196,N_3840,N_3821);
xnor U4197 (N_4197,N_3944,N_3899);
nand U4198 (N_4198,N_3999,N_3873);
nand U4199 (N_4199,N_3983,N_3849);
xor U4200 (N_4200,N_4190,N_4156);
nor U4201 (N_4201,N_4193,N_4154);
or U4202 (N_4202,N_4102,N_4145);
or U4203 (N_4203,N_4045,N_4078);
and U4204 (N_4204,N_4137,N_4014);
and U4205 (N_4205,N_4148,N_4094);
and U4206 (N_4206,N_4079,N_4088);
or U4207 (N_4207,N_4076,N_4050);
xnor U4208 (N_4208,N_4127,N_4051);
nand U4209 (N_4209,N_4100,N_4036);
and U4210 (N_4210,N_4135,N_4116);
or U4211 (N_4211,N_4044,N_4095);
or U4212 (N_4212,N_4133,N_4114);
and U4213 (N_4213,N_4058,N_4169);
or U4214 (N_4214,N_4093,N_4172);
or U4215 (N_4215,N_4181,N_4056);
xnor U4216 (N_4216,N_4042,N_4144);
or U4217 (N_4217,N_4164,N_4035);
nor U4218 (N_4218,N_4166,N_4011);
or U4219 (N_4219,N_4119,N_4087);
and U4220 (N_4220,N_4084,N_4184);
xor U4221 (N_4221,N_4165,N_4023);
nand U4222 (N_4222,N_4092,N_4168);
and U4223 (N_4223,N_4068,N_4009);
xnor U4224 (N_4224,N_4183,N_4066);
or U4225 (N_4225,N_4186,N_4090);
or U4226 (N_4226,N_4097,N_4101);
or U4227 (N_4227,N_4140,N_4053);
or U4228 (N_4228,N_4065,N_4001);
or U4229 (N_4229,N_4175,N_4083);
nor U4230 (N_4230,N_4091,N_4073);
or U4231 (N_4231,N_4107,N_4086);
or U4232 (N_4232,N_4059,N_4173);
or U4233 (N_4233,N_4039,N_4010);
xor U4234 (N_4234,N_4016,N_4006);
and U4235 (N_4235,N_4198,N_4069);
nor U4236 (N_4236,N_4103,N_4197);
nand U4237 (N_4237,N_4162,N_4124);
nand U4238 (N_4238,N_4054,N_4134);
nand U4239 (N_4239,N_4177,N_4021);
nand U4240 (N_4240,N_4109,N_4012);
xor U4241 (N_4241,N_4117,N_4070);
xnor U4242 (N_4242,N_4128,N_4029);
nand U4243 (N_4243,N_4192,N_4061);
xnor U4244 (N_4244,N_4017,N_4120);
nand U4245 (N_4245,N_4167,N_4024);
nand U4246 (N_4246,N_4188,N_4060);
xor U4247 (N_4247,N_4149,N_4112);
nand U4248 (N_4248,N_4081,N_4152);
nor U4249 (N_4249,N_4161,N_4003);
xor U4250 (N_4250,N_4046,N_4047);
nand U4251 (N_4251,N_4104,N_4130);
nor U4252 (N_4252,N_4026,N_4196);
and U4253 (N_4253,N_4187,N_4142);
xnor U4254 (N_4254,N_4085,N_4067);
nor U4255 (N_4255,N_4038,N_4031);
nand U4256 (N_4256,N_4160,N_4063);
or U4257 (N_4257,N_4015,N_4143);
and U4258 (N_4258,N_4163,N_4020);
or U4259 (N_4259,N_4132,N_4032);
nor U4260 (N_4260,N_4077,N_4136);
xnor U4261 (N_4261,N_4176,N_4155);
xnor U4262 (N_4262,N_4121,N_4055);
and U4263 (N_4263,N_4158,N_4062);
nand U4264 (N_4264,N_4041,N_4180);
xor U4265 (N_4265,N_4048,N_4111);
or U4266 (N_4266,N_4075,N_4005);
or U4267 (N_4267,N_4096,N_4071);
and U4268 (N_4268,N_4000,N_4125);
xor U4269 (N_4269,N_4129,N_4185);
and U4270 (N_4270,N_4150,N_4191);
xor U4271 (N_4271,N_4139,N_4033);
or U4272 (N_4272,N_4199,N_4131);
nand U4273 (N_4273,N_4195,N_4153);
nand U4274 (N_4274,N_4189,N_4151);
xnor U4275 (N_4275,N_4122,N_4034);
xor U4276 (N_4276,N_4182,N_4064);
nand U4277 (N_4277,N_4040,N_4080);
nor U4278 (N_4278,N_4007,N_4105);
or U4279 (N_4279,N_4108,N_4146);
xnor U4280 (N_4280,N_4004,N_4049);
or U4281 (N_4281,N_4170,N_4030);
nand U4282 (N_4282,N_4052,N_4106);
nor U4283 (N_4283,N_4002,N_4194);
nor U4284 (N_4284,N_4126,N_4123);
xnor U4285 (N_4285,N_4171,N_4179);
nand U4286 (N_4286,N_4099,N_4115);
xor U4287 (N_4287,N_4043,N_4022);
xnor U4288 (N_4288,N_4028,N_4074);
and U4289 (N_4289,N_4098,N_4008);
nor U4290 (N_4290,N_4025,N_4037);
nor U4291 (N_4291,N_4057,N_4019);
xor U4292 (N_4292,N_4027,N_4113);
and U4293 (N_4293,N_4013,N_4018);
nor U4294 (N_4294,N_4174,N_4159);
xor U4295 (N_4295,N_4138,N_4082);
nand U4296 (N_4296,N_4178,N_4157);
nor U4297 (N_4297,N_4147,N_4110);
nand U4298 (N_4298,N_4072,N_4141);
nand U4299 (N_4299,N_4089,N_4118);
nand U4300 (N_4300,N_4122,N_4092);
or U4301 (N_4301,N_4135,N_4076);
nor U4302 (N_4302,N_4120,N_4095);
and U4303 (N_4303,N_4163,N_4077);
and U4304 (N_4304,N_4091,N_4067);
xor U4305 (N_4305,N_4008,N_4015);
and U4306 (N_4306,N_4199,N_4109);
nand U4307 (N_4307,N_4056,N_4053);
nand U4308 (N_4308,N_4090,N_4062);
and U4309 (N_4309,N_4174,N_4023);
xnor U4310 (N_4310,N_4100,N_4041);
xor U4311 (N_4311,N_4199,N_4161);
and U4312 (N_4312,N_4104,N_4066);
nand U4313 (N_4313,N_4105,N_4123);
nor U4314 (N_4314,N_4009,N_4032);
and U4315 (N_4315,N_4070,N_4018);
or U4316 (N_4316,N_4175,N_4142);
nand U4317 (N_4317,N_4061,N_4060);
and U4318 (N_4318,N_4143,N_4039);
and U4319 (N_4319,N_4047,N_4097);
and U4320 (N_4320,N_4079,N_4143);
and U4321 (N_4321,N_4038,N_4028);
or U4322 (N_4322,N_4160,N_4086);
nor U4323 (N_4323,N_4038,N_4157);
or U4324 (N_4324,N_4030,N_4184);
and U4325 (N_4325,N_4076,N_4191);
and U4326 (N_4326,N_4031,N_4144);
xor U4327 (N_4327,N_4006,N_4091);
xor U4328 (N_4328,N_4060,N_4133);
nor U4329 (N_4329,N_4069,N_4148);
and U4330 (N_4330,N_4131,N_4088);
nor U4331 (N_4331,N_4155,N_4072);
nand U4332 (N_4332,N_4076,N_4103);
xor U4333 (N_4333,N_4088,N_4057);
nand U4334 (N_4334,N_4090,N_4089);
or U4335 (N_4335,N_4126,N_4048);
or U4336 (N_4336,N_4090,N_4170);
nand U4337 (N_4337,N_4094,N_4198);
nor U4338 (N_4338,N_4165,N_4147);
xnor U4339 (N_4339,N_4158,N_4044);
xor U4340 (N_4340,N_4131,N_4139);
nor U4341 (N_4341,N_4163,N_4049);
xnor U4342 (N_4342,N_4052,N_4154);
and U4343 (N_4343,N_4022,N_4135);
nor U4344 (N_4344,N_4103,N_4184);
xor U4345 (N_4345,N_4157,N_4083);
nor U4346 (N_4346,N_4036,N_4073);
or U4347 (N_4347,N_4042,N_4093);
and U4348 (N_4348,N_4027,N_4023);
and U4349 (N_4349,N_4055,N_4136);
or U4350 (N_4350,N_4132,N_4157);
nor U4351 (N_4351,N_4145,N_4159);
nand U4352 (N_4352,N_4186,N_4151);
nand U4353 (N_4353,N_4194,N_4195);
nand U4354 (N_4354,N_4181,N_4062);
and U4355 (N_4355,N_4076,N_4165);
nand U4356 (N_4356,N_4058,N_4030);
or U4357 (N_4357,N_4159,N_4148);
nand U4358 (N_4358,N_4044,N_4181);
xnor U4359 (N_4359,N_4033,N_4044);
nand U4360 (N_4360,N_4034,N_4045);
nor U4361 (N_4361,N_4160,N_4085);
or U4362 (N_4362,N_4029,N_4162);
and U4363 (N_4363,N_4031,N_4171);
nor U4364 (N_4364,N_4191,N_4048);
xnor U4365 (N_4365,N_4084,N_4080);
xnor U4366 (N_4366,N_4049,N_4081);
and U4367 (N_4367,N_4170,N_4106);
nor U4368 (N_4368,N_4104,N_4007);
nor U4369 (N_4369,N_4126,N_4061);
nor U4370 (N_4370,N_4128,N_4160);
xnor U4371 (N_4371,N_4179,N_4045);
and U4372 (N_4372,N_4041,N_4162);
or U4373 (N_4373,N_4085,N_4150);
nand U4374 (N_4374,N_4082,N_4101);
xnor U4375 (N_4375,N_4053,N_4111);
nand U4376 (N_4376,N_4181,N_4061);
nor U4377 (N_4377,N_4042,N_4135);
nor U4378 (N_4378,N_4011,N_4017);
xor U4379 (N_4379,N_4094,N_4077);
xor U4380 (N_4380,N_4001,N_4109);
nor U4381 (N_4381,N_4030,N_4136);
nand U4382 (N_4382,N_4061,N_4140);
and U4383 (N_4383,N_4167,N_4179);
nand U4384 (N_4384,N_4080,N_4145);
or U4385 (N_4385,N_4069,N_4053);
or U4386 (N_4386,N_4195,N_4173);
or U4387 (N_4387,N_4146,N_4063);
nor U4388 (N_4388,N_4176,N_4118);
or U4389 (N_4389,N_4164,N_4124);
nor U4390 (N_4390,N_4035,N_4063);
nand U4391 (N_4391,N_4064,N_4046);
xnor U4392 (N_4392,N_4161,N_4118);
nor U4393 (N_4393,N_4081,N_4033);
nor U4394 (N_4394,N_4167,N_4128);
or U4395 (N_4395,N_4084,N_4186);
nor U4396 (N_4396,N_4011,N_4163);
and U4397 (N_4397,N_4086,N_4173);
xnor U4398 (N_4398,N_4106,N_4005);
nor U4399 (N_4399,N_4008,N_4175);
or U4400 (N_4400,N_4272,N_4273);
nor U4401 (N_4401,N_4240,N_4275);
xor U4402 (N_4402,N_4386,N_4307);
and U4403 (N_4403,N_4348,N_4263);
and U4404 (N_4404,N_4347,N_4207);
nand U4405 (N_4405,N_4370,N_4242);
nand U4406 (N_4406,N_4327,N_4278);
xnor U4407 (N_4407,N_4335,N_4393);
nor U4408 (N_4408,N_4267,N_4294);
and U4409 (N_4409,N_4374,N_4320);
nand U4410 (N_4410,N_4352,N_4329);
and U4411 (N_4411,N_4222,N_4380);
and U4412 (N_4412,N_4336,N_4289);
or U4413 (N_4413,N_4300,N_4389);
or U4414 (N_4414,N_4350,N_4297);
nor U4415 (N_4415,N_4322,N_4353);
and U4416 (N_4416,N_4392,N_4293);
and U4417 (N_4417,N_4303,N_4285);
or U4418 (N_4418,N_4270,N_4344);
nor U4419 (N_4419,N_4355,N_4203);
xnor U4420 (N_4420,N_4243,N_4257);
nor U4421 (N_4421,N_4260,N_4360);
and U4422 (N_4422,N_4249,N_4206);
nand U4423 (N_4423,N_4286,N_4202);
or U4424 (N_4424,N_4213,N_4395);
or U4425 (N_4425,N_4215,N_4258);
nand U4426 (N_4426,N_4204,N_4230);
nand U4427 (N_4427,N_4354,N_4311);
nor U4428 (N_4428,N_4201,N_4217);
and U4429 (N_4429,N_4391,N_4342);
nand U4430 (N_4430,N_4276,N_4209);
or U4431 (N_4431,N_4387,N_4364);
nand U4432 (N_4432,N_4341,N_4382);
nor U4433 (N_4433,N_4223,N_4340);
nand U4434 (N_4434,N_4359,N_4264);
nor U4435 (N_4435,N_4237,N_4261);
xor U4436 (N_4436,N_4325,N_4372);
or U4437 (N_4437,N_4390,N_4259);
nor U4438 (N_4438,N_4229,N_4277);
xor U4439 (N_4439,N_4255,N_4271);
or U4440 (N_4440,N_4324,N_4385);
or U4441 (N_4441,N_4226,N_4314);
or U4442 (N_4442,N_4358,N_4315);
nor U4443 (N_4443,N_4346,N_4361);
or U4444 (N_4444,N_4274,N_4239);
nand U4445 (N_4445,N_4279,N_4396);
nor U4446 (N_4446,N_4231,N_4366);
and U4447 (N_4447,N_4345,N_4247);
nand U4448 (N_4448,N_4253,N_4357);
nand U4449 (N_4449,N_4210,N_4304);
and U4450 (N_4450,N_4312,N_4218);
nor U4451 (N_4451,N_4228,N_4319);
nor U4452 (N_4452,N_4337,N_4291);
nor U4453 (N_4453,N_4284,N_4282);
or U4454 (N_4454,N_4266,N_4292);
xor U4455 (N_4455,N_4214,N_4373);
nor U4456 (N_4456,N_4248,N_4356);
xnor U4457 (N_4457,N_4318,N_4212);
nor U4458 (N_4458,N_4349,N_4371);
nor U4459 (N_4459,N_4262,N_4323);
nand U4460 (N_4460,N_4306,N_4332);
or U4461 (N_4461,N_4316,N_4219);
and U4462 (N_4462,N_4268,N_4220);
and U4463 (N_4463,N_4383,N_4238);
or U4464 (N_4464,N_4254,N_4388);
nand U4465 (N_4465,N_4211,N_4295);
and U4466 (N_4466,N_4317,N_4368);
xor U4467 (N_4467,N_4299,N_4375);
or U4468 (N_4468,N_4321,N_4227);
nand U4469 (N_4469,N_4398,N_4296);
nor U4470 (N_4470,N_4365,N_4328);
xor U4471 (N_4471,N_4280,N_4379);
xnor U4472 (N_4472,N_4235,N_4330);
xor U4473 (N_4473,N_4378,N_4308);
nor U4474 (N_4474,N_4265,N_4241);
nor U4475 (N_4475,N_4250,N_4331);
xnor U4476 (N_4476,N_4287,N_4338);
nor U4477 (N_4477,N_4252,N_4394);
nor U4478 (N_4478,N_4281,N_4234);
or U4479 (N_4479,N_4313,N_4298);
nor U4480 (N_4480,N_4399,N_4246);
nand U4481 (N_4481,N_4205,N_4236);
nand U4482 (N_4482,N_4351,N_4326);
xnor U4483 (N_4483,N_4343,N_4305);
xnor U4484 (N_4484,N_4251,N_4269);
and U4485 (N_4485,N_4256,N_4339);
xnor U4486 (N_4486,N_4244,N_4288);
or U4487 (N_4487,N_4216,N_4310);
nor U4488 (N_4488,N_4384,N_4302);
nand U4489 (N_4489,N_4301,N_4363);
xor U4490 (N_4490,N_4200,N_4334);
and U4491 (N_4491,N_4290,N_4233);
nand U4492 (N_4492,N_4232,N_4225);
nand U4493 (N_4493,N_4221,N_4283);
xnor U4494 (N_4494,N_4309,N_4367);
nor U4495 (N_4495,N_4224,N_4397);
nor U4496 (N_4496,N_4377,N_4369);
nand U4497 (N_4497,N_4381,N_4376);
xnor U4498 (N_4498,N_4208,N_4245);
nor U4499 (N_4499,N_4362,N_4333);
nor U4500 (N_4500,N_4204,N_4212);
nor U4501 (N_4501,N_4372,N_4305);
xor U4502 (N_4502,N_4346,N_4246);
and U4503 (N_4503,N_4359,N_4299);
nor U4504 (N_4504,N_4285,N_4260);
xnor U4505 (N_4505,N_4380,N_4248);
xor U4506 (N_4506,N_4375,N_4294);
xor U4507 (N_4507,N_4357,N_4292);
xor U4508 (N_4508,N_4299,N_4320);
and U4509 (N_4509,N_4333,N_4389);
or U4510 (N_4510,N_4320,N_4338);
and U4511 (N_4511,N_4361,N_4340);
or U4512 (N_4512,N_4227,N_4283);
nor U4513 (N_4513,N_4255,N_4218);
nor U4514 (N_4514,N_4236,N_4348);
nor U4515 (N_4515,N_4299,N_4240);
xor U4516 (N_4516,N_4210,N_4301);
nor U4517 (N_4517,N_4399,N_4269);
or U4518 (N_4518,N_4228,N_4397);
nor U4519 (N_4519,N_4203,N_4379);
nand U4520 (N_4520,N_4355,N_4374);
or U4521 (N_4521,N_4348,N_4377);
nand U4522 (N_4522,N_4211,N_4383);
or U4523 (N_4523,N_4330,N_4342);
or U4524 (N_4524,N_4321,N_4398);
or U4525 (N_4525,N_4227,N_4221);
xor U4526 (N_4526,N_4226,N_4299);
and U4527 (N_4527,N_4276,N_4274);
xnor U4528 (N_4528,N_4381,N_4201);
nor U4529 (N_4529,N_4271,N_4243);
nor U4530 (N_4530,N_4386,N_4337);
xnor U4531 (N_4531,N_4246,N_4221);
xnor U4532 (N_4532,N_4254,N_4251);
nor U4533 (N_4533,N_4304,N_4384);
and U4534 (N_4534,N_4370,N_4201);
xor U4535 (N_4535,N_4360,N_4253);
xor U4536 (N_4536,N_4370,N_4257);
xnor U4537 (N_4537,N_4363,N_4361);
nor U4538 (N_4538,N_4201,N_4280);
nor U4539 (N_4539,N_4288,N_4223);
and U4540 (N_4540,N_4252,N_4385);
and U4541 (N_4541,N_4311,N_4255);
nor U4542 (N_4542,N_4217,N_4225);
or U4543 (N_4543,N_4269,N_4317);
or U4544 (N_4544,N_4252,N_4215);
nand U4545 (N_4545,N_4334,N_4252);
or U4546 (N_4546,N_4267,N_4262);
or U4547 (N_4547,N_4370,N_4280);
xnor U4548 (N_4548,N_4266,N_4303);
nor U4549 (N_4549,N_4255,N_4220);
and U4550 (N_4550,N_4393,N_4338);
nand U4551 (N_4551,N_4221,N_4366);
nand U4552 (N_4552,N_4291,N_4367);
nor U4553 (N_4553,N_4302,N_4366);
or U4554 (N_4554,N_4391,N_4264);
nand U4555 (N_4555,N_4288,N_4352);
nand U4556 (N_4556,N_4369,N_4287);
nand U4557 (N_4557,N_4228,N_4275);
nor U4558 (N_4558,N_4228,N_4284);
nand U4559 (N_4559,N_4275,N_4368);
nor U4560 (N_4560,N_4248,N_4262);
xnor U4561 (N_4561,N_4317,N_4375);
nand U4562 (N_4562,N_4352,N_4374);
nand U4563 (N_4563,N_4294,N_4291);
and U4564 (N_4564,N_4334,N_4390);
nand U4565 (N_4565,N_4389,N_4395);
nand U4566 (N_4566,N_4201,N_4215);
nor U4567 (N_4567,N_4202,N_4327);
and U4568 (N_4568,N_4332,N_4260);
nand U4569 (N_4569,N_4330,N_4218);
and U4570 (N_4570,N_4363,N_4212);
xnor U4571 (N_4571,N_4246,N_4380);
nand U4572 (N_4572,N_4314,N_4376);
or U4573 (N_4573,N_4276,N_4306);
xnor U4574 (N_4574,N_4274,N_4291);
nand U4575 (N_4575,N_4210,N_4356);
xnor U4576 (N_4576,N_4204,N_4269);
or U4577 (N_4577,N_4325,N_4251);
xor U4578 (N_4578,N_4245,N_4390);
nand U4579 (N_4579,N_4324,N_4232);
or U4580 (N_4580,N_4345,N_4368);
or U4581 (N_4581,N_4316,N_4202);
xor U4582 (N_4582,N_4288,N_4311);
xnor U4583 (N_4583,N_4286,N_4220);
nand U4584 (N_4584,N_4294,N_4321);
nand U4585 (N_4585,N_4255,N_4305);
xnor U4586 (N_4586,N_4365,N_4245);
or U4587 (N_4587,N_4228,N_4323);
or U4588 (N_4588,N_4344,N_4214);
and U4589 (N_4589,N_4323,N_4326);
xor U4590 (N_4590,N_4217,N_4232);
and U4591 (N_4591,N_4228,N_4393);
and U4592 (N_4592,N_4277,N_4395);
and U4593 (N_4593,N_4348,N_4363);
nor U4594 (N_4594,N_4397,N_4313);
or U4595 (N_4595,N_4399,N_4282);
or U4596 (N_4596,N_4296,N_4234);
xor U4597 (N_4597,N_4327,N_4201);
and U4598 (N_4598,N_4330,N_4216);
nor U4599 (N_4599,N_4264,N_4202);
or U4600 (N_4600,N_4460,N_4507);
or U4601 (N_4601,N_4474,N_4417);
nor U4602 (N_4602,N_4458,N_4412);
and U4603 (N_4603,N_4542,N_4595);
or U4604 (N_4604,N_4587,N_4598);
nand U4605 (N_4605,N_4448,N_4485);
and U4606 (N_4606,N_4555,N_4517);
or U4607 (N_4607,N_4423,N_4584);
nand U4608 (N_4608,N_4492,N_4528);
or U4609 (N_4609,N_4436,N_4403);
or U4610 (N_4610,N_4416,N_4575);
or U4611 (N_4611,N_4464,N_4490);
or U4612 (N_4612,N_4547,N_4481);
xor U4613 (N_4613,N_4411,N_4499);
nand U4614 (N_4614,N_4443,N_4553);
or U4615 (N_4615,N_4467,N_4573);
nand U4616 (N_4616,N_4459,N_4535);
or U4617 (N_4617,N_4432,N_4599);
nand U4618 (N_4618,N_4591,N_4552);
xnor U4619 (N_4619,N_4583,N_4494);
nor U4620 (N_4620,N_4454,N_4581);
nand U4621 (N_4621,N_4433,N_4408);
nor U4622 (N_4622,N_4424,N_4472);
and U4623 (N_4623,N_4419,N_4512);
or U4624 (N_4624,N_4468,N_4400);
and U4625 (N_4625,N_4502,N_4557);
nor U4626 (N_4626,N_4452,N_4427);
or U4627 (N_4627,N_4461,N_4405);
and U4628 (N_4628,N_4441,N_4420);
and U4629 (N_4629,N_4504,N_4544);
xor U4630 (N_4630,N_4520,N_4519);
xnor U4631 (N_4631,N_4550,N_4445);
or U4632 (N_4632,N_4561,N_4551);
nand U4633 (N_4633,N_4563,N_4487);
xor U4634 (N_4634,N_4523,N_4439);
or U4635 (N_4635,N_4466,N_4526);
nand U4636 (N_4636,N_4497,N_4482);
nand U4637 (N_4637,N_4508,N_4421);
nor U4638 (N_4638,N_4469,N_4567);
and U4639 (N_4639,N_4594,N_4515);
nand U4640 (N_4640,N_4522,N_4404);
nand U4641 (N_4641,N_4437,N_4409);
or U4642 (N_4642,N_4518,N_4429);
nor U4643 (N_4643,N_4509,N_4566);
xor U4644 (N_4644,N_4489,N_4449);
or U4645 (N_4645,N_4446,N_4435);
and U4646 (N_4646,N_4414,N_4440);
or U4647 (N_4647,N_4462,N_4498);
or U4648 (N_4648,N_4546,N_4442);
nor U4649 (N_4649,N_4418,N_4564);
xnor U4650 (N_4650,N_4471,N_4456);
xor U4651 (N_4651,N_4401,N_4510);
nand U4652 (N_4652,N_4493,N_4577);
or U4653 (N_4653,N_4534,N_4568);
xor U4654 (N_4654,N_4455,N_4480);
nand U4655 (N_4655,N_4506,N_4422);
nor U4656 (N_4656,N_4559,N_4428);
and U4657 (N_4657,N_4415,N_4450);
nor U4658 (N_4658,N_4505,N_4463);
nor U4659 (N_4659,N_4576,N_4501);
nor U4660 (N_4660,N_4539,N_4596);
nand U4661 (N_4661,N_4530,N_4500);
xor U4662 (N_4662,N_4570,N_4457);
xor U4663 (N_4663,N_4590,N_4572);
or U4664 (N_4664,N_4558,N_4438);
nand U4665 (N_4665,N_4549,N_4538);
nor U4666 (N_4666,N_4537,N_4470);
nand U4667 (N_4667,N_4444,N_4407);
and U4668 (N_4668,N_4543,N_4545);
nor U4669 (N_4669,N_4483,N_4488);
nor U4670 (N_4670,N_4541,N_4475);
or U4671 (N_4671,N_4425,N_4516);
or U4672 (N_4672,N_4571,N_4486);
xnor U4673 (N_4673,N_4413,N_4513);
xor U4674 (N_4674,N_4511,N_4521);
xnor U4675 (N_4675,N_4406,N_4548);
xor U4676 (N_4676,N_4465,N_4426);
nand U4677 (N_4677,N_4592,N_4560);
or U4678 (N_4678,N_4430,N_4525);
xor U4679 (N_4679,N_4589,N_4484);
nand U4680 (N_4680,N_4491,N_4579);
and U4681 (N_4681,N_4478,N_4479);
nor U4682 (N_4682,N_4410,N_4476);
xor U4683 (N_4683,N_4451,N_4585);
and U4684 (N_4684,N_4434,N_4524);
nor U4685 (N_4685,N_4569,N_4582);
or U4686 (N_4686,N_4540,N_4402);
nor U4687 (N_4687,N_4496,N_4473);
or U4688 (N_4688,N_4533,N_4477);
xor U4689 (N_4689,N_4586,N_4554);
nand U4690 (N_4690,N_4447,N_4562);
nor U4691 (N_4691,N_4503,N_4574);
nor U4692 (N_4692,N_4514,N_4529);
nor U4693 (N_4693,N_4565,N_4431);
and U4694 (N_4694,N_4527,N_4556);
xnor U4695 (N_4695,N_4593,N_4532);
xnor U4696 (N_4696,N_4580,N_4531);
nand U4697 (N_4697,N_4536,N_4597);
nand U4698 (N_4698,N_4453,N_4495);
or U4699 (N_4699,N_4588,N_4578);
and U4700 (N_4700,N_4574,N_4417);
and U4701 (N_4701,N_4547,N_4418);
or U4702 (N_4702,N_4441,N_4451);
xor U4703 (N_4703,N_4534,N_4515);
nand U4704 (N_4704,N_4431,N_4408);
or U4705 (N_4705,N_4558,N_4485);
or U4706 (N_4706,N_4470,N_4521);
xnor U4707 (N_4707,N_4494,N_4599);
xnor U4708 (N_4708,N_4562,N_4535);
or U4709 (N_4709,N_4547,N_4509);
and U4710 (N_4710,N_4540,N_4428);
nand U4711 (N_4711,N_4580,N_4491);
and U4712 (N_4712,N_4576,N_4519);
and U4713 (N_4713,N_4402,N_4450);
and U4714 (N_4714,N_4429,N_4535);
nand U4715 (N_4715,N_4490,N_4452);
and U4716 (N_4716,N_4441,N_4424);
and U4717 (N_4717,N_4584,N_4569);
xor U4718 (N_4718,N_4530,N_4589);
or U4719 (N_4719,N_4474,N_4581);
and U4720 (N_4720,N_4454,N_4429);
and U4721 (N_4721,N_4570,N_4548);
nor U4722 (N_4722,N_4584,N_4469);
or U4723 (N_4723,N_4556,N_4595);
xnor U4724 (N_4724,N_4446,N_4504);
xnor U4725 (N_4725,N_4426,N_4436);
nand U4726 (N_4726,N_4542,N_4428);
xor U4727 (N_4727,N_4415,N_4544);
or U4728 (N_4728,N_4404,N_4549);
and U4729 (N_4729,N_4447,N_4469);
and U4730 (N_4730,N_4472,N_4490);
and U4731 (N_4731,N_4408,N_4547);
nand U4732 (N_4732,N_4451,N_4521);
or U4733 (N_4733,N_4454,N_4587);
xor U4734 (N_4734,N_4461,N_4525);
xnor U4735 (N_4735,N_4472,N_4448);
or U4736 (N_4736,N_4512,N_4403);
and U4737 (N_4737,N_4539,N_4572);
nand U4738 (N_4738,N_4459,N_4426);
and U4739 (N_4739,N_4474,N_4448);
and U4740 (N_4740,N_4447,N_4436);
xor U4741 (N_4741,N_4411,N_4590);
and U4742 (N_4742,N_4518,N_4489);
and U4743 (N_4743,N_4480,N_4436);
or U4744 (N_4744,N_4432,N_4499);
or U4745 (N_4745,N_4549,N_4589);
nand U4746 (N_4746,N_4593,N_4583);
and U4747 (N_4747,N_4579,N_4515);
or U4748 (N_4748,N_4538,N_4560);
nand U4749 (N_4749,N_4532,N_4575);
nor U4750 (N_4750,N_4465,N_4596);
or U4751 (N_4751,N_4429,N_4422);
nand U4752 (N_4752,N_4552,N_4434);
xnor U4753 (N_4753,N_4512,N_4554);
xnor U4754 (N_4754,N_4534,N_4550);
or U4755 (N_4755,N_4421,N_4536);
or U4756 (N_4756,N_4562,N_4491);
nand U4757 (N_4757,N_4574,N_4587);
nand U4758 (N_4758,N_4583,N_4422);
and U4759 (N_4759,N_4450,N_4467);
or U4760 (N_4760,N_4412,N_4442);
or U4761 (N_4761,N_4457,N_4400);
and U4762 (N_4762,N_4436,N_4568);
and U4763 (N_4763,N_4510,N_4502);
nor U4764 (N_4764,N_4561,N_4539);
xnor U4765 (N_4765,N_4513,N_4524);
nor U4766 (N_4766,N_4564,N_4531);
or U4767 (N_4767,N_4506,N_4475);
xnor U4768 (N_4768,N_4432,N_4404);
nor U4769 (N_4769,N_4546,N_4563);
or U4770 (N_4770,N_4468,N_4485);
and U4771 (N_4771,N_4537,N_4465);
xor U4772 (N_4772,N_4510,N_4597);
or U4773 (N_4773,N_4593,N_4493);
nand U4774 (N_4774,N_4479,N_4577);
xnor U4775 (N_4775,N_4434,N_4579);
nor U4776 (N_4776,N_4546,N_4568);
nand U4777 (N_4777,N_4569,N_4573);
and U4778 (N_4778,N_4542,N_4585);
or U4779 (N_4779,N_4540,N_4465);
xor U4780 (N_4780,N_4517,N_4535);
nor U4781 (N_4781,N_4564,N_4437);
or U4782 (N_4782,N_4507,N_4543);
nand U4783 (N_4783,N_4580,N_4403);
xor U4784 (N_4784,N_4550,N_4441);
nand U4785 (N_4785,N_4416,N_4446);
and U4786 (N_4786,N_4401,N_4459);
nand U4787 (N_4787,N_4412,N_4422);
nand U4788 (N_4788,N_4504,N_4563);
nand U4789 (N_4789,N_4457,N_4579);
xor U4790 (N_4790,N_4522,N_4578);
and U4791 (N_4791,N_4533,N_4532);
nand U4792 (N_4792,N_4582,N_4487);
nand U4793 (N_4793,N_4537,N_4471);
and U4794 (N_4794,N_4586,N_4557);
xnor U4795 (N_4795,N_4508,N_4439);
or U4796 (N_4796,N_4572,N_4507);
nor U4797 (N_4797,N_4584,N_4589);
and U4798 (N_4798,N_4442,N_4468);
nor U4799 (N_4799,N_4458,N_4439);
nor U4800 (N_4800,N_4675,N_4766);
nand U4801 (N_4801,N_4791,N_4605);
nor U4802 (N_4802,N_4775,N_4660);
or U4803 (N_4803,N_4755,N_4787);
or U4804 (N_4804,N_4654,N_4745);
nor U4805 (N_4805,N_4757,N_4729);
or U4806 (N_4806,N_4698,N_4730);
or U4807 (N_4807,N_4752,N_4602);
nor U4808 (N_4808,N_4686,N_4677);
nor U4809 (N_4809,N_4748,N_4667);
or U4810 (N_4810,N_4792,N_4645);
and U4811 (N_4811,N_4740,N_4636);
nor U4812 (N_4812,N_4621,N_4674);
xnor U4813 (N_4813,N_4708,N_4603);
nor U4814 (N_4814,N_4756,N_4696);
nand U4815 (N_4815,N_4718,N_4710);
and U4816 (N_4816,N_4651,N_4687);
and U4817 (N_4817,N_4716,N_4774);
xnor U4818 (N_4818,N_4615,N_4772);
and U4819 (N_4819,N_4678,N_4711);
nand U4820 (N_4820,N_4689,N_4731);
nand U4821 (N_4821,N_4793,N_4709);
nor U4822 (N_4822,N_4688,N_4797);
and U4823 (N_4823,N_4768,N_4706);
nor U4824 (N_4824,N_4773,N_4692);
and U4825 (N_4825,N_4609,N_4619);
nor U4826 (N_4826,N_4650,N_4758);
nor U4827 (N_4827,N_4653,N_4722);
or U4828 (N_4828,N_4760,N_4765);
and U4829 (N_4829,N_4632,N_4707);
nor U4830 (N_4830,N_4777,N_4601);
xnor U4831 (N_4831,N_4781,N_4785);
nand U4832 (N_4832,N_4702,N_4783);
and U4833 (N_4833,N_4664,N_4700);
or U4834 (N_4834,N_4633,N_4735);
or U4835 (N_4835,N_4694,N_4670);
xor U4836 (N_4836,N_4759,N_4701);
xor U4837 (N_4837,N_4727,N_4693);
xor U4838 (N_4838,N_4613,N_4648);
xor U4839 (N_4839,N_4604,N_4637);
nand U4840 (N_4840,N_4618,N_4738);
xnor U4841 (N_4841,N_4724,N_4754);
xnor U4842 (N_4842,N_4662,N_4733);
and U4843 (N_4843,N_4771,N_4719);
nand U4844 (N_4844,N_4690,N_4607);
xor U4845 (N_4845,N_4764,N_4794);
nand U4846 (N_4846,N_4649,N_4642);
nand U4847 (N_4847,N_4681,N_4737);
and U4848 (N_4848,N_4717,N_4635);
and U4849 (N_4849,N_4665,N_4634);
and U4850 (N_4850,N_4741,N_4600);
nor U4851 (N_4851,N_4795,N_4610);
or U4852 (N_4852,N_4616,N_4747);
nand U4853 (N_4853,N_4663,N_4713);
nor U4854 (N_4854,N_4780,N_4620);
nand U4855 (N_4855,N_4631,N_4624);
and U4856 (N_4856,N_4695,N_4626);
or U4857 (N_4857,N_4625,N_4629);
and U4858 (N_4858,N_4611,N_4714);
xnor U4859 (N_4859,N_4685,N_4638);
or U4860 (N_4860,N_4657,N_4782);
or U4861 (N_4861,N_4778,N_4796);
nand U4862 (N_4862,N_4723,N_4788);
xnor U4863 (N_4863,N_4646,N_4715);
nor U4864 (N_4864,N_4680,N_4669);
nand U4865 (N_4865,N_4753,N_4767);
xnor U4866 (N_4866,N_4750,N_4655);
nor U4867 (N_4867,N_4732,N_4789);
nor U4868 (N_4868,N_4744,N_4627);
xor U4869 (N_4869,N_4679,N_4652);
xor U4870 (N_4870,N_4671,N_4683);
nor U4871 (N_4871,N_4672,N_4691);
and U4872 (N_4872,N_4612,N_4630);
and U4873 (N_4873,N_4704,N_4786);
xnor U4874 (N_4874,N_4673,N_4628);
nand U4875 (N_4875,N_4762,N_4703);
nor U4876 (N_4876,N_4726,N_4658);
nand U4877 (N_4877,N_4721,N_4712);
nand U4878 (N_4878,N_4640,N_4705);
xnor U4879 (N_4879,N_4656,N_4622);
xnor U4880 (N_4880,N_4614,N_4682);
xor U4881 (N_4881,N_4668,N_4697);
or U4882 (N_4882,N_4725,N_4799);
xnor U4883 (N_4883,N_4720,N_4769);
nor U4884 (N_4884,N_4798,N_4666);
xnor U4885 (N_4885,N_4770,N_4643);
and U4886 (N_4886,N_4623,N_4746);
and U4887 (N_4887,N_4606,N_4751);
nand U4888 (N_4888,N_4742,N_4776);
nor U4889 (N_4889,N_4644,N_4661);
or U4890 (N_4890,N_4790,N_4608);
nand U4891 (N_4891,N_4728,N_4641);
nor U4892 (N_4892,N_4734,N_4617);
or U4893 (N_4893,N_4736,N_4659);
or U4894 (N_4894,N_4699,N_4743);
xnor U4895 (N_4895,N_4676,N_4779);
and U4896 (N_4896,N_4763,N_4761);
nand U4897 (N_4897,N_4739,N_4647);
or U4898 (N_4898,N_4639,N_4784);
nand U4899 (N_4899,N_4684,N_4749);
nor U4900 (N_4900,N_4653,N_4751);
or U4901 (N_4901,N_4609,N_4755);
nand U4902 (N_4902,N_4765,N_4723);
or U4903 (N_4903,N_4663,N_4638);
and U4904 (N_4904,N_4741,N_4690);
nand U4905 (N_4905,N_4759,N_4720);
xnor U4906 (N_4906,N_4793,N_4670);
nor U4907 (N_4907,N_4604,N_4788);
or U4908 (N_4908,N_4690,N_4625);
nand U4909 (N_4909,N_4613,N_4713);
or U4910 (N_4910,N_4652,N_4678);
nor U4911 (N_4911,N_4642,N_4782);
and U4912 (N_4912,N_4715,N_4749);
nand U4913 (N_4913,N_4680,N_4774);
or U4914 (N_4914,N_4600,N_4697);
nor U4915 (N_4915,N_4698,N_4664);
or U4916 (N_4916,N_4693,N_4760);
xor U4917 (N_4917,N_4739,N_4796);
and U4918 (N_4918,N_4615,N_4768);
nand U4919 (N_4919,N_4729,N_4610);
xor U4920 (N_4920,N_4774,N_4683);
and U4921 (N_4921,N_4658,N_4612);
and U4922 (N_4922,N_4734,N_4682);
or U4923 (N_4923,N_4635,N_4622);
or U4924 (N_4924,N_4609,N_4677);
or U4925 (N_4925,N_4700,N_4647);
nand U4926 (N_4926,N_4683,N_4737);
nand U4927 (N_4927,N_4769,N_4749);
and U4928 (N_4928,N_4752,N_4680);
or U4929 (N_4929,N_4690,N_4756);
and U4930 (N_4930,N_4648,N_4771);
nor U4931 (N_4931,N_4701,N_4650);
or U4932 (N_4932,N_4771,N_4797);
or U4933 (N_4933,N_4625,N_4631);
and U4934 (N_4934,N_4770,N_4670);
and U4935 (N_4935,N_4713,N_4773);
and U4936 (N_4936,N_4697,N_4690);
or U4937 (N_4937,N_4663,N_4708);
xor U4938 (N_4938,N_4624,N_4763);
nand U4939 (N_4939,N_4651,N_4608);
nand U4940 (N_4940,N_4639,N_4721);
nand U4941 (N_4941,N_4718,N_4783);
nor U4942 (N_4942,N_4605,N_4778);
xnor U4943 (N_4943,N_4783,N_4696);
or U4944 (N_4944,N_4700,N_4717);
xor U4945 (N_4945,N_4711,N_4613);
xor U4946 (N_4946,N_4701,N_4643);
nand U4947 (N_4947,N_4720,N_4660);
xor U4948 (N_4948,N_4744,N_4692);
nand U4949 (N_4949,N_4620,N_4672);
xnor U4950 (N_4950,N_4706,N_4731);
or U4951 (N_4951,N_4702,N_4695);
xor U4952 (N_4952,N_4778,N_4666);
xor U4953 (N_4953,N_4690,N_4719);
and U4954 (N_4954,N_4792,N_4680);
nand U4955 (N_4955,N_4634,N_4734);
nor U4956 (N_4956,N_4717,N_4776);
or U4957 (N_4957,N_4616,N_4687);
or U4958 (N_4958,N_4766,N_4776);
nor U4959 (N_4959,N_4662,N_4611);
or U4960 (N_4960,N_4661,N_4781);
or U4961 (N_4961,N_4646,N_4737);
xnor U4962 (N_4962,N_4779,N_4770);
or U4963 (N_4963,N_4610,N_4721);
nor U4964 (N_4964,N_4643,N_4627);
xnor U4965 (N_4965,N_4605,N_4701);
or U4966 (N_4966,N_4696,N_4749);
nand U4967 (N_4967,N_4639,N_4746);
nand U4968 (N_4968,N_4640,N_4628);
and U4969 (N_4969,N_4715,N_4674);
nor U4970 (N_4970,N_4717,N_4753);
or U4971 (N_4971,N_4715,N_4738);
nor U4972 (N_4972,N_4627,N_4750);
and U4973 (N_4973,N_4610,N_4662);
xnor U4974 (N_4974,N_4615,N_4731);
nor U4975 (N_4975,N_4741,N_4776);
and U4976 (N_4976,N_4611,N_4722);
nor U4977 (N_4977,N_4789,N_4781);
or U4978 (N_4978,N_4667,N_4669);
and U4979 (N_4979,N_4723,N_4748);
or U4980 (N_4980,N_4647,N_4632);
or U4981 (N_4981,N_4680,N_4725);
nand U4982 (N_4982,N_4785,N_4651);
or U4983 (N_4983,N_4713,N_4639);
nor U4984 (N_4984,N_4640,N_4721);
and U4985 (N_4985,N_4726,N_4707);
nand U4986 (N_4986,N_4775,N_4671);
and U4987 (N_4987,N_4624,N_4797);
nor U4988 (N_4988,N_4664,N_4694);
and U4989 (N_4989,N_4678,N_4621);
nand U4990 (N_4990,N_4715,N_4751);
or U4991 (N_4991,N_4706,N_4689);
nand U4992 (N_4992,N_4791,N_4722);
xor U4993 (N_4993,N_4627,N_4696);
or U4994 (N_4994,N_4611,N_4747);
nand U4995 (N_4995,N_4679,N_4673);
xnor U4996 (N_4996,N_4730,N_4741);
xnor U4997 (N_4997,N_4654,N_4641);
nand U4998 (N_4998,N_4727,N_4692);
or U4999 (N_4999,N_4722,N_4645);
xnor U5000 (N_5000,N_4962,N_4940);
xor U5001 (N_5001,N_4979,N_4907);
nor U5002 (N_5002,N_4822,N_4914);
or U5003 (N_5003,N_4938,N_4836);
and U5004 (N_5004,N_4811,N_4883);
xor U5005 (N_5005,N_4876,N_4925);
and U5006 (N_5006,N_4890,N_4936);
or U5007 (N_5007,N_4964,N_4818);
nor U5008 (N_5008,N_4981,N_4951);
and U5009 (N_5009,N_4928,N_4860);
xnor U5010 (N_5010,N_4939,N_4909);
xor U5011 (N_5011,N_4934,N_4892);
or U5012 (N_5012,N_4901,N_4868);
nand U5013 (N_5013,N_4812,N_4872);
or U5014 (N_5014,N_4803,N_4800);
xor U5015 (N_5015,N_4986,N_4884);
xor U5016 (N_5016,N_4852,N_4902);
and U5017 (N_5017,N_4982,N_4987);
nor U5018 (N_5018,N_4926,N_4966);
and U5019 (N_5019,N_4993,N_4952);
nand U5020 (N_5020,N_4996,N_4817);
or U5021 (N_5021,N_4947,N_4871);
xnor U5022 (N_5022,N_4911,N_4841);
and U5023 (N_5023,N_4999,N_4848);
xnor U5024 (N_5024,N_4894,N_4815);
xor U5025 (N_5025,N_4851,N_4921);
nand U5026 (N_5026,N_4932,N_4915);
nor U5027 (N_5027,N_4943,N_4916);
or U5028 (N_5028,N_4912,N_4942);
and U5029 (N_5029,N_4953,N_4823);
and U5030 (N_5030,N_4839,N_4863);
nor U5031 (N_5031,N_4968,N_4950);
and U5032 (N_5032,N_4956,N_4917);
nor U5033 (N_5033,N_4857,N_4870);
or U5034 (N_5034,N_4819,N_4930);
or U5035 (N_5035,N_4880,N_4989);
nor U5036 (N_5036,N_4831,N_4960);
and U5037 (N_5037,N_4820,N_4903);
and U5038 (N_5038,N_4824,N_4924);
nand U5039 (N_5039,N_4963,N_4927);
nor U5040 (N_5040,N_4865,N_4975);
nor U5041 (N_5041,N_4816,N_4957);
nand U5042 (N_5042,N_4898,N_4959);
xor U5043 (N_5043,N_4881,N_4899);
and U5044 (N_5044,N_4829,N_4904);
or U5045 (N_5045,N_4888,N_4854);
nand U5046 (N_5046,N_4882,N_4843);
or U5047 (N_5047,N_4923,N_4978);
and U5048 (N_5048,N_4837,N_4809);
and U5049 (N_5049,N_4906,N_4828);
xnor U5050 (N_5050,N_4976,N_4826);
nand U5051 (N_5051,N_4922,N_4985);
nor U5052 (N_5052,N_4849,N_4858);
nand U5053 (N_5053,N_4929,N_4842);
and U5054 (N_5054,N_4980,N_4897);
nand U5055 (N_5055,N_4995,N_4965);
xnor U5056 (N_5056,N_4905,N_4887);
xnor U5057 (N_5057,N_4998,N_4955);
and U5058 (N_5058,N_4850,N_4967);
or U5059 (N_5059,N_4885,N_4873);
nor U5060 (N_5060,N_4974,N_4814);
and U5061 (N_5061,N_4830,N_4855);
nand U5062 (N_5062,N_4895,N_4886);
xnor U5063 (N_5063,N_4845,N_4838);
nand U5064 (N_5064,N_4807,N_4954);
nand U5065 (N_5065,N_4918,N_4946);
nor U5066 (N_5066,N_4935,N_4810);
nand U5067 (N_5067,N_4853,N_4844);
nor U5068 (N_5068,N_4835,N_4866);
xor U5069 (N_5069,N_4879,N_4862);
nor U5070 (N_5070,N_4802,N_4988);
or U5071 (N_5071,N_4861,N_4958);
xnor U5072 (N_5072,N_4948,N_4867);
nor U5073 (N_5073,N_4878,N_4973);
xor U5074 (N_5074,N_4847,N_4827);
or U5075 (N_5075,N_4994,N_4913);
xnor U5076 (N_5076,N_4971,N_4908);
xnor U5077 (N_5077,N_4821,N_4889);
nor U5078 (N_5078,N_4991,N_4977);
nor U5079 (N_5079,N_4896,N_4856);
nor U5080 (N_5080,N_4840,N_4970);
nand U5081 (N_5081,N_4983,N_4945);
nand U5082 (N_5082,N_4997,N_4910);
nor U5083 (N_5083,N_4875,N_4806);
xnor U5084 (N_5084,N_4808,N_4920);
or U5085 (N_5085,N_4832,N_4801);
or U5086 (N_5086,N_4990,N_4825);
nor U5087 (N_5087,N_4933,N_4961);
and U5088 (N_5088,N_4877,N_4941);
or U5089 (N_5089,N_4813,N_4984);
nor U5090 (N_5090,N_4864,N_4944);
nor U5091 (N_5091,N_4893,N_4846);
and U5092 (N_5092,N_4937,N_4805);
xnor U5093 (N_5093,N_4834,N_4874);
nor U5094 (N_5094,N_4859,N_4804);
nand U5095 (N_5095,N_4972,N_4891);
and U5096 (N_5096,N_4949,N_4869);
nor U5097 (N_5097,N_4931,N_4969);
xnor U5098 (N_5098,N_4919,N_4833);
and U5099 (N_5099,N_4992,N_4900);
nor U5100 (N_5100,N_4827,N_4937);
nor U5101 (N_5101,N_4962,N_4832);
xnor U5102 (N_5102,N_4929,N_4932);
nand U5103 (N_5103,N_4905,N_4813);
and U5104 (N_5104,N_4910,N_4918);
and U5105 (N_5105,N_4875,N_4813);
xor U5106 (N_5106,N_4990,N_4917);
nor U5107 (N_5107,N_4840,N_4804);
and U5108 (N_5108,N_4841,N_4986);
and U5109 (N_5109,N_4854,N_4910);
nor U5110 (N_5110,N_4834,N_4885);
xnor U5111 (N_5111,N_4843,N_4874);
or U5112 (N_5112,N_4819,N_4848);
and U5113 (N_5113,N_4849,N_4982);
nand U5114 (N_5114,N_4905,N_4965);
or U5115 (N_5115,N_4833,N_4990);
nor U5116 (N_5116,N_4891,N_4990);
xor U5117 (N_5117,N_4882,N_4826);
and U5118 (N_5118,N_4874,N_4804);
nand U5119 (N_5119,N_4987,N_4901);
or U5120 (N_5120,N_4932,N_4956);
nand U5121 (N_5121,N_4860,N_4833);
nor U5122 (N_5122,N_4905,N_4895);
nand U5123 (N_5123,N_4983,N_4932);
nor U5124 (N_5124,N_4956,N_4974);
nor U5125 (N_5125,N_4804,N_4955);
nor U5126 (N_5126,N_4844,N_4978);
nand U5127 (N_5127,N_4963,N_4995);
or U5128 (N_5128,N_4944,N_4816);
nand U5129 (N_5129,N_4877,N_4888);
or U5130 (N_5130,N_4978,N_4845);
nor U5131 (N_5131,N_4967,N_4949);
and U5132 (N_5132,N_4867,N_4876);
nor U5133 (N_5133,N_4974,N_4822);
xnor U5134 (N_5134,N_4986,N_4810);
or U5135 (N_5135,N_4953,N_4910);
nor U5136 (N_5136,N_4978,N_4901);
nand U5137 (N_5137,N_4810,N_4979);
and U5138 (N_5138,N_4959,N_4897);
and U5139 (N_5139,N_4882,N_4960);
nand U5140 (N_5140,N_4975,N_4925);
and U5141 (N_5141,N_4961,N_4884);
nand U5142 (N_5142,N_4977,N_4948);
nand U5143 (N_5143,N_4943,N_4841);
nor U5144 (N_5144,N_4985,N_4987);
nand U5145 (N_5145,N_4999,N_4860);
or U5146 (N_5146,N_4891,N_4977);
or U5147 (N_5147,N_4938,N_4828);
nor U5148 (N_5148,N_4827,N_4980);
nor U5149 (N_5149,N_4852,N_4967);
and U5150 (N_5150,N_4868,N_4898);
and U5151 (N_5151,N_4870,N_4858);
xnor U5152 (N_5152,N_4825,N_4977);
nand U5153 (N_5153,N_4918,N_4931);
or U5154 (N_5154,N_4864,N_4885);
nor U5155 (N_5155,N_4918,N_4811);
and U5156 (N_5156,N_4856,N_4957);
nor U5157 (N_5157,N_4855,N_4820);
xnor U5158 (N_5158,N_4928,N_4962);
or U5159 (N_5159,N_4919,N_4950);
nand U5160 (N_5160,N_4985,N_4968);
nand U5161 (N_5161,N_4943,N_4920);
xor U5162 (N_5162,N_4951,N_4805);
nor U5163 (N_5163,N_4822,N_4953);
or U5164 (N_5164,N_4909,N_4811);
and U5165 (N_5165,N_4829,N_4999);
or U5166 (N_5166,N_4816,N_4831);
or U5167 (N_5167,N_4814,N_4943);
nand U5168 (N_5168,N_4937,N_4940);
nand U5169 (N_5169,N_4837,N_4801);
and U5170 (N_5170,N_4847,N_4918);
or U5171 (N_5171,N_4962,N_4810);
nand U5172 (N_5172,N_4895,N_4979);
or U5173 (N_5173,N_4847,N_4890);
or U5174 (N_5174,N_4966,N_4815);
and U5175 (N_5175,N_4949,N_4834);
and U5176 (N_5176,N_4941,N_4908);
or U5177 (N_5177,N_4968,N_4860);
nand U5178 (N_5178,N_4962,N_4980);
nand U5179 (N_5179,N_4960,N_4935);
nor U5180 (N_5180,N_4881,N_4953);
nor U5181 (N_5181,N_4824,N_4896);
xnor U5182 (N_5182,N_4984,N_4881);
xnor U5183 (N_5183,N_4849,N_4804);
and U5184 (N_5184,N_4879,N_4950);
nor U5185 (N_5185,N_4990,N_4822);
xor U5186 (N_5186,N_4838,N_4861);
xor U5187 (N_5187,N_4875,N_4932);
nand U5188 (N_5188,N_4978,N_4898);
nor U5189 (N_5189,N_4901,N_4889);
or U5190 (N_5190,N_4891,N_4958);
and U5191 (N_5191,N_4835,N_4810);
nand U5192 (N_5192,N_4860,N_4925);
nand U5193 (N_5193,N_4933,N_4925);
nand U5194 (N_5194,N_4863,N_4910);
nor U5195 (N_5195,N_4949,N_4895);
and U5196 (N_5196,N_4800,N_4857);
and U5197 (N_5197,N_4946,N_4806);
nand U5198 (N_5198,N_4893,N_4847);
xor U5199 (N_5199,N_4807,N_4875);
nor U5200 (N_5200,N_5098,N_5033);
and U5201 (N_5201,N_5097,N_5070);
nor U5202 (N_5202,N_5106,N_5157);
and U5203 (N_5203,N_5173,N_5117);
nand U5204 (N_5204,N_5199,N_5057);
nor U5205 (N_5205,N_5022,N_5136);
xor U5206 (N_5206,N_5130,N_5104);
nor U5207 (N_5207,N_5187,N_5049);
nand U5208 (N_5208,N_5135,N_5000);
and U5209 (N_5209,N_5094,N_5195);
or U5210 (N_5210,N_5036,N_5112);
nor U5211 (N_5211,N_5066,N_5184);
xnor U5212 (N_5212,N_5023,N_5061);
and U5213 (N_5213,N_5031,N_5099);
xor U5214 (N_5214,N_5155,N_5085);
nor U5215 (N_5215,N_5043,N_5147);
nor U5216 (N_5216,N_5191,N_5142);
and U5217 (N_5217,N_5185,N_5072);
or U5218 (N_5218,N_5109,N_5039);
or U5219 (N_5219,N_5197,N_5041);
and U5220 (N_5220,N_5037,N_5071);
and U5221 (N_5221,N_5101,N_5038);
nand U5222 (N_5222,N_5081,N_5013);
nand U5223 (N_5223,N_5080,N_5167);
xnor U5224 (N_5224,N_5119,N_5161);
nand U5225 (N_5225,N_5144,N_5140);
and U5226 (N_5226,N_5074,N_5190);
nand U5227 (N_5227,N_5151,N_5143);
xor U5228 (N_5228,N_5132,N_5152);
and U5229 (N_5229,N_5020,N_5055);
xnor U5230 (N_5230,N_5133,N_5028);
nand U5231 (N_5231,N_5058,N_5016);
xor U5232 (N_5232,N_5088,N_5146);
and U5233 (N_5233,N_5174,N_5054);
nor U5234 (N_5234,N_5123,N_5069);
xor U5235 (N_5235,N_5125,N_5165);
nand U5236 (N_5236,N_5150,N_5047);
xnor U5237 (N_5237,N_5068,N_5181);
and U5238 (N_5238,N_5025,N_5192);
nor U5239 (N_5239,N_5095,N_5158);
or U5240 (N_5240,N_5021,N_5170);
nand U5241 (N_5241,N_5179,N_5018);
and U5242 (N_5242,N_5188,N_5105);
nand U5243 (N_5243,N_5107,N_5126);
nor U5244 (N_5244,N_5169,N_5073);
xor U5245 (N_5245,N_5108,N_5059);
and U5246 (N_5246,N_5160,N_5003);
nor U5247 (N_5247,N_5011,N_5046);
and U5248 (N_5248,N_5177,N_5089);
nand U5249 (N_5249,N_5086,N_5114);
nand U5250 (N_5250,N_5153,N_5005);
and U5251 (N_5251,N_5141,N_5079);
and U5252 (N_5252,N_5149,N_5015);
or U5253 (N_5253,N_5134,N_5026);
or U5254 (N_5254,N_5122,N_5002);
nand U5255 (N_5255,N_5029,N_5064);
nand U5256 (N_5256,N_5045,N_5034);
nand U5257 (N_5257,N_5024,N_5035);
nor U5258 (N_5258,N_5012,N_5083);
and U5259 (N_5259,N_5127,N_5082);
nor U5260 (N_5260,N_5096,N_5164);
nor U5261 (N_5261,N_5138,N_5111);
xor U5262 (N_5262,N_5113,N_5154);
or U5263 (N_5263,N_5006,N_5198);
nand U5264 (N_5264,N_5093,N_5010);
xor U5265 (N_5265,N_5182,N_5186);
xor U5266 (N_5266,N_5103,N_5051);
nor U5267 (N_5267,N_5168,N_5076);
nor U5268 (N_5268,N_5062,N_5116);
and U5269 (N_5269,N_5156,N_5183);
and U5270 (N_5270,N_5092,N_5008);
or U5271 (N_5271,N_5178,N_5032);
xor U5272 (N_5272,N_5060,N_5087);
xor U5273 (N_5273,N_5148,N_5189);
and U5274 (N_5274,N_5129,N_5194);
nor U5275 (N_5275,N_5131,N_5090);
nand U5276 (N_5276,N_5159,N_5056);
and U5277 (N_5277,N_5100,N_5175);
nand U5278 (N_5278,N_5166,N_5102);
or U5279 (N_5279,N_5004,N_5172);
nor U5280 (N_5280,N_5176,N_5007);
xnor U5281 (N_5281,N_5115,N_5137);
nand U5282 (N_5282,N_5063,N_5139);
xnor U5283 (N_5283,N_5030,N_5044);
xor U5284 (N_5284,N_5145,N_5118);
nand U5285 (N_5285,N_5065,N_5040);
xor U5286 (N_5286,N_5001,N_5027);
or U5287 (N_5287,N_5120,N_5162);
or U5288 (N_5288,N_5017,N_5019);
and U5289 (N_5289,N_5067,N_5084);
nand U5290 (N_5290,N_5196,N_5077);
nor U5291 (N_5291,N_5050,N_5052);
xnor U5292 (N_5292,N_5048,N_5042);
and U5293 (N_5293,N_5014,N_5091);
or U5294 (N_5294,N_5009,N_5180);
or U5295 (N_5295,N_5193,N_5075);
or U5296 (N_5296,N_5163,N_5078);
xor U5297 (N_5297,N_5128,N_5121);
or U5298 (N_5298,N_5110,N_5053);
or U5299 (N_5299,N_5124,N_5171);
xor U5300 (N_5300,N_5117,N_5185);
and U5301 (N_5301,N_5024,N_5009);
nand U5302 (N_5302,N_5018,N_5157);
nor U5303 (N_5303,N_5180,N_5087);
nor U5304 (N_5304,N_5105,N_5050);
nand U5305 (N_5305,N_5144,N_5077);
nand U5306 (N_5306,N_5081,N_5017);
nand U5307 (N_5307,N_5071,N_5142);
nand U5308 (N_5308,N_5117,N_5045);
or U5309 (N_5309,N_5035,N_5037);
or U5310 (N_5310,N_5051,N_5012);
nand U5311 (N_5311,N_5150,N_5014);
or U5312 (N_5312,N_5036,N_5090);
and U5313 (N_5313,N_5173,N_5162);
nor U5314 (N_5314,N_5077,N_5145);
nor U5315 (N_5315,N_5056,N_5193);
or U5316 (N_5316,N_5100,N_5177);
nand U5317 (N_5317,N_5093,N_5168);
nand U5318 (N_5318,N_5031,N_5040);
or U5319 (N_5319,N_5135,N_5056);
and U5320 (N_5320,N_5166,N_5025);
xnor U5321 (N_5321,N_5174,N_5159);
or U5322 (N_5322,N_5141,N_5185);
nand U5323 (N_5323,N_5116,N_5032);
or U5324 (N_5324,N_5042,N_5179);
nand U5325 (N_5325,N_5011,N_5140);
or U5326 (N_5326,N_5073,N_5092);
or U5327 (N_5327,N_5154,N_5149);
xnor U5328 (N_5328,N_5199,N_5089);
xor U5329 (N_5329,N_5091,N_5153);
nand U5330 (N_5330,N_5167,N_5067);
xnor U5331 (N_5331,N_5083,N_5042);
or U5332 (N_5332,N_5140,N_5069);
nand U5333 (N_5333,N_5047,N_5080);
nor U5334 (N_5334,N_5001,N_5085);
and U5335 (N_5335,N_5045,N_5064);
xor U5336 (N_5336,N_5003,N_5028);
nor U5337 (N_5337,N_5182,N_5056);
nor U5338 (N_5338,N_5180,N_5092);
nor U5339 (N_5339,N_5028,N_5157);
nor U5340 (N_5340,N_5182,N_5168);
nor U5341 (N_5341,N_5194,N_5037);
and U5342 (N_5342,N_5177,N_5088);
nand U5343 (N_5343,N_5171,N_5130);
and U5344 (N_5344,N_5131,N_5170);
nor U5345 (N_5345,N_5151,N_5174);
nor U5346 (N_5346,N_5003,N_5197);
nand U5347 (N_5347,N_5065,N_5084);
xnor U5348 (N_5348,N_5127,N_5133);
nand U5349 (N_5349,N_5151,N_5088);
and U5350 (N_5350,N_5160,N_5063);
nand U5351 (N_5351,N_5063,N_5110);
nor U5352 (N_5352,N_5125,N_5007);
or U5353 (N_5353,N_5039,N_5093);
nand U5354 (N_5354,N_5191,N_5129);
nand U5355 (N_5355,N_5052,N_5191);
or U5356 (N_5356,N_5168,N_5041);
xor U5357 (N_5357,N_5073,N_5127);
xnor U5358 (N_5358,N_5161,N_5156);
xor U5359 (N_5359,N_5020,N_5141);
and U5360 (N_5360,N_5049,N_5119);
or U5361 (N_5361,N_5198,N_5149);
or U5362 (N_5362,N_5180,N_5057);
and U5363 (N_5363,N_5141,N_5101);
nand U5364 (N_5364,N_5163,N_5184);
and U5365 (N_5365,N_5133,N_5155);
or U5366 (N_5366,N_5027,N_5161);
nand U5367 (N_5367,N_5036,N_5131);
and U5368 (N_5368,N_5066,N_5112);
nand U5369 (N_5369,N_5190,N_5165);
xnor U5370 (N_5370,N_5044,N_5125);
and U5371 (N_5371,N_5179,N_5058);
xor U5372 (N_5372,N_5117,N_5188);
and U5373 (N_5373,N_5149,N_5118);
and U5374 (N_5374,N_5092,N_5157);
nand U5375 (N_5375,N_5065,N_5020);
nor U5376 (N_5376,N_5056,N_5150);
and U5377 (N_5377,N_5012,N_5146);
and U5378 (N_5378,N_5166,N_5012);
nor U5379 (N_5379,N_5138,N_5190);
and U5380 (N_5380,N_5015,N_5073);
and U5381 (N_5381,N_5049,N_5088);
and U5382 (N_5382,N_5142,N_5173);
and U5383 (N_5383,N_5157,N_5162);
nand U5384 (N_5384,N_5092,N_5006);
and U5385 (N_5385,N_5059,N_5169);
or U5386 (N_5386,N_5024,N_5040);
nor U5387 (N_5387,N_5029,N_5088);
and U5388 (N_5388,N_5126,N_5153);
or U5389 (N_5389,N_5184,N_5102);
nor U5390 (N_5390,N_5040,N_5193);
xnor U5391 (N_5391,N_5008,N_5091);
and U5392 (N_5392,N_5088,N_5057);
nand U5393 (N_5393,N_5180,N_5160);
nor U5394 (N_5394,N_5059,N_5171);
nor U5395 (N_5395,N_5076,N_5162);
or U5396 (N_5396,N_5133,N_5137);
or U5397 (N_5397,N_5167,N_5186);
and U5398 (N_5398,N_5019,N_5007);
nand U5399 (N_5399,N_5183,N_5167);
and U5400 (N_5400,N_5381,N_5289);
and U5401 (N_5401,N_5338,N_5311);
nor U5402 (N_5402,N_5258,N_5242);
nand U5403 (N_5403,N_5327,N_5254);
and U5404 (N_5404,N_5382,N_5268);
nand U5405 (N_5405,N_5355,N_5253);
and U5406 (N_5406,N_5214,N_5251);
and U5407 (N_5407,N_5287,N_5349);
or U5408 (N_5408,N_5307,N_5261);
nor U5409 (N_5409,N_5284,N_5292);
or U5410 (N_5410,N_5236,N_5389);
nor U5411 (N_5411,N_5309,N_5354);
nand U5412 (N_5412,N_5276,N_5310);
and U5413 (N_5413,N_5370,N_5286);
nor U5414 (N_5414,N_5345,N_5364);
nor U5415 (N_5415,N_5323,N_5264);
nand U5416 (N_5416,N_5350,N_5288);
nor U5417 (N_5417,N_5290,N_5369);
and U5418 (N_5418,N_5352,N_5234);
xnor U5419 (N_5419,N_5379,N_5213);
or U5420 (N_5420,N_5315,N_5239);
or U5421 (N_5421,N_5380,N_5241);
nor U5422 (N_5422,N_5348,N_5321);
or U5423 (N_5423,N_5215,N_5223);
and U5424 (N_5424,N_5332,N_5334);
nor U5425 (N_5425,N_5372,N_5391);
xnor U5426 (N_5426,N_5283,N_5351);
or U5427 (N_5427,N_5298,N_5237);
nand U5428 (N_5428,N_5277,N_5358);
xor U5429 (N_5429,N_5388,N_5207);
xor U5430 (N_5430,N_5296,N_5312);
nor U5431 (N_5431,N_5291,N_5361);
nor U5432 (N_5432,N_5255,N_5273);
or U5433 (N_5433,N_5328,N_5337);
nor U5434 (N_5434,N_5246,N_5227);
nor U5435 (N_5435,N_5385,N_5233);
or U5436 (N_5436,N_5275,N_5397);
xor U5437 (N_5437,N_5357,N_5330);
or U5438 (N_5438,N_5209,N_5220);
nand U5439 (N_5439,N_5205,N_5384);
and U5440 (N_5440,N_5272,N_5386);
and U5441 (N_5441,N_5243,N_5247);
and U5442 (N_5442,N_5200,N_5300);
xnor U5443 (N_5443,N_5210,N_5342);
or U5444 (N_5444,N_5232,N_5263);
nor U5445 (N_5445,N_5318,N_5353);
or U5446 (N_5446,N_5396,N_5340);
and U5447 (N_5447,N_5219,N_5375);
or U5448 (N_5448,N_5260,N_5371);
nand U5449 (N_5449,N_5324,N_5265);
or U5450 (N_5450,N_5212,N_5302);
nand U5451 (N_5451,N_5269,N_5305);
and U5452 (N_5452,N_5203,N_5383);
nor U5453 (N_5453,N_5295,N_5285);
xnor U5454 (N_5454,N_5250,N_5344);
and U5455 (N_5455,N_5377,N_5218);
xnor U5456 (N_5456,N_5313,N_5336);
nand U5457 (N_5457,N_5293,N_5240);
or U5458 (N_5458,N_5303,N_5206);
xnor U5459 (N_5459,N_5230,N_5201);
and U5460 (N_5460,N_5221,N_5238);
xnor U5461 (N_5461,N_5398,N_5235);
xnor U5462 (N_5462,N_5399,N_5297);
nand U5463 (N_5463,N_5231,N_5360);
nand U5464 (N_5464,N_5224,N_5356);
and U5465 (N_5465,N_5266,N_5267);
or U5466 (N_5466,N_5308,N_5346);
and U5467 (N_5467,N_5274,N_5217);
nor U5468 (N_5468,N_5204,N_5359);
nand U5469 (N_5469,N_5331,N_5393);
nor U5470 (N_5470,N_5279,N_5339);
nand U5471 (N_5471,N_5343,N_5363);
xnor U5472 (N_5472,N_5395,N_5365);
nand U5473 (N_5473,N_5262,N_5368);
nor U5474 (N_5474,N_5228,N_5333);
or U5475 (N_5475,N_5304,N_5325);
or U5476 (N_5476,N_5367,N_5322);
nand U5477 (N_5477,N_5362,N_5335);
nand U5478 (N_5478,N_5392,N_5211);
or U5479 (N_5479,N_5249,N_5245);
nand U5480 (N_5480,N_5376,N_5347);
or U5481 (N_5481,N_5259,N_5378);
or U5482 (N_5482,N_5225,N_5301);
nor U5483 (N_5483,N_5256,N_5299);
or U5484 (N_5484,N_5341,N_5373);
xnor U5485 (N_5485,N_5229,N_5320);
xor U5486 (N_5486,N_5248,N_5390);
nand U5487 (N_5487,N_5282,N_5366);
xor U5488 (N_5488,N_5281,N_5294);
nand U5489 (N_5489,N_5271,N_5316);
nand U5490 (N_5490,N_5394,N_5257);
and U5491 (N_5491,N_5319,N_5326);
xnor U5492 (N_5492,N_5306,N_5387);
or U5493 (N_5493,N_5280,N_5329);
and U5494 (N_5494,N_5278,N_5314);
nand U5495 (N_5495,N_5317,N_5222);
or U5496 (N_5496,N_5374,N_5202);
xor U5497 (N_5497,N_5208,N_5216);
and U5498 (N_5498,N_5270,N_5244);
or U5499 (N_5499,N_5226,N_5252);
xnor U5500 (N_5500,N_5221,N_5231);
xnor U5501 (N_5501,N_5292,N_5209);
and U5502 (N_5502,N_5363,N_5210);
and U5503 (N_5503,N_5276,N_5398);
nand U5504 (N_5504,N_5324,N_5256);
and U5505 (N_5505,N_5385,N_5336);
and U5506 (N_5506,N_5346,N_5329);
and U5507 (N_5507,N_5245,N_5390);
or U5508 (N_5508,N_5341,N_5384);
nand U5509 (N_5509,N_5267,N_5312);
nor U5510 (N_5510,N_5238,N_5285);
and U5511 (N_5511,N_5370,N_5345);
nand U5512 (N_5512,N_5378,N_5360);
or U5513 (N_5513,N_5246,N_5313);
xor U5514 (N_5514,N_5354,N_5227);
or U5515 (N_5515,N_5347,N_5250);
nand U5516 (N_5516,N_5294,N_5340);
or U5517 (N_5517,N_5212,N_5283);
nor U5518 (N_5518,N_5319,N_5232);
nand U5519 (N_5519,N_5297,N_5212);
xnor U5520 (N_5520,N_5270,N_5204);
nand U5521 (N_5521,N_5362,N_5320);
xnor U5522 (N_5522,N_5208,N_5232);
xnor U5523 (N_5523,N_5244,N_5241);
or U5524 (N_5524,N_5363,N_5275);
or U5525 (N_5525,N_5211,N_5222);
or U5526 (N_5526,N_5234,N_5380);
nor U5527 (N_5527,N_5353,N_5350);
or U5528 (N_5528,N_5236,N_5230);
and U5529 (N_5529,N_5208,N_5229);
or U5530 (N_5530,N_5208,N_5381);
nand U5531 (N_5531,N_5308,N_5266);
or U5532 (N_5532,N_5247,N_5335);
nor U5533 (N_5533,N_5356,N_5319);
or U5534 (N_5534,N_5224,N_5293);
nand U5535 (N_5535,N_5272,N_5259);
nand U5536 (N_5536,N_5394,N_5336);
nand U5537 (N_5537,N_5311,N_5393);
and U5538 (N_5538,N_5280,N_5258);
nand U5539 (N_5539,N_5206,N_5371);
nor U5540 (N_5540,N_5374,N_5227);
nor U5541 (N_5541,N_5355,N_5283);
and U5542 (N_5542,N_5295,N_5350);
or U5543 (N_5543,N_5308,N_5254);
nor U5544 (N_5544,N_5288,N_5342);
or U5545 (N_5545,N_5255,N_5318);
xnor U5546 (N_5546,N_5270,N_5389);
nand U5547 (N_5547,N_5280,N_5307);
and U5548 (N_5548,N_5229,N_5308);
or U5549 (N_5549,N_5314,N_5237);
xor U5550 (N_5550,N_5330,N_5273);
nor U5551 (N_5551,N_5340,N_5275);
xor U5552 (N_5552,N_5345,N_5331);
nand U5553 (N_5553,N_5337,N_5290);
xor U5554 (N_5554,N_5290,N_5207);
or U5555 (N_5555,N_5340,N_5214);
or U5556 (N_5556,N_5345,N_5321);
or U5557 (N_5557,N_5279,N_5289);
nor U5558 (N_5558,N_5360,N_5317);
or U5559 (N_5559,N_5240,N_5311);
nor U5560 (N_5560,N_5357,N_5221);
xor U5561 (N_5561,N_5337,N_5348);
nor U5562 (N_5562,N_5298,N_5342);
and U5563 (N_5563,N_5242,N_5224);
xor U5564 (N_5564,N_5381,N_5398);
nor U5565 (N_5565,N_5366,N_5269);
or U5566 (N_5566,N_5307,N_5237);
or U5567 (N_5567,N_5341,N_5215);
nor U5568 (N_5568,N_5380,N_5310);
xnor U5569 (N_5569,N_5212,N_5323);
xor U5570 (N_5570,N_5233,N_5264);
xor U5571 (N_5571,N_5230,N_5227);
nand U5572 (N_5572,N_5325,N_5239);
nand U5573 (N_5573,N_5289,N_5379);
nor U5574 (N_5574,N_5204,N_5342);
nand U5575 (N_5575,N_5325,N_5326);
nand U5576 (N_5576,N_5278,N_5297);
xnor U5577 (N_5577,N_5383,N_5387);
and U5578 (N_5578,N_5258,N_5345);
or U5579 (N_5579,N_5356,N_5359);
nand U5580 (N_5580,N_5335,N_5220);
and U5581 (N_5581,N_5219,N_5222);
nand U5582 (N_5582,N_5295,N_5356);
xor U5583 (N_5583,N_5211,N_5225);
nand U5584 (N_5584,N_5386,N_5299);
or U5585 (N_5585,N_5363,N_5319);
or U5586 (N_5586,N_5208,N_5222);
nand U5587 (N_5587,N_5206,N_5276);
nand U5588 (N_5588,N_5259,N_5265);
and U5589 (N_5589,N_5390,N_5304);
xnor U5590 (N_5590,N_5369,N_5234);
nand U5591 (N_5591,N_5373,N_5258);
nor U5592 (N_5592,N_5213,N_5334);
nand U5593 (N_5593,N_5230,N_5328);
and U5594 (N_5594,N_5222,N_5264);
and U5595 (N_5595,N_5377,N_5245);
nor U5596 (N_5596,N_5348,N_5242);
xor U5597 (N_5597,N_5332,N_5389);
nor U5598 (N_5598,N_5270,N_5351);
nor U5599 (N_5599,N_5229,N_5316);
nor U5600 (N_5600,N_5455,N_5558);
and U5601 (N_5601,N_5509,N_5561);
and U5602 (N_5602,N_5546,N_5465);
xnor U5603 (N_5603,N_5550,N_5543);
xor U5604 (N_5604,N_5457,N_5479);
nand U5605 (N_5605,N_5521,N_5427);
nand U5606 (N_5606,N_5433,N_5447);
nand U5607 (N_5607,N_5437,N_5575);
nor U5608 (N_5608,N_5483,N_5404);
nand U5609 (N_5609,N_5421,N_5517);
nand U5610 (N_5610,N_5554,N_5560);
nor U5611 (N_5611,N_5400,N_5444);
nand U5612 (N_5612,N_5480,N_5574);
nor U5613 (N_5613,N_5488,N_5428);
nor U5614 (N_5614,N_5467,N_5583);
nor U5615 (N_5615,N_5458,N_5571);
nor U5616 (N_5616,N_5596,N_5473);
and U5617 (N_5617,N_5470,N_5584);
or U5618 (N_5618,N_5541,N_5585);
or U5619 (N_5619,N_5476,N_5530);
xnor U5620 (N_5620,N_5567,N_5401);
nor U5621 (N_5621,N_5409,N_5524);
xnor U5622 (N_5622,N_5454,N_5462);
or U5623 (N_5623,N_5557,N_5415);
xnor U5624 (N_5624,N_5597,N_5406);
nand U5625 (N_5625,N_5526,N_5496);
and U5626 (N_5626,N_5568,N_5474);
nand U5627 (N_5627,N_5591,N_5592);
nor U5628 (N_5628,N_5424,N_5579);
xor U5629 (N_5629,N_5547,N_5408);
nand U5630 (N_5630,N_5414,N_5477);
nand U5631 (N_5631,N_5525,N_5410);
and U5632 (N_5632,N_5553,N_5468);
nor U5633 (N_5633,N_5441,N_5412);
xnor U5634 (N_5634,N_5580,N_5593);
and U5635 (N_5635,N_5495,N_5538);
and U5636 (N_5636,N_5403,N_5508);
nor U5637 (N_5637,N_5570,N_5576);
xor U5638 (N_5638,N_5563,N_5544);
or U5639 (N_5639,N_5586,N_5481);
xor U5640 (N_5640,N_5516,N_5569);
nor U5641 (N_5641,N_5535,N_5588);
and U5642 (N_5642,N_5402,N_5599);
and U5643 (N_5643,N_5528,N_5518);
xor U5644 (N_5644,N_5595,N_5534);
xnor U5645 (N_5645,N_5461,N_5527);
or U5646 (N_5646,N_5456,N_5514);
and U5647 (N_5647,N_5502,N_5519);
nor U5648 (N_5648,N_5464,N_5411);
and U5649 (N_5649,N_5540,N_5449);
or U5650 (N_5650,N_5416,N_5469);
or U5651 (N_5651,N_5536,N_5426);
and U5652 (N_5652,N_5503,N_5513);
and U5653 (N_5653,N_5445,N_5434);
xor U5654 (N_5654,N_5450,N_5548);
nand U5655 (N_5655,N_5598,N_5432);
nor U5656 (N_5656,N_5566,N_5435);
nor U5657 (N_5657,N_5531,N_5451);
nor U5658 (N_5658,N_5523,N_5407);
or U5659 (N_5659,N_5499,N_5505);
nand U5660 (N_5660,N_5562,N_5556);
nor U5661 (N_5661,N_5493,N_5590);
or U5662 (N_5662,N_5551,N_5439);
and U5663 (N_5663,N_5511,N_5417);
nand U5664 (N_5664,N_5565,N_5506);
nor U5665 (N_5665,N_5478,N_5504);
and U5666 (N_5666,N_5436,N_5448);
nand U5667 (N_5667,N_5491,N_5472);
xor U5668 (N_5668,N_5405,N_5532);
nor U5669 (N_5669,N_5498,N_5440);
nand U5670 (N_5670,N_5510,N_5552);
xor U5671 (N_5671,N_5520,N_5475);
nor U5672 (N_5672,N_5539,N_5581);
xor U5673 (N_5673,N_5484,N_5522);
and U5674 (N_5674,N_5471,N_5438);
or U5675 (N_5675,N_5431,N_5494);
nand U5676 (N_5676,N_5422,N_5559);
or U5677 (N_5677,N_5549,N_5490);
or U5678 (N_5678,N_5497,N_5446);
or U5679 (N_5679,N_5459,N_5529);
nor U5680 (N_5680,N_5442,N_5545);
or U5681 (N_5681,N_5564,N_5485);
or U5682 (N_5682,N_5453,N_5418);
xor U5683 (N_5683,N_5413,N_5466);
nand U5684 (N_5684,N_5429,N_5430);
xor U5685 (N_5685,N_5452,N_5537);
and U5686 (N_5686,N_5589,N_5515);
and U5687 (N_5687,N_5501,N_5463);
nand U5688 (N_5688,N_5507,N_5533);
and U5689 (N_5689,N_5542,N_5486);
and U5690 (N_5690,N_5573,N_5578);
xor U5691 (N_5691,N_5420,N_5419);
or U5692 (N_5692,N_5577,N_5500);
and U5693 (N_5693,N_5594,N_5512);
and U5694 (N_5694,N_5460,N_5587);
xnor U5695 (N_5695,N_5443,N_5489);
xnor U5696 (N_5696,N_5425,N_5582);
nand U5697 (N_5697,N_5492,N_5482);
nor U5698 (N_5698,N_5423,N_5572);
xor U5699 (N_5699,N_5487,N_5555);
nor U5700 (N_5700,N_5528,N_5496);
xor U5701 (N_5701,N_5528,N_5588);
or U5702 (N_5702,N_5535,N_5447);
and U5703 (N_5703,N_5480,N_5544);
nand U5704 (N_5704,N_5524,N_5533);
xnor U5705 (N_5705,N_5547,N_5431);
nor U5706 (N_5706,N_5511,N_5524);
xnor U5707 (N_5707,N_5441,N_5547);
nand U5708 (N_5708,N_5520,N_5497);
nand U5709 (N_5709,N_5493,N_5448);
xnor U5710 (N_5710,N_5408,N_5598);
nand U5711 (N_5711,N_5531,N_5548);
nand U5712 (N_5712,N_5426,N_5590);
xor U5713 (N_5713,N_5444,N_5452);
nand U5714 (N_5714,N_5528,N_5413);
nor U5715 (N_5715,N_5439,N_5400);
or U5716 (N_5716,N_5508,N_5570);
nand U5717 (N_5717,N_5517,N_5427);
nand U5718 (N_5718,N_5460,N_5442);
nand U5719 (N_5719,N_5465,N_5556);
and U5720 (N_5720,N_5588,N_5444);
nor U5721 (N_5721,N_5469,N_5453);
xnor U5722 (N_5722,N_5524,N_5529);
nor U5723 (N_5723,N_5577,N_5587);
or U5724 (N_5724,N_5468,N_5428);
and U5725 (N_5725,N_5538,N_5544);
nand U5726 (N_5726,N_5542,N_5445);
xor U5727 (N_5727,N_5431,N_5532);
nand U5728 (N_5728,N_5488,N_5582);
nand U5729 (N_5729,N_5474,N_5571);
xnor U5730 (N_5730,N_5539,N_5470);
or U5731 (N_5731,N_5525,N_5426);
nor U5732 (N_5732,N_5584,N_5525);
or U5733 (N_5733,N_5423,N_5403);
nor U5734 (N_5734,N_5551,N_5584);
xnor U5735 (N_5735,N_5530,N_5527);
or U5736 (N_5736,N_5569,N_5526);
nor U5737 (N_5737,N_5474,N_5468);
and U5738 (N_5738,N_5503,N_5408);
or U5739 (N_5739,N_5428,N_5506);
xnor U5740 (N_5740,N_5553,N_5481);
nor U5741 (N_5741,N_5594,N_5414);
or U5742 (N_5742,N_5499,N_5512);
xor U5743 (N_5743,N_5484,N_5551);
xor U5744 (N_5744,N_5410,N_5464);
and U5745 (N_5745,N_5484,N_5586);
and U5746 (N_5746,N_5587,N_5571);
and U5747 (N_5747,N_5514,N_5495);
nand U5748 (N_5748,N_5581,N_5578);
nand U5749 (N_5749,N_5515,N_5556);
xor U5750 (N_5750,N_5575,N_5561);
or U5751 (N_5751,N_5471,N_5537);
nor U5752 (N_5752,N_5415,N_5544);
xor U5753 (N_5753,N_5523,N_5489);
and U5754 (N_5754,N_5567,N_5463);
nand U5755 (N_5755,N_5531,N_5513);
xor U5756 (N_5756,N_5458,N_5587);
xnor U5757 (N_5757,N_5459,N_5553);
or U5758 (N_5758,N_5440,N_5459);
nor U5759 (N_5759,N_5532,N_5577);
and U5760 (N_5760,N_5491,N_5583);
nor U5761 (N_5761,N_5448,N_5485);
and U5762 (N_5762,N_5565,N_5597);
nor U5763 (N_5763,N_5518,N_5421);
or U5764 (N_5764,N_5548,N_5436);
nand U5765 (N_5765,N_5526,N_5495);
nand U5766 (N_5766,N_5505,N_5464);
nand U5767 (N_5767,N_5433,N_5449);
xnor U5768 (N_5768,N_5421,N_5419);
xor U5769 (N_5769,N_5498,N_5580);
nand U5770 (N_5770,N_5414,N_5431);
nor U5771 (N_5771,N_5582,N_5555);
xor U5772 (N_5772,N_5425,N_5423);
nor U5773 (N_5773,N_5585,N_5457);
nor U5774 (N_5774,N_5532,N_5596);
and U5775 (N_5775,N_5509,N_5539);
or U5776 (N_5776,N_5594,N_5530);
or U5777 (N_5777,N_5486,N_5410);
or U5778 (N_5778,N_5494,N_5502);
xor U5779 (N_5779,N_5529,N_5487);
xor U5780 (N_5780,N_5475,N_5420);
or U5781 (N_5781,N_5512,N_5482);
xor U5782 (N_5782,N_5400,N_5561);
or U5783 (N_5783,N_5425,N_5571);
nor U5784 (N_5784,N_5521,N_5532);
or U5785 (N_5785,N_5457,N_5456);
xnor U5786 (N_5786,N_5448,N_5494);
and U5787 (N_5787,N_5404,N_5505);
nor U5788 (N_5788,N_5595,N_5561);
xnor U5789 (N_5789,N_5485,N_5595);
nand U5790 (N_5790,N_5439,N_5576);
or U5791 (N_5791,N_5481,N_5408);
or U5792 (N_5792,N_5529,N_5561);
xor U5793 (N_5793,N_5405,N_5439);
xor U5794 (N_5794,N_5486,N_5473);
nor U5795 (N_5795,N_5467,N_5559);
nor U5796 (N_5796,N_5526,N_5475);
nand U5797 (N_5797,N_5405,N_5538);
and U5798 (N_5798,N_5578,N_5445);
and U5799 (N_5799,N_5483,N_5505);
xnor U5800 (N_5800,N_5631,N_5740);
nor U5801 (N_5801,N_5684,N_5669);
xor U5802 (N_5802,N_5626,N_5788);
nor U5803 (N_5803,N_5752,N_5687);
nand U5804 (N_5804,N_5686,N_5668);
nand U5805 (N_5805,N_5710,N_5660);
nor U5806 (N_5806,N_5758,N_5612);
or U5807 (N_5807,N_5798,N_5627);
and U5808 (N_5808,N_5601,N_5779);
xnor U5809 (N_5809,N_5621,N_5782);
xnor U5810 (N_5810,N_5716,N_5711);
nand U5811 (N_5811,N_5655,N_5757);
xnor U5812 (N_5812,N_5776,N_5677);
or U5813 (N_5813,N_5754,N_5661);
nand U5814 (N_5814,N_5709,N_5731);
nand U5815 (N_5815,N_5727,N_5733);
and U5816 (N_5816,N_5653,N_5694);
xor U5817 (N_5817,N_5795,N_5648);
or U5818 (N_5818,N_5741,N_5714);
or U5819 (N_5819,N_5768,N_5794);
nand U5820 (N_5820,N_5652,N_5633);
nand U5821 (N_5821,N_5718,N_5778);
nor U5822 (N_5822,N_5624,N_5753);
xnor U5823 (N_5823,N_5755,N_5681);
or U5824 (N_5824,N_5750,N_5725);
or U5825 (N_5825,N_5712,N_5766);
nand U5826 (N_5826,N_5691,N_5748);
xnor U5827 (N_5827,N_5719,N_5615);
and U5828 (N_5828,N_5680,N_5708);
nand U5829 (N_5829,N_5673,N_5721);
and U5830 (N_5830,N_5724,N_5628);
nor U5831 (N_5831,N_5722,N_5701);
xor U5832 (N_5832,N_5606,N_5796);
or U5833 (N_5833,N_5780,N_5616);
or U5834 (N_5834,N_5678,N_5646);
nand U5835 (N_5835,N_5785,N_5697);
and U5836 (N_5836,N_5705,N_5634);
nor U5837 (N_5837,N_5743,N_5690);
xor U5838 (N_5838,N_5702,N_5650);
or U5839 (N_5839,N_5645,N_5742);
nand U5840 (N_5840,N_5617,N_5632);
or U5841 (N_5841,N_5786,N_5734);
nand U5842 (N_5842,N_5608,N_5699);
and U5843 (N_5843,N_5791,N_5771);
and U5844 (N_5844,N_5656,N_5738);
and U5845 (N_5845,N_5641,N_5670);
and U5846 (N_5846,N_5777,N_5797);
or U5847 (N_5847,N_5792,N_5689);
nor U5848 (N_5848,N_5720,N_5671);
nand U5849 (N_5849,N_5623,N_5726);
or U5850 (N_5850,N_5762,N_5605);
xor U5851 (N_5851,N_5604,N_5676);
or U5852 (N_5852,N_5625,N_5602);
and U5853 (N_5853,N_5629,N_5775);
nor U5854 (N_5854,N_5774,N_5630);
nor U5855 (N_5855,N_5763,N_5644);
xor U5856 (N_5856,N_5772,N_5667);
and U5857 (N_5857,N_5713,N_5735);
and U5858 (N_5858,N_5639,N_5603);
nor U5859 (N_5859,N_5703,N_5751);
nand U5860 (N_5860,N_5783,N_5654);
nor U5861 (N_5861,N_5736,N_5643);
nor U5862 (N_5862,N_5695,N_5679);
and U5863 (N_5863,N_5651,N_5730);
xor U5864 (N_5864,N_5787,N_5642);
and U5865 (N_5865,N_5773,N_5607);
nand U5866 (N_5866,N_5657,N_5662);
nand U5867 (N_5867,N_5760,N_5715);
or U5868 (N_5868,N_5672,N_5683);
and U5869 (N_5869,N_5620,N_5622);
or U5870 (N_5870,N_5746,N_5682);
xnor U5871 (N_5871,N_5728,N_5614);
or U5872 (N_5872,N_5675,N_5636);
xnor U5873 (N_5873,N_5613,N_5663);
nor U5874 (N_5874,N_5619,N_5756);
xnor U5875 (N_5875,N_5764,N_5693);
and U5876 (N_5876,N_5658,N_5781);
xor U5877 (N_5877,N_5640,N_5732);
xor U5878 (N_5878,N_5737,N_5749);
or U5879 (N_5879,N_5745,N_5692);
and U5880 (N_5880,N_5717,N_5793);
and U5881 (N_5881,N_5609,N_5784);
nor U5882 (N_5882,N_5665,N_5739);
nor U5883 (N_5883,N_5666,N_5649);
and U5884 (N_5884,N_5659,N_5765);
nand U5885 (N_5885,N_5638,N_5767);
or U5886 (N_5886,N_5759,N_5729);
nand U5887 (N_5887,N_5664,N_5685);
and U5888 (N_5888,N_5610,N_5700);
xnor U5889 (N_5889,N_5789,N_5723);
nand U5890 (N_5890,N_5790,N_5704);
xor U5891 (N_5891,N_5647,N_5674);
xnor U5892 (N_5892,N_5744,N_5600);
nand U5893 (N_5893,N_5747,N_5618);
nand U5894 (N_5894,N_5698,N_5688);
xnor U5895 (N_5895,N_5611,N_5706);
xnor U5896 (N_5896,N_5769,N_5770);
nand U5897 (N_5897,N_5761,N_5637);
nor U5898 (N_5898,N_5707,N_5696);
nand U5899 (N_5899,N_5635,N_5799);
and U5900 (N_5900,N_5610,N_5634);
xnor U5901 (N_5901,N_5788,N_5675);
nor U5902 (N_5902,N_5694,N_5664);
and U5903 (N_5903,N_5647,N_5735);
xnor U5904 (N_5904,N_5770,N_5679);
or U5905 (N_5905,N_5670,N_5654);
xor U5906 (N_5906,N_5633,N_5662);
or U5907 (N_5907,N_5797,N_5705);
nor U5908 (N_5908,N_5685,N_5780);
xor U5909 (N_5909,N_5711,N_5654);
and U5910 (N_5910,N_5697,N_5692);
xor U5911 (N_5911,N_5798,N_5665);
and U5912 (N_5912,N_5660,N_5761);
or U5913 (N_5913,N_5710,N_5706);
and U5914 (N_5914,N_5622,N_5608);
xor U5915 (N_5915,N_5710,N_5653);
xor U5916 (N_5916,N_5712,N_5784);
or U5917 (N_5917,N_5728,N_5769);
or U5918 (N_5918,N_5740,N_5608);
nand U5919 (N_5919,N_5628,N_5765);
and U5920 (N_5920,N_5746,N_5749);
xnor U5921 (N_5921,N_5615,N_5728);
or U5922 (N_5922,N_5751,N_5778);
nand U5923 (N_5923,N_5742,N_5736);
xnor U5924 (N_5924,N_5657,N_5785);
or U5925 (N_5925,N_5614,N_5787);
and U5926 (N_5926,N_5623,N_5714);
and U5927 (N_5927,N_5653,N_5716);
or U5928 (N_5928,N_5686,N_5743);
or U5929 (N_5929,N_5610,N_5702);
and U5930 (N_5930,N_5672,N_5649);
nor U5931 (N_5931,N_5795,N_5714);
nor U5932 (N_5932,N_5737,N_5705);
nor U5933 (N_5933,N_5724,N_5723);
or U5934 (N_5934,N_5622,N_5742);
nand U5935 (N_5935,N_5729,N_5702);
nand U5936 (N_5936,N_5717,N_5600);
or U5937 (N_5937,N_5708,N_5718);
and U5938 (N_5938,N_5738,N_5681);
or U5939 (N_5939,N_5752,N_5644);
xnor U5940 (N_5940,N_5677,N_5756);
and U5941 (N_5941,N_5763,N_5677);
or U5942 (N_5942,N_5726,N_5765);
and U5943 (N_5943,N_5676,N_5771);
nor U5944 (N_5944,N_5636,N_5688);
nor U5945 (N_5945,N_5793,N_5633);
nor U5946 (N_5946,N_5777,N_5626);
nand U5947 (N_5947,N_5610,N_5686);
or U5948 (N_5948,N_5653,N_5736);
nand U5949 (N_5949,N_5629,N_5615);
or U5950 (N_5950,N_5711,N_5796);
nand U5951 (N_5951,N_5706,N_5737);
xnor U5952 (N_5952,N_5772,N_5792);
nand U5953 (N_5953,N_5601,N_5697);
and U5954 (N_5954,N_5653,N_5745);
and U5955 (N_5955,N_5793,N_5738);
xor U5956 (N_5956,N_5793,N_5799);
nand U5957 (N_5957,N_5736,N_5669);
nand U5958 (N_5958,N_5759,N_5624);
nor U5959 (N_5959,N_5600,N_5614);
xnor U5960 (N_5960,N_5782,N_5676);
nand U5961 (N_5961,N_5742,N_5719);
nand U5962 (N_5962,N_5625,N_5662);
nor U5963 (N_5963,N_5636,N_5779);
and U5964 (N_5964,N_5618,N_5705);
nand U5965 (N_5965,N_5675,N_5621);
nor U5966 (N_5966,N_5744,N_5710);
and U5967 (N_5967,N_5603,N_5621);
xor U5968 (N_5968,N_5771,N_5672);
nor U5969 (N_5969,N_5702,N_5726);
or U5970 (N_5970,N_5665,N_5611);
or U5971 (N_5971,N_5672,N_5775);
and U5972 (N_5972,N_5649,N_5734);
or U5973 (N_5973,N_5617,N_5618);
nor U5974 (N_5974,N_5688,N_5743);
or U5975 (N_5975,N_5719,N_5681);
nor U5976 (N_5976,N_5633,N_5731);
xnor U5977 (N_5977,N_5757,N_5607);
and U5978 (N_5978,N_5724,N_5771);
xnor U5979 (N_5979,N_5757,N_5723);
and U5980 (N_5980,N_5743,N_5631);
and U5981 (N_5981,N_5765,N_5703);
or U5982 (N_5982,N_5675,N_5745);
xnor U5983 (N_5983,N_5625,N_5710);
xnor U5984 (N_5984,N_5676,N_5704);
nor U5985 (N_5985,N_5758,N_5602);
and U5986 (N_5986,N_5668,N_5780);
nand U5987 (N_5987,N_5627,N_5675);
and U5988 (N_5988,N_5666,N_5781);
nor U5989 (N_5989,N_5665,N_5634);
nand U5990 (N_5990,N_5774,N_5605);
nand U5991 (N_5991,N_5611,N_5612);
xnor U5992 (N_5992,N_5661,N_5694);
nand U5993 (N_5993,N_5798,N_5671);
and U5994 (N_5994,N_5797,N_5742);
nor U5995 (N_5995,N_5702,N_5684);
nor U5996 (N_5996,N_5726,N_5614);
xnor U5997 (N_5997,N_5680,N_5648);
or U5998 (N_5998,N_5751,N_5632);
or U5999 (N_5999,N_5692,N_5612);
nor U6000 (N_6000,N_5957,N_5906);
nor U6001 (N_6001,N_5827,N_5968);
or U6002 (N_6002,N_5850,N_5887);
xor U6003 (N_6003,N_5839,N_5872);
nor U6004 (N_6004,N_5944,N_5992);
nand U6005 (N_6005,N_5825,N_5803);
xnor U6006 (N_6006,N_5878,N_5978);
nand U6007 (N_6007,N_5970,N_5877);
nand U6008 (N_6008,N_5858,N_5908);
xor U6009 (N_6009,N_5880,N_5816);
and U6010 (N_6010,N_5929,N_5910);
or U6011 (N_6011,N_5871,N_5949);
nand U6012 (N_6012,N_5857,N_5826);
nand U6013 (N_6013,N_5817,N_5930);
nand U6014 (N_6014,N_5917,N_5953);
xor U6015 (N_6015,N_5864,N_5937);
or U6016 (N_6016,N_5875,N_5855);
nor U6017 (N_6017,N_5959,N_5915);
and U6018 (N_6018,N_5940,N_5832);
and U6019 (N_6019,N_5873,N_5868);
nor U6020 (N_6020,N_5982,N_5971);
and U6021 (N_6021,N_5923,N_5942);
xor U6022 (N_6022,N_5810,N_5834);
nor U6023 (N_6023,N_5984,N_5919);
nor U6024 (N_6024,N_5932,N_5913);
and U6025 (N_6025,N_5933,N_5936);
or U6026 (N_6026,N_5896,N_5876);
and U6027 (N_6027,N_5842,N_5965);
nor U6028 (N_6028,N_5861,N_5838);
and U6029 (N_6029,N_5852,N_5867);
or U6030 (N_6030,N_5843,N_5883);
nand U6031 (N_6031,N_5831,N_5829);
nor U6032 (N_6032,N_5946,N_5980);
nor U6033 (N_6033,N_5954,N_5907);
xnor U6034 (N_6034,N_5848,N_5931);
nand U6035 (N_6035,N_5987,N_5830);
nor U6036 (N_6036,N_5902,N_5859);
xnor U6037 (N_6037,N_5952,N_5879);
nand U6038 (N_6038,N_5962,N_5882);
or U6039 (N_6039,N_5837,N_5967);
and U6040 (N_6040,N_5836,N_5988);
xor U6041 (N_6041,N_5972,N_5966);
nand U6042 (N_6042,N_5922,N_5976);
nand U6043 (N_6043,N_5812,N_5860);
or U6044 (N_6044,N_5844,N_5921);
xor U6045 (N_6045,N_5806,N_5963);
nand U6046 (N_6046,N_5820,N_5846);
nor U6047 (N_6047,N_5991,N_5822);
nor U6048 (N_6048,N_5893,N_5849);
and U6049 (N_6049,N_5890,N_5847);
or U6050 (N_6050,N_5851,N_5905);
xnor U6051 (N_6051,N_5808,N_5979);
xnor U6052 (N_6052,N_5989,N_5969);
nor U6053 (N_6053,N_5824,N_5863);
or U6054 (N_6054,N_5918,N_5909);
or U6055 (N_6055,N_5973,N_5956);
nand U6056 (N_6056,N_5948,N_5994);
nor U6057 (N_6057,N_5927,N_5993);
nor U6058 (N_6058,N_5961,N_5925);
and U6059 (N_6059,N_5802,N_5951);
or U6060 (N_6060,N_5960,N_5955);
xor U6061 (N_6061,N_5815,N_5828);
nand U6062 (N_6062,N_5914,N_5841);
nor U6063 (N_6063,N_5935,N_5904);
nand U6064 (N_6064,N_5939,N_5894);
or U6065 (N_6065,N_5801,N_5854);
or U6066 (N_6066,N_5881,N_5945);
xor U6067 (N_6067,N_5998,N_5821);
xor U6068 (N_6068,N_5974,N_5884);
xor U6069 (N_6069,N_5856,N_5862);
and U6070 (N_6070,N_5888,N_5977);
and U6071 (N_6071,N_5809,N_5813);
or U6072 (N_6072,N_5901,N_5840);
xor U6073 (N_6073,N_5985,N_5804);
xnor U6074 (N_6074,N_5920,N_5981);
xor U6075 (N_6075,N_5912,N_5916);
nand U6076 (N_6076,N_5995,N_5892);
nor U6077 (N_6077,N_5990,N_5958);
xnor U6078 (N_6078,N_5996,N_5823);
and U6079 (N_6079,N_5866,N_5924);
nor U6080 (N_6080,N_5899,N_5835);
and U6081 (N_6081,N_5975,N_5898);
or U6082 (N_6082,N_5999,N_5964);
and U6083 (N_6083,N_5889,N_5983);
nand U6084 (N_6084,N_5947,N_5853);
nand U6085 (N_6085,N_5903,N_5865);
nand U6086 (N_6086,N_5986,N_5934);
xor U6087 (N_6087,N_5870,N_5805);
or U6088 (N_6088,N_5874,N_5997);
and U6089 (N_6089,N_5833,N_5885);
or U6090 (N_6090,N_5911,N_5926);
nor U6091 (N_6091,N_5818,N_5814);
nand U6092 (N_6092,N_5941,N_5869);
nor U6093 (N_6093,N_5811,N_5950);
and U6094 (N_6094,N_5819,N_5845);
nor U6095 (N_6095,N_5943,N_5891);
and U6096 (N_6096,N_5897,N_5807);
nand U6097 (N_6097,N_5800,N_5886);
nor U6098 (N_6098,N_5928,N_5938);
nand U6099 (N_6099,N_5900,N_5895);
nand U6100 (N_6100,N_5964,N_5931);
and U6101 (N_6101,N_5979,N_5970);
nand U6102 (N_6102,N_5963,N_5999);
or U6103 (N_6103,N_5846,N_5849);
xnor U6104 (N_6104,N_5869,N_5983);
and U6105 (N_6105,N_5818,N_5954);
nand U6106 (N_6106,N_5858,N_5984);
nor U6107 (N_6107,N_5884,N_5936);
or U6108 (N_6108,N_5958,N_5903);
nor U6109 (N_6109,N_5843,N_5861);
nor U6110 (N_6110,N_5914,N_5868);
nor U6111 (N_6111,N_5880,N_5841);
or U6112 (N_6112,N_5929,N_5976);
and U6113 (N_6113,N_5988,N_5831);
nor U6114 (N_6114,N_5830,N_5861);
or U6115 (N_6115,N_5934,N_5973);
or U6116 (N_6116,N_5952,N_5863);
xnor U6117 (N_6117,N_5814,N_5962);
or U6118 (N_6118,N_5971,N_5892);
nor U6119 (N_6119,N_5831,N_5889);
or U6120 (N_6120,N_5896,N_5975);
nand U6121 (N_6121,N_5925,N_5880);
or U6122 (N_6122,N_5871,N_5965);
nor U6123 (N_6123,N_5968,N_5849);
and U6124 (N_6124,N_5856,N_5886);
and U6125 (N_6125,N_5939,N_5876);
and U6126 (N_6126,N_5894,N_5944);
or U6127 (N_6127,N_5975,N_5845);
xnor U6128 (N_6128,N_5818,N_5901);
or U6129 (N_6129,N_5864,N_5834);
xor U6130 (N_6130,N_5979,N_5947);
nor U6131 (N_6131,N_5854,N_5947);
nand U6132 (N_6132,N_5994,N_5863);
and U6133 (N_6133,N_5889,N_5975);
and U6134 (N_6134,N_5984,N_5830);
or U6135 (N_6135,N_5862,N_5994);
nand U6136 (N_6136,N_5976,N_5982);
and U6137 (N_6137,N_5942,N_5913);
nor U6138 (N_6138,N_5945,N_5871);
xor U6139 (N_6139,N_5917,N_5913);
nand U6140 (N_6140,N_5973,N_5802);
nor U6141 (N_6141,N_5996,N_5999);
or U6142 (N_6142,N_5842,N_5900);
nor U6143 (N_6143,N_5998,N_5948);
nand U6144 (N_6144,N_5882,N_5827);
and U6145 (N_6145,N_5862,N_5948);
nand U6146 (N_6146,N_5819,N_5841);
and U6147 (N_6147,N_5981,N_5929);
nor U6148 (N_6148,N_5854,N_5868);
and U6149 (N_6149,N_5895,N_5903);
nand U6150 (N_6150,N_5983,N_5964);
xor U6151 (N_6151,N_5845,N_5997);
and U6152 (N_6152,N_5919,N_5815);
or U6153 (N_6153,N_5952,N_5956);
nand U6154 (N_6154,N_5905,N_5800);
nand U6155 (N_6155,N_5860,N_5926);
nor U6156 (N_6156,N_5915,N_5840);
xor U6157 (N_6157,N_5888,N_5928);
or U6158 (N_6158,N_5833,N_5990);
xor U6159 (N_6159,N_5860,N_5976);
xnor U6160 (N_6160,N_5835,N_5840);
and U6161 (N_6161,N_5957,N_5881);
or U6162 (N_6162,N_5860,N_5936);
and U6163 (N_6163,N_5844,N_5882);
nand U6164 (N_6164,N_5903,N_5917);
and U6165 (N_6165,N_5858,N_5842);
xnor U6166 (N_6166,N_5898,N_5879);
nand U6167 (N_6167,N_5988,N_5983);
xnor U6168 (N_6168,N_5907,N_5897);
xor U6169 (N_6169,N_5987,N_5808);
xnor U6170 (N_6170,N_5838,N_5824);
and U6171 (N_6171,N_5984,N_5814);
or U6172 (N_6172,N_5946,N_5990);
xor U6173 (N_6173,N_5964,N_5970);
or U6174 (N_6174,N_5952,N_5914);
nor U6175 (N_6175,N_5897,N_5848);
and U6176 (N_6176,N_5853,N_5897);
nand U6177 (N_6177,N_5824,N_5847);
xnor U6178 (N_6178,N_5912,N_5836);
nor U6179 (N_6179,N_5851,N_5817);
xnor U6180 (N_6180,N_5975,N_5861);
nand U6181 (N_6181,N_5837,N_5951);
and U6182 (N_6182,N_5894,N_5951);
xor U6183 (N_6183,N_5946,N_5873);
or U6184 (N_6184,N_5894,N_5873);
or U6185 (N_6185,N_5880,N_5909);
nand U6186 (N_6186,N_5933,N_5830);
and U6187 (N_6187,N_5921,N_5968);
nand U6188 (N_6188,N_5840,N_5974);
nor U6189 (N_6189,N_5839,N_5938);
and U6190 (N_6190,N_5824,N_5861);
nand U6191 (N_6191,N_5956,N_5852);
or U6192 (N_6192,N_5852,N_5880);
or U6193 (N_6193,N_5862,N_5958);
xor U6194 (N_6194,N_5821,N_5845);
nand U6195 (N_6195,N_5856,N_5889);
nand U6196 (N_6196,N_5891,N_5913);
xnor U6197 (N_6197,N_5967,N_5853);
xnor U6198 (N_6198,N_5975,N_5918);
nand U6199 (N_6199,N_5806,N_5938);
or U6200 (N_6200,N_6079,N_6015);
or U6201 (N_6201,N_6135,N_6088);
nor U6202 (N_6202,N_6098,N_6138);
and U6203 (N_6203,N_6169,N_6106);
and U6204 (N_6204,N_6097,N_6113);
nand U6205 (N_6205,N_6148,N_6140);
nand U6206 (N_6206,N_6174,N_6153);
xnor U6207 (N_6207,N_6134,N_6013);
xnor U6208 (N_6208,N_6066,N_6073);
nor U6209 (N_6209,N_6063,N_6028);
or U6210 (N_6210,N_6077,N_6023);
and U6211 (N_6211,N_6190,N_6195);
and U6212 (N_6212,N_6121,N_6049);
and U6213 (N_6213,N_6147,N_6046);
xor U6214 (N_6214,N_6176,N_6105);
nor U6215 (N_6215,N_6014,N_6152);
and U6216 (N_6216,N_6025,N_6196);
or U6217 (N_6217,N_6091,N_6149);
and U6218 (N_6218,N_6089,N_6166);
or U6219 (N_6219,N_6090,N_6055);
nor U6220 (N_6220,N_6050,N_6018);
nand U6221 (N_6221,N_6053,N_6067);
nor U6222 (N_6222,N_6110,N_6033);
nand U6223 (N_6223,N_6127,N_6052);
and U6224 (N_6224,N_6096,N_6158);
xnor U6225 (N_6225,N_6032,N_6144);
and U6226 (N_6226,N_6146,N_6099);
or U6227 (N_6227,N_6188,N_6094);
and U6228 (N_6228,N_6160,N_6086);
nand U6229 (N_6229,N_6056,N_6122);
nand U6230 (N_6230,N_6012,N_6080);
xor U6231 (N_6231,N_6048,N_6093);
nor U6232 (N_6232,N_6005,N_6186);
nand U6233 (N_6233,N_6156,N_6092);
or U6234 (N_6234,N_6078,N_6103);
nor U6235 (N_6235,N_6114,N_6065);
and U6236 (N_6236,N_6167,N_6154);
xor U6237 (N_6237,N_6071,N_6136);
or U6238 (N_6238,N_6031,N_6051);
and U6239 (N_6239,N_6117,N_6082);
xor U6240 (N_6240,N_6130,N_6062);
nand U6241 (N_6241,N_6026,N_6112);
or U6242 (N_6242,N_6145,N_6116);
nand U6243 (N_6243,N_6183,N_6177);
nor U6244 (N_6244,N_6139,N_6179);
xor U6245 (N_6245,N_6009,N_6192);
or U6246 (N_6246,N_6151,N_6128);
nor U6247 (N_6247,N_6197,N_6115);
xor U6248 (N_6248,N_6075,N_6059);
and U6249 (N_6249,N_6194,N_6021);
nor U6250 (N_6250,N_6161,N_6107);
nand U6251 (N_6251,N_6001,N_6104);
xor U6252 (N_6252,N_6034,N_6108);
nor U6253 (N_6253,N_6070,N_6164);
and U6254 (N_6254,N_6159,N_6058);
nor U6255 (N_6255,N_6004,N_6042);
xnor U6256 (N_6256,N_6087,N_6187);
or U6257 (N_6257,N_6168,N_6143);
or U6258 (N_6258,N_6074,N_6095);
xor U6259 (N_6259,N_6171,N_6123);
nor U6260 (N_6260,N_6100,N_6109);
and U6261 (N_6261,N_6175,N_6180);
xor U6262 (N_6262,N_6060,N_6120);
and U6263 (N_6263,N_6007,N_6006);
xnor U6264 (N_6264,N_6011,N_6173);
nor U6265 (N_6265,N_6020,N_6030);
and U6266 (N_6266,N_6081,N_6111);
and U6267 (N_6267,N_6157,N_6172);
nor U6268 (N_6268,N_6054,N_6125);
nand U6269 (N_6269,N_6185,N_6039);
xnor U6270 (N_6270,N_6170,N_6118);
nand U6271 (N_6271,N_6163,N_6017);
and U6272 (N_6272,N_6131,N_6102);
nor U6273 (N_6273,N_6044,N_6191);
xor U6274 (N_6274,N_6182,N_6178);
nor U6275 (N_6275,N_6045,N_6041);
xnor U6276 (N_6276,N_6000,N_6162);
nor U6277 (N_6277,N_6010,N_6141);
or U6278 (N_6278,N_6019,N_6069);
nor U6279 (N_6279,N_6008,N_6016);
and U6280 (N_6280,N_6198,N_6035);
xor U6281 (N_6281,N_6037,N_6129);
and U6282 (N_6282,N_6003,N_6083);
and U6283 (N_6283,N_6181,N_6085);
nand U6284 (N_6284,N_6165,N_6072);
nor U6285 (N_6285,N_6057,N_6189);
and U6286 (N_6286,N_6061,N_6047);
xnor U6287 (N_6287,N_6150,N_6038);
nand U6288 (N_6288,N_6043,N_6027);
nor U6289 (N_6289,N_6184,N_6036);
xor U6290 (N_6290,N_6126,N_6022);
nand U6291 (N_6291,N_6040,N_6119);
xor U6292 (N_6292,N_6193,N_6142);
xnor U6293 (N_6293,N_6084,N_6155);
xnor U6294 (N_6294,N_6199,N_6064);
nand U6295 (N_6295,N_6133,N_6137);
xor U6296 (N_6296,N_6132,N_6076);
or U6297 (N_6297,N_6024,N_6029);
and U6298 (N_6298,N_6124,N_6002);
or U6299 (N_6299,N_6101,N_6068);
or U6300 (N_6300,N_6152,N_6190);
nand U6301 (N_6301,N_6069,N_6129);
xor U6302 (N_6302,N_6022,N_6147);
and U6303 (N_6303,N_6170,N_6080);
nor U6304 (N_6304,N_6003,N_6037);
xnor U6305 (N_6305,N_6161,N_6053);
nor U6306 (N_6306,N_6130,N_6045);
nor U6307 (N_6307,N_6157,N_6178);
nor U6308 (N_6308,N_6097,N_6013);
and U6309 (N_6309,N_6012,N_6139);
or U6310 (N_6310,N_6052,N_6019);
or U6311 (N_6311,N_6160,N_6132);
nand U6312 (N_6312,N_6000,N_6152);
xnor U6313 (N_6313,N_6153,N_6125);
nor U6314 (N_6314,N_6007,N_6112);
xor U6315 (N_6315,N_6181,N_6098);
or U6316 (N_6316,N_6001,N_6062);
or U6317 (N_6317,N_6142,N_6132);
nand U6318 (N_6318,N_6076,N_6005);
nand U6319 (N_6319,N_6144,N_6183);
or U6320 (N_6320,N_6004,N_6011);
xnor U6321 (N_6321,N_6182,N_6091);
xor U6322 (N_6322,N_6104,N_6164);
xnor U6323 (N_6323,N_6116,N_6136);
nor U6324 (N_6324,N_6009,N_6054);
and U6325 (N_6325,N_6151,N_6058);
xnor U6326 (N_6326,N_6029,N_6107);
or U6327 (N_6327,N_6077,N_6144);
and U6328 (N_6328,N_6011,N_6191);
nand U6329 (N_6329,N_6144,N_6033);
nand U6330 (N_6330,N_6169,N_6069);
or U6331 (N_6331,N_6198,N_6091);
xor U6332 (N_6332,N_6100,N_6133);
xnor U6333 (N_6333,N_6180,N_6088);
or U6334 (N_6334,N_6046,N_6112);
xor U6335 (N_6335,N_6038,N_6081);
or U6336 (N_6336,N_6011,N_6036);
and U6337 (N_6337,N_6076,N_6168);
nor U6338 (N_6338,N_6022,N_6075);
or U6339 (N_6339,N_6136,N_6093);
nand U6340 (N_6340,N_6125,N_6061);
nor U6341 (N_6341,N_6113,N_6063);
and U6342 (N_6342,N_6009,N_6098);
nand U6343 (N_6343,N_6024,N_6003);
xor U6344 (N_6344,N_6175,N_6130);
xor U6345 (N_6345,N_6025,N_6179);
nand U6346 (N_6346,N_6036,N_6165);
xor U6347 (N_6347,N_6174,N_6082);
nand U6348 (N_6348,N_6125,N_6157);
nor U6349 (N_6349,N_6075,N_6183);
xnor U6350 (N_6350,N_6086,N_6083);
and U6351 (N_6351,N_6010,N_6009);
and U6352 (N_6352,N_6152,N_6066);
nand U6353 (N_6353,N_6083,N_6064);
nand U6354 (N_6354,N_6191,N_6122);
nor U6355 (N_6355,N_6088,N_6032);
and U6356 (N_6356,N_6123,N_6010);
xor U6357 (N_6357,N_6174,N_6103);
nor U6358 (N_6358,N_6143,N_6178);
or U6359 (N_6359,N_6075,N_6070);
xnor U6360 (N_6360,N_6132,N_6163);
and U6361 (N_6361,N_6091,N_6145);
xnor U6362 (N_6362,N_6120,N_6054);
nor U6363 (N_6363,N_6108,N_6083);
xor U6364 (N_6364,N_6023,N_6179);
and U6365 (N_6365,N_6008,N_6005);
or U6366 (N_6366,N_6121,N_6005);
xor U6367 (N_6367,N_6155,N_6021);
or U6368 (N_6368,N_6064,N_6172);
xor U6369 (N_6369,N_6010,N_6116);
and U6370 (N_6370,N_6029,N_6133);
nor U6371 (N_6371,N_6163,N_6130);
and U6372 (N_6372,N_6041,N_6004);
nor U6373 (N_6373,N_6066,N_6176);
and U6374 (N_6374,N_6040,N_6051);
and U6375 (N_6375,N_6057,N_6192);
nand U6376 (N_6376,N_6189,N_6156);
and U6377 (N_6377,N_6040,N_6033);
nand U6378 (N_6378,N_6055,N_6199);
or U6379 (N_6379,N_6038,N_6146);
nor U6380 (N_6380,N_6004,N_6087);
xnor U6381 (N_6381,N_6153,N_6175);
xnor U6382 (N_6382,N_6025,N_6096);
nor U6383 (N_6383,N_6030,N_6014);
or U6384 (N_6384,N_6166,N_6017);
nand U6385 (N_6385,N_6057,N_6037);
nor U6386 (N_6386,N_6140,N_6176);
and U6387 (N_6387,N_6122,N_6115);
and U6388 (N_6388,N_6022,N_6150);
or U6389 (N_6389,N_6089,N_6069);
xnor U6390 (N_6390,N_6196,N_6100);
xnor U6391 (N_6391,N_6134,N_6179);
xnor U6392 (N_6392,N_6082,N_6014);
and U6393 (N_6393,N_6063,N_6006);
nor U6394 (N_6394,N_6031,N_6035);
nor U6395 (N_6395,N_6147,N_6033);
nand U6396 (N_6396,N_6063,N_6129);
or U6397 (N_6397,N_6017,N_6187);
nor U6398 (N_6398,N_6073,N_6034);
xor U6399 (N_6399,N_6199,N_6133);
xnor U6400 (N_6400,N_6300,N_6223);
nand U6401 (N_6401,N_6297,N_6206);
nor U6402 (N_6402,N_6352,N_6234);
and U6403 (N_6403,N_6256,N_6391);
and U6404 (N_6404,N_6366,N_6321);
nor U6405 (N_6405,N_6273,N_6389);
nand U6406 (N_6406,N_6235,N_6261);
nand U6407 (N_6407,N_6298,N_6302);
and U6408 (N_6408,N_6210,N_6381);
xnor U6409 (N_6409,N_6284,N_6359);
or U6410 (N_6410,N_6271,N_6283);
and U6411 (N_6411,N_6386,N_6227);
nor U6412 (N_6412,N_6328,N_6238);
or U6413 (N_6413,N_6342,N_6335);
or U6414 (N_6414,N_6334,N_6254);
xnor U6415 (N_6415,N_6351,N_6205);
nand U6416 (N_6416,N_6211,N_6353);
xnor U6417 (N_6417,N_6267,N_6365);
nor U6418 (N_6418,N_6207,N_6364);
xnor U6419 (N_6419,N_6320,N_6277);
and U6420 (N_6420,N_6348,N_6383);
nor U6421 (N_6421,N_6293,N_6220);
or U6422 (N_6422,N_6382,N_6219);
nand U6423 (N_6423,N_6215,N_6289);
and U6424 (N_6424,N_6209,N_6332);
or U6425 (N_6425,N_6248,N_6319);
nand U6426 (N_6426,N_6200,N_6322);
nor U6427 (N_6427,N_6270,N_6286);
nor U6428 (N_6428,N_6245,N_6392);
nand U6429 (N_6429,N_6253,N_6349);
xor U6430 (N_6430,N_6327,N_6340);
xnor U6431 (N_6431,N_6344,N_6380);
xnor U6432 (N_6432,N_6263,N_6295);
or U6433 (N_6433,N_6232,N_6318);
or U6434 (N_6434,N_6279,N_6280);
xnor U6435 (N_6435,N_6376,N_6323);
nand U6436 (N_6436,N_6216,N_6268);
or U6437 (N_6437,N_6208,N_6287);
nor U6438 (N_6438,N_6292,N_6251);
and U6439 (N_6439,N_6363,N_6202);
and U6440 (N_6440,N_6356,N_6372);
nand U6441 (N_6441,N_6237,N_6399);
nor U6442 (N_6442,N_6369,N_6355);
nor U6443 (N_6443,N_6246,N_6395);
nand U6444 (N_6444,N_6257,N_6324);
nand U6445 (N_6445,N_6299,N_6229);
nor U6446 (N_6446,N_6255,N_6370);
xnor U6447 (N_6447,N_6244,N_6367);
xnor U6448 (N_6448,N_6350,N_6201);
nor U6449 (N_6449,N_6228,N_6294);
or U6450 (N_6450,N_6288,N_6306);
xnor U6451 (N_6451,N_6230,N_6265);
nand U6452 (N_6452,N_6374,N_6260);
and U6453 (N_6453,N_6379,N_6213);
nand U6454 (N_6454,N_6221,N_6331);
or U6455 (N_6455,N_6338,N_6343);
and U6456 (N_6456,N_6358,N_6240);
and U6457 (N_6457,N_6275,N_6247);
and U6458 (N_6458,N_6314,N_6266);
nor U6459 (N_6459,N_6225,N_6317);
xnor U6460 (N_6460,N_6282,N_6378);
nand U6461 (N_6461,N_6347,N_6290);
xor U6462 (N_6462,N_6345,N_6249);
and U6463 (N_6463,N_6308,N_6360);
and U6464 (N_6464,N_6291,N_6337);
nand U6465 (N_6465,N_6354,N_6312);
xor U6466 (N_6466,N_6394,N_6276);
or U6467 (N_6467,N_6385,N_6224);
or U6468 (N_6468,N_6393,N_6264);
xnor U6469 (N_6469,N_6218,N_6203);
and U6470 (N_6470,N_6330,N_6250);
nor U6471 (N_6471,N_6362,N_6329);
nor U6472 (N_6472,N_6313,N_6336);
xor U6473 (N_6473,N_6285,N_6357);
nand U6474 (N_6474,N_6239,N_6231);
and U6475 (N_6475,N_6303,N_6388);
xnor U6476 (N_6476,N_6361,N_6305);
nand U6477 (N_6477,N_6346,N_6241);
and U6478 (N_6478,N_6296,N_6269);
or U6479 (N_6479,N_6242,N_6390);
nor U6480 (N_6480,N_6222,N_6278);
and U6481 (N_6481,N_6301,N_6368);
nor U6482 (N_6482,N_6204,N_6371);
and U6483 (N_6483,N_6310,N_6236);
nor U6484 (N_6484,N_6326,N_6373);
nand U6485 (N_6485,N_6384,N_6387);
and U6486 (N_6486,N_6259,N_6339);
nand U6487 (N_6487,N_6341,N_6281);
or U6488 (N_6488,N_6311,N_6375);
or U6489 (N_6489,N_6397,N_6377);
nand U6490 (N_6490,N_6316,N_6258);
or U6491 (N_6491,N_6243,N_6226);
nor U6492 (N_6492,N_6262,N_6333);
and U6493 (N_6493,N_6212,N_6272);
xnor U6494 (N_6494,N_6398,N_6274);
and U6495 (N_6495,N_6309,N_6315);
and U6496 (N_6496,N_6307,N_6214);
and U6497 (N_6497,N_6396,N_6217);
xnor U6498 (N_6498,N_6325,N_6233);
xor U6499 (N_6499,N_6252,N_6304);
nor U6500 (N_6500,N_6361,N_6381);
and U6501 (N_6501,N_6395,N_6354);
or U6502 (N_6502,N_6248,N_6212);
nand U6503 (N_6503,N_6288,N_6325);
nand U6504 (N_6504,N_6214,N_6373);
nand U6505 (N_6505,N_6291,N_6323);
nor U6506 (N_6506,N_6347,N_6233);
xnor U6507 (N_6507,N_6243,N_6354);
xor U6508 (N_6508,N_6336,N_6222);
and U6509 (N_6509,N_6285,N_6387);
xor U6510 (N_6510,N_6308,N_6330);
nand U6511 (N_6511,N_6314,N_6390);
or U6512 (N_6512,N_6351,N_6301);
xor U6513 (N_6513,N_6295,N_6292);
nor U6514 (N_6514,N_6260,N_6326);
or U6515 (N_6515,N_6358,N_6294);
or U6516 (N_6516,N_6336,N_6317);
or U6517 (N_6517,N_6300,N_6214);
and U6518 (N_6518,N_6361,N_6258);
nand U6519 (N_6519,N_6335,N_6225);
xnor U6520 (N_6520,N_6369,N_6316);
or U6521 (N_6521,N_6365,N_6346);
xnor U6522 (N_6522,N_6206,N_6285);
nand U6523 (N_6523,N_6266,N_6214);
and U6524 (N_6524,N_6399,N_6363);
and U6525 (N_6525,N_6263,N_6247);
nand U6526 (N_6526,N_6305,N_6307);
nor U6527 (N_6527,N_6232,N_6207);
nor U6528 (N_6528,N_6269,N_6267);
nand U6529 (N_6529,N_6370,N_6271);
or U6530 (N_6530,N_6328,N_6232);
nor U6531 (N_6531,N_6280,N_6276);
nand U6532 (N_6532,N_6341,N_6297);
and U6533 (N_6533,N_6224,N_6256);
xnor U6534 (N_6534,N_6322,N_6243);
nor U6535 (N_6535,N_6286,N_6336);
nand U6536 (N_6536,N_6390,N_6343);
nor U6537 (N_6537,N_6356,N_6388);
or U6538 (N_6538,N_6360,N_6247);
or U6539 (N_6539,N_6224,N_6247);
nor U6540 (N_6540,N_6335,N_6253);
xnor U6541 (N_6541,N_6275,N_6277);
or U6542 (N_6542,N_6213,N_6237);
and U6543 (N_6543,N_6330,N_6209);
and U6544 (N_6544,N_6377,N_6226);
nand U6545 (N_6545,N_6288,N_6357);
or U6546 (N_6546,N_6265,N_6393);
xor U6547 (N_6547,N_6216,N_6350);
xnor U6548 (N_6548,N_6232,N_6396);
xnor U6549 (N_6549,N_6383,N_6316);
and U6550 (N_6550,N_6221,N_6377);
nor U6551 (N_6551,N_6388,N_6396);
nor U6552 (N_6552,N_6383,N_6275);
or U6553 (N_6553,N_6351,N_6392);
or U6554 (N_6554,N_6353,N_6232);
and U6555 (N_6555,N_6260,N_6259);
xor U6556 (N_6556,N_6211,N_6292);
and U6557 (N_6557,N_6205,N_6393);
nor U6558 (N_6558,N_6389,N_6224);
nor U6559 (N_6559,N_6221,N_6367);
and U6560 (N_6560,N_6350,N_6311);
nand U6561 (N_6561,N_6384,N_6320);
and U6562 (N_6562,N_6357,N_6313);
xnor U6563 (N_6563,N_6285,N_6364);
nand U6564 (N_6564,N_6349,N_6222);
or U6565 (N_6565,N_6281,N_6398);
xor U6566 (N_6566,N_6322,N_6384);
and U6567 (N_6567,N_6398,N_6250);
nand U6568 (N_6568,N_6367,N_6263);
and U6569 (N_6569,N_6239,N_6299);
or U6570 (N_6570,N_6261,N_6266);
xor U6571 (N_6571,N_6215,N_6354);
nand U6572 (N_6572,N_6334,N_6246);
nand U6573 (N_6573,N_6373,N_6205);
nor U6574 (N_6574,N_6332,N_6243);
nor U6575 (N_6575,N_6325,N_6345);
nand U6576 (N_6576,N_6364,N_6348);
nand U6577 (N_6577,N_6390,N_6354);
nor U6578 (N_6578,N_6230,N_6314);
and U6579 (N_6579,N_6350,N_6304);
and U6580 (N_6580,N_6257,N_6262);
xor U6581 (N_6581,N_6397,N_6375);
or U6582 (N_6582,N_6342,N_6341);
nor U6583 (N_6583,N_6208,N_6376);
xnor U6584 (N_6584,N_6359,N_6324);
or U6585 (N_6585,N_6356,N_6326);
nor U6586 (N_6586,N_6229,N_6227);
nor U6587 (N_6587,N_6381,N_6273);
and U6588 (N_6588,N_6383,N_6281);
xor U6589 (N_6589,N_6238,N_6209);
xor U6590 (N_6590,N_6212,N_6252);
and U6591 (N_6591,N_6329,N_6346);
xor U6592 (N_6592,N_6362,N_6281);
nor U6593 (N_6593,N_6230,N_6386);
xnor U6594 (N_6594,N_6226,N_6288);
nor U6595 (N_6595,N_6340,N_6288);
nand U6596 (N_6596,N_6296,N_6340);
or U6597 (N_6597,N_6226,N_6255);
and U6598 (N_6598,N_6236,N_6357);
nand U6599 (N_6599,N_6283,N_6314);
nand U6600 (N_6600,N_6498,N_6460);
and U6601 (N_6601,N_6590,N_6444);
nand U6602 (N_6602,N_6584,N_6540);
xor U6603 (N_6603,N_6575,N_6457);
xor U6604 (N_6604,N_6423,N_6499);
and U6605 (N_6605,N_6555,N_6529);
nor U6606 (N_6606,N_6548,N_6491);
nor U6607 (N_6607,N_6557,N_6585);
nor U6608 (N_6608,N_6583,N_6400);
nand U6609 (N_6609,N_6580,N_6445);
xnor U6610 (N_6610,N_6416,N_6441);
xnor U6611 (N_6611,N_6438,N_6576);
nor U6612 (N_6612,N_6511,N_6595);
nand U6613 (N_6613,N_6542,N_6483);
or U6614 (N_6614,N_6593,N_6524);
or U6615 (N_6615,N_6408,N_6456);
nand U6616 (N_6616,N_6541,N_6410);
nor U6617 (N_6617,N_6481,N_6545);
or U6618 (N_6618,N_6465,N_6485);
or U6619 (N_6619,N_6428,N_6577);
nor U6620 (N_6620,N_6538,N_6547);
xnor U6621 (N_6621,N_6488,N_6490);
and U6622 (N_6622,N_6403,N_6494);
or U6623 (N_6623,N_6554,N_6594);
and U6624 (N_6624,N_6436,N_6437);
or U6625 (N_6625,N_6500,N_6573);
and U6626 (N_6626,N_6472,N_6478);
nand U6627 (N_6627,N_6451,N_6505);
and U6628 (N_6628,N_6516,N_6533);
and U6629 (N_6629,N_6429,N_6598);
or U6630 (N_6630,N_6515,N_6487);
or U6631 (N_6631,N_6424,N_6562);
and U6632 (N_6632,N_6462,N_6473);
nand U6633 (N_6633,N_6558,N_6471);
and U6634 (N_6634,N_6502,N_6574);
nor U6635 (N_6635,N_6519,N_6448);
nand U6636 (N_6636,N_6537,N_6479);
or U6637 (N_6637,N_6435,N_6442);
or U6638 (N_6638,N_6470,N_6482);
and U6639 (N_6639,N_6418,N_6534);
nand U6640 (N_6640,N_6597,N_6586);
or U6641 (N_6641,N_6405,N_6521);
or U6642 (N_6642,N_6546,N_6459);
nand U6643 (N_6643,N_6404,N_6570);
nand U6644 (N_6644,N_6421,N_6560);
nand U6645 (N_6645,N_6526,N_6552);
and U6646 (N_6646,N_6440,N_6422);
xnor U6647 (N_6647,N_6561,N_6406);
xor U6648 (N_6648,N_6464,N_6592);
nand U6649 (N_6649,N_6420,N_6582);
or U6650 (N_6650,N_6528,N_6531);
and U6651 (N_6651,N_6484,N_6467);
xor U6652 (N_6652,N_6507,N_6588);
xnor U6653 (N_6653,N_6544,N_6508);
nand U6654 (N_6654,N_6402,N_6477);
nand U6655 (N_6655,N_6503,N_6599);
nand U6656 (N_6656,N_6455,N_6453);
and U6657 (N_6657,N_6536,N_6543);
nand U6658 (N_6658,N_6587,N_6463);
or U6659 (N_6659,N_6581,N_6553);
nor U6660 (N_6660,N_6504,N_6564);
and U6661 (N_6661,N_6468,N_6497);
xnor U6662 (N_6662,N_6413,N_6427);
nand U6663 (N_6663,N_6571,N_6419);
or U6664 (N_6664,N_6530,N_6443);
and U6665 (N_6665,N_6452,N_6458);
nand U6666 (N_6666,N_6596,N_6409);
nand U6667 (N_6667,N_6486,N_6425);
nand U6668 (N_6668,N_6407,N_6514);
nand U6669 (N_6669,N_6550,N_6417);
nor U6670 (N_6670,N_6551,N_6495);
nor U6671 (N_6671,N_6591,N_6589);
nor U6672 (N_6672,N_6509,N_6517);
nand U6673 (N_6673,N_6556,N_6432);
nand U6674 (N_6674,N_6414,N_6539);
nor U6675 (N_6675,N_6518,N_6527);
and U6676 (N_6676,N_6522,N_6450);
nand U6677 (N_6677,N_6431,N_6506);
nand U6678 (N_6678,N_6520,N_6535);
or U6679 (N_6679,N_6565,N_6513);
and U6680 (N_6680,N_6447,N_6569);
and U6681 (N_6681,N_6559,N_6525);
or U6682 (N_6682,N_6496,N_6532);
or U6683 (N_6683,N_6492,N_6563);
or U6684 (N_6684,N_6430,N_6523);
and U6685 (N_6685,N_6568,N_6449);
nor U6686 (N_6686,N_6475,N_6426);
nand U6687 (N_6687,N_6434,N_6411);
or U6688 (N_6688,N_6466,N_6461);
or U6689 (N_6689,N_6439,N_6578);
nor U6690 (N_6690,N_6412,N_6480);
or U6691 (N_6691,N_6549,N_6415);
nand U6692 (N_6692,N_6433,N_6501);
nand U6693 (N_6693,N_6454,N_6493);
and U6694 (N_6694,N_6401,N_6566);
nor U6695 (N_6695,N_6446,N_6510);
or U6696 (N_6696,N_6469,N_6489);
nand U6697 (N_6697,N_6512,N_6567);
and U6698 (N_6698,N_6474,N_6572);
and U6699 (N_6699,N_6476,N_6579);
or U6700 (N_6700,N_6474,N_6526);
xor U6701 (N_6701,N_6459,N_6475);
or U6702 (N_6702,N_6502,N_6404);
or U6703 (N_6703,N_6538,N_6470);
and U6704 (N_6704,N_6415,N_6428);
and U6705 (N_6705,N_6499,N_6408);
nand U6706 (N_6706,N_6474,N_6549);
and U6707 (N_6707,N_6407,N_6474);
nor U6708 (N_6708,N_6497,N_6550);
nand U6709 (N_6709,N_6563,N_6538);
and U6710 (N_6710,N_6566,N_6419);
and U6711 (N_6711,N_6593,N_6579);
nand U6712 (N_6712,N_6465,N_6525);
nor U6713 (N_6713,N_6424,N_6587);
and U6714 (N_6714,N_6583,N_6467);
nor U6715 (N_6715,N_6556,N_6535);
and U6716 (N_6716,N_6583,N_6553);
nand U6717 (N_6717,N_6525,N_6557);
nor U6718 (N_6718,N_6490,N_6587);
nor U6719 (N_6719,N_6431,N_6429);
xnor U6720 (N_6720,N_6438,N_6570);
xor U6721 (N_6721,N_6436,N_6450);
or U6722 (N_6722,N_6551,N_6482);
or U6723 (N_6723,N_6418,N_6444);
xnor U6724 (N_6724,N_6564,N_6432);
nor U6725 (N_6725,N_6438,N_6496);
or U6726 (N_6726,N_6434,N_6499);
xor U6727 (N_6727,N_6431,N_6490);
or U6728 (N_6728,N_6538,N_6477);
nand U6729 (N_6729,N_6419,N_6586);
and U6730 (N_6730,N_6465,N_6517);
nand U6731 (N_6731,N_6567,N_6403);
xnor U6732 (N_6732,N_6535,N_6551);
xnor U6733 (N_6733,N_6587,N_6539);
and U6734 (N_6734,N_6501,N_6406);
xnor U6735 (N_6735,N_6480,N_6411);
nor U6736 (N_6736,N_6579,N_6483);
or U6737 (N_6737,N_6431,N_6475);
xnor U6738 (N_6738,N_6492,N_6521);
nand U6739 (N_6739,N_6517,N_6539);
and U6740 (N_6740,N_6573,N_6529);
xnor U6741 (N_6741,N_6430,N_6469);
nand U6742 (N_6742,N_6450,N_6503);
nor U6743 (N_6743,N_6421,N_6576);
and U6744 (N_6744,N_6460,N_6599);
nor U6745 (N_6745,N_6451,N_6500);
and U6746 (N_6746,N_6597,N_6522);
and U6747 (N_6747,N_6508,N_6568);
nand U6748 (N_6748,N_6540,N_6528);
and U6749 (N_6749,N_6409,N_6473);
and U6750 (N_6750,N_6409,N_6515);
and U6751 (N_6751,N_6517,N_6596);
and U6752 (N_6752,N_6498,N_6519);
nand U6753 (N_6753,N_6537,N_6431);
nand U6754 (N_6754,N_6492,N_6517);
nor U6755 (N_6755,N_6554,N_6501);
and U6756 (N_6756,N_6437,N_6466);
or U6757 (N_6757,N_6565,N_6551);
and U6758 (N_6758,N_6598,N_6446);
nand U6759 (N_6759,N_6527,N_6564);
xnor U6760 (N_6760,N_6422,N_6516);
or U6761 (N_6761,N_6555,N_6542);
or U6762 (N_6762,N_6540,N_6583);
nand U6763 (N_6763,N_6581,N_6416);
or U6764 (N_6764,N_6525,N_6480);
nor U6765 (N_6765,N_6488,N_6475);
nor U6766 (N_6766,N_6501,N_6472);
xor U6767 (N_6767,N_6506,N_6430);
and U6768 (N_6768,N_6432,N_6415);
nor U6769 (N_6769,N_6526,N_6576);
nor U6770 (N_6770,N_6568,N_6435);
nor U6771 (N_6771,N_6512,N_6586);
and U6772 (N_6772,N_6469,N_6456);
nor U6773 (N_6773,N_6518,N_6536);
or U6774 (N_6774,N_6445,N_6558);
or U6775 (N_6775,N_6513,N_6546);
or U6776 (N_6776,N_6408,N_6438);
xnor U6777 (N_6777,N_6402,N_6425);
xnor U6778 (N_6778,N_6597,N_6537);
and U6779 (N_6779,N_6502,N_6531);
or U6780 (N_6780,N_6586,N_6488);
xnor U6781 (N_6781,N_6531,N_6540);
and U6782 (N_6782,N_6504,N_6461);
nand U6783 (N_6783,N_6545,N_6562);
nand U6784 (N_6784,N_6559,N_6456);
nor U6785 (N_6785,N_6455,N_6414);
nand U6786 (N_6786,N_6424,N_6473);
or U6787 (N_6787,N_6513,N_6461);
xnor U6788 (N_6788,N_6530,N_6579);
xnor U6789 (N_6789,N_6551,N_6568);
xnor U6790 (N_6790,N_6412,N_6407);
or U6791 (N_6791,N_6593,N_6423);
and U6792 (N_6792,N_6478,N_6566);
or U6793 (N_6793,N_6521,N_6512);
or U6794 (N_6794,N_6511,N_6476);
and U6795 (N_6795,N_6537,N_6493);
or U6796 (N_6796,N_6412,N_6550);
or U6797 (N_6797,N_6590,N_6551);
nor U6798 (N_6798,N_6564,N_6553);
nand U6799 (N_6799,N_6484,N_6479);
xor U6800 (N_6800,N_6691,N_6778);
and U6801 (N_6801,N_6641,N_6638);
or U6802 (N_6802,N_6602,N_6694);
or U6803 (N_6803,N_6623,N_6788);
nor U6804 (N_6804,N_6758,N_6724);
xnor U6805 (N_6805,N_6634,N_6682);
nor U6806 (N_6806,N_6662,N_6692);
and U6807 (N_6807,N_6684,N_6637);
or U6808 (N_6808,N_6755,N_6765);
and U6809 (N_6809,N_6636,N_6734);
or U6810 (N_6810,N_6631,N_6657);
and U6811 (N_6811,N_6675,N_6674);
or U6812 (N_6812,N_6799,N_6663);
or U6813 (N_6813,N_6644,N_6654);
nand U6814 (N_6814,N_6647,N_6613);
xor U6815 (N_6815,N_6779,N_6665);
or U6816 (N_6816,N_6748,N_6706);
nor U6817 (N_6817,N_6655,N_6639);
or U6818 (N_6818,N_6702,N_6699);
nand U6819 (N_6819,N_6646,N_6786);
xor U6820 (N_6820,N_6696,N_6718);
xnor U6821 (N_6821,N_6793,N_6652);
nand U6822 (N_6822,N_6608,N_6769);
xnor U6823 (N_6823,N_6751,N_6754);
nor U6824 (N_6824,N_6749,N_6732);
nand U6825 (N_6825,N_6610,N_6743);
nand U6826 (N_6826,N_6740,N_6686);
and U6827 (N_6827,N_6775,N_6745);
nor U6828 (N_6828,N_6773,N_6629);
xor U6829 (N_6829,N_6677,N_6739);
nor U6830 (N_6830,N_6719,N_6771);
xor U6831 (N_6831,N_6622,N_6603);
xnor U6832 (N_6832,N_6703,N_6667);
or U6833 (N_6833,N_6716,N_6700);
nor U6834 (N_6834,N_6625,N_6762);
nor U6835 (N_6835,N_6624,N_6656);
xnor U6836 (N_6836,N_6756,N_6760);
and U6837 (N_6837,N_6709,N_6768);
xnor U6838 (N_6838,N_6673,N_6661);
and U6839 (N_6839,N_6707,N_6681);
nor U6840 (N_6840,N_6725,N_6776);
nor U6841 (N_6841,N_6791,N_6780);
or U6842 (N_6842,N_6723,N_6733);
or U6843 (N_6843,N_6697,N_6600);
nand U6844 (N_6844,N_6666,N_6632);
and U6845 (N_6845,N_6615,N_6676);
nor U6846 (N_6846,N_6651,N_6738);
xor U6847 (N_6847,N_6757,N_6790);
or U6848 (N_6848,N_6648,N_6658);
and U6849 (N_6849,N_6616,N_6742);
xor U6850 (N_6850,N_6714,N_6766);
xor U6851 (N_6851,N_6736,N_6649);
nand U6852 (N_6852,N_6704,N_6785);
or U6853 (N_6853,N_6764,N_6630);
xnor U6854 (N_6854,N_6690,N_6787);
nor U6855 (N_6855,N_6669,N_6687);
and U6856 (N_6856,N_6782,N_6671);
nor U6857 (N_6857,N_6761,N_6672);
nand U6858 (N_6858,N_6789,N_6731);
xnor U6859 (N_6859,N_6712,N_6640);
nand U6860 (N_6860,N_6607,N_6685);
nand U6861 (N_6861,N_6767,N_6772);
nand U6862 (N_6862,N_6601,N_6794);
and U6863 (N_6863,N_6750,N_6659);
or U6864 (N_6864,N_6653,N_6660);
nand U6865 (N_6865,N_6701,N_6688);
nand U6866 (N_6866,N_6606,N_6617);
or U6867 (N_6867,N_6722,N_6620);
and U6868 (N_6868,N_6693,N_6727);
xor U6869 (N_6869,N_6643,N_6628);
and U6870 (N_6870,N_6650,N_6753);
or U6871 (N_6871,N_6633,N_6670);
or U6872 (N_6872,N_6747,N_6777);
xnor U6873 (N_6873,N_6664,N_6679);
and U6874 (N_6874,N_6797,N_6604);
or U6875 (N_6875,N_6726,N_6710);
and U6876 (N_6876,N_6774,N_6626);
and U6877 (N_6877,N_6619,N_6781);
nand U6878 (N_6878,N_6605,N_6770);
xnor U6879 (N_6879,N_6695,N_6735);
and U6880 (N_6880,N_6642,N_6698);
and U6881 (N_6881,N_6721,N_6784);
nand U6882 (N_6882,N_6711,N_6713);
and U6883 (N_6883,N_6728,N_6614);
xnor U6884 (N_6884,N_6729,N_6618);
and U6885 (N_6885,N_6609,N_6645);
xor U6886 (N_6886,N_6708,N_6720);
nand U6887 (N_6887,N_6741,N_6752);
nand U6888 (N_6888,N_6759,N_6611);
nand U6889 (N_6889,N_6798,N_6612);
or U6890 (N_6890,N_6689,N_6717);
xor U6891 (N_6891,N_6678,N_6621);
xor U6892 (N_6892,N_6792,N_6737);
and U6893 (N_6893,N_6746,N_6705);
xor U6894 (N_6894,N_6627,N_6668);
or U6895 (N_6895,N_6796,N_6635);
nand U6896 (N_6896,N_6783,N_6763);
xor U6897 (N_6897,N_6683,N_6795);
and U6898 (N_6898,N_6680,N_6715);
nand U6899 (N_6899,N_6730,N_6744);
nand U6900 (N_6900,N_6748,N_6798);
nor U6901 (N_6901,N_6777,N_6665);
nand U6902 (N_6902,N_6731,N_6771);
and U6903 (N_6903,N_6651,N_6741);
or U6904 (N_6904,N_6633,N_6730);
xor U6905 (N_6905,N_6756,N_6649);
xnor U6906 (N_6906,N_6663,N_6775);
nor U6907 (N_6907,N_6669,N_6617);
or U6908 (N_6908,N_6704,N_6713);
xnor U6909 (N_6909,N_6768,N_6760);
nor U6910 (N_6910,N_6763,N_6764);
and U6911 (N_6911,N_6697,N_6772);
xor U6912 (N_6912,N_6765,N_6672);
and U6913 (N_6913,N_6679,N_6769);
nand U6914 (N_6914,N_6652,N_6687);
or U6915 (N_6915,N_6649,N_6769);
nor U6916 (N_6916,N_6761,N_6734);
and U6917 (N_6917,N_6699,N_6656);
and U6918 (N_6918,N_6719,N_6650);
nand U6919 (N_6919,N_6686,N_6673);
and U6920 (N_6920,N_6662,N_6619);
nand U6921 (N_6921,N_6677,N_6795);
nor U6922 (N_6922,N_6723,N_6646);
nor U6923 (N_6923,N_6775,N_6628);
and U6924 (N_6924,N_6796,N_6609);
nand U6925 (N_6925,N_6755,N_6651);
xnor U6926 (N_6926,N_6676,N_6662);
nor U6927 (N_6927,N_6676,N_6604);
and U6928 (N_6928,N_6699,N_6685);
xor U6929 (N_6929,N_6627,N_6678);
and U6930 (N_6930,N_6683,N_6623);
nand U6931 (N_6931,N_6792,N_6666);
and U6932 (N_6932,N_6667,N_6702);
nand U6933 (N_6933,N_6658,N_6679);
xor U6934 (N_6934,N_6688,N_6649);
and U6935 (N_6935,N_6633,N_6767);
or U6936 (N_6936,N_6648,N_6674);
xnor U6937 (N_6937,N_6644,N_6689);
and U6938 (N_6938,N_6645,N_6661);
nand U6939 (N_6939,N_6643,N_6755);
xnor U6940 (N_6940,N_6692,N_6799);
and U6941 (N_6941,N_6799,N_6693);
nor U6942 (N_6942,N_6784,N_6698);
nor U6943 (N_6943,N_6635,N_6770);
nand U6944 (N_6944,N_6761,N_6753);
nand U6945 (N_6945,N_6702,N_6719);
nand U6946 (N_6946,N_6614,N_6763);
nor U6947 (N_6947,N_6669,N_6644);
or U6948 (N_6948,N_6791,N_6680);
nor U6949 (N_6949,N_6723,N_6644);
or U6950 (N_6950,N_6776,N_6792);
and U6951 (N_6951,N_6707,N_6600);
nand U6952 (N_6952,N_6771,N_6642);
xor U6953 (N_6953,N_6775,N_6692);
xor U6954 (N_6954,N_6665,N_6751);
and U6955 (N_6955,N_6779,N_6655);
nand U6956 (N_6956,N_6764,N_6790);
and U6957 (N_6957,N_6623,N_6799);
or U6958 (N_6958,N_6776,N_6730);
nor U6959 (N_6959,N_6765,N_6684);
nand U6960 (N_6960,N_6688,N_6640);
and U6961 (N_6961,N_6641,N_6619);
and U6962 (N_6962,N_6781,N_6724);
nor U6963 (N_6963,N_6639,N_6631);
nor U6964 (N_6964,N_6737,N_6632);
xor U6965 (N_6965,N_6665,N_6615);
nor U6966 (N_6966,N_6791,N_6636);
and U6967 (N_6967,N_6761,N_6759);
nand U6968 (N_6968,N_6724,N_6763);
nand U6969 (N_6969,N_6669,N_6721);
xor U6970 (N_6970,N_6678,N_6699);
nor U6971 (N_6971,N_6682,N_6670);
xnor U6972 (N_6972,N_6747,N_6630);
nor U6973 (N_6973,N_6746,N_6716);
or U6974 (N_6974,N_6638,N_6602);
and U6975 (N_6975,N_6690,N_6623);
and U6976 (N_6976,N_6695,N_6603);
or U6977 (N_6977,N_6604,N_6694);
nor U6978 (N_6978,N_6799,N_6779);
nor U6979 (N_6979,N_6674,N_6733);
xor U6980 (N_6980,N_6700,N_6682);
xor U6981 (N_6981,N_6672,N_6715);
or U6982 (N_6982,N_6630,N_6738);
and U6983 (N_6983,N_6775,N_6726);
or U6984 (N_6984,N_6795,N_6679);
nand U6985 (N_6985,N_6705,N_6785);
nand U6986 (N_6986,N_6612,N_6744);
or U6987 (N_6987,N_6791,N_6655);
nor U6988 (N_6988,N_6604,N_6644);
nand U6989 (N_6989,N_6653,N_6710);
nand U6990 (N_6990,N_6769,N_6718);
and U6991 (N_6991,N_6653,N_6782);
and U6992 (N_6992,N_6668,N_6726);
or U6993 (N_6993,N_6644,N_6625);
or U6994 (N_6994,N_6638,N_6696);
or U6995 (N_6995,N_6661,N_6707);
and U6996 (N_6996,N_6738,N_6717);
nand U6997 (N_6997,N_6637,N_6731);
and U6998 (N_6998,N_6680,N_6616);
nand U6999 (N_6999,N_6789,N_6643);
and U7000 (N_7000,N_6941,N_6996);
or U7001 (N_7001,N_6891,N_6961);
nor U7002 (N_7002,N_6859,N_6863);
nand U7003 (N_7003,N_6936,N_6944);
nor U7004 (N_7004,N_6997,N_6933);
nor U7005 (N_7005,N_6845,N_6907);
nand U7006 (N_7006,N_6934,N_6802);
nor U7007 (N_7007,N_6877,N_6966);
or U7008 (N_7008,N_6890,N_6828);
xnor U7009 (N_7009,N_6968,N_6826);
or U7010 (N_7010,N_6956,N_6894);
and U7011 (N_7011,N_6927,N_6811);
xnor U7012 (N_7012,N_6977,N_6861);
or U7013 (N_7013,N_6914,N_6888);
and U7014 (N_7014,N_6827,N_6825);
and U7015 (N_7015,N_6878,N_6946);
nand U7016 (N_7016,N_6900,N_6882);
nand U7017 (N_7017,N_6880,N_6959);
or U7018 (N_7018,N_6831,N_6816);
xnor U7019 (N_7019,N_6841,N_6805);
nand U7020 (N_7020,N_6897,N_6987);
nor U7021 (N_7021,N_6820,N_6875);
nor U7022 (N_7022,N_6969,N_6860);
and U7023 (N_7023,N_6804,N_6868);
nor U7024 (N_7024,N_6840,N_6857);
nand U7025 (N_7025,N_6916,N_6912);
or U7026 (N_7026,N_6832,N_6869);
and U7027 (N_7027,N_6919,N_6847);
nor U7028 (N_7028,N_6846,N_6906);
nor U7029 (N_7029,N_6932,N_6807);
xor U7030 (N_7030,N_6808,N_6978);
or U7031 (N_7031,N_6853,N_6979);
xnor U7032 (N_7032,N_6823,N_6953);
xor U7033 (N_7033,N_6922,N_6871);
xor U7034 (N_7034,N_6948,N_6901);
and U7035 (N_7035,N_6949,N_6943);
and U7036 (N_7036,N_6848,N_6814);
nand U7037 (N_7037,N_6862,N_6817);
or U7038 (N_7038,N_6809,N_6965);
nand U7039 (N_7039,N_6874,N_6958);
nand U7040 (N_7040,N_6990,N_6818);
and U7041 (N_7041,N_6992,N_6926);
nor U7042 (N_7042,N_6833,N_6837);
xnor U7043 (N_7043,N_6954,N_6852);
xor U7044 (N_7044,N_6854,N_6812);
or U7045 (N_7045,N_6980,N_6838);
nor U7046 (N_7046,N_6885,N_6994);
and U7047 (N_7047,N_6908,N_6952);
xnor U7048 (N_7048,N_6824,N_6917);
or U7049 (N_7049,N_6849,N_6950);
xnor U7050 (N_7050,N_6879,N_6829);
or U7051 (N_7051,N_6989,N_6887);
and U7052 (N_7052,N_6867,N_6813);
or U7053 (N_7053,N_6999,N_6905);
or U7054 (N_7054,N_6881,N_6865);
or U7055 (N_7055,N_6986,N_6975);
nor U7056 (N_7056,N_6973,N_6971);
nand U7057 (N_7057,N_6844,N_6850);
or U7058 (N_7058,N_6985,N_6902);
and U7059 (N_7059,N_6864,N_6876);
nand U7060 (N_7060,N_6929,N_6892);
nor U7061 (N_7061,N_6895,N_6858);
and U7062 (N_7062,N_6972,N_6851);
or U7063 (N_7063,N_6872,N_6931);
nand U7064 (N_7064,N_6898,N_6920);
nand U7065 (N_7065,N_6967,N_6945);
or U7066 (N_7066,N_6884,N_6842);
nor U7067 (N_7067,N_6839,N_6909);
nor U7068 (N_7068,N_6955,N_6939);
or U7069 (N_7069,N_6899,N_6964);
nand U7070 (N_7070,N_6800,N_6836);
nor U7071 (N_7071,N_6930,N_6821);
or U7072 (N_7072,N_6960,N_6886);
xnor U7073 (N_7073,N_6998,N_6951);
nand U7074 (N_7074,N_6963,N_6935);
xor U7075 (N_7075,N_6957,N_6947);
or U7076 (N_7076,N_6915,N_6988);
xor U7077 (N_7077,N_6910,N_6806);
nor U7078 (N_7078,N_6984,N_6983);
xnor U7079 (N_7079,N_6938,N_6893);
and U7080 (N_7080,N_6982,N_6819);
or U7081 (N_7081,N_6896,N_6942);
nor U7082 (N_7082,N_6801,N_6913);
xnor U7083 (N_7083,N_6928,N_6830);
nand U7084 (N_7084,N_6883,N_6835);
nand U7085 (N_7085,N_6903,N_6918);
and U7086 (N_7086,N_6843,N_6923);
or U7087 (N_7087,N_6870,N_6873);
and U7088 (N_7088,N_6995,N_6991);
nand U7089 (N_7089,N_6810,N_6911);
or U7090 (N_7090,N_6921,N_6856);
nand U7091 (N_7091,N_6962,N_6974);
xor U7092 (N_7092,N_6904,N_6803);
and U7093 (N_7093,N_6866,N_6822);
xor U7094 (N_7094,N_6976,N_6889);
xor U7095 (N_7095,N_6855,N_6925);
or U7096 (N_7096,N_6981,N_6970);
or U7097 (N_7097,N_6834,N_6937);
and U7098 (N_7098,N_6815,N_6940);
nor U7099 (N_7099,N_6993,N_6924);
nor U7100 (N_7100,N_6878,N_6975);
nand U7101 (N_7101,N_6990,N_6888);
and U7102 (N_7102,N_6982,N_6930);
nand U7103 (N_7103,N_6861,N_6974);
nand U7104 (N_7104,N_6817,N_6901);
nand U7105 (N_7105,N_6823,N_6931);
nor U7106 (N_7106,N_6900,N_6887);
and U7107 (N_7107,N_6822,N_6932);
and U7108 (N_7108,N_6987,N_6864);
or U7109 (N_7109,N_6998,N_6827);
or U7110 (N_7110,N_6946,N_6834);
xnor U7111 (N_7111,N_6954,N_6819);
nor U7112 (N_7112,N_6953,N_6910);
nor U7113 (N_7113,N_6927,N_6935);
and U7114 (N_7114,N_6952,N_6897);
or U7115 (N_7115,N_6856,N_6946);
or U7116 (N_7116,N_6910,N_6918);
xnor U7117 (N_7117,N_6863,N_6994);
and U7118 (N_7118,N_6815,N_6859);
nand U7119 (N_7119,N_6843,N_6968);
or U7120 (N_7120,N_6913,N_6955);
nand U7121 (N_7121,N_6925,N_6983);
xor U7122 (N_7122,N_6915,N_6849);
nor U7123 (N_7123,N_6856,N_6908);
and U7124 (N_7124,N_6850,N_6978);
xnor U7125 (N_7125,N_6929,N_6802);
nor U7126 (N_7126,N_6842,N_6875);
nand U7127 (N_7127,N_6936,N_6938);
or U7128 (N_7128,N_6971,N_6949);
xor U7129 (N_7129,N_6891,N_6962);
nor U7130 (N_7130,N_6857,N_6807);
nand U7131 (N_7131,N_6945,N_6975);
xnor U7132 (N_7132,N_6874,N_6879);
nor U7133 (N_7133,N_6900,N_6868);
nor U7134 (N_7134,N_6880,N_6958);
xor U7135 (N_7135,N_6862,N_6880);
nor U7136 (N_7136,N_6840,N_6800);
and U7137 (N_7137,N_6829,N_6921);
nor U7138 (N_7138,N_6955,N_6857);
or U7139 (N_7139,N_6896,N_6818);
nand U7140 (N_7140,N_6802,N_6951);
nor U7141 (N_7141,N_6998,N_6956);
and U7142 (N_7142,N_6990,N_6814);
and U7143 (N_7143,N_6803,N_6914);
xor U7144 (N_7144,N_6908,N_6948);
nand U7145 (N_7145,N_6918,N_6924);
and U7146 (N_7146,N_6830,N_6851);
or U7147 (N_7147,N_6931,N_6815);
nand U7148 (N_7148,N_6864,N_6840);
or U7149 (N_7149,N_6960,N_6949);
and U7150 (N_7150,N_6840,N_6809);
nor U7151 (N_7151,N_6833,N_6991);
xnor U7152 (N_7152,N_6815,N_6973);
or U7153 (N_7153,N_6923,N_6831);
xnor U7154 (N_7154,N_6948,N_6925);
or U7155 (N_7155,N_6873,N_6813);
or U7156 (N_7156,N_6987,N_6872);
nand U7157 (N_7157,N_6834,N_6825);
nor U7158 (N_7158,N_6831,N_6842);
or U7159 (N_7159,N_6903,N_6821);
or U7160 (N_7160,N_6880,N_6889);
and U7161 (N_7161,N_6860,N_6858);
xnor U7162 (N_7162,N_6933,N_6864);
nor U7163 (N_7163,N_6855,N_6847);
and U7164 (N_7164,N_6943,N_6845);
nand U7165 (N_7165,N_6862,N_6884);
and U7166 (N_7166,N_6916,N_6904);
xor U7167 (N_7167,N_6824,N_6964);
or U7168 (N_7168,N_6830,N_6915);
or U7169 (N_7169,N_6993,N_6831);
or U7170 (N_7170,N_6819,N_6834);
nor U7171 (N_7171,N_6840,N_6962);
and U7172 (N_7172,N_6975,N_6845);
and U7173 (N_7173,N_6962,N_6802);
or U7174 (N_7174,N_6832,N_6937);
nand U7175 (N_7175,N_6956,N_6940);
and U7176 (N_7176,N_6803,N_6945);
xnor U7177 (N_7177,N_6859,N_6906);
nor U7178 (N_7178,N_6950,N_6973);
and U7179 (N_7179,N_6946,N_6990);
nor U7180 (N_7180,N_6959,N_6974);
xnor U7181 (N_7181,N_6841,N_6803);
and U7182 (N_7182,N_6865,N_6982);
nand U7183 (N_7183,N_6908,N_6863);
xor U7184 (N_7184,N_6991,N_6960);
nor U7185 (N_7185,N_6997,N_6974);
or U7186 (N_7186,N_6941,N_6809);
or U7187 (N_7187,N_6980,N_6993);
nor U7188 (N_7188,N_6869,N_6973);
xnor U7189 (N_7189,N_6812,N_6863);
or U7190 (N_7190,N_6854,N_6976);
and U7191 (N_7191,N_6854,N_6848);
xnor U7192 (N_7192,N_6990,N_6868);
and U7193 (N_7193,N_6808,N_6960);
and U7194 (N_7194,N_6833,N_6891);
nand U7195 (N_7195,N_6999,N_6930);
nand U7196 (N_7196,N_6988,N_6960);
or U7197 (N_7197,N_6862,N_6980);
and U7198 (N_7198,N_6860,N_6981);
nor U7199 (N_7199,N_6945,N_6853);
and U7200 (N_7200,N_7039,N_7059);
nor U7201 (N_7201,N_7085,N_7162);
and U7202 (N_7202,N_7092,N_7163);
and U7203 (N_7203,N_7000,N_7107);
or U7204 (N_7204,N_7108,N_7012);
nor U7205 (N_7205,N_7063,N_7167);
and U7206 (N_7206,N_7029,N_7055);
and U7207 (N_7207,N_7173,N_7149);
nand U7208 (N_7208,N_7024,N_7174);
nand U7209 (N_7209,N_7037,N_7090);
nand U7210 (N_7210,N_7035,N_7195);
or U7211 (N_7211,N_7193,N_7150);
or U7212 (N_7212,N_7114,N_7156);
or U7213 (N_7213,N_7031,N_7030);
nand U7214 (N_7214,N_7138,N_7026);
and U7215 (N_7215,N_7040,N_7001);
and U7216 (N_7216,N_7151,N_7176);
nor U7217 (N_7217,N_7079,N_7099);
nor U7218 (N_7218,N_7147,N_7111);
and U7219 (N_7219,N_7160,N_7142);
xor U7220 (N_7220,N_7082,N_7008);
nor U7221 (N_7221,N_7127,N_7089);
nor U7222 (N_7222,N_7102,N_7074);
nand U7223 (N_7223,N_7178,N_7096);
xor U7224 (N_7224,N_7006,N_7105);
xnor U7225 (N_7225,N_7103,N_7093);
or U7226 (N_7226,N_7018,N_7194);
nor U7227 (N_7227,N_7170,N_7014);
and U7228 (N_7228,N_7051,N_7075);
nand U7229 (N_7229,N_7036,N_7116);
nor U7230 (N_7230,N_7118,N_7058);
nor U7231 (N_7231,N_7146,N_7081);
or U7232 (N_7232,N_7027,N_7153);
xnor U7233 (N_7233,N_7190,N_7130);
xnor U7234 (N_7234,N_7175,N_7067);
and U7235 (N_7235,N_7033,N_7154);
and U7236 (N_7236,N_7155,N_7041);
nand U7237 (N_7237,N_7091,N_7186);
nor U7238 (N_7238,N_7177,N_7080);
nand U7239 (N_7239,N_7045,N_7183);
or U7240 (N_7240,N_7199,N_7043);
or U7241 (N_7241,N_7181,N_7070);
or U7242 (N_7242,N_7021,N_7143);
and U7243 (N_7243,N_7047,N_7123);
nor U7244 (N_7244,N_7159,N_7066);
nand U7245 (N_7245,N_7022,N_7073);
and U7246 (N_7246,N_7017,N_7166);
and U7247 (N_7247,N_7015,N_7097);
xnor U7248 (N_7248,N_7078,N_7019);
or U7249 (N_7249,N_7110,N_7124);
nor U7250 (N_7250,N_7044,N_7122);
xnor U7251 (N_7251,N_7060,N_7023);
nand U7252 (N_7252,N_7144,N_7064);
nor U7253 (N_7253,N_7084,N_7148);
nand U7254 (N_7254,N_7061,N_7007);
and U7255 (N_7255,N_7071,N_7121);
nand U7256 (N_7256,N_7129,N_7168);
or U7257 (N_7257,N_7113,N_7010);
xor U7258 (N_7258,N_7098,N_7069);
nor U7259 (N_7259,N_7157,N_7101);
or U7260 (N_7260,N_7077,N_7002);
and U7261 (N_7261,N_7196,N_7003);
or U7262 (N_7262,N_7137,N_7020);
nor U7263 (N_7263,N_7005,N_7100);
or U7264 (N_7264,N_7197,N_7125);
nor U7265 (N_7265,N_7048,N_7042);
nor U7266 (N_7266,N_7187,N_7013);
and U7267 (N_7267,N_7141,N_7094);
or U7268 (N_7268,N_7095,N_7140);
and U7269 (N_7269,N_7068,N_7028);
and U7270 (N_7270,N_7057,N_7112);
and U7271 (N_7271,N_7120,N_7182);
or U7272 (N_7272,N_7052,N_7164);
xor U7273 (N_7273,N_7161,N_7172);
and U7274 (N_7274,N_7139,N_7128);
nand U7275 (N_7275,N_7188,N_7185);
or U7276 (N_7276,N_7032,N_7198);
nand U7277 (N_7277,N_7191,N_7050);
xor U7278 (N_7278,N_7009,N_7109);
nand U7279 (N_7279,N_7158,N_7034);
and U7280 (N_7280,N_7106,N_7038);
or U7281 (N_7281,N_7076,N_7152);
or U7282 (N_7282,N_7165,N_7119);
nand U7283 (N_7283,N_7016,N_7132);
and U7284 (N_7284,N_7025,N_7088);
nand U7285 (N_7285,N_7145,N_7115);
or U7286 (N_7286,N_7126,N_7046);
nor U7287 (N_7287,N_7086,N_7136);
and U7288 (N_7288,N_7133,N_7072);
and U7289 (N_7289,N_7062,N_7169);
or U7290 (N_7290,N_7171,N_7049);
and U7291 (N_7291,N_7054,N_7189);
and U7292 (N_7292,N_7134,N_7131);
or U7293 (N_7293,N_7180,N_7104);
or U7294 (N_7294,N_7083,N_7184);
xor U7295 (N_7295,N_7192,N_7011);
or U7296 (N_7296,N_7087,N_7179);
and U7297 (N_7297,N_7065,N_7117);
and U7298 (N_7298,N_7004,N_7053);
or U7299 (N_7299,N_7056,N_7135);
or U7300 (N_7300,N_7077,N_7110);
or U7301 (N_7301,N_7094,N_7068);
nand U7302 (N_7302,N_7010,N_7051);
nand U7303 (N_7303,N_7088,N_7149);
nor U7304 (N_7304,N_7082,N_7182);
and U7305 (N_7305,N_7007,N_7172);
or U7306 (N_7306,N_7036,N_7012);
xnor U7307 (N_7307,N_7062,N_7043);
and U7308 (N_7308,N_7188,N_7014);
xnor U7309 (N_7309,N_7046,N_7181);
xor U7310 (N_7310,N_7011,N_7047);
or U7311 (N_7311,N_7130,N_7042);
xnor U7312 (N_7312,N_7004,N_7107);
nand U7313 (N_7313,N_7097,N_7069);
xnor U7314 (N_7314,N_7182,N_7193);
nand U7315 (N_7315,N_7161,N_7030);
nand U7316 (N_7316,N_7125,N_7112);
and U7317 (N_7317,N_7066,N_7168);
and U7318 (N_7318,N_7167,N_7133);
nand U7319 (N_7319,N_7030,N_7084);
or U7320 (N_7320,N_7063,N_7027);
nand U7321 (N_7321,N_7160,N_7111);
xnor U7322 (N_7322,N_7173,N_7168);
or U7323 (N_7323,N_7101,N_7102);
nand U7324 (N_7324,N_7003,N_7135);
or U7325 (N_7325,N_7063,N_7135);
xor U7326 (N_7326,N_7199,N_7083);
nor U7327 (N_7327,N_7030,N_7013);
or U7328 (N_7328,N_7087,N_7170);
nor U7329 (N_7329,N_7134,N_7044);
nand U7330 (N_7330,N_7150,N_7066);
xnor U7331 (N_7331,N_7171,N_7086);
xor U7332 (N_7332,N_7087,N_7050);
nand U7333 (N_7333,N_7186,N_7126);
or U7334 (N_7334,N_7024,N_7067);
or U7335 (N_7335,N_7019,N_7199);
nor U7336 (N_7336,N_7152,N_7108);
and U7337 (N_7337,N_7185,N_7063);
xnor U7338 (N_7338,N_7079,N_7016);
nor U7339 (N_7339,N_7138,N_7120);
nor U7340 (N_7340,N_7181,N_7125);
nand U7341 (N_7341,N_7174,N_7132);
or U7342 (N_7342,N_7182,N_7048);
xor U7343 (N_7343,N_7128,N_7007);
nand U7344 (N_7344,N_7132,N_7071);
nor U7345 (N_7345,N_7118,N_7157);
and U7346 (N_7346,N_7127,N_7059);
xnor U7347 (N_7347,N_7116,N_7131);
or U7348 (N_7348,N_7027,N_7059);
or U7349 (N_7349,N_7108,N_7060);
and U7350 (N_7350,N_7005,N_7091);
xnor U7351 (N_7351,N_7014,N_7196);
nand U7352 (N_7352,N_7119,N_7015);
or U7353 (N_7353,N_7014,N_7044);
or U7354 (N_7354,N_7036,N_7007);
nor U7355 (N_7355,N_7003,N_7101);
or U7356 (N_7356,N_7073,N_7051);
and U7357 (N_7357,N_7055,N_7067);
or U7358 (N_7358,N_7003,N_7174);
and U7359 (N_7359,N_7137,N_7191);
or U7360 (N_7360,N_7117,N_7124);
and U7361 (N_7361,N_7094,N_7023);
xor U7362 (N_7362,N_7028,N_7073);
or U7363 (N_7363,N_7049,N_7048);
xnor U7364 (N_7364,N_7180,N_7101);
nor U7365 (N_7365,N_7099,N_7097);
or U7366 (N_7366,N_7038,N_7182);
and U7367 (N_7367,N_7010,N_7034);
nand U7368 (N_7368,N_7021,N_7181);
nor U7369 (N_7369,N_7065,N_7018);
nor U7370 (N_7370,N_7114,N_7000);
or U7371 (N_7371,N_7088,N_7114);
nor U7372 (N_7372,N_7142,N_7040);
nor U7373 (N_7373,N_7138,N_7021);
nor U7374 (N_7374,N_7187,N_7195);
nand U7375 (N_7375,N_7040,N_7108);
nor U7376 (N_7376,N_7149,N_7148);
nand U7377 (N_7377,N_7117,N_7111);
nand U7378 (N_7378,N_7111,N_7012);
and U7379 (N_7379,N_7052,N_7030);
nor U7380 (N_7380,N_7095,N_7158);
nand U7381 (N_7381,N_7140,N_7145);
xnor U7382 (N_7382,N_7192,N_7073);
xor U7383 (N_7383,N_7101,N_7067);
nor U7384 (N_7384,N_7058,N_7040);
nand U7385 (N_7385,N_7009,N_7148);
nor U7386 (N_7386,N_7050,N_7033);
xor U7387 (N_7387,N_7027,N_7060);
nand U7388 (N_7388,N_7089,N_7072);
nand U7389 (N_7389,N_7041,N_7070);
and U7390 (N_7390,N_7040,N_7081);
nand U7391 (N_7391,N_7087,N_7140);
or U7392 (N_7392,N_7056,N_7119);
xnor U7393 (N_7393,N_7105,N_7113);
xnor U7394 (N_7394,N_7106,N_7175);
nand U7395 (N_7395,N_7128,N_7166);
nor U7396 (N_7396,N_7085,N_7076);
or U7397 (N_7397,N_7139,N_7188);
or U7398 (N_7398,N_7063,N_7122);
or U7399 (N_7399,N_7180,N_7120);
and U7400 (N_7400,N_7205,N_7298);
xor U7401 (N_7401,N_7270,N_7347);
xor U7402 (N_7402,N_7326,N_7366);
nor U7403 (N_7403,N_7387,N_7377);
xnor U7404 (N_7404,N_7224,N_7314);
or U7405 (N_7405,N_7203,N_7350);
xnor U7406 (N_7406,N_7223,N_7333);
nand U7407 (N_7407,N_7250,N_7291);
nand U7408 (N_7408,N_7266,N_7212);
xnor U7409 (N_7409,N_7358,N_7289);
xnor U7410 (N_7410,N_7395,N_7344);
xor U7411 (N_7411,N_7254,N_7336);
or U7412 (N_7412,N_7339,N_7319);
nor U7413 (N_7413,N_7240,N_7308);
and U7414 (N_7414,N_7248,N_7269);
or U7415 (N_7415,N_7249,N_7315);
nor U7416 (N_7416,N_7374,N_7389);
or U7417 (N_7417,N_7274,N_7391);
nand U7418 (N_7418,N_7258,N_7290);
xnor U7419 (N_7419,N_7257,N_7352);
and U7420 (N_7420,N_7247,N_7268);
xnor U7421 (N_7421,N_7342,N_7292);
nor U7422 (N_7422,N_7293,N_7362);
nand U7423 (N_7423,N_7295,N_7375);
nand U7424 (N_7424,N_7369,N_7200);
or U7425 (N_7425,N_7312,N_7235);
and U7426 (N_7426,N_7243,N_7379);
and U7427 (N_7427,N_7394,N_7372);
nor U7428 (N_7428,N_7202,N_7299);
nand U7429 (N_7429,N_7383,N_7259);
or U7430 (N_7430,N_7204,N_7286);
nand U7431 (N_7431,N_7337,N_7330);
and U7432 (N_7432,N_7334,N_7359);
and U7433 (N_7433,N_7311,N_7281);
and U7434 (N_7434,N_7360,N_7316);
nor U7435 (N_7435,N_7239,N_7231);
and U7436 (N_7436,N_7279,N_7300);
xor U7437 (N_7437,N_7216,N_7246);
xnor U7438 (N_7438,N_7277,N_7368);
and U7439 (N_7439,N_7267,N_7381);
xor U7440 (N_7440,N_7304,N_7303);
xnor U7441 (N_7441,N_7367,N_7296);
xnor U7442 (N_7442,N_7214,N_7263);
and U7443 (N_7443,N_7228,N_7227);
nand U7444 (N_7444,N_7215,N_7338);
nand U7445 (N_7445,N_7354,N_7241);
xnor U7446 (N_7446,N_7313,N_7213);
xor U7447 (N_7447,N_7260,N_7388);
and U7448 (N_7448,N_7222,N_7329);
nand U7449 (N_7449,N_7221,N_7349);
xnor U7450 (N_7450,N_7265,N_7218);
or U7451 (N_7451,N_7219,N_7232);
or U7452 (N_7452,N_7317,N_7272);
nand U7453 (N_7453,N_7220,N_7201);
or U7454 (N_7454,N_7365,N_7230);
or U7455 (N_7455,N_7208,N_7264);
or U7456 (N_7456,N_7361,N_7211);
and U7457 (N_7457,N_7373,N_7210);
nand U7458 (N_7458,N_7238,N_7332);
nor U7459 (N_7459,N_7364,N_7229);
and U7460 (N_7460,N_7399,N_7207);
or U7461 (N_7461,N_7237,N_7288);
xnor U7462 (N_7462,N_7262,N_7380);
or U7463 (N_7463,N_7357,N_7234);
nor U7464 (N_7464,N_7318,N_7294);
nor U7465 (N_7465,N_7353,N_7306);
nor U7466 (N_7466,N_7284,N_7341);
xnor U7467 (N_7467,N_7278,N_7209);
nor U7468 (N_7468,N_7370,N_7385);
and U7469 (N_7469,N_7226,N_7255);
xnor U7470 (N_7470,N_7297,N_7310);
nand U7471 (N_7471,N_7331,N_7305);
and U7472 (N_7472,N_7327,N_7307);
or U7473 (N_7473,N_7275,N_7233);
xor U7474 (N_7474,N_7309,N_7371);
xor U7475 (N_7475,N_7252,N_7351);
nand U7476 (N_7476,N_7217,N_7242);
or U7477 (N_7477,N_7384,N_7378);
xor U7478 (N_7478,N_7322,N_7398);
nand U7479 (N_7479,N_7386,N_7396);
nor U7480 (N_7480,N_7282,N_7345);
or U7481 (N_7481,N_7397,N_7206);
and U7482 (N_7482,N_7356,N_7261);
nand U7483 (N_7483,N_7287,N_7244);
xor U7484 (N_7484,N_7225,N_7343);
and U7485 (N_7485,N_7325,N_7245);
nor U7486 (N_7486,N_7253,N_7324);
nor U7487 (N_7487,N_7251,N_7256);
nand U7488 (N_7488,N_7302,N_7276);
nand U7489 (N_7489,N_7363,N_7348);
and U7490 (N_7490,N_7271,N_7335);
nand U7491 (N_7491,N_7340,N_7301);
nor U7492 (N_7492,N_7346,N_7390);
or U7493 (N_7493,N_7321,N_7283);
nand U7494 (N_7494,N_7285,N_7355);
xor U7495 (N_7495,N_7328,N_7393);
or U7496 (N_7496,N_7280,N_7323);
nor U7497 (N_7497,N_7382,N_7392);
or U7498 (N_7498,N_7236,N_7376);
xnor U7499 (N_7499,N_7320,N_7273);
and U7500 (N_7500,N_7251,N_7343);
and U7501 (N_7501,N_7222,N_7396);
nor U7502 (N_7502,N_7212,N_7299);
and U7503 (N_7503,N_7334,N_7245);
nor U7504 (N_7504,N_7354,N_7306);
or U7505 (N_7505,N_7316,N_7248);
or U7506 (N_7506,N_7382,N_7204);
and U7507 (N_7507,N_7366,N_7252);
xnor U7508 (N_7508,N_7363,N_7372);
nor U7509 (N_7509,N_7301,N_7396);
nand U7510 (N_7510,N_7323,N_7321);
nor U7511 (N_7511,N_7320,N_7289);
xnor U7512 (N_7512,N_7283,N_7362);
and U7513 (N_7513,N_7286,N_7383);
nor U7514 (N_7514,N_7235,N_7351);
or U7515 (N_7515,N_7277,N_7263);
nor U7516 (N_7516,N_7264,N_7382);
nor U7517 (N_7517,N_7369,N_7263);
nor U7518 (N_7518,N_7243,N_7315);
or U7519 (N_7519,N_7318,N_7393);
and U7520 (N_7520,N_7252,N_7316);
or U7521 (N_7521,N_7337,N_7340);
and U7522 (N_7522,N_7292,N_7366);
xnor U7523 (N_7523,N_7366,N_7257);
nor U7524 (N_7524,N_7376,N_7383);
or U7525 (N_7525,N_7258,N_7351);
nor U7526 (N_7526,N_7246,N_7277);
and U7527 (N_7527,N_7218,N_7371);
nand U7528 (N_7528,N_7347,N_7253);
nand U7529 (N_7529,N_7345,N_7357);
nor U7530 (N_7530,N_7325,N_7298);
xnor U7531 (N_7531,N_7240,N_7201);
nor U7532 (N_7532,N_7344,N_7204);
nor U7533 (N_7533,N_7270,N_7282);
nand U7534 (N_7534,N_7302,N_7327);
nor U7535 (N_7535,N_7349,N_7297);
nor U7536 (N_7536,N_7355,N_7323);
nand U7537 (N_7537,N_7215,N_7235);
and U7538 (N_7538,N_7334,N_7299);
and U7539 (N_7539,N_7324,N_7276);
nand U7540 (N_7540,N_7379,N_7355);
and U7541 (N_7541,N_7323,N_7319);
or U7542 (N_7542,N_7397,N_7285);
nand U7543 (N_7543,N_7216,N_7242);
and U7544 (N_7544,N_7362,N_7253);
or U7545 (N_7545,N_7212,N_7355);
xor U7546 (N_7546,N_7323,N_7339);
or U7547 (N_7547,N_7386,N_7368);
and U7548 (N_7548,N_7341,N_7206);
nor U7549 (N_7549,N_7258,N_7260);
nor U7550 (N_7550,N_7345,N_7350);
or U7551 (N_7551,N_7282,N_7210);
xor U7552 (N_7552,N_7307,N_7398);
nor U7553 (N_7553,N_7242,N_7369);
and U7554 (N_7554,N_7300,N_7297);
nand U7555 (N_7555,N_7213,N_7397);
nor U7556 (N_7556,N_7342,N_7247);
xor U7557 (N_7557,N_7386,N_7286);
or U7558 (N_7558,N_7321,N_7343);
nand U7559 (N_7559,N_7314,N_7351);
and U7560 (N_7560,N_7204,N_7323);
and U7561 (N_7561,N_7259,N_7265);
nor U7562 (N_7562,N_7394,N_7230);
and U7563 (N_7563,N_7302,N_7230);
xor U7564 (N_7564,N_7327,N_7256);
nor U7565 (N_7565,N_7212,N_7354);
nand U7566 (N_7566,N_7334,N_7318);
xnor U7567 (N_7567,N_7262,N_7236);
or U7568 (N_7568,N_7330,N_7265);
nand U7569 (N_7569,N_7309,N_7304);
nand U7570 (N_7570,N_7274,N_7314);
nor U7571 (N_7571,N_7388,N_7308);
nand U7572 (N_7572,N_7281,N_7328);
xnor U7573 (N_7573,N_7274,N_7220);
and U7574 (N_7574,N_7229,N_7215);
and U7575 (N_7575,N_7324,N_7373);
xor U7576 (N_7576,N_7371,N_7372);
xnor U7577 (N_7577,N_7373,N_7357);
or U7578 (N_7578,N_7304,N_7240);
xor U7579 (N_7579,N_7269,N_7245);
nand U7580 (N_7580,N_7358,N_7369);
xnor U7581 (N_7581,N_7215,N_7397);
nand U7582 (N_7582,N_7369,N_7235);
nand U7583 (N_7583,N_7241,N_7388);
nand U7584 (N_7584,N_7289,N_7394);
or U7585 (N_7585,N_7245,N_7263);
nand U7586 (N_7586,N_7391,N_7226);
or U7587 (N_7587,N_7371,N_7287);
nand U7588 (N_7588,N_7231,N_7228);
nor U7589 (N_7589,N_7352,N_7217);
nand U7590 (N_7590,N_7303,N_7250);
nor U7591 (N_7591,N_7385,N_7247);
and U7592 (N_7592,N_7330,N_7240);
or U7593 (N_7593,N_7364,N_7231);
xor U7594 (N_7594,N_7300,N_7227);
or U7595 (N_7595,N_7364,N_7345);
and U7596 (N_7596,N_7222,N_7321);
nor U7597 (N_7597,N_7223,N_7205);
nor U7598 (N_7598,N_7310,N_7314);
and U7599 (N_7599,N_7320,N_7305);
or U7600 (N_7600,N_7443,N_7445);
nor U7601 (N_7601,N_7418,N_7483);
nor U7602 (N_7602,N_7538,N_7495);
and U7603 (N_7603,N_7539,N_7488);
nand U7604 (N_7604,N_7407,N_7459);
nor U7605 (N_7605,N_7440,N_7437);
nand U7606 (N_7606,N_7468,N_7569);
and U7607 (N_7607,N_7419,N_7500);
nor U7608 (N_7608,N_7586,N_7560);
or U7609 (N_7609,N_7401,N_7400);
nand U7610 (N_7610,N_7518,N_7472);
and U7611 (N_7611,N_7572,N_7589);
xor U7612 (N_7612,N_7416,N_7411);
xnor U7613 (N_7613,N_7446,N_7458);
and U7614 (N_7614,N_7563,N_7480);
and U7615 (N_7615,N_7596,N_7566);
nand U7616 (N_7616,N_7575,N_7425);
and U7617 (N_7617,N_7512,N_7581);
xnor U7618 (N_7618,N_7421,N_7436);
or U7619 (N_7619,N_7417,N_7453);
or U7620 (N_7620,N_7490,N_7456);
nand U7621 (N_7621,N_7404,N_7501);
xnor U7622 (N_7622,N_7576,N_7460);
or U7623 (N_7623,N_7561,N_7502);
and U7624 (N_7624,N_7597,N_7565);
nor U7625 (N_7625,N_7499,N_7476);
nor U7626 (N_7626,N_7588,N_7598);
and U7627 (N_7627,N_7537,N_7442);
and U7628 (N_7628,N_7454,N_7599);
and U7629 (N_7629,N_7414,N_7415);
xnor U7630 (N_7630,N_7571,N_7543);
and U7631 (N_7631,N_7494,N_7550);
xor U7632 (N_7632,N_7595,N_7420);
xnor U7633 (N_7633,N_7583,N_7525);
nand U7634 (N_7634,N_7528,N_7529);
and U7635 (N_7635,N_7405,N_7463);
nand U7636 (N_7636,N_7481,N_7562);
and U7637 (N_7637,N_7582,N_7424);
nor U7638 (N_7638,N_7467,N_7465);
nand U7639 (N_7639,N_7558,N_7574);
nand U7640 (N_7640,N_7451,N_7505);
xor U7641 (N_7641,N_7409,N_7428);
nand U7642 (N_7642,N_7448,N_7457);
xor U7643 (N_7643,N_7504,N_7497);
nand U7644 (N_7644,N_7520,N_7506);
and U7645 (N_7645,N_7542,N_7473);
nand U7646 (N_7646,N_7461,N_7439);
or U7647 (N_7647,N_7489,N_7491);
nor U7648 (N_7648,N_7475,N_7515);
xnor U7649 (N_7649,N_7464,N_7485);
xor U7650 (N_7650,N_7477,N_7547);
nand U7651 (N_7651,N_7568,N_7553);
xor U7652 (N_7652,N_7555,N_7482);
or U7653 (N_7653,N_7503,N_7513);
xor U7654 (N_7654,N_7527,N_7402);
nand U7655 (N_7655,N_7554,N_7498);
or U7656 (N_7656,N_7590,N_7549);
or U7657 (N_7657,N_7429,N_7523);
and U7658 (N_7658,N_7447,N_7544);
and U7659 (N_7659,N_7423,N_7536);
or U7660 (N_7660,N_7531,N_7511);
nand U7661 (N_7661,N_7517,N_7470);
and U7662 (N_7662,N_7551,N_7533);
or U7663 (N_7663,N_7514,N_7532);
xor U7664 (N_7664,N_7435,N_7430);
xnor U7665 (N_7665,N_7557,N_7434);
or U7666 (N_7666,N_7594,N_7508);
or U7667 (N_7667,N_7541,N_7530);
and U7668 (N_7668,N_7432,N_7493);
nor U7669 (N_7669,N_7535,N_7593);
or U7670 (N_7670,N_7492,N_7585);
xor U7671 (N_7671,N_7471,N_7486);
and U7672 (N_7672,N_7408,N_7534);
and U7673 (N_7673,N_7570,N_7526);
nand U7674 (N_7674,N_7478,N_7487);
and U7675 (N_7675,N_7496,N_7591);
xnor U7676 (N_7676,N_7444,N_7556);
nor U7677 (N_7677,N_7559,N_7573);
xnor U7678 (N_7678,N_7579,N_7412);
nor U7679 (N_7679,N_7507,N_7433);
xor U7680 (N_7680,N_7431,N_7592);
nand U7681 (N_7681,N_7509,N_7438);
and U7682 (N_7682,N_7450,N_7462);
xor U7683 (N_7683,N_7422,N_7427);
nand U7684 (N_7684,N_7545,N_7546);
nand U7685 (N_7685,N_7577,N_7426);
or U7686 (N_7686,N_7466,N_7455);
or U7687 (N_7687,N_7548,N_7584);
xnor U7688 (N_7688,N_7410,N_7403);
nand U7689 (N_7689,N_7452,N_7567);
nor U7690 (N_7690,N_7522,N_7484);
xnor U7691 (N_7691,N_7449,N_7441);
or U7692 (N_7692,N_7413,N_7524);
or U7693 (N_7693,N_7587,N_7519);
and U7694 (N_7694,N_7580,N_7406);
xor U7695 (N_7695,N_7474,N_7516);
xor U7696 (N_7696,N_7469,N_7479);
and U7697 (N_7697,N_7521,N_7564);
nand U7698 (N_7698,N_7510,N_7552);
or U7699 (N_7699,N_7540,N_7578);
or U7700 (N_7700,N_7561,N_7401);
or U7701 (N_7701,N_7487,N_7406);
nand U7702 (N_7702,N_7439,N_7417);
nor U7703 (N_7703,N_7552,N_7520);
nor U7704 (N_7704,N_7410,N_7454);
nand U7705 (N_7705,N_7557,N_7401);
nor U7706 (N_7706,N_7432,N_7474);
nor U7707 (N_7707,N_7509,N_7417);
xnor U7708 (N_7708,N_7461,N_7559);
xor U7709 (N_7709,N_7575,N_7557);
nor U7710 (N_7710,N_7568,N_7595);
nor U7711 (N_7711,N_7573,N_7548);
or U7712 (N_7712,N_7549,N_7579);
nand U7713 (N_7713,N_7561,N_7518);
and U7714 (N_7714,N_7492,N_7434);
and U7715 (N_7715,N_7524,N_7539);
and U7716 (N_7716,N_7519,N_7412);
nor U7717 (N_7717,N_7472,N_7474);
and U7718 (N_7718,N_7464,N_7434);
xor U7719 (N_7719,N_7446,N_7592);
and U7720 (N_7720,N_7541,N_7574);
xor U7721 (N_7721,N_7409,N_7568);
nor U7722 (N_7722,N_7559,N_7419);
or U7723 (N_7723,N_7546,N_7547);
and U7724 (N_7724,N_7405,N_7480);
nor U7725 (N_7725,N_7420,N_7425);
and U7726 (N_7726,N_7481,N_7441);
nor U7727 (N_7727,N_7527,N_7565);
nand U7728 (N_7728,N_7574,N_7466);
nand U7729 (N_7729,N_7497,N_7488);
and U7730 (N_7730,N_7526,N_7450);
and U7731 (N_7731,N_7455,N_7479);
and U7732 (N_7732,N_7538,N_7542);
xnor U7733 (N_7733,N_7517,N_7574);
xor U7734 (N_7734,N_7583,N_7427);
nand U7735 (N_7735,N_7596,N_7597);
xnor U7736 (N_7736,N_7548,N_7528);
and U7737 (N_7737,N_7589,N_7416);
nor U7738 (N_7738,N_7517,N_7516);
and U7739 (N_7739,N_7562,N_7455);
nand U7740 (N_7740,N_7555,N_7437);
xnor U7741 (N_7741,N_7437,N_7414);
xor U7742 (N_7742,N_7513,N_7423);
nor U7743 (N_7743,N_7547,N_7500);
or U7744 (N_7744,N_7479,N_7543);
nand U7745 (N_7745,N_7402,N_7414);
xor U7746 (N_7746,N_7422,N_7576);
nand U7747 (N_7747,N_7598,N_7597);
nor U7748 (N_7748,N_7587,N_7528);
nand U7749 (N_7749,N_7503,N_7562);
or U7750 (N_7750,N_7557,N_7536);
nand U7751 (N_7751,N_7518,N_7500);
or U7752 (N_7752,N_7587,N_7538);
xnor U7753 (N_7753,N_7402,N_7577);
or U7754 (N_7754,N_7567,N_7465);
nor U7755 (N_7755,N_7427,N_7460);
xnor U7756 (N_7756,N_7483,N_7536);
xor U7757 (N_7757,N_7585,N_7530);
xnor U7758 (N_7758,N_7598,N_7539);
and U7759 (N_7759,N_7555,N_7439);
or U7760 (N_7760,N_7503,N_7480);
or U7761 (N_7761,N_7422,N_7477);
or U7762 (N_7762,N_7549,N_7447);
nor U7763 (N_7763,N_7547,N_7464);
nor U7764 (N_7764,N_7526,N_7485);
and U7765 (N_7765,N_7549,N_7432);
xnor U7766 (N_7766,N_7559,N_7563);
or U7767 (N_7767,N_7547,N_7431);
xor U7768 (N_7768,N_7528,N_7431);
and U7769 (N_7769,N_7498,N_7424);
nand U7770 (N_7770,N_7548,N_7431);
or U7771 (N_7771,N_7582,N_7551);
xor U7772 (N_7772,N_7471,N_7477);
or U7773 (N_7773,N_7535,N_7487);
xnor U7774 (N_7774,N_7480,N_7417);
xnor U7775 (N_7775,N_7593,N_7434);
xor U7776 (N_7776,N_7529,N_7426);
nand U7777 (N_7777,N_7572,N_7483);
nand U7778 (N_7778,N_7576,N_7440);
xnor U7779 (N_7779,N_7491,N_7472);
or U7780 (N_7780,N_7483,N_7577);
nand U7781 (N_7781,N_7454,N_7525);
nand U7782 (N_7782,N_7463,N_7545);
xnor U7783 (N_7783,N_7563,N_7436);
nand U7784 (N_7784,N_7442,N_7590);
nor U7785 (N_7785,N_7565,N_7548);
xor U7786 (N_7786,N_7578,N_7431);
and U7787 (N_7787,N_7415,N_7491);
xor U7788 (N_7788,N_7455,N_7426);
nand U7789 (N_7789,N_7463,N_7462);
xor U7790 (N_7790,N_7565,N_7493);
nand U7791 (N_7791,N_7519,N_7441);
or U7792 (N_7792,N_7579,N_7403);
nand U7793 (N_7793,N_7572,N_7480);
nand U7794 (N_7794,N_7553,N_7458);
nand U7795 (N_7795,N_7513,N_7474);
nor U7796 (N_7796,N_7462,N_7431);
nand U7797 (N_7797,N_7483,N_7544);
or U7798 (N_7798,N_7487,N_7529);
nor U7799 (N_7799,N_7550,N_7405);
nor U7800 (N_7800,N_7796,N_7670);
nor U7801 (N_7801,N_7698,N_7658);
nor U7802 (N_7802,N_7765,N_7706);
xor U7803 (N_7803,N_7692,N_7641);
xor U7804 (N_7804,N_7666,N_7775);
and U7805 (N_7805,N_7678,N_7680);
or U7806 (N_7806,N_7699,N_7713);
or U7807 (N_7807,N_7710,N_7615);
and U7808 (N_7808,N_7746,N_7601);
and U7809 (N_7809,N_7629,N_7628);
and U7810 (N_7810,N_7669,N_7744);
nand U7811 (N_7811,N_7657,N_7738);
xnor U7812 (N_7812,N_7704,N_7762);
and U7813 (N_7813,N_7603,N_7777);
nand U7814 (N_7814,N_7697,N_7650);
xnor U7815 (N_7815,N_7694,N_7696);
nor U7816 (N_7816,N_7779,N_7683);
nand U7817 (N_7817,N_7639,N_7723);
or U7818 (N_7818,N_7667,N_7722);
and U7819 (N_7819,N_7621,N_7761);
xnor U7820 (N_7820,N_7663,N_7613);
xor U7821 (N_7821,N_7673,N_7788);
and U7822 (N_7822,N_7693,N_7612);
nand U7823 (N_7823,N_7703,N_7783);
nor U7824 (N_7824,N_7770,N_7748);
xor U7825 (N_7825,N_7634,N_7790);
nor U7826 (N_7826,N_7707,N_7773);
nor U7827 (N_7827,N_7672,N_7757);
xor U7828 (N_7828,N_7646,N_7600);
or U7829 (N_7829,N_7712,N_7637);
nand U7830 (N_7830,N_7732,N_7671);
nand U7831 (N_7831,N_7763,N_7635);
nor U7832 (N_7832,N_7774,N_7797);
and U7833 (N_7833,N_7660,N_7614);
or U7834 (N_7834,N_7617,N_7794);
or U7835 (N_7835,N_7632,N_7688);
or U7836 (N_7836,N_7681,N_7709);
nor U7837 (N_7837,N_7686,N_7760);
or U7838 (N_7838,N_7750,N_7656);
and U7839 (N_7839,N_7653,N_7647);
and U7840 (N_7840,N_7636,N_7605);
xnor U7841 (N_7841,N_7778,N_7714);
nor U7842 (N_7842,N_7684,N_7737);
nor U7843 (N_7843,N_7786,N_7745);
or U7844 (N_7844,N_7649,N_7608);
nor U7845 (N_7845,N_7791,N_7662);
xnor U7846 (N_7846,N_7741,N_7611);
nor U7847 (N_7847,N_7652,N_7640);
nor U7848 (N_7848,N_7715,N_7785);
nand U7849 (N_7849,N_7767,N_7659);
or U7850 (N_7850,N_7645,N_7727);
nand U7851 (N_7851,N_7734,N_7701);
and U7852 (N_7852,N_7695,N_7622);
xnor U7853 (N_7853,N_7609,N_7759);
xor U7854 (N_7854,N_7771,N_7766);
xnor U7855 (N_7855,N_7716,N_7780);
nor U7856 (N_7856,N_7730,N_7633);
or U7857 (N_7857,N_7643,N_7642);
and U7858 (N_7858,N_7674,N_7793);
and U7859 (N_7859,N_7784,N_7644);
nor U7860 (N_7860,N_7720,N_7756);
nand U7861 (N_7861,N_7717,N_7736);
nand U7862 (N_7862,N_7625,N_7795);
nor U7863 (N_7863,N_7731,N_7626);
and U7864 (N_7864,N_7725,N_7690);
nor U7865 (N_7865,N_7739,N_7792);
xor U7866 (N_7866,N_7751,N_7787);
nand U7867 (N_7867,N_7638,N_7768);
nor U7868 (N_7868,N_7618,N_7616);
xor U7869 (N_7869,N_7679,N_7799);
xor U7870 (N_7870,N_7675,N_7747);
and U7871 (N_7871,N_7721,N_7664);
nand U7872 (N_7872,N_7781,N_7718);
or U7873 (N_7873,N_7606,N_7753);
nand U7874 (N_7874,N_7798,N_7677);
or U7875 (N_7875,N_7602,N_7772);
xor U7876 (N_7876,N_7676,N_7607);
xnor U7877 (N_7877,N_7789,N_7654);
and U7878 (N_7878,N_7700,N_7687);
and U7879 (N_7879,N_7729,N_7719);
and U7880 (N_7880,N_7758,N_7702);
and U7881 (N_7881,N_7776,N_7631);
nand U7882 (N_7882,N_7769,N_7752);
nor U7883 (N_7883,N_7754,N_7742);
xor U7884 (N_7884,N_7661,N_7764);
nor U7885 (N_7885,N_7623,N_7735);
and U7886 (N_7886,N_7749,N_7627);
nand U7887 (N_7887,N_7620,N_7743);
and U7888 (N_7888,N_7691,N_7651);
and U7889 (N_7889,N_7711,N_7705);
nand U7890 (N_7890,N_7708,N_7728);
nand U7891 (N_7891,N_7755,N_7624);
nor U7892 (N_7892,N_7733,N_7648);
and U7893 (N_7893,N_7782,N_7619);
nor U7894 (N_7894,N_7668,N_7682);
or U7895 (N_7895,N_7610,N_7655);
xnor U7896 (N_7896,N_7630,N_7740);
nand U7897 (N_7897,N_7604,N_7724);
nor U7898 (N_7898,N_7726,N_7685);
or U7899 (N_7899,N_7689,N_7665);
xnor U7900 (N_7900,N_7714,N_7659);
nand U7901 (N_7901,N_7743,N_7765);
nor U7902 (N_7902,N_7654,N_7703);
xor U7903 (N_7903,N_7757,N_7785);
and U7904 (N_7904,N_7620,N_7765);
xnor U7905 (N_7905,N_7660,N_7609);
nor U7906 (N_7906,N_7654,N_7725);
nand U7907 (N_7907,N_7678,N_7740);
xor U7908 (N_7908,N_7604,N_7673);
or U7909 (N_7909,N_7731,N_7676);
and U7910 (N_7910,N_7644,N_7739);
nor U7911 (N_7911,N_7715,N_7716);
or U7912 (N_7912,N_7628,N_7600);
and U7913 (N_7913,N_7713,N_7781);
nand U7914 (N_7914,N_7629,N_7670);
or U7915 (N_7915,N_7772,N_7600);
or U7916 (N_7916,N_7629,N_7633);
nand U7917 (N_7917,N_7627,N_7606);
and U7918 (N_7918,N_7649,N_7701);
or U7919 (N_7919,N_7680,N_7760);
or U7920 (N_7920,N_7771,N_7656);
nor U7921 (N_7921,N_7785,N_7608);
xor U7922 (N_7922,N_7689,N_7638);
xor U7923 (N_7923,N_7701,N_7797);
and U7924 (N_7924,N_7797,N_7616);
nand U7925 (N_7925,N_7642,N_7698);
nor U7926 (N_7926,N_7647,N_7671);
and U7927 (N_7927,N_7617,N_7603);
nand U7928 (N_7928,N_7704,N_7618);
xor U7929 (N_7929,N_7621,N_7627);
nor U7930 (N_7930,N_7770,N_7772);
or U7931 (N_7931,N_7697,N_7639);
and U7932 (N_7932,N_7660,N_7684);
nor U7933 (N_7933,N_7744,N_7633);
and U7934 (N_7934,N_7793,N_7702);
nand U7935 (N_7935,N_7773,N_7665);
nor U7936 (N_7936,N_7635,N_7663);
nor U7937 (N_7937,N_7794,N_7636);
or U7938 (N_7938,N_7718,N_7647);
nand U7939 (N_7939,N_7705,N_7662);
nor U7940 (N_7940,N_7789,N_7745);
xor U7941 (N_7941,N_7781,N_7659);
nand U7942 (N_7942,N_7716,N_7718);
nor U7943 (N_7943,N_7722,N_7621);
and U7944 (N_7944,N_7778,N_7715);
or U7945 (N_7945,N_7709,N_7706);
nor U7946 (N_7946,N_7705,N_7791);
and U7947 (N_7947,N_7617,N_7761);
xnor U7948 (N_7948,N_7693,N_7728);
or U7949 (N_7949,N_7656,N_7794);
or U7950 (N_7950,N_7777,N_7710);
or U7951 (N_7951,N_7654,N_7709);
nor U7952 (N_7952,N_7667,N_7726);
xnor U7953 (N_7953,N_7792,N_7755);
or U7954 (N_7954,N_7657,N_7651);
xnor U7955 (N_7955,N_7763,N_7776);
xnor U7956 (N_7956,N_7628,N_7625);
or U7957 (N_7957,N_7605,N_7736);
or U7958 (N_7958,N_7623,N_7674);
nor U7959 (N_7959,N_7762,N_7786);
and U7960 (N_7960,N_7614,N_7777);
and U7961 (N_7961,N_7729,N_7602);
and U7962 (N_7962,N_7785,N_7774);
and U7963 (N_7963,N_7604,N_7703);
nor U7964 (N_7964,N_7722,N_7798);
or U7965 (N_7965,N_7667,N_7671);
and U7966 (N_7966,N_7779,N_7602);
and U7967 (N_7967,N_7682,N_7713);
or U7968 (N_7968,N_7639,N_7620);
nor U7969 (N_7969,N_7630,N_7680);
xnor U7970 (N_7970,N_7662,N_7784);
nor U7971 (N_7971,N_7783,N_7689);
or U7972 (N_7972,N_7739,N_7795);
nor U7973 (N_7973,N_7722,N_7700);
xnor U7974 (N_7974,N_7654,N_7683);
and U7975 (N_7975,N_7765,N_7758);
nor U7976 (N_7976,N_7692,N_7619);
nor U7977 (N_7977,N_7700,N_7661);
nor U7978 (N_7978,N_7766,N_7687);
or U7979 (N_7979,N_7632,N_7610);
nor U7980 (N_7980,N_7784,N_7724);
nor U7981 (N_7981,N_7783,N_7603);
or U7982 (N_7982,N_7671,N_7698);
nor U7983 (N_7983,N_7643,N_7777);
nor U7984 (N_7984,N_7649,N_7749);
and U7985 (N_7985,N_7782,N_7769);
xnor U7986 (N_7986,N_7792,N_7686);
nand U7987 (N_7987,N_7719,N_7782);
xor U7988 (N_7988,N_7617,N_7786);
nor U7989 (N_7989,N_7767,N_7777);
nand U7990 (N_7990,N_7698,N_7741);
nand U7991 (N_7991,N_7757,N_7751);
xnor U7992 (N_7992,N_7781,N_7649);
nand U7993 (N_7993,N_7707,N_7695);
nand U7994 (N_7994,N_7704,N_7634);
and U7995 (N_7995,N_7693,N_7712);
and U7996 (N_7996,N_7750,N_7622);
xnor U7997 (N_7997,N_7796,N_7791);
nor U7998 (N_7998,N_7748,N_7714);
nand U7999 (N_7999,N_7764,N_7788);
nand U8000 (N_8000,N_7808,N_7938);
nand U8001 (N_8001,N_7959,N_7936);
and U8002 (N_8002,N_7885,N_7926);
nor U8003 (N_8003,N_7937,N_7825);
and U8004 (N_8004,N_7854,N_7864);
or U8005 (N_8005,N_7816,N_7848);
or U8006 (N_8006,N_7916,N_7985);
nand U8007 (N_8007,N_7987,N_7895);
and U8008 (N_8008,N_7993,N_7878);
nand U8009 (N_8009,N_7939,N_7844);
xor U8010 (N_8010,N_7857,N_7845);
nor U8011 (N_8011,N_7929,N_7822);
nor U8012 (N_8012,N_7823,N_7982);
xor U8013 (N_8013,N_7968,N_7973);
nand U8014 (N_8014,N_7818,N_7974);
or U8015 (N_8015,N_7839,N_7914);
or U8016 (N_8016,N_7947,N_7998);
and U8017 (N_8017,N_7986,N_7874);
nor U8018 (N_8018,N_7897,N_7828);
and U8019 (N_8019,N_7882,N_7837);
xnor U8020 (N_8020,N_7963,N_7852);
and U8021 (N_8021,N_7975,N_7856);
or U8022 (N_8022,N_7924,N_7892);
and U8023 (N_8023,N_7912,N_7909);
nor U8024 (N_8024,N_7957,N_7863);
or U8025 (N_8025,N_7832,N_7930);
xor U8026 (N_8026,N_7813,N_7950);
and U8027 (N_8027,N_7884,N_7902);
and U8028 (N_8028,N_7996,N_7880);
xnor U8029 (N_8029,N_7978,N_7908);
nand U8030 (N_8030,N_7964,N_7955);
or U8031 (N_8031,N_7980,N_7949);
nand U8032 (N_8032,N_7875,N_7919);
nand U8033 (N_8033,N_7969,N_7981);
and U8034 (N_8034,N_7960,N_7802);
and U8035 (N_8035,N_7846,N_7862);
nand U8036 (N_8036,N_7925,N_7858);
xor U8037 (N_8037,N_7948,N_7977);
and U8038 (N_8038,N_7941,N_7876);
and U8039 (N_8039,N_7867,N_7850);
nand U8040 (N_8040,N_7965,N_7951);
xnor U8041 (N_8041,N_7992,N_7915);
and U8042 (N_8042,N_7967,N_7803);
xor U8043 (N_8043,N_7983,N_7944);
nand U8044 (N_8044,N_7801,N_7994);
and U8045 (N_8045,N_7971,N_7866);
nand U8046 (N_8046,N_7810,N_7942);
and U8047 (N_8047,N_7997,N_7806);
nor U8048 (N_8048,N_7905,N_7860);
and U8049 (N_8049,N_7855,N_7952);
or U8050 (N_8050,N_7946,N_7879);
nand U8051 (N_8051,N_7899,N_7827);
nor U8052 (N_8052,N_7907,N_7889);
nor U8053 (N_8053,N_7826,N_7901);
nor U8054 (N_8054,N_7920,N_7958);
nor U8055 (N_8055,N_7881,N_7928);
nand U8056 (N_8056,N_7972,N_7887);
and U8057 (N_8057,N_7976,N_7868);
or U8058 (N_8058,N_7811,N_7872);
xor U8059 (N_8059,N_7888,N_7898);
nor U8060 (N_8060,N_7851,N_7979);
xor U8061 (N_8061,N_7989,N_7804);
nand U8062 (N_8062,N_7849,N_7913);
nor U8063 (N_8063,N_7865,N_7900);
nand U8064 (N_8064,N_7841,N_7814);
nand U8065 (N_8065,N_7800,N_7896);
nand U8066 (N_8066,N_7940,N_7954);
nand U8067 (N_8067,N_7932,N_7861);
nand U8068 (N_8068,N_7931,N_7830);
nor U8069 (N_8069,N_7836,N_7923);
nor U8070 (N_8070,N_7821,N_7945);
and U8071 (N_8071,N_7935,N_7918);
xor U8072 (N_8072,N_7877,N_7921);
and U8073 (N_8073,N_7999,N_7873);
nor U8074 (N_8074,N_7893,N_7812);
nand U8075 (N_8075,N_7838,N_7995);
or U8076 (N_8076,N_7934,N_7831);
and U8077 (N_8077,N_7890,N_7817);
xor U8078 (N_8078,N_7953,N_7962);
xnor U8079 (N_8079,N_7966,N_7943);
or U8080 (N_8080,N_7815,N_7933);
nand U8081 (N_8081,N_7886,N_7956);
and U8082 (N_8082,N_7805,N_7984);
nor U8083 (N_8083,N_7835,N_7961);
nor U8084 (N_8084,N_7869,N_7883);
nor U8085 (N_8085,N_7809,N_7904);
or U8086 (N_8086,N_7847,N_7894);
nand U8087 (N_8087,N_7807,N_7988);
or U8088 (N_8088,N_7829,N_7824);
nor U8089 (N_8089,N_7840,N_7871);
nor U8090 (N_8090,N_7922,N_7990);
or U8091 (N_8091,N_7833,N_7917);
xor U8092 (N_8092,N_7820,N_7891);
nor U8093 (N_8093,N_7911,N_7870);
nor U8094 (N_8094,N_7842,N_7991);
or U8095 (N_8095,N_7927,N_7910);
xnor U8096 (N_8096,N_7819,N_7843);
or U8097 (N_8097,N_7970,N_7903);
xor U8098 (N_8098,N_7853,N_7906);
nand U8099 (N_8099,N_7859,N_7834);
nand U8100 (N_8100,N_7965,N_7980);
or U8101 (N_8101,N_7895,N_7970);
nor U8102 (N_8102,N_7996,N_7824);
nor U8103 (N_8103,N_7952,N_7896);
nor U8104 (N_8104,N_7835,N_7871);
nand U8105 (N_8105,N_7929,N_7906);
nand U8106 (N_8106,N_7884,N_7907);
nand U8107 (N_8107,N_7978,N_7822);
xor U8108 (N_8108,N_7994,N_7802);
xor U8109 (N_8109,N_7898,N_7843);
xnor U8110 (N_8110,N_7884,N_7896);
or U8111 (N_8111,N_7902,N_7939);
and U8112 (N_8112,N_7891,N_7906);
nand U8113 (N_8113,N_7908,N_7867);
nor U8114 (N_8114,N_7861,N_7809);
xnor U8115 (N_8115,N_7888,N_7940);
and U8116 (N_8116,N_7895,N_7853);
nand U8117 (N_8117,N_7900,N_7983);
and U8118 (N_8118,N_7932,N_7801);
and U8119 (N_8119,N_7958,N_7971);
xor U8120 (N_8120,N_7824,N_7831);
xor U8121 (N_8121,N_7978,N_7944);
nand U8122 (N_8122,N_7983,N_7963);
and U8123 (N_8123,N_7825,N_7927);
and U8124 (N_8124,N_7901,N_7914);
nand U8125 (N_8125,N_7816,N_7861);
or U8126 (N_8126,N_7989,N_7935);
or U8127 (N_8127,N_7855,N_7890);
or U8128 (N_8128,N_7959,N_7906);
or U8129 (N_8129,N_7947,N_7863);
and U8130 (N_8130,N_7835,N_7840);
and U8131 (N_8131,N_7992,N_7905);
xnor U8132 (N_8132,N_7937,N_7836);
xor U8133 (N_8133,N_7802,N_7978);
xnor U8134 (N_8134,N_7828,N_7802);
xor U8135 (N_8135,N_7942,N_7863);
and U8136 (N_8136,N_7895,N_7856);
xnor U8137 (N_8137,N_7998,N_7916);
xor U8138 (N_8138,N_7825,N_7832);
or U8139 (N_8139,N_7998,N_7893);
or U8140 (N_8140,N_7872,N_7813);
nand U8141 (N_8141,N_7972,N_7812);
nor U8142 (N_8142,N_7998,N_7920);
nand U8143 (N_8143,N_7849,N_7945);
or U8144 (N_8144,N_7997,N_7966);
nand U8145 (N_8145,N_7851,N_7871);
and U8146 (N_8146,N_7887,N_7940);
nor U8147 (N_8147,N_7930,N_7961);
nand U8148 (N_8148,N_7820,N_7906);
nand U8149 (N_8149,N_7995,N_7816);
nor U8150 (N_8150,N_7901,N_7994);
xnor U8151 (N_8151,N_7842,N_7829);
and U8152 (N_8152,N_7855,N_7893);
nor U8153 (N_8153,N_7976,N_7834);
nand U8154 (N_8154,N_7869,N_7840);
and U8155 (N_8155,N_7829,N_7856);
nand U8156 (N_8156,N_7827,N_7986);
nand U8157 (N_8157,N_7855,N_7847);
nand U8158 (N_8158,N_7819,N_7870);
and U8159 (N_8159,N_7877,N_7900);
nand U8160 (N_8160,N_7873,N_7978);
nor U8161 (N_8161,N_7907,N_7978);
nor U8162 (N_8162,N_7998,N_7800);
nor U8163 (N_8163,N_7984,N_7858);
or U8164 (N_8164,N_7869,N_7952);
nand U8165 (N_8165,N_7986,N_7802);
xnor U8166 (N_8166,N_7882,N_7904);
xor U8167 (N_8167,N_7840,N_7939);
nand U8168 (N_8168,N_7803,N_7816);
xnor U8169 (N_8169,N_7870,N_7868);
nor U8170 (N_8170,N_7827,N_7883);
nor U8171 (N_8171,N_7866,N_7807);
or U8172 (N_8172,N_7994,N_7890);
and U8173 (N_8173,N_7842,N_7875);
xor U8174 (N_8174,N_7916,N_7983);
or U8175 (N_8175,N_7913,N_7950);
nand U8176 (N_8176,N_7831,N_7995);
nor U8177 (N_8177,N_7936,N_7836);
xor U8178 (N_8178,N_7834,N_7818);
or U8179 (N_8179,N_7995,N_7864);
xnor U8180 (N_8180,N_7834,N_7831);
nor U8181 (N_8181,N_7966,N_7916);
or U8182 (N_8182,N_7842,N_7928);
nand U8183 (N_8183,N_7868,N_7907);
nor U8184 (N_8184,N_7847,N_7808);
nand U8185 (N_8185,N_7807,N_7849);
xor U8186 (N_8186,N_7983,N_7859);
nand U8187 (N_8187,N_7999,N_7980);
and U8188 (N_8188,N_7866,N_7802);
and U8189 (N_8189,N_7858,N_7924);
nor U8190 (N_8190,N_7867,N_7954);
nand U8191 (N_8191,N_7978,N_7888);
or U8192 (N_8192,N_7891,N_7853);
nor U8193 (N_8193,N_7821,N_7990);
nor U8194 (N_8194,N_7964,N_7936);
nor U8195 (N_8195,N_7898,N_7969);
and U8196 (N_8196,N_7916,N_7878);
nor U8197 (N_8197,N_7947,N_7938);
nand U8198 (N_8198,N_7858,N_7849);
or U8199 (N_8199,N_7868,N_7846);
or U8200 (N_8200,N_8117,N_8055);
and U8201 (N_8201,N_8161,N_8033);
nor U8202 (N_8202,N_8164,N_8029);
nand U8203 (N_8203,N_8036,N_8076);
or U8204 (N_8204,N_8183,N_8054);
or U8205 (N_8205,N_8166,N_8048);
and U8206 (N_8206,N_8063,N_8195);
and U8207 (N_8207,N_8101,N_8157);
xor U8208 (N_8208,N_8069,N_8008);
xnor U8209 (N_8209,N_8023,N_8169);
nor U8210 (N_8210,N_8049,N_8094);
or U8211 (N_8211,N_8077,N_8090);
and U8212 (N_8212,N_8188,N_8072);
and U8213 (N_8213,N_8056,N_8139);
and U8214 (N_8214,N_8122,N_8022);
nor U8215 (N_8215,N_8159,N_8154);
and U8216 (N_8216,N_8126,N_8129);
xor U8217 (N_8217,N_8071,N_8019);
and U8218 (N_8218,N_8024,N_8107);
nor U8219 (N_8219,N_8050,N_8011);
nand U8220 (N_8220,N_8026,N_8199);
nand U8221 (N_8221,N_8184,N_8091);
xnor U8222 (N_8222,N_8124,N_8088);
nor U8223 (N_8223,N_8138,N_8046);
xnor U8224 (N_8224,N_8189,N_8162);
and U8225 (N_8225,N_8194,N_8001);
and U8226 (N_8226,N_8173,N_8143);
nor U8227 (N_8227,N_8160,N_8016);
nor U8228 (N_8228,N_8137,N_8178);
and U8229 (N_8229,N_8070,N_8153);
and U8230 (N_8230,N_8105,N_8040);
nor U8231 (N_8231,N_8074,N_8096);
and U8232 (N_8232,N_8131,N_8085);
or U8233 (N_8233,N_8065,N_8197);
nor U8234 (N_8234,N_8167,N_8191);
nor U8235 (N_8235,N_8052,N_8079);
or U8236 (N_8236,N_8186,N_8089);
xor U8237 (N_8237,N_8015,N_8087);
or U8238 (N_8238,N_8141,N_8192);
or U8239 (N_8239,N_8041,N_8047);
xnor U8240 (N_8240,N_8039,N_8032);
nor U8241 (N_8241,N_8151,N_8140);
and U8242 (N_8242,N_8013,N_8163);
xnor U8243 (N_8243,N_8042,N_8142);
xor U8244 (N_8244,N_8007,N_8043);
or U8245 (N_8245,N_8181,N_8004);
nor U8246 (N_8246,N_8044,N_8168);
nor U8247 (N_8247,N_8171,N_8100);
and U8248 (N_8248,N_8187,N_8034);
nand U8249 (N_8249,N_8095,N_8185);
nand U8250 (N_8250,N_8083,N_8175);
nor U8251 (N_8251,N_8064,N_8182);
nand U8252 (N_8252,N_8067,N_8086);
or U8253 (N_8253,N_8146,N_8093);
nor U8254 (N_8254,N_8104,N_8002);
nand U8255 (N_8255,N_8196,N_8062);
nand U8256 (N_8256,N_8156,N_8014);
xnor U8257 (N_8257,N_8118,N_8025);
nand U8258 (N_8258,N_8111,N_8073);
nor U8259 (N_8259,N_8198,N_8174);
or U8260 (N_8260,N_8149,N_8123);
and U8261 (N_8261,N_8028,N_8098);
and U8262 (N_8262,N_8158,N_8106);
xor U8263 (N_8263,N_8078,N_8132);
nand U8264 (N_8264,N_8080,N_8119);
nand U8265 (N_8265,N_8128,N_8010);
or U8266 (N_8266,N_8003,N_8155);
and U8267 (N_8267,N_8103,N_8190);
and U8268 (N_8268,N_8099,N_8031);
nor U8269 (N_8269,N_8021,N_8136);
nand U8270 (N_8270,N_8000,N_8006);
xnor U8271 (N_8271,N_8017,N_8113);
and U8272 (N_8272,N_8179,N_8012);
or U8273 (N_8273,N_8152,N_8145);
nor U8274 (N_8274,N_8005,N_8170);
nor U8275 (N_8275,N_8059,N_8027);
xor U8276 (N_8276,N_8084,N_8120);
xor U8277 (N_8277,N_8193,N_8121);
or U8278 (N_8278,N_8125,N_8102);
nor U8279 (N_8279,N_8045,N_8148);
and U8280 (N_8280,N_8110,N_8057);
nor U8281 (N_8281,N_8147,N_8112);
or U8282 (N_8282,N_8127,N_8134);
nor U8283 (N_8283,N_8066,N_8176);
xor U8284 (N_8284,N_8038,N_8116);
nor U8285 (N_8285,N_8061,N_8109);
or U8286 (N_8286,N_8114,N_8075);
nor U8287 (N_8287,N_8150,N_8115);
nand U8288 (N_8288,N_8130,N_8135);
nor U8289 (N_8289,N_8053,N_8068);
nand U8290 (N_8290,N_8009,N_8097);
nor U8291 (N_8291,N_8108,N_8060);
xnor U8292 (N_8292,N_8180,N_8058);
or U8293 (N_8293,N_8051,N_8030);
nand U8294 (N_8294,N_8144,N_8082);
and U8295 (N_8295,N_8035,N_8172);
xor U8296 (N_8296,N_8092,N_8081);
or U8297 (N_8297,N_8177,N_8037);
xor U8298 (N_8298,N_8018,N_8165);
nand U8299 (N_8299,N_8133,N_8020);
nand U8300 (N_8300,N_8122,N_8094);
and U8301 (N_8301,N_8024,N_8018);
xnor U8302 (N_8302,N_8123,N_8124);
nor U8303 (N_8303,N_8098,N_8185);
xor U8304 (N_8304,N_8003,N_8115);
or U8305 (N_8305,N_8178,N_8122);
xnor U8306 (N_8306,N_8101,N_8131);
nand U8307 (N_8307,N_8040,N_8156);
xor U8308 (N_8308,N_8050,N_8017);
nand U8309 (N_8309,N_8083,N_8180);
nor U8310 (N_8310,N_8160,N_8173);
and U8311 (N_8311,N_8119,N_8174);
nor U8312 (N_8312,N_8198,N_8134);
nor U8313 (N_8313,N_8191,N_8146);
xor U8314 (N_8314,N_8003,N_8173);
and U8315 (N_8315,N_8033,N_8159);
nand U8316 (N_8316,N_8115,N_8093);
or U8317 (N_8317,N_8076,N_8080);
and U8318 (N_8318,N_8148,N_8083);
nor U8319 (N_8319,N_8167,N_8130);
and U8320 (N_8320,N_8140,N_8056);
nand U8321 (N_8321,N_8143,N_8129);
or U8322 (N_8322,N_8086,N_8185);
nand U8323 (N_8323,N_8109,N_8041);
nor U8324 (N_8324,N_8114,N_8088);
xnor U8325 (N_8325,N_8105,N_8041);
nand U8326 (N_8326,N_8031,N_8054);
and U8327 (N_8327,N_8029,N_8060);
xnor U8328 (N_8328,N_8183,N_8002);
or U8329 (N_8329,N_8016,N_8007);
nand U8330 (N_8330,N_8139,N_8135);
xnor U8331 (N_8331,N_8146,N_8086);
nor U8332 (N_8332,N_8061,N_8132);
nand U8333 (N_8333,N_8152,N_8131);
nor U8334 (N_8334,N_8088,N_8091);
xnor U8335 (N_8335,N_8029,N_8151);
or U8336 (N_8336,N_8164,N_8090);
and U8337 (N_8337,N_8077,N_8015);
and U8338 (N_8338,N_8020,N_8034);
xor U8339 (N_8339,N_8133,N_8083);
nor U8340 (N_8340,N_8106,N_8024);
or U8341 (N_8341,N_8066,N_8192);
and U8342 (N_8342,N_8192,N_8129);
or U8343 (N_8343,N_8102,N_8196);
or U8344 (N_8344,N_8076,N_8037);
nor U8345 (N_8345,N_8103,N_8092);
xor U8346 (N_8346,N_8012,N_8110);
or U8347 (N_8347,N_8059,N_8176);
or U8348 (N_8348,N_8054,N_8131);
and U8349 (N_8349,N_8035,N_8137);
xor U8350 (N_8350,N_8109,N_8055);
or U8351 (N_8351,N_8145,N_8046);
or U8352 (N_8352,N_8188,N_8170);
xor U8353 (N_8353,N_8036,N_8037);
nand U8354 (N_8354,N_8028,N_8037);
xor U8355 (N_8355,N_8161,N_8119);
and U8356 (N_8356,N_8059,N_8093);
xor U8357 (N_8357,N_8125,N_8004);
xor U8358 (N_8358,N_8053,N_8186);
or U8359 (N_8359,N_8190,N_8159);
nand U8360 (N_8360,N_8091,N_8154);
or U8361 (N_8361,N_8131,N_8060);
xor U8362 (N_8362,N_8130,N_8160);
or U8363 (N_8363,N_8190,N_8049);
xor U8364 (N_8364,N_8054,N_8058);
nor U8365 (N_8365,N_8028,N_8065);
and U8366 (N_8366,N_8182,N_8188);
nand U8367 (N_8367,N_8162,N_8033);
xnor U8368 (N_8368,N_8140,N_8103);
xor U8369 (N_8369,N_8034,N_8179);
or U8370 (N_8370,N_8026,N_8115);
and U8371 (N_8371,N_8018,N_8075);
and U8372 (N_8372,N_8144,N_8133);
nor U8373 (N_8373,N_8147,N_8002);
and U8374 (N_8374,N_8146,N_8132);
xnor U8375 (N_8375,N_8102,N_8128);
nor U8376 (N_8376,N_8161,N_8105);
or U8377 (N_8377,N_8124,N_8101);
xnor U8378 (N_8378,N_8151,N_8173);
nor U8379 (N_8379,N_8016,N_8136);
nand U8380 (N_8380,N_8155,N_8176);
xor U8381 (N_8381,N_8049,N_8158);
and U8382 (N_8382,N_8053,N_8134);
nand U8383 (N_8383,N_8086,N_8101);
xor U8384 (N_8384,N_8067,N_8021);
nor U8385 (N_8385,N_8059,N_8184);
or U8386 (N_8386,N_8127,N_8080);
or U8387 (N_8387,N_8140,N_8089);
and U8388 (N_8388,N_8080,N_8042);
or U8389 (N_8389,N_8083,N_8119);
nor U8390 (N_8390,N_8016,N_8088);
and U8391 (N_8391,N_8042,N_8000);
nor U8392 (N_8392,N_8089,N_8100);
nor U8393 (N_8393,N_8088,N_8077);
and U8394 (N_8394,N_8093,N_8038);
xor U8395 (N_8395,N_8121,N_8191);
nand U8396 (N_8396,N_8130,N_8028);
xnor U8397 (N_8397,N_8028,N_8120);
and U8398 (N_8398,N_8195,N_8188);
nand U8399 (N_8399,N_8096,N_8097);
nor U8400 (N_8400,N_8284,N_8265);
nand U8401 (N_8401,N_8289,N_8229);
or U8402 (N_8402,N_8232,N_8283);
xnor U8403 (N_8403,N_8331,N_8336);
xnor U8404 (N_8404,N_8372,N_8330);
nand U8405 (N_8405,N_8376,N_8340);
xnor U8406 (N_8406,N_8354,N_8290);
or U8407 (N_8407,N_8378,N_8225);
nand U8408 (N_8408,N_8363,N_8367);
and U8409 (N_8409,N_8361,N_8273);
nor U8410 (N_8410,N_8388,N_8242);
nor U8411 (N_8411,N_8302,N_8239);
and U8412 (N_8412,N_8356,N_8324);
nand U8413 (N_8413,N_8384,N_8275);
nor U8414 (N_8414,N_8262,N_8332);
nand U8415 (N_8415,N_8291,N_8227);
xnor U8416 (N_8416,N_8256,N_8261);
and U8417 (N_8417,N_8205,N_8292);
nor U8418 (N_8418,N_8301,N_8358);
or U8419 (N_8419,N_8266,N_8231);
xnor U8420 (N_8420,N_8311,N_8206);
or U8421 (N_8421,N_8385,N_8263);
xnor U8422 (N_8422,N_8369,N_8269);
xnor U8423 (N_8423,N_8396,N_8219);
or U8424 (N_8424,N_8217,N_8207);
xnor U8425 (N_8425,N_8334,N_8306);
nor U8426 (N_8426,N_8296,N_8240);
and U8427 (N_8427,N_8399,N_8276);
and U8428 (N_8428,N_8203,N_8391);
nor U8429 (N_8429,N_8286,N_8257);
xnor U8430 (N_8430,N_8395,N_8319);
xor U8431 (N_8431,N_8341,N_8373);
xnor U8432 (N_8432,N_8245,N_8345);
nor U8433 (N_8433,N_8236,N_8312);
nand U8434 (N_8434,N_8221,N_8270);
xor U8435 (N_8435,N_8244,N_8326);
and U8436 (N_8436,N_8338,N_8264);
nand U8437 (N_8437,N_8374,N_8359);
nor U8438 (N_8438,N_8309,N_8315);
nor U8439 (N_8439,N_8218,N_8299);
nand U8440 (N_8440,N_8387,N_8327);
xnor U8441 (N_8441,N_8249,N_8212);
and U8442 (N_8442,N_8343,N_8277);
and U8443 (N_8443,N_8235,N_8288);
and U8444 (N_8444,N_8254,N_8226);
and U8445 (N_8445,N_8382,N_8375);
nand U8446 (N_8446,N_8344,N_8352);
and U8447 (N_8447,N_8377,N_8200);
nor U8448 (N_8448,N_8279,N_8335);
nand U8449 (N_8449,N_8246,N_8348);
nand U8450 (N_8450,N_8365,N_8328);
or U8451 (N_8451,N_8379,N_8251);
nor U8452 (N_8452,N_8323,N_8223);
or U8453 (N_8453,N_8322,N_8281);
or U8454 (N_8454,N_8268,N_8271);
xor U8455 (N_8455,N_8282,N_8259);
nand U8456 (N_8456,N_8342,N_8287);
and U8457 (N_8457,N_8213,N_8305);
nand U8458 (N_8458,N_8278,N_8307);
nand U8459 (N_8459,N_8353,N_8211);
and U8460 (N_8460,N_8329,N_8320);
and U8461 (N_8461,N_8339,N_8222);
xor U8462 (N_8462,N_8383,N_8233);
and U8463 (N_8463,N_8390,N_8253);
xnor U8464 (N_8464,N_8314,N_8398);
and U8465 (N_8465,N_8337,N_8208);
nand U8466 (N_8466,N_8298,N_8201);
or U8467 (N_8467,N_8243,N_8394);
xor U8468 (N_8468,N_8370,N_8228);
or U8469 (N_8469,N_8308,N_8230);
and U8470 (N_8470,N_8333,N_8393);
xnor U8471 (N_8471,N_8220,N_8355);
xnor U8472 (N_8472,N_8380,N_8368);
or U8473 (N_8473,N_8247,N_8310);
nor U8474 (N_8474,N_8209,N_8317);
and U8475 (N_8475,N_8347,N_8272);
and U8476 (N_8476,N_8285,N_8294);
and U8477 (N_8477,N_8321,N_8397);
nand U8478 (N_8478,N_8295,N_8234);
nand U8479 (N_8479,N_8293,N_8357);
xnor U8480 (N_8480,N_8258,N_8366);
or U8481 (N_8481,N_8381,N_8304);
nand U8482 (N_8482,N_8215,N_8202);
and U8483 (N_8483,N_8260,N_8350);
xnor U8484 (N_8484,N_8250,N_8252);
nand U8485 (N_8485,N_8204,N_8237);
and U8486 (N_8486,N_8346,N_8362);
or U8487 (N_8487,N_8316,N_8297);
nand U8488 (N_8488,N_8224,N_8280);
nand U8489 (N_8489,N_8255,N_8364);
and U8490 (N_8490,N_8392,N_8371);
or U8491 (N_8491,N_8300,N_8216);
nand U8492 (N_8492,N_8325,N_8389);
xor U8493 (N_8493,N_8360,N_8274);
nand U8494 (N_8494,N_8386,N_8210);
or U8495 (N_8495,N_8238,N_8349);
xnor U8496 (N_8496,N_8241,N_8313);
xor U8497 (N_8497,N_8214,N_8248);
xnor U8498 (N_8498,N_8303,N_8318);
xnor U8499 (N_8499,N_8267,N_8351);
and U8500 (N_8500,N_8274,N_8319);
nor U8501 (N_8501,N_8355,N_8241);
nand U8502 (N_8502,N_8344,N_8345);
nand U8503 (N_8503,N_8283,N_8336);
nor U8504 (N_8504,N_8367,N_8284);
or U8505 (N_8505,N_8312,N_8348);
nor U8506 (N_8506,N_8308,N_8292);
and U8507 (N_8507,N_8339,N_8274);
or U8508 (N_8508,N_8205,N_8273);
nand U8509 (N_8509,N_8238,N_8372);
xor U8510 (N_8510,N_8334,N_8370);
and U8511 (N_8511,N_8225,N_8322);
nand U8512 (N_8512,N_8230,N_8251);
nand U8513 (N_8513,N_8244,N_8241);
xor U8514 (N_8514,N_8250,N_8379);
nor U8515 (N_8515,N_8249,N_8282);
nand U8516 (N_8516,N_8313,N_8286);
and U8517 (N_8517,N_8252,N_8247);
nor U8518 (N_8518,N_8302,N_8266);
and U8519 (N_8519,N_8220,N_8358);
xor U8520 (N_8520,N_8230,N_8368);
or U8521 (N_8521,N_8236,N_8310);
nor U8522 (N_8522,N_8390,N_8279);
and U8523 (N_8523,N_8217,N_8353);
xor U8524 (N_8524,N_8222,N_8206);
or U8525 (N_8525,N_8395,N_8309);
nand U8526 (N_8526,N_8312,N_8335);
xnor U8527 (N_8527,N_8214,N_8231);
and U8528 (N_8528,N_8223,N_8227);
nor U8529 (N_8529,N_8309,N_8217);
nor U8530 (N_8530,N_8359,N_8332);
or U8531 (N_8531,N_8363,N_8343);
xnor U8532 (N_8532,N_8277,N_8328);
nor U8533 (N_8533,N_8236,N_8263);
and U8534 (N_8534,N_8336,N_8338);
or U8535 (N_8535,N_8386,N_8219);
nor U8536 (N_8536,N_8378,N_8203);
or U8537 (N_8537,N_8294,N_8269);
or U8538 (N_8538,N_8203,N_8331);
nand U8539 (N_8539,N_8315,N_8249);
and U8540 (N_8540,N_8396,N_8209);
and U8541 (N_8541,N_8268,N_8299);
nand U8542 (N_8542,N_8328,N_8200);
or U8543 (N_8543,N_8270,N_8283);
xor U8544 (N_8544,N_8255,N_8289);
and U8545 (N_8545,N_8278,N_8255);
and U8546 (N_8546,N_8322,N_8329);
and U8547 (N_8547,N_8278,N_8377);
xnor U8548 (N_8548,N_8306,N_8323);
xnor U8549 (N_8549,N_8293,N_8292);
xor U8550 (N_8550,N_8202,N_8247);
or U8551 (N_8551,N_8250,N_8325);
or U8552 (N_8552,N_8214,N_8207);
nor U8553 (N_8553,N_8370,N_8231);
xor U8554 (N_8554,N_8261,N_8277);
nor U8555 (N_8555,N_8368,N_8324);
or U8556 (N_8556,N_8354,N_8225);
and U8557 (N_8557,N_8209,N_8371);
nor U8558 (N_8558,N_8206,N_8307);
or U8559 (N_8559,N_8307,N_8317);
nor U8560 (N_8560,N_8224,N_8349);
and U8561 (N_8561,N_8221,N_8352);
xnor U8562 (N_8562,N_8268,N_8327);
and U8563 (N_8563,N_8255,N_8335);
or U8564 (N_8564,N_8255,N_8258);
nor U8565 (N_8565,N_8377,N_8390);
or U8566 (N_8566,N_8211,N_8358);
nor U8567 (N_8567,N_8380,N_8266);
xor U8568 (N_8568,N_8313,N_8206);
nor U8569 (N_8569,N_8365,N_8295);
nor U8570 (N_8570,N_8250,N_8335);
and U8571 (N_8571,N_8383,N_8326);
or U8572 (N_8572,N_8215,N_8383);
xnor U8573 (N_8573,N_8363,N_8281);
nor U8574 (N_8574,N_8251,N_8219);
or U8575 (N_8575,N_8292,N_8204);
nand U8576 (N_8576,N_8254,N_8333);
nand U8577 (N_8577,N_8344,N_8308);
xnor U8578 (N_8578,N_8376,N_8215);
and U8579 (N_8579,N_8292,N_8355);
xnor U8580 (N_8580,N_8300,N_8346);
or U8581 (N_8581,N_8215,N_8314);
or U8582 (N_8582,N_8327,N_8323);
and U8583 (N_8583,N_8387,N_8323);
nand U8584 (N_8584,N_8269,N_8357);
nor U8585 (N_8585,N_8306,N_8246);
or U8586 (N_8586,N_8306,N_8304);
nand U8587 (N_8587,N_8283,N_8276);
nand U8588 (N_8588,N_8340,N_8375);
and U8589 (N_8589,N_8331,N_8393);
nor U8590 (N_8590,N_8292,N_8256);
nor U8591 (N_8591,N_8224,N_8389);
nand U8592 (N_8592,N_8267,N_8329);
and U8593 (N_8593,N_8278,N_8376);
nand U8594 (N_8594,N_8315,N_8327);
or U8595 (N_8595,N_8355,N_8320);
or U8596 (N_8596,N_8272,N_8353);
xor U8597 (N_8597,N_8306,N_8322);
nor U8598 (N_8598,N_8228,N_8216);
or U8599 (N_8599,N_8212,N_8382);
or U8600 (N_8600,N_8536,N_8485);
or U8601 (N_8601,N_8591,N_8466);
or U8602 (N_8602,N_8562,N_8581);
nor U8603 (N_8603,N_8507,N_8588);
nor U8604 (N_8604,N_8446,N_8432);
nor U8605 (N_8605,N_8472,N_8559);
nor U8606 (N_8606,N_8506,N_8564);
nor U8607 (N_8607,N_8508,N_8513);
and U8608 (N_8608,N_8554,N_8582);
xnor U8609 (N_8609,N_8463,N_8565);
or U8610 (N_8610,N_8442,N_8469);
nor U8611 (N_8611,N_8594,N_8545);
and U8612 (N_8612,N_8471,N_8455);
and U8613 (N_8613,N_8447,N_8589);
xor U8614 (N_8614,N_8460,N_8423);
nor U8615 (N_8615,N_8422,N_8538);
and U8616 (N_8616,N_8547,N_8498);
or U8617 (N_8617,N_8541,N_8491);
nor U8618 (N_8618,N_8456,N_8576);
nand U8619 (N_8619,N_8402,N_8476);
and U8620 (N_8620,N_8492,N_8549);
nand U8621 (N_8621,N_8431,N_8477);
nand U8622 (N_8622,N_8465,N_8521);
and U8623 (N_8623,N_8482,N_8544);
nor U8624 (N_8624,N_8522,N_8494);
or U8625 (N_8625,N_8468,N_8493);
nor U8626 (N_8626,N_8410,N_8577);
xnor U8627 (N_8627,N_8443,N_8599);
nand U8628 (N_8628,N_8424,N_8523);
nor U8629 (N_8629,N_8504,N_8478);
nand U8630 (N_8630,N_8555,N_8527);
xnor U8631 (N_8631,N_8407,N_8474);
and U8632 (N_8632,N_8433,N_8445);
nand U8633 (N_8633,N_8571,N_8440);
or U8634 (N_8634,N_8550,N_8490);
xnor U8635 (N_8635,N_8542,N_8454);
xor U8636 (N_8636,N_8537,N_8426);
or U8637 (N_8637,N_8596,N_8458);
or U8638 (N_8638,N_8451,N_8479);
and U8639 (N_8639,N_8430,N_8462);
nand U8640 (N_8640,N_8553,N_8401);
or U8641 (N_8641,N_8519,N_8517);
nor U8642 (N_8642,N_8501,N_8572);
xor U8643 (N_8643,N_8461,N_8529);
nor U8644 (N_8644,N_8467,N_8450);
nor U8645 (N_8645,N_8510,N_8487);
nor U8646 (N_8646,N_8453,N_8546);
or U8647 (N_8647,N_8409,N_8425);
or U8648 (N_8648,N_8563,N_8568);
or U8649 (N_8649,N_8595,N_8444);
nand U8650 (N_8650,N_8417,N_8558);
and U8651 (N_8651,N_8452,N_8509);
xnor U8652 (N_8652,N_8540,N_8497);
nand U8653 (N_8653,N_8459,N_8570);
xnor U8654 (N_8654,N_8464,N_8584);
or U8655 (N_8655,N_8526,N_8560);
xor U8656 (N_8656,N_8434,N_8480);
nand U8657 (N_8657,N_8449,N_8505);
and U8658 (N_8658,N_8548,N_8512);
nor U8659 (N_8659,N_8539,N_8475);
or U8660 (N_8660,N_8415,N_8436);
and U8661 (N_8661,N_8439,N_8535);
and U8662 (N_8662,N_8585,N_8590);
xnor U8663 (N_8663,N_8525,N_8533);
xnor U8664 (N_8664,N_8406,N_8551);
and U8665 (N_8665,N_8496,N_8421);
nor U8666 (N_8666,N_8473,N_8520);
nand U8667 (N_8667,N_8413,N_8567);
xor U8668 (N_8668,N_8502,N_8470);
nor U8669 (N_8669,N_8484,N_8578);
nor U8670 (N_8670,N_8514,N_8429);
xnor U8671 (N_8671,N_8499,N_8404);
xor U8672 (N_8672,N_8457,N_8597);
nand U8673 (N_8673,N_8552,N_8580);
nand U8674 (N_8674,N_8486,N_8441);
nand U8675 (N_8675,N_8575,N_8411);
nand U8676 (N_8676,N_8481,N_8403);
or U8677 (N_8677,N_8598,N_8518);
or U8678 (N_8678,N_8414,N_8524);
nand U8679 (N_8679,N_8556,N_8573);
xor U8680 (N_8680,N_8574,N_8516);
or U8681 (N_8681,N_8412,N_8561);
and U8682 (N_8682,N_8534,N_8435);
nand U8683 (N_8683,N_8528,N_8437);
or U8684 (N_8684,N_8587,N_8503);
xor U8685 (N_8685,N_8488,N_8483);
nor U8686 (N_8686,N_8408,N_8489);
xnor U8687 (N_8687,N_8448,N_8515);
nor U8688 (N_8688,N_8586,N_8416);
nand U8689 (N_8689,N_8592,N_8583);
nor U8690 (N_8690,N_8495,N_8419);
nand U8691 (N_8691,N_8420,N_8405);
nor U8692 (N_8692,N_8427,N_8418);
nor U8693 (N_8693,N_8428,N_8557);
or U8694 (N_8694,N_8566,N_8530);
nor U8695 (N_8695,N_8543,N_8569);
nor U8696 (N_8696,N_8511,N_8400);
and U8697 (N_8697,N_8593,N_8532);
nand U8698 (N_8698,N_8579,N_8438);
nand U8699 (N_8699,N_8531,N_8500);
and U8700 (N_8700,N_8463,N_8480);
nand U8701 (N_8701,N_8546,N_8505);
nand U8702 (N_8702,N_8471,N_8546);
or U8703 (N_8703,N_8493,N_8574);
nor U8704 (N_8704,N_8503,N_8541);
xnor U8705 (N_8705,N_8500,N_8444);
xnor U8706 (N_8706,N_8496,N_8448);
or U8707 (N_8707,N_8468,N_8585);
or U8708 (N_8708,N_8570,N_8421);
or U8709 (N_8709,N_8456,N_8497);
nor U8710 (N_8710,N_8406,N_8435);
or U8711 (N_8711,N_8460,N_8504);
and U8712 (N_8712,N_8500,N_8419);
nand U8713 (N_8713,N_8507,N_8406);
nor U8714 (N_8714,N_8443,N_8560);
xnor U8715 (N_8715,N_8597,N_8539);
or U8716 (N_8716,N_8435,N_8518);
and U8717 (N_8717,N_8493,N_8505);
or U8718 (N_8718,N_8486,N_8407);
and U8719 (N_8719,N_8464,N_8536);
and U8720 (N_8720,N_8480,N_8599);
xor U8721 (N_8721,N_8590,N_8503);
xor U8722 (N_8722,N_8426,N_8440);
or U8723 (N_8723,N_8463,N_8458);
nand U8724 (N_8724,N_8524,N_8495);
xnor U8725 (N_8725,N_8455,N_8557);
or U8726 (N_8726,N_8582,N_8455);
and U8727 (N_8727,N_8486,N_8550);
nor U8728 (N_8728,N_8562,N_8410);
xor U8729 (N_8729,N_8456,N_8527);
and U8730 (N_8730,N_8492,N_8503);
nor U8731 (N_8731,N_8447,N_8538);
and U8732 (N_8732,N_8582,N_8436);
xnor U8733 (N_8733,N_8423,N_8535);
nor U8734 (N_8734,N_8460,N_8418);
or U8735 (N_8735,N_8483,N_8512);
nand U8736 (N_8736,N_8550,N_8451);
and U8737 (N_8737,N_8569,N_8403);
or U8738 (N_8738,N_8561,N_8467);
nand U8739 (N_8739,N_8424,N_8576);
nor U8740 (N_8740,N_8563,N_8579);
and U8741 (N_8741,N_8449,N_8560);
or U8742 (N_8742,N_8509,N_8596);
nand U8743 (N_8743,N_8597,N_8403);
or U8744 (N_8744,N_8418,N_8564);
nand U8745 (N_8745,N_8538,N_8533);
nor U8746 (N_8746,N_8444,N_8416);
nor U8747 (N_8747,N_8436,N_8450);
nand U8748 (N_8748,N_8404,N_8591);
and U8749 (N_8749,N_8515,N_8446);
nand U8750 (N_8750,N_8464,N_8501);
and U8751 (N_8751,N_8440,N_8478);
and U8752 (N_8752,N_8475,N_8549);
xor U8753 (N_8753,N_8583,N_8472);
xnor U8754 (N_8754,N_8581,N_8455);
and U8755 (N_8755,N_8520,N_8407);
nand U8756 (N_8756,N_8417,N_8573);
nand U8757 (N_8757,N_8514,N_8426);
and U8758 (N_8758,N_8470,N_8488);
or U8759 (N_8759,N_8577,N_8573);
and U8760 (N_8760,N_8464,N_8579);
nand U8761 (N_8761,N_8504,N_8446);
xor U8762 (N_8762,N_8595,N_8598);
or U8763 (N_8763,N_8459,N_8568);
and U8764 (N_8764,N_8520,N_8546);
nand U8765 (N_8765,N_8453,N_8569);
and U8766 (N_8766,N_8588,N_8558);
or U8767 (N_8767,N_8501,N_8550);
nor U8768 (N_8768,N_8555,N_8433);
or U8769 (N_8769,N_8496,N_8430);
nand U8770 (N_8770,N_8412,N_8493);
nand U8771 (N_8771,N_8445,N_8545);
and U8772 (N_8772,N_8474,N_8497);
and U8773 (N_8773,N_8527,N_8498);
nand U8774 (N_8774,N_8494,N_8431);
nor U8775 (N_8775,N_8517,N_8547);
or U8776 (N_8776,N_8440,N_8492);
xnor U8777 (N_8777,N_8439,N_8528);
nor U8778 (N_8778,N_8448,N_8433);
xor U8779 (N_8779,N_8496,N_8460);
nor U8780 (N_8780,N_8448,N_8589);
nor U8781 (N_8781,N_8571,N_8420);
or U8782 (N_8782,N_8454,N_8500);
or U8783 (N_8783,N_8440,N_8443);
nand U8784 (N_8784,N_8488,N_8435);
xor U8785 (N_8785,N_8533,N_8445);
nand U8786 (N_8786,N_8502,N_8410);
nand U8787 (N_8787,N_8557,N_8587);
or U8788 (N_8788,N_8428,N_8509);
nand U8789 (N_8789,N_8521,N_8519);
nand U8790 (N_8790,N_8504,N_8450);
xnor U8791 (N_8791,N_8565,N_8522);
nand U8792 (N_8792,N_8440,N_8507);
xor U8793 (N_8793,N_8560,N_8509);
and U8794 (N_8794,N_8417,N_8501);
or U8795 (N_8795,N_8473,N_8578);
and U8796 (N_8796,N_8531,N_8591);
xor U8797 (N_8797,N_8420,N_8459);
nor U8798 (N_8798,N_8522,N_8537);
nand U8799 (N_8799,N_8575,N_8455);
or U8800 (N_8800,N_8744,N_8696);
nand U8801 (N_8801,N_8625,N_8761);
xor U8802 (N_8802,N_8776,N_8795);
nor U8803 (N_8803,N_8675,N_8605);
xor U8804 (N_8804,N_8689,N_8611);
and U8805 (N_8805,N_8666,N_8698);
xor U8806 (N_8806,N_8691,N_8711);
nor U8807 (N_8807,N_8630,N_8749);
or U8808 (N_8808,N_8649,N_8647);
and U8809 (N_8809,N_8615,N_8642);
nand U8810 (N_8810,N_8786,N_8633);
or U8811 (N_8811,N_8750,N_8646);
xnor U8812 (N_8812,N_8716,N_8687);
or U8813 (N_8813,N_8632,N_8620);
nor U8814 (N_8814,N_8703,N_8758);
or U8815 (N_8815,N_8670,N_8650);
nand U8816 (N_8816,N_8678,N_8715);
xnor U8817 (N_8817,N_8797,N_8606);
nand U8818 (N_8818,N_8737,N_8741);
nand U8819 (N_8819,N_8626,N_8773);
or U8820 (N_8820,N_8681,N_8644);
xor U8821 (N_8821,N_8731,N_8634);
nor U8822 (N_8822,N_8778,N_8693);
nand U8823 (N_8823,N_8709,N_8748);
and U8824 (N_8824,N_8683,N_8610);
nor U8825 (N_8825,N_8622,N_8706);
nor U8826 (N_8826,N_8617,N_8686);
xor U8827 (N_8827,N_8672,N_8657);
nand U8828 (N_8828,N_8674,N_8631);
or U8829 (N_8829,N_8743,N_8738);
or U8830 (N_8830,N_8679,N_8710);
xnor U8831 (N_8831,N_8727,N_8665);
or U8832 (N_8832,N_8600,N_8668);
and U8833 (N_8833,N_8636,N_8601);
xnor U8834 (N_8834,N_8729,N_8638);
nand U8835 (N_8835,N_8669,N_8671);
and U8836 (N_8836,N_8684,N_8713);
and U8837 (N_8837,N_8720,N_8781);
xnor U8838 (N_8838,N_8777,N_8762);
and U8839 (N_8839,N_8708,N_8690);
or U8840 (N_8840,N_8725,N_8624);
or U8841 (N_8841,N_8753,N_8712);
nand U8842 (N_8842,N_8787,N_8699);
nor U8843 (N_8843,N_8627,N_8798);
nor U8844 (N_8844,N_8635,N_8747);
and U8845 (N_8845,N_8697,N_8779);
nand U8846 (N_8846,N_8785,N_8742);
or U8847 (N_8847,N_8789,N_8759);
nand U8848 (N_8848,N_8602,N_8724);
or U8849 (N_8849,N_8756,N_8730);
nand U8850 (N_8850,N_8767,N_8770);
xnor U8851 (N_8851,N_8794,N_8769);
nand U8852 (N_8852,N_8662,N_8721);
nand U8853 (N_8853,N_8760,N_8658);
xnor U8854 (N_8854,N_8692,N_8718);
nor U8855 (N_8855,N_8780,N_8663);
nor U8856 (N_8856,N_8677,N_8673);
or U8857 (N_8857,N_8659,N_8700);
or U8858 (N_8858,N_8765,N_8655);
nand U8859 (N_8859,N_8603,N_8736);
xnor U8860 (N_8860,N_8734,N_8604);
nand U8861 (N_8861,N_8704,N_8764);
xnor U8862 (N_8862,N_8701,N_8754);
nand U8863 (N_8863,N_8637,N_8739);
nor U8864 (N_8864,N_8643,N_8719);
or U8865 (N_8865,N_8608,N_8714);
nand U8866 (N_8866,N_8616,N_8746);
or U8867 (N_8867,N_8768,N_8628);
and U8868 (N_8868,N_8735,N_8774);
or U8869 (N_8869,N_8792,N_8694);
nor U8870 (N_8870,N_8645,N_8619);
nor U8871 (N_8871,N_8685,N_8752);
xnor U8872 (N_8872,N_8717,N_8783);
and U8873 (N_8873,N_8707,N_8676);
xnor U8874 (N_8874,N_8784,N_8682);
and U8875 (N_8875,N_8656,N_8641);
nor U8876 (N_8876,N_8629,N_8660);
or U8877 (N_8877,N_8680,N_8618);
and U8878 (N_8878,N_8621,N_8702);
or U8879 (N_8879,N_8688,N_8791);
nand U8880 (N_8880,N_8723,N_8790);
nand U8881 (N_8881,N_8782,N_8733);
xor U8882 (N_8882,N_8654,N_8772);
nor U8883 (N_8883,N_8664,N_8651);
nor U8884 (N_8884,N_8607,N_8775);
or U8885 (N_8885,N_8640,N_8653);
nor U8886 (N_8886,N_8623,N_8757);
nor U8887 (N_8887,N_8751,N_8652);
or U8888 (N_8888,N_8661,N_8755);
nor U8889 (N_8889,N_8614,N_8612);
or U8890 (N_8890,N_8740,N_8609);
and U8891 (N_8891,N_8799,N_8788);
nand U8892 (N_8892,N_8763,N_8728);
or U8893 (N_8893,N_8648,N_8793);
or U8894 (N_8894,N_8705,N_8613);
nand U8895 (N_8895,N_8732,N_8722);
and U8896 (N_8896,N_8745,N_8766);
xor U8897 (N_8897,N_8726,N_8639);
and U8898 (N_8898,N_8771,N_8796);
or U8899 (N_8899,N_8667,N_8695);
nand U8900 (N_8900,N_8716,N_8754);
or U8901 (N_8901,N_8600,N_8689);
nand U8902 (N_8902,N_8697,N_8681);
nand U8903 (N_8903,N_8623,N_8641);
nor U8904 (N_8904,N_8651,N_8745);
xor U8905 (N_8905,N_8673,N_8624);
and U8906 (N_8906,N_8626,N_8659);
and U8907 (N_8907,N_8618,N_8786);
and U8908 (N_8908,N_8724,N_8603);
and U8909 (N_8909,N_8786,N_8780);
and U8910 (N_8910,N_8707,N_8622);
xor U8911 (N_8911,N_8798,N_8796);
xnor U8912 (N_8912,N_8737,N_8641);
xor U8913 (N_8913,N_8668,N_8769);
or U8914 (N_8914,N_8641,N_8742);
or U8915 (N_8915,N_8783,N_8662);
nor U8916 (N_8916,N_8615,N_8687);
or U8917 (N_8917,N_8660,N_8623);
nor U8918 (N_8918,N_8734,N_8707);
or U8919 (N_8919,N_8720,N_8753);
nor U8920 (N_8920,N_8667,N_8603);
nand U8921 (N_8921,N_8723,N_8768);
nor U8922 (N_8922,N_8787,N_8617);
xor U8923 (N_8923,N_8797,N_8651);
or U8924 (N_8924,N_8632,N_8628);
nand U8925 (N_8925,N_8681,N_8636);
or U8926 (N_8926,N_8669,N_8732);
and U8927 (N_8927,N_8704,N_8637);
or U8928 (N_8928,N_8759,N_8694);
and U8929 (N_8929,N_8702,N_8685);
and U8930 (N_8930,N_8644,N_8735);
and U8931 (N_8931,N_8601,N_8669);
or U8932 (N_8932,N_8682,N_8600);
nor U8933 (N_8933,N_8722,N_8738);
or U8934 (N_8934,N_8671,N_8771);
or U8935 (N_8935,N_8619,N_8689);
nand U8936 (N_8936,N_8767,N_8750);
xnor U8937 (N_8937,N_8786,N_8679);
xnor U8938 (N_8938,N_8760,N_8674);
and U8939 (N_8939,N_8661,N_8713);
xnor U8940 (N_8940,N_8641,N_8790);
nor U8941 (N_8941,N_8617,N_8786);
and U8942 (N_8942,N_8600,N_8656);
or U8943 (N_8943,N_8708,N_8683);
nor U8944 (N_8944,N_8652,N_8648);
nor U8945 (N_8945,N_8734,N_8735);
and U8946 (N_8946,N_8715,N_8780);
nand U8947 (N_8947,N_8748,N_8796);
and U8948 (N_8948,N_8690,N_8799);
or U8949 (N_8949,N_8750,N_8724);
nand U8950 (N_8950,N_8692,N_8708);
and U8951 (N_8951,N_8679,N_8724);
nand U8952 (N_8952,N_8794,N_8643);
and U8953 (N_8953,N_8622,N_8733);
xnor U8954 (N_8954,N_8640,N_8682);
or U8955 (N_8955,N_8734,N_8611);
and U8956 (N_8956,N_8731,N_8603);
nand U8957 (N_8957,N_8702,N_8731);
and U8958 (N_8958,N_8683,N_8778);
xnor U8959 (N_8959,N_8703,N_8634);
and U8960 (N_8960,N_8769,N_8627);
or U8961 (N_8961,N_8602,N_8680);
nor U8962 (N_8962,N_8679,N_8603);
xor U8963 (N_8963,N_8749,N_8653);
xnor U8964 (N_8964,N_8656,N_8670);
or U8965 (N_8965,N_8653,N_8726);
or U8966 (N_8966,N_8742,N_8765);
and U8967 (N_8967,N_8657,N_8648);
xor U8968 (N_8968,N_8636,N_8757);
nand U8969 (N_8969,N_8693,N_8620);
and U8970 (N_8970,N_8661,N_8796);
xor U8971 (N_8971,N_8689,N_8669);
nor U8972 (N_8972,N_8671,N_8622);
xor U8973 (N_8973,N_8693,N_8787);
or U8974 (N_8974,N_8786,N_8638);
nor U8975 (N_8975,N_8671,N_8732);
xnor U8976 (N_8976,N_8758,N_8618);
or U8977 (N_8977,N_8787,N_8605);
and U8978 (N_8978,N_8736,N_8795);
nand U8979 (N_8979,N_8646,N_8708);
nand U8980 (N_8980,N_8658,N_8656);
or U8981 (N_8981,N_8760,N_8751);
and U8982 (N_8982,N_8751,N_8735);
nor U8983 (N_8983,N_8683,N_8692);
xnor U8984 (N_8984,N_8671,N_8657);
xnor U8985 (N_8985,N_8617,N_8775);
and U8986 (N_8986,N_8755,N_8770);
and U8987 (N_8987,N_8617,N_8751);
and U8988 (N_8988,N_8755,N_8762);
and U8989 (N_8989,N_8798,N_8688);
nand U8990 (N_8990,N_8636,N_8796);
nand U8991 (N_8991,N_8692,N_8665);
or U8992 (N_8992,N_8653,N_8745);
or U8993 (N_8993,N_8699,N_8799);
nor U8994 (N_8994,N_8718,N_8703);
or U8995 (N_8995,N_8608,N_8758);
xor U8996 (N_8996,N_8671,N_8786);
or U8997 (N_8997,N_8662,N_8645);
or U8998 (N_8998,N_8694,N_8703);
xor U8999 (N_8999,N_8716,N_8777);
xor U9000 (N_9000,N_8828,N_8855);
or U9001 (N_9001,N_8933,N_8850);
xor U9002 (N_9002,N_8977,N_8927);
nor U9003 (N_9003,N_8836,N_8808);
xnor U9004 (N_9004,N_8817,N_8875);
nand U9005 (N_9005,N_8894,N_8822);
and U9006 (N_9006,N_8849,N_8955);
nor U9007 (N_9007,N_8802,N_8967);
nand U9008 (N_9008,N_8991,N_8961);
and U9009 (N_9009,N_8962,N_8803);
nor U9010 (N_9010,N_8976,N_8919);
nor U9011 (N_9011,N_8999,N_8966);
nor U9012 (N_9012,N_8869,N_8917);
and U9013 (N_9013,N_8852,N_8901);
xor U9014 (N_9014,N_8951,N_8932);
or U9015 (N_9015,N_8959,N_8982);
and U9016 (N_9016,N_8859,N_8916);
nand U9017 (N_9017,N_8837,N_8840);
nand U9018 (N_9018,N_8847,N_8903);
xor U9019 (N_9019,N_8863,N_8921);
nor U9020 (N_9020,N_8853,N_8807);
and U9021 (N_9021,N_8924,N_8805);
or U9022 (N_9022,N_8947,N_8856);
and U9023 (N_9023,N_8884,N_8820);
and U9024 (N_9024,N_8886,N_8978);
nand U9025 (N_9025,N_8812,N_8821);
and U9026 (N_9026,N_8825,N_8888);
xnor U9027 (N_9027,N_8938,N_8896);
nand U9028 (N_9028,N_8876,N_8922);
xor U9029 (N_9029,N_8920,N_8819);
and U9030 (N_9030,N_8858,N_8814);
and U9031 (N_9031,N_8890,N_8910);
or U9032 (N_9032,N_8969,N_8879);
or U9033 (N_9033,N_8842,N_8833);
xor U9034 (N_9034,N_8936,N_8897);
nor U9035 (N_9035,N_8801,N_8873);
xor U9036 (N_9036,N_8971,N_8867);
nand U9037 (N_9037,N_8827,N_8979);
or U9038 (N_9038,N_8800,N_8957);
and U9039 (N_9039,N_8815,N_8809);
or U9040 (N_9040,N_8887,N_8945);
and U9041 (N_9041,N_8874,N_8811);
or U9042 (N_9042,N_8974,N_8987);
nand U9043 (N_9043,N_8988,N_8895);
and U9044 (N_9044,N_8841,N_8900);
nand U9045 (N_9045,N_8871,N_8968);
and U9046 (N_9046,N_8806,N_8989);
nand U9047 (N_9047,N_8904,N_8816);
xor U9048 (N_9048,N_8829,N_8844);
nor U9049 (N_9049,N_8992,N_8878);
nand U9050 (N_9050,N_8960,N_8914);
xnor U9051 (N_9051,N_8983,N_8993);
nor U9052 (N_9052,N_8860,N_8926);
nand U9053 (N_9053,N_8835,N_8889);
nand U9054 (N_9054,N_8905,N_8866);
nand U9055 (N_9055,N_8834,N_8946);
and U9056 (N_9056,N_8832,N_8881);
xnor U9057 (N_9057,N_8891,N_8880);
xor U9058 (N_9058,N_8915,N_8824);
nor U9059 (N_9059,N_8804,N_8943);
nor U9060 (N_9060,N_8956,N_8865);
nand U9061 (N_9061,N_8870,N_8831);
and U9062 (N_9062,N_8911,N_8954);
nor U9063 (N_9063,N_8830,N_8985);
and U9064 (N_9064,N_8838,N_8975);
nor U9065 (N_9065,N_8918,N_8913);
nor U9066 (N_9066,N_8931,N_8963);
and U9067 (N_9067,N_8908,N_8925);
xnor U9068 (N_9068,N_8845,N_8818);
nor U9069 (N_9069,N_8883,N_8810);
nand U9070 (N_9070,N_8882,N_8912);
xor U9071 (N_9071,N_8851,N_8861);
xor U9072 (N_9072,N_8980,N_8964);
nor U9073 (N_9073,N_8848,N_8984);
or U9074 (N_9074,N_8990,N_8864);
xor U9075 (N_9075,N_8942,N_8941);
and U9076 (N_9076,N_8839,N_8872);
and U9077 (N_9077,N_8854,N_8935);
xor U9078 (N_9078,N_8902,N_8940);
nor U9079 (N_9079,N_8937,N_8868);
or U9080 (N_9080,N_8973,N_8929);
nor U9081 (N_9081,N_8892,N_8986);
or U9082 (N_9082,N_8965,N_8996);
or U9083 (N_9083,N_8948,N_8899);
xor U9084 (N_9084,N_8952,N_8862);
nand U9085 (N_9085,N_8998,N_8898);
nand U9086 (N_9086,N_8823,N_8906);
nand U9087 (N_9087,N_8939,N_8981);
nand U9088 (N_9088,N_8923,N_8934);
nand U9089 (N_9089,N_8893,N_8949);
or U9090 (N_9090,N_8970,N_8843);
nor U9091 (N_9091,N_8907,N_8953);
or U9092 (N_9092,N_8995,N_8846);
or U9093 (N_9093,N_8909,N_8928);
nor U9094 (N_9094,N_8950,N_8930);
nand U9095 (N_9095,N_8857,N_8994);
and U9096 (N_9096,N_8972,N_8813);
or U9097 (N_9097,N_8877,N_8826);
and U9098 (N_9098,N_8944,N_8997);
and U9099 (N_9099,N_8885,N_8958);
and U9100 (N_9100,N_8906,N_8927);
nor U9101 (N_9101,N_8806,N_8851);
xnor U9102 (N_9102,N_8986,N_8850);
nand U9103 (N_9103,N_8817,N_8922);
nor U9104 (N_9104,N_8915,N_8879);
nor U9105 (N_9105,N_8963,N_8853);
and U9106 (N_9106,N_8831,N_8959);
nand U9107 (N_9107,N_8927,N_8941);
nand U9108 (N_9108,N_8859,N_8809);
and U9109 (N_9109,N_8821,N_8903);
nor U9110 (N_9110,N_8867,N_8855);
xor U9111 (N_9111,N_8992,N_8993);
nor U9112 (N_9112,N_8835,N_8984);
and U9113 (N_9113,N_8885,N_8825);
xor U9114 (N_9114,N_8885,N_8818);
nand U9115 (N_9115,N_8834,N_8996);
nor U9116 (N_9116,N_8900,N_8899);
nor U9117 (N_9117,N_8880,N_8828);
nand U9118 (N_9118,N_8949,N_8879);
xor U9119 (N_9119,N_8819,N_8802);
or U9120 (N_9120,N_8839,N_8859);
nand U9121 (N_9121,N_8937,N_8902);
and U9122 (N_9122,N_8899,N_8920);
or U9123 (N_9123,N_8987,N_8894);
nand U9124 (N_9124,N_8928,N_8865);
and U9125 (N_9125,N_8819,N_8997);
nand U9126 (N_9126,N_8886,N_8928);
nor U9127 (N_9127,N_8897,N_8984);
or U9128 (N_9128,N_8854,N_8846);
nor U9129 (N_9129,N_8985,N_8915);
or U9130 (N_9130,N_8979,N_8848);
nor U9131 (N_9131,N_8917,N_8960);
xnor U9132 (N_9132,N_8890,N_8857);
nor U9133 (N_9133,N_8955,N_8967);
and U9134 (N_9134,N_8861,N_8846);
xnor U9135 (N_9135,N_8995,N_8860);
nand U9136 (N_9136,N_8962,N_8982);
and U9137 (N_9137,N_8988,N_8960);
xnor U9138 (N_9138,N_8848,N_8906);
or U9139 (N_9139,N_8817,N_8809);
and U9140 (N_9140,N_8864,N_8927);
nor U9141 (N_9141,N_8980,N_8863);
nand U9142 (N_9142,N_8997,N_8993);
or U9143 (N_9143,N_8979,N_8846);
nor U9144 (N_9144,N_8920,N_8914);
nand U9145 (N_9145,N_8956,N_8998);
and U9146 (N_9146,N_8803,N_8976);
xnor U9147 (N_9147,N_8988,N_8949);
nor U9148 (N_9148,N_8967,N_8940);
and U9149 (N_9149,N_8850,N_8895);
nor U9150 (N_9150,N_8997,N_8878);
xnor U9151 (N_9151,N_8969,N_8931);
nand U9152 (N_9152,N_8888,N_8940);
nand U9153 (N_9153,N_8838,N_8841);
xor U9154 (N_9154,N_8975,N_8996);
xor U9155 (N_9155,N_8930,N_8841);
xnor U9156 (N_9156,N_8861,N_8911);
and U9157 (N_9157,N_8953,N_8971);
or U9158 (N_9158,N_8886,N_8883);
or U9159 (N_9159,N_8940,N_8984);
nor U9160 (N_9160,N_8810,N_8982);
and U9161 (N_9161,N_8851,N_8899);
nand U9162 (N_9162,N_8955,N_8839);
and U9163 (N_9163,N_8988,N_8897);
nor U9164 (N_9164,N_8935,N_8927);
nand U9165 (N_9165,N_8993,N_8904);
or U9166 (N_9166,N_8979,N_8906);
nor U9167 (N_9167,N_8815,N_8966);
nand U9168 (N_9168,N_8829,N_8880);
or U9169 (N_9169,N_8931,N_8844);
and U9170 (N_9170,N_8904,N_8925);
nand U9171 (N_9171,N_8809,N_8876);
xor U9172 (N_9172,N_8909,N_8985);
nand U9173 (N_9173,N_8969,N_8808);
xor U9174 (N_9174,N_8876,N_8834);
nor U9175 (N_9175,N_8893,N_8908);
xor U9176 (N_9176,N_8942,N_8996);
nand U9177 (N_9177,N_8985,N_8811);
xor U9178 (N_9178,N_8903,N_8914);
xnor U9179 (N_9179,N_8921,N_8967);
nand U9180 (N_9180,N_8919,N_8995);
or U9181 (N_9181,N_8807,N_8992);
and U9182 (N_9182,N_8836,N_8868);
nand U9183 (N_9183,N_8887,N_8802);
and U9184 (N_9184,N_8949,N_8978);
or U9185 (N_9185,N_8950,N_8850);
and U9186 (N_9186,N_8934,N_8872);
and U9187 (N_9187,N_8966,N_8898);
nand U9188 (N_9188,N_8817,N_8851);
nand U9189 (N_9189,N_8879,N_8840);
nand U9190 (N_9190,N_8885,N_8875);
nor U9191 (N_9191,N_8963,N_8924);
or U9192 (N_9192,N_8991,N_8988);
xnor U9193 (N_9193,N_8910,N_8987);
or U9194 (N_9194,N_8829,N_8920);
or U9195 (N_9195,N_8991,N_8892);
nand U9196 (N_9196,N_8925,N_8863);
and U9197 (N_9197,N_8888,N_8812);
or U9198 (N_9198,N_8937,N_8896);
or U9199 (N_9199,N_8970,N_8927);
xor U9200 (N_9200,N_9168,N_9187);
and U9201 (N_9201,N_9128,N_9073);
xnor U9202 (N_9202,N_9133,N_9102);
nand U9203 (N_9203,N_9194,N_9126);
nor U9204 (N_9204,N_9107,N_9189);
xnor U9205 (N_9205,N_9183,N_9105);
xnor U9206 (N_9206,N_9069,N_9104);
nand U9207 (N_9207,N_9060,N_9023);
xnor U9208 (N_9208,N_9031,N_9117);
nor U9209 (N_9209,N_9096,N_9108);
and U9210 (N_9210,N_9182,N_9174);
xor U9211 (N_9211,N_9160,N_9161);
or U9212 (N_9212,N_9064,N_9081);
nor U9213 (N_9213,N_9180,N_9147);
nand U9214 (N_9214,N_9097,N_9058);
nor U9215 (N_9215,N_9028,N_9088);
or U9216 (N_9216,N_9125,N_9151);
xor U9217 (N_9217,N_9042,N_9170);
nand U9218 (N_9218,N_9080,N_9066);
nor U9219 (N_9219,N_9008,N_9148);
nand U9220 (N_9220,N_9124,N_9186);
nor U9221 (N_9221,N_9195,N_9113);
or U9222 (N_9222,N_9038,N_9007);
xor U9223 (N_9223,N_9114,N_9067);
xor U9224 (N_9224,N_9002,N_9109);
nand U9225 (N_9225,N_9049,N_9163);
xnor U9226 (N_9226,N_9142,N_9188);
nor U9227 (N_9227,N_9062,N_9127);
or U9228 (N_9228,N_9177,N_9011);
nand U9229 (N_9229,N_9025,N_9162);
nand U9230 (N_9230,N_9044,N_9120);
and U9231 (N_9231,N_9087,N_9098);
and U9232 (N_9232,N_9015,N_9006);
xnor U9233 (N_9233,N_9090,N_9199);
nand U9234 (N_9234,N_9101,N_9022);
or U9235 (N_9235,N_9196,N_9138);
and U9236 (N_9236,N_9178,N_9035);
xnor U9237 (N_9237,N_9130,N_9020);
and U9238 (N_9238,N_9070,N_9018);
nand U9239 (N_9239,N_9164,N_9167);
and U9240 (N_9240,N_9034,N_9071);
xnor U9241 (N_9241,N_9179,N_9121);
and U9242 (N_9242,N_9143,N_9092);
or U9243 (N_9243,N_9003,N_9047);
nand U9244 (N_9244,N_9145,N_9085);
xnor U9245 (N_9245,N_9116,N_9019);
nand U9246 (N_9246,N_9041,N_9154);
nor U9247 (N_9247,N_9061,N_9155);
xnor U9248 (N_9248,N_9026,N_9144);
nor U9249 (N_9249,N_9048,N_9135);
nand U9250 (N_9250,N_9001,N_9198);
and U9251 (N_9251,N_9118,N_9051);
nor U9252 (N_9252,N_9173,N_9110);
nand U9253 (N_9253,N_9190,N_9095);
xnor U9254 (N_9254,N_9165,N_9140);
nand U9255 (N_9255,N_9193,N_9156);
xnor U9256 (N_9256,N_9146,N_9065);
nor U9257 (N_9257,N_9119,N_9059);
or U9258 (N_9258,N_9129,N_9057);
or U9259 (N_9259,N_9150,N_9084);
or U9260 (N_9260,N_9106,N_9141);
nand U9261 (N_9261,N_9152,N_9139);
or U9262 (N_9262,N_9158,N_9037);
xor U9263 (N_9263,N_9030,N_9175);
xnor U9264 (N_9264,N_9082,N_9004);
or U9265 (N_9265,N_9149,N_9075);
nor U9266 (N_9266,N_9115,N_9040);
xor U9267 (N_9267,N_9172,N_9086);
or U9268 (N_9268,N_9103,N_9014);
xor U9269 (N_9269,N_9094,N_9181);
nand U9270 (N_9270,N_9024,N_9132);
or U9271 (N_9271,N_9077,N_9013);
xor U9272 (N_9272,N_9089,N_9054);
or U9273 (N_9273,N_9111,N_9033);
and U9274 (N_9274,N_9052,N_9184);
xor U9275 (N_9275,N_9032,N_9046);
nand U9276 (N_9276,N_9039,N_9159);
and U9277 (N_9277,N_9122,N_9136);
xnor U9278 (N_9278,N_9123,N_9072);
or U9279 (N_9279,N_9171,N_9076);
nor U9280 (N_9280,N_9063,N_9005);
nand U9281 (N_9281,N_9191,N_9137);
nand U9282 (N_9282,N_9027,N_9043);
and U9283 (N_9283,N_9021,N_9029);
or U9284 (N_9284,N_9166,N_9078);
xor U9285 (N_9285,N_9053,N_9079);
xor U9286 (N_9286,N_9045,N_9000);
and U9287 (N_9287,N_9192,N_9012);
or U9288 (N_9288,N_9050,N_9185);
and U9289 (N_9289,N_9099,N_9010);
and U9290 (N_9290,N_9153,N_9197);
nor U9291 (N_9291,N_9017,N_9068);
or U9292 (N_9292,N_9131,N_9093);
nand U9293 (N_9293,N_9112,N_9055);
xnor U9294 (N_9294,N_9074,N_9016);
and U9295 (N_9295,N_9036,N_9009);
xor U9296 (N_9296,N_9176,N_9169);
xnor U9297 (N_9297,N_9091,N_9083);
or U9298 (N_9298,N_9134,N_9100);
nor U9299 (N_9299,N_9157,N_9056);
or U9300 (N_9300,N_9031,N_9030);
nand U9301 (N_9301,N_9177,N_9195);
xor U9302 (N_9302,N_9150,N_9180);
nor U9303 (N_9303,N_9137,N_9141);
and U9304 (N_9304,N_9157,N_9152);
or U9305 (N_9305,N_9001,N_9009);
xor U9306 (N_9306,N_9072,N_9157);
xnor U9307 (N_9307,N_9179,N_9126);
and U9308 (N_9308,N_9011,N_9184);
nor U9309 (N_9309,N_9121,N_9143);
xor U9310 (N_9310,N_9120,N_9115);
or U9311 (N_9311,N_9009,N_9171);
xor U9312 (N_9312,N_9134,N_9042);
xor U9313 (N_9313,N_9058,N_9072);
xor U9314 (N_9314,N_9057,N_9124);
nand U9315 (N_9315,N_9153,N_9041);
or U9316 (N_9316,N_9130,N_9102);
and U9317 (N_9317,N_9055,N_9177);
or U9318 (N_9318,N_9040,N_9023);
or U9319 (N_9319,N_9048,N_9197);
or U9320 (N_9320,N_9137,N_9192);
and U9321 (N_9321,N_9049,N_9145);
and U9322 (N_9322,N_9025,N_9081);
nand U9323 (N_9323,N_9105,N_9149);
and U9324 (N_9324,N_9002,N_9008);
nand U9325 (N_9325,N_9093,N_9160);
and U9326 (N_9326,N_9156,N_9052);
and U9327 (N_9327,N_9123,N_9097);
xor U9328 (N_9328,N_9007,N_9188);
xor U9329 (N_9329,N_9150,N_9093);
nor U9330 (N_9330,N_9115,N_9036);
or U9331 (N_9331,N_9094,N_9147);
xor U9332 (N_9332,N_9142,N_9028);
xnor U9333 (N_9333,N_9178,N_9058);
and U9334 (N_9334,N_9163,N_9199);
nor U9335 (N_9335,N_9160,N_9164);
and U9336 (N_9336,N_9071,N_9177);
or U9337 (N_9337,N_9199,N_9026);
xor U9338 (N_9338,N_9163,N_9039);
xnor U9339 (N_9339,N_9114,N_9075);
nand U9340 (N_9340,N_9084,N_9198);
nor U9341 (N_9341,N_9167,N_9031);
nand U9342 (N_9342,N_9120,N_9180);
nor U9343 (N_9343,N_9154,N_9097);
or U9344 (N_9344,N_9111,N_9120);
or U9345 (N_9345,N_9172,N_9141);
nand U9346 (N_9346,N_9190,N_9141);
xor U9347 (N_9347,N_9087,N_9145);
and U9348 (N_9348,N_9151,N_9111);
and U9349 (N_9349,N_9135,N_9195);
xnor U9350 (N_9350,N_9198,N_9073);
nand U9351 (N_9351,N_9042,N_9004);
nand U9352 (N_9352,N_9122,N_9047);
and U9353 (N_9353,N_9074,N_9012);
and U9354 (N_9354,N_9197,N_9113);
nand U9355 (N_9355,N_9082,N_9038);
xor U9356 (N_9356,N_9041,N_9132);
xnor U9357 (N_9357,N_9010,N_9186);
and U9358 (N_9358,N_9048,N_9189);
or U9359 (N_9359,N_9157,N_9113);
nor U9360 (N_9360,N_9073,N_9036);
or U9361 (N_9361,N_9135,N_9086);
nor U9362 (N_9362,N_9140,N_9099);
nor U9363 (N_9363,N_9042,N_9078);
and U9364 (N_9364,N_9169,N_9115);
nor U9365 (N_9365,N_9005,N_9127);
and U9366 (N_9366,N_9005,N_9115);
nand U9367 (N_9367,N_9016,N_9164);
xnor U9368 (N_9368,N_9043,N_9006);
nor U9369 (N_9369,N_9066,N_9130);
nand U9370 (N_9370,N_9036,N_9143);
and U9371 (N_9371,N_9161,N_9067);
xnor U9372 (N_9372,N_9034,N_9020);
or U9373 (N_9373,N_9052,N_9113);
and U9374 (N_9374,N_9180,N_9124);
xnor U9375 (N_9375,N_9043,N_9080);
and U9376 (N_9376,N_9199,N_9007);
and U9377 (N_9377,N_9143,N_9011);
and U9378 (N_9378,N_9178,N_9118);
nor U9379 (N_9379,N_9180,N_9176);
nor U9380 (N_9380,N_9043,N_9010);
nor U9381 (N_9381,N_9034,N_9053);
and U9382 (N_9382,N_9069,N_9009);
or U9383 (N_9383,N_9032,N_9043);
and U9384 (N_9384,N_9155,N_9079);
nand U9385 (N_9385,N_9029,N_9133);
nor U9386 (N_9386,N_9056,N_9156);
nand U9387 (N_9387,N_9120,N_9073);
nor U9388 (N_9388,N_9018,N_9151);
and U9389 (N_9389,N_9108,N_9077);
xnor U9390 (N_9390,N_9126,N_9036);
nand U9391 (N_9391,N_9178,N_9008);
and U9392 (N_9392,N_9140,N_9003);
nand U9393 (N_9393,N_9158,N_9011);
and U9394 (N_9394,N_9142,N_9064);
or U9395 (N_9395,N_9100,N_9178);
xnor U9396 (N_9396,N_9158,N_9104);
nor U9397 (N_9397,N_9009,N_9093);
or U9398 (N_9398,N_9047,N_9192);
or U9399 (N_9399,N_9110,N_9049);
and U9400 (N_9400,N_9316,N_9327);
nor U9401 (N_9401,N_9380,N_9294);
and U9402 (N_9402,N_9278,N_9246);
nor U9403 (N_9403,N_9296,N_9350);
nor U9404 (N_9404,N_9284,N_9309);
nor U9405 (N_9405,N_9210,N_9207);
xor U9406 (N_9406,N_9337,N_9388);
xor U9407 (N_9407,N_9370,N_9311);
xnor U9408 (N_9408,N_9382,N_9303);
or U9409 (N_9409,N_9218,N_9213);
nand U9410 (N_9410,N_9354,N_9360);
nand U9411 (N_9411,N_9236,N_9399);
xor U9412 (N_9412,N_9286,N_9390);
xor U9413 (N_9413,N_9392,N_9243);
nor U9414 (N_9414,N_9355,N_9203);
nand U9415 (N_9415,N_9344,N_9290);
or U9416 (N_9416,N_9206,N_9221);
xnor U9417 (N_9417,N_9330,N_9228);
or U9418 (N_9418,N_9306,N_9367);
or U9419 (N_9419,N_9345,N_9312);
and U9420 (N_9420,N_9342,N_9340);
or U9421 (N_9421,N_9348,N_9300);
nor U9422 (N_9422,N_9292,N_9394);
and U9423 (N_9423,N_9200,N_9255);
xnor U9424 (N_9424,N_9211,N_9365);
or U9425 (N_9425,N_9209,N_9372);
and U9426 (N_9426,N_9289,N_9371);
nand U9427 (N_9427,N_9377,N_9277);
and U9428 (N_9428,N_9285,N_9224);
xnor U9429 (N_9429,N_9352,N_9253);
or U9430 (N_9430,N_9265,N_9346);
and U9431 (N_9431,N_9279,N_9287);
nor U9432 (N_9432,N_9230,N_9222);
and U9433 (N_9433,N_9334,N_9232);
or U9434 (N_9434,N_9214,N_9322);
nor U9435 (N_9435,N_9263,N_9387);
nand U9436 (N_9436,N_9288,N_9304);
and U9437 (N_9437,N_9329,N_9216);
and U9438 (N_9438,N_9381,N_9358);
xnor U9439 (N_9439,N_9204,N_9299);
nand U9440 (N_9440,N_9269,N_9326);
nand U9441 (N_9441,N_9368,N_9267);
nor U9442 (N_9442,N_9349,N_9212);
nor U9443 (N_9443,N_9217,N_9275);
and U9444 (N_9444,N_9320,N_9356);
nand U9445 (N_9445,N_9220,N_9283);
xor U9446 (N_9446,N_9362,N_9266);
or U9447 (N_9447,N_9389,N_9302);
nor U9448 (N_9448,N_9341,N_9258);
and U9449 (N_9449,N_9386,N_9351);
xnor U9450 (N_9450,N_9391,N_9225);
nor U9451 (N_9451,N_9291,N_9229);
xnor U9452 (N_9452,N_9215,N_9332);
nor U9453 (N_9453,N_9314,N_9256);
xnor U9454 (N_9454,N_9357,N_9364);
or U9455 (N_9455,N_9301,N_9202);
and U9456 (N_9456,N_9262,N_9318);
nor U9457 (N_9457,N_9251,N_9393);
nor U9458 (N_9458,N_9325,N_9383);
and U9459 (N_9459,N_9223,N_9295);
nand U9460 (N_9460,N_9384,N_9369);
nor U9461 (N_9461,N_9310,N_9321);
and U9462 (N_9462,N_9235,N_9379);
and U9463 (N_9463,N_9239,N_9260);
and U9464 (N_9464,N_9244,N_9282);
xnor U9465 (N_9465,N_9201,N_9385);
and U9466 (N_9466,N_9378,N_9343);
xnor U9467 (N_9467,N_9363,N_9315);
nand U9468 (N_9468,N_9397,N_9293);
or U9469 (N_9469,N_9333,N_9234);
and U9470 (N_9470,N_9247,N_9298);
nand U9471 (N_9471,N_9323,N_9338);
nor U9472 (N_9472,N_9297,N_9317);
and U9473 (N_9473,N_9280,N_9264);
xor U9474 (N_9474,N_9281,N_9273);
nor U9475 (N_9475,N_9359,N_9259);
or U9476 (N_9476,N_9336,N_9366);
and U9477 (N_9477,N_9328,N_9257);
nand U9478 (N_9478,N_9254,N_9252);
nand U9479 (N_9479,N_9231,N_9249);
nand U9480 (N_9480,N_9233,N_9353);
xor U9481 (N_9481,N_9347,N_9271);
nand U9482 (N_9482,N_9208,N_9374);
xnor U9483 (N_9483,N_9361,N_9324);
or U9484 (N_9484,N_9227,N_9270);
or U9485 (N_9485,N_9331,N_9339);
xor U9486 (N_9486,N_9242,N_9319);
and U9487 (N_9487,N_9272,N_9226);
and U9488 (N_9488,N_9237,N_9240);
and U9489 (N_9489,N_9250,N_9276);
or U9490 (N_9490,N_9308,N_9375);
xor U9491 (N_9491,N_9335,N_9268);
xor U9492 (N_9492,N_9274,N_9398);
or U9493 (N_9493,N_9307,N_9245);
and U9494 (N_9494,N_9205,N_9396);
nand U9495 (N_9495,N_9241,N_9248);
or U9496 (N_9496,N_9376,N_9313);
xnor U9497 (N_9497,N_9373,N_9261);
nor U9498 (N_9498,N_9395,N_9238);
or U9499 (N_9499,N_9219,N_9305);
or U9500 (N_9500,N_9209,N_9249);
xnor U9501 (N_9501,N_9297,N_9337);
or U9502 (N_9502,N_9262,N_9250);
and U9503 (N_9503,N_9255,N_9267);
or U9504 (N_9504,N_9244,N_9319);
nand U9505 (N_9505,N_9390,N_9244);
or U9506 (N_9506,N_9230,N_9281);
xor U9507 (N_9507,N_9323,N_9268);
nand U9508 (N_9508,N_9363,N_9343);
or U9509 (N_9509,N_9354,N_9273);
nor U9510 (N_9510,N_9383,N_9284);
or U9511 (N_9511,N_9349,N_9247);
or U9512 (N_9512,N_9259,N_9260);
and U9513 (N_9513,N_9311,N_9347);
nand U9514 (N_9514,N_9331,N_9209);
and U9515 (N_9515,N_9303,N_9315);
or U9516 (N_9516,N_9230,N_9232);
xor U9517 (N_9517,N_9273,N_9233);
nor U9518 (N_9518,N_9382,N_9210);
nand U9519 (N_9519,N_9204,N_9266);
nand U9520 (N_9520,N_9394,N_9368);
and U9521 (N_9521,N_9315,N_9397);
and U9522 (N_9522,N_9245,N_9324);
or U9523 (N_9523,N_9248,N_9251);
nor U9524 (N_9524,N_9373,N_9384);
nor U9525 (N_9525,N_9390,N_9214);
or U9526 (N_9526,N_9244,N_9300);
xor U9527 (N_9527,N_9350,N_9326);
and U9528 (N_9528,N_9206,N_9307);
xor U9529 (N_9529,N_9227,N_9250);
nor U9530 (N_9530,N_9383,N_9267);
xor U9531 (N_9531,N_9322,N_9330);
or U9532 (N_9532,N_9364,N_9303);
nand U9533 (N_9533,N_9286,N_9248);
or U9534 (N_9534,N_9242,N_9206);
and U9535 (N_9535,N_9274,N_9280);
xor U9536 (N_9536,N_9355,N_9398);
or U9537 (N_9537,N_9359,N_9381);
or U9538 (N_9538,N_9302,N_9258);
nor U9539 (N_9539,N_9224,N_9302);
nor U9540 (N_9540,N_9372,N_9303);
nand U9541 (N_9541,N_9238,N_9284);
xnor U9542 (N_9542,N_9361,N_9259);
and U9543 (N_9543,N_9265,N_9316);
xor U9544 (N_9544,N_9379,N_9278);
nand U9545 (N_9545,N_9227,N_9324);
or U9546 (N_9546,N_9250,N_9207);
xnor U9547 (N_9547,N_9389,N_9253);
and U9548 (N_9548,N_9336,N_9359);
nand U9549 (N_9549,N_9216,N_9246);
nor U9550 (N_9550,N_9247,N_9345);
xor U9551 (N_9551,N_9260,N_9312);
xor U9552 (N_9552,N_9348,N_9396);
or U9553 (N_9553,N_9297,N_9334);
xor U9554 (N_9554,N_9262,N_9396);
nand U9555 (N_9555,N_9335,N_9208);
and U9556 (N_9556,N_9233,N_9209);
nor U9557 (N_9557,N_9361,N_9391);
nand U9558 (N_9558,N_9351,N_9368);
and U9559 (N_9559,N_9309,N_9236);
nor U9560 (N_9560,N_9346,N_9201);
or U9561 (N_9561,N_9303,N_9306);
and U9562 (N_9562,N_9317,N_9237);
or U9563 (N_9563,N_9398,N_9334);
nand U9564 (N_9564,N_9373,N_9236);
xor U9565 (N_9565,N_9373,N_9370);
nor U9566 (N_9566,N_9239,N_9266);
nand U9567 (N_9567,N_9382,N_9290);
or U9568 (N_9568,N_9211,N_9260);
nor U9569 (N_9569,N_9272,N_9218);
nor U9570 (N_9570,N_9298,N_9309);
xnor U9571 (N_9571,N_9356,N_9298);
nand U9572 (N_9572,N_9211,N_9200);
xor U9573 (N_9573,N_9269,N_9255);
and U9574 (N_9574,N_9316,N_9213);
xor U9575 (N_9575,N_9227,N_9234);
nor U9576 (N_9576,N_9365,N_9246);
and U9577 (N_9577,N_9310,N_9226);
and U9578 (N_9578,N_9256,N_9378);
nand U9579 (N_9579,N_9294,N_9275);
and U9580 (N_9580,N_9291,N_9307);
xor U9581 (N_9581,N_9365,N_9393);
nor U9582 (N_9582,N_9246,N_9219);
or U9583 (N_9583,N_9326,N_9368);
nand U9584 (N_9584,N_9329,N_9235);
nor U9585 (N_9585,N_9257,N_9352);
and U9586 (N_9586,N_9214,N_9315);
xor U9587 (N_9587,N_9236,N_9288);
nand U9588 (N_9588,N_9203,N_9359);
and U9589 (N_9589,N_9307,N_9371);
nor U9590 (N_9590,N_9268,N_9242);
nor U9591 (N_9591,N_9237,N_9315);
or U9592 (N_9592,N_9250,N_9366);
and U9593 (N_9593,N_9336,N_9223);
and U9594 (N_9594,N_9311,N_9385);
nor U9595 (N_9595,N_9241,N_9222);
or U9596 (N_9596,N_9290,N_9232);
nand U9597 (N_9597,N_9273,N_9249);
and U9598 (N_9598,N_9346,N_9220);
and U9599 (N_9599,N_9342,N_9219);
and U9600 (N_9600,N_9513,N_9461);
and U9601 (N_9601,N_9418,N_9584);
nor U9602 (N_9602,N_9597,N_9453);
xor U9603 (N_9603,N_9467,N_9507);
nand U9604 (N_9604,N_9493,N_9408);
xnor U9605 (N_9605,N_9494,N_9447);
or U9606 (N_9606,N_9577,N_9471);
xnor U9607 (N_9607,N_9451,N_9519);
nand U9608 (N_9608,N_9481,N_9582);
or U9609 (N_9609,N_9557,N_9559);
and U9610 (N_9610,N_9535,N_9544);
xor U9611 (N_9611,N_9543,N_9539);
xor U9612 (N_9612,N_9427,N_9587);
xnor U9613 (N_9613,N_9522,N_9483);
or U9614 (N_9614,N_9527,N_9537);
xor U9615 (N_9615,N_9458,N_9508);
nand U9616 (N_9616,N_9448,N_9541);
nand U9617 (N_9617,N_9407,N_9533);
and U9618 (N_9618,N_9431,N_9436);
nor U9619 (N_9619,N_9433,N_9429);
nand U9620 (N_9620,N_9492,N_9503);
xor U9621 (N_9621,N_9498,N_9567);
xor U9622 (N_9622,N_9509,N_9596);
xnor U9623 (N_9623,N_9488,N_9469);
nor U9624 (N_9624,N_9401,N_9554);
nor U9625 (N_9625,N_9578,N_9406);
nand U9626 (N_9626,N_9443,N_9504);
or U9627 (N_9627,N_9588,N_9564);
xnor U9628 (N_9628,N_9430,N_9415);
nand U9629 (N_9629,N_9590,N_9550);
xor U9630 (N_9630,N_9529,N_9473);
xor U9631 (N_9631,N_9548,N_9512);
xor U9632 (N_9632,N_9437,N_9482);
or U9633 (N_9633,N_9593,N_9547);
and U9634 (N_9634,N_9403,N_9570);
nor U9635 (N_9635,N_9560,N_9466);
nor U9636 (N_9636,N_9419,N_9514);
nand U9637 (N_9637,N_9475,N_9417);
nand U9638 (N_9638,N_9532,N_9538);
nand U9639 (N_9639,N_9555,N_9495);
nand U9640 (N_9640,N_9574,N_9591);
xnor U9641 (N_9641,N_9424,N_9456);
xnor U9642 (N_9642,N_9580,N_9553);
nor U9643 (N_9643,N_9439,N_9490);
nand U9644 (N_9644,N_9594,N_9520);
nand U9645 (N_9645,N_9511,N_9523);
nor U9646 (N_9646,N_9500,N_9434);
nor U9647 (N_9647,N_9413,N_9402);
xnor U9648 (N_9648,N_9455,N_9472);
nand U9649 (N_9649,N_9556,N_9528);
or U9650 (N_9650,N_9485,N_9510);
nand U9651 (N_9651,N_9505,N_9474);
nor U9652 (N_9652,N_9484,N_9480);
xor U9653 (N_9653,N_9506,N_9573);
xor U9654 (N_9654,N_9586,N_9581);
nor U9655 (N_9655,N_9525,N_9477);
xnor U9656 (N_9656,N_9585,N_9426);
nand U9657 (N_9657,N_9470,N_9499);
nand U9658 (N_9658,N_9515,N_9598);
xnor U9659 (N_9659,N_9502,N_9568);
xor U9660 (N_9660,N_9440,N_9491);
or U9661 (N_9661,N_9445,N_9411);
nor U9662 (N_9662,N_9501,N_9536);
nor U9663 (N_9663,N_9579,N_9422);
nor U9664 (N_9664,N_9476,N_9416);
xor U9665 (N_9665,N_9432,N_9563);
xor U9666 (N_9666,N_9400,N_9454);
xnor U9667 (N_9667,N_9576,N_9420);
nor U9668 (N_9668,N_9446,N_9468);
and U9669 (N_9669,N_9517,N_9478);
xnor U9670 (N_9670,N_9518,N_9489);
nor U9671 (N_9671,N_9438,N_9558);
and U9672 (N_9672,N_9409,N_9425);
nand U9673 (N_9673,N_9531,N_9449);
nand U9674 (N_9674,N_9545,N_9496);
nor U9675 (N_9675,N_9516,N_9442);
nand U9676 (N_9676,N_9524,N_9459);
and U9677 (N_9677,N_9464,N_9521);
xnor U9678 (N_9678,N_9479,N_9463);
and U9679 (N_9679,N_9428,N_9583);
xor U9680 (N_9680,N_9465,N_9552);
nand U9681 (N_9681,N_9423,N_9569);
nand U9682 (N_9682,N_9452,N_9542);
or U9683 (N_9683,N_9572,N_9414);
and U9684 (N_9684,N_9487,N_9566);
nand U9685 (N_9685,N_9497,N_9526);
nand U9686 (N_9686,N_9450,N_9441);
xor U9687 (N_9687,N_9595,N_9486);
and U9688 (N_9688,N_9410,N_9540);
nand U9689 (N_9689,N_9592,N_9444);
or U9690 (N_9690,N_9546,N_9404);
or U9691 (N_9691,N_9421,N_9412);
nand U9692 (N_9692,N_9549,N_9530);
xnor U9693 (N_9693,N_9405,N_9575);
and U9694 (N_9694,N_9534,N_9460);
and U9695 (N_9695,N_9571,N_9562);
and U9696 (N_9696,N_9561,N_9565);
or U9697 (N_9697,N_9457,N_9599);
xnor U9698 (N_9698,N_9551,N_9435);
nand U9699 (N_9699,N_9589,N_9462);
nand U9700 (N_9700,N_9437,N_9448);
nand U9701 (N_9701,N_9402,N_9578);
nor U9702 (N_9702,N_9596,N_9473);
xor U9703 (N_9703,N_9509,N_9438);
nand U9704 (N_9704,N_9472,N_9444);
xor U9705 (N_9705,N_9536,N_9595);
nor U9706 (N_9706,N_9587,N_9584);
nor U9707 (N_9707,N_9567,N_9435);
and U9708 (N_9708,N_9417,N_9501);
nor U9709 (N_9709,N_9514,N_9506);
or U9710 (N_9710,N_9411,N_9556);
xor U9711 (N_9711,N_9558,N_9485);
xor U9712 (N_9712,N_9593,N_9415);
and U9713 (N_9713,N_9595,N_9517);
nand U9714 (N_9714,N_9550,N_9546);
nand U9715 (N_9715,N_9544,N_9452);
xor U9716 (N_9716,N_9462,N_9419);
nor U9717 (N_9717,N_9473,N_9551);
and U9718 (N_9718,N_9518,N_9448);
nand U9719 (N_9719,N_9535,N_9555);
and U9720 (N_9720,N_9449,N_9530);
and U9721 (N_9721,N_9526,N_9563);
nor U9722 (N_9722,N_9446,N_9560);
nand U9723 (N_9723,N_9486,N_9481);
nand U9724 (N_9724,N_9560,N_9509);
or U9725 (N_9725,N_9478,N_9490);
or U9726 (N_9726,N_9589,N_9479);
or U9727 (N_9727,N_9456,N_9494);
nand U9728 (N_9728,N_9483,N_9523);
nand U9729 (N_9729,N_9529,N_9400);
and U9730 (N_9730,N_9421,N_9467);
and U9731 (N_9731,N_9490,N_9453);
or U9732 (N_9732,N_9458,N_9568);
and U9733 (N_9733,N_9467,N_9557);
or U9734 (N_9734,N_9538,N_9474);
and U9735 (N_9735,N_9527,N_9581);
or U9736 (N_9736,N_9525,N_9485);
nor U9737 (N_9737,N_9431,N_9533);
nand U9738 (N_9738,N_9563,N_9513);
xor U9739 (N_9739,N_9472,N_9452);
xnor U9740 (N_9740,N_9595,N_9504);
or U9741 (N_9741,N_9475,N_9556);
nand U9742 (N_9742,N_9476,N_9525);
nor U9743 (N_9743,N_9500,N_9589);
or U9744 (N_9744,N_9540,N_9567);
nand U9745 (N_9745,N_9564,N_9433);
or U9746 (N_9746,N_9483,N_9531);
nor U9747 (N_9747,N_9485,N_9591);
xor U9748 (N_9748,N_9536,N_9514);
xnor U9749 (N_9749,N_9526,N_9410);
nor U9750 (N_9750,N_9514,N_9478);
xor U9751 (N_9751,N_9400,N_9521);
nor U9752 (N_9752,N_9430,N_9591);
and U9753 (N_9753,N_9511,N_9564);
and U9754 (N_9754,N_9427,N_9529);
or U9755 (N_9755,N_9555,N_9471);
nand U9756 (N_9756,N_9422,N_9514);
and U9757 (N_9757,N_9582,N_9578);
or U9758 (N_9758,N_9433,N_9516);
nor U9759 (N_9759,N_9545,N_9558);
nand U9760 (N_9760,N_9486,N_9537);
nand U9761 (N_9761,N_9418,N_9566);
xnor U9762 (N_9762,N_9531,N_9410);
nor U9763 (N_9763,N_9564,N_9524);
nor U9764 (N_9764,N_9465,N_9508);
nor U9765 (N_9765,N_9534,N_9589);
nand U9766 (N_9766,N_9476,N_9420);
and U9767 (N_9767,N_9424,N_9585);
and U9768 (N_9768,N_9577,N_9434);
nand U9769 (N_9769,N_9589,N_9402);
nand U9770 (N_9770,N_9439,N_9417);
xnor U9771 (N_9771,N_9538,N_9462);
and U9772 (N_9772,N_9450,N_9563);
and U9773 (N_9773,N_9564,N_9449);
and U9774 (N_9774,N_9483,N_9570);
nor U9775 (N_9775,N_9508,N_9467);
and U9776 (N_9776,N_9442,N_9525);
and U9777 (N_9777,N_9480,N_9573);
and U9778 (N_9778,N_9558,N_9503);
xnor U9779 (N_9779,N_9497,N_9505);
or U9780 (N_9780,N_9533,N_9568);
nand U9781 (N_9781,N_9498,N_9474);
or U9782 (N_9782,N_9519,N_9572);
xnor U9783 (N_9783,N_9550,N_9431);
or U9784 (N_9784,N_9467,N_9541);
and U9785 (N_9785,N_9476,N_9474);
and U9786 (N_9786,N_9567,N_9487);
nor U9787 (N_9787,N_9412,N_9540);
nand U9788 (N_9788,N_9467,N_9538);
nand U9789 (N_9789,N_9560,N_9556);
nor U9790 (N_9790,N_9545,N_9429);
or U9791 (N_9791,N_9576,N_9595);
or U9792 (N_9792,N_9575,N_9419);
and U9793 (N_9793,N_9400,N_9416);
or U9794 (N_9794,N_9591,N_9494);
nand U9795 (N_9795,N_9440,N_9400);
xnor U9796 (N_9796,N_9494,N_9485);
nand U9797 (N_9797,N_9461,N_9493);
nand U9798 (N_9798,N_9402,N_9552);
xnor U9799 (N_9799,N_9460,N_9598);
nor U9800 (N_9800,N_9637,N_9753);
nand U9801 (N_9801,N_9738,N_9727);
xor U9802 (N_9802,N_9726,N_9613);
nor U9803 (N_9803,N_9788,N_9716);
nor U9804 (N_9804,N_9799,N_9611);
nor U9805 (N_9805,N_9686,N_9772);
nand U9806 (N_9806,N_9707,N_9740);
and U9807 (N_9807,N_9660,N_9700);
nor U9808 (N_9808,N_9781,N_9650);
and U9809 (N_9809,N_9617,N_9705);
nand U9810 (N_9810,N_9688,N_9604);
or U9811 (N_9811,N_9677,N_9794);
or U9812 (N_9812,N_9666,N_9678);
xor U9813 (N_9813,N_9640,N_9724);
xnor U9814 (N_9814,N_9722,N_9693);
xor U9815 (N_9815,N_9602,N_9624);
nand U9816 (N_9816,N_9658,N_9786);
and U9817 (N_9817,N_9618,N_9751);
or U9818 (N_9818,N_9718,N_9605);
nor U9819 (N_9819,N_9736,N_9748);
nand U9820 (N_9820,N_9619,N_9723);
and U9821 (N_9821,N_9679,N_9770);
nor U9822 (N_9822,N_9649,N_9743);
xor U9823 (N_9823,N_9681,N_9787);
and U9824 (N_9824,N_9627,N_9702);
and U9825 (N_9825,N_9701,N_9714);
nand U9826 (N_9826,N_9720,N_9737);
nor U9827 (N_9827,N_9766,N_9725);
and U9828 (N_9828,N_9768,N_9783);
nand U9829 (N_9829,N_9663,N_9610);
nand U9830 (N_9830,N_9721,N_9710);
nor U9831 (N_9831,N_9691,N_9767);
and U9832 (N_9832,N_9796,N_9790);
xnor U9833 (N_9833,N_9667,N_9730);
nand U9834 (N_9834,N_9782,N_9762);
nand U9835 (N_9835,N_9797,N_9784);
xor U9836 (N_9836,N_9630,N_9747);
or U9837 (N_9837,N_9659,N_9646);
nand U9838 (N_9838,N_9697,N_9655);
and U9839 (N_9839,N_9636,N_9749);
nor U9840 (N_9840,N_9715,N_9795);
nor U9841 (N_9841,N_9684,N_9651);
xnor U9842 (N_9842,N_9616,N_9798);
or U9843 (N_9843,N_9759,N_9623);
nand U9844 (N_9844,N_9661,N_9756);
nand U9845 (N_9845,N_9670,N_9614);
and U9846 (N_9846,N_9744,N_9750);
xnor U9847 (N_9847,N_9741,N_9791);
nand U9848 (N_9848,N_9669,N_9779);
and U9849 (N_9849,N_9694,N_9746);
or U9850 (N_9850,N_9696,N_9755);
xor U9851 (N_9851,N_9785,N_9774);
or U9852 (N_9852,N_9682,N_9633);
nor U9853 (N_9853,N_9675,N_9628);
and U9854 (N_9854,N_9769,N_9625);
xor U9855 (N_9855,N_9644,N_9608);
nand U9856 (N_9856,N_9639,N_9763);
or U9857 (N_9857,N_9695,N_9776);
nand U9858 (N_9858,N_9754,N_9600);
or U9859 (N_9859,N_9671,N_9733);
nand U9860 (N_9860,N_9777,N_9728);
nand U9861 (N_9861,N_9745,N_9668);
xnor U9862 (N_9862,N_9778,N_9664);
nand U9863 (N_9863,N_9615,N_9752);
xor U9864 (N_9864,N_9775,N_9674);
nand U9865 (N_9865,N_9757,N_9621);
xor U9866 (N_9866,N_9711,N_9732);
and U9867 (N_9867,N_9719,N_9672);
nand U9868 (N_9868,N_9656,N_9680);
xor U9869 (N_9869,N_9789,N_9626);
nor U9870 (N_9870,N_9689,N_9687);
nand U9871 (N_9871,N_9676,N_9735);
xor U9872 (N_9872,N_9638,N_9706);
nor U9873 (N_9873,N_9758,N_9601);
and U9874 (N_9874,N_9662,N_9642);
xor U9875 (N_9875,N_9641,N_9606);
nor U9876 (N_9876,N_9652,N_9761);
or U9877 (N_9877,N_9692,N_9739);
xor U9878 (N_9878,N_9734,N_9629);
or U9879 (N_9879,N_9653,N_9742);
xor U9880 (N_9880,N_9632,N_9622);
or U9881 (N_9881,N_9773,N_9709);
nor U9882 (N_9882,N_9620,N_9713);
or U9883 (N_9883,N_9780,N_9673);
or U9884 (N_9884,N_9771,N_9654);
xnor U9885 (N_9885,N_9708,N_9731);
xnor U9886 (N_9886,N_9685,N_9603);
or U9887 (N_9887,N_9764,N_9712);
xnor U9888 (N_9888,N_9648,N_9631);
xor U9889 (N_9889,N_9643,N_9698);
nor U9890 (N_9890,N_9729,N_9635);
or U9891 (N_9891,N_9690,N_9793);
and U9892 (N_9892,N_9765,N_9634);
nand U9893 (N_9893,N_9703,N_9665);
xnor U9894 (N_9894,N_9607,N_9645);
xnor U9895 (N_9895,N_9657,N_9704);
nand U9896 (N_9896,N_9699,N_9717);
nor U9897 (N_9897,N_9612,N_9683);
nand U9898 (N_9898,N_9760,N_9609);
nor U9899 (N_9899,N_9792,N_9647);
nor U9900 (N_9900,N_9607,N_9610);
or U9901 (N_9901,N_9660,N_9725);
and U9902 (N_9902,N_9789,N_9700);
and U9903 (N_9903,N_9626,N_9622);
nand U9904 (N_9904,N_9623,N_9743);
nand U9905 (N_9905,N_9709,N_9641);
nand U9906 (N_9906,N_9768,N_9664);
xor U9907 (N_9907,N_9706,N_9702);
xor U9908 (N_9908,N_9634,N_9699);
nor U9909 (N_9909,N_9786,N_9775);
xor U9910 (N_9910,N_9631,N_9611);
nor U9911 (N_9911,N_9646,N_9624);
xnor U9912 (N_9912,N_9731,N_9610);
xnor U9913 (N_9913,N_9629,N_9611);
nand U9914 (N_9914,N_9689,N_9663);
xnor U9915 (N_9915,N_9744,N_9760);
or U9916 (N_9916,N_9773,N_9725);
or U9917 (N_9917,N_9648,N_9699);
nand U9918 (N_9918,N_9777,N_9617);
nor U9919 (N_9919,N_9766,N_9738);
and U9920 (N_9920,N_9661,N_9713);
and U9921 (N_9921,N_9796,N_9676);
xnor U9922 (N_9922,N_9765,N_9618);
and U9923 (N_9923,N_9642,N_9736);
xor U9924 (N_9924,N_9662,N_9651);
xnor U9925 (N_9925,N_9718,N_9717);
and U9926 (N_9926,N_9678,N_9743);
nor U9927 (N_9927,N_9630,N_9655);
xnor U9928 (N_9928,N_9612,N_9768);
nand U9929 (N_9929,N_9647,N_9616);
nor U9930 (N_9930,N_9684,N_9754);
or U9931 (N_9931,N_9761,N_9634);
nor U9932 (N_9932,N_9705,N_9723);
and U9933 (N_9933,N_9710,N_9731);
xnor U9934 (N_9934,N_9777,N_9722);
nand U9935 (N_9935,N_9700,N_9750);
or U9936 (N_9936,N_9773,N_9623);
or U9937 (N_9937,N_9757,N_9710);
nand U9938 (N_9938,N_9648,N_9725);
nor U9939 (N_9939,N_9645,N_9704);
nand U9940 (N_9940,N_9686,N_9765);
nand U9941 (N_9941,N_9658,N_9709);
nand U9942 (N_9942,N_9614,N_9782);
or U9943 (N_9943,N_9667,N_9612);
nand U9944 (N_9944,N_9757,N_9687);
xnor U9945 (N_9945,N_9694,N_9619);
nand U9946 (N_9946,N_9662,N_9641);
xnor U9947 (N_9947,N_9640,N_9799);
and U9948 (N_9948,N_9611,N_9626);
or U9949 (N_9949,N_9793,N_9624);
or U9950 (N_9950,N_9649,N_9674);
or U9951 (N_9951,N_9761,N_9716);
xnor U9952 (N_9952,N_9757,N_9729);
xor U9953 (N_9953,N_9628,N_9790);
or U9954 (N_9954,N_9768,N_9785);
nor U9955 (N_9955,N_9783,N_9761);
xor U9956 (N_9956,N_9709,N_9721);
and U9957 (N_9957,N_9676,N_9669);
nor U9958 (N_9958,N_9719,N_9610);
and U9959 (N_9959,N_9651,N_9627);
or U9960 (N_9960,N_9640,N_9697);
and U9961 (N_9961,N_9655,N_9665);
nand U9962 (N_9962,N_9675,N_9763);
nand U9963 (N_9963,N_9681,N_9702);
nand U9964 (N_9964,N_9601,N_9687);
xor U9965 (N_9965,N_9769,N_9732);
or U9966 (N_9966,N_9711,N_9759);
or U9967 (N_9967,N_9728,N_9748);
nand U9968 (N_9968,N_9641,N_9779);
and U9969 (N_9969,N_9675,N_9737);
or U9970 (N_9970,N_9691,N_9710);
or U9971 (N_9971,N_9610,N_9603);
and U9972 (N_9972,N_9723,N_9616);
nand U9973 (N_9973,N_9659,N_9640);
or U9974 (N_9974,N_9730,N_9706);
or U9975 (N_9975,N_9617,N_9765);
xor U9976 (N_9976,N_9734,N_9622);
or U9977 (N_9977,N_9706,N_9756);
or U9978 (N_9978,N_9791,N_9689);
xnor U9979 (N_9979,N_9764,N_9746);
xnor U9980 (N_9980,N_9783,N_9771);
and U9981 (N_9981,N_9647,N_9753);
and U9982 (N_9982,N_9609,N_9632);
nand U9983 (N_9983,N_9769,N_9632);
nand U9984 (N_9984,N_9670,N_9625);
and U9985 (N_9985,N_9762,N_9622);
nor U9986 (N_9986,N_9691,N_9716);
nand U9987 (N_9987,N_9614,N_9641);
or U9988 (N_9988,N_9600,N_9780);
and U9989 (N_9989,N_9638,N_9780);
and U9990 (N_9990,N_9697,N_9678);
and U9991 (N_9991,N_9602,N_9672);
nor U9992 (N_9992,N_9677,N_9669);
nand U9993 (N_9993,N_9643,N_9751);
and U9994 (N_9994,N_9731,N_9623);
nand U9995 (N_9995,N_9612,N_9725);
or U9996 (N_9996,N_9679,N_9647);
nand U9997 (N_9997,N_9780,N_9795);
and U9998 (N_9998,N_9725,N_9722);
nand U9999 (N_9999,N_9643,N_9624);
or U10000 (N_10000,N_9906,N_9968);
nor U10001 (N_10001,N_9976,N_9869);
nand U10002 (N_10002,N_9817,N_9847);
and U10003 (N_10003,N_9953,N_9830);
and U10004 (N_10004,N_9999,N_9842);
xnor U10005 (N_10005,N_9899,N_9850);
and U10006 (N_10006,N_9997,N_9972);
and U10007 (N_10007,N_9913,N_9879);
nor U10008 (N_10008,N_9813,N_9810);
nand U10009 (N_10009,N_9861,N_9802);
xor U10010 (N_10010,N_9880,N_9803);
or U10011 (N_10011,N_9852,N_9915);
nand U10012 (N_10012,N_9874,N_9979);
or U10013 (N_10013,N_9975,N_9833);
nor U10014 (N_10014,N_9834,N_9855);
or U10015 (N_10015,N_9991,N_9926);
xnor U10016 (N_10016,N_9934,N_9839);
or U10017 (N_10017,N_9912,N_9942);
or U10018 (N_10018,N_9966,N_9962);
xor U10019 (N_10019,N_9807,N_9887);
or U10020 (N_10020,N_9994,N_9846);
nand U10021 (N_10021,N_9933,N_9875);
nand U10022 (N_10022,N_9947,N_9925);
xor U10023 (N_10023,N_9808,N_9851);
and U10024 (N_10024,N_9963,N_9967);
and U10025 (N_10025,N_9965,N_9897);
nand U10026 (N_10026,N_9878,N_9911);
or U10027 (N_10027,N_9903,N_9956);
xor U10028 (N_10028,N_9800,N_9987);
nand U10029 (N_10029,N_9922,N_9931);
xor U10030 (N_10030,N_9998,N_9908);
xor U10031 (N_10031,N_9923,N_9992);
and U10032 (N_10032,N_9876,N_9973);
xor U10033 (N_10033,N_9881,N_9832);
xor U10034 (N_10034,N_9954,N_9894);
nand U10035 (N_10035,N_9980,N_9857);
xnor U10036 (N_10036,N_9905,N_9872);
xnor U10037 (N_10037,N_9820,N_9946);
nor U10038 (N_10038,N_9882,N_9936);
xor U10039 (N_10039,N_9841,N_9910);
and U10040 (N_10040,N_9868,N_9893);
nand U10041 (N_10041,N_9836,N_9819);
xor U10042 (N_10042,N_9930,N_9918);
nand U10043 (N_10043,N_9805,N_9939);
and U10044 (N_10044,N_9928,N_9891);
nor U10045 (N_10045,N_9951,N_9920);
nor U10046 (N_10046,N_9971,N_9974);
or U10047 (N_10047,N_9843,N_9858);
nand U10048 (N_10048,N_9990,N_9945);
nor U10049 (N_10049,N_9826,N_9900);
nand U10050 (N_10050,N_9961,N_9943);
nor U10051 (N_10051,N_9982,N_9827);
xor U10052 (N_10052,N_9937,N_9902);
or U10053 (N_10053,N_9977,N_9921);
nand U10054 (N_10054,N_9909,N_9960);
xor U10055 (N_10055,N_9995,N_9949);
nor U10056 (N_10056,N_9884,N_9811);
xnor U10057 (N_10057,N_9856,N_9862);
nor U10058 (N_10058,N_9993,N_9890);
or U10059 (N_10059,N_9941,N_9835);
nand U10060 (N_10060,N_9831,N_9818);
or U10061 (N_10061,N_9837,N_9886);
nor U10062 (N_10062,N_9932,N_9981);
and U10063 (N_10063,N_9950,N_9948);
xnor U10064 (N_10064,N_9804,N_9801);
xnor U10065 (N_10065,N_9929,N_9938);
nor U10066 (N_10066,N_9940,N_9848);
nand U10067 (N_10067,N_9959,N_9889);
and U10068 (N_10068,N_9863,N_9895);
xnor U10069 (N_10069,N_9957,N_9806);
xor U10070 (N_10070,N_9989,N_9907);
nand U10071 (N_10071,N_9904,N_9883);
nand U10072 (N_10072,N_9867,N_9916);
nand U10073 (N_10073,N_9944,N_9854);
or U10074 (N_10074,N_9914,N_9969);
or U10075 (N_10075,N_9935,N_9825);
and U10076 (N_10076,N_9823,N_9892);
nor U10077 (N_10077,N_9927,N_9919);
nand U10078 (N_10078,N_9838,N_9814);
nand U10079 (N_10079,N_9986,N_9970);
xnor U10080 (N_10080,N_9898,N_9844);
nor U10081 (N_10081,N_9865,N_9901);
xnor U10082 (N_10082,N_9870,N_9984);
nor U10083 (N_10083,N_9849,N_9821);
nor U10084 (N_10084,N_9809,N_9952);
nor U10085 (N_10085,N_9828,N_9958);
nor U10086 (N_10086,N_9822,N_9829);
and U10087 (N_10087,N_9866,N_9985);
or U10088 (N_10088,N_9978,N_9859);
or U10089 (N_10089,N_9864,N_9996);
and U10090 (N_10090,N_9873,N_9896);
nor U10091 (N_10091,N_9845,N_9871);
or U10092 (N_10092,N_9860,N_9924);
nor U10093 (N_10093,N_9840,N_9988);
nor U10094 (N_10094,N_9955,N_9964);
nor U10095 (N_10095,N_9815,N_9853);
xnor U10096 (N_10096,N_9885,N_9877);
nor U10097 (N_10097,N_9816,N_9812);
and U10098 (N_10098,N_9917,N_9983);
xor U10099 (N_10099,N_9888,N_9824);
and U10100 (N_10100,N_9968,N_9877);
nand U10101 (N_10101,N_9850,N_9978);
xnor U10102 (N_10102,N_9848,N_9974);
or U10103 (N_10103,N_9802,N_9881);
xor U10104 (N_10104,N_9931,N_9896);
or U10105 (N_10105,N_9844,N_9831);
nor U10106 (N_10106,N_9843,N_9913);
or U10107 (N_10107,N_9922,N_9980);
and U10108 (N_10108,N_9968,N_9806);
or U10109 (N_10109,N_9830,N_9856);
nor U10110 (N_10110,N_9917,N_9868);
xor U10111 (N_10111,N_9896,N_9814);
nor U10112 (N_10112,N_9943,N_9848);
nand U10113 (N_10113,N_9859,N_9935);
nand U10114 (N_10114,N_9919,N_9814);
nand U10115 (N_10115,N_9895,N_9834);
or U10116 (N_10116,N_9835,N_9812);
or U10117 (N_10117,N_9868,N_9822);
and U10118 (N_10118,N_9956,N_9975);
nor U10119 (N_10119,N_9837,N_9848);
nand U10120 (N_10120,N_9949,N_9940);
or U10121 (N_10121,N_9899,N_9808);
and U10122 (N_10122,N_9952,N_9855);
nor U10123 (N_10123,N_9860,N_9929);
and U10124 (N_10124,N_9900,N_9955);
and U10125 (N_10125,N_9934,N_9922);
and U10126 (N_10126,N_9969,N_9809);
or U10127 (N_10127,N_9978,N_9985);
xnor U10128 (N_10128,N_9859,N_9822);
nand U10129 (N_10129,N_9929,N_9807);
or U10130 (N_10130,N_9806,N_9898);
or U10131 (N_10131,N_9872,N_9856);
nand U10132 (N_10132,N_9930,N_9973);
and U10133 (N_10133,N_9848,N_9813);
and U10134 (N_10134,N_9895,N_9877);
xor U10135 (N_10135,N_9891,N_9885);
and U10136 (N_10136,N_9916,N_9905);
and U10137 (N_10137,N_9874,N_9918);
and U10138 (N_10138,N_9804,N_9883);
or U10139 (N_10139,N_9985,N_9837);
xnor U10140 (N_10140,N_9979,N_9982);
and U10141 (N_10141,N_9876,N_9997);
xor U10142 (N_10142,N_9804,N_9843);
or U10143 (N_10143,N_9839,N_9891);
nor U10144 (N_10144,N_9946,N_9905);
and U10145 (N_10145,N_9830,N_9917);
xor U10146 (N_10146,N_9870,N_9921);
or U10147 (N_10147,N_9858,N_9981);
xnor U10148 (N_10148,N_9974,N_9920);
or U10149 (N_10149,N_9896,N_9939);
nor U10150 (N_10150,N_9934,N_9873);
xor U10151 (N_10151,N_9852,N_9950);
and U10152 (N_10152,N_9929,N_9987);
or U10153 (N_10153,N_9937,N_9846);
nand U10154 (N_10154,N_9922,N_9930);
xor U10155 (N_10155,N_9977,N_9844);
and U10156 (N_10156,N_9875,N_9804);
or U10157 (N_10157,N_9998,N_9976);
nor U10158 (N_10158,N_9998,N_9888);
nor U10159 (N_10159,N_9861,N_9864);
nand U10160 (N_10160,N_9930,N_9877);
nand U10161 (N_10161,N_9903,N_9997);
nor U10162 (N_10162,N_9969,N_9859);
nor U10163 (N_10163,N_9975,N_9977);
nand U10164 (N_10164,N_9913,N_9995);
nor U10165 (N_10165,N_9873,N_9979);
and U10166 (N_10166,N_9800,N_9834);
nand U10167 (N_10167,N_9820,N_9843);
xnor U10168 (N_10168,N_9956,N_9872);
and U10169 (N_10169,N_9855,N_9965);
nand U10170 (N_10170,N_9893,N_9975);
and U10171 (N_10171,N_9993,N_9861);
nor U10172 (N_10172,N_9926,N_9857);
and U10173 (N_10173,N_9884,N_9842);
and U10174 (N_10174,N_9936,N_9834);
or U10175 (N_10175,N_9863,N_9978);
and U10176 (N_10176,N_9813,N_9800);
or U10177 (N_10177,N_9832,N_9965);
nor U10178 (N_10178,N_9981,N_9839);
xor U10179 (N_10179,N_9835,N_9826);
xor U10180 (N_10180,N_9817,N_9846);
nand U10181 (N_10181,N_9930,N_9872);
xor U10182 (N_10182,N_9893,N_9853);
xor U10183 (N_10183,N_9801,N_9967);
or U10184 (N_10184,N_9903,N_9805);
nand U10185 (N_10185,N_9810,N_9821);
nand U10186 (N_10186,N_9802,N_9974);
or U10187 (N_10187,N_9974,N_9898);
nand U10188 (N_10188,N_9987,N_9997);
xor U10189 (N_10189,N_9941,N_9816);
or U10190 (N_10190,N_9815,N_9900);
and U10191 (N_10191,N_9900,N_9989);
nand U10192 (N_10192,N_9959,N_9898);
or U10193 (N_10193,N_9812,N_9903);
xor U10194 (N_10194,N_9945,N_9846);
nand U10195 (N_10195,N_9967,N_9812);
nand U10196 (N_10196,N_9982,N_9873);
or U10197 (N_10197,N_9865,N_9837);
nor U10198 (N_10198,N_9862,N_9946);
xnor U10199 (N_10199,N_9888,N_9841);
nor U10200 (N_10200,N_10161,N_10143);
nand U10201 (N_10201,N_10162,N_10017);
nor U10202 (N_10202,N_10196,N_10120);
and U10203 (N_10203,N_10054,N_10199);
xnor U10204 (N_10204,N_10057,N_10156);
nor U10205 (N_10205,N_10087,N_10109);
nor U10206 (N_10206,N_10159,N_10106);
and U10207 (N_10207,N_10139,N_10023);
or U10208 (N_10208,N_10119,N_10135);
nand U10209 (N_10209,N_10146,N_10140);
xor U10210 (N_10210,N_10194,N_10163);
or U10211 (N_10211,N_10151,N_10021);
and U10212 (N_10212,N_10168,N_10075);
nand U10213 (N_10213,N_10197,N_10027);
nor U10214 (N_10214,N_10050,N_10175);
or U10215 (N_10215,N_10052,N_10051);
nand U10216 (N_10216,N_10071,N_10125);
xor U10217 (N_10217,N_10022,N_10015);
xnor U10218 (N_10218,N_10005,N_10011);
and U10219 (N_10219,N_10033,N_10186);
nand U10220 (N_10220,N_10141,N_10129);
and U10221 (N_10221,N_10095,N_10074);
nor U10222 (N_10222,N_10133,N_10184);
nand U10223 (N_10223,N_10097,N_10082);
xnor U10224 (N_10224,N_10032,N_10116);
nor U10225 (N_10225,N_10165,N_10157);
and U10226 (N_10226,N_10076,N_10100);
nand U10227 (N_10227,N_10180,N_10152);
and U10228 (N_10228,N_10073,N_10193);
nor U10229 (N_10229,N_10118,N_10144);
nor U10230 (N_10230,N_10093,N_10070);
nand U10231 (N_10231,N_10006,N_10124);
nor U10232 (N_10232,N_10062,N_10060);
and U10233 (N_10233,N_10134,N_10067);
nand U10234 (N_10234,N_10115,N_10037);
and U10235 (N_10235,N_10080,N_10104);
xnor U10236 (N_10236,N_10101,N_10049);
nor U10237 (N_10237,N_10189,N_10167);
or U10238 (N_10238,N_10108,N_10012);
and U10239 (N_10239,N_10092,N_10053);
nand U10240 (N_10240,N_10088,N_10113);
and U10241 (N_10241,N_10166,N_10036);
and U10242 (N_10242,N_10055,N_10091);
or U10243 (N_10243,N_10096,N_10081);
nand U10244 (N_10244,N_10103,N_10013);
nor U10245 (N_10245,N_10130,N_10182);
xor U10246 (N_10246,N_10153,N_10046);
xor U10247 (N_10247,N_10177,N_10179);
nor U10248 (N_10248,N_10077,N_10024);
nor U10249 (N_10249,N_10066,N_10138);
xnor U10250 (N_10250,N_10126,N_10031);
and U10251 (N_10251,N_10065,N_10034);
nand U10252 (N_10252,N_10147,N_10185);
nor U10253 (N_10253,N_10114,N_10112);
nor U10254 (N_10254,N_10018,N_10132);
nand U10255 (N_10255,N_10010,N_10121);
nor U10256 (N_10256,N_10009,N_10188);
xnor U10257 (N_10257,N_10145,N_10063);
and U10258 (N_10258,N_10154,N_10061);
and U10259 (N_10259,N_10086,N_10028);
xnor U10260 (N_10260,N_10000,N_10117);
and U10261 (N_10261,N_10084,N_10020);
nor U10262 (N_10262,N_10045,N_10122);
or U10263 (N_10263,N_10150,N_10002);
xnor U10264 (N_10264,N_10001,N_10072);
xor U10265 (N_10265,N_10110,N_10131);
nor U10266 (N_10266,N_10158,N_10160);
or U10267 (N_10267,N_10098,N_10048);
and U10268 (N_10268,N_10187,N_10085);
nand U10269 (N_10269,N_10004,N_10105);
or U10270 (N_10270,N_10079,N_10191);
xor U10271 (N_10271,N_10016,N_10178);
and U10272 (N_10272,N_10190,N_10025);
nand U10273 (N_10273,N_10170,N_10181);
and U10274 (N_10274,N_10083,N_10195);
nor U10275 (N_10275,N_10127,N_10149);
nor U10276 (N_10276,N_10058,N_10123);
xnor U10277 (N_10277,N_10089,N_10044);
nor U10278 (N_10278,N_10094,N_10111);
xor U10279 (N_10279,N_10099,N_10029);
and U10280 (N_10280,N_10068,N_10174);
or U10281 (N_10281,N_10090,N_10040);
or U10282 (N_10282,N_10183,N_10192);
nor U10283 (N_10283,N_10038,N_10198);
and U10284 (N_10284,N_10148,N_10026);
nand U10285 (N_10285,N_10155,N_10069);
nor U10286 (N_10286,N_10019,N_10007);
nor U10287 (N_10287,N_10102,N_10056);
xnor U10288 (N_10288,N_10176,N_10107);
or U10289 (N_10289,N_10035,N_10014);
nand U10290 (N_10290,N_10042,N_10137);
nand U10291 (N_10291,N_10171,N_10169);
or U10292 (N_10292,N_10030,N_10142);
nand U10293 (N_10293,N_10003,N_10128);
and U10294 (N_10294,N_10172,N_10064);
nand U10295 (N_10295,N_10047,N_10078);
and U10296 (N_10296,N_10039,N_10043);
nand U10297 (N_10297,N_10164,N_10041);
nor U10298 (N_10298,N_10008,N_10136);
xor U10299 (N_10299,N_10173,N_10059);
and U10300 (N_10300,N_10036,N_10000);
and U10301 (N_10301,N_10165,N_10093);
and U10302 (N_10302,N_10058,N_10061);
xor U10303 (N_10303,N_10081,N_10163);
xor U10304 (N_10304,N_10036,N_10018);
or U10305 (N_10305,N_10108,N_10037);
or U10306 (N_10306,N_10027,N_10038);
nor U10307 (N_10307,N_10133,N_10050);
nor U10308 (N_10308,N_10042,N_10142);
or U10309 (N_10309,N_10038,N_10033);
nor U10310 (N_10310,N_10013,N_10191);
or U10311 (N_10311,N_10175,N_10171);
nor U10312 (N_10312,N_10067,N_10086);
xor U10313 (N_10313,N_10161,N_10030);
xnor U10314 (N_10314,N_10022,N_10099);
nand U10315 (N_10315,N_10057,N_10190);
or U10316 (N_10316,N_10077,N_10055);
nand U10317 (N_10317,N_10109,N_10021);
nor U10318 (N_10318,N_10026,N_10054);
or U10319 (N_10319,N_10067,N_10018);
and U10320 (N_10320,N_10099,N_10177);
nor U10321 (N_10321,N_10151,N_10121);
and U10322 (N_10322,N_10159,N_10015);
xor U10323 (N_10323,N_10188,N_10015);
nor U10324 (N_10324,N_10124,N_10015);
xnor U10325 (N_10325,N_10098,N_10161);
or U10326 (N_10326,N_10084,N_10095);
xor U10327 (N_10327,N_10155,N_10024);
xnor U10328 (N_10328,N_10030,N_10136);
xnor U10329 (N_10329,N_10011,N_10068);
and U10330 (N_10330,N_10165,N_10194);
and U10331 (N_10331,N_10142,N_10018);
or U10332 (N_10332,N_10177,N_10162);
nand U10333 (N_10333,N_10064,N_10094);
and U10334 (N_10334,N_10123,N_10177);
nand U10335 (N_10335,N_10053,N_10170);
xor U10336 (N_10336,N_10113,N_10188);
nand U10337 (N_10337,N_10076,N_10173);
nand U10338 (N_10338,N_10191,N_10073);
and U10339 (N_10339,N_10070,N_10063);
xor U10340 (N_10340,N_10084,N_10037);
and U10341 (N_10341,N_10027,N_10096);
nor U10342 (N_10342,N_10034,N_10056);
nor U10343 (N_10343,N_10166,N_10195);
xnor U10344 (N_10344,N_10044,N_10095);
nor U10345 (N_10345,N_10015,N_10034);
nor U10346 (N_10346,N_10056,N_10189);
and U10347 (N_10347,N_10116,N_10103);
nor U10348 (N_10348,N_10157,N_10013);
or U10349 (N_10349,N_10184,N_10092);
nand U10350 (N_10350,N_10048,N_10022);
or U10351 (N_10351,N_10071,N_10072);
nand U10352 (N_10352,N_10153,N_10022);
nand U10353 (N_10353,N_10186,N_10035);
or U10354 (N_10354,N_10011,N_10036);
and U10355 (N_10355,N_10175,N_10158);
and U10356 (N_10356,N_10168,N_10042);
nor U10357 (N_10357,N_10085,N_10041);
nor U10358 (N_10358,N_10059,N_10189);
nor U10359 (N_10359,N_10004,N_10077);
and U10360 (N_10360,N_10119,N_10018);
xor U10361 (N_10361,N_10120,N_10042);
nand U10362 (N_10362,N_10049,N_10103);
nor U10363 (N_10363,N_10130,N_10017);
or U10364 (N_10364,N_10190,N_10182);
xor U10365 (N_10365,N_10159,N_10055);
xnor U10366 (N_10366,N_10038,N_10106);
and U10367 (N_10367,N_10098,N_10019);
nor U10368 (N_10368,N_10186,N_10178);
and U10369 (N_10369,N_10019,N_10080);
and U10370 (N_10370,N_10004,N_10146);
nand U10371 (N_10371,N_10021,N_10030);
or U10372 (N_10372,N_10007,N_10163);
nor U10373 (N_10373,N_10037,N_10154);
or U10374 (N_10374,N_10116,N_10008);
or U10375 (N_10375,N_10128,N_10092);
and U10376 (N_10376,N_10114,N_10070);
nor U10377 (N_10377,N_10040,N_10029);
and U10378 (N_10378,N_10023,N_10134);
nand U10379 (N_10379,N_10033,N_10018);
xnor U10380 (N_10380,N_10053,N_10091);
and U10381 (N_10381,N_10149,N_10178);
or U10382 (N_10382,N_10085,N_10130);
nor U10383 (N_10383,N_10054,N_10051);
nand U10384 (N_10384,N_10019,N_10048);
nand U10385 (N_10385,N_10005,N_10151);
and U10386 (N_10386,N_10040,N_10139);
and U10387 (N_10387,N_10165,N_10158);
nand U10388 (N_10388,N_10006,N_10155);
and U10389 (N_10389,N_10053,N_10136);
and U10390 (N_10390,N_10112,N_10177);
and U10391 (N_10391,N_10152,N_10038);
and U10392 (N_10392,N_10032,N_10178);
or U10393 (N_10393,N_10197,N_10012);
nand U10394 (N_10394,N_10126,N_10166);
xnor U10395 (N_10395,N_10011,N_10119);
nand U10396 (N_10396,N_10131,N_10045);
and U10397 (N_10397,N_10100,N_10066);
xor U10398 (N_10398,N_10189,N_10126);
and U10399 (N_10399,N_10114,N_10073);
nor U10400 (N_10400,N_10342,N_10392);
nor U10401 (N_10401,N_10347,N_10361);
nand U10402 (N_10402,N_10216,N_10237);
or U10403 (N_10403,N_10353,N_10238);
nand U10404 (N_10404,N_10358,N_10296);
nand U10405 (N_10405,N_10313,N_10396);
or U10406 (N_10406,N_10359,N_10217);
xor U10407 (N_10407,N_10256,N_10289);
and U10408 (N_10408,N_10239,N_10212);
and U10409 (N_10409,N_10262,N_10287);
nand U10410 (N_10410,N_10235,N_10299);
nand U10411 (N_10411,N_10246,N_10297);
xnor U10412 (N_10412,N_10382,N_10326);
nand U10413 (N_10413,N_10261,N_10288);
and U10414 (N_10414,N_10276,N_10220);
or U10415 (N_10415,N_10318,N_10316);
and U10416 (N_10416,N_10337,N_10380);
or U10417 (N_10417,N_10335,N_10245);
and U10418 (N_10418,N_10257,N_10203);
or U10419 (N_10419,N_10323,N_10312);
and U10420 (N_10420,N_10362,N_10320);
xor U10421 (N_10421,N_10329,N_10258);
or U10422 (N_10422,N_10305,N_10395);
and U10423 (N_10423,N_10300,N_10332);
xnor U10424 (N_10424,N_10346,N_10241);
or U10425 (N_10425,N_10221,N_10207);
xor U10426 (N_10426,N_10298,N_10222);
and U10427 (N_10427,N_10371,N_10247);
or U10428 (N_10428,N_10315,N_10374);
or U10429 (N_10429,N_10321,N_10253);
and U10430 (N_10430,N_10236,N_10223);
nor U10431 (N_10431,N_10204,N_10213);
or U10432 (N_10432,N_10279,N_10356);
and U10433 (N_10433,N_10202,N_10377);
xnor U10434 (N_10434,N_10277,N_10309);
and U10435 (N_10435,N_10384,N_10341);
and U10436 (N_10436,N_10366,N_10254);
xnor U10437 (N_10437,N_10283,N_10381);
xnor U10438 (N_10438,N_10227,N_10215);
or U10439 (N_10439,N_10306,N_10280);
nand U10440 (N_10440,N_10263,N_10225);
xor U10441 (N_10441,N_10228,N_10230);
xor U10442 (N_10442,N_10242,N_10345);
xnor U10443 (N_10443,N_10375,N_10268);
and U10444 (N_10444,N_10360,N_10340);
nor U10445 (N_10445,N_10229,N_10385);
nor U10446 (N_10446,N_10387,N_10363);
and U10447 (N_10447,N_10378,N_10388);
and U10448 (N_10448,N_10324,N_10301);
or U10449 (N_10449,N_10255,N_10325);
and U10450 (N_10450,N_10267,N_10368);
or U10451 (N_10451,N_10249,N_10372);
and U10452 (N_10452,N_10354,N_10350);
nand U10453 (N_10453,N_10344,N_10349);
and U10454 (N_10454,N_10339,N_10351);
or U10455 (N_10455,N_10328,N_10302);
nor U10456 (N_10456,N_10333,N_10369);
and U10457 (N_10457,N_10248,N_10376);
nor U10458 (N_10458,N_10226,N_10367);
nor U10459 (N_10459,N_10281,N_10206);
and U10460 (N_10460,N_10365,N_10370);
xnor U10461 (N_10461,N_10210,N_10291);
and U10462 (N_10462,N_10303,N_10201);
and U10463 (N_10463,N_10269,N_10355);
or U10464 (N_10464,N_10211,N_10373);
and U10465 (N_10465,N_10244,N_10391);
or U10466 (N_10466,N_10292,N_10271);
or U10467 (N_10467,N_10294,N_10250);
or U10468 (N_10468,N_10322,N_10352);
nor U10469 (N_10469,N_10272,N_10314);
and U10470 (N_10470,N_10334,N_10266);
or U10471 (N_10471,N_10398,N_10307);
xnor U10472 (N_10472,N_10264,N_10209);
nand U10473 (N_10473,N_10331,N_10393);
xor U10474 (N_10474,N_10286,N_10295);
and U10475 (N_10475,N_10310,N_10214);
or U10476 (N_10476,N_10319,N_10265);
and U10477 (N_10477,N_10243,N_10275);
or U10478 (N_10478,N_10386,N_10327);
and U10479 (N_10479,N_10338,N_10251);
xnor U10480 (N_10480,N_10308,N_10304);
nor U10481 (N_10481,N_10336,N_10232);
and U10482 (N_10482,N_10397,N_10390);
and U10483 (N_10483,N_10357,N_10274);
or U10484 (N_10484,N_10219,N_10311);
and U10485 (N_10485,N_10224,N_10284);
and U10486 (N_10486,N_10273,N_10285);
and U10487 (N_10487,N_10317,N_10252);
and U10488 (N_10488,N_10348,N_10379);
nor U10489 (N_10489,N_10394,N_10200);
or U10490 (N_10490,N_10234,N_10231);
nand U10491 (N_10491,N_10364,N_10270);
xnor U10492 (N_10492,N_10259,N_10218);
xor U10493 (N_10493,N_10343,N_10233);
nand U10494 (N_10494,N_10205,N_10389);
and U10495 (N_10495,N_10330,N_10399);
nor U10496 (N_10496,N_10240,N_10260);
nor U10497 (N_10497,N_10278,N_10293);
nor U10498 (N_10498,N_10208,N_10383);
and U10499 (N_10499,N_10282,N_10290);
xnor U10500 (N_10500,N_10319,N_10252);
xor U10501 (N_10501,N_10331,N_10245);
nor U10502 (N_10502,N_10283,N_10266);
xor U10503 (N_10503,N_10266,N_10383);
nor U10504 (N_10504,N_10219,N_10388);
nand U10505 (N_10505,N_10384,N_10262);
or U10506 (N_10506,N_10368,N_10292);
or U10507 (N_10507,N_10308,N_10336);
nor U10508 (N_10508,N_10237,N_10258);
nor U10509 (N_10509,N_10262,N_10305);
xor U10510 (N_10510,N_10390,N_10280);
and U10511 (N_10511,N_10271,N_10216);
nand U10512 (N_10512,N_10286,N_10332);
or U10513 (N_10513,N_10397,N_10333);
xnor U10514 (N_10514,N_10275,N_10319);
or U10515 (N_10515,N_10399,N_10268);
xnor U10516 (N_10516,N_10302,N_10295);
and U10517 (N_10517,N_10362,N_10228);
xnor U10518 (N_10518,N_10306,N_10261);
xnor U10519 (N_10519,N_10348,N_10287);
nand U10520 (N_10520,N_10341,N_10391);
and U10521 (N_10521,N_10220,N_10312);
or U10522 (N_10522,N_10292,N_10391);
nand U10523 (N_10523,N_10339,N_10237);
nor U10524 (N_10524,N_10255,N_10353);
or U10525 (N_10525,N_10244,N_10327);
or U10526 (N_10526,N_10277,N_10374);
nor U10527 (N_10527,N_10261,N_10234);
or U10528 (N_10528,N_10301,N_10348);
and U10529 (N_10529,N_10255,N_10203);
and U10530 (N_10530,N_10286,N_10241);
and U10531 (N_10531,N_10394,N_10338);
nor U10532 (N_10532,N_10225,N_10224);
nand U10533 (N_10533,N_10215,N_10253);
nand U10534 (N_10534,N_10279,N_10243);
and U10535 (N_10535,N_10212,N_10253);
and U10536 (N_10536,N_10341,N_10235);
xor U10537 (N_10537,N_10357,N_10254);
and U10538 (N_10538,N_10252,N_10246);
and U10539 (N_10539,N_10281,N_10276);
and U10540 (N_10540,N_10398,N_10313);
nand U10541 (N_10541,N_10399,N_10252);
or U10542 (N_10542,N_10293,N_10342);
nor U10543 (N_10543,N_10219,N_10348);
and U10544 (N_10544,N_10270,N_10290);
or U10545 (N_10545,N_10202,N_10221);
or U10546 (N_10546,N_10351,N_10218);
xor U10547 (N_10547,N_10214,N_10255);
and U10548 (N_10548,N_10340,N_10267);
or U10549 (N_10549,N_10225,N_10353);
nor U10550 (N_10550,N_10332,N_10273);
or U10551 (N_10551,N_10206,N_10370);
nand U10552 (N_10552,N_10293,N_10390);
and U10553 (N_10553,N_10373,N_10317);
or U10554 (N_10554,N_10236,N_10224);
and U10555 (N_10555,N_10320,N_10387);
xnor U10556 (N_10556,N_10353,N_10380);
xor U10557 (N_10557,N_10329,N_10334);
and U10558 (N_10558,N_10246,N_10342);
nor U10559 (N_10559,N_10296,N_10242);
nor U10560 (N_10560,N_10331,N_10246);
and U10561 (N_10561,N_10276,N_10296);
nand U10562 (N_10562,N_10371,N_10273);
or U10563 (N_10563,N_10359,N_10371);
and U10564 (N_10564,N_10279,N_10316);
or U10565 (N_10565,N_10279,N_10340);
xor U10566 (N_10566,N_10374,N_10270);
xnor U10567 (N_10567,N_10234,N_10314);
or U10568 (N_10568,N_10351,N_10364);
nand U10569 (N_10569,N_10290,N_10388);
and U10570 (N_10570,N_10238,N_10213);
nor U10571 (N_10571,N_10219,N_10380);
nand U10572 (N_10572,N_10346,N_10252);
nand U10573 (N_10573,N_10268,N_10214);
and U10574 (N_10574,N_10264,N_10229);
xnor U10575 (N_10575,N_10242,N_10233);
nand U10576 (N_10576,N_10268,N_10336);
nand U10577 (N_10577,N_10276,N_10268);
and U10578 (N_10578,N_10291,N_10286);
nand U10579 (N_10579,N_10336,N_10287);
xnor U10580 (N_10580,N_10218,N_10326);
or U10581 (N_10581,N_10379,N_10243);
or U10582 (N_10582,N_10243,N_10281);
or U10583 (N_10583,N_10296,N_10277);
nor U10584 (N_10584,N_10231,N_10270);
nand U10585 (N_10585,N_10323,N_10265);
nand U10586 (N_10586,N_10356,N_10320);
xnor U10587 (N_10587,N_10356,N_10263);
nand U10588 (N_10588,N_10246,N_10220);
xor U10589 (N_10589,N_10205,N_10393);
nand U10590 (N_10590,N_10263,N_10292);
nor U10591 (N_10591,N_10319,N_10211);
xor U10592 (N_10592,N_10379,N_10373);
or U10593 (N_10593,N_10224,N_10364);
nand U10594 (N_10594,N_10357,N_10363);
nor U10595 (N_10595,N_10331,N_10204);
and U10596 (N_10596,N_10251,N_10346);
and U10597 (N_10597,N_10367,N_10215);
and U10598 (N_10598,N_10226,N_10323);
xor U10599 (N_10599,N_10209,N_10218);
nor U10600 (N_10600,N_10405,N_10568);
xnor U10601 (N_10601,N_10547,N_10514);
xnor U10602 (N_10602,N_10455,N_10584);
xor U10603 (N_10603,N_10432,N_10565);
or U10604 (N_10604,N_10556,N_10437);
nor U10605 (N_10605,N_10444,N_10548);
nand U10606 (N_10606,N_10517,N_10597);
xor U10607 (N_10607,N_10567,N_10577);
nor U10608 (N_10608,N_10500,N_10454);
nor U10609 (N_10609,N_10477,N_10491);
nand U10610 (N_10610,N_10490,N_10442);
nand U10611 (N_10611,N_10531,N_10504);
or U10612 (N_10612,N_10403,N_10559);
and U10613 (N_10613,N_10428,N_10520);
nand U10614 (N_10614,N_10507,N_10519);
or U10615 (N_10615,N_10553,N_10552);
xnor U10616 (N_10616,N_10571,N_10449);
nor U10617 (N_10617,N_10511,N_10594);
nand U10618 (N_10618,N_10440,N_10588);
or U10619 (N_10619,N_10536,N_10471);
nand U10620 (N_10620,N_10558,N_10469);
nor U10621 (N_10621,N_10581,N_10421);
xor U10622 (N_10622,N_10410,N_10466);
nor U10623 (N_10623,N_10516,N_10554);
nor U10624 (N_10624,N_10537,N_10586);
xnor U10625 (N_10625,N_10578,N_10473);
or U10626 (N_10626,N_10420,N_10475);
nand U10627 (N_10627,N_10435,N_10484);
or U10628 (N_10628,N_10515,N_10546);
or U10629 (N_10629,N_10541,N_10417);
nand U10630 (N_10630,N_10443,N_10446);
or U10631 (N_10631,N_10412,N_10564);
nand U10632 (N_10632,N_10599,N_10439);
or U10633 (N_10633,N_10427,N_10463);
nor U10634 (N_10634,N_10423,N_10573);
or U10635 (N_10635,N_10487,N_10465);
and U10636 (N_10636,N_10489,N_10575);
or U10637 (N_10637,N_10415,N_10461);
or U10638 (N_10638,N_10524,N_10512);
or U10639 (N_10639,N_10596,N_10464);
and U10640 (N_10640,N_10457,N_10431);
nor U10641 (N_10641,N_10572,N_10458);
nor U10642 (N_10642,N_10555,N_10562);
or U10643 (N_10643,N_10496,N_10425);
and U10644 (N_10644,N_10462,N_10509);
nor U10645 (N_10645,N_10402,N_10445);
nand U10646 (N_10646,N_10503,N_10563);
and U10647 (N_10647,N_10585,N_10478);
nor U10648 (N_10648,N_10545,N_10406);
or U10649 (N_10649,N_10583,N_10413);
nand U10650 (N_10650,N_10485,N_10540);
nor U10651 (N_10651,N_10570,N_10522);
or U10652 (N_10652,N_10539,N_10538);
nor U10653 (N_10653,N_10416,N_10459);
nor U10654 (N_10654,N_10419,N_10560);
nor U10655 (N_10655,N_10476,N_10430);
nand U10656 (N_10656,N_10441,N_10498);
and U10657 (N_10657,N_10530,N_10506);
nor U10658 (N_10658,N_10479,N_10591);
nor U10659 (N_10659,N_10401,N_10598);
and U10660 (N_10660,N_10521,N_10549);
xnor U10661 (N_10661,N_10529,N_10486);
or U10662 (N_10662,N_10448,N_10502);
nor U10663 (N_10663,N_10580,N_10480);
nor U10664 (N_10664,N_10424,N_10470);
nand U10665 (N_10665,N_10468,N_10418);
nand U10666 (N_10666,N_10535,N_10408);
nand U10667 (N_10667,N_10482,N_10561);
nand U10668 (N_10668,N_10542,N_10497);
nand U10669 (N_10669,N_10422,N_10447);
nor U10670 (N_10670,N_10550,N_10579);
nand U10671 (N_10671,N_10429,N_10544);
nand U10672 (N_10672,N_10557,N_10495);
or U10673 (N_10673,N_10436,N_10513);
nor U10674 (N_10674,N_10518,N_10407);
nor U10675 (N_10675,N_10569,N_10523);
nor U10676 (N_10676,N_10404,N_10438);
nor U10677 (N_10677,N_10499,N_10574);
or U10678 (N_10678,N_10501,N_10409);
nand U10679 (N_10679,N_10526,N_10426);
nor U10680 (N_10680,N_10453,N_10593);
xnor U10681 (N_10681,N_10534,N_10488);
nor U10682 (N_10682,N_10576,N_10450);
xor U10683 (N_10683,N_10505,N_10411);
and U10684 (N_10684,N_10527,N_10492);
and U10685 (N_10685,N_10460,N_10434);
or U10686 (N_10686,N_10582,N_10551);
xor U10687 (N_10687,N_10433,N_10474);
xor U10688 (N_10688,N_10528,N_10494);
nand U10689 (N_10689,N_10595,N_10543);
or U10690 (N_10690,N_10566,N_10533);
nand U10691 (N_10691,N_10532,N_10525);
and U10692 (N_10692,N_10508,N_10451);
xnor U10693 (N_10693,N_10589,N_10510);
xor U10694 (N_10694,N_10414,N_10472);
nor U10695 (N_10695,N_10493,N_10590);
nor U10696 (N_10696,N_10452,N_10456);
or U10697 (N_10697,N_10400,N_10483);
and U10698 (N_10698,N_10467,N_10587);
or U10699 (N_10699,N_10592,N_10481);
xnor U10700 (N_10700,N_10589,N_10532);
or U10701 (N_10701,N_10498,N_10460);
xor U10702 (N_10702,N_10487,N_10535);
and U10703 (N_10703,N_10529,N_10497);
or U10704 (N_10704,N_10531,N_10400);
xor U10705 (N_10705,N_10596,N_10537);
and U10706 (N_10706,N_10537,N_10405);
nand U10707 (N_10707,N_10487,N_10590);
nor U10708 (N_10708,N_10438,N_10538);
or U10709 (N_10709,N_10445,N_10527);
or U10710 (N_10710,N_10587,N_10475);
and U10711 (N_10711,N_10550,N_10492);
nand U10712 (N_10712,N_10580,N_10404);
xor U10713 (N_10713,N_10436,N_10400);
or U10714 (N_10714,N_10487,N_10466);
nor U10715 (N_10715,N_10433,N_10414);
and U10716 (N_10716,N_10571,N_10455);
and U10717 (N_10717,N_10466,N_10559);
nand U10718 (N_10718,N_10490,N_10509);
xor U10719 (N_10719,N_10404,N_10526);
xnor U10720 (N_10720,N_10571,N_10560);
nor U10721 (N_10721,N_10422,N_10401);
and U10722 (N_10722,N_10447,N_10487);
or U10723 (N_10723,N_10577,N_10575);
and U10724 (N_10724,N_10546,N_10598);
or U10725 (N_10725,N_10519,N_10571);
nand U10726 (N_10726,N_10428,N_10489);
nor U10727 (N_10727,N_10561,N_10402);
or U10728 (N_10728,N_10482,N_10525);
xnor U10729 (N_10729,N_10575,N_10568);
xnor U10730 (N_10730,N_10507,N_10548);
or U10731 (N_10731,N_10570,N_10444);
or U10732 (N_10732,N_10560,N_10443);
or U10733 (N_10733,N_10446,N_10571);
nor U10734 (N_10734,N_10570,N_10568);
nand U10735 (N_10735,N_10570,N_10510);
and U10736 (N_10736,N_10400,N_10571);
and U10737 (N_10737,N_10454,N_10538);
and U10738 (N_10738,N_10522,N_10590);
nor U10739 (N_10739,N_10501,N_10455);
or U10740 (N_10740,N_10515,N_10410);
or U10741 (N_10741,N_10408,N_10506);
and U10742 (N_10742,N_10574,N_10549);
nor U10743 (N_10743,N_10580,N_10432);
nor U10744 (N_10744,N_10505,N_10551);
nor U10745 (N_10745,N_10498,N_10525);
and U10746 (N_10746,N_10540,N_10504);
nand U10747 (N_10747,N_10455,N_10508);
nor U10748 (N_10748,N_10525,N_10573);
nand U10749 (N_10749,N_10430,N_10554);
or U10750 (N_10750,N_10401,N_10520);
nor U10751 (N_10751,N_10592,N_10469);
nand U10752 (N_10752,N_10535,N_10509);
or U10753 (N_10753,N_10468,N_10582);
xnor U10754 (N_10754,N_10429,N_10504);
nor U10755 (N_10755,N_10565,N_10515);
nand U10756 (N_10756,N_10452,N_10497);
xor U10757 (N_10757,N_10403,N_10539);
nor U10758 (N_10758,N_10526,N_10584);
nor U10759 (N_10759,N_10542,N_10595);
nor U10760 (N_10760,N_10583,N_10562);
and U10761 (N_10761,N_10492,N_10501);
and U10762 (N_10762,N_10588,N_10554);
nor U10763 (N_10763,N_10586,N_10492);
or U10764 (N_10764,N_10568,N_10469);
xnor U10765 (N_10765,N_10410,N_10431);
and U10766 (N_10766,N_10429,N_10546);
nand U10767 (N_10767,N_10540,N_10432);
nand U10768 (N_10768,N_10517,N_10416);
or U10769 (N_10769,N_10551,N_10589);
xor U10770 (N_10770,N_10472,N_10567);
nand U10771 (N_10771,N_10585,N_10510);
nand U10772 (N_10772,N_10417,N_10484);
nor U10773 (N_10773,N_10516,N_10437);
or U10774 (N_10774,N_10470,N_10584);
and U10775 (N_10775,N_10538,N_10473);
nor U10776 (N_10776,N_10561,N_10533);
nor U10777 (N_10777,N_10494,N_10579);
or U10778 (N_10778,N_10594,N_10531);
and U10779 (N_10779,N_10414,N_10501);
nor U10780 (N_10780,N_10480,N_10592);
and U10781 (N_10781,N_10536,N_10558);
xor U10782 (N_10782,N_10460,N_10480);
and U10783 (N_10783,N_10442,N_10527);
and U10784 (N_10784,N_10500,N_10447);
nand U10785 (N_10785,N_10502,N_10423);
nand U10786 (N_10786,N_10473,N_10478);
nor U10787 (N_10787,N_10544,N_10524);
nand U10788 (N_10788,N_10467,N_10585);
nor U10789 (N_10789,N_10567,N_10534);
or U10790 (N_10790,N_10425,N_10570);
nand U10791 (N_10791,N_10541,N_10550);
xor U10792 (N_10792,N_10595,N_10407);
and U10793 (N_10793,N_10517,N_10545);
nor U10794 (N_10794,N_10480,N_10573);
nand U10795 (N_10795,N_10556,N_10403);
or U10796 (N_10796,N_10430,N_10496);
nor U10797 (N_10797,N_10479,N_10476);
and U10798 (N_10798,N_10502,N_10442);
and U10799 (N_10799,N_10596,N_10568);
or U10800 (N_10800,N_10603,N_10638);
or U10801 (N_10801,N_10715,N_10664);
nor U10802 (N_10802,N_10666,N_10692);
and U10803 (N_10803,N_10689,N_10799);
or U10804 (N_10804,N_10651,N_10703);
and U10805 (N_10805,N_10759,N_10648);
or U10806 (N_10806,N_10627,N_10660);
nor U10807 (N_10807,N_10657,N_10626);
and U10808 (N_10808,N_10676,N_10702);
nor U10809 (N_10809,N_10613,N_10643);
nor U10810 (N_10810,N_10795,N_10693);
or U10811 (N_10811,N_10671,N_10680);
xor U10812 (N_10812,N_10734,N_10719);
nand U10813 (N_10813,N_10681,N_10729);
and U10814 (N_10814,N_10611,N_10764);
nand U10815 (N_10815,N_10695,N_10788);
and U10816 (N_10816,N_10622,N_10767);
xor U10817 (N_10817,N_10748,N_10645);
and U10818 (N_10818,N_10683,N_10667);
or U10819 (N_10819,N_10737,N_10757);
nand U10820 (N_10820,N_10725,N_10605);
nand U10821 (N_10821,N_10754,N_10650);
nand U10822 (N_10822,N_10608,N_10717);
xnor U10823 (N_10823,N_10750,N_10762);
and U10824 (N_10824,N_10728,N_10712);
nand U10825 (N_10825,N_10674,N_10639);
or U10826 (N_10826,N_10735,N_10632);
or U10827 (N_10827,N_10721,N_10615);
or U10828 (N_10828,N_10786,N_10624);
or U10829 (N_10829,N_10709,N_10656);
nand U10830 (N_10830,N_10704,N_10701);
nand U10831 (N_10831,N_10647,N_10787);
nand U10832 (N_10832,N_10773,N_10600);
nand U10833 (N_10833,N_10746,N_10636);
nand U10834 (N_10834,N_10637,N_10714);
nand U10835 (N_10835,N_10687,N_10634);
and U10836 (N_10836,N_10672,N_10768);
and U10837 (N_10837,N_10760,N_10630);
xnor U10838 (N_10838,N_10783,N_10614);
or U10839 (N_10839,N_10744,N_10722);
xnor U10840 (N_10840,N_10619,N_10677);
nor U10841 (N_10841,N_10780,N_10742);
nor U10842 (N_10842,N_10606,N_10623);
or U10843 (N_10843,N_10752,N_10662);
or U10844 (N_10844,N_10694,N_10708);
or U10845 (N_10845,N_10724,N_10755);
or U10846 (N_10846,N_10775,N_10751);
xor U10847 (N_10847,N_10690,N_10732);
nand U10848 (N_10848,N_10670,N_10716);
nand U10849 (N_10849,N_10733,N_10731);
nand U10850 (N_10850,N_10718,N_10763);
nor U10851 (N_10851,N_10642,N_10779);
xor U10852 (N_10852,N_10659,N_10641);
xor U10853 (N_10853,N_10743,N_10796);
nand U10854 (N_10854,N_10798,N_10635);
xor U10855 (N_10855,N_10723,N_10730);
or U10856 (N_10856,N_10761,N_10617);
nand U10857 (N_10857,N_10685,N_10663);
xnor U10858 (N_10858,N_10785,N_10697);
xnor U10859 (N_10859,N_10777,N_10612);
nor U10860 (N_10860,N_10726,N_10640);
or U10861 (N_10861,N_10609,N_10747);
xnor U10862 (N_10862,N_10698,N_10668);
nand U10863 (N_10863,N_10625,N_10713);
xor U10864 (N_10864,N_10602,N_10684);
or U10865 (N_10865,N_10601,N_10688);
xor U10866 (N_10866,N_10618,N_10629);
nand U10867 (N_10867,N_10654,N_10792);
xor U10868 (N_10868,N_10706,N_10628);
xor U10869 (N_10869,N_10772,N_10720);
or U10870 (N_10870,N_10631,N_10644);
nand U10871 (N_10871,N_10679,N_10793);
xnor U10872 (N_10872,N_10710,N_10749);
nor U10873 (N_10873,N_10661,N_10711);
and U10874 (N_10874,N_10782,N_10705);
and U10875 (N_10875,N_10691,N_10784);
nor U10876 (N_10876,N_10739,N_10652);
or U10877 (N_10877,N_10673,N_10769);
or U10878 (N_10878,N_10736,N_10610);
nand U10879 (N_10879,N_10707,N_10604);
nand U10880 (N_10880,N_10655,N_10649);
xor U10881 (N_10881,N_10620,N_10616);
or U10882 (N_10882,N_10794,N_10665);
nor U10883 (N_10883,N_10646,N_10621);
nor U10884 (N_10884,N_10653,N_10682);
or U10885 (N_10885,N_10789,N_10770);
or U10886 (N_10886,N_10774,N_10778);
xor U10887 (N_10887,N_10727,N_10765);
nand U10888 (N_10888,N_10766,N_10633);
or U10889 (N_10889,N_10699,N_10776);
xnor U10890 (N_10890,N_10658,N_10758);
and U10891 (N_10891,N_10738,N_10741);
or U10892 (N_10892,N_10675,N_10696);
nand U10893 (N_10893,N_10753,N_10700);
or U10894 (N_10894,N_10745,N_10607);
and U10895 (N_10895,N_10686,N_10756);
and U10896 (N_10896,N_10797,N_10791);
nor U10897 (N_10897,N_10771,N_10740);
and U10898 (N_10898,N_10669,N_10790);
or U10899 (N_10899,N_10678,N_10781);
or U10900 (N_10900,N_10650,N_10783);
nand U10901 (N_10901,N_10664,N_10632);
nor U10902 (N_10902,N_10744,N_10607);
nand U10903 (N_10903,N_10641,N_10648);
nand U10904 (N_10904,N_10769,N_10787);
and U10905 (N_10905,N_10771,N_10722);
or U10906 (N_10906,N_10748,N_10786);
nand U10907 (N_10907,N_10699,N_10711);
nand U10908 (N_10908,N_10685,N_10655);
xnor U10909 (N_10909,N_10607,N_10644);
or U10910 (N_10910,N_10768,N_10670);
nand U10911 (N_10911,N_10662,N_10708);
xor U10912 (N_10912,N_10625,N_10623);
xnor U10913 (N_10913,N_10631,N_10683);
or U10914 (N_10914,N_10798,N_10661);
xor U10915 (N_10915,N_10696,N_10724);
nor U10916 (N_10916,N_10710,N_10669);
xnor U10917 (N_10917,N_10775,N_10695);
and U10918 (N_10918,N_10707,N_10626);
and U10919 (N_10919,N_10652,N_10602);
nor U10920 (N_10920,N_10729,N_10627);
and U10921 (N_10921,N_10698,N_10665);
xor U10922 (N_10922,N_10778,N_10646);
xor U10923 (N_10923,N_10659,N_10751);
or U10924 (N_10924,N_10729,N_10611);
xor U10925 (N_10925,N_10623,N_10744);
and U10926 (N_10926,N_10720,N_10613);
xnor U10927 (N_10927,N_10745,N_10673);
nand U10928 (N_10928,N_10767,N_10727);
or U10929 (N_10929,N_10652,N_10634);
or U10930 (N_10930,N_10653,N_10678);
nand U10931 (N_10931,N_10637,N_10747);
xnor U10932 (N_10932,N_10654,N_10645);
nor U10933 (N_10933,N_10768,N_10709);
nor U10934 (N_10934,N_10786,N_10717);
or U10935 (N_10935,N_10722,N_10742);
nor U10936 (N_10936,N_10787,N_10749);
xnor U10937 (N_10937,N_10635,N_10647);
xnor U10938 (N_10938,N_10780,N_10637);
and U10939 (N_10939,N_10689,N_10679);
nor U10940 (N_10940,N_10689,N_10645);
or U10941 (N_10941,N_10698,N_10704);
or U10942 (N_10942,N_10668,N_10683);
xnor U10943 (N_10943,N_10774,N_10667);
nand U10944 (N_10944,N_10752,N_10743);
nor U10945 (N_10945,N_10752,N_10750);
nor U10946 (N_10946,N_10678,N_10724);
xor U10947 (N_10947,N_10621,N_10730);
nand U10948 (N_10948,N_10645,N_10749);
nand U10949 (N_10949,N_10618,N_10665);
xor U10950 (N_10950,N_10758,N_10709);
nand U10951 (N_10951,N_10744,N_10619);
and U10952 (N_10952,N_10712,N_10683);
xor U10953 (N_10953,N_10762,N_10679);
and U10954 (N_10954,N_10667,N_10635);
and U10955 (N_10955,N_10636,N_10624);
nand U10956 (N_10956,N_10797,N_10780);
nand U10957 (N_10957,N_10731,N_10715);
or U10958 (N_10958,N_10645,N_10729);
nand U10959 (N_10959,N_10772,N_10742);
nand U10960 (N_10960,N_10785,N_10793);
and U10961 (N_10961,N_10693,N_10762);
nor U10962 (N_10962,N_10757,N_10638);
and U10963 (N_10963,N_10609,N_10722);
nand U10964 (N_10964,N_10709,N_10624);
or U10965 (N_10965,N_10787,N_10691);
nand U10966 (N_10966,N_10709,N_10776);
and U10967 (N_10967,N_10696,N_10725);
or U10968 (N_10968,N_10710,N_10647);
or U10969 (N_10969,N_10629,N_10632);
nor U10970 (N_10970,N_10787,N_10701);
or U10971 (N_10971,N_10637,N_10795);
nand U10972 (N_10972,N_10672,N_10664);
or U10973 (N_10973,N_10722,N_10734);
and U10974 (N_10974,N_10615,N_10618);
nor U10975 (N_10975,N_10748,N_10659);
nor U10976 (N_10976,N_10757,N_10729);
or U10977 (N_10977,N_10695,N_10786);
and U10978 (N_10978,N_10658,N_10608);
nor U10979 (N_10979,N_10655,N_10741);
or U10980 (N_10980,N_10673,N_10737);
xnor U10981 (N_10981,N_10625,N_10742);
nor U10982 (N_10982,N_10600,N_10727);
or U10983 (N_10983,N_10722,N_10693);
xor U10984 (N_10984,N_10619,N_10785);
and U10985 (N_10985,N_10604,N_10779);
or U10986 (N_10986,N_10688,N_10727);
nor U10987 (N_10987,N_10688,N_10738);
or U10988 (N_10988,N_10661,N_10726);
and U10989 (N_10989,N_10662,N_10685);
nand U10990 (N_10990,N_10621,N_10733);
xnor U10991 (N_10991,N_10721,N_10722);
xor U10992 (N_10992,N_10783,N_10675);
or U10993 (N_10993,N_10701,N_10769);
nand U10994 (N_10994,N_10782,N_10779);
or U10995 (N_10995,N_10635,N_10755);
and U10996 (N_10996,N_10777,N_10789);
and U10997 (N_10997,N_10704,N_10745);
nor U10998 (N_10998,N_10730,N_10709);
nand U10999 (N_10999,N_10680,N_10738);
or U11000 (N_11000,N_10910,N_10813);
or U11001 (N_11001,N_10821,N_10810);
xnor U11002 (N_11002,N_10830,N_10927);
xor U11003 (N_11003,N_10890,N_10893);
or U11004 (N_11004,N_10994,N_10923);
or U11005 (N_11005,N_10820,N_10998);
or U11006 (N_11006,N_10997,N_10861);
nor U11007 (N_11007,N_10873,N_10804);
or U11008 (N_11008,N_10898,N_10843);
nor U11009 (N_11009,N_10960,N_10956);
xor U11010 (N_11010,N_10812,N_10881);
or U11011 (N_11011,N_10986,N_10906);
and U11012 (N_11012,N_10982,N_10918);
and U11013 (N_11013,N_10930,N_10967);
or U11014 (N_11014,N_10925,N_10825);
nor U11015 (N_11015,N_10844,N_10934);
or U11016 (N_11016,N_10985,N_10860);
or U11017 (N_11017,N_10884,N_10917);
or U11018 (N_11018,N_10837,N_10838);
nand U11019 (N_11019,N_10809,N_10903);
xnor U11020 (N_11020,N_10991,N_10950);
nand U11021 (N_11021,N_10892,N_10871);
nand U11022 (N_11022,N_10858,N_10990);
or U11023 (N_11023,N_10978,N_10851);
and U11024 (N_11024,N_10944,N_10977);
or U11025 (N_11025,N_10912,N_10822);
nor U11026 (N_11026,N_10931,N_10815);
or U11027 (N_11027,N_10849,N_10886);
nand U11028 (N_11028,N_10996,N_10993);
xor U11029 (N_11029,N_10942,N_10916);
and U11030 (N_11030,N_10801,N_10802);
or U11031 (N_11031,N_10966,N_10816);
nor U11032 (N_11032,N_10938,N_10952);
nand U11033 (N_11033,N_10839,N_10899);
xor U11034 (N_11034,N_10870,N_10932);
nor U11035 (N_11035,N_10852,N_10907);
and U11036 (N_11036,N_10829,N_10827);
or U11037 (N_11037,N_10808,N_10949);
nor U11038 (N_11038,N_10919,N_10875);
nand U11039 (N_11039,N_10921,N_10805);
xnor U11040 (N_11040,N_10963,N_10866);
or U11041 (N_11041,N_10885,N_10826);
xnor U11042 (N_11042,N_10882,N_10999);
nand U11043 (N_11043,N_10926,N_10976);
or U11044 (N_11044,N_10980,N_10846);
nand U11045 (N_11045,N_10811,N_10803);
nand U11046 (N_11046,N_10888,N_10833);
nor U11047 (N_11047,N_10902,N_10909);
nand U11048 (N_11048,N_10981,N_10989);
and U11049 (N_11049,N_10883,N_10862);
and U11050 (N_11050,N_10865,N_10937);
or U11051 (N_11051,N_10965,N_10962);
xor U11052 (N_11052,N_10891,N_10971);
or U11053 (N_11053,N_10834,N_10835);
nand U11054 (N_11054,N_10877,N_10841);
or U11055 (N_11055,N_10900,N_10988);
or U11056 (N_11056,N_10894,N_10880);
and U11057 (N_11057,N_10824,N_10823);
nand U11058 (N_11058,N_10868,N_10855);
and U11059 (N_11059,N_10992,N_10854);
xnor U11060 (N_11060,N_10897,N_10800);
nor U11061 (N_11061,N_10896,N_10817);
or U11062 (N_11062,N_10979,N_10943);
xor U11063 (N_11063,N_10878,N_10922);
and U11064 (N_11064,N_10818,N_10845);
nor U11065 (N_11065,N_10983,N_10941);
xor U11066 (N_11066,N_10972,N_10864);
nand U11067 (N_11067,N_10961,N_10975);
nand U11068 (N_11068,N_10876,N_10928);
or U11069 (N_11069,N_10969,N_10904);
xnor U11070 (N_11070,N_10895,N_10853);
nand U11071 (N_11071,N_10887,N_10819);
xor U11072 (N_11072,N_10933,N_10908);
and U11073 (N_11073,N_10832,N_10939);
nor U11074 (N_11074,N_10947,N_10920);
nor U11075 (N_11075,N_10955,N_10872);
nand U11076 (N_11076,N_10807,N_10879);
nor U11077 (N_11077,N_10954,N_10945);
xnor U11078 (N_11078,N_10848,N_10842);
or U11079 (N_11079,N_10957,N_10905);
nand U11080 (N_11080,N_10970,N_10959);
xor U11081 (N_11081,N_10857,N_10814);
and U11082 (N_11082,N_10914,N_10915);
nand U11083 (N_11083,N_10867,N_10847);
and U11084 (N_11084,N_10948,N_10987);
nor U11085 (N_11085,N_10935,N_10850);
nand U11086 (N_11086,N_10901,N_10968);
xnor U11087 (N_11087,N_10911,N_10836);
nand U11088 (N_11088,N_10940,N_10929);
and U11089 (N_11089,N_10924,N_10889);
or U11090 (N_11090,N_10840,N_10828);
and U11091 (N_11091,N_10856,N_10806);
nor U11092 (N_11092,N_10874,N_10913);
nand U11093 (N_11093,N_10973,N_10936);
and U11094 (N_11094,N_10995,N_10946);
and U11095 (N_11095,N_10951,N_10958);
nor U11096 (N_11096,N_10863,N_10984);
nor U11097 (N_11097,N_10869,N_10859);
nand U11098 (N_11098,N_10831,N_10953);
nand U11099 (N_11099,N_10974,N_10964);
and U11100 (N_11100,N_10965,N_10938);
nor U11101 (N_11101,N_10901,N_10998);
or U11102 (N_11102,N_10834,N_10958);
nor U11103 (N_11103,N_10967,N_10991);
and U11104 (N_11104,N_10979,N_10882);
nor U11105 (N_11105,N_10874,N_10818);
nand U11106 (N_11106,N_10905,N_10879);
and U11107 (N_11107,N_10871,N_10911);
nor U11108 (N_11108,N_10917,N_10906);
nor U11109 (N_11109,N_10921,N_10934);
nand U11110 (N_11110,N_10905,N_10864);
nand U11111 (N_11111,N_10905,N_10916);
nand U11112 (N_11112,N_10899,N_10989);
and U11113 (N_11113,N_10946,N_10955);
nor U11114 (N_11114,N_10934,N_10944);
and U11115 (N_11115,N_10885,N_10831);
or U11116 (N_11116,N_10893,N_10863);
nor U11117 (N_11117,N_10935,N_10828);
or U11118 (N_11118,N_10863,N_10938);
or U11119 (N_11119,N_10827,N_10938);
or U11120 (N_11120,N_10944,N_10930);
xnor U11121 (N_11121,N_10847,N_10921);
nand U11122 (N_11122,N_10883,N_10998);
xor U11123 (N_11123,N_10990,N_10955);
nand U11124 (N_11124,N_10904,N_10944);
nand U11125 (N_11125,N_10967,N_10852);
or U11126 (N_11126,N_10850,N_10827);
and U11127 (N_11127,N_10979,N_10840);
and U11128 (N_11128,N_10927,N_10835);
or U11129 (N_11129,N_10971,N_10899);
nor U11130 (N_11130,N_10939,N_10969);
xor U11131 (N_11131,N_10902,N_10854);
nor U11132 (N_11132,N_10844,N_10953);
nand U11133 (N_11133,N_10919,N_10977);
nand U11134 (N_11134,N_10932,N_10842);
or U11135 (N_11135,N_10836,N_10893);
xor U11136 (N_11136,N_10860,N_10871);
or U11137 (N_11137,N_10984,N_10850);
nand U11138 (N_11138,N_10906,N_10992);
or U11139 (N_11139,N_10886,N_10958);
and U11140 (N_11140,N_10938,N_10954);
xor U11141 (N_11141,N_10979,N_10868);
nor U11142 (N_11142,N_10964,N_10895);
nand U11143 (N_11143,N_10874,N_10801);
and U11144 (N_11144,N_10977,N_10841);
and U11145 (N_11145,N_10947,N_10979);
xor U11146 (N_11146,N_10962,N_10826);
xor U11147 (N_11147,N_10879,N_10840);
nor U11148 (N_11148,N_10999,N_10932);
nor U11149 (N_11149,N_10854,N_10917);
nor U11150 (N_11150,N_10926,N_10897);
or U11151 (N_11151,N_10881,N_10892);
or U11152 (N_11152,N_10959,N_10993);
or U11153 (N_11153,N_10832,N_10838);
and U11154 (N_11154,N_10816,N_10993);
nand U11155 (N_11155,N_10903,N_10843);
xnor U11156 (N_11156,N_10861,N_10839);
xor U11157 (N_11157,N_10999,N_10935);
or U11158 (N_11158,N_10837,N_10925);
and U11159 (N_11159,N_10833,N_10862);
or U11160 (N_11160,N_10997,N_10946);
nor U11161 (N_11161,N_10801,N_10902);
and U11162 (N_11162,N_10917,N_10843);
or U11163 (N_11163,N_10876,N_10917);
and U11164 (N_11164,N_10997,N_10969);
xor U11165 (N_11165,N_10968,N_10989);
and U11166 (N_11166,N_10808,N_10929);
or U11167 (N_11167,N_10904,N_10837);
or U11168 (N_11168,N_10815,N_10864);
and U11169 (N_11169,N_10920,N_10962);
and U11170 (N_11170,N_10921,N_10845);
nor U11171 (N_11171,N_10814,N_10892);
xnor U11172 (N_11172,N_10871,N_10833);
xor U11173 (N_11173,N_10886,N_10938);
and U11174 (N_11174,N_10866,N_10979);
or U11175 (N_11175,N_10932,N_10991);
nor U11176 (N_11176,N_10937,N_10815);
nor U11177 (N_11177,N_10883,N_10959);
and U11178 (N_11178,N_10969,N_10837);
nor U11179 (N_11179,N_10945,N_10951);
xor U11180 (N_11180,N_10969,N_10967);
nand U11181 (N_11181,N_10896,N_10814);
nor U11182 (N_11182,N_10895,N_10953);
or U11183 (N_11183,N_10994,N_10887);
nand U11184 (N_11184,N_10838,N_10805);
nand U11185 (N_11185,N_10936,N_10825);
nand U11186 (N_11186,N_10987,N_10868);
xnor U11187 (N_11187,N_10846,N_10945);
xnor U11188 (N_11188,N_10923,N_10858);
or U11189 (N_11189,N_10987,N_10889);
and U11190 (N_11190,N_10905,N_10906);
or U11191 (N_11191,N_10975,N_10900);
xnor U11192 (N_11192,N_10921,N_10851);
nor U11193 (N_11193,N_10822,N_10934);
and U11194 (N_11194,N_10986,N_10977);
or U11195 (N_11195,N_10902,N_10860);
xor U11196 (N_11196,N_10991,N_10866);
and U11197 (N_11197,N_10894,N_10810);
nor U11198 (N_11198,N_10842,N_10809);
nor U11199 (N_11199,N_10803,N_10960);
and U11200 (N_11200,N_11122,N_11042);
nand U11201 (N_11201,N_11162,N_11074);
xnor U11202 (N_11202,N_11168,N_11089);
or U11203 (N_11203,N_11081,N_11032);
or U11204 (N_11204,N_11060,N_11041);
and U11205 (N_11205,N_11038,N_11163);
and U11206 (N_11206,N_11183,N_11148);
xor U11207 (N_11207,N_11078,N_11124);
and U11208 (N_11208,N_11141,N_11109);
nor U11209 (N_11209,N_11145,N_11147);
or U11210 (N_11210,N_11154,N_11180);
nand U11211 (N_11211,N_11049,N_11054);
xnor U11212 (N_11212,N_11098,N_11050);
xnor U11213 (N_11213,N_11065,N_11146);
or U11214 (N_11214,N_11090,N_11169);
xnor U11215 (N_11215,N_11138,N_11048);
nor U11216 (N_11216,N_11184,N_11193);
or U11217 (N_11217,N_11111,N_11157);
and U11218 (N_11218,N_11057,N_11121);
nand U11219 (N_11219,N_11051,N_11113);
nand U11220 (N_11220,N_11129,N_11118);
nor U11221 (N_11221,N_11108,N_11080);
or U11222 (N_11222,N_11008,N_11178);
nor U11223 (N_11223,N_11039,N_11126);
nor U11224 (N_11224,N_11006,N_11059);
or U11225 (N_11225,N_11047,N_11067);
nand U11226 (N_11226,N_11190,N_11029);
nor U11227 (N_11227,N_11053,N_11114);
or U11228 (N_11228,N_11132,N_11037);
nor U11229 (N_11229,N_11196,N_11177);
or U11230 (N_11230,N_11088,N_11068);
or U11231 (N_11231,N_11024,N_11174);
and U11232 (N_11232,N_11061,N_11159);
nor U11233 (N_11233,N_11071,N_11179);
xor U11234 (N_11234,N_11131,N_11171);
or U11235 (N_11235,N_11079,N_11085);
or U11236 (N_11236,N_11160,N_11191);
nor U11237 (N_11237,N_11007,N_11073);
xor U11238 (N_11238,N_11117,N_11104);
or U11239 (N_11239,N_11064,N_11046);
xor U11240 (N_11240,N_11173,N_11086);
nor U11241 (N_11241,N_11103,N_11170);
nand U11242 (N_11242,N_11033,N_11014);
and U11243 (N_11243,N_11052,N_11130);
and U11244 (N_11244,N_11087,N_11189);
nor U11245 (N_11245,N_11077,N_11076);
and U11246 (N_11246,N_11015,N_11075);
xor U11247 (N_11247,N_11156,N_11022);
xnor U11248 (N_11248,N_11155,N_11101);
nor U11249 (N_11249,N_11153,N_11186);
nand U11250 (N_11250,N_11020,N_11062);
nand U11251 (N_11251,N_11019,N_11083);
and U11252 (N_11252,N_11112,N_11198);
xnor U11253 (N_11253,N_11181,N_11150);
nor U11254 (N_11254,N_11120,N_11166);
and U11255 (N_11255,N_11151,N_11093);
or U11256 (N_11256,N_11139,N_11110);
nand U11257 (N_11257,N_11031,N_11106);
nand U11258 (N_11258,N_11123,N_11009);
or U11259 (N_11259,N_11143,N_11188);
and U11260 (N_11260,N_11199,N_11070);
and U11261 (N_11261,N_11099,N_11058);
xnor U11262 (N_11262,N_11040,N_11107);
and U11263 (N_11263,N_11100,N_11197);
nand U11264 (N_11264,N_11152,N_11069);
xor U11265 (N_11265,N_11195,N_11045);
nand U11266 (N_11266,N_11096,N_11004);
xor U11267 (N_11267,N_11000,N_11094);
nand U11268 (N_11268,N_11115,N_11167);
nor U11269 (N_11269,N_11025,N_11063);
nand U11270 (N_11270,N_11149,N_11092);
and U11271 (N_11271,N_11140,N_11165);
or U11272 (N_11272,N_11119,N_11030);
nand U11273 (N_11273,N_11172,N_11185);
nand U11274 (N_11274,N_11017,N_11043);
nand U11275 (N_11275,N_11035,N_11161);
or U11276 (N_11276,N_11158,N_11005);
nand U11277 (N_11277,N_11036,N_11002);
xnor U11278 (N_11278,N_11026,N_11134);
and U11279 (N_11279,N_11137,N_11095);
xnor U11280 (N_11280,N_11082,N_11192);
nor U11281 (N_11281,N_11066,N_11133);
or U11282 (N_11282,N_11128,N_11044);
xnor U11283 (N_11283,N_11116,N_11135);
and U11284 (N_11284,N_11136,N_11016);
xor U11285 (N_11285,N_11011,N_11175);
nand U11286 (N_11286,N_11102,N_11164);
or U11287 (N_11287,N_11144,N_11125);
and U11288 (N_11288,N_11097,N_11072);
xor U11289 (N_11289,N_11003,N_11021);
or U11290 (N_11290,N_11127,N_11142);
nand U11291 (N_11291,N_11084,N_11187);
nor U11292 (N_11292,N_11018,N_11027);
xnor U11293 (N_11293,N_11176,N_11034);
and U11294 (N_11294,N_11013,N_11012);
or U11295 (N_11295,N_11105,N_11001);
or U11296 (N_11296,N_11055,N_11182);
or U11297 (N_11297,N_11091,N_11010);
nand U11298 (N_11298,N_11023,N_11056);
or U11299 (N_11299,N_11028,N_11194);
or U11300 (N_11300,N_11199,N_11086);
nor U11301 (N_11301,N_11104,N_11175);
xnor U11302 (N_11302,N_11007,N_11019);
and U11303 (N_11303,N_11084,N_11149);
xnor U11304 (N_11304,N_11186,N_11040);
xnor U11305 (N_11305,N_11016,N_11000);
and U11306 (N_11306,N_11080,N_11024);
xor U11307 (N_11307,N_11018,N_11067);
and U11308 (N_11308,N_11128,N_11122);
nand U11309 (N_11309,N_11025,N_11130);
nor U11310 (N_11310,N_11019,N_11119);
xor U11311 (N_11311,N_11021,N_11024);
nor U11312 (N_11312,N_11008,N_11034);
or U11313 (N_11313,N_11134,N_11043);
or U11314 (N_11314,N_11145,N_11175);
or U11315 (N_11315,N_11122,N_11079);
xnor U11316 (N_11316,N_11087,N_11117);
nand U11317 (N_11317,N_11092,N_11002);
nand U11318 (N_11318,N_11036,N_11148);
nor U11319 (N_11319,N_11088,N_11156);
xor U11320 (N_11320,N_11161,N_11104);
and U11321 (N_11321,N_11198,N_11027);
nand U11322 (N_11322,N_11037,N_11177);
nor U11323 (N_11323,N_11126,N_11046);
or U11324 (N_11324,N_11072,N_11176);
nand U11325 (N_11325,N_11007,N_11075);
nor U11326 (N_11326,N_11190,N_11094);
or U11327 (N_11327,N_11018,N_11166);
nor U11328 (N_11328,N_11130,N_11047);
nand U11329 (N_11329,N_11169,N_11199);
nand U11330 (N_11330,N_11026,N_11019);
xor U11331 (N_11331,N_11137,N_11066);
nand U11332 (N_11332,N_11186,N_11045);
and U11333 (N_11333,N_11153,N_11007);
xnor U11334 (N_11334,N_11133,N_11103);
nand U11335 (N_11335,N_11108,N_11130);
or U11336 (N_11336,N_11148,N_11020);
or U11337 (N_11337,N_11010,N_11100);
nand U11338 (N_11338,N_11017,N_11053);
nand U11339 (N_11339,N_11195,N_11176);
nor U11340 (N_11340,N_11008,N_11083);
nor U11341 (N_11341,N_11072,N_11135);
nand U11342 (N_11342,N_11195,N_11121);
or U11343 (N_11343,N_11184,N_11018);
nor U11344 (N_11344,N_11147,N_11051);
xor U11345 (N_11345,N_11053,N_11154);
nor U11346 (N_11346,N_11063,N_11097);
xor U11347 (N_11347,N_11052,N_11045);
or U11348 (N_11348,N_11068,N_11095);
nand U11349 (N_11349,N_11119,N_11045);
nand U11350 (N_11350,N_11156,N_11150);
nand U11351 (N_11351,N_11167,N_11044);
nor U11352 (N_11352,N_11181,N_11014);
xor U11353 (N_11353,N_11036,N_11068);
nor U11354 (N_11354,N_11103,N_11199);
nor U11355 (N_11355,N_11074,N_11133);
nor U11356 (N_11356,N_11062,N_11154);
nand U11357 (N_11357,N_11085,N_11001);
nor U11358 (N_11358,N_11097,N_11152);
and U11359 (N_11359,N_11198,N_11067);
nand U11360 (N_11360,N_11169,N_11189);
nand U11361 (N_11361,N_11042,N_11132);
xnor U11362 (N_11362,N_11099,N_11055);
nor U11363 (N_11363,N_11005,N_11054);
nor U11364 (N_11364,N_11014,N_11124);
xnor U11365 (N_11365,N_11088,N_11131);
nand U11366 (N_11366,N_11149,N_11117);
and U11367 (N_11367,N_11193,N_11175);
nor U11368 (N_11368,N_11126,N_11088);
and U11369 (N_11369,N_11076,N_11014);
and U11370 (N_11370,N_11101,N_11034);
or U11371 (N_11371,N_11157,N_11095);
nor U11372 (N_11372,N_11077,N_11184);
nor U11373 (N_11373,N_11098,N_11007);
and U11374 (N_11374,N_11090,N_11103);
nor U11375 (N_11375,N_11031,N_11083);
nand U11376 (N_11376,N_11054,N_11085);
or U11377 (N_11377,N_11013,N_11103);
or U11378 (N_11378,N_11079,N_11097);
nand U11379 (N_11379,N_11079,N_11048);
nor U11380 (N_11380,N_11077,N_11109);
and U11381 (N_11381,N_11025,N_11062);
xor U11382 (N_11382,N_11193,N_11154);
xor U11383 (N_11383,N_11076,N_11179);
nand U11384 (N_11384,N_11123,N_11032);
or U11385 (N_11385,N_11087,N_11069);
or U11386 (N_11386,N_11112,N_11064);
nor U11387 (N_11387,N_11039,N_11115);
or U11388 (N_11388,N_11077,N_11187);
or U11389 (N_11389,N_11007,N_11006);
nor U11390 (N_11390,N_11054,N_11146);
or U11391 (N_11391,N_11052,N_11113);
nand U11392 (N_11392,N_11173,N_11056);
nor U11393 (N_11393,N_11040,N_11005);
or U11394 (N_11394,N_11145,N_11130);
or U11395 (N_11395,N_11016,N_11092);
nor U11396 (N_11396,N_11117,N_11193);
or U11397 (N_11397,N_11133,N_11188);
or U11398 (N_11398,N_11080,N_11198);
xnor U11399 (N_11399,N_11041,N_11016);
nor U11400 (N_11400,N_11397,N_11231);
nand U11401 (N_11401,N_11334,N_11272);
and U11402 (N_11402,N_11376,N_11352);
or U11403 (N_11403,N_11227,N_11234);
nor U11404 (N_11404,N_11396,N_11359);
xor U11405 (N_11405,N_11384,N_11329);
nand U11406 (N_11406,N_11244,N_11220);
and U11407 (N_11407,N_11389,N_11293);
or U11408 (N_11408,N_11277,N_11282);
and U11409 (N_11409,N_11200,N_11321);
or U11410 (N_11410,N_11323,N_11288);
nand U11411 (N_11411,N_11203,N_11335);
xor U11412 (N_11412,N_11229,N_11266);
xnor U11413 (N_11413,N_11371,N_11320);
or U11414 (N_11414,N_11224,N_11363);
or U11415 (N_11415,N_11238,N_11305);
nand U11416 (N_11416,N_11211,N_11242);
and U11417 (N_11417,N_11348,N_11303);
nand U11418 (N_11418,N_11315,N_11361);
nand U11419 (N_11419,N_11215,N_11398);
and U11420 (N_11420,N_11258,N_11367);
and U11421 (N_11421,N_11331,N_11327);
or U11422 (N_11422,N_11252,N_11365);
or U11423 (N_11423,N_11373,N_11294);
or U11424 (N_11424,N_11391,N_11357);
nand U11425 (N_11425,N_11233,N_11217);
nor U11426 (N_11426,N_11353,N_11387);
and U11427 (N_11427,N_11390,N_11237);
xnor U11428 (N_11428,N_11333,N_11248);
nand U11429 (N_11429,N_11308,N_11222);
nand U11430 (N_11430,N_11374,N_11386);
nand U11431 (N_11431,N_11276,N_11311);
nor U11432 (N_11432,N_11296,N_11239);
or U11433 (N_11433,N_11351,N_11306);
nor U11434 (N_11434,N_11226,N_11241);
nor U11435 (N_11435,N_11360,N_11221);
xor U11436 (N_11436,N_11350,N_11301);
nor U11437 (N_11437,N_11219,N_11279);
xor U11438 (N_11438,N_11297,N_11206);
and U11439 (N_11439,N_11307,N_11265);
and U11440 (N_11440,N_11340,N_11326);
and U11441 (N_11441,N_11338,N_11364);
and U11442 (N_11442,N_11383,N_11328);
and U11443 (N_11443,N_11393,N_11349);
xor U11444 (N_11444,N_11332,N_11375);
and U11445 (N_11445,N_11264,N_11245);
and U11446 (N_11446,N_11314,N_11309);
nor U11447 (N_11447,N_11366,N_11204);
nor U11448 (N_11448,N_11287,N_11341);
or U11449 (N_11449,N_11310,N_11232);
or U11450 (N_11450,N_11300,N_11324);
or U11451 (N_11451,N_11262,N_11270);
and U11452 (N_11452,N_11322,N_11213);
nand U11453 (N_11453,N_11259,N_11261);
xnor U11454 (N_11454,N_11243,N_11380);
nor U11455 (N_11455,N_11370,N_11210);
xor U11456 (N_11456,N_11281,N_11236);
and U11457 (N_11457,N_11263,N_11369);
or U11458 (N_11458,N_11385,N_11269);
xor U11459 (N_11459,N_11207,N_11345);
nand U11460 (N_11460,N_11355,N_11325);
nand U11461 (N_11461,N_11368,N_11280);
nor U11462 (N_11462,N_11285,N_11223);
and U11463 (N_11463,N_11388,N_11377);
and U11464 (N_11464,N_11313,N_11399);
nor U11465 (N_11465,N_11249,N_11292);
or U11466 (N_11466,N_11208,N_11278);
xor U11467 (N_11467,N_11286,N_11275);
xor U11468 (N_11468,N_11358,N_11316);
and U11469 (N_11469,N_11283,N_11228);
nor U11470 (N_11470,N_11319,N_11235);
and U11471 (N_11471,N_11312,N_11336);
xor U11472 (N_11472,N_11284,N_11247);
or U11473 (N_11473,N_11212,N_11342);
and U11474 (N_11474,N_11347,N_11392);
nor U11475 (N_11475,N_11395,N_11225);
nor U11476 (N_11476,N_11382,N_11271);
and U11477 (N_11477,N_11250,N_11254);
or U11478 (N_11478,N_11230,N_11214);
nand U11479 (N_11479,N_11257,N_11291);
and U11480 (N_11480,N_11379,N_11216);
and U11481 (N_11481,N_11318,N_11381);
or U11482 (N_11482,N_11267,N_11201);
xnor U11483 (N_11483,N_11302,N_11330);
nor U11484 (N_11484,N_11202,N_11251);
and U11485 (N_11485,N_11295,N_11260);
or U11486 (N_11486,N_11304,N_11255);
nand U11487 (N_11487,N_11253,N_11372);
or U11488 (N_11488,N_11343,N_11290);
or U11489 (N_11489,N_11246,N_11378);
nand U11490 (N_11490,N_11256,N_11354);
and U11491 (N_11491,N_11289,N_11205);
nand U11492 (N_11492,N_11273,N_11218);
nor U11493 (N_11493,N_11346,N_11394);
or U11494 (N_11494,N_11209,N_11240);
nor U11495 (N_11495,N_11298,N_11344);
and U11496 (N_11496,N_11317,N_11339);
and U11497 (N_11497,N_11337,N_11362);
nor U11498 (N_11498,N_11274,N_11268);
nand U11499 (N_11499,N_11299,N_11356);
nor U11500 (N_11500,N_11364,N_11265);
nor U11501 (N_11501,N_11369,N_11299);
nand U11502 (N_11502,N_11212,N_11336);
nor U11503 (N_11503,N_11238,N_11352);
xnor U11504 (N_11504,N_11337,N_11225);
or U11505 (N_11505,N_11267,N_11308);
or U11506 (N_11506,N_11241,N_11397);
and U11507 (N_11507,N_11352,N_11298);
xnor U11508 (N_11508,N_11253,N_11302);
nor U11509 (N_11509,N_11241,N_11239);
xor U11510 (N_11510,N_11212,N_11256);
xor U11511 (N_11511,N_11218,N_11388);
xor U11512 (N_11512,N_11385,N_11312);
and U11513 (N_11513,N_11339,N_11262);
or U11514 (N_11514,N_11350,N_11360);
and U11515 (N_11515,N_11210,N_11238);
or U11516 (N_11516,N_11379,N_11386);
and U11517 (N_11517,N_11384,N_11311);
and U11518 (N_11518,N_11219,N_11316);
and U11519 (N_11519,N_11225,N_11223);
or U11520 (N_11520,N_11360,N_11306);
nor U11521 (N_11521,N_11360,N_11203);
xor U11522 (N_11522,N_11341,N_11211);
xor U11523 (N_11523,N_11289,N_11393);
or U11524 (N_11524,N_11385,N_11329);
nor U11525 (N_11525,N_11248,N_11266);
nand U11526 (N_11526,N_11356,N_11338);
and U11527 (N_11527,N_11334,N_11250);
xor U11528 (N_11528,N_11312,N_11307);
xor U11529 (N_11529,N_11309,N_11331);
or U11530 (N_11530,N_11381,N_11209);
nand U11531 (N_11531,N_11258,N_11224);
nand U11532 (N_11532,N_11316,N_11393);
and U11533 (N_11533,N_11283,N_11223);
and U11534 (N_11534,N_11277,N_11342);
or U11535 (N_11535,N_11383,N_11381);
or U11536 (N_11536,N_11265,N_11354);
xnor U11537 (N_11537,N_11358,N_11238);
nand U11538 (N_11538,N_11337,N_11234);
nand U11539 (N_11539,N_11371,N_11219);
nand U11540 (N_11540,N_11349,N_11341);
nor U11541 (N_11541,N_11310,N_11247);
or U11542 (N_11542,N_11245,N_11217);
nor U11543 (N_11543,N_11284,N_11306);
and U11544 (N_11544,N_11312,N_11213);
and U11545 (N_11545,N_11351,N_11282);
and U11546 (N_11546,N_11228,N_11297);
or U11547 (N_11547,N_11307,N_11206);
nand U11548 (N_11548,N_11214,N_11332);
or U11549 (N_11549,N_11267,N_11221);
xnor U11550 (N_11550,N_11240,N_11311);
nand U11551 (N_11551,N_11225,N_11387);
xnor U11552 (N_11552,N_11255,N_11218);
nand U11553 (N_11553,N_11206,N_11347);
nand U11554 (N_11554,N_11236,N_11277);
and U11555 (N_11555,N_11399,N_11255);
nand U11556 (N_11556,N_11380,N_11379);
and U11557 (N_11557,N_11356,N_11217);
nor U11558 (N_11558,N_11301,N_11334);
nand U11559 (N_11559,N_11383,N_11335);
nand U11560 (N_11560,N_11327,N_11357);
or U11561 (N_11561,N_11314,N_11255);
or U11562 (N_11562,N_11336,N_11241);
and U11563 (N_11563,N_11384,N_11383);
nor U11564 (N_11564,N_11274,N_11311);
xor U11565 (N_11565,N_11281,N_11352);
xnor U11566 (N_11566,N_11388,N_11259);
xor U11567 (N_11567,N_11383,N_11308);
nor U11568 (N_11568,N_11224,N_11207);
nand U11569 (N_11569,N_11261,N_11240);
and U11570 (N_11570,N_11353,N_11303);
and U11571 (N_11571,N_11282,N_11241);
nor U11572 (N_11572,N_11388,N_11290);
or U11573 (N_11573,N_11287,N_11315);
nor U11574 (N_11574,N_11217,N_11256);
nand U11575 (N_11575,N_11314,N_11229);
or U11576 (N_11576,N_11206,N_11310);
nor U11577 (N_11577,N_11218,N_11349);
or U11578 (N_11578,N_11237,N_11234);
nand U11579 (N_11579,N_11211,N_11284);
xnor U11580 (N_11580,N_11363,N_11368);
xnor U11581 (N_11581,N_11250,N_11289);
nand U11582 (N_11582,N_11291,N_11232);
nand U11583 (N_11583,N_11339,N_11383);
nand U11584 (N_11584,N_11233,N_11324);
nor U11585 (N_11585,N_11221,N_11209);
nor U11586 (N_11586,N_11283,N_11271);
or U11587 (N_11587,N_11359,N_11229);
xnor U11588 (N_11588,N_11317,N_11244);
and U11589 (N_11589,N_11285,N_11359);
or U11590 (N_11590,N_11267,N_11377);
xnor U11591 (N_11591,N_11368,N_11320);
xor U11592 (N_11592,N_11232,N_11264);
or U11593 (N_11593,N_11361,N_11236);
nand U11594 (N_11594,N_11271,N_11202);
and U11595 (N_11595,N_11205,N_11391);
nor U11596 (N_11596,N_11303,N_11352);
nand U11597 (N_11597,N_11354,N_11297);
nand U11598 (N_11598,N_11297,N_11258);
nand U11599 (N_11599,N_11340,N_11248);
or U11600 (N_11600,N_11496,N_11418);
or U11601 (N_11601,N_11474,N_11565);
xnor U11602 (N_11602,N_11514,N_11497);
and U11603 (N_11603,N_11573,N_11488);
and U11604 (N_11604,N_11542,N_11559);
xnor U11605 (N_11605,N_11508,N_11574);
nand U11606 (N_11606,N_11509,N_11447);
or U11607 (N_11607,N_11520,N_11417);
or U11608 (N_11608,N_11435,N_11554);
and U11609 (N_11609,N_11547,N_11470);
and U11610 (N_11610,N_11431,N_11584);
nor U11611 (N_11611,N_11410,N_11482);
nor U11612 (N_11612,N_11445,N_11458);
or U11613 (N_11613,N_11551,N_11558);
nor U11614 (N_11614,N_11515,N_11400);
nand U11615 (N_11615,N_11402,N_11427);
nand U11616 (N_11616,N_11484,N_11540);
nand U11617 (N_11617,N_11587,N_11500);
and U11618 (N_11618,N_11531,N_11543);
nand U11619 (N_11619,N_11529,N_11533);
xor U11620 (N_11620,N_11592,N_11564);
or U11621 (N_11621,N_11528,N_11442);
and U11622 (N_11622,N_11459,N_11495);
or U11623 (N_11623,N_11426,N_11538);
or U11624 (N_11624,N_11476,N_11589);
nand U11625 (N_11625,N_11582,N_11523);
and U11626 (N_11626,N_11440,N_11443);
and U11627 (N_11627,N_11594,N_11535);
xnor U11628 (N_11628,N_11408,N_11439);
nand U11629 (N_11629,N_11499,N_11463);
nor U11630 (N_11630,N_11469,N_11438);
xnor U11631 (N_11631,N_11461,N_11557);
and U11632 (N_11632,N_11599,N_11448);
and U11633 (N_11633,N_11422,N_11518);
or U11634 (N_11634,N_11598,N_11567);
xnor U11635 (N_11635,N_11583,N_11429);
nand U11636 (N_11636,N_11433,N_11492);
nor U11637 (N_11637,N_11591,N_11585);
xor U11638 (N_11638,N_11477,N_11552);
and U11639 (N_11639,N_11485,N_11483);
or U11640 (N_11640,N_11536,N_11539);
xnor U11641 (N_11641,N_11544,N_11446);
xor U11642 (N_11642,N_11479,N_11452);
xnor U11643 (N_11643,N_11546,N_11511);
and U11644 (N_11644,N_11512,N_11545);
xnor U11645 (N_11645,N_11489,N_11526);
nor U11646 (N_11646,N_11510,N_11401);
or U11647 (N_11647,N_11444,N_11471);
nand U11648 (N_11648,N_11527,N_11586);
nand U11649 (N_11649,N_11480,N_11541);
or U11650 (N_11650,N_11569,N_11490);
or U11651 (N_11651,N_11441,N_11454);
or U11652 (N_11652,N_11516,N_11424);
or U11653 (N_11653,N_11420,N_11414);
and U11654 (N_11654,N_11406,N_11428);
nand U11655 (N_11655,N_11421,N_11593);
or U11656 (N_11656,N_11416,N_11419);
and U11657 (N_11657,N_11505,N_11524);
nor U11658 (N_11658,N_11556,N_11522);
nor U11659 (N_11659,N_11525,N_11430);
nor U11660 (N_11660,N_11519,N_11596);
nand U11661 (N_11661,N_11534,N_11494);
xor U11662 (N_11662,N_11561,N_11578);
xnor U11663 (N_11663,N_11560,N_11481);
nor U11664 (N_11664,N_11464,N_11453);
nor U11665 (N_11665,N_11436,N_11403);
xor U11666 (N_11666,N_11507,N_11532);
or U11667 (N_11667,N_11577,N_11570);
nand U11668 (N_11668,N_11455,N_11575);
nor U11669 (N_11669,N_11576,N_11579);
xor U11670 (N_11670,N_11562,N_11450);
nor U11671 (N_11671,N_11491,N_11503);
nor U11672 (N_11672,N_11563,N_11595);
nor U11673 (N_11673,N_11456,N_11486);
or U11674 (N_11674,N_11457,N_11572);
nor U11675 (N_11675,N_11548,N_11404);
and U11676 (N_11676,N_11590,N_11537);
xor U11677 (N_11677,N_11415,N_11502);
xnor U11678 (N_11678,N_11478,N_11409);
and U11679 (N_11679,N_11405,N_11550);
or U11680 (N_11680,N_11501,N_11504);
nand U11681 (N_11681,N_11498,N_11449);
nand U11682 (N_11682,N_11521,N_11566);
nor U11683 (N_11683,N_11423,N_11467);
xor U11684 (N_11684,N_11506,N_11517);
and U11685 (N_11685,N_11468,N_11475);
and U11686 (N_11686,N_11412,N_11465);
or U11687 (N_11687,N_11581,N_11588);
xnor U11688 (N_11688,N_11472,N_11568);
nor U11689 (N_11689,N_11437,N_11411);
xor U11690 (N_11690,N_11462,N_11434);
nor U11691 (N_11691,N_11597,N_11413);
and U11692 (N_11692,N_11580,N_11493);
and U11693 (N_11693,N_11513,N_11451);
or U11694 (N_11694,N_11555,N_11571);
nand U11695 (N_11695,N_11473,N_11460);
nand U11696 (N_11696,N_11407,N_11432);
nor U11697 (N_11697,N_11553,N_11530);
and U11698 (N_11698,N_11487,N_11425);
xor U11699 (N_11699,N_11466,N_11549);
and U11700 (N_11700,N_11475,N_11410);
nor U11701 (N_11701,N_11421,N_11599);
nor U11702 (N_11702,N_11466,N_11488);
or U11703 (N_11703,N_11445,N_11426);
nand U11704 (N_11704,N_11574,N_11539);
xor U11705 (N_11705,N_11420,N_11464);
xnor U11706 (N_11706,N_11571,N_11497);
nand U11707 (N_11707,N_11527,N_11415);
nor U11708 (N_11708,N_11566,N_11501);
nand U11709 (N_11709,N_11462,N_11533);
or U11710 (N_11710,N_11587,N_11515);
and U11711 (N_11711,N_11517,N_11487);
xor U11712 (N_11712,N_11468,N_11474);
nor U11713 (N_11713,N_11466,N_11512);
and U11714 (N_11714,N_11585,N_11473);
and U11715 (N_11715,N_11538,N_11569);
and U11716 (N_11716,N_11425,N_11453);
nand U11717 (N_11717,N_11525,N_11551);
nor U11718 (N_11718,N_11596,N_11433);
nor U11719 (N_11719,N_11441,N_11464);
or U11720 (N_11720,N_11406,N_11529);
nor U11721 (N_11721,N_11457,N_11418);
xor U11722 (N_11722,N_11559,N_11503);
and U11723 (N_11723,N_11464,N_11542);
and U11724 (N_11724,N_11444,N_11578);
nand U11725 (N_11725,N_11457,N_11596);
or U11726 (N_11726,N_11546,N_11573);
nand U11727 (N_11727,N_11559,N_11535);
xor U11728 (N_11728,N_11427,N_11544);
nor U11729 (N_11729,N_11407,N_11546);
nor U11730 (N_11730,N_11463,N_11545);
and U11731 (N_11731,N_11416,N_11438);
or U11732 (N_11732,N_11471,N_11460);
xor U11733 (N_11733,N_11536,N_11513);
nor U11734 (N_11734,N_11431,N_11583);
nor U11735 (N_11735,N_11591,N_11455);
nor U11736 (N_11736,N_11478,N_11560);
or U11737 (N_11737,N_11445,N_11563);
or U11738 (N_11738,N_11581,N_11444);
or U11739 (N_11739,N_11509,N_11485);
xnor U11740 (N_11740,N_11487,N_11544);
xor U11741 (N_11741,N_11497,N_11414);
xor U11742 (N_11742,N_11488,N_11448);
nand U11743 (N_11743,N_11516,N_11431);
and U11744 (N_11744,N_11573,N_11424);
or U11745 (N_11745,N_11545,N_11419);
or U11746 (N_11746,N_11584,N_11543);
nor U11747 (N_11747,N_11456,N_11471);
nor U11748 (N_11748,N_11459,N_11453);
nor U11749 (N_11749,N_11447,N_11401);
xor U11750 (N_11750,N_11406,N_11409);
xor U11751 (N_11751,N_11480,N_11593);
or U11752 (N_11752,N_11453,N_11402);
xor U11753 (N_11753,N_11510,N_11454);
nor U11754 (N_11754,N_11556,N_11468);
or U11755 (N_11755,N_11494,N_11466);
nor U11756 (N_11756,N_11557,N_11428);
nor U11757 (N_11757,N_11489,N_11458);
xnor U11758 (N_11758,N_11431,N_11599);
and U11759 (N_11759,N_11590,N_11587);
xnor U11760 (N_11760,N_11453,N_11415);
nor U11761 (N_11761,N_11523,N_11488);
or U11762 (N_11762,N_11455,N_11596);
or U11763 (N_11763,N_11469,N_11509);
and U11764 (N_11764,N_11427,N_11573);
xor U11765 (N_11765,N_11401,N_11506);
nand U11766 (N_11766,N_11552,N_11410);
xnor U11767 (N_11767,N_11436,N_11482);
and U11768 (N_11768,N_11456,N_11424);
xor U11769 (N_11769,N_11450,N_11516);
nand U11770 (N_11770,N_11460,N_11463);
nor U11771 (N_11771,N_11465,N_11470);
and U11772 (N_11772,N_11480,N_11573);
xnor U11773 (N_11773,N_11466,N_11476);
nand U11774 (N_11774,N_11482,N_11542);
nand U11775 (N_11775,N_11422,N_11517);
xor U11776 (N_11776,N_11462,N_11584);
nand U11777 (N_11777,N_11481,N_11509);
nand U11778 (N_11778,N_11513,N_11573);
xnor U11779 (N_11779,N_11453,N_11519);
or U11780 (N_11780,N_11405,N_11404);
or U11781 (N_11781,N_11507,N_11430);
nor U11782 (N_11782,N_11584,N_11490);
nand U11783 (N_11783,N_11460,N_11494);
and U11784 (N_11784,N_11500,N_11440);
and U11785 (N_11785,N_11526,N_11486);
and U11786 (N_11786,N_11426,N_11508);
and U11787 (N_11787,N_11573,N_11539);
and U11788 (N_11788,N_11510,N_11555);
or U11789 (N_11789,N_11561,N_11564);
or U11790 (N_11790,N_11459,N_11545);
and U11791 (N_11791,N_11422,N_11567);
nor U11792 (N_11792,N_11502,N_11480);
xor U11793 (N_11793,N_11550,N_11469);
nor U11794 (N_11794,N_11512,N_11521);
and U11795 (N_11795,N_11481,N_11597);
xor U11796 (N_11796,N_11462,N_11544);
or U11797 (N_11797,N_11431,N_11408);
and U11798 (N_11798,N_11448,N_11494);
nor U11799 (N_11799,N_11417,N_11434);
nor U11800 (N_11800,N_11634,N_11668);
or U11801 (N_11801,N_11722,N_11730);
or U11802 (N_11802,N_11766,N_11797);
and U11803 (N_11803,N_11674,N_11620);
or U11804 (N_11804,N_11779,N_11669);
or U11805 (N_11805,N_11784,N_11778);
nand U11806 (N_11806,N_11792,N_11717);
or U11807 (N_11807,N_11738,N_11733);
nor U11808 (N_11808,N_11694,N_11764);
nand U11809 (N_11809,N_11752,N_11746);
or U11810 (N_11810,N_11613,N_11624);
xnor U11811 (N_11811,N_11719,N_11604);
nand U11812 (N_11812,N_11796,N_11704);
xor U11813 (N_11813,N_11737,N_11725);
or U11814 (N_11814,N_11711,N_11653);
xnor U11815 (N_11815,N_11633,N_11603);
xor U11816 (N_11816,N_11677,N_11697);
nor U11817 (N_11817,N_11756,N_11747);
and U11818 (N_11818,N_11724,N_11742);
and U11819 (N_11819,N_11696,N_11661);
xor U11820 (N_11820,N_11606,N_11729);
or U11821 (N_11821,N_11637,N_11642);
xor U11822 (N_11822,N_11767,N_11650);
xnor U11823 (N_11823,N_11675,N_11611);
xnor U11824 (N_11824,N_11723,N_11614);
and U11825 (N_11825,N_11617,N_11786);
xor U11826 (N_11826,N_11664,N_11726);
or U11827 (N_11827,N_11749,N_11732);
or U11828 (N_11828,N_11753,N_11718);
nor U11829 (N_11829,N_11710,N_11676);
nand U11830 (N_11830,N_11631,N_11644);
xor U11831 (N_11831,N_11689,N_11693);
and U11832 (N_11832,N_11640,N_11685);
or U11833 (N_11833,N_11657,N_11731);
nor U11834 (N_11834,N_11682,N_11795);
or U11835 (N_11835,N_11680,N_11673);
nand U11836 (N_11836,N_11759,N_11755);
nand U11837 (N_11837,N_11748,N_11788);
xor U11838 (N_11838,N_11616,N_11662);
nor U11839 (N_11839,N_11715,N_11625);
nand U11840 (N_11840,N_11769,N_11785);
nand U11841 (N_11841,N_11713,N_11622);
nand U11842 (N_11842,N_11745,N_11765);
and U11843 (N_11843,N_11774,N_11686);
xnor U11844 (N_11844,N_11720,N_11787);
nor U11845 (N_11845,N_11751,N_11762);
and U11846 (N_11846,N_11660,N_11708);
nand U11847 (N_11847,N_11651,N_11630);
and U11848 (N_11848,N_11670,N_11618);
nand U11849 (N_11849,N_11735,N_11702);
xor U11850 (N_11850,N_11703,N_11645);
xor U11851 (N_11851,N_11690,N_11798);
nor U11852 (N_11852,N_11684,N_11705);
or U11853 (N_11853,N_11727,N_11679);
or U11854 (N_11854,N_11609,N_11760);
and U11855 (N_11855,N_11707,N_11646);
nand U11856 (N_11856,N_11655,N_11750);
nand U11857 (N_11857,N_11687,N_11627);
or U11858 (N_11858,N_11605,N_11615);
xor U11859 (N_11859,N_11681,N_11799);
or U11860 (N_11860,N_11648,N_11728);
nand U11861 (N_11861,N_11643,N_11761);
and U11862 (N_11862,N_11772,N_11656);
nor U11863 (N_11863,N_11639,N_11663);
xnor U11864 (N_11864,N_11626,N_11744);
or U11865 (N_11865,N_11698,N_11619);
or U11866 (N_11866,N_11736,N_11775);
or U11867 (N_11867,N_11629,N_11781);
or U11868 (N_11868,N_11768,N_11601);
or U11869 (N_11869,N_11665,N_11741);
or U11870 (N_11870,N_11659,N_11699);
or U11871 (N_11871,N_11773,N_11740);
xor U11872 (N_11872,N_11636,N_11793);
nor U11873 (N_11873,N_11712,N_11638);
nor U11874 (N_11874,N_11734,N_11654);
or U11875 (N_11875,N_11612,N_11754);
xor U11876 (N_11876,N_11794,N_11692);
nor U11877 (N_11877,N_11623,N_11666);
nand U11878 (N_11878,N_11780,N_11678);
xor U11879 (N_11879,N_11671,N_11658);
or U11880 (N_11880,N_11701,N_11641);
nand U11881 (N_11881,N_11610,N_11683);
or U11882 (N_11882,N_11714,N_11791);
nand U11883 (N_11883,N_11652,N_11672);
nor U11884 (N_11884,N_11743,N_11770);
or U11885 (N_11885,N_11782,N_11700);
and U11886 (N_11886,N_11757,N_11789);
xnor U11887 (N_11887,N_11649,N_11709);
and U11888 (N_11888,N_11608,N_11632);
nand U11889 (N_11889,N_11635,N_11695);
xnor U11890 (N_11890,N_11721,N_11739);
and U11891 (N_11891,N_11771,N_11776);
xnor U11892 (N_11892,N_11688,N_11758);
nor U11893 (N_11893,N_11706,N_11607);
nand U11894 (N_11894,N_11716,N_11691);
nand U11895 (N_11895,N_11667,N_11602);
xnor U11896 (N_11896,N_11647,N_11621);
and U11897 (N_11897,N_11777,N_11628);
nor U11898 (N_11898,N_11600,N_11763);
nor U11899 (N_11899,N_11790,N_11783);
nand U11900 (N_11900,N_11712,N_11605);
or U11901 (N_11901,N_11750,N_11664);
and U11902 (N_11902,N_11683,N_11682);
nor U11903 (N_11903,N_11621,N_11659);
nor U11904 (N_11904,N_11718,N_11601);
nor U11905 (N_11905,N_11726,N_11747);
or U11906 (N_11906,N_11692,N_11738);
nor U11907 (N_11907,N_11606,N_11678);
nor U11908 (N_11908,N_11693,N_11641);
and U11909 (N_11909,N_11720,N_11750);
and U11910 (N_11910,N_11768,N_11747);
or U11911 (N_11911,N_11663,N_11626);
or U11912 (N_11912,N_11631,N_11747);
nor U11913 (N_11913,N_11646,N_11621);
xnor U11914 (N_11914,N_11735,N_11671);
or U11915 (N_11915,N_11654,N_11640);
or U11916 (N_11916,N_11764,N_11704);
or U11917 (N_11917,N_11602,N_11775);
and U11918 (N_11918,N_11799,N_11739);
xnor U11919 (N_11919,N_11730,N_11712);
nand U11920 (N_11920,N_11751,N_11649);
nand U11921 (N_11921,N_11664,N_11712);
and U11922 (N_11922,N_11623,N_11787);
xor U11923 (N_11923,N_11715,N_11790);
nor U11924 (N_11924,N_11646,N_11687);
nor U11925 (N_11925,N_11706,N_11742);
or U11926 (N_11926,N_11771,N_11600);
nor U11927 (N_11927,N_11602,N_11687);
or U11928 (N_11928,N_11716,N_11718);
and U11929 (N_11929,N_11639,N_11694);
and U11930 (N_11930,N_11656,N_11650);
and U11931 (N_11931,N_11769,N_11735);
or U11932 (N_11932,N_11685,N_11681);
or U11933 (N_11933,N_11761,N_11741);
nor U11934 (N_11934,N_11795,N_11711);
and U11935 (N_11935,N_11762,N_11642);
xnor U11936 (N_11936,N_11713,N_11641);
xnor U11937 (N_11937,N_11770,N_11740);
nor U11938 (N_11938,N_11654,N_11792);
or U11939 (N_11939,N_11716,N_11614);
or U11940 (N_11940,N_11768,N_11663);
xor U11941 (N_11941,N_11635,N_11683);
nand U11942 (N_11942,N_11613,N_11610);
nor U11943 (N_11943,N_11606,N_11649);
nand U11944 (N_11944,N_11779,N_11730);
nor U11945 (N_11945,N_11652,N_11766);
and U11946 (N_11946,N_11614,N_11629);
nor U11947 (N_11947,N_11679,N_11648);
or U11948 (N_11948,N_11743,N_11695);
nand U11949 (N_11949,N_11612,N_11636);
nand U11950 (N_11950,N_11649,N_11613);
nand U11951 (N_11951,N_11794,N_11622);
nor U11952 (N_11952,N_11644,N_11702);
nor U11953 (N_11953,N_11635,N_11647);
and U11954 (N_11954,N_11677,N_11657);
nand U11955 (N_11955,N_11656,N_11734);
and U11956 (N_11956,N_11717,N_11708);
nor U11957 (N_11957,N_11663,N_11615);
nor U11958 (N_11958,N_11798,N_11672);
and U11959 (N_11959,N_11791,N_11741);
nor U11960 (N_11960,N_11635,N_11617);
and U11961 (N_11961,N_11645,N_11704);
and U11962 (N_11962,N_11618,N_11757);
xor U11963 (N_11963,N_11799,N_11771);
nor U11964 (N_11964,N_11627,N_11744);
or U11965 (N_11965,N_11687,N_11651);
or U11966 (N_11966,N_11620,N_11613);
nand U11967 (N_11967,N_11694,N_11666);
and U11968 (N_11968,N_11738,N_11735);
or U11969 (N_11969,N_11710,N_11788);
nand U11970 (N_11970,N_11735,N_11618);
nor U11971 (N_11971,N_11656,N_11713);
nor U11972 (N_11972,N_11786,N_11722);
nor U11973 (N_11973,N_11798,N_11768);
nand U11974 (N_11974,N_11633,N_11777);
and U11975 (N_11975,N_11698,N_11679);
nor U11976 (N_11976,N_11741,N_11725);
nor U11977 (N_11977,N_11693,N_11622);
xor U11978 (N_11978,N_11664,N_11683);
nor U11979 (N_11979,N_11799,N_11668);
nor U11980 (N_11980,N_11616,N_11785);
nor U11981 (N_11981,N_11620,N_11700);
nand U11982 (N_11982,N_11780,N_11663);
nand U11983 (N_11983,N_11612,N_11630);
nor U11984 (N_11984,N_11778,N_11666);
nand U11985 (N_11985,N_11736,N_11657);
or U11986 (N_11986,N_11611,N_11628);
xnor U11987 (N_11987,N_11662,N_11698);
and U11988 (N_11988,N_11649,N_11686);
nor U11989 (N_11989,N_11686,N_11788);
nand U11990 (N_11990,N_11649,N_11703);
nand U11991 (N_11991,N_11613,N_11733);
xnor U11992 (N_11992,N_11625,N_11689);
or U11993 (N_11993,N_11723,N_11655);
nand U11994 (N_11994,N_11786,N_11798);
nand U11995 (N_11995,N_11752,N_11761);
xor U11996 (N_11996,N_11648,N_11770);
nand U11997 (N_11997,N_11645,N_11665);
and U11998 (N_11998,N_11603,N_11709);
nor U11999 (N_11999,N_11671,N_11646);
nand U12000 (N_12000,N_11884,N_11853);
nor U12001 (N_12001,N_11813,N_11972);
and U12002 (N_12002,N_11838,N_11941);
or U12003 (N_12003,N_11800,N_11849);
nand U12004 (N_12004,N_11866,N_11848);
and U12005 (N_12005,N_11876,N_11870);
nor U12006 (N_12006,N_11911,N_11913);
nor U12007 (N_12007,N_11820,N_11825);
xor U12008 (N_12008,N_11917,N_11852);
nor U12009 (N_12009,N_11802,N_11973);
nor U12010 (N_12010,N_11915,N_11827);
nor U12011 (N_12011,N_11992,N_11997);
xor U12012 (N_12012,N_11879,N_11961);
or U12013 (N_12013,N_11830,N_11841);
or U12014 (N_12014,N_11880,N_11981);
or U12015 (N_12015,N_11909,N_11847);
xor U12016 (N_12016,N_11971,N_11975);
and U12017 (N_12017,N_11896,N_11988);
and U12018 (N_12018,N_11935,N_11956);
nand U12019 (N_12019,N_11931,N_11989);
or U12020 (N_12020,N_11892,N_11860);
xnor U12021 (N_12021,N_11927,N_11906);
nand U12022 (N_12022,N_11871,N_11952);
xnor U12023 (N_12023,N_11899,N_11829);
xor U12024 (N_12024,N_11861,N_11891);
nor U12025 (N_12025,N_11869,N_11976);
nand U12026 (N_12026,N_11995,N_11882);
xor U12027 (N_12027,N_11805,N_11816);
nand U12028 (N_12028,N_11863,N_11819);
nor U12029 (N_12029,N_11812,N_11960);
nand U12030 (N_12030,N_11977,N_11859);
or U12031 (N_12031,N_11902,N_11910);
xor U12032 (N_12032,N_11814,N_11945);
nor U12033 (N_12033,N_11803,N_11983);
and U12034 (N_12034,N_11929,N_11883);
nand U12035 (N_12035,N_11986,N_11926);
or U12036 (N_12036,N_11806,N_11933);
nand U12037 (N_12037,N_11950,N_11949);
or U12038 (N_12038,N_11923,N_11900);
and U12039 (N_12039,N_11834,N_11856);
and U12040 (N_12040,N_11990,N_11804);
nand U12041 (N_12041,N_11938,N_11835);
xnor U12042 (N_12042,N_11984,N_11937);
or U12043 (N_12043,N_11998,N_11842);
nor U12044 (N_12044,N_11948,N_11874);
nand U12045 (N_12045,N_11897,N_11886);
or U12046 (N_12046,N_11831,N_11940);
nor U12047 (N_12047,N_11914,N_11822);
xor U12048 (N_12048,N_11969,N_11947);
nand U12049 (N_12049,N_11817,N_11895);
nor U12050 (N_12050,N_11979,N_11888);
nor U12051 (N_12051,N_11936,N_11894);
and U12052 (N_12052,N_11890,N_11836);
or U12053 (N_12053,N_11964,N_11924);
or U12054 (N_12054,N_11832,N_11957);
and U12055 (N_12055,N_11922,N_11996);
xnor U12056 (N_12056,N_11875,N_11908);
or U12057 (N_12057,N_11942,N_11864);
and U12058 (N_12058,N_11865,N_11881);
or U12059 (N_12059,N_11967,N_11999);
nor U12060 (N_12060,N_11867,N_11928);
and U12061 (N_12061,N_11982,N_11809);
and U12062 (N_12062,N_11858,N_11919);
or U12063 (N_12063,N_11843,N_11953);
nand U12064 (N_12064,N_11925,N_11833);
nor U12065 (N_12065,N_11965,N_11893);
nand U12066 (N_12066,N_11962,N_11846);
xor U12067 (N_12067,N_11815,N_11966);
and U12068 (N_12068,N_11872,N_11857);
nand U12069 (N_12069,N_11921,N_11974);
nor U12070 (N_12070,N_11807,N_11920);
or U12071 (N_12071,N_11844,N_11934);
or U12072 (N_12072,N_11885,N_11845);
and U12073 (N_12073,N_11877,N_11887);
and U12074 (N_12074,N_11963,N_11932);
nor U12075 (N_12075,N_11978,N_11912);
xnor U12076 (N_12076,N_11823,N_11901);
nor U12077 (N_12077,N_11905,N_11801);
or U12078 (N_12078,N_11980,N_11955);
and U12079 (N_12079,N_11918,N_11868);
and U12080 (N_12080,N_11951,N_11855);
nand U12081 (N_12081,N_11946,N_11811);
xnor U12082 (N_12082,N_11878,N_11821);
nor U12083 (N_12083,N_11898,N_11907);
xnor U12084 (N_12084,N_11828,N_11808);
nand U12085 (N_12085,N_11824,N_11854);
xor U12086 (N_12086,N_11959,N_11818);
nand U12087 (N_12087,N_11954,N_11944);
nand U12088 (N_12088,N_11994,N_11939);
and U12089 (N_12089,N_11916,N_11991);
and U12090 (N_12090,N_11810,N_11889);
xnor U12091 (N_12091,N_11840,N_11943);
or U12092 (N_12092,N_11826,N_11970);
xnor U12093 (N_12093,N_11993,N_11850);
and U12094 (N_12094,N_11930,N_11873);
nand U12095 (N_12095,N_11851,N_11985);
nor U12096 (N_12096,N_11987,N_11862);
xor U12097 (N_12097,N_11958,N_11903);
or U12098 (N_12098,N_11968,N_11839);
or U12099 (N_12099,N_11904,N_11837);
nand U12100 (N_12100,N_11844,N_11886);
nand U12101 (N_12101,N_11874,N_11805);
nor U12102 (N_12102,N_11851,N_11897);
nand U12103 (N_12103,N_11903,N_11963);
xor U12104 (N_12104,N_11882,N_11806);
nor U12105 (N_12105,N_11951,N_11814);
or U12106 (N_12106,N_11907,N_11838);
or U12107 (N_12107,N_11960,N_11908);
nor U12108 (N_12108,N_11894,N_11899);
nand U12109 (N_12109,N_11896,N_11827);
nor U12110 (N_12110,N_11910,N_11911);
nor U12111 (N_12111,N_11817,N_11890);
nand U12112 (N_12112,N_11865,N_11812);
nor U12113 (N_12113,N_11809,N_11918);
nand U12114 (N_12114,N_11820,N_11810);
and U12115 (N_12115,N_11940,N_11888);
nor U12116 (N_12116,N_11920,N_11959);
nor U12117 (N_12117,N_11984,N_11902);
nor U12118 (N_12118,N_11914,N_11841);
or U12119 (N_12119,N_11897,N_11927);
or U12120 (N_12120,N_11946,N_11864);
nor U12121 (N_12121,N_11860,N_11842);
and U12122 (N_12122,N_11890,N_11857);
or U12123 (N_12123,N_11914,N_11866);
and U12124 (N_12124,N_11871,N_11910);
and U12125 (N_12125,N_11985,N_11997);
and U12126 (N_12126,N_11943,N_11948);
xor U12127 (N_12127,N_11990,N_11860);
and U12128 (N_12128,N_11917,N_11925);
nor U12129 (N_12129,N_11829,N_11954);
nand U12130 (N_12130,N_11989,N_11847);
xor U12131 (N_12131,N_11846,N_11919);
nand U12132 (N_12132,N_11922,N_11816);
nand U12133 (N_12133,N_11815,N_11949);
nor U12134 (N_12134,N_11966,N_11839);
nand U12135 (N_12135,N_11975,N_11890);
or U12136 (N_12136,N_11840,N_11972);
nand U12137 (N_12137,N_11970,N_11945);
and U12138 (N_12138,N_11983,N_11945);
and U12139 (N_12139,N_11817,N_11876);
nand U12140 (N_12140,N_11871,N_11839);
nand U12141 (N_12141,N_11854,N_11840);
nand U12142 (N_12142,N_11954,N_11809);
nand U12143 (N_12143,N_11887,N_11953);
or U12144 (N_12144,N_11970,N_11815);
and U12145 (N_12145,N_11953,N_11942);
or U12146 (N_12146,N_11894,N_11848);
xor U12147 (N_12147,N_11802,N_11917);
or U12148 (N_12148,N_11815,N_11845);
and U12149 (N_12149,N_11887,N_11902);
xnor U12150 (N_12150,N_11828,N_11998);
nand U12151 (N_12151,N_11856,N_11989);
xnor U12152 (N_12152,N_11948,N_11891);
nor U12153 (N_12153,N_11849,N_11931);
and U12154 (N_12154,N_11801,N_11981);
nor U12155 (N_12155,N_11950,N_11823);
xor U12156 (N_12156,N_11840,N_11968);
xor U12157 (N_12157,N_11823,N_11919);
nand U12158 (N_12158,N_11947,N_11994);
nand U12159 (N_12159,N_11928,N_11915);
and U12160 (N_12160,N_11981,N_11865);
and U12161 (N_12161,N_11926,N_11830);
nor U12162 (N_12162,N_11844,N_11978);
nor U12163 (N_12163,N_11913,N_11815);
nand U12164 (N_12164,N_11807,N_11906);
nand U12165 (N_12165,N_11960,N_11846);
xnor U12166 (N_12166,N_11964,N_11910);
nand U12167 (N_12167,N_11955,N_11928);
nand U12168 (N_12168,N_11931,N_11948);
nor U12169 (N_12169,N_11903,N_11876);
and U12170 (N_12170,N_11847,N_11873);
or U12171 (N_12171,N_11997,N_11962);
nor U12172 (N_12172,N_11991,N_11883);
and U12173 (N_12173,N_11899,N_11919);
xor U12174 (N_12174,N_11819,N_11916);
and U12175 (N_12175,N_11823,N_11825);
or U12176 (N_12176,N_11807,N_11888);
or U12177 (N_12177,N_11831,N_11970);
nor U12178 (N_12178,N_11905,N_11982);
nand U12179 (N_12179,N_11987,N_11990);
or U12180 (N_12180,N_11932,N_11953);
nand U12181 (N_12181,N_11879,N_11930);
and U12182 (N_12182,N_11995,N_11879);
xnor U12183 (N_12183,N_11887,N_11815);
xnor U12184 (N_12184,N_11851,N_11946);
or U12185 (N_12185,N_11840,N_11984);
nand U12186 (N_12186,N_11880,N_11846);
xnor U12187 (N_12187,N_11877,N_11981);
or U12188 (N_12188,N_11908,N_11810);
and U12189 (N_12189,N_11934,N_11892);
nand U12190 (N_12190,N_11882,N_11896);
nor U12191 (N_12191,N_11902,N_11826);
nor U12192 (N_12192,N_11858,N_11864);
nor U12193 (N_12193,N_11976,N_11922);
nand U12194 (N_12194,N_11948,N_11830);
or U12195 (N_12195,N_11920,N_11952);
xnor U12196 (N_12196,N_11963,N_11883);
or U12197 (N_12197,N_11933,N_11935);
nor U12198 (N_12198,N_11904,N_11966);
nand U12199 (N_12199,N_11920,N_11893);
nor U12200 (N_12200,N_12136,N_12104);
or U12201 (N_12201,N_12096,N_12081);
and U12202 (N_12202,N_12109,N_12032);
and U12203 (N_12203,N_12196,N_12190);
xor U12204 (N_12204,N_12059,N_12174);
and U12205 (N_12205,N_12095,N_12045);
nand U12206 (N_12206,N_12108,N_12089);
nand U12207 (N_12207,N_12145,N_12103);
nor U12208 (N_12208,N_12031,N_12087);
or U12209 (N_12209,N_12036,N_12038);
or U12210 (N_12210,N_12053,N_12051);
or U12211 (N_12211,N_12181,N_12193);
nor U12212 (N_12212,N_12184,N_12101);
and U12213 (N_12213,N_12026,N_12017);
nor U12214 (N_12214,N_12061,N_12188);
nor U12215 (N_12215,N_12154,N_12177);
or U12216 (N_12216,N_12117,N_12100);
nand U12217 (N_12217,N_12033,N_12025);
and U12218 (N_12218,N_12069,N_12010);
nand U12219 (N_12219,N_12133,N_12137);
and U12220 (N_12220,N_12163,N_12146);
xnor U12221 (N_12221,N_12028,N_12044);
xor U12222 (N_12222,N_12191,N_12124);
or U12223 (N_12223,N_12007,N_12122);
and U12224 (N_12224,N_12116,N_12167);
or U12225 (N_12225,N_12049,N_12016);
or U12226 (N_12226,N_12097,N_12077);
nand U12227 (N_12227,N_12186,N_12004);
nand U12228 (N_12228,N_12121,N_12119);
or U12229 (N_12229,N_12132,N_12060);
nor U12230 (N_12230,N_12135,N_12088);
xnor U12231 (N_12231,N_12005,N_12080);
and U12232 (N_12232,N_12166,N_12083);
nor U12233 (N_12233,N_12029,N_12009);
nand U12234 (N_12234,N_12098,N_12012);
and U12235 (N_12235,N_12041,N_12013);
and U12236 (N_12236,N_12195,N_12185);
nand U12237 (N_12237,N_12157,N_12047);
or U12238 (N_12238,N_12140,N_12072);
nand U12239 (N_12239,N_12042,N_12054);
nand U12240 (N_12240,N_12134,N_12147);
and U12241 (N_12241,N_12006,N_12015);
and U12242 (N_12242,N_12023,N_12086);
and U12243 (N_12243,N_12148,N_12156);
or U12244 (N_12244,N_12114,N_12065);
or U12245 (N_12245,N_12192,N_12102);
or U12246 (N_12246,N_12161,N_12068);
nor U12247 (N_12247,N_12175,N_12112);
or U12248 (N_12248,N_12180,N_12058);
nor U12249 (N_12249,N_12000,N_12173);
or U12250 (N_12250,N_12050,N_12057);
nand U12251 (N_12251,N_12062,N_12123);
and U12252 (N_12252,N_12037,N_12090);
or U12253 (N_12253,N_12118,N_12091);
nand U12254 (N_12254,N_12008,N_12022);
xnor U12255 (N_12255,N_12046,N_12106);
and U12256 (N_12256,N_12170,N_12011);
nand U12257 (N_12257,N_12143,N_12189);
or U12258 (N_12258,N_12152,N_12043);
nor U12259 (N_12259,N_12092,N_12130);
and U12260 (N_12260,N_12052,N_12099);
nand U12261 (N_12261,N_12162,N_12021);
nand U12262 (N_12262,N_12027,N_12018);
and U12263 (N_12263,N_12056,N_12076);
xor U12264 (N_12264,N_12153,N_12197);
nand U12265 (N_12265,N_12107,N_12070);
xor U12266 (N_12266,N_12149,N_12158);
xnor U12267 (N_12267,N_12194,N_12078);
nand U12268 (N_12268,N_12111,N_12071);
or U12269 (N_12269,N_12066,N_12179);
and U12270 (N_12270,N_12084,N_12129);
nand U12271 (N_12271,N_12079,N_12126);
xnor U12272 (N_12272,N_12125,N_12142);
and U12273 (N_12273,N_12055,N_12183);
xor U12274 (N_12274,N_12105,N_12082);
and U12275 (N_12275,N_12030,N_12172);
nor U12276 (N_12276,N_12113,N_12128);
nand U12277 (N_12277,N_12198,N_12003);
and U12278 (N_12278,N_12073,N_12160);
or U12279 (N_12279,N_12064,N_12176);
xor U12280 (N_12280,N_12131,N_12164);
nor U12281 (N_12281,N_12063,N_12035);
nand U12282 (N_12282,N_12139,N_12085);
nor U12283 (N_12283,N_12110,N_12002);
nand U12284 (N_12284,N_12074,N_12020);
nor U12285 (N_12285,N_12155,N_12094);
nand U12286 (N_12286,N_12138,N_12014);
xor U12287 (N_12287,N_12151,N_12019);
nand U12288 (N_12288,N_12168,N_12039);
and U12289 (N_12289,N_12187,N_12075);
nor U12290 (N_12290,N_12127,N_12024);
and U12291 (N_12291,N_12034,N_12182);
nor U12292 (N_12292,N_12169,N_12093);
nor U12293 (N_12293,N_12144,N_12001);
nand U12294 (N_12294,N_12141,N_12048);
or U12295 (N_12295,N_12040,N_12115);
nor U12296 (N_12296,N_12067,N_12178);
and U12297 (N_12297,N_12171,N_12120);
nand U12298 (N_12298,N_12159,N_12199);
and U12299 (N_12299,N_12165,N_12150);
nor U12300 (N_12300,N_12070,N_12128);
nor U12301 (N_12301,N_12187,N_12029);
and U12302 (N_12302,N_12002,N_12025);
or U12303 (N_12303,N_12042,N_12107);
and U12304 (N_12304,N_12143,N_12132);
or U12305 (N_12305,N_12164,N_12000);
xor U12306 (N_12306,N_12091,N_12111);
xor U12307 (N_12307,N_12149,N_12141);
and U12308 (N_12308,N_12134,N_12172);
nand U12309 (N_12309,N_12018,N_12010);
nor U12310 (N_12310,N_12118,N_12135);
or U12311 (N_12311,N_12076,N_12052);
and U12312 (N_12312,N_12065,N_12130);
xor U12313 (N_12313,N_12083,N_12175);
xor U12314 (N_12314,N_12187,N_12106);
nand U12315 (N_12315,N_12037,N_12157);
nand U12316 (N_12316,N_12184,N_12051);
and U12317 (N_12317,N_12127,N_12066);
xor U12318 (N_12318,N_12007,N_12023);
nor U12319 (N_12319,N_12013,N_12199);
or U12320 (N_12320,N_12088,N_12114);
xnor U12321 (N_12321,N_12175,N_12178);
xnor U12322 (N_12322,N_12039,N_12085);
nor U12323 (N_12323,N_12133,N_12061);
and U12324 (N_12324,N_12023,N_12012);
nor U12325 (N_12325,N_12067,N_12164);
nor U12326 (N_12326,N_12153,N_12111);
nand U12327 (N_12327,N_12021,N_12086);
nand U12328 (N_12328,N_12096,N_12122);
nand U12329 (N_12329,N_12114,N_12085);
or U12330 (N_12330,N_12013,N_12162);
or U12331 (N_12331,N_12019,N_12030);
xor U12332 (N_12332,N_12094,N_12187);
or U12333 (N_12333,N_12145,N_12031);
or U12334 (N_12334,N_12175,N_12126);
nand U12335 (N_12335,N_12143,N_12134);
nand U12336 (N_12336,N_12029,N_12083);
or U12337 (N_12337,N_12045,N_12000);
xnor U12338 (N_12338,N_12063,N_12111);
xor U12339 (N_12339,N_12189,N_12043);
nor U12340 (N_12340,N_12118,N_12085);
xor U12341 (N_12341,N_12113,N_12083);
or U12342 (N_12342,N_12145,N_12117);
nand U12343 (N_12343,N_12089,N_12195);
and U12344 (N_12344,N_12182,N_12031);
nand U12345 (N_12345,N_12015,N_12106);
nand U12346 (N_12346,N_12148,N_12072);
nor U12347 (N_12347,N_12119,N_12010);
nor U12348 (N_12348,N_12159,N_12176);
nand U12349 (N_12349,N_12134,N_12079);
or U12350 (N_12350,N_12089,N_12117);
and U12351 (N_12351,N_12022,N_12096);
xnor U12352 (N_12352,N_12068,N_12140);
nor U12353 (N_12353,N_12186,N_12103);
xor U12354 (N_12354,N_12125,N_12156);
and U12355 (N_12355,N_12040,N_12060);
xor U12356 (N_12356,N_12114,N_12167);
and U12357 (N_12357,N_12115,N_12181);
nand U12358 (N_12358,N_12179,N_12149);
and U12359 (N_12359,N_12123,N_12164);
nor U12360 (N_12360,N_12048,N_12028);
nand U12361 (N_12361,N_12052,N_12158);
and U12362 (N_12362,N_12019,N_12087);
xnor U12363 (N_12363,N_12112,N_12137);
or U12364 (N_12364,N_12197,N_12021);
or U12365 (N_12365,N_12045,N_12086);
xnor U12366 (N_12366,N_12014,N_12170);
xor U12367 (N_12367,N_12118,N_12107);
xor U12368 (N_12368,N_12087,N_12173);
nand U12369 (N_12369,N_12195,N_12112);
or U12370 (N_12370,N_12068,N_12190);
xnor U12371 (N_12371,N_12164,N_12125);
nor U12372 (N_12372,N_12021,N_12100);
and U12373 (N_12373,N_12029,N_12196);
xnor U12374 (N_12374,N_12095,N_12100);
and U12375 (N_12375,N_12015,N_12134);
or U12376 (N_12376,N_12026,N_12136);
and U12377 (N_12377,N_12156,N_12183);
nor U12378 (N_12378,N_12155,N_12086);
or U12379 (N_12379,N_12167,N_12031);
and U12380 (N_12380,N_12178,N_12040);
xor U12381 (N_12381,N_12156,N_12112);
and U12382 (N_12382,N_12087,N_12199);
xnor U12383 (N_12383,N_12105,N_12054);
xor U12384 (N_12384,N_12032,N_12057);
nand U12385 (N_12385,N_12034,N_12149);
nor U12386 (N_12386,N_12004,N_12062);
or U12387 (N_12387,N_12070,N_12111);
xor U12388 (N_12388,N_12020,N_12055);
or U12389 (N_12389,N_12132,N_12019);
nand U12390 (N_12390,N_12087,N_12197);
nand U12391 (N_12391,N_12036,N_12071);
nand U12392 (N_12392,N_12111,N_12143);
nand U12393 (N_12393,N_12080,N_12144);
and U12394 (N_12394,N_12181,N_12034);
nand U12395 (N_12395,N_12132,N_12134);
xnor U12396 (N_12396,N_12197,N_12110);
nor U12397 (N_12397,N_12008,N_12051);
and U12398 (N_12398,N_12065,N_12113);
nand U12399 (N_12399,N_12101,N_12147);
nor U12400 (N_12400,N_12227,N_12389);
nor U12401 (N_12401,N_12326,N_12375);
xnor U12402 (N_12402,N_12296,N_12216);
xor U12403 (N_12403,N_12323,N_12218);
xor U12404 (N_12404,N_12336,N_12374);
or U12405 (N_12405,N_12351,N_12278);
xnor U12406 (N_12406,N_12258,N_12328);
xnor U12407 (N_12407,N_12263,N_12314);
or U12408 (N_12408,N_12357,N_12260);
xnor U12409 (N_12409,N_12319,N_12293);
or U12410 (N_12410,N_12324,N_12322);
nor U12411 (N_12411,N_12238,N_12366);
or U12412 (N_12412,N_12367,N_12231);
and U12413 (N_12413,N_12264,N_12399);
nand U12414 (N_12414,N_12330,N_12362);
xnor U12415 (N_12415,N_12377,N_12368);
xor U12416 (N_12416,N_12267,N_12237);
and U12417 (N_12417,N_12276,N_12348);
nor U12418 (N_12418,N_12302,N_12215);
xor U12419 (N_12419,N_12266,N_12243);
nor U12420 (N_12420,N_12245,N_12200);
or U12421 (N_12421,N_12307,N_12361);
nor U12422 (N_12422,N_12391,N_12311);
and U12423 (N_12423,N_12233,N_12294);
or U12424 (N_12424,N_12340,N_12378);
xor U12425 (N_12425,N_12207,N_12273);
nand U12426 (N_12426,N_12398,N_12371);
nand U12427 (N_12427,N_12315,N_12269);
nor U12428 (N_12428,N_12249,N_12261);
xor U12429 (N_12429,N_12363,N_12262);
or U12430 (N_12430,N_12277,N_12345);
or U12431 (N_12431,N_12338,N_12313);
nand U12432 (N_12432,N_12346,N_12203);
xor U12433 (N_12433,N_12220,N_12270);
and U12434 (N_12434,N_12337,N_12225);
xnor U12435 (N_12435,N_12365,N_12205);
or U12436 (N_12436,N_12382,N_12316);
and U12437 (N_12437,N_12224,N_12221);
nand U12438 (N_12438,N_12247,N_12309);
xnor U12439 (N_12439,N_12254,N_12219);
or U12440 (N_12440,N_12303,N_12201);
and U12441 (N_12441,N_12331,N_12385);
nand U12442 (N_12442,N_12255,N_12356);
and U12443 (N_12443,N_12397,N_12279);
xnor U12444 (N_12444,N_12308,N_12395);
or U12445 (N_12445,N_12268,N_12212);
or U12446 (N_12446,N_12252,N_12253);
nand U12447 (N_12447,N_12259,N_12214);
nor U12448 (N_12448,N_12388,N_12244);
xor U12449 (N_12449,N_12274,N_12290);
nand U12450 (N_12450,N_12226,N_12240);
and U12451 (N_12451,N_12297,N_12206);
nor U12452 (N_12452,N_12347,N_12343);
nor U12453 (N_12453,N_12280,N_12333);
nand U12454 (N_12454,N_12381,N_12256);
and U12455 (N_12455,N_12287,N_12235);
or U12456 (N_12456,N_12339,N_12236);
nand U12457 (N_12457,N_12204,N_12292);
nand U12458 (N_12458,N_12284,N_12310);
nor U12459 (N_12459,N_12370,N_12288);
nor U12460 (N_12460,N_12291,N_12379);
nand U12461 (N_12461,N_12289,N_12305);
xor U12462 (N_12462,N_12239,N_12329);
nand U12463 (N_12463,N_12283,N_12282);
or U12464 (N_12464,N_12392,N_12369);
or U12465 (N_12465,N_12223,N_12286);
or U12466 (N_12466,N_12275,N_12210);
nand U12467 (N_12467,N_12222,N_12334);
xnor U12468 (N_12468,N_12230,N_12271);
nor U12469 (N_12469,N_12390,N_12335);
nor U12470 (N_12470,N_12228,N_12384);
nand U12471 (N_12471,N_12349,N_12301);
and U12472 (N_12472,N_12248,N_12342);
nand U12473 (N_12473,N_12359,N_12354);
or U12474 (N_12474,N_12250,N_12380);
nand U12475 (N_12475,N_12383,N_12320);
or U12476 (N_12476,N_12299,N_12358);
nand U12477 (N_12477,N_12304,N_12373);
or U12478 (N_12478,N_12318,N_12229);
or U12479 (N_12479,N_12393,N_12242);
xnor U12480 (N_12480,N_12202,N_12396);
and U12481 (N_12481,N_12281,N_12352);
or U12482 (N_12482,N_12325,N_12265);
nand U12483 (N_12483,N_12217,N_12211);
nand U12484 (N_12484,N_12355,N_12232);
or U12485 (N_12485,N_12353,N_12394);
or U12486 (N_12486,N_12298,N_12312);
nor U12487 (N_12487,N_12234,N_12350);
xnor U12488 (N_12488,N_12387,N_12295);
nand U12489 (N_12489,N_12300,N_12386);
or U12490 (N_12490,N_12241,N_12306);
nor U12491 (N_12491,N_12327,N_12360);
xnor U12492 (N_12492,N_12257,N_12376);
and U12493 (N_12493,N_12209,N_12332);
nand U12494 (N_12494,N_12208,N_12317);
nor U12495 (N_12495,N_12213,N_12251);
nand U12496 (N_12496,N_12372,N_12246);
xor U12497 (N_12497,N_12321,N_12344);
nand U12498 (N_12498,N_12341,N_12364);
nand U12499 (N_12499,N_12272,N_12285);
or U12500 (N_12500,N_12326,N_12365);
nor U12501 (N_12501,N_12270,N_12324);
nand U12502 (N_12502,N_12215,N_12319);
nand U12503 (N_12503,N_12212,N_12274);
nor U12504 (N_12504,N_12285,N_12317);
xnor U12505 (N_12505,N_12314,N_12299);
and U12506 (N_12506,N_12227,N_12254);
nor U12507 (N_12507,N_12313,N_12303);
xnor U12508 (N_12508,N_12384,N_12259);
or U12509 (N_12509,N_12320,N_12359);
or U12510 (N_12510,N_12359,N_12266);
and U12511 (N_12511,N_12218,N_12368);
nand U12512 (N_12512,N_12264,N_12340);
or U12513 (N_12513,N_12217,N_12378);
xnor U12514 (N_12514,N_12344,N_12304);
nor U12515 (N_12515,N_12327,N_12387);
nand U12516 (N_12516,N_12232,N_12276);
nand U12517 (N_12517,N_12394,N_12258);
nor U12518 (N_12518,N_12363,N_12245);
nor U12519 (N_12519,N_12357,N_12339);
and U12520 (N_12520,N_12303,N_12325);
nand U12521 (N_12521,N_12220,N_12254);
and U12522 (N_12522,N_12302,N_12309);
and U12523 (N_12523,N_12294,N_12372);
or U12524 (N_12524,N_12232,N_12354);
nand U12525 (N_12525,N_12235,N_12399);
and U12526 (N_12526,N_12320,N_12246);
nand U12527 (N_12527,N_12308,N_12209);
or U12528 (N_12528,N_12234,N_12271);
nor U12529 (N_12529,N_12285,N_12344);
or U12530 (N_12530,N_12305,N_12230);
xor U12531 (N_12531,N_12362,N_12368);
nor U12532 (N_12532,N_12224,N_12345);
or U12533 (N_12533,N_12357,N_12340);
and U12534 (N_12534,N_12261,N_12378);
or U12535 (N_12535,N_12310,N_12324);
nor U12536 (N_12536,N_12230,N_12297);
or U12537 (N_12537,N_12220,N_12396);
and U12538 (N_12538,N_12368,N_12397);
nand U12539 (N_12539,N_12385,N_12259);
nor U12540 (N_12540,N_12230,N_12375);
nand U12541 (N_12541,N_12250,N_12286);
and U12542 (N_12542,N_12373,N_12327);
or U12543 (N_12543,N_12242,N_12248);
nor U12544 (N_12544,N_12202,N_12276);
nand U12545 (N_12545,N_12372,N_12314);
and U12546 (N_12546,N_12376,N_12293);
or U12547 (N_12547,N_12311,N_12248);
xor U12548 (N_12548,N_12286,N_12282);
and U12549 (N_12549,N_12253,N_12294);
xnor U12550 (N_12550,N_12301,N_12285);
xnor U12551 (N_12551,N_12250,N_12212);
nor U12552 (N_12552,N_12315,N_12241);
nor U12553 (N_12553,N_12357,N_12352);
and U12554 (N_12554,N_12248,N_12334);
nand U12555 (N_12555,N_12270,N_12217);
and U12556 (N_12556,N_12393,N_12348);
nand U12557 (N_12557,N_12395,N_12223);
nand U12558 (N_12558,N_12219,N_12336);
and U12559 (N_12559,N_12331,N_12275);
xnor U12560 (N_12560,N_12366,N_12332);
or U12561 (N_12561,N_12220,N_12345);
or U12562 (N_12562,N_12368,N_12391);
or U12563 (N_12563,N_12202,N_12352);
nor U12564 (N_12564,N_12212,N_12289);
xnor U12565 (N_12565,N_12282,N_12387);
and U12566 (N_12566,N_12311,N_12356);
xnor U12567 (N_12567,N_12377,N_12289);
or U12568 (N_12568,N_12229,N_12279);
and U12569 (N_12569,N_12288,N_12258);
or U12570 (N_12570,N_12264,N_12379);
xor U12571 (N_12571,N_12270,N_12207);
xnor U12572 (N_12572,N_12241,N_12379);
or U12573 (N_12573,N_12261,N_12346);
nand U12574 (N_12574,N_12369,N_12221);
and U12575 (N_12575,N_12210,N_12221);
nor U12576 (N_12576,N_12260,N_12226);
nand U12577 (N_12577,N_12297,N_12326);
or U12578 (N_12578,N_12266,N_12271);
nor U12579 (N_12579,N_12298,N_12246);
and U12580 (N_12580,N_12282,N_12257);
nand U12581 (N_12581,N_12283,N_12254);
and U12582 (N_12582,N_12396,N_12358);
nor U12583 (N_12583,N_12341,N_12346);
nand U12584 (N_12584,N_12273,N_12270);
xnor U12585 (N_12585,N_12340,N_12393);
nand U12586 (N_12586,N_12249,N_12342);
or U12587 (N_12587,N_12279,N_12298);
and U12588 (N_12588,N_12223,N_12268);
and U12589 (N_12589,N_12379,N_12372);
and U12590 (N_12590,N_12384,N_12271);
nor U12591 (N_12591,N_12365,N_12213);
nand U12592 (N_12592,N_12330,N_12263);
nand U12593 (N_12593,N_12234,N_12260);
and U12594 (N_12594,N_12301,N_12336);
xnor U12595 (N_12595,N_12298,N_12268);
and U12596 (N_12596,N_12258,N_12357);
or U12597 (N_12597,N_12340,N_12383);
xor U12598 (N_12598,N_12325,N_12388);
nand U12599 (N_12599,N_12360,N_12307);
or U12600 (N_12600,N_12415,N_12430);
and U12601 (N_12601,N_12429,N_12534);
and U12602 (N_12602,N_12458,N_12570);
nor U12603 (N_12603,N_12431,N_12549);
nand U12604 (N_12604,N_12420,N_12590);
and U12605 (N_12605,N_12409,N_12428);
or U12606 (N_12606,N_12524,N_12426);
or U12607 (N_12607,N_12538,N_12452);
and U12608 (N_12608,N_12439,N_12487);
nor U12609 (N_12609,N_12578,N_12472);
xnor U12610 (N_12610,N_12521,N_12464);
nor U12611 (N_12611,N_12574,N_12517);
xor U12612 (N_12612,N_12540,N_12412);
xor U12613 (N_12613,N_12539,N_12599);
nand U12614 (N_12614,N_12558,N_12489);
nor U12615 (N_12615,N_12440,N_12403);
and U12616 (N_12616,N_12594,N_12511);
xnor U12617 (N_12617,N_12408,N_12579);
and U12618 (N_12618,N_12566,N_12484);
or U12619 (N_12619,N_12438,N_12477);
or U12620 (N_12620,N_12462,N_12567);
xor U12621 (N_12621,N_12500,N_12402);
nor U12622 (N_12622,N_12564,N_12481);
nand U12623 (N_12623,N_12554,N_12488);
nand U12624 (N_12624,N_12444,N_12585);
nand U12625 (N_12625,N_12407,N_12469);
or U12626 (N_12626,N_12492,N_12457);
and U12627 (N_12627,N_12503,N_12432);
xor U12628 (N_12628,N_12419,N_12421);
or U12629 (N_12629,N_12433,N_12441);
or U12630 (N_12630,N_12411,N_12552);
xnor U12631 (N_12631,N_12446,N_12571);
nand U12632 (N_12632,N_12595,N_12589);
or U12633 (N_12633,N_12475,N_12507);
nand U12634 (N_12634,N_12543,N_12596);
nor U12635 (N_12635,N_12496,N_12527);
nor U12636 (N_12636,N_12453,N_12536);
nor U12637 (N_12637,N_12580,N_12545);
nand U12638 (N_12638,N_12400,N_12401);
nand U12639 (N_12639,N_12502,N_12519);
nand U12640 (N_12640,N_12541,N_12513);
nand U12641 (N_12641,N_12542,N_12476);
xor U12642 (N_12642,N_12576,N_12530);
nor U12643 (N_12643,N_12504,N_12532);
or U12644 (N_12644,N_12510,N_12417);
nor U12645 (N_12645,N_12461,N_12449);
and U12646 (N_12646,N_12582,N_12598);
or U12647 (N_12647,N_12531,N_12568);
xnor U12648 (N_12648,N_12563,N_12495);
and U12649 (N_12649,N_12480,N_12592);
xor U12650 (N_12650,N_12575,N_12544);
or U12651 (N_12651,N_12494,N_12465);
xor U12652 (N_12652,N_12424,N_12479);
or U12653 (N_12653,N_12437,N_12447);
nor U12654 (N_12654,N_12474,N_12587);
nand U12655 (N_12655,N_12478,N_12434);
and U12656 (N_12656,N_12451,N_12445);
and U12657 (N_12657,N_12525,N_12581);
and U12658 (N_12658,N_12456,N_12562);
nand U12659 (N_12659,N_12499,N_12498);
nor U12660 (N_12660,N_12505,N_12435);
or U12661 (N_12661,N_12588,N_12482);
nand U12662 (N_12662,N_12463,N_12526);
nand U12663 (N_12663,N_12506,N_12512);
nand U12664 (N_12664,N_12454,N_12572);
xor U12665 (N_12665,N_12556,N_12597);
nand U12666 (N_12666,N_12548,N_12425);
xor U12667 (N_12667,N_12561,N_12547);
and U12668 (N_12668,N_12491,N_12553);
nand U12669 (N_12669,N_12422,N_12450);
nand U12670 (N_12670,N_12523,N_12467);
or U12671 (N_12671,N_12518,N_12528);
nor U12672 (N_12672,N_12546,N_12473);
nand U12673 (N_12673,N_12577,N_12586);
nand U12674 (N_12674,N_12485,N_12406);
nand U12675 (N_12675,N_12559,N_12466);
and U12676 (N_12676,N_12460,N_12529);
nor U12677 (N_12677,N_12483,N_12497);
and U12678 (N_12678,N_12442,N_12509);
and U12679 (N_12679,N_12501,N_12416);
and U12680 (N_12680,N_12423,N_12516);
nand U12681 (N_12681,N_12573,N_12560);
nand U12682 (N_12682,N_12593,N_12535);
and U12683 (N_12683,N_12569,N_12583);
and U12684 (N_12684,N_12515,N_12427);
nor U12685 (N_12685,N_12533,N_12443);
or U12686 (N_12686,N_12459,N_12404);
nor U12687 (N_12687,N_12520,N_12514);
xnor U12688 (N_12688,N_12468,N_12584);
or U12689 (N_12689,N_12490,N_12414);
xor U12690 (N_12690,N_12448,N_12508);
nor U12691 (N_12691,N_12455,N_12551);
nor U12692 (N_12692,N_12550,N_12493);
and U12693 (N_12693,N_12591,N_12522);
nand U12694 (N_12694,N_12413,N_12565);
and U12695 (N_12695,N_12486,N_12537);
nand U12696 (N_12696,N_12471,N_12470);
or U12697 (N_12697,N_12555,N_12436);
nor U12698 (N_12698,N_12557,N_12405);
nor U12699 (N_12699,N_12410,N_12418);
nand U12700 (N_12700,N_12439,N_12585);
and U12701 (N_12701,N_12568,N_12403);
nor U12702 (N_12702,N_12575,N_12541);
and U12703 (N_12703,N_12516,N_12496);
or U12704 (N_12704,N_12539,N_12587);
xnor U12705 (N_12705,N_12401,N_12561);
nand U12706 (N_12706,N_12563,N_12566);
or U12707 (N_12707,N_12409,N_12488);
nor U12708 (N_12708,N_12411,N_12500);
nand U12709 (N_12709,N_12485,N_12481);
or U12710 (N_12710,N_12439,N_12586);
nor U12711 (N_12711,N_12555,N_12574);
nor U12712 (N_12712,N_12558,N_12437);
and U12713 (N_12713,N_12502,N_12496);
or U12714 (N_12714,N_12489,N_12562);
nand U12715 (N_12715,N_12439,N_12435);
and U12716 (N_12716,N_12582,N_12492);
nor U12717 (N_12717,N_12517,N_12489);
nor U12718 (N_12718,N_12435,N_12506);
nor U12719 (N_12719,N_12572,N_12539);
nand U12720 (N_12720,N_12442,N_12406);
nor U12721 (N_12721,N_12407,N_12596);
nor U12722 (N_12722,N_12515,N_12571);
and U12723 (N_12723,N_12502,N_12530);
and U12724 (N_12724,N_12469,N_12556);
or U12725 (N_12725,N_12507,N_12533);
nand U12726 (N_12726,N_12491,N_12480);
nand U12727 (N_12727,N_12597,N_12530);
nor U12728 (N_12728,N_12460,N_12566);
nand U12729 (N_12729,N_12497,N_12489);
and U12730 (N_12730,N_12472,N_12528);
xnor U12731 (N_12731,N_12507,N_12513);
nand U12732 (N_12732,N_12436,N_12569);
and U12733 (N_12733,N_12452,N_12505);
or U12734 (N_12734,N_12454,N_12556);
nor U12735 (N_12735,N_12440,N_12450);
nand U12736 (N_12736,N_12577,N_12561);
nand U12737 (N_12737,N_12593,N_12528);
xor U12738 (N_12738,N_12556,N_12587);
or U12739 (N_12739,N_12572,N_12486);
and U12740 (N_12740,N_12491,N_12568);
and U12741 (N_12741,N_12472,N_12440);
or U12742 (N_12742,N_12483,N_12420);
and U12743 (N_12743,N_12583,N_12479);
and U12744 (N_12744,N_12427,N_12550);
xnor U12745 (N_12745,N_12554,N_12573);
nand U12746 (N_12746,N_12595,N_12415);
and U12747 (N_12747,N_12500,N_12513);
nor U12748 (N_12748,N_12510,N_12468);
nand U12749 (N_12749,N_12561,N_12418);
and U12750 (N_12750,N_12579,N_12543);
nand U12751 (N_12751,N_12590,N_12419);
and U12752 (N_12752,N_12412,N_12435);
xnor U12753 (N_12753,N_12421,N_12464);
or U12754 (N_12754,N_12426,N_12536);
or U12755 (N_12755,N_12447,N_12460);
or U12756 (N_12756,N_12463,N_12400);
and U12757 (N_12757,N_12550,N_12464);
nor U12758 (N_12758,N_12571,N_12536);
or U12759 (N_12759,N_12429,N_12491);
or U12760 (N_12760,N_12452,N_12533);
and U12761 (N_12761,N_12500,N_12520);
nor U12762 (N_12762,N_12456,N_12419);
nor U12763 (N_12763,N_12578,N_12498);
xnor U12764 (N_12764,N_12416,N_12468);
or U12765 (N_12765,N_12438,N_12468);
and U12766 (N_12766,N_12460,N_12469);
or U12767 (N_12767,N_12581,N_12532);
or U12768 (N_12768,N_12565,N_12471);
and U12769 (N_12769,N_12465,N_12509);
and U12770 (N_12770,N_12544,N_12533);
nand U12771 (N_12771,N_12528,N_12534);
xor U12772 (N_12772,N_12506,N_12423);
xor U12773 (N_12773,N_12487,N_12454);
and U12774 (N_12774,N_12449,N_12552);
and U12775 (N_12775,N_12506,N_12470);
or U12776 (N_12776,N_12588,N_12473);
xnor U12777 (N_12777,N_12504,N_12426);
xnor U12778 (N_12778,N_12495,N_12411);
or U12779 (N_12779,N_12462,N_12451);
or U12780 (N_12780,N_12400,N_12498);
and U12781 (N_12781,N_12455,N_12421);
xnor U12782 (N_12782,N_12497,N_12531);
or U12783 (N_12783,N_12599,N_12466);
nor U12784 (N_12784,N_12464,N_12403);
nand U12785 (N_12785,N_12473,N_12466);
and U12786 (N_12786,N_12509,N_12431);
and U12787 (N_12787,N_12526,N_12482);
xnor U12788 (N_12788,N_12511,N_12429);
nand U12789 (N_12789,N_12414,N_12549);
or U12790 (N_12790,N_12560,N_12594);
xnor U12791 (N_12791,N_12419,N_12513);
nor U12792 (N_12792,N_12557,N_12502);
nand U12793 (N_12793,N_12581,N_12483);
nor U12794 (N_12794,N_12447,N_12405);
nor U12795 (N_12795,N_12471,N_12511);
and U12796 (N_12796,N_12547,N_12537);
nor U12797 (N_12797,N_12507,N_12470);
and U12798 (N_12798,N_12409,N_12486);
and U12799 (N_12799,N_12405,N_12473);
and U12800 (N_12800,N_12685,N_12671);
or U12801 (N_12801,N_12678,N_12626);
or U12802 (N_12802,N_12665,N_12780);
or U12803 (N_12803,N_12703,N_12660);
nor U12804 (N_12804,N_12726,N_12607);
nand U12805 (N_12805,N_12604,N_12794);
nor U12806 (N_12806,N_12619,N_12750);
nor U12807 (N_12807,N_12624,N_12782);
xor U12808 (N_12808,N_12630,N_12729);
and U12809 (N_12809,N_12783,N_12767);
xnor U12810 (N_12810,N_12734,N_12719);
nor U12811 (N_12811,N_12778,N_12658);
xor U12812 (N_12812,N_12736,N_12768);
and U12813 (N_12813,N_12614,N_12643);
nor U12814 (N_12814,N_12668,N_12664);
xnor U12815 (N_12815,N_12642,N_12702);
xnor U12816 (N_12816,N_12789,N_12681);
nor U12817 (N_12817,N_12762,N_12717);
nand U12818 (N_12818,N_12733,N_12779);
and U12819 (N_12819,N_12752,N_12628);
xnor U12820 (N_12820,N_12636,N_12603);
or U12821 (N_12821,N_12649,N_12606);
and U12822 (N_12822,N_12797,N_12600);
or U12823 (N_12823,N_12730,N_12735);
nor U12824 (N_12824,N_12674,N_12633);
and U12825 (N_12825,N_12713,N_12682);
nor U12826 (N_12826,N_12712,N_12722);
and U12827 (N_12827,N_12670,N_12708);
xnor U12828 (N_12828,N_12621,N_12721);
nand U12829 (N_12829,N_12724,N_12666);
or U12830 (N_12830,N_12707,N_12749);
nor U12831 (N_12831,N_12739,N_12781);
or U12832 (N_12832,N_12646,N_12746);
nand U12833 (N_12833,N_12798,N_12645);
nand U12834 (N_12834,N_12617,N_12623);
nor U12835 (N_12835,N_12747,N_12743);
xnor U12836 (N_12836,N_12709,N_12676);
xor U12837 (N_12837,N_12696,N_12662);
nand U12838 (N_12838,N_12745,N_12710);
or U12839 (N_12839,N_12799,N_12715);
or U12840 (N_12840,N_12615,N_12706);
nor U12841 (N_12841,N_12700,N_12756);
nor U12842 (N_12842,N_12686,N_12687);
nor U12843 (N_12843,N_12693,N_12785);
xor U12844 (N_12844,N_12601,N_12644);
nand U12845 (N_12845,N_12656,N_12701);
or U12846 (N_12846,N_12788,N_12769);
xor U12847 (N_12847,N_12766,N_12631);
xnor U12848 (N_12848,N_12753,N_12773);
nor U12849 (N_12849,N_12611,N_12759);
or U12850 (N_12850,N_12692,N_12669);
xor U12851 (N_12851,N_12791,N_12772);
nor U12852 (N_12852,N_12697,N_12672);
and U12853 (N_12853,N_12770,N_12684);
nand U12854 (N_12854,N_12758,N_12629);
xnor U12855 (N_12855,N_12732,N_12775);
nor U12856 (N_12856,N_12680,N_12638);
or U12857 (N_12857,N_12690,N_12663);
xnor U12858 (N_12858,N_12716,N_12725);
nand U12859 (N_12859,N_12764,N_12667);
nand U12860 (N_12860,N_12659,N_12741);
xor U12861 (N_12861,N_12618,N_12748);
or U12862 (N_12862,N_12627,N_12647);
or U12863 (N_12863,N_12795,N_12634);
and U12864 (N_12864,N_12771,N_12784);
and U12865 (N_12865,N_12723,N_12639);
xnor U12866 (N_12866,N_12792,N_12657);
or U12867 (N_12867,N_12738,N_12728);
xor U12868 (N_12868,N_12737,N_12613);
and U12869 (N_12869,N_12760,N_12776);
xnor U12870 (N_12870,N_12742,N_12637);
nor U12871 (N_12871,N_12605,N_12622);
or U12872 (N_12872,N_12757,N_12793);
and U12873 (N_12873,N_12786,N_12694);
and U12874 (N_12874,N_12661,N_12689);
and U12875 (N_12875,N_12744,N_12691);
or U12876 (N_12876,N_12616,N_12673);
and U12877 (N_12877,N_12777,N_12731);
or U12878 (N_12878,N_12612,N_12765);
nand U12879 (N_12879,N_12763,N_12740);
and U12880 (N_12880,N_12608,N_12695);
or U12881 (N_12881,N_12755,N_12754);
nor U12882 (N_12882,N_12675,N_12610);
or U12883 (N_12883,N_12654,N_12640);
nor U12884 (N_12884,N_12698,N_12727);
nor U12885 (N_12885,N_12796,N_12704);
or U12886 (N_12886,N_12632,N_12774);
nand U12887 (N_12887,N_12761,N_12679);
nand U12888 (N_12888,N_12718,N_12705);
nor U12889 (N_12889,N_12650,N_12651);
nor U12890 (N_12890,N_12787,N_12714);
nand U12891 (N_12891,N_12688,N_12620);
or U12892 (N_12892,N_12641,N_12653);
and U12893 (N_12893,N_12751,N_12635);
xor U12894 (N_12894,N_12790,N_12609);
and U12895 (N_12895,N_12683,N_12652);
and U12896 (N_12896,N_12602,N_12720);
nor U12897 (N_12897,N_12625,N_12655);
or U12898 (N_12898,N_12677,N_12699);
and U12899 (N_12899,N_12711,N_12648);
nor U12900 (N_12900,N_12710,N_12777);
and U12901 (N_12901,N_12791,N_12627);
nand U12902 (N_12902,N_12705,N_12697);
and U12903 (N_12903,N_12696,N_12660);
or U12904 (N_12904,N_12644,N_12658);
xor U12905 (N_12905,N_12708,N_12707);
nand U12906 (N_12906,N_12694,N_12779);
and U12907 (N_12907,N_12648,N_12707);
nor U12908 (N_12908,N_12716,N_12666);
and U12909 (N_12909,N_12627,N_12761);
xnor U12910 (N_12910,N_12794,N_12695);
nand U12911 (N_12911,N_12682,N_12752);
nor U12912 (N_12912,N_12645,N_12667);
nor U12913 (N_12913,N_12762,N_12783);
and U12914 (N_12914,N_12709,N_12602);
xnor U12915 (N_12915,N_12624,N_12600);
or U12916 (N_12916,N_12670,N_12687);
xor U12917 (N_12917,N_12684,N_12715);
or U12918 (N_12918,N_12720,N_12770);
nor U12919 (N_12919,N_12666,N_12604);
xnor U12920 (N_12920,N_12798,N_12788);
nor U12921 (N_12921,N_12713,N_12652);
nand U12922 (N_12922,N_12782,N_12757);
xnor U12923 (N_12923,N_12634,N_12779);
nand U12924 (N_12924,N_12638,N_12796);
and U12925 (N_12925,N_12722,N_12733);
nor U12926 (N_12926,N_12627,N_12642);
nand U12927 (N_12927,N_12688,N_12747);
and U12928 (N_12928,N_12775,N_12640);
and U12929 (N_12929,N_12691,N_12707);
and U12930 (N_12930,N_12770,N_12682);
xor U12931 (N_12931,N_12760,N_12680);
or U12932 (N_12932,N_12738,N_12763);
nand U12933 (N_12933,N_12650,N_12694);
or U12934 (N_12934,N_12609,N_12638);
nand U12935 (N_12935,N_12733,N_12606);
nor U12936 (N_12936,N_12688,N_12636);
nand U12937 (N_12937,N_12696,N_12794);
nand U12938 (N_12938,N_12659,N_12667);
and U12939 (N_12939,N_12759,N_12687);
nand U12940 (N_12940,N_12714,N_12703);
and U12941 (N_12941,N_12736,N_12684);
xnor U12942 (N_12942,N_12790,N_12636);
or U12943 (N_12943,N_12618,N_12605);
nor U12944 (N_12944,N_12712,N_12628);
and U12945 (N_12945,N_12637,N_12720);
xor U12946 (N_12946,N_12718,N_12655);
and U12947 (N_12947,N_12609,N_12764);
and U12948 (N_12948,N_12746,N_12629);
xnor U12949 (N_12949,N_12650,N_12750);
or U12950 (N_12950,N_12631,N_12712);
nand U12951 (N_12951,N_12772,N_12682);
nor U12952 (N_12952,N_12632,N_12796);
and U12953 (N_12953,N_12616,N_12760);
or U12954 (N_12954,N_12659,N_12682);
nand U12955 (N_12955,N_12715,N_12778);
nor U12956 (N_12956,N_12748,N_12778);
and U12957 (N_12957,N_12684,N_12649);
or U12958 (N_12958,N_12732,N_12728);
nand U12959 (N_12959,N_12773,N_12786);
and U12960 (N_12960,N_12682,N_12730);
nor U12961 (N_12961,N_12730,N_12616);
and U12962 (N_12962,N_12603,N_12664);
nor U12963 (N_12963,N_12604,N_12605);
and U12964 (N_12964,N_12714,N_12798);
or U12965 (N_12965,N_12750,N_12747);
or U12966 (N_12966,N_12607,N_12605);
or U12967 (N_12967,N_12728,N_12652);
xnor U12968 (N_12968,N_12603,N_12744);
or U12969 (N_12969,N_12656,N_12643);
nand U12970 (N_12970,N_12611,N_12709);
nor U12971 (N_12971,N_12612,N_12685);
xnor U12972 (N_12972,N_12770,N_12731);
nor U12973 (N_12973,N_12641,N_12780);
or U12974 (N_12974,N_12718,N_12628);
nand U12975 (N_12975,N_12775,N_12636);
xnor U12976 (N_12976,N_12704,N_12687);
nor U12977 (N_12977,N_12705,N_12750);
or U12978 (N_12978,N_12711,N_12783);
nand U12979 (N_12979,N_12795,N_12659);
nor U12980 (N_12980,N_12756,N_12705);
and U12981 (N_12981,N_12799,N_12653);
nor U12982 (N_12982,N_12685,N_12676);
and U12983 (N_12983,N_12654,N_12634);
nand U12984 (N_12984,N_12787,N_12729);
nor U12985 (N_12985,N_12649,N_12773);
nand U12986 (N_12986,N_12765,N_12709);
and U12987 (N_12987,N_12650,N_12764);
xnor U12988 (N_12988,N_12722,N_12743);
nor U12989 (N_12989,N_12709,N_12734);
nand U12990 (N_12990,N_12760,N_12786);
and U12991 (N_12991,N_12761,N_12736);
and U12992 (N_12992,N_12664,N_12635);
and U12993 (N_12993,N_12756,N_12792);
nand U12994 (N_12994,N_12728,N_12699);
nor U12995 (N_12995,N_12774,N_12748);
xnor U12996 (N_12996,N_12670,N_12774);
xor U12997 (N_12997,N_12614,N_12734);
nand U12998 (N_12998,N_12725,N_12759);
or U12999 (N_12999,N_12649,N_12659);
and U13000 (N_13000,N_12964,N_12828);
nand U13001 (N_13001,N_12839,N_12884);
or U13002 (N_13002,N_12879,N_12933);
xor U13003 (N_13003,N_12892,N_12917);
nand U13004 (N_13004,N_12972,N_12926);
xnor U13005 (N_13005,N_12919,N_12912);
and U13006 (N_13006,N_12890,N_12947);
nand U13007 (N_13007,N_12959,N_12812);
nand U13008 (N_13008,N_12814,N_12853);
or U13009 (N_13009,N_12843,N_12968);
or U13010 (N_13010,N_12872,N_12992);
nor U13011 (N_13011,N_12916,N_12988);
xor U13012 (N_13012,N_12954,N_12813);
nand U13013 (N_13013,N_12880,N_12990);
or U13014 (N_13014,N_12823,N_12845);
nor U13015 (N_13015,N_12909,N_12913);
nand U13016 (N_13016,N_12818,N_12961);
nor U13017 (N_13017,N_12866,N_12971);
and U13018 (N_13018,N_12967,N_12918);
nand U13019 (N_13019,N_12958,N_12855);
nand U13020 (N_13020,N_12978,N_12973);
xnor U13021 (N_13021,N_12851,N_12861);
xnor U13022 (N_13022,N_12834,N_12897);
xor U13023 (N_13023,N_12952,N_12910);
nor U13024 (N_13024,N_12960,N_12935);
or U13025 (N_13025,N_12955,N_12877);
and U13026 (N_13026,N_12966,N_12941);
nand U13027 (N_13027,N_12948,N_12943);
nor U13028 (N_13028,N_12822,N_12827);
nor U13029 (N_13029,N_12956,N_12894);
xor U13030 (N_13030,N_12929,N_12805);
nor U13031 (N_13031,N_12907,N_12920);
or U13032 (N_13032,N_12859,N_12840);
nand U13033 (N_13033,N_12825,N_12835);
nand U13034 (N_13034,N_12923,N_12831);
or U13035 (N_13035,N_12821,N_12854);
xor U13036 (N_13036,N_12815,N_12934);
or U13037 (N_13037,N_12870,N_12932);
xor U13038 (N_13038,N_12982,N_12829);
or U13039 (N_13039,N_12881,N_12819);
and U13040 (N_13040,N_12882,N_12950);
xnor U13041 (N_13041,N_12974,N_12915);
xnor U13042 (N_13042,N_12985,N_12981);
nor U13043 (N_13043,N_12945,N_12969);
nor U13044 (N_13044,N_12875,N_12849);
xor U13045 (N_13045,N_12807,N_12963);
xor U13046 (N_13046,N_12864,N_12977);
xor U13047 (N_13047,N_12886,N_12832);
nor U13048 (N_13048,N_12804,N_12997);
xnor U13049 (N_13049,N_12984,N_12893);
xnor U13050 (N_13050,N_12946,N_12937);
nor U13051 (N_13051,N_12836,N_12820);
xor U13052 (N_13052,N_12924,N_12994);
nor U13053 (N_13053,N_12824,N_12962);
nor U13054 (N_13054,N_12806,N_12979);
nor U13055 (N_13055,N_12904,N_12993);
nor U13056 (N_13056,N_12878,N_12908);
or U13057 (N_13057,N_12848,N_12888);
or U13058 (N_13058,N_12949,N_12808);
and U13059 (N_13059,N_12899,N_12970);
or U13060 (N_13060,N_12914,N_12802);
xnor U13061 (N_13061,N_12930,N_12857);
xor U13062 (N_13062,N_12896,N_12965);
xnor U13063 (N_13063,N_12906,N_12800);
nor U13064 (N_13064,N_12856,N_12844);
nand U13065 (N_13065,N_12922,N_12957);
or U13066 (N_13066,N_12816,N_12873);
nand U13067 (N_13067,N_12951,N_12989);
xnor U13068 (N_13068,N_12987,N_12903);
and U13069 (N_13069,N_12931,N_12865);
nor U13070 (N_13070,N_12858,N_12983);
nor U13071 (N_13071,N_12811,N_12868);
nand U13072 (N_13072,N_12911,N_12841);
nor U13073 (N_13073,N_12837,N_12901);
or U13074 (N_13074,N_12801,N_12826);
or U13075 (N_13075,N_12921,N_12852);
or U13076 (N_13076,N_12928,N_12939);
nor U13077 (N_13077,N_12867,N_12871);
nor U13078 (N_13078,N_12838,N_12869);
nor U13079 (N_13079,N_12944,N_12887);
nor U13080 (N_13080,N_12891,N_12810);
nand U13081 (N_13081,N_12998,N_12833);
nor U13082 (N_13082,N_12938,N_12883);
or U13083 (N_13083,N_12986,N_12927);
xor U13084 (N_13084,N_12847,N_12940);
xnor U13085 (N_13085,N_12850,N_12942);
nand U13086 (N_13086,N_12830,N_12900);
or U13087 (N_13087,N_12936,N_12889);
and U13088 (N_13088,N_12999,N_12803);
xnor U13089 (N_13089,N_12846,N_12953);
xnor U13090 (N_13090,N_12975,N_12860);
or U13091 (N_13091,N_12876,N_12902);
nand U13092 (N_13092,N_12925,N_12980);
and U13093 (N_13093,N_12991,N_12874);
nand U13094 (N_13094,N_12817,N_12905);
or U13095 (N_13095,N_12842,N_12885);
and U13096 (N_13096,N_12863,N_12898);
or U13097 (N_13097,N_12995,N_12976);
or U13098 (N_13098,N_12809,N_12996);
nand U13099 (N_13099,N_12862,N_12895);
xor U13100 (N_13100,N_12825,N_12841);
nor U13101 (N_13101,N_12963,N_12837);
or U13102 (N_13102,N_12967,N_12883);
xor U13103 (N_13103,N_12934,N_12832);
and U13104 (N_13104,N_12838,N_12842);
and U13105 (N_13105,N_12853,N_12835);
xnor U13106 (N_13106,N_12964,N_12986);
nor U13107 (N_13107,N_12982,N_12986);
nor U13108 (N_13108,N_12935,N_12873);
nor U13109 (N_13109,N_12982,N_12841);
xor U13110 (N_13110,N_12832,N_12811);
or U13111 (N_13111,N_12845,N_12916);
xnor U13112 (N_13112,N_12932,N_12969);
nor U13113 (N_13113,N_12855,N_12866);
and U13114 (N_13114,N_12927,N_12873);
and U13115 (N_13115,N_12949,N_12885);
nor U13116 (N_13116,N_12942,N_12852);
xnor U13117 (N_13117,N_12996,N_12956);
or U13118 (N_13118,N_12925,N_12916);
nor U13119 (N_13119,N_12954,N_12971);
nor U13120 (N_13120,N_12854,N_12848);
nor U13121 (N_13121,N_12959,N_12925);
xnor U13122 (N_13122,N_12901,N_12874);
nand U13123 (N_13123,N_12841,N_12882);
xnor U13124 (N_13124,N_12993,N_12984);
xor U13125 (N_13125,N_12924,N_12996);
and U13126 (N_13126,N_12975,N_12853);
nand U13127 (N_13127,N_12855,N_12844);
nor U13128 (N_13128,N_12842,N_12874);
nand U13129 (N_13129,N_12816,N_12832);
nand U13130 (N_13130,N_12931,N_12867);
nand U13131 (N_13131,N_12843,N_12943);
and U13132 (N_13132,N_12981,N_12888);
nand U13133 (N_13133,N_12903,N_12853);
xor U13134 (N_13134,N_12912,N_12973);
xnor U13135 (N_13135,N_12916,N_12942);
nor U13136 (N_13136,N_12832,N_12904);
nor U13137 (N_13137,N_12987,N_12938);
nand U13138 (N_13138,N_12824,N_12964);
nand U13139 (N_13139,N_12966,N_12912);
and U13140 (N_13140,N_12809,N_12934);
nor U13141 (N_13141,N_12813,N_12891);
xnor U13142 (N_13142,N_12824,N_12916);
xnor U13143 (N_13143,N_12819,N_12850);
nand U13144 (N_13144,N_12998,N_12860);
and U13145 (N_13145,N_12994,N_12969);
or U13146 (N_13146,N_12973,N_12848);
and U13147 (N_13147,N_12983,N_12870);
and U13148 (N_13148,N_12916,N_12972);
nand U13149 (N_13149,N_12964,N_12901);
and U13150 (N_13150,N_12815,N_12928);
or U13151 (N_13151,N_12822,N_12991);
and U13152 (N_13152,N_12808,N_12894);
or U13153 (N_13153,N_12998,N_12827);
xor U13154 (N_13154,N_12955,N_12855);
nor U13155 (N_13155,N_12880,N_12967);
nand U13156 (N_13156,N_12931,N_12903);
xor U13157 (N_13157,N_12942,N_12893);
or U13158 (N_13158,N_12876,N_12984);
and U13159 (N_13159,N_12814,N_12845);
and U13160 (N_13160,N_12869,N_12959);
xor U13161 (N_13161,N_12956,N_12938);
and U13162 (N_13162,N_12873,N_12946);
and U13163 (N_13163,N_12992,N_12978);
nor U13164 (N_13164,N_12850,N_12965);
nor U13165 (N_13165,N_12928,N_12970);
xnor U13166 (N_13166,N_12824,N_12883);
nor U13167 (N_13167,N_12997,N_12911);
xor U13168 (N_13168,N_12868,N_12807);
and U13169 (N_13169,N_12975,N_12907);
nand U13170 (N_13170,N_12989,N_12901);
nor U13171 (N_13171,N_12942,N_12855);
nand U13172 (N_13172,N_12813,N_12915);
nor U13173 (N_13173,N_12975,N_12810);
nor U13174 (N_13174,N_12804,N_12865);
and U13175 (N_13175,N_12934,N_12866);
and U13176 (N_13176,N_12877,N_12990);
xor U13177 (N_13177,N_12912,N_12892);
xor U13178 (N_13178,N_12985,N_12902);
or U13179 (N_13179,N_12934,N_12910);
nor U13180 (N_13180,N_12953,N_12837);
nand U13181 (N_13181,N_12896,N_12999);
and U13182 (N_13182,N_12802,N_12951);
nor U13183 (N_13183,N_12863,N_12960);
and U13184 (N_13184,N_12909,N_12959);
or U13185 (N_13185,N_12829,N_12834);
nor U13186 (N_13186,N_12945,N_12816);
nor U13187 (N_13187,N_12827,N_12826);
nor U13188 (N_13188,N_12916,N_12937);
nor U13189 (N_13189,N_12813,N_12910);
and U13190 (N_13190,N_12822,N_12964);
xnor U13191 (N_13191,N_12813,N_12876);
nor U13192 (N_13192,N_12985,N_12943);
and U13193 (N_13193,N_12872,N_12861);
nor U13194 (N_13194,N_12992,N_12991);
xor U13195 (N_13195,N_12999,N_12965);
nor U13196 (N_13196,N_12827,N_12803);
and U13197 (N_13197,N_12914,N_12982);
nand U13198 (N_13198,N_12895,N_12851);
nand U13199 (N_13199,N_12819,N_12835);
and U13200 (N_13200,N_13109,N_13011);
xor U13201 (N_13201,N_13181,N_13035);
xor U13202 (N_13202,N_13072,N_13089);
nand U13203 (N_13203,N_13069,N_13194);
nor U13204 (N_13204,N_13047,N_13138);
nor U13205 (N_13205,N_13091,N_13110);
and U13206 (N_13206,N_13193,N_13192);
nand U13207 (N_13207,N_13198,N_13134);
nor U13208 (N_13208,N_13133,N_13088);
nor U13209 (N_13209,N_13187,N_13175);
or U13210 (N_13210,N_13043,N_13008);
or U13211 (N_13211,N_13017,N_13151);
nor U13212 (N_13212,N_13006,N_13136);
nor U13213 (N_13213,N_13118,N_13122);
or U13214 (N_13214,N_13016,N_13082);
xor U13215 (N_13215,N_13195,N_13038);
xor U13216 (N_13216,N_13165,N_13179);
nand U13217 (N_13217,N_13084,N_13028);
and U13218 (N_13218,N_13097,N_13183);
nor U13219 (N_13219,N_13056,N_13111);
nand U13220 (N_13220,N_13106,N_13157);
nand U13221 (N_13221,N_13046,N_13108);
or U13222 (N_13222,N_13124,N_13184);
nor U13223 (N_13223,N_13182,N_13103);
xor U13224 (N_13224,N_13155,N_13126);
xor U13225 (N_13225,N_13015,N_13197);
xor U13226 (N_13226,N_13003,N_13114);
or U13227 (N_13227,N_13079,N_13098);
and U13228 (N_13228,N_13123,N_13077);
nor U13229 (N_13229,N_13050,N_13113);
xor U13230 (N_13230,N_13009,N_13099);
xnor U13231 (N_13231,N_13093,N_13018);
and U13232 (N_13232,N_13086,N_13154);
nand U13233 (N_13233,N_13125,N_13068);
and U13234 (N_13234,N_13166,N_13051);
nor U13235 (N_13235,N_13104,N_13039);
nand U13236 (N_13236,N_13169,N_13066);
nand U13237 (N_13237,N_13170,N_13145);
nor U13238 (N_13238,N_13112,N_13080);
and U13239 (N_13239,N_13027,N_13115);
nor U13240 (N_13240,N_13004,N_13160);
and U13241 (N_13241,N_13119,N_13020);
and U13242 (N_13242,N_13025,N_13094);
nand U13243 (N_13243,N_13161,N_13162);
nand U13244 (N_13244,N_13012,N_13107);
and U13245 (N_13245,N_13022,N_13167);
nand U13246 (N_13246,N_13152,N_13054);
nor U13247 (N_13247,N_13031,N_13085);
nor U13248 (N_13248,N_13007,N_13135);
xnor U13249 (N_13249,N_13100,N_13021);
nand U13250 (N_13250,N_13023,N_13001);
xnor U13251 (N_13251,N_13164,N_13173);
and U13252 (N_13252,N_13137,N_13143);
xor U13253 (N_13253,N_13096,N_13042);
nand U13254 (N_13254,N_13055,N_13188);
and U13255 (N_13255,N_13177,N_13074);
xnor U13256 (N_13256,N_13142,N_13024);
nor U13257 (N_13257,N_13057,N_13064);
or U13258 (N_13258,N_13146,N_13159);
and U13259 (N_13259,N_13190,N_13095);
nand U13260 (N_13260,N_13034,N_13002);
and U13261 (N_13261,N_13102,N_13153);
nand U13262 (N_13262,N_13090,N_13156);
and U13263 (N_13263,N_13185,N_13014);
or U13264 (N_13264,N_13144,N_13150);
nor U13265 (N_13265,N_13073,N_13148);
or U13266 (N_13266,N_13130,N_13058);
and U13267 (N_13267,N_13172,N_13129);
nor U13268 (N_13268,N_13070,N_13147);
and U13269 (N_13269,N_13128,N_13180);
or U13270 (N_13270,N_13076,N_13045);
or U13271 (N_13271,N_13174,N_13120);
and U13272 (N_13272,N_13067,N_13116);
xnor U13273 (N_13273,N_13013,N_13037);
or U13274 (N_13274,N_13105,N_13117);
nand U13275 (N_13275,N_13127,N_13078);
nand U13276 (N_13276,N_13032,N_13041);
or U13277 (N_13277,N_13000,N_13065);
nor U13278 (N_13278,N_13092,N_13189);
and U13279 (N_13279,N_13040,N_13049);
xnor U13280 (N_13280,N_13176,N_13158);
or U13281 (N_13281,N_13171,N_13071);
nor U13282 (N_13282,N_13121,N_13062);
or U13283 (N_13283,N_13178,N_13063);
nand U13284 (N_13284,N_13061,N_13048);
xor U13285 (N_13285,N_13059,N_13060);
nand U13286 (N_13286,N_13141,N_13199);
nor U13287 (N_13287,N_13030,N_13101);
or U13288 (N_13288,N_13044,N_13026);
nor U13289 (N_13289,N_13191,N_13029);
nand U13290 (N_13290,N_13186,N_13087);
and U13291 (N_13291,N_13081,N_13036);
or U13292 (N_13292,N_13140,N_13033);
nor U13293 (N_13293,N_13149,N_13075);
nor U13294 (N_13294,N_13163,N_13052);
nand U13295 (N_13295,N_13010,N_13139);
nor U13296 (N_13296,N_13132,N_13083);
and U13297 (N_13297,N_13005,N_13019);
or U13298 (N_13298,N_13131,N_13196);
or U13299 (N_13299,N_13053,N_13168);
and U13300 (N_13300,N_13104,N_13091);
nor U13301 (N_13301,N_13071,N_13115);
and U13302 (N_13302,N_13090,N_13035);
and U13303 (N_13303,N_13139,N_13005);
nor U13304 (N_13304,N_13126,N_13004);
nor U13305 (N_13305,N_13006,N_13043);
nand U13306 (N_13306,N_13118,N_13111);
nand U13307 (N_13307,N_13131,N_13190);
nor U13308 (N_13308,N_13005,N_13041);
nand U13309 (N_13309,N_13095,N_13096);
nor U13310 (N_13310,N_13187,N_13196);
xor U13311 (N_13311,N_13088,N_13011);
or U13312 (N_13312,N_13121,N_13166);
xor U13313 (N_13313,N_13188,N_13068);
nand U13314 (N_13314,N_13083,N_13002);
and U13315 (N_13315,N_13040,N_13129);
or U13316 (N_13316,N_13081,N_13139);
nand U13317 (N_13317,N_13043,N_13141);
xor U13318 (N_13318,N_13021,N_13041);
xor U13319 (N_13319,N_13161,N_13062);
xnor U13320 (N_13320,N_13041,N_13075);
nor U13321 (N_13321,N_13086,N_13072);
nand U13322 (N_13322,N_13158,N_13054);
nor U13323 (N_13323,N_13165,N_13008);
nand U13324 (N_13324,N_13109,N_13180);
or U13325 (N_13325,N_13152,N_13041);
and U13326 (N_13326,N_13009,N_13188);
nor U13327 (N_13327,N_13029,N_13149);
nand U13328 (N_13328,N_13101,N_13087);
or U13329 (N_13329,N_13047,N_13114);
nand U13330 (N_13330,N_13061,N_13145);
or U13331 (N_13331,N_13013,N_13083);
or U13332 (N_13332,N_13137,N_13032);
and U13333 (N_13333,N_13072,N_13116);
xnor U13334 (N_13334,N_13055,N_13026);
nor U13335 (N_13335,N_13196,N_13026);
or U13336 (N_13336,N_13156,N_13004);
or U13337 (N_13337,N_13057,N_13182);
or U13338 (N_13338,N_13008,N_13153);
or U13339 (N_13339,N_13144,N_13179);
or U13340 (N_13340,N_13083,N_13197);
nand U13341 (N_13341,N_13094,N_13103);
nor U13342 (N_13342,N_13013,N_13177);
nand U13343 (N_13343,N_13005,N_13185);
nand U13344 (N_13344,N_13122,N_13101);
nor U13345 (N_13345,N_13030,N_13077);
xor U13346 (N_13346,N_13096,N_13019);
xor U13347 (N_13347,N_13006,N_13044);
or U13348 (N_13348,N_13041,N_13088);
or U13349 (N_13349,N_13098,N_13130);
nand U13350 (N_13350,N_13073,N_13053);
and U13351 (N_13351,N_13067,N_13023);
and U13352 (N_13352,N_13050,N_13015);
xnor U13353 (N_13353,N_13082,N_13158);
xnor U13354 (N_13354,N_13093,N_13164);
nand U13355 (N_13355,N_13087,N_13045);
and U13356 (N_13356,N_13156,N_13006);
nor U13357 (N_13357,N_13153,N_13179);
and U13358 (N_13358,N_13109,N_13034);
or U13359 (N_13359,N_13147,N_13024);
xor U13360 (N_13360,N_13038,N_13179);
or U13361 (N_13361,N_13096,N_13100);
nand U13362 (N_13362,N_13101,N_13029);
nor U13363 (N_13363,N_13002,N_13035);
or U13364 (N_13364,N_13093,N_13003);
nor U13365 (N_13365,N_13184,N_13080);
nor U13366 (N_13366,N_13062,N_13013);
nand U13367 (N_13367,N_13191,N_13069);
xnor U13368 (N_13368,N_13181,N_13001);
nand U13369 (N_13369,N_13063,N_13013);
or U13370 (N_13370,N_13060,N_13062);
and U13371 (N_13371,N_13045,N_13199);
and U13372 (N_13372,N_13184,N_13098);
nor U13373 (N_13373,N_13033,N_13149);
xor U13374 (N_13374,N_13199,N_13109);
nor U13375 (N_13375,N_13020,N_13183);
nand U13376 (N_13376,N_13128,N_13147);
nor U13377 (N_13377,N_13010,N_13076);
nand U13378 (N_13378,N_13019,N_13172);
or U13379 (N_13379,N_13029,N_13121);
and U13380 (N_13380,N_13116,N_13134);
or U13381 (N_13381,N_13158,N_13053);
nor U13382 (N_13382,N_13048,N_13170);
nand U13383 (N_13383,N_13082,N_13020);
and U13384 (N_13384,N_13091,N_13011);
nand U13385 (N_13385,N_13064,N_13161);
and U13386 (N_13386,N_13048,N_13180);
nand U13387 (N_13387,N_13022,N_13081);
or U13388 (N_13388,N_13013,N_13030);
nor U13389 (N_13389,N_13097,N_13059);
and U13390 (N_13390,N_13021,N_13195);
xnor U13391 (N_13391,N_13190,N_13152);
nor U13392 (N_13392,N_13023,N_13097);
xor U13393 (N_13393,N_13059,N_13151);
or U13394 (N_13394,N_13181,N_13053);
and U13395 (N_13395,N_13186,N_13016);
or U13396 (N_13396,N_13144,N_13167);
or U13397 (N_13397,N_13006,N_13180);
nor U13398 (N_13398,N_13036,N_13142);
nor U13399 (N_13399,N_13179,N_13168);
nand U13400 (N_13400,N_13339,N_13212);
nor U13401 (N_13401,N_13273,N_13360);
xor U13402 (N_13402,N_13229,N_13261);
nor U13403 (N_13403,N_13393,N_13399);
and U13404 (N_13404,N_13363,N_13347);
xor U13405 (N_13405,N_13291,N_13263);
nand U13406 (N_13406,N_13293,N_13242);
and U13407 (N_13407,N_13377,N_13378);
nor U13408 (N_13408,N_13376,N_13221);
xor U13409 (N_13409,N_13231,N_13294);
xnor U13410 (N_13410,N_13201,N_13253);
nand U13411 (N_13411,N_13236,N_13310);
and U13412 (N_13412,N_13218,N_13353);
nor U13413 (N_13413,N_13292,N_13262);
nor U13414 (N_13414,N_13367,N_13256);
or U13415 (N_13415,N_13252,N_13316);
nand U13416 (N_13416,N_13366,N_13220);
or U13417 (N_13417,N_13286,N_13235);
nand U13418 (N_13418,N_13333,N_13359);
nand U13419 (N_13419,N_13223,N_13217);
or U13420 (N_13420,N_13375,N_13288);
or U13421 (N_13421,N_13248,N_13299);
or U13422 (N_13422,N_13207,N_13318);
nand U13423 (N_13423,N_13216,N_13264);
or U13424 (N_13424,N_13204,N_13249);
xor U13425 (N_13425,N_13331,N_13370);
nand U13426 (N_13426,N_13283,N_13228);
or U13427 (N_13427,N_13381,N_13372);
and U13428 (N_13428,N_13386,N_13319);
nor U13429 (N_13429,N_13308,N_13341);
xor U13430 (N_13430,N_13277,N_13224);
nand U13431 (N_13431,N_13227,N_13343);
and U13432 (N_13432,N_13361,N_13305);
nor U13433 (N_13433,N_13210,N_13285);
nand U13434 (N_13434,N_13374,N_13255);
xor U13435 (N_13435,N_13352,N_13321);
xor U13436 (N_13436,N_13320,N_13222);
nor U13437 (N_13437,N_13251,N_13245);
nor U13438 (N_13438,N_13358,N_13289);
and U13439 (N_13439,N_13274,N_13209);
nand U13440 (N_13440,N_13259,N_13270);
and U13441 (N_13441,N_13208,N_13284);
and U13442 (N_13442,N_13260,N_13240);
or U13443 (N_13443,N_13338,N_13392);
and U13444 (N_13444,N_13250,N_13297);
nor U13445 (N_13445,N_13272,N_13369);
xnor U13446 (N_13446,N_13247,N_13327);
xor U13447 (N_13447,N_13205,N_13267);
nor U13448 (N_13448,N_13282,N_13345);
nor U13449 (N_13449,N_13398,N_13281);
nor U13450 (N_13450,N_13233,N_13306);
xnor U13451 (N_13451,N_13239,N_13388);
nor U13452 (N_13452,N_13324,N_13258);
nand U13453 (N_13453,N_13389,N_13328);
and U13454 (N_13454,N_13332,N_13265);
nand U13455 (N_13455,N_13275,N_13266);
and U13456 (N_13456,N_13384,N_13203);
or U13457 (N_13457,N_13215,N_13200);
nand U13458 (N_13458,N_13295,N_13298);
and U13459 (N_13459,N_13241,N_13314);
or U13460 (N_13460,N_13350,N_13368);
or U13461 (N_13461,N_13391,N_13315);
xor U13462 (N_13462,N_13226,N_13271);
xnor U13463 (N_13463,N_13278,N_13257);
nand U13464 (N_13464,N_13354,N_13219);
and U13465 (N_13465,N_13355,N_13346);
nand U13466 (N_13466,N_13206,N_13351);
xnor U13467 (N_13467,N_13307,N_13385);
or U13468 (N_13468,N_13342,N_13357);
or U13469 (N_13469,N_13335,N_13337);
and U13470 (N_13470,N_13237,N_13234);
nor U13471 (N_13471,N_13243,N_13397);
nor U13472 (N_13472,N_13344,N_13287);
or U13473 (N_13473,N_13390,N_13323);
or U13474 (N_13474,N_13276,N_13396);
xor U13475 (N_13475,N_13312,N_13365);
nor U13476 (N_13476,N_13364,N_13225);
nand U13477 (N_13477,N_13371,N_13334);
and U13478 (N_13478,N_13395,N_13309);
and U13479 (N_13479,N_13211,N_13348);
xnor U13480 (N_13480,N_13254,N_13340);
and U13481 (N_13481,N_13296,N_13300);
and U13482 (N_13482,N_13246,N_13325);
nand U13483 (N_13483,N_13244,N_13379);
nor U13484 (N_13484,N_13387,N_13304);
and U13485 (N_13485,N_13301,N_13214);
and U13486 (N_13486,N_13317,N_13349);
or U13487 (N_13487,N_13329,N_13269);
xnor U13488 (N_13488,N_13322,N_13238);
xor U13489 (N_13489,N_13336,N_13362);
or U13490 (N_13490,N_13311,N_13394);
xnor U13491 (N_13491,N_13382,N_13202);
nand U13492 (N_13492,N_13380,N_13302);
or U13493 (N_13493,N_13303,N_13232);
and U13494 (N_13494,N_13383,N_13330);
xnor U13495 (N_13495,N_13230,N_13213);
or U13496 (N_13496,N_13373,N_13356);
or U13497 (N_13497,N_13279,N_13268);
and U13498 (N_13498,N_13280,N_13313);
xor U13499 (N_13499,N_13290,N_13326);
or U13500 (N_13500,N_13397,N_13231);
and U13501 (N_13501,N_13365,N_13379);
nor U13502 (N_13502,N_13255,N_13277);
or U13503 (N_13503,N_13210,N_13321);
or U13504 (N_13504,N_13310,N_13306);
or U13505 (N_13505,N_13362,N_13232);
xor U13506 (N_13506,N_13394,N_13341);
and U13507 (N_13507,N_13393,N_13228);
and U13508 (N_13508,N_13336,N_13315);
or U13509 (N_13509,N_13232,N_13384);
and U13510 (N_13510,N_13322,N_13320);
nand U13511 (N_13511,N_13251,N_13211);
nor U13512 (N_13512,N_13300,N_13291);
or U13513 (N_13513,N_13350,N_13247);
and U13514 (N_13514,N_13374,N_13273);
and U13515 (N_13515,N_13262,N_13316);
nor U13516 (N_13516,N_13386,N_13262);
xnor U13517 (N_13517,N_13208,N_13361);
xor U13518 (N_13518,N_13244,N_13391);
xor U13519 (N_13519,N_13261,N_13303);
and U13520 (N_13520,N_13352,N_13259);
or U13521 (N_13521,N_13265,N_13237);
or U13522 (N_13522,N_13377,N_13292);
nand U13523 (N_13523,N_13399,N_13349);
and U13524 (N_13524,N_13322,N_13351);
xnor U13525 (N_13525,N_13304,N_13389);
nand U13526 (N_13526,N_13393,N_13335);
nand U13527 (N_13527,N_13284,N_13292);
and U13528 (N_13528,N_13318,N_13371);
xnor U13529 (N_13529,N_13239,N_13307);
or U13530 (N_13530,N_13283,N_13243);
and U13531 (N_13531,N_13272,N_13301);
nor U13532 (N_13532,N_13382,N_13281);
nor U13533 (N_13533,N_13253,N_13237);
xnor U13534 (N_13534,N_13234,N_13312);
nand U13535 (N_13535,N_13266,N_13368);
nor U13536 (N_13536,N_13234,N_13212);
or U13537 (N_13537,N_13282,N_13289);
xor U13538 (N_13538,N_13364,N_13382);
and U13539 (N_13539,N_13384,N_13337);
and U13540 (N_13540,N_13319,N_13292);
nor U13541 (N_13541,N_13358,N_13336);
nor U13542 (N_13542,N_13367,N_13343);
or U13543 (N_13543,N_13268,N_13326);
nor U13544 (N_13544,N_13305,N_13300);
xnor U13545 (N_13545,N_13217,N_13209);
xor U13546 (N_13546,N_13314,N_13367);
nand U13547 (N_13547,N_13207,N_13337);
nor U13548 (N_13548,N_13234,N_13216);
and U13549 (N_13549,N_13273,N_13366);
or U13550 (N_13550,N_13397,N_13263);
and U13551 (N_13551,N_13340,N_13381);
nor U13552 (N_13552,N_13244,N_13388);
or U13553 (N_13553,N_13299,N_13258);
nor U13554 (N_13554,N_13391,N_13278);
nor U13555 (N_13555,N_13323,N_13214);
and U13556 (N_13556,N_13330,N_13372);
xnor U13557 (N_13557,N_13280,N_13329);
nand U13558 (N_13558,N_13324,N_13353);
nor U13559 (N_13559,N_13243,N_13336);
nand U13560 (N_13560,N_13320,N_13365);
xor U13561 (N_13561,N_13314,N_13216);
xor U13562 (N_13562,N_13284,N_13210);
nand U13563 (N_13563,N_13364,N_13297);
xnor U13564 (N_13564,N_13204,N_13202);
and U13565 (N_13565,N_13349,N_13388);
and U13566 (N_13566,N_13338,N_13303);
nor U13567 (N_13567,N_13311,N_13356);
xor U13568 (N_13568,N_13274,N_13386);
or U13569 (N_13569,N_13289,N_13216);
nor U13570 (N_13570,N_13345,N_13362);
and U13571 (N_13571,N_13354,N_13271);
nor U13572 (N_13572,N_13388,N_13264);
nor U13573 (N_13573,N_13392,N_13275);
or U13574 (N_13574,N_13374,N_13263);
nand U13575 (N_13575,N_13214,N_13384);
nor U13576 (N_13576,N_13345,N_13390);
and U13577 (N_13577,N_13214,N_13256);
nor U13578 (N_13578,N_13316,N_13366);
nor U13579 (N_13579,N_13296,N_13241);
and U13580 (N_13580,N_13390,N_13386);
nand U13581 (N_13581,N_13351,N_13318);
nand U13582 (N_13582,N_13366,N_13203);
xnor U13583 (N_13583,N_13279,N_13381);
and U13584 (N_13584,N_13349,N_13292);
or U13585 (N_13585,N_13293,N_13367);
nand U13586 (N_13586,N_13362,N_13281);
nand U13587 (N_13587,N_13259,N_13341);
nor U13588 (N_13588,N_13289,N_13384);
nor U13589 (N_13589,N_13290,N_13284);
xnor U13590 (N_13590,N_13342,N_13280);
nor U13591 (N_13591,N_13332,N_13399);
nand U13592 (N_13592,N_13348,N_13281);
and U13593 (N_13593,N_13243,N_13238);
xor U13594 (N_13594,N_13279,N_13311);
nor U13595 (N_13595,N_13333,N_13373);
nor U13596 (N_13596,N_13328,N_13237);
and U13597 (N_13597,N_13295,N_13281);
or U13598 (N_13598,N_13297,N_13304);
xnor U13599 (N_13599,N_13370,N_13384);
nand U13600 (N_13600,N_13515,N_13548);
nor U13601 (N_13601,N_13583,N_13563);
or U13602 (N_13602,N_13547,N_13592);
or U13603 (N_13603,N_13467,N_13407);
and U13604 (N_13604,N_13520,N_13527);
or U13605 (N_13605,N_13537,N_13517);
nand U13606 (N_13606,N_13492,N_13476);
or U13607 (N_13607,N_13509,N_13514);
and U13608 (N_13608,N_13420,N_13403);
or U13609 (N_13609,N_13469,N_13432);
xor U13610 (N_13610,N_13493,N_13594);
and U13611 (N_13611,N_13573,N_13513);
nand U13612 (N_13612,N_13512,N_13472);
or U13613 (N_13613,N_13498,N_13522);
nor U13614 (N_13614,N_13518,N_13506);
nand U13615 (N_13615,N_13541,N_13599);
and U13616 (N_13616,N_13598,N_13468);
and U13617 (N_13617,N_13443,N_13474);
and U13618 (N_13618,N_13505,N_13502);
nand U13619 (N_13619,N_13429,N_13544);
or U13620 (N_13620,N_13579,N_13508);
or U13621 (N_13621,N_13501,N_13442);
nor U13622 (N_13622,N_13570,N_13409);
xor U13623 (N_13623,N_13511,N_13595);
nand U13624 (N_13624,N_13435,N_13434);
nor U13625 (N_13625,N_13597,N_13414);
nand U13626 (N_13626,N_13559,N_13466);
nor U13627 (N_13627,N_13450,N_13452);
xnor U13628 (N_13628,N_13456,N_13567);
and U13629 (N_13629,N_13422,N_13487);
and U13630 (N_13630,N_13525,N_13484);
xnor U13631 (N_13631,N_13555,N_13480);
and U13632 (N_13632,N_13596,N_13556);
or U13633 (N_13633,N_13499,N_13489);
nor U13634 (N_13634,N_13451,N_13540);
and U13635 (N_13635,N_13551,N_13530);
nand U13636 (N_13636,N_13460,N_13523);
xnor U13637 (N_13637,N_13411,N_13496);
or U13638 (N_13638,N_13449,N_13459);
or U13639 (N_13639,N_13538,N_13528);
and U13640 (N_13640,N_13478,N_13533);
nor U13641 (N_13641,N_13462,N_13419);
nand U13642 (N_13642,N_13590,N_13486);
and U13643 (N_13643,N_13574,N_13457);
xnor U13644 (N_13644,N_13483,N_13539);
xor U13645 (N_13645,N_13562,N_13535);
xor U13646 (N_13646,N_13545,N_13529);
and U13647 (N_13647,N_13550,N_13446);
xnor U13648 (N_13648,N_13591,N_13582);
nand U13649 (N_13649,N_13497,N_13417);
and U13650 (N_13650,N_13471,N_13588);
nor U13651 (N_13651,N_13437,N_13448);
nor U13652 (N_13652,N_13561,N_13521);
nand U13653 (N_13653,N_13500,N_13586);
nor U13654 (N_13654,N_13477,N_13423);
nor U13655 (N_13655,N_13569,N_13461);
or U13656 (N_13656,N_13421,N_13571);
and U13657 (N_13657,N_13416,N_13589);
or U13658 (N_13658,N_13404,N_13475);
nor U13659 (N_13659,N_13464,N_13406);
nand U13660 (N_13660,N_13585,N_13433);
or U13661 (N_13661,N_13543,N_13482);
nand U13662 (N_13662,N_13441,N_13453);
nor U13663 (N_13663,N_13568,N_13572);
nor U13664 (N_13664,N_13454,N_13532);
xnor U13665 (N_13665,N_13410,N_13577);
xor U13666 (N_13666,N_13405,N_13425);
nand U13667 (N_13667,N_13536,N_13549);
nor U13668 (N_13668,N_13491,N_13408);
nor U13669 (N_13669,N_13495,N_13430);
nor U13670 (N_13670,N_13402,N_13488);
and U13671 (N_13671,N_13584,N_13439);
and U13672 (N_13672,N_13552,N_13415);
or U13673 (N_13673,N_13564,N_13560);
and U13674 (N_13674,N_13554,N_13566);
nand U13675 (N_13675,N_13581,N_13427);
or U13676 (N_13676,N_13445,N_13444);
and U13677 (N_13677,N_13401,N_13455);
or U13678 (N_13678,N_13526,N_13575);
and U13679 (N_13679,N_13542,N_13558);
or U13680 (N_13680,N_13470,N_13481);
nand U13681 (N_13681,N_13490,N_13447);
nor U13682 (N_13682,N_13458,N_13565);
and U13683 (N_13683,N_13438,N_13557);
xnor U13684 (N_13684,N_13440,N_13412);
nor U13685 (N_13685,N_13413,N_13428);
nor U13686 (N_13686,N_13426,N_13519);
or U13687 (N_13687,N_13576,N_13485);
xor U13688 (N_13688,N_13473,N_13510);
nand U13689 (N_13689,N_13593,N_13424);
nor U13690 (N_13690,N_13531,N_13546);
and U13691 (N_13691,N_13507,N_13431);
nand U13692 (N_13692,N_13534,N_13418);
nor U13693 (N_13693,N_13479,N_13580);
or U13694 (N_13694,N_13465,N_13494);
nand U13695 (N_13695,N_13516,N_13578);
xor U13696 (N_13696,N_13400,N_13463);
or U13697 (N_13697,N_13524,N_13587);
xor U13698 (N_13698,N_13553,N_13504);
and U13699 (N_13699,N_13436,N_13503);
nor U13700 (N_13700,N_13440,N_13537);
and U13701 (N_13701,N_13486,N_13425);
nor U13702 (N_13702,N_13506,N_13572);
nor U13703 (N_13703,N_13425,N_13550);
nand U13704 (N_13704,N_13556,N_13526);
nor U13705 (N_13705,N_13552,N_13419);
and U13706 (N_13706,N_13431,N_13549);
or U13707 (N_13707,N_13457,N_13502);
or U13708 (N_13708,N_13497,N_13462);
nor U13709 (N_13709,N_13553,N_13409);
xnor U13710 (N_13710,N_13462,N_13516);
or U13711 (N_13711,N_13485,N_13443);
xor U13712 (N_13712,N_13400,N_13531);
nand U13713 (N_13713,N_13414,N_13521);
nand U13714 (N_13714,N_13498,N_13573);
nor U13715 (N_13715,N_13474,N_13550);
xor U13716 (N_13716,N_13563,N_13407);
or U13717 (N_13717,N_13580,N_13520);
nor U13718 (N_13718,N_13523,N_13533);
nor U13719 (N_13719,N_13474,N_13597);
nand U13720 (N_13720,N_13596,N_13430);
or U13721 (N_13721,N_13425,N_13536);
xnor U13722 (N_13722,N_13440,N_13429);
nor U13723 (N_13723,N_13554,N_13591);
and U13724 (N_13724,N_13495,N_13477);
xnor U13725 (N_13725,N_13417,N_13415);
nor U13726 (N_13726,N_13566,N_13477);
xor U13727 (N_13727,N_13542,N_13537);
nor U13728 (N_13728,N_13596,N_13576);
nand U13729 (N_13729,N_13548,N_13465);
xnor U13730 (N_13730,N_13599,N_13415);
nand U13731 (N_13731,N_13416,N_13510);
or U13732 (N_13732,N_13543,N_13450);
nor U13733 (N_13733,N_13425,N_13539);
xnor U13734 (N_13734,N_13508,N_13400);
nor U13735 (N_13735,N_13570,N_13486);
nor U13736 (N_13736,N_13427,N_13504);
nand U13737 (N_13737,N_13454,N_13522);
nor U13738 (N_13738,N_13463,N_13516);
and U13739 (N_13739,N_13508,N_13541);
nand U13740 (N_13740,N_13416,N_13455);
and U13741 (N_13741,N_13510,N_13530);
and U13742 (N_13742,N_13512,N_13513);
or U13743 (N_13743,N_13584,N_13461);
xnor U13744 (N_13744,N_13493,N_13429);
nand U13745 (N_13745,N_13517,N_13598);
nand U13746 (N_13746,N_13580,N_13569);
or U13747 (N_13747,N_13413,N_13471);
xnor U13748 (N_13748,N_13403,N_13585);
and U13749 (N_13749,N_13463,N_13484);
or U13750 (N_13750,N_13443,N_13402);
nand U13751 (N_13751,N_13424,N_13420);
nor U13752 (N_13752,N_13495,N_13405);
nand U13753 (N_13753,N_13589,N_13442);
nor U13754 (N_13754,N_13531,N_13508);
xnor U13755 (N_13755,N_13426,N_13476);
xor U13756 (N_13756,N_13498,N_13428);
or U13757 (N_13757,N_13499,N_13564);
or U13758 (N_13758,N_13585,N_13410);
xnor U13759 (N_13759,N_13505,N_13448);
nor U13760 (N_13760,N_13529,N_13585);
or U13761 (N_13761,N_13556,N_13506);
and U13762 (N_13762,N_13417,N_13532);
nand U13763 (N_13763,N_13554,N_13469);
and U13764 (N_13764,N_13410,N_13502);
nand U13765 (N_13765,N_13533,N_13554);
or U13766 (N_13766,N_13422,N_13548);
xor U13767 (N_13767,N_13430,N_13438);
xnor U13768 (N_13768,N_13477,N_13470);
nor U13769 (N_13769,N_13542,N_13526);
or U13770 (N_13770,N_13418,N_13438);
nor U13771 (N_13771,N_13449,N_13445);
and U13772 (N_13772,N_13473,N_13509);
xor U13773 (N_13773,N_13542,N_13500);
and U13774 (N_13774,N_13594,N_13556);
nand U13775 (N_13775,N_13401,N_13523);
nor U13776 (N_13776,N_13471,N_13474);
nor U13777 (N_13777,N_13534,N_13487);
or U13778 (N_13778,N_13582,N_13515);
or U13779 (N_13779,N_13593,N_13498);
or U13780 (N_13780,N_13408,N_13422);
nand U13781 (N_13781,N_13505,N_13406);
and U13782 (N_13782,N_13566,N_13592);
or U13783 (N_13783,N_13569,N_13400);
xor U13784 (N_13784,N_13410,N_13504);
or U13785 (N_13785,N_13505,N_13536);
nand U13786 (N_13786,N_13441,N_13471);
nor U13787 (N_13787,N_13418,N_13424);
and U13788 (N_13788,N_13566,N_13486);
or U13789 (N_13789,N_13585,N_13540);
and U13790 (N_13790,N_13494,N_13538);
nor U13791 (N_13791,N_13403,N_13451);
nor U13792 (N_13792,N_13599,N_13445);
and U13793 (N_13793,N_13554,N_13439);
nand U13794 (N_13794,N_13560,N_13576);
nor U13795 (N_13795,N_13555,N_13485);
nor U13796 (N_13796,N_13532,N_13469);
nand U13797 (N_13797,N_13418,N_13421);
nor U13798 (N_13798,N_13466,N_13458);
nor U13799 (N_13799,N_13446,N_13402);
nand U13800 (N_13800,N_13760,N_13725);
nand U13801 (N_13801,N_13790,N_13716);
nor U13802 (N_13802,N_13612,N_13719);
xor U13803 (N_13803,N_13742,N_13770);
xor U13804 (N_13804,N_13767,N_13643);
or U13805 (N_13805,N_13667,N_13759);
and U13806 (N_13806,N_13700,N_13642);
nand U13807 (N_13807,N_13669,N_13785);
xnor U13808 (N_13808,N_13644,N_13679);
nor U13809 (N_13809,N_13798,N_13714);
nand U13810 (N_13810,N_13784,N_13633);
xor U13811 (N_13811,N_13608,N_13629);
nand U13812 (N_13812,N_13726,N_13634);
nor U13813 (N_13813,N_13752,N_13695);
nor U13814 (N_13814,N_13781,N_13645);
nand U13815 (N_13815,N_13748,N_13733);
nand U13816 (N_13816,N_13666,N_13706);
and U13817 (N_13817,N_13616,N_13604);
nand U13818 (N_13818,N_13722,N_13686);
nor U13819 (N_13819,N_13709,N_13736);
xnor U13820 (N_13820,N_13731,N_13796);
or U13821 (N_13821,N_13625,N_13793);
nor U13822 (N_13822,N_13647,N_13772);
nor U13823 (N_13823,N_13649,N_13693);
nand U13824 (N_13824,N_13658,N_13626);
nand U13825 (N_13825,N_13741,N_13628);
and U13826 (N_13826,N_13677,N_13680);
and U13827 (N_13827,N_13653,N_13678);
or U13828 (N_13828,N_13743,N_13690);
and U13829 (N_13829,N_13708,N_13755);
and U13830 (N_13830,N_13768,N_13681);
or U13831 (N_13831,N_13664,N_13746);
nand U13832 (N_13832,N_13799,N_13747);
xnor U13833 (N_13833,N_13648,N_13766);
and U13834 (N_13834,N_13623,N_13756);
or U13835 (N_13835,N_13780,N_13704);
nor U13836 (N_13836,N_13745,N_13650);
or U13837 (N_13837,N_13638,N_13788);
and U13838 (N_13838,N_13603,N_13710);
nand U13839 (N_13839,N_13783,N_13778);
xor U13840 (N_13840,N_13791,N_13620);
nand U13841 (N_13841,N_13771,N_13663);
nand U13842 (N_13842,N_13734,N_13671);
nor U13843 (N_13843,N_13676,N_13682);
or U13844 (N_13844,N_13773,N_13737);
and U13845 (N_13845,N_13674,N_13769);
nand U13846 (N_13846,N_13735,N_13703);
or U13847 (N_13847,N_13684,N_13758);
and U13848 (N_13848,N_13786,N_13635);
and U13849 (N_13849,N_13740,N_13609);
or U13850 (N_13850,N_13797,N_13683);
xor U13851 (N_13851,N_13654,N_13673);
xor U13852 (N_13852,N_13662,N_13622);
or U13853 (N_13853,N_13611,N_13613);
xor U13854 (N_13854,N_13665,N_13640);
xnor U13855 (N_13855,N_13765,N_13692);
or U13856 (N_13856,N_13723,N_13761);
and U13857 (N_13857,N_13792,N_13621);
nor U13858 (N_13858,N_13721,N_13701);
nor U13859 (N_13859,N_13659,N_13729);
or U13860 (N_13860,N_13685,N_13661);
nand U13861 (N_13861,N_13689,N_13672);
xnor U13862 (N_13862,N_13787,N_13660);
xnor U13863 (N_13863,N_13618,N_13631);
xor U13864 (N_13864,N_13606,N_13641);
nand U13865 (N_13865,N_13627,N_13774);
and U13866 (N_13866,N_13712,N_13789);
xnor U13867 (N_13867,N_13657,N_13637);
nand U13868 (N_13868,N_13764,N_13615);
xnor U13869 (N_13869,N_13750,N_13711);
xor U13870 (N_13870,N_13795,N_13697);
and U13871 (N_13871,N_13757,N_13738);
xor U13872 (N_13872,N_13718,N_13610);
and U13873 (N_13873,N_13698,N_13688);
nand U13874 (N_13874,N_13632,N_13702);
or U13875 (N_13875,N_13646,N_13724);
nor U13876 (N_13876,N_13600,N_13687);
nand U13877 (N_13877,N_13730,N_13668);
xnor U13878 (N_13878,N_13744,N_13636);
xnor U13879 (N_13879,N_13776,N_13762);
nor U13880 (N_13880,N_13670,N_13619);
xor U13881 (N_13881,N_13732,N_13777);
xnor U13882 (N_13882,N_13630,N_13779);
or U13883 (N_13883,N_13602,N_13720);
and U13884 (N_13884,N_13694,N_13775);
and U13885 (N_13885,N_13624,N_13754);
nand U13886 (N_13886,N_13751,N_13705);
xor U13887 (N_13887,N_13617,N_13607);
nor U13888 (N_13888,N_13691,N_13656);
nor U13889 (N_13889,N_13717,N_13639);
nand U13890 (N_13890,N_13675,N_13651);
nor U13891 (N_13891,N_13601,N_13605);
nand U13892 (N_13892,N_13739,N_13727);
xnor U13893 (N_13893,N_13655,N_13763);
nand U13894 (N_13894,N_13696,N_13753);
nand U13895 (N_13895,N_13699,N_13794);
xnor U13896 (N_13896,N_13782,N_13749);
nor U13897 (N_13897,N_13707,N_13614);
xnor U13898 (N_13898,N_13715,N_13652);
and U13899 (N_13899,N_13728,N_13713);
xnor U13900 (N_13900,N_13727,N_13780);
or U13901 (N_13901,N_13752,N_13742);
nand U13902 (N_13902,N_13714,N_13753);
xnor U13903 (N_13903,N_13653,N_13667);
nor U13904 (N_13904,N_13680,N_13604);
nand U13905 (N_13905,N_13609,N_13663);
xnor U13906 (N_13906,N_13697,N_13671);
xor U13907 (N_13907,N_13759,N_13792);
nand U13908 (N_13908,N_13715,N_13765);
xnor U13909 (N_13909,N_13614,N_13709);
and U13910 (N_13910,N_13687,N_13653);
xnor U13911 (N_13911,N_13632,N_13676);
nor U13912 (N_13912,N_13630,N_13747);
or U13913 (N_13913,N_13646,N_13756);
xor U13914 (N_13914,N_13777,N_13689);
nor U13915 (N_13915,N_13686,N_13757);
or U13916 (N_13916,N_13679,N_13670);
and U13917 (N_13917,N_13784,N_13772);
and U13918 (N_13918,N_13750,N_13626);
xor U13919 (N_13919,N_13771,N_13730);
and U13920 (N_13920,N_13685,N_13611);
and U13921 (N_13921,N_13639,N_13663);
xnor U13922 (N_13922,N_13779,N_13681);
xor U13923 (N_13923,N_13607,N_13624);
nor U13924 (N_13924,N_13698,N_13779);
and U13925 (N_13925,N_13679,N_13735);
and U13926 (N_13926,N_13606,N_13609);
nor U13927 (N_13927,N_13652,N_13641);
or U13928 (N_13928,N_13676,N_13770);
and U13929 (N_13929,N_13721,N_13739);
nand U13930 (N_13930,N_13617,N_13659);
nand U13931 (N_13931,N_13714,N_13602);
or U13932 (N_13932,N_13670,N_13748);
nor U13933 (N_13933,N_13691,N_13724);
nor U13934 (N_13934,N_13647,N_13724);
nor U13935 (N_13935,N_13632,N_13759);
xor U13936 (N_13936,N_13610,N_13637);
nand U13937 (N_13937,N_13738,N_13775);
xnor U13938 (N_13938,N_13639,N_13786);
and U13939 (N_13939,N_13744,N_13619);
and U13940 (N_13940,N_13624,N_13733);
and U13941 (N_13941,N_13749,N_13654);
xnor U13942 (N_13942,N_13791,N_13676);
nor U13943 (N_13943,N_13670,N_13676);
and U13944 (N_13944,N_13719,N_13758);
and U13945 (N_13945,N_13650,N_13776);
nor U13946 (N_13946,N_13612,N_13661);
nor U13947 (N_13947,N_13706,N_13606);
and U13948 (N_13948,N_13648,N_13771);
or U13949 (N_13949,N_13680,N_13693);
or U13950 (N_13950,N_13628,N_13712);
or U13951 (N_13951,N_13603,N_13707);
and U13952 (N_13952,N_13689,N_13791);
and U13953 (N_13953,N_13633,N_13767);
xnor U13954 (N_13954,N_13692,N_13655);
nand U13955 (N_13955,N_13618,N_13689);
xor U13956 (N_13956,N_13686,N_13786);
nor U13957 (N_13957,N_13689,N_13638);
nor U13958 (N_13958,N_13687,N_13633);
nor U13959 (N_13959,N_13799,N_13655);
nor U13960 (N_13960,N_13685,N_13797);
nand U13961 (N_13961,N_13621,N_13645);
and U13962 (N_13962,N_13633,N_13638);
or U13963 (N_13963,N_13739,N_13617);
and U13964 (N_13964,N_13792,N_13614);
or U13965 (N_13965,N_13645,N_13768);
xor U13966 (N_13966,N_13648,N_13695);
xor U13967 (N_13967,N_13657,N_13799);
xor U13968 (N_13968,N_13719,N_13600);
nand U13969 (N_13969,N_13753,N_13717);
and U13970 (N_13970,N_13775,N_13782);
and U13971 (N_13971,N_13759,N_13633);
nand U13972 (N_13972,N_13604,N_13606);
nand U13973 (N_13973,N_13706,N_13742);
and U13974 (N_13974,N_13698,N_13742);
nand U13975 (N_13975,N_13710,N_13709);
xor U13976 (N_13976,N_13729,N_13769);
nor U13977 (N_13977,N_13645,N_13766);
nor U13978 (N_13978,N_13781,N_13720);
and U13979 (N_13979,N_13735,N_13762);
xor U13980 (N_13980,N_13793,N_13784);
xnor U13981 (N_13981,N_13748,N_13799);
xor U13982 (N_13982,N_13735,N_13625);
nand U13983 (N_13983,N_13676,N_13608);
or U13984 (N_13984,N_13773,N_13641);
xor U13985 (N_13985,N_13715,N_13795);
nor U13986 (N_13986,N_13764,N_13675);
nand U13987 (N_13987,N_13691,N_13701);
or U13988 (N_13988,N_13767,N_13600);
xor U13989 (N_13989,N_13732,N_13653);
nor U13990 (N_13990,N_13718,N_13673);
xor U13991 (N_13991,N_13636,N_13651);
or U13992 (N_13992,N_13625,N_13643);
or U13993 (N_13993,N_13613,N_13602);
or U13994 (N_13994,N_13699,N_13781);
xor U13995 (N_13995,N_13785,N_13759);
or U13996 (N_13996,N_13752,N_13628);
or U13997 (N_13997,N_13744,N_13695);
xnor U13998 (N_13998,N_13642,N_13779);
xnor U13999 (N_13999,N_13627,N_13733);
nor U14000 (N_14000,N_13825,N_13910);
xor U14001 (N_14001,N_13943,N_13922);
nand U14002 (N_14002,N_13934,N_13906);
or U14003 (N_14003,N_13917,N_13974);
nand U14004 (N_14004,N_13975,N_13959);
nor U14005 (N_14005,N_13942,N_13815);
nor U14006 (N_14006,N_13872,N_13987);
nor U14007 (N_14007,N_13938,N_13805);
nor U14008 (N_14008,N_13864,N_13903);
xnor U14009 (N_14009,N_13929,N_13931);
nand U14010 (N_14010,N_13892,N_13822);
xnor U14011 (N_14011,N_13996,N_13867);
nor U14012 (N_14012,N_13842,N_13871);
and U14013 (N_14013,N_13961,N_13878);
nand U14014 (N_14014,N_13868,N_13880);
or U14015 (N_14015,N_13849,N_13951);
xor U14016 (N_14016,N_13851,N_13828);
xnor U14017 (N_14017,N_13809,N_13870);
or U14018 (N_14018,N_13863,N_13835);
xor U14019 (N_14019,N_13887,N_13855);
nand U14020 (N_14020,N_13821,N_13995);
or U14021 (N_14021,N_13832,N_13891);
or U14022 (N_14022,N_13981,N_13955);
nor U14023 (N_14023,N_13911,N_13806);
xnor U14024 (N_14024,N_13904,N_13896);
or U14025 (N_14025,N_13920,N_13834);
nor U14026 (N_14026,N_13944,N_13950);
nand U14027 (N_14027,N_13889,N_13823);
or U14028 (N_14028,N_13883,N_13977);
nand U14029 (N_14029,N_13893,N_13853);
nor U14030 (N_14030,N_13994,N_13940);
nor U14031 (N_14031,N_13845,N_13901);
xnor U14032 (N_14032,N_13965,N_13972);
and U14033 (N_14033,N_13874,N_13916);
nor U14034 (N_14034,N_13984,N_13895);
nand U14035 (N_14035,N_13949,N_13924);
xor U14036 (N_14036,N_13927,N_13860);
and U14037 (N_14037,N_13824,N_13812);
and U14038 (N_14038,N_13861,N_13939);
or U14039 (N_14039,N_13915,N_13960);
and U14040 (N_14040,N_13902,N_13877);
and U14041 (N_14041,N_13964,N_13914);
and U14042 (N_14042,N_13847,N_13808);
and U14043 (N_14043,N_13999,N_13813);
or U14044 (N_14044,N_13881,N_13919);
nor U14045 (N_14045,N_13963,N_13869);
nor U14046 (N_14046,N_13801,N_13804);
or U14047 (N_14047,N_13894,N_13875);
or U14048 (N_14048,N_13907,N_13876);
nand U14049 (N_14049,N_13856,N_13852);
or U14050 (N_14050,N_13811,N_13800);
nor U14051 (N_14051,N_13831,N_13935);
and U14052 (N_14052,N_13958,N_13971);
or U14053 (N_14053,N_13836,N_13978);
or U14054 (N_14054,N_13865,N_13839);
or U14055 (N_14055,N_13820,N_13854);
or U14056 (N_14056,N_13802,N_13862);
and U14057 (N_14057,N_13945,N_13866);
nand U14058 (N_14058,N_13918,N_13885);
nand U14059 (N_14059,N_13969,N_13946);
or U14060 (N_14060,N_13898,N_13843);
nor U14061 (N_14061,N_13956,N_13816);
nand U14062 (N_14062,N_13980,N_13970);
xnor U14063 (N_14063,N_13957,N_13810);
or U14064 (N_14064,N_13899,N_13827);
xnor U14065 (N_14065,N_13953,N_13982);
xnor U14066 (N_14066,N_13993,N_13879);
nand U14067 (N_14067,N_13859,N_13841);
nor U14068 (N_14068,N_13826,N_13905);
and U14069 (N_14069,N_13846,N_13992);
nand U14070 (N_14070,N_13890,N_13986);
and U14071 (N_14071,N_13967,N_13807);
and U14072 (N_14072,N_13913,N_13998);
or U14073 (N_14073,N_13858,N_13844);
or U14074 (N_14074,N_13928,N_13988);
nor U14075 (N_14075,N_13990,N_13897);
xor U14076 (N_14076,N_13968,N_13962);
nor U14077 (N_14077,N_13830,N_13973);
nor U14078 (N_14078,N_13803,N_13948);
nand U14079 (N_14079,N_13900,N_13840);
nand U14080 (N_14080,N_13884,N_13936);
or U14081 (N_14081,N_13912,N_13925);
nand U14082 (N_14082,N_13985,N_13882);
nand U14083 (N_14083,N_13923,N_13833);
xor U14084 (N_14084,N_13908,N_13850);
nand U14085 (N_14085,N_13966,N_13997);
nor U14086 (N_14086,N_13983,N_13930);
and U14087 (N_14087,N_13837,N_13932);
and U14088 (N_14088,N_13829,N_13989);
xor U14089 (N_14089,N_13873,N_13976);
nand U14090 (N_14090,N_13921,N_13886);
xnor U14091 (N_14091,N_13819,N_13909);
or U14092 (N_14092,N_13947,N_13857);
xnor U14093 (N_14093,N_13818,N_13817);
or U14094 (N_14094,N_13979,N_13937);
nor U14095 (N_14095,N_13941,N_13991);
nand U14096 (N_14096,N_13848,N_13926);
xor U14097 (N_14097,N_13954,N_13933);
nor U14098 (N_14098,N_13838,N_13952);
or U14099 (N_14099,N_13888,N_13814);
or U14100 (N_14100,N_13906,N_13942);
and U14101 (N_14101,N_13812,N_13864);
and U14102 (N_14102,N_13890,N_13940);
xnor U14103 (N_14103,N_13974,N_13916);
xnor U14104 (N_14104,N_13821,N_13814);
nor U14105 (N_14105,N_13932,N_13936);
nor U14106 (N_14106,N_13966,N_13808);
or U14107 (N_14107,N_13911,N_13803);
xor U14108 (N_14108,N_13922,N_13915);
or U14109 (N_14109,N_13840,N_13868);
nor U14110 (N_14110,N_13847,N_13830);
nand U14111 (N_14111,N_13889,N_13873);
nand U14112 (N_14112,N_13942,N_13946);
or U14113 (N_14113,N_13800,N_13995);
or U14114 (N_14114,N_13871,N_13917);
and U14115 (N_14115,N_13987,N_13975);
xnor U14116 (N_14116,N_13871,N_13839);
or U14117 (N_14117,N_13978,N_13926);
nand U14118 (N_14118,N_13924,N_13876);
or U14119 (N_14119,N_13825,N_13940);
or U14120 (N_14120,N_13969,N_13871);
nand U14121 (N_14121,N_13953,N_13963);
and U14122 (N_14122,N_13844,N_13940);
xnor U14123 (N_14123,N_13929,N_13878);
nand U14124 (N_14124,N_13817,N_13931);
xor U14125 (N_14125,N_13908,N_13991);
and U14126 (N_14126,N_13876,N_13980);
and U14127 (N_14127,N_13975,N_13876);
nand U14128 (N_14128,N_13837,N_13880);
nor U14129 (N_14129,N_13889,N_13931);
xnor U14130 (N_14130,N_13917,N_13904);
and U14131 (N_14131,N_13963,N_13922);
nand U14132 (N_14132,N_13850,N_13941);
or U14133 (N_14133,N_13910,N_13801);
and U14134 (N_14134,N_13881,N_13829);
xnor U14135 (N_14135,N_13938,N_13898);
nor U14136 (N_14136,N_13986,N_13926);
xor U14137 (N_14137,N_13882,N_13900);
and U14138 (N_14138,N_13978,N_13878);
nand U14139 (N_14139,N_13975,N_13823);
and U14140 (N_14140,N_13807,N_13856);
nand U14141 (N_14141,N_13874,N_13873);
nand U14142 (N_14142,N_13935,N_13940);
and U14143 (N_14143,N_13807,N_13867);
and U14144 (N_14144,N_13818,N_13898);
nor U14145 (N_14145,N_13871,N_13803);
nor U14146 (N_14146,N_13947,N_13829);
xor U14147 (N_14147,N_13832,N_13905);
or U14148 (N_14148,N_13965,N_13818);
nand U14149 (N_14149,N_13945,N_13890);
or U14150 (N_14150,N_13951,N_13839);
and U14151 (N_14151,N_13828,N_13834);
nor U14152 (N_14152,N_13970,N_13917);
xor U14153 (N_14153,N_13963,N_13841);
xnor U14154 (N_14154,N_13982,N_13956);
nand U14155 (N_14155,N_13920,N_13836);
or U14156 (N_14156,N_13910,N_13824);
or U14157 (N_14157,N_13814,N_13806);
and U14158 (N_14158,N_13952,N_13881);
nor U14159 (N_14159,N_13969,N_13825);
or U14160 (N_14160,N_13965,N_13953);
nor U14161 (N_14161,N_13876,N_13943);
and U14162 (N_14162,N_13818,N_13934);
or U14163 (N_14163,N_13937,N_13872);
xor U14164 (N_14164,N_13995,N_13999);
nand U14165 (N_14165,N_13952,N_13996);
nor U14166 (N_14166,N_13838,N_13828);
xor U14167 (N_14167,N_13879,N_13962);
xnor U14168 (N_14168,N_13935,N_13806);
or U14169 (N_14169,N_13989,N_13819);
or U14170 (N_14170,N_13962,N_13917);
or U14171 (N_14171,N_13985,N_13896);
xnor U14172 (N_14172,N_13844,N_13990);
nor U14173 (N_14173,N_13828,N_13940);
nor U14174 (N_14174,N_13832,N_13947);
xnor U14175 (N_14175,N_13885,N_13803);
and U14176 (N_14176,N_13881,N_13958);
nor U14177 (N_14177,N_13931,N_13863);
xor U14178 (N_14178,N_13847,N_13832);
xor U14179 (N_14179,N_13898,N_13915);
or U14180 (N_14180,N_13966,N_13957);
nand U14181 (N_14181,N_13986,N_13887);
xor U14182 (N_14182,N_13860,N_13982);
and U14183 (N_14183,N_13835,N_13903);
xor U14184 (N_14184,N_13974,N_13913);
xnor U14185 (N_14185,N_13966,N_13944);
nor U14186 (N_14186,N_13839,N_13941);
and U14187 (N_14187,N_13938,N_13822);
xor U14188 (N_14188,N_13967,N_13866);
and U14189 (N_14189,N_13960,N_13877);
or U14190 (N_14190,N_13967,N_13809);
and U14191 (N_14191,N_13863,N_13891);
xnor U14192 (N_14192,N_13932,N_13925);
nor U14193 (N_14193,N_13878,N_13849);
nor U14194 (N_14194,N_13814,N_13877);
nand U14195 (N_14195,N_13834,N_13849);
or U14196 (N_14196,N_13884,N_13845);
or U14197 (N_14197,N_13970,N_13816);
nor U14198 (N_14198,N_13811,N_13969);
xnor U14199 (N_14199,N_13942,N_13929);
nand U14200 (N_14200,N_14143,N_14146);
and U14201 (N_14201,N_14193,N_14161);
nand U14202 (N_14202,N_14113,N_14011);
or U14203 (N_14203,N_14179,N_14150);
nor U14204 (N_14204,N_14153,N_14010);
and U14205 (N_14205,N_14194,N_14196);
or U14206 (N_14206,N_14139,N_14170);
and U14207 (N_14207,N_14030,N_14026);
or U14208 (N_14208,N_14105,N_14035);
nand U14209 (N_14209,N_14068,N_14076);
and U14210 (N_14210,N_14132,N_14158);
or U14211 (N_14211,N_14195,N_14180);
xnor U14212 (N_14212,N_14122,N_14008);
and U14213 (N_14213,N_14007,N_14108);
xnor U14214 (N_14214,N_14014,N_14031);
and U14215 (N_14215,N_14072,N_14175);
and U14216 (N_14216,N_14156,N_14051);
nor U14217 (N_14217,N_14095,N_14097);
or U14218 (N_14218,N_14155,N_14100);
nand U14219 (N_14219,N_14082,N_14015);
or U14220 (N_14220,N_14021,N_14079);
nand U14221 (N_14221,N_14178,N_14002);
or U14222 (N_14222,N_14165,N_14020);
or U14223 (N_14223,N_14096,N_14001);
nor U14224 (N_14224,N_14157,N_14086);
nor U14225 (N_14225,N_14027,N_14053);
and U14226 (N_14226,N_14044,N_14177);
or U14227 (N_14227,N_14160,N_14118);
or U14228 (N_14228,N_14028,N_14070);
nand U14229 (N_14229,N_14092,N_14018);
and U14230 (N_14230,N_14109,N_14116);
nand U14231 (N_14231,N_14149,N_14163);
nor U14232 (N_14232,N_14059,N_14073);
nor U14233 (N_14233,N_14136,N_14060);
or U14234 (N_14234,N_14110,N_14087);
nor U14235 (N_14235,N_14058,N_14172);
or U14236 (N_14236,N_14084,N_14098);
or U14237 (N_14237,N_14111,N_14106);
nor U14238 (N_14238,N_14065,N_14046);
nor U14239 (N_14239,N_14140,N_14151);
or U14240 (N_14240,N_14071,N_14183);
xor U14241 (N_14241,N_14101,N_14089);
and U14242 (N_14242,N_14074,N_14012);
xor U14243 (N_14243,N_14174,N_14131);
xnor U14244 (N_14244,N_14091,N_14167);
or U14245 (N_14245,N_14077,N_14025);
nand U14246 (N_14246,N_14009,N_14123);
nand U14247 (N_14247,N_14085,N_14048);
or U14248 (N_14248,N_14016,N_14148);
and U14249 (N_14249,N_14152,N_14080);
and U14250 (N_14250,N_14003,N_14061);
nor U14251 (N_14251,N_14176,N_14164);
nor U14252 (N_14252,N_14188,N_14049);
xor U14253 (N_14253,N_14057,N_14173);
xnor U14254 (N_14254,N_14099,N_14038);
nand U14255 (N_14255,N_14128,N_14135);
xor U14256 (N_14256,N_14050,N_14024);
xnor U14257 (N_14257,N_14120,N_14137);
or U14258 (N_14258,N_14019,N_14119);
or U14259 (N_14259,N_14034,N_14181);
xor U14260 (N_14260,N_14088,N_14184);
xor U14261 (N_14261,N_14017,N_14117);
nand U14262 (N_14262,N_14121,N_14032);
or U14263 (N_14263,N_14067,N_14093);
or U14264 (N_14264,N_14166,N_14189);
xnor U14265 (N_14265,N_14129,N_14090);
or U14266 (N_14266,N_14125,N_14102);
and U14267 (N_14267,N_14199,N_14141);
nor U14268 (N_14268,N_14138,N_14124);
xnor U14269 (N_14269,N_14169,N_14022);
or U14270 (N_14270,N_14147,N_14043);
xor U14271 (N_14271,N_14168,N_14190);
nand U14272 (N_14272,N_14083,N_14039);
xnor U14273 (N_14273,N_14023,N_14197);
xor U14274 (N_14274,N_14130,N_14064);
nor U14275 (N_14275,N_14144,N_14006);
or U14276 (N_14276,N_14126,N_14115);
nand U14277 (N_14277,N_14052,N_14114);
or U14278 (N_14278,N_14191,N_14103);
nand U14279 (N_14279,N_14062,N_14094);
and U14280 (N_14280,N_14036,N_14133);
or U14281 (N_14281,N_14054,N_14004);
xor U14282 (N_14282,N_14005,N_14055);
nand U14283 (N_14283,N_14040,N_14187);
nand U14284 (N_14284,N_14142,N_14063);
nand U14285 (N_14285,N_14047,N_14075);
xnor U14286 (N_14286,N_14186,N_14045);
nand U14287 (N_14287,N_14033,N_14171);
or U14288 (N_14288,N_14037,N_14145);
nand U14289 (N_14289,N_14182,N_14107);
nor U14290 (N_14290,N_14192,N_14104);
and U14291 (N_14291,N_14081,N_14000);
and U14292 (N_14292,N_14162,N_14069);
nand U14293 (N_14293,N_14127,N_14134);
nand U14294 (N_14294,N_14029,N_14185);
xor U14295 (N_14295,N_14066,N_14159);
nand U14296 (N_14296,N_14042,N_14078);
nand U14297 (N_14297,N_14154,N_14112);
and U14298 (N_14298,N_14013,N_14198);
xor U14299 (N_14299,N_14056,N_14041);
nor U14300 (N_14300,N_14088,N_14189);
and U14301 (N_14301,N_14179,N_14146);
or U14302 (N_14302,N_14114,N_14112);
and U14303 (N_14303,N_14126,N_14055);
nand U14304 (N_14304,N_14173,N_14024);
nand U14305 (N_14305,N_14091,N_14180);
nand U14306 (N_14306,N_14114,N_14116);
and U14307 (N_14307,N_14197,N_14027);
xnor U14308 (N_14308,N_14173,N_14184);
nand U14309 (N_14309,N_14067,N_14152);
nand U14310 (N_14310,N_14127,N_14097);
or U14311 (N_14311,N_14160,N_14145);
and U14312 (N_14312,N_14111,N_14140);
nand U14313 (N_14313,N_14008,N_14019);
and U14314 (N_14314,N_14170,N_14035);
or U14315 (N_14315,N_14177,N_14059);
xnor U14316 (N_14316,N_14157,N_14106);
or U14317 (N_14317,N_14114,N_14162);
nor U14318 (N_14318,N_14009,N_14138);
and U14319 (N_14319,N_14042,N_14125);
and U14320 (N_14320,N_14056,N_14125);
or U14321 (N_14321,N_14145,N_14147);
nor U14322 (N_14322,N_14094,N_14090);
or U14323 (N_14323,N_14056,N_14127);
or U14324 (N_14324,N_14138,N_14163);
nor U14325 (N_14325,N_14181,N_14015);
and U14326 (N_14326,N_14017,N_14034);
and U14327 (N_14327,N_14104,N_14169);
xor U14328 (N_14328,N_14146,N_14172);
nor U14329 (N_14329,N_14163,N_14170);
xnor U14330 (N_14330,N_14007,N_14063);
nor U14331 (N_14331,N_14194,N_14087);
and U14332 (N_14332,N_14049,N_14124);
and U14333 (N_14333,N_14108,N_14140);
xor U14334 (N_14334,N_14099,N_14148);
nor U14335 (N_14335,N_14126,N_14194);
nor U14336 (N_14336,N_14022,N_14104);
xor U14337 (N_14337,N_14042,N_14117);
or U14338 (N_14338,N_14053,N_14048);
or U14339 (N_14339,N_14170,N_14172);
or U14340 (N_14340,N_14078,N_14070);
xnor U14341 (N_14341,N_14070,N_14172);
nor U14342 (N_14342,N_14140,N_14073);
or U14343 (N_14343,N_14170,N_14155);
nor U14344 (N_14344,N_14081,N_14156);
and U14345 (N_14345,N_14057,N_14079);
and U14346 (N_14346,N_14017,N_14142);
nand U14347 (N_14347,N_14199,N_14191);
nor U14348 (N_14348,N_14151,N_14188);
nor U14349 (N_14349,N_14188,N_14182);
xor U14350 (N_14350,N_14029,N_14117);
xnor U14351 (N_14351,N_14019,N_14061);
nand U14352 (N_14352,N_14022,N_14187);
nor U14353 (N_14353,N_14128,N_14192);
nand U14354 (N_14354,N_14033,N_14054);
xor U14355 (N_14355,N_14041,N_14149);
and U14356 (N_14356,N_14095,N_14026);
xor U14357 (N_14357,N_14191,N_14018);
or U14358 (N_14358,N_14085,N_14004);
nor U14359 (N_14359,N_14138,N_14043);
or U14360 (N_14360,N_14183,N_14065);
nand U14361 (N_14361,N_14052,N_14010);
or U14362 (N_14362,N_14075,N_14063);
nand U14363 (N_14363,N_14072,N_14077);
nand U14364 (N_14364,N_14114,N_14164);
xnor U14365 (N_14365,N_14035,N_14185);
nor U14366 (N_14366,N_14085,N_14178);
nor U14367 (N_14367,N_14127,N_14148);
nand U14368 (N_14368,N_14035,N_14162);
and U14369 (N_14369,N_14117,N_14158);
nor U14370 (N_14370,N_14125,N_14111);
xnor U14371 (N_14371,N_14108,N_14122);
or U14372 (N_14372,N_14149,N_14091);
or U14373 (N_14373,N_14166,N_14132);
and U14374 (N_14374,N_14178,N_14016);
nor U14375 (N_14375,N_14166,N_14056);
nor U14376 (N_14376,N_14029,N_14033);
nand U14377 (N_14377,N_14045,N_14123);
or U14378 (N_14378,N_14015,N_14080);
xnor U14379 (N_14379,N_14091,N_14061);
xnor U14380 (N_14380,N_14003,N_14158);
nand U14381 (N_14381,N_14066,N_14056);
xor U14382 (N_14382,N_14199,N_14174);
nor U14383 (N_14383,N_14011,N_14048);
nor U14384 (N_14384,N_14123,N_14006);
or U14385 (N_14385,N_14199,N_14160);
nand U14386 (N_14386,N_14169,N_14085);
and U14387 (N_14387,N_14060,N_14009);
or U14388 (N_14388,N_14038,N_14186);
or U14389 (N_14389,N_14001,N_14117);
nand U14390 (N_14390,N_14067,N_14153);
xnor U14391 (N_14391,N_14108,N_14154);
nor U14392 (N_14392,N_14163,N_14166);
and U14393 (N_14393,N_14093,N_14170);
and U14394 (N_14394,N_14045,N_14003);
xnor U14395 (N_14395,N_14098,N_14184);
or U14396 (N_14396,N_14059,N_14064);
nand U14397 (N_14397,N_14146,N_14112);
and U14398 (N_14398,N_14146,N_14183);
nor U14399 (N_14399,N_14118,N_14154);
nor U14400 (N_14400,N_14394,N_14356);
and U14401 (N_14401,N_14368,N_14295);
xnor U14402 (N_14402,N_14333,N_14290);
and U14403 (N_14403,N_14375,N_14223);
nand U14404 (N_14404,N_14253,N_14244);
nand U14405 (N_14405,N_14396,N_14353);
and U14406 (N_14406,N_14322,N_14226);
or U14407 (N_14407,N_14267,N_14329);
xor U14408 (N_14408,N_14235,N_14330);
nand U14409 (N_14409,N_14385,N_14377);
xnor U14410 (N_14410,N_14337,N_14204);
nor U14411 (N_14411,N_14286,N_14374);
nand U14412 (N_14412,N_14276,N_14307);
or U14413 (N_14413,N_14380,N_14240);
xnor U14414 (N_14414,N_14263,N_14225);
or U14415 (N_14415,N_14316,N_14249);
xnor U14416 (N_14416,N_14345,N_14305);
or U14417 (N_14417,N_14291,N_14234);
and U14418 (N_14418,N_14216,N_14293);
xnor U14419 (N_14419,N_14268,N_14357);
nor U14420 (N_14420,N_14334,N_14231);
or U14421 (N_14421,N_14228,N_14261);
xor U14422 (N_14422,N_14362,N_14203);
nor U14423 (N_14423,N_14237,N_14217);
nand U14424 (N_14424,N_14210,N_14222);
nor U14425 (N_14425,N_14346,N_14221);
and U14426 (N_14426,N_14300,N_14298);
or U14427 (N_14427,N_14314,N_14215);
nor U14428 (N_14428,N_14227,N_14365);
or U14429 (N_14429,N_14370,N_14219);
or U14430 (N_14430,N_14369,N_14278);
or U14431 (N_14431,N_14259,N_14390);
nor U14432 (N_14432,N_14381,N_14304);
nor U14433 (N_14433,N_14342,N_14250);
nand U14434 (N_14434,N_14206,N_14399);
or U14435 (N_14435,N_14328,N_14306);
or U14436 (N_14436,N_14313,N_14326);
nor U14437 (N_14437,N_14245,N_14288);
nor U14438 (N_14438,N_14379,N_14323);
nand U14439 (N_14439,N_14281,N_14387);
xnor U14440 (N_14440,N_14280,N_14247);
or U14441 (N_14441,N_14277,N_14297);
or U14442 (N_14442,N_14287,N_14332);
nor U14443 (N_14443,N_14207,N_14208);
xnor U14444 (N_14444,N_14397,N_14335);
and U14445 (N_14445,N_14248,N_14376);
xor U14446 (N_14446,N_14309,N_14318);
nand U14447 (N_14447,N_14212,N_14378);
nand U14448 (N_14448,N_14275,N_14236);
and U14449 (N_14449,N_14200,N_14258);
xor U14450 (N_14450,N_14327,N_14325);
nand U14451 (N_14451,N_14270,N_14364);
xor U14452 (N_14452,N_14349,N_14324);
nand U14453 (N_14453,N_14283,N_14255);
nand U14454 (N_14454,N_14320,N_14229);
and U14455 (N_14455,N_14382,N_14285);
and U14456 (N_14456,N_14266,N_14232);
nand U14457 (N_14457,N_14395,N_14224);
xnor U14458 (N_14458,N_14384,N_14359);
and U14459 (N_14459,N_14254,N_14386);
and U14460 (N_14460,N_14372,N_14282);
nand U14461 (N_14461,N_14238,N_14319);
or U14462 (N_14462,N_14292,N_14284);
and U14463 (N_14463,N_14242,N_14302);
xor U14464 (N_14464,N_14312,N_14271);
nor U14465 (N_14465,N_14246,N_14347);
xor U14466 (N_14466,N_14398,N_14344);
or U14467 (N_14467,N_14256,N_14257);
or U14468 (N_14468,N_14252,N_14358);
nor U14469 (N_14469,N_14391,N_14388);
nor U14470 (N_14470,N_14363,N_14321);
or U14471 (N_14471,N_14354,N_14355);
and U14472 (N_14472,N_14243,N_14209);
nand U14473 (N_14473,N_14213,N_14274);
and U14474 (N_14474,N_14339,N_14299);
nor U14475 (N_14475,N_14220,N_14366);
nand U14476 (N_14476,N_14373,N_14211);
nand U14477 (N_14477,N_14301,N_14241);
and U14478 (N_14478,N_14340,N_14296);
or U14479 (N_14479,N_14294,N_14230);
nand U14480 (N_14480,N_14352,N_14205);
nor U14481 (N_14481,N_14289,N_14343);
and U14482 (N_14482,N_14361,N_14273);
and U14483 (N_14483,N_14239,N_14317);
nand U14484 (N_14484,N_14233,N_14311);
nand U14485 (N_14485,N_14279,N_14350);
nand U14486 (N_14486,N_14389,N_14310);
nor U14487 (N_14487,N_14315,N_14393);
nand U14488 (N_14488,N_14269,N_14341);
xnor U14489 (N_14489,N_14308,N_14202);
xor U14490 (N_14490,N_14264,N_14367);
nand U14491 (N_14491,N_14303,N_14383);
or U14492 (N_14492,N_14214,N_14218);
and U14493 (N_14493,N_14351,N_14260);
and U14494 (N_14494,N_14262,N_14272);
nand U14495 (N_14495,N_14336,N_14201);
and U14496 (N_14496,N_14348,N_14331);
xnor U14497 (N_14497,N_14360,N_14338);
or U14498 (N_14498,N_14371,N_14251);
or U14499 (N_14499,N_14392,N_14265);
nand U14500 (N_14500,N_14329,N_14370);
nor U14501 (N_14501,N_14390,N_14397);
nand U14502 (N_14502,N_14201,N_14242);
nand U14503 (N_14503,N_14355,N_14267);
xor U14504 (N_14504,N_14370,N_14232);
nand U14505 (N_14505,N_14355,N_14212);
and U14506 (N_14506,N_14246,N_14344);
xor U14507 (N_14507,N_14329,N_14365);
nor U14508 (N_14508,N_14359,N_14315);
nor U14509 (N_14509,N_14218,N_14233);
nor U14510 (N_14510,N_14387,N_14200);
or U14511 (N_14511,N_14399,N_14370);
nand U14512 (N_14512,N_14380,N_14332);
and U14513 (N_14513,N_14231,N_14206);
nor U14514 (N_14514,N_14218,N_14213);
nand U14515 (N_14515,N_14309,N_14287);
xor U14516 (N_14516,N_14223,N_14384);
or U14517 (N_14517,N_14321,N_14390);
and U14518 (N_14518,N_14222,N_14205);
and U14519 (N_14519,N_14241,N_14362);
and U14520 (N_14520,N_14289,N_14287);
nor U14521 (N_14521,N_14358,N_14298);
nand U14522 (N_14522,N_14375,N_14217);
and U14523 (N_14523,N_14307,N_14206);
nor U14524 (N_14524,N_14207,N_14320);
and U14525 (N_14525,N_14239,N_14237);
nor U14526 (N_14526,N_14203,N_14332);
nor U14527 (N_14527,N_14276,N_14384);
or U14528 (N_14528,N_14342,N_14387);
nand U14529 (N_14529,N_14378,N_14237);
nand U14530 (N_14530,N_14310,N_14293);
and U14531 (N_14531,N_14290,N_14241);
or U14532 (N_14532,N_14333,N_14268);
nand U14533 (N_14533,N_14215,N_14244);
and U14534 (N_14534,N_14262,N_14275);
and U14535 (N_14535,N_14228,N_14247);
nor U14536 (N_14536,N_14358,N_14349);
or U14537 (N_14537,N_14249,N_14271);
and U14538 (N_14538,N_14211,N_14245);
or U14539 (N_14539,N_14367,N_14342);
nand U14540 (N_14540,N_14202,N_14347);
nor U14541 (N_14541,N_14254,N_14387);
nor U14542 (N_14542,N_14272,N_14270);
xor U14543 (N_14543,N_14249,N_14272);
nand U14544 (N_14544,N_14262,N_14269);
xnor U14545 (N_14545,N_14209,N_14323);
nand U14546 (N_14546,N_14237,N_14320);
or U14547 (N_14547,N_14313,N_14323);
or U14548 (N_14548,N_14390,N_14200);
xor U14549 (N_14549,N_14317,N_14250);
and U14550 (N_14550,N_14210,N_14232);
or U14551 (N_14551,N_14228,N_14249);
and U14552 (N_14552,N_14284,N_14262);
nand U14553 (N_14553,N_14313,N_14201);
and U14554 (N_14554,N_14246,N_14225);
or U14555 (N_14555,N_14245,N_14316);
nand U14556 (N_14556,N_14338,N_14339);
nand U14557 (N_14557,N_14219,N_14309);
nor U14558 (N_14558,N_14292,N_14300);
or U14559 (N_14559,N_14274,N_14336);
and U14560 (N_14560,N_14207,N_14369);
nor U14561 (N_14561,N_14309,N_14201);
xnor U14562 (N_14562,N_14287,N_14268);
nor U14563 (N_14563,N_14271,N_14399);
and U14564 (N_14564,N_14321,N_14343);
nand U14565 (N_14565,N_14365,N_14213);
nand U14566 (N_14566,N_14388,N_14324);
xor U14567 (N_14567,N_14298,N_14383);
or U14568 (N_14568,N_14210,N_14331);
xor U14569 (N_14569,N_14397,N_14276);
xnor U14570 (N_14570,N_14230,N_14276);
nand U14571 (N_14571,N_14358,N_14369);
nand U14572 (N_14572,N_14271,N_14263);
and U14573 (N_14573,N_14246,N_14348);
or U14574 (N_14574,N_14325,N_14306);
nand U14575 (N_14575,N_14388,N_14297);
nand U14576 (N_14576,N_14350,N_14209);
and U14577 (N_14577,N_14264,N_14340);
nand U14578 (N_14578,N_14315,N_14294);
or U14579 (N_14579,N_14382,N_14243);
nor U14580 (N_14580,N_14270,N_14317);
and U14581 (N_14581,N_14346,N_14323);
xor U14582 (N_14582,N_14243,N_14344);
or U14583 (N_14583,N_14336,N_14378);
and U14584 (N_14584,N_14342,N_14307);
and U14585 (N_14585,N_14254,N_14338);
nand U14586 (N_14586,N_14383,N_14367);
or U14587 (N_14587,N_14342,N_14377);
and U14588 (N_14588,N_14371,N_14350);
nor U14589 (N_14589,N_14338,N_14207);
and U14590 (N_14590,N_14385,N_14222);
xnor U14591 (N_14591,N_14243,N_14273);
nor U14592 (N_14592,N_14216,N_14350);
nor U14593 (N_14593,N_14310,N_14372);
or U14594 (N_14594,N_14313,N_14234);
and U14595 (N_14595,N_14232,N_14378);
nor U14596 (N_14596,N_14289,N_14204);
nor U14597 (N_14597,N_14200,N_14364);
and U14598 (N_14598,N_14232,N_14227);
nand U14599 (N_14599,N_14264,N_14232);
nor U14600 (N_14600,N_14564,N_14494);
and U14601 (N_14601,N_14440,N_14505);
nor U14602 (N_14602,N_14421,N_14442);
xnor U14603 (N_14603,N_14575,N_14512);
nand U14604 (N_14604,N_14410,N_14450);
or U14605 (N_14605,N_14419,N_14490);
xnor U14606 (N_14606,N_14471,N_14425);
or U14607 (N_14607,N_14456,N_14547);
or U14608 (N_14608,N_14417,N_14412);
xor U14609 (N_14609,N_14488,N_14546);
xnor U14610 (N_14610,N_14508,N_14521);
nand U14611 (N_14611,N_14594,N_14593);
nor U14612 (N_14612,N_14481,N_14476);
nor U14613 (N_14613,N_14431,N_14441);
or U14614 (N_14614,N_14571,N_14407);
nand U14615 (N_14615,N_14543,N_14541);
nor U14616 (N_14616,N_14432,N_14578);
or U14617 (N_14617,N_14466,N_14592);
xnor U14618 (N_14618,N_14401,N_14573);
or U14619 (N_14619,N_14597,N_14402);
nor U14620 (N_14620,N_14428,N_14460);
nand U14621 (N_14621,N_14485,N_14523);
or U14622 (N_14622,N_14453,N_14411);
nand U14623 (N_14623,N_14409,N_14400);
and U14624 (N_14624,N_14538,N_14520);
nor U14625 (N_14625,N_14513,N_14550);
or U14626 (N_14626,N_14473,N_14534);
xor U14627 (N_14627,N_14530,N_14516);
nand U14628 (N_14628,N_14559,N_14536);
and U14629 (N_14629,N_14483,N_14581);
nor U14630 (N_14630,N_14415,N_14562);
and U14631 (N_14631,N_14438,N_14449);
nand U14632 (N_14632,N_14423,N_14542);
nand U14633 (N_14633,N_14586,N_14463);
or U14634 (N_14634,N_14405,N_14497);
nand U14635 (N_14635,N_14587,N_14489);
nand U14636 (N_14636,N_14548,N_14468);
and U14637 (N_14637,N_14580,N_14467);
or U14638 (N_14638,N_14435,N_14424);
nor U14639 (N_14639,N_14519,N_14566);
nor U14640 (N_14640,N_14452,N_14555);
and U14641 (N_14641,N_14461,N_14565);
xor U14642 (N_14642,N_14487,N_14444);
nand U14643 (N_14643,N_14585,N_14527);
and U14644 (N_14644,N_14591,N_14501);
or U14645 (N_14645,N_14579,N_14455);
or U14646 (N_14646,N_14525,N_14554);
nand U14647 (N_14647,N_14563,N_14574);
or U14648 (N_14648,N_14443,N_14598);
and U14649 (N_14649,N_14545,N_14504);
nor U14650 (N_14650,N_14569,N_14478);
xor U14651 (N_14651,N_14433,N_14493);
or U14652 (N_14652,N_14560,N_14552);
or U14653 (N_14653,N_14445,N_14499);
or U14654 (N_14654,N_14406,N_14526);
xnor U14655 (N_14655,N_14539,N_14517);
xor U14656 (N_14656,N_14568,N_14482);
and U14657 (N_14657,N_14522,N_14479);
or U14658 (N_14658,N_14510,N_14589);
and U14659 (N_14659,N_14414,N_14544);
nand U14660 (N_14660,N_14549,N_14426);
or U14661 (N_14661,N_14457,N_14459);
and U14662 (N_14662,N_14429,N_14469);
or U14663 (N_14663,N_14420,N_14439);
xnor U14664 (N_14664,N_14588,N_14533);
nor U14665 (N_14665,N_14599,N_14561);
xor U14666 (N_14666,N_14515,N_14447);
nor U14667 (N_14667,N_14422,N_14446);
nand U14668 (N_14668,N_14524,N_14430);
nor U14669 (N_14669,N_14413,N_14558);
nor U14670 (N_14670,N_14503,N_14458);
or U14671 (N_14671,N_14448,N_14496);
nor U14672 (N_14672,N_14436,N_14535);
nand U14673 (N_14673,N_14557,N_14480);
and U14674 (N_14674,N_14434,N_14492);
or U14675 (N_14675,N_14418,N_14511);
and U14676 (N_14676,N_14537,N_14470);
and U14677 (N_14677,N_14451,N_14403);
xor U14678 (N_14678,N_14408,N_14582);
nand U14679 (N_14679,N_14572,N_14491);
xor U14680 (N_14680,N_14454,N_14477);
and U14681 (N_14681,N_14509,N_14553);
nor U14682 (N_14682,N_14486,N_14529);
nand U14683 (N_14683,N_14500,N_14551);
or U14684 (N_14684,N_14576,N_14498);
xor U14685 (N_14685,N_14556,N_14518);
or U14686 (N_14686,N_14514,N_14570);
xor U14687 (N_14687,N_14528,N_14475);
nor U14688 (N_14688,N_14474,N_14495);
and U14689 (N_14689,N_14404,N_14567);
nor U14690 (N_14690,N_14506,N_14531);
nand U14691 (N_14691,N_14577,N_14502);
or U14692 (N_14692,N_14596,N_14507);
or U14693 (N_14693,N_14540,N_14465);
nand U14694 (N_14694,N_14472,N_14584);
or U14695 (N_14695,N_14427,N_14532);
or U14696 (N_14696,N_14416,N_14464);
nor U14697 (N_14697,N_14462,N_14595);
xor U14698 (N_14698,N_14583,N_14590);
nor U14699 (N_14699,N_14437,N_14484);
nand U14700 (N_14700,N_14563,N_14465);
or U14701 (N_14701,N_14476,N_14421);
nor U14702 (N_14702,N_14476,N_14550);
or U14703 (N_14703,N_14403,N_14561);
or U14704 (N_14704,N_14555,N_14432);
or U14705 (N_14705,N_14409,N_14520);
or U14706 (N_14706,N_14480,N_14469);
or U14707 (N_14707,N_14589,N_14468);
nor U14708 (N_14708,N_14583,N_14434);
or U14709 (N_14709,N_14572,N_14551);
xor U14710 (N_14710,N_14404,N_14415);
xnor U14711 (N_14711,N_14543,N_14418);
nand U14712 (N_14712,N_14513,N_14448);
or U14713 (N_14713,N_14504,N_14516);
nand U14714 (N_14714,N_14472,N_14554);
and U14715 (N_14715,N_14498,N_14590);
nor U14716 (N_14716,N_14521,N_14445);
xor U14717 (N_14717,N_14550,N_14459);
nor U14718 (N_14718,N_14555,N_14492);
xor U14719 (N_14719,N_14418,N_14479);
nor U14720 (N_14720,N_14489,N_14585);
and U14721 (N_14721,N_14514,N_14409);
xnor U14722 (N_14722,N_14418,N_14438);
or U14723 (N_14723,N_14554,N_14581);
xnor U14724 (N_14724,N_14431,N_14414);
and U14725 (N_14725,N_14560,N_14464);
or U14726 (N_14726,N_14505,N_14571);
and U14727 (N_14727,N_14473,N_14485);
or U14728 (N_14728,N_14426,N_14478);
or U14729 (N_14729,N_14546,N_14541);
xnor U14730 (N_14730,N_14412,N_14434);
or U14731 (N_14731,N_14541,N_14435);
nor U14732 (N_14732,N_14461,N_14429);
or U14733 (N_14733,N_14404,N_14560);
and U14734 (N_14734,N_14487,N_14513);
xnor U14735 (N_14735,N_14405,N_14585);
nand U14736 (N_14736,N_14451,N_14595);
or U14737 (N_14737,N_14416,N_14447);
and U14738 (N_14738,N_14438,N_14434);
nand U14739 (N_14739,N_14589,N_14530);
xor U14740 (N_14740,N_14416,N_14440);
nand U14741 (N_14741,N_14506,N_14543);
xor U14742 (N_14742,N_14504,N_14591);
and U14743 (N_14743,N_14581,N_14591);
nor U14744 (N_14744,N_14483,N_14403);
xnor U14745 (N_14745,N_14401,N_14470);
or U14746 (N_14746,N_14584,N_14548);
and U14747 (N_14747,N_14556,N_14408);
nand U14748 (N_14748,N_14445,N_14503);
xnor U14749 (N_14749,N_14431,N_14572);
or U14750 (N_14750,N_14483,N_14538);
or U14751 (N_14751,N_14425,N_14511);
and U14752 (N_14752,N_14439,N_14414);
nand U14753 (N_14753,N_14400,N_14441);
and U14754 (N_14754,N_14556,N_14502);
or U14755 (N_14755,N_14513,N_14489);
or U14756 (N_14756,N_14448,N_14575);
nor U14757 (N_14757,N_14405,N_14567);
and U14758 (N_14758,N_14556,N_14539);
or U14759 (N_14759,N_14571,N_14585);
and U14760 (N_14760,N_14429,N_14443);
xnor U14761 (N_14761,N_14519,N_14400);
nand U14762 (N_14762,N_14561,N_14425);
nor U14763 (N_14763,N_14475,N_14437);
xor U14764 (N_14764,N_14447,N_14476);
and U14765 (N_14765,N_14404,N_14553);
or U14766 (N_14766,N_14448,N_14447);
xnor U14767 (N_14767,N_14455,N_14448);
xnor U14768 (N_14768,N_14514,N_14480);
or U14769 (N_14769,N_14591,N_14416);
or U14770 (N_14770,N_14541,N_14530);
or U14771 (N_14771,N_14545,N_14585);
and U14772 (N_14772,N_14588,N_14465);
nor U14773 (N_14773,N_14539,N_14599);
or U14774 (N_14774,N_14405,N_14410);
xor U14775 (N_14775,N_14416,N_14483);
nand U14776 (N_14776,N_14485,N_14566);
xnor U14777 (N_14777,N_14491,N_14490);
and U14778 (N_14778,N_14531,N_14454);
or U14779 (N_14779,N_14481,N_14523);
nor U14780 (N_14780,N_14579,N_14440);
and U14781 (N_14781,N_14415,N_14454);
nand U14782 (N_14782,N_14538,N_14569);
nor U14783 (N_14783,N_14483,N_14458);
xor U14784 (N_14784,N_14518,N_14532);
or U14785 (N_14785,N_14599,N_14589);
or U14786 (N_14786,N_14467,N_14440);
and U14787 (N_14787,N_14534,N_14596);
xor U14788 (N_14788,N_14572,N_14535);
or U14789 (N_14789,N_14518,N_14585);
nor U14790 (N_14790,N_14408,N_14529);
nand U14791 (N_14791,N_14419,N_14410);
xnor U14792 (N_14792,N_14547,N_14525);
xnor U14793 (N_14793,N_14451,N_14444);
nor U14794 (N_14794,N_14586,N_14539);
or U14795 (N_14795,N_14562,N_14409);
nor U14796 (N_14796,N_14539,N_14519);
nor U14797 (N_14797,N_14446,N_14517);
xnor U14798 (N_14798,N_14457,N_14506);
and U14799 (N_14799,N_14560,N_14524);
nor U14800 (N_14800,N_14732,N_14683);
xor U14801 (N_14801,N_14630,N_14711);
nor U14802 (N_14802,N_14617,N_14627);
and U14803 (N_14803,N_14760,N_14784);
nor U14804 (N_14804,N_14748,N_14766);
and U14805 (N_14805,N_14753,N_14657);
and U14806 (N_14806,N_14684,N_14749);
and U14807 (N_14807,N_14704,N_14678);
or U14808 (N_14808,N_14738,N_14792);
nand U14809 (N_14809,N_14620,N_14687);
nor U14810 (N_14810,N_14779,N_14622);
nor U14811 (N_14811,N_14716,N_14680);
xnor U14812 (N_14812,N_14707,N_14718);
and U14813 (N_14813,N_14772,N_14747);
nand U14814 (N_14814,N_14626,N_14669);
nor U14815 (N_14815,N_14629,N_14603);
xnor U14816 (N_14816,N_14606,N_14673);
xnor U14817 (N_14817,N_14639,N_14795);
nor U14818 (N_14818,N_14650,N_14615);
and U14819 (N_14819,N_14758,N_14752);
and U14820 (N_14820,N_14782,N_14697);
nor U14821 (N_14821,N_14778,N_14663);
and U14822 (N_14822,N_14667,N_14636);
nand U14823 (N_14823,N_14654,N_14776);
xor U14824 (N_14824,N_14659,N_14698);
nand U14825 (N_14825,N_14668,N_14725);
and U14826 (N_14826,N_14709,N_14604);
or U14827 (N_14827,N_14655,N_14702);
nand U14828 (N_14828,N_14643,N_14767);
and U14829 (N_14829,N_14658,N_14641);
xor U14830 (N_14830,N_14787,N_14731);
or U14831 (N_14831,N_14780,N_14789);
and U14832 (N_14832,N_14605,N_14723);
nand U14833 (N_14833,N_14777,N_14773);
or U14834 (N_14834,N_14688,N_14715);
or U14835 (N_14835,N_14649,N_14693);
xnor U14836 (N_14836,N_14645,N_14610);
nand U14837 (N_14837,N_14638,N_14726);
nor U14838 (N_14838,N_14708,N_14700);
xor U14839 (N_14839,N_14652,N_14741);
or U14840 (N_14840,N_14679,N_14611);
xnor U14841 (N_14841,N_14646,N_14785);
or U14842 (N_14842,N_14637,N_14689);
xor U14843 (N_14843,N_14736,N_14794);
nand U14844 (N_14844,N_14665,N_14653);
and U14845 (N_14845,N_14607,N_14775);
xnor U14846 (N_14846,N_14694,N_14692);
nor U14847 (N_14847,N_14751,N_14737);
nor U14848 (N_14848,N_14757,N_14759);
nand U14849 (N_14849,N_14619,N_14633);
nor U14850 (N_14850,N_14632,N_14685);
nand U14851 (N_14851,N_14691,N_14635);
or U14852 (N_14852,N_14746,N_14722);
xnor U14853 (N_14853,N_14743,N_14786);
and U14854 (N_14854,N_14634,N_14733);
nand U14855 (N_14855,N_14656,N_14661);
and U14856 (N_14856,N_14642,N_14647);
and U14857 (N_14857,N_14706,N_14671);
or U14858 (N_14858,N_14769,N_14681);
and U14859 (N_14859,N_14625,N_14721);
and U14860 (N_14860,N_14601,N_14717);
xor U14861 (N_14861,N_14628,N_14799);
or U14862 (N_14862,N_14712,N_14768);
or U14863 (N_14863,N_14770,N_14763);
xor U14864 (N_14864,N_14695,N_14796);
xnor U14865 (N_14865,N_14613,N_14682);
or U14866 (N_14866,N_14745,N_14624);
and U14867 (N_14867,N_14616,N_14724);
or U14868 (N_14868,N_14674,N_14790);
and U14869 (N_14869,N_14644,N_14664);
or U14870 (N_14870,N_14612,N_14686);
nand U14871 (N_14871,N_14788,N_14609);
nor U14872 (N_14872,N_14705,N_14623);
xnor U14873 (N_14873,N_14740,N_14713);
or U14874 (N_14874,N_14774,N_14666);
or U14875 (N_14875,N_14648,N_14793);
or U14876 (N_14876,N_14640,N_14672);
or U14877 (N_14877,N_14734,N_14600);
nor U14878 (N_14878,N_14728,N_14703);
and U14879 (N_14879,N_14631,N_14727);
nor U14880 (N_14880,N_14755,N_14765);
nand U14881 (N_14881,N_14739,N_14730);
or U14882 (N_14882,N_14675,N_14742);
or U14883 (N_14883,N_14690,N_14735);
or U14884 (N_14884,N_14662,N_14791);
and U14885 (N_14885,N_14719,N_14602);
nand U14886 (N_14886,N_14677,N_14618);
and U14887 (N_14887,N_14754,N_14762);
nand U14888 (N_14888,N_14714,N_14750);
xor U14889 (N_14889,N_14710,N_14670);
or U14890 (N_14890,N_14651,N_14699);
and U14891 (N_14891,N_14720,N_14756);
xnor U14892 (N_14892,N_14798,N_14797);
and U14893 (N_14893,N_14783,N_14621);
or U14894 (N_14894,N_14744,N_14761);
nand U14895 (N_14895,N_14614,N_14608);
and U14896 (N_14896,N_14676,N_14701);
nor U14897 (N_14897,N_14660,N_14764);
or U14898 (N_14898,N_14781,N_14696);
xnor U14899 (N_14899,N_14771,N_14729);
nand U14900 (N_14900,N_14649,N_14617);
nor U14901 (N_14901,N_14620,N_14629);
nand U14902 (N_14902,N_14670,N_14725);
or U14903 (N_14903,N_14626,N_14786);
nor U14904 (N_14904,N_14715,N_14716);
xor U14905 (N_14905,N_14649,N_14715);
xnor U14906 (N_14906,N_14601,N_14701);
nand U14907 (N_14907,N_14711,N_14652);
or U14908 (N_14908,N_14770,N_14731);
nor U14909 (N_14909,N_14651,N_14613);
xor U14910 (N_14910,N_14796,N_14768);
nor U14911 (N_14911,N_14706,N_14769);
xnor U14912 (N_14912,N_14662,N_14616);
nor U14913 (N_14913,N_14728,N_14790);
nor U14914 (N_14914,N_14617,N_14670);
nand U14915 (N_14915,N_14706,N_14679);
nor U14916 (N_14916,N_14687,N_14728);
and U14917 (N_14917,N_14740,N_14731);
and U14918 (N_14918,N_14678,N_14755);
nor U14919 (N_14919,N_14729,N_14777);
and U14920 (N_14920,N_14661,N_14718);
xor U14921 (N_14921,N_14710,N_14688);
nor U14922 (N_14922,N_14600,N_14623);
nand U14923 (N_14923,N_14679,N_14796);
or U14924 (N_14924,N_14744,N_14607);
nand U14925 (N_14925,N_14651,N_14746);
nand U14926 (N_14926,N_14767,N_14704);
or U14927 (N_14927,N_14770,N_14784);
or U14928 (N_14928,N_14744,N_14692);
nand U14929 (N_14929,N_14613,N_14768);
xnor U14930 (N_14930,N_14630,N_14770);
or U14931 (N_14931,N_14647,N_14652);
and U14932 (N_14932,N_14781,N_14727);
and U14933 (N_14933,N_14615,N_14637);
or U14934 (N_14934,N_14686,N_14723);
or U14935 (N_14935,N_14685,N_14614);
nor U14936 (N_14936,N_14747,N_14637);
nand U14937 (N_14937,N_14794,N_14652);
xnor U14938 (N_14938,N_14628,N_14711);
and U14939 (N_14939,N_14684,N_14786);
or U14940 (N_14940,N_14674,N_14609);
nor U14941 (N_14941,N_14650,N_14610);
nand U14942 (N_14942,N_14763,N_14759);
or U14943 (N_14943,N_14640,N_14737);
or U14944 (N_14944,N_14656,N_14673);
nor U14945 (N_14945,N_14665,N_14613);
xor U14946 (N_14946,N_14644,N_14678);
nand U14947 (N_14947,N_14772,N_14665);
or U14948 (N_14948,N_14751,N_14765);
nand U14949 (N_14949,N_14662,N_14613);
xor U14950 (N_14950,N_14744,N_14631);
or U14951 (N_14951,N_14762,N_14721);
nand U14952 (N_14952,N_14718,N_14617);
nor U14953 (N_14953,N_14756,N_14620);
or U14954 (N_14954,N_14778,N_14792);
xor U14955 (N_14955,N_14782,N_14667);
and U14956 (N_14956,N_14712,N_14679);
xnor U14957 (N_14957,N_14759,N_14716);
nand U14958 (N_14958,N_14619,N_14641);
nand U14959 (N_14959,N_14745,N_14677);
nor U14960 (N_14960,N_14715,N_14653);
and U14961 (N_14961,N_14740,N_14704);
nor U14962 (N_14962,N_14789,N_14791);
or U14963 (N_14963,N_14697,N_14656);
and U14964 (N_14964,N_14663,N_14724);
and U14965 (N_14965,N_14756,N_14637);
nor U14966 (N_14966,N_14799,N_14765);
and U14967 (N_14967,N_14622,N_14680);
nor U14968 (N_14968,N_14612,N_14766);
or U14969 (N_14969,N_14726,N_14740);
and U14970 (N_14970,N_14703,N_14743);
nor U14971 (N_14971,N_14615,N_14619);
and U14972 (N_14972,N_14645,N_14743);
nand U14973 (N_14973,N_14757,N_14751);
nor U14974 (N_14974,N_14661,N_14638);
xnor U14975 (N_14975,N_14629,N_14740);
nor U14976 (N_14976,N_14719,N_14771);
xnor U14977 (N_14977,N_14782,N_14714);
nand U14978 (N_14978,N_14790,N_14623);
nand U14979 (N_14979,N_14736,N_14622);
nand U14980 (N_14980,N_14741,N_14650);
or U14981 (N_14981,N_14715,N_14767);
nand U14982 (N_14982,N_14650,N_14695);
xnor U14983 (N_14983,N_14614,N_14787);
xor U14984 (N_14984,N_14658,N_14799);
or U14985 (N_14985,N_14720,N_14678);
nand U14986 (N_14986,N_14737,N_14740);
and U14987 (N_14987,N_14640,N_14794);
or U14988 (N_14988,N_14731,N_14700);
or U14989 (N_14989,N_14665,N_14626);
nor U14990 (N_14990,N_14698,N_14616);
nand U14991 (N_14991,N_14654,N_14743);
nand U14992 (N_14992,N_14622,N_14791);
or U14993 (N_14993,N_14601,N_14600);
and U14994 (N_14994,N_14689,N_14666);
nor U14995 (N_14995,N_14644,N_14689);
nand U14996 (N_14996,N_14718,N_14758);
or U14997 (N_14997,N_14627,N_14638);
or U14998 (N_14998,N_14752,N_14763);
nor U14999 (N_14999,N_14696,N_14643);
nor U15000 (N_15000,N_14841,N_14804);
xor U15001 (N_15001,N_14884,N_14970);
nor U15002 (N_15002,N_14950,N_14948);
and U15003 (N_15003,N_14860,N_14941);
and U15004 (N_15004,N_14971,N_14988);
nor U15005 (N_15005,N_14832,N_14972);
and U15006 (N_15006,N_14815,N_14886);
and U15007 (N_15007,N_14842,N_14887);
xor U15008 (N_15008,N_14938,N_14836);
xnor U15009 (N_15009,N_14867,N_14866);
nand U15010 (N_15010,N_14831,N_14893);
xnor U15011 (N_15011,N_14837,N_14913);
or U15012 (N_15012,N_14964,N_14818);
and U15013 (N_15013,N_14924,N_14874);
xnor U15014 (N_15014,N_14931,N_14914);
xnor U15015 (N_15015,N_14888,N_14973);
and U15016 (N_15016,N_14822,N_14902);
nand U15017 (N_15017,N_14949,N_14813);
xor U15018 (N_15018,N_14922,N_14967);
xor U15019 (N_15019,N_14895,N_14909);
or U15020 (N_15020,N_14911,N_14805);
nor U15021 (N_15021,N_14863,N_14828);
nand U15022 (N_15022,N_14944,N_14963);
nand U15023 (N_15023,N_14891,N_14894);
nand U15024 (N_15024,N_14843,N_14977);
nand U15025 (N_15025,N_14984,N_14945);
and U15026 (N_15026,N_14932,N_14905);
nand U15027 (N_15027,N_14900,N_14845);
nor U15028 (N_15028,N_14985,N_14853);
xor U15029 (N_15029,N_14846,N_14904);
and U15030 (N_15030,N_14821,N_14835);
nand U15031 (N_15031,N_14961,N_14898);
and U15032 (N_15032,N_14890,N_14829);
nor U15033 (N_15033,N_14801,N_14864);
nor U15034 (N_15034,N_14879,N_14810);
or U15035 (N_15035,N_14875,N_14926);
nand U15036 (N_15036,N_14855,N_14889);
nor U15037 (N_15037,N_14965,N_14929);
nand U15038 (N_15038,N_14800,N_14915);
nor U15039 (N_15039,N_14910,N_14980);
and U15040 (N_15040,N_14998,N_14881);
nor U15041 (N_15041,N_14858,N_14999);
or U15042 (N_15042,N_14908,N_14856);
or U15043 (N_15043,N_14947,N_14877);
nand U15044 (N_15044,N_14943,N_14920);
xor U15045 (N_15045,N_14953,N_14921);
nor U15046 (N_15046,N_14834,N_14848);
nand U15047 (N_15047,N_14959,N_14820);
nor U15048 (N_15048,N_14859,N_14878);
nand U15049 (N_15049,N_14816,N_14951);
nand U15050 (N_15050,N_14954,N_14880);
and U15051 (N_15051,N_14826,N_14817);
nor U15052 (N_15052,N_14833,N_14897);
xor U15053 (N_15053,N_14814,N_14892);
nand U15054 (N_15054,N_14838,N_14987);
and U15055 (N_15055,N_14896,N_14823);
nand U15056 (N_15056,N_14839,N_14849);
and U15057 (N_15057,N_14871,N_14869);
xor U15058 (N_15058,N_14942,N_14882);
or U15059 (N_15059,N_14995,N_14937);
nand U15060 (N_15060,N_14803,N_14812);
and U15061 (N_15061,N_14997,N_14824);
xnor U15062 (N_15062,N_14940,N_14991);
or U15063 (N_15063,N_14806,N_14809);
and U15064 (N_15064,N_14907,N_14807);
nor U15065 (N_15065,N_14974,N_14919);
and U15066 (N_15066,N_14962,N_14851);
and U15067 (N_15067,N_14865,N_14982);
nand U15068 (N_15068,N_14957,N_14969);
nand U15069 (N_15069,N_14899,N_14830);
xor U15070 (N_15070,N_14936,N_14876);
and U15071 (N_15071,N_14811,N_14976);
nand U15072 (N_15072,N_14989,N_14872);
nor U15073 (N_15073,N_14935,N_14825);
xnor U15074 (N_15074,N_14960,N_14968);
nand U15075 (N_15075,N_14903,N_14994);
xor U15076 (N_15076,N_14983,N_14992);
nor U15077 (N_15077,N_14917,N_14990);
and U15078 (N_15078,N_14955,N_14981);
nand U15079 (N_15079,N_14912,N_14946);
or U15080 (N_15080,N_14808,N_14956);
nor U15081 (N_15081,N_14850,N_14934);
xor U15082 (N_15082,N_14870,N_14854);
nand U15083 (N_15083,N_14862,N_14802);
xor U15084 (N_15084,N_14901,N_14883);
and U15085 (N_15085,N_14916,N_14925);
or U15086 (N_15086,N_14939,N_14930);
nand U15087 (N_15087,N_14861,N_14986);
or U15088 (N_15088,N_14933,N_14996);
nand U15089 (N_15089,N_14885,N_14918);
or U15090 (N_15090,N_14844,N_14840);
and U15091 (N_15091,N_14975,N_14958);
xor U15092 (N_15092,N_14819,N_14906);
nor U15093 (N_15093,N_14852,N_14952);
nor U15094 (N_15094,N_14857,N_14827);
xor U15095 (N_15095,N_14928,N_14927);
nor U15096 (N_15096,N_14979,N_14923);
nand U15097 (N_15097,N_14847,N_14978);
nand U15098 (N_15098,N_14966,N_14868);
nor U15099 (N_15099,N_14873,N_14993);
or U15100 (N_15100,N_14856,N_14895);
xnor U15101 (N_15101,N_14814,N_14851);
or U15102 (N_15102,N_14821,N_14932);
xnor U15103 (N_15103,N_14905,N_14990);
nor U15104 (N_15104,N_14949,N_14830);
xor U15105 (N_15105,N_14877,N_14802);
and U15106 (N_15106,N_14874,N_14846);
xnor U15107 (N_15107,N_14871,N_14823);
nor U15108 (N_15108,N_14872,N_14825);
and U15109 (N_15109,N_14930,N_14800);
and U15110 (N_15110,N_14857,N_14833);
nor U15111 (N_15111,N_14834,N_14999);
xnor U15112 (N_15112,N_14862,N_14968);
xor U15113 (N_15113,N_14856,N_14934);
nor U15114 (N_15114,N_14932,N_14872);
or U15115 (N_15115,N_14884,N_14845);
and U15116 (N_15116,N_14868,N_14864);
or U15117 (N_15117,N_14998,N_14865);
and U15118 (N_15118,N_14853,N_14814);
and U15119 (N_15119,N_14974,N_14830);
nand U15120 (N_15120,N_14921,N_14896);
or U15121 (N_15121,N_14808,N_14899);
nor U15122 (N_15122,N_14881,N_14901);
xnor U15123 (N_15123,N_14861,N_14884);
nand U15124 (N_15124,N_14815,N_14805);
nor U15125 (N_15125,N_14982,N_14905);
xnor U15126 (N_15126,N_14898,N_14992);
and U15127 (N_15127,N_14930,N_14924);
xnor U15128 (N_15128,N_14925,N_14879);
nor U15129 (N_15129,N_14918,N_14942);
nor U15130 (N_15130,N_14957,N_14932);
xnor U15131 (N_15131,N_14979,N_14816);
or U15132 (N_15132,N_14837,N_14936);
or U15133 (N_15133,N_14883,N_14960);
nand U15134 (N_15134,N_14937,N_14900);
or U15135 (N_15135,N_14873,N_14810);
nand U15136 (N_15136,N_14877,N_14985);
or U15137 (N_15137,N_14974,N_14998);
and U15138 (N_15138,N_14936,N_14992);
and U15139 (N_15139,N_14892,N_14947);
nand U15140 (N_15140,N_14924,N_14945);
nor U15141 (N_15141,N_14941,N_14997);
and U15142 (N_15142,N_14839,N_14809);
or U15143 (N_15143,N_14953,N_14959);
or U15144 (N_15144,N_14969,N_14937);
nand U15145 (N_15145,N_14956,N_14854);
xnor U15146 (N_15146,N_14919,N_14912);
xnor U15147 (N_15147,N_14924,N_14828);
nor U15148 (N_15148,N_14964,N_14963);
or U15149 (N_15149,N_14811,N_14951);
xor U15150 (N_15150,N_14985,N_14959);
nor U15151 (N_15151,N_14825,N_14936);
nor U15152 (N_15152,N_14881,N_14904);
nor U15153 (N_15153,N_14829,N_14977);
xnor U15154 (N_15154,N_14808,N_14945);
and U15155 (N_15155,N_14964,N_14980);
xor U15156 (N_15156,N_14876,N_14976);
xor U15157 (N_15157,N_14849,N_14892);
xnor U15158 (N_15158,N_14891,N_14918);
nor U15159 (N_15159,N_14931,N_14890);
and U15160 (N_15160,N_14987,N_14904);
xnor U15161 (N_15161,N_14850,N_14856);
xnor U15162 (N_15162,N_14884,N_14915);
or U15163 (N_15163,N_14926,N_14815);
or U15164 (N_15164,N_14878,N_14991);
or U15165 (N_15165,N_14815,N_14943);
or U15166 (N_15166,N_14823,N_14926);
and U15167 (N_15167,N_14946,N_14860);
nor U15168 (N_15168,N_14826,N_14888);
or U15169 (N_15169,N_14816,N_14843);
nor U15170 (N_15170,N_14976,N_14940);
nor U15171 (N_15171,N_14869,N_14891);
and U15172 (N_15172,N_14875,N_14851);
xor U15173 (N_15173,N_14992,N_14903);
nor U15174 (N_15174,N_14838,N_14909);
nand U15175 (N_15175,N_14977,N_14820);
xnor U15176 (N_15176,N_14935,N_14944);
or U15177 (N_15177,N_14872,N_14925);
nand U15178 (N_15178,N_14977,N_14807);
xor U15179 (N_15179,N_14873,N_14859);
or U15180 (N_15180,N_14826,N_14937);
or U15181 (N_15181,N_14834,N_14971);
and U15182 (N_15182,N_14856,N_14893);
and U15183 (N_15183,N_14941,N_14908);
and U15184 (N_15184,N_14860,N_14808);
nand U15185 (N_15185,N_14822,N_14895);
xnor U15186 (N_15186,N_14816,N_14929);
xnor U15187 (N_15187,N_14933,N_14965);
or U15188 (N_15188,N_14830,N_14802);
xor U15189 (N_15189,N_14886,N_14889);
xor U15190 (N_15190,N_14846,N_14839);
and U15191 (N_15191,N_14952,N_14824);
nor U15192 (N_15192,N_14800,N_14820);
nand U15193 (N_15193,N_14970,N_14881);
or U15194 (N_15194,N_14869,N_14857);
and U15195 (N_15195,N_14860,N_14870);
and U15196 (N_15196,N_14993,N_14905);
nand U15197 (N_15197,N_14966,N_14982);
or U15198 (N_15198,N_14903,N_14913);
or U15199 (N_15199,N_14985,N_14979);
nand U15200 (N_15200,N_15189,N_15100);
and U15201 (N_15201,N_15000,N_15198);
nor U15202 (N_15202,N_15167,N_15011);
nor U15203 (N_15203,N_15036,N_15015);
or U15204 (N_15204,N_15009,N_15027);
nor U15205 (N_15205,N_15058,N_15172);
xor U15206 (N_15206,N_15098,N_15071);
nand U15207 (N_15207,N_15076,N_15032);
nand U15208 (N_15208,N_15166,N_15038);
or U15209 (N_15209,N_15079,N_15113);
xnor U15210 (N_15210,N_15059,N_15074);
nor U15211 (N_15211,N_15126,N_15083);
or U15212 (N_15212,N_15073,N_15193);
nor U15213 (N_15213,N_15134,N_15022);
or U15214 (N_15214,N_15163,N_15066);
xor U15215 (N_15215,N_15170,N_15116);
xor U15216 (N_15216,N_15191,N_15169);
and U15217 (N_15217,N_15041,N_15147);
nand U15218 (N_15218,N_15174,N_15008);
or U15219 (N_15219,N_15110,N_15108);
or U15220 (N_15220,N_15107,N_15149);
xor U15221 (N_15221,N_15117,N_15195);
nor U15222 (N_15222,N_15093,N_15124);
nand U15223 (N_15223,N_15096,N_15137);
nand U15224 (N_15224,N_15104,N_15077);
nor U15225 (N_15225,N_15070,N_15190);
and U15226 (N_15226,N_15075,N_15141);
xor U15227 (N_15227,N_15173,N_15086);
or U15228 (N_15228,N_15092,N_15161);
xnor U15229 (N_15229,N_15154,N_15055);
or U15230 (N_15230,N_15181,N_15177);
or U15231 (N_15231,N_15188,N_15040);
xnor U15232 (N_15232,N_15001,N_15025);
or U15233 (N_15233,N_15136,N_15153);
xor U15234 (N_15234,N_15048,N_15056);
nor U15235 (N_15235,N_15034,N_15033);
xnor U15236 (N_15236,N_15168,N_15016);
xnor U15237 (N_15237,N_15120,N_15186);
nor U15238 (N_15238,N_15155,N_15006);
and U15239 (N_15239,N_15044,N_15157);
and U15240 (N_15240,N_15180,N_15084);
and U15241 (N_15241,N_15158,N_15050);
and U15242 (N_15242,N_15176,N_15131);
and U15243 (N_15243,N_15132,N_15165);
nand U15244 (N_15244,N_15045,N_15114);
or U15245 (N_15245,N_15065,N_15199);
nand U15246 (N_15246,N_15028,N_15089);
nand U15247 (N_15247,N_15078,N_15042);
nor U15248 (N_15248,N_15024,N_15021);
xor U15249 (N_15249,N_15194,N_15017);
or U15250 (N_15250,N_15182,N_15128);
or U15251 (N_15251,N_15064,N_15004);
and U15252 (N_15252,N_15002,N_15106);
and U15253 (N_15253,N_15103,N_15109);
or U15254 (N_15254,N_15111,N_15019);
or U15255 (N_15255,N_15068,N_15095);
xor U15256 (N_15256,N_15018,N_15192);
xnor U15257 (N_15257,N_15178,N_15007);
xnor U15258 (N_15258,N_15184,N_15102);
xnor U15259 (N_15259,N_15010,N_15197);
or U15260 (N_15260,N_15049,N_15123);
nand U15261 (N_15261,N_15130,N_15088);
or U15262 (N_15262,N_15080,N_15031);
and U15263 (N_15263,N_15175,N_15003);
nand U15264 (N_15264,N_15133,N_15105);
or U15265 (N_15265,N_15087,N_15118);
nor U15266 (N_15266,N_15138,N_15051);
and U15267 (N_15267,N_15023,N_15090);
nand U15268 (N_15268,N_15035,N_15037);
nor U15269 (N_15269,N_15187,N_15145);
or U15270 (N_15270,N_15030,N_15020);
or U15271 (N_15271,N_15144,N_15125);
xnor U15272 (N_15272,N_15060,N_15013);
nand U15273 (N_15273,N_15014,N_15143);
nor U15274 (N_15274,N_15069,N_15135);
or U15275 (N_15275,N_15121,N_15085);
nor U15276 (N_15276,N_15129,N_15062);
and U15277 (N_15277,N_15179,N_15052);
or U15278 (N_15278,N_15139,N_15043);
xnor U15279 (N_15279,N_15127,N_15082);
or U15280 (N_15280,N_15122,N_15164);
nand U15281 (N_15281,N_15142,N_15150);
or U15282 (N_15282,N_15053,N_15146);
nor U15283 (N_15283,N_15171,N_15054);
nor U15284 (N_15284,N_15047,N_15094);
nor U15285 (N_15285,N_15183,N_15026);
nor U15286 (N_15286,N_15159,N_15160);
or U15287 (N_15287,N_15151,N_15152);
or U15288 (N_15288,N_15115,N_15012);
or U15289 (N_15289,N_15185,N_15119);
xor U15290 (N_15290,N_15067,N_15005);
xor U15291 (N_15291,N_15101,N_15063);
or U15292 (N_15292,N_15196,N_15091);
nor U15293 (N_15293,N_15148,N_15029);
xor U15294 (N_15294,N_15081,N_15039);
and U15295 (N_15295,N_15140,N_15046);
nand U15296 (N_15296,N_15097,N_15072);
and U15297 (N_15297,N_15057,N_15099);
xnor U15298 (N_15298,N_15162,N_15156);
nor U15299 (N_15299,N_15061,N_15112);
nor U15300 (N_15300,N_15089,N_15074);
or U15301 (N_15301,N_15098,N_15073);
nor U15302 (N_15302,N_15010,N_15102);
nor U15303 (N_15303,N_15149,N_15038);
nor U15304 (N_15304,N_15124,N_15106);
or U15305 (N_15305,N_15018,N_15011);
or U15306 (N_15306,N_15008,N_15036);
nand U15307 (N_15307,N_15026,N_15147);
nand U15308 (N_15308,N_15101,N_15138);
xnor U15309 (N_15309,N_15092,N_15063);
or U15310 (N_15310,N_15163,N_15087);
nor U15311 (N_15311,N_15030,N_15198);
or U15312 (N_15312,N_15167,N_15012);
xnor U15313 (N_15313,N_15169,N_15062);
nand U15314 (N_15314,N_15187,N_15045);
xor U15315 (N_15315,N_15037,N_15144);
nand U15316 (N_15316,N_15040,N_15121);
nand U15317 (N_15317,N_15068,N_15128);
nand U15318 (N_15318,N_15048,N_15097);
nand U15319 (N_15319,N_15118,N_15113);
nor U15320 (N_15320,N_15165,N_15191);
nand U15321 (N_15321,N_15159,N_15190);
and U15322 (N_15322,N_15094,N_15020);
nand U15323 (N_15323,N_15079,N_15029);
or U15324 (N_15324,N_15199,N_15142);
nor U15325 (N_15325,N_15128,N_15078);
and U15326 (N_15326,N_15118,N_15085);
nand U15327 (N_15327,N_15105,N_15026);
or U15328 (N_15328,N_15032,N_15051);
nor U15329 (N_15329,N_15028,N_15147);
nand U15330 (N_15330,N_15012,N_15062);
and U15331 (N_15331,N_15066,N_15072);
or U15332 (N_15332,N_15114,N_15074);
nand U15333 (N_15333,N_15021,N_15016);
nor U15334 (N_15334,N_15108,N_15050);
and U15335 (N_15335,N_15169,N_15141);
nand U15336 (N_15336,N_15029,N_15114);
nor U15337 (N_15337,N_15074,N_15118);
xnor U15338 (N_15338,N_15087,N_15116);
or U15339 (N_15339,N_15022,N_15025);
and U15340 (N_15340,N_15166,N_15150);
nor U15341 (N_15341,N_15005,N_15079);
nor U15342 (N_15342,N_15088,N_15127);
or U15343 (N_15343,N_15177,N_15064);
nor U15344 (N_15344,N_15034,N_15092);
nand U15345 (N_15345,N_15010,N_15069);
xnor U15346 (N_15346,N_15101,N_15162);
xnor U15347 (N_15347,N_15116,N_15171);
or U15348 (N_15348,N_15078,N_15043);
nor U15349 (N_15349,N_15010,N_15095);
nor U15350 (N_15350,N_15101,N_15038);
nand U15351 (N_15351,N_15104,N_15006);
or U15352 (N_15352,N_15097,N_15078);
or U15353 (N_15353,N_15159,N_15055);
xor U15354 (N_15354,N_15000,N_15005);
and U15355 (N_15355,N_15196,N_15168);
xnor U15356 (N_15356,N_15095,N_15088);
or U15357 (N_15357,N_15161,N_15014);
and U15358 (N_15358,N_15087,N_15059);
nand U15359 (N_15359,N_15035,N_15025);
nand U15360 (N_15360,N_15189,N_15137);
nor U15361 (N_15361,N_15020,N_15066);
nor U15362 (N_15362,N_15114,N_15109);
nor U15363 (N_15363,N_15125,N_15024);
xor U15364 (N_15364,N_15147,N_15197);
nand U15365 (N_15365,N_15050,N_15113);
and U15366 (N_15366,N_15100,N_15109);
and U15367 (N_15367,N_15128,N_15053);
nand U15368 (N_15368,N_15073,N_15028);
xnor U15369 (N_15369,N_15029,N_15095);
xor U15370 (N_15370,N_15152,N_15091);
or U15371 (N_15371,N_15080,N_15094);
and U15372 (N_15372,N_15199,N_15113);
and U15373 (N_15373,N_15027,N_15196);
xnor U15374 (N_15374,N_15193,N_15106);
nand U15375 (N_15375,N_15039,N_15022);
nor U15376 (N_15376,N_15073,N_15048);
or U15377 (N_15377,N_15030,N_15048);
nor U15378 (N_15378,N_15110,N_15097);
xor U15379 (N_15379,N_15050,N_15103);
and U15380 (N_15380,N_15109,N_15142);
xor U15381 (N_15381,N_15183,N_15172);
xnor U15382 (N_15382,N_15070,N_15063);
xor U15383 (N_15383,N_15169,N_15006);
xor U15384 (N_15384,N_15020,N_15077);
or U15385 (N_15385,N_15126,N_15116);
nand U15386 (N_15386,N_15036,N_15026);
or U15387 (N_15387,N_15036,N_15171);
xor U15388 (N_15388,N_15049,N_15091);
nor U15389 (N_15389,N_15016,N_15127);
nor U15390 (N_15390,N_15061,N_15133);
xor U15391 (N_15391,N_15135,N_15192);
nand U15392 (N_15392,N_15067,N_15173);
xor U15393 (N_15393,N_15178,N_15124);
or U15394 (N_15394,N_15182,N_15014);
and U15395 (N_15395,N_15181,N_15178);
nor U15396 (N_15396,N_15030,N_15111);
xnor U15397 (N_15397,N_15149,N_15011);
or U15398 (N_15398,N_15109,N_15186);
and U15399 (N_15399,N_15088,N_15155);
nand U15400 (N_15400,N_15346,N_15317);
or U15401 (N_15401,N_15328,N_15367);
and U15402 (N_15402,N_15208,N_15362);
or U15403 (N_15403,N_15300,N_15283);
nand U15404 (N_15404,N_15270,N_15333);
or U15405 (N_15405,N_15298,N_15206);
nand U15406 (N_15406,N_15343,N_15309);
and U15407 (N_15407,N_15369,N_15393);
nand U15408 (N_15408,N_15353,N_15341);
xnor U15409 (N_15409,N_15245,N_15234);
nor U15410 (N_15410,N_15320,N_15335);
nand U15411 (N_15411,N_15292,N_15390);
or U15412 (N_15412,N_15248,N_15288);
nor U15413 (N_15413,N_15297,N_15258);
or U15414 (N_15414,N_15267,N_15228);
or U15415 (N_15415,N_15312,N_15289);
nand U15416 (N_15416,N_15392,N_15397);
or U15417 (N_15417,N_15259,N_15386);
xnor U15418 (N_15418,N_15381,N_15327);
nand U15419 (N_15419,N_15365,N_15332);
nand U15420 (N_15420,N_15374,N_15242);
nor U15421 (N_15421,N_15360,N_15231);
nand U15422 (N_15422,N_15273,N_15344);
or U15423 (N_15423,N_15255,N_15268);
or U15424 (N_15424,N_15329,N_15314);
nand U15425 (N_15425,N_15239,N_15337);
xor U15426 (N_15426,N_15313,N_15265);
and U15427 (N_15427,N_15303,N_15290);
and U15428 (N_15428,N_15287,N_15241);
and U15429 (N_15429,N_15200,N_15230);
nand U15430 (N_15430,N_15395,N_15366);
nor U15431 (N_15431,N_15282,N_15201);
nand U15432 (N_15432,N_15348,N_15210);
nor U15433 (N_15433,N_15378,N_15250);
or U15434 (N_15434,N_15304,N_15319);
xor U15435 (N_15435,N_15339,N_15363);
xor U15436 (N_15436,N_15269,N_15247);
nor U15437 (N_15437,N_15243,N_15235);
or U15438 (N_15438,N_15316,N_15254);
nor U15439 (N_15439,N_15264,N_15331);
or U15440 (N_15440,N_15311,N_15203);
nor U15441 (N_15441,N_15222,N_15285);
xor U15442 (N_15442,N_15275,N_15351);
nand U15443 (N_15443,N_15356,N_15215);
xor U15444 (N_15444,N_15226,N_15322);
xnor U15445 (N_15445,N_15295,N_15213);
and U15446 (N_15446,N_15349,N_15217);
xnor U15447 (N_15447,N_15240,N_15315);
nor U15448 (N_15448,N_15384,N_15318);
and U15449 (N_15449,N_15387,N_15350);
nand U15450 (N_15450,N_15352,N_15361);
nand U15451 (N_15451,N_15294,N_15375);
nand U15452 (N_15452,N_15212,N_15355);
xor U15453 (N_15453,N_15370,N_15225);
nor U15454 (N_15454,N_15336,N_15347);
or U15455 (N_15455,N_15205,N_15244);
nand U15456 (N_15456,N_15389,N_15207);
or U15457 (N_15457,N_15261,N_15237);
nand U15458 (N_15458,N_15305,N_15321);
and U15459 (N_15459,N_15330,N_15204);
nor U15460 (N_15460,N_15278,N_15396);
xor U15461 (N_15461,N_15280,N_15246);
nand U15462 (N_15462,N_15345,N_15307);
or U15463 (N_15463,N_15286,N_15296);
xnor U15464 (N_15464,N_15236,N_15372);
xor U15465 (N_15465,N_15232,N_15227);
and U15466 (N_15466,N_15249,N_15377);
and U15467 (N_15467,N_15379,N_15284);
nand U15468 (N_15468,N_15233,N_15383);
and U15469 (N_15469,N_15334,N_15260);
nand U15470 (N_15470,N_15299,N_15263);
or U15471 (N_15471,N_15388,N_15373);
nand U15472 (N_15472,N_15272,N_15358);
nand U15473 (N_15473,N_15324,N_15216);
nor U15474 (N_15474,N_15224,N_15223);
nand U15475 (N_15475,N_15323,N_15238);
xnor U15476 (N_15476,N_15209,N_15340);
nand U15477 (N_15477,N_15262,N_15376);
or U15478 (N_15478,N_15291,N_15325);
and U15479 (N_15479,N_15221,N_15253);
and U15480 (N_15480,N_15256,N_15281);
nand U15481 (N_15481,N_15211,N_15391);
nor U15482 (N_15482,N_15357,N_15398);
nor U15483 (N_15483,N_15382,N_15354);
or U15484 (N_15484,N_15306,N_15338);
nor U15485 (N_15485,N_15380,N_15214);
xnor U15486 (N_15486,N_15302,N_15271);
xor U15487 (N_15487,N_15252,N_15385);
xor U15488 (N_15488,N_15251,N_15277);
and U15489 (N_15489,N_15326,N_15257);
xor U15490 (N_15490,N_15359,N_15293);
and U15491 (N_15491,N_15394,N_15229);
nand U15492 (N_15492,N_15218,N_15301);
nor U15493 (N_15493,N_15220,N_15364);
xnor U15494 (N_15494,N_15399,N_15371);
or U15495 (N_15495,N_15276,N_15310);
xor U15496 (N_15496,N_15274,N_15279);
or U15497 (N_15497,N_15202,N_15368);
nor U15498 (N_15498,N_15342,N_15308);
nand U15499 (N_15499,N_15219,N_15266);
nor U15500 (N_15500,N_15243,N_15297);
nor U15501 (N_15501,N_15218,N_15366);
xor U15502 (N_15502,N_15240,N_15319);
xnor U15503 (N_15503,N_15287,N_15377);
nor U15504 (N_15504,N_15302,N_15317);
or U15505 (N_15505,N_15353,N_15278);
or U15506 (N_15506,N_15334,N_15204);
xnor U15507 (N_15507,N_15313,N_15222);
nor U15508 (N_15508,N_15267,N_15301);
or U15509 (N_15509,N_15311,N_15264);
xor U15510 (N_15510,N_15240,N_15212);
or U15511 (N_15511,N_15395,N_15212);
or U15512 (N_15512,N_15323,N_15342);
nor U15513 (N_15513,N_15296,N_15298);
and U15514 (N_15514,N_15289,N_15314);
nor U15515 (N_15515,N_15272,N_15293);
nand U15516 (N_15516,N_15230,N_15228);
and U15517 (N_15517,N_15263,N_15215);
xor U15518 (N_15518,N_15396,N_15237);
or U15519 (N_15519,N_15378,N_15240);
xnor U15520 (N_15520,N_15355,N_15223);
or U15521 (N_15521,N_15237,N_15293);
xnor U15522 (N_15522,N_15254,N_15358);
or U15523 (N_15523,N_15395,N_15254);
nor U15524 (N_15524,N_15288,N_15292);
nand U15525 (N_15525,N_15204,N_15305);
nor U15526 (N_15526,N_15325,N_15296);
xnor U15527 (N_15527,N_15365,N_15253);
or U15528 (N_15528,N_15337,N_15260);
nor U15529 (N_15529,N_15288,N_15362);
nand U15530 (N_15530,N_15209,N_15339);
nand U15531 (N_15531,N_15397,N_15219);
nand U15532 (N_15532,N_15322,N_15201);
nor U15533 (N_15533,N_15335,N_15243);
xnor U15534 (N_15534,N_15376,N_15390);
nor U15535 (N_15535,N_15360,N_15365);
or U15536 (N_15536,N_15292,N_15257);
and U15537 (N_15537,N_15389,N_15321);
or U15538 (N_15538,N_15321,N_15336);
nand U15539 (N_15539,N_15343,N_15382);
xnor U15540 (N_15540,N_15388,N_15220);
xor U15541 (N_15541,N_15343,N_15236);
nor U15542 (N_15542,N_15231,N_15343);
xnor U15543 (N_15543,N_15224,N_15236);
and U15544 (N_15544,N_15366,N_15276);
or U15545 (N_15545,N_15391,N_15360);
or U15546 (N_15546,N_15308,N_15201);
and U15547 (N_15547,N_15385,N_15351);
xnor U15548 (N_15548,N_15237,N_15314);
nor U15549 (N_15549,N_15326,N_15359);
nand U15550 (N_15550,N_15271,N_15367);
and U15551 (N_15551,N_15236,N_15256);
xor U15552 (N_15552,N_15234,N_15267);
nand U15553 (N_15553,N_15364,N_15382);
nor U15554 (N_15554,N_15309,N_15326);
nand U15555 (N_15555,N_15280,N_15356);
or U15556 (N_15556,N_15370,N_15351);
or U15557 (N_15557,N_15355,N_15201);
nor U15558 (N_15558,N_15232,N_15398);
nor U15559 (N_15559,N_15201,N_15276);
nand U15560 (N_15560,N_15321,N_15362);
and U15561 (N_15561,N_15330,N_15253);
or U15562 (N_15562,N_15280,N_15386);
xor U15563 (N_15563,N_15346,N_15390);
nor U15564 (N_15564,N_15358,N_15263);
xnor U15565 (N_15565,N_15348,N_15247);
or U15566 (N_15566,N_15266,N_15272);
or U15567 (N_15567,N_15205,N_15256);
xnor U15568 (N_15568,N_15350,N_15397);
and U15569 (N_15569,N_15291,N_15314);
nor U15570 (N_15570,N_15223,N_15204);
and U15571 (N_15571,N_15308,N_15286);
xor U15572 (N_15572,N_15214,N_15282);
or U15573 (N_15573,N_15318,N_15362);
or U15574 (N_15574,N_15246,N_15398);
and U15575 (N_15575,N_15325,N_15249);
nor U15576 (N_15576,N_15249,N_15330);
nor U15577 (N_15577,N_15331,N_15257);
and U15578 (N_15578,N_15350,N_15341);
and U15579 (N_15579,N_15214,N_15264);
nor U15580 (N_15580,N_15277,N_15285);
nor U15581 (N_15581,N_15223,N_15329);
nand U15582 (N_15582,N_15321,N_15391);
or U15583 (N_15583,N_15291,N_15227);
xor U15584 (N_15584,N_15374,N_15250);
and U15585 (N_15585,N_15257,N_15362);
xnor U15586 (N_15586,N_15302,N_15237);
or U15587 (N_15587,N_15311,N_15289);
and U15588 (N_15588,N_15335,N_15284);
or U15589 (N_15589,N_15315,N_15357);
nor U15590 (N_15590,N_15223,N_15288);
nand U15591 (N_15591,N_15288,N_15221);
xor U15592 (N_15592,N_15313,N_15203);
or U15593 (N_15593,N_15220,N_15345);
or U15594 (N_15594,N_15204,N_15358);
and U15595 (N_15595,N_15234,N_15336);
nand U15596 (N_15596,N_15312,N_15317);
nand U15597 (N_15597,N_15373,N_15285);
xnor U15598 (N_15598,N_15257,N_15325);
nand U15599 (N_15599,N_15235,N_15390);
nor U15600 (N_15600,N_15423,N_15543);
nand U15601 (N_15601,N_15501,N_15442);
or U15602 (N_15602,N_15558,N_15524);
or U15603 (N_15603,N_15517,N_15460);
and U15604 (N_15604,N_15400,N_15450);
xor U15605 (N_15605,N_15463,N_15504);
nand U15606 (N_15606,N_15557,N_15457);
and U15607 (N_15607,N_15537,N_15401);
and U15608 (N_15608,N_15597,N_15403);
nand U15609 (N_15609,N_15506,N_15451);
or U15610 (N_15610,N_15592,N_15563);
xnor U15611 (N_15611,N_15479,N_15418);
nor U15612 (N_15612,N_15512,N_15413);
nand U15613 (N_15613,N_15476,N_15435);
nand U15614 (N_15614,N_15415,N_15478);
nor U15615 (N_15615,N_15470,N_15477);
nor U15616 (N_15616,N_15409,N_15410);
nor U15617 (N_15617,N_15514,N_15575);
nor U15618 (N_15618,N_15532,N_15586);
and U15619 (N_15619,N_15591,N_15579);
and U15620 (N_15620,N_15493,N_15578);
nor U15621 (N_15621,N_15588,N_15509);
nand U15622 (N_15622,N_15553,N_15444);
nor U15623 (N_15623,N_15468,N_15582);
or U15624 (N_15624,N_15564,N_15437);
nor U15625 (N_15625,N_15590,N_15533);
nor U15626 (N_15626,N_15500,N_15552);
and U15627 (N_15627,N_15443,N_15492);
or U15628 (N_15628,N_15521,N_15416);
xor U15629 (N_15629,N_15561,N_15518);
nor U15630 (N_15630,N_15507,N_15599);
and U15631 (N_15631,N_15421,N_15522);
nand U15632 (N_15632,N_15471,N_15449);
nor U15633 (N_15633,N_15595,N_15598);
or U15634 (N_15634,N_15488,N_15498);
nand U15635 (N_15635,N_15546,N_15448);
or U15636 (N_15636,N_15411,N_15464);
and U15637 (N_15637,N_15528,N_15534);
nand U15638 (N_15638,N_15475,N_15473);
nand U15639 (N_15639,N_15513,N_15540);
and U15640 (N_15640,N_15531,N_15490);
nand U15641 (N_15641,N_15458,N_15407);
nor U15642 (N_15642,N_15527,N_15529);
or U15643 (N_15643,N_15583,N_15412);
xnor U15644 (N_15644,N_15550,N_15565);
xnor U15645 (N_15645,N_15420,N_15538);
and U15646 (N_15646,N_15589,N_15480);
or U15647 (N_15647,N_15545,N_15580);
or U15648 (N_15648,N_15526,N_15472);
or U15649 (N_15649,N_15431,N_15520);
or U15650 (N_15650,N_15519,N_15581);
xor U15651 (N_15651,N_15574,N_15573);
and U15652 (N_15652,N_15454,N_15441);
nand U15653 (N_15653,N_15515,N_15426);
or U15654 (N_15654,N_15474,N_15505);
and U15655 (N_15655,N_15456,N_15497);
nor U15656 (N_15656,N_15429,N_15495);
nand U15657 (N_15657,N_15424,N_15419);
xor U15658 (N_15658,N_15459,N_15568);
xor U15659 (N_15659,N_15484,N_15503);
xnor U15660 (N_15660,N_15494,N_15428);
or U15661 (N_15661,N_15406,N_15562);
nand U15662 (N_15662,N_15511,N_15486);
and U15663 (N_15663,N_15402,N_15465);
and U15664 (N_15664,N_15542,N_15438);
or U15665 (N_15665,N_15499,N_15425);
and U15666 (N_15666,N_15487,N_15452);
nand U15667 (N_15667,N_15571,N_15439);
or U15668 (N_15668,N_15466,N_15485);
or U15669 (N_15669,N_15567,N_15434);
or U15670 (N_15670,N_15516,N_15445);
or U15671 (N_15671,N_15530,N_15523);
or U15672 (N_15672,N_15572,N_15404);
nand U15673 (N_15673,N_15483,N_15548);
xor U15674 (N_15674,N_15559,N_15585);
xor U15675 (N_15675,N_15570,N_15440);
nor U15676 (N_15676,N_15481,N_15560);
xnor U15677 (N_15677,N_15569,N_15455);
nand U15678 (N_15678,N_15414,N_15405);
xor U15679 (N_15679,N_15549,N_15482);
or U15680 (N_15680,N_15436,N_15510);
and U15681 (N_15681,N_15417,N_15467);
and U15682 (N_15682,N_15469,N_15489);
or U15683 (N_15683,N_15408,N_15547);
nand U15684 (N_15684,N_15566,N_15496);
or U15685 (N_15685,N_15554,N_15462);
nand U15686 (N_15686,N_15432,N_15535);
or U15687 (N_15687,N_15461,N_15584);
xnor U15688 (N_15688,N_15525,N_15422);
nor U15689 (N_15689,N_15502,N_15491);
or U15690 (N_15690,N_15596,N_15577);
nand U15691 (N_15691,N_15593,N_15427);
nor U15692 (N_15692,N_15576,N_15541);
xnor U15693 (N_15693,N_15433,N_15447);
xnor U15694 (N_15694,N_15551,N_15430);
or U15695 (N_15695,N_15594,N_15555);
and U15696 (N_15696,N_15556,N_15587);
and U15697 (N_15697,N_15544,N_15508);
nor U15698 (N_15698,N_15539,N_15453);
nor U15699 (N_15699,N_15446,N_15536);
xor U15700 (N_15700,N_15546,N_15594);
or U15701 (N_15701,N_15546,N_15436);
xnor U15702 (N_15702,N_15424,N_15571);
and U15703 (N_15703,N_15534,N_15502);
xnor U15704 (N_15704,N_15576,N_15538);
or U15705 (N_15705,N_15501,N_15580);
nor U15706 (N_15706,N_15447,N_15529);
xnor U15707 (N_15707,N_15521,N_15482);
or U15708 (N_15708,N_15406,N_15463);
xor U15709 (N_15709,N_15498,N_15435);
xor U15710 (N_15710,N_15548,N_15405);
nor U15711 (N_15711,N_15484,N_15409);
nand U15712 (N_15712,N_15536,N_15424);
nor U15713 (N_15713,N_15507,N_15497);
nand U15714 (N_15714,N_15541,N_15529);
and U15715 (N_15715,N_15466,N_15429);
xor U15716 (N_15716,N_15563,N_15593);
or U15717 (N_15717,N_15525,N_15488);
or U15718 (N_15718,N_15409,N_15426);
and U15719 (N_15719,N_15416,N_15583);
nor U15720 (N_15720,N_15569,N_15599);
and U15721 (N_15721,N_15568,N_15592);
nor U15722 (N_15722,N_15453,N_15526);
nor U15723 (N_15723,N_15579,N_15477);
nor U15724 (N_15724,N_15413,N_15522);
xor U15725 (N_15725,N_15469,N_15451);
nor U15726 (N_15726,N_15443,N_15575);
and U15727 (N_15727,N_15469,N_15417);
and U15728 (N_15728,N_15457,N_15579);
or U15729 (N_15729,N_15438,N_15581);
xor U15730 (N_15730,N_15421,N_15513);
nor U15731 (N_15731,N_15573,N_15435);
nor U15732 (N_15732,N_15471,N_15419);
nand U15733 (N_15733,N_15569,N_15495);
nor U15734 (N_15734,N_15515,N_15473);
nor U15735 (N_15735,N_15448,N_15566);
nor U15736 (N_15736,N_15506,N_15512);
xnor U15737 (N_15737,N_15419,N_15510);
nor U15738 (N_15738,N_15547,N_15562);
nor U15739 (N_15739,N_15426,N_15536);
or U15740 (N_15740,N_15585,N_15545);
xor U15741 (N_15741,N_15480,N_15439);
nand U15742 (N_15742,N_15450,N_15448);
nor U15743 (N_15743,N_15401,N_15407);
nand U15744 (N_15744,N_15513,N_15554);
and U15745 (N_15745,N_15421,N_15539);
xor U15746 (N_15746,N_15481,N_15544);
xor U15747 (N_15747,N_15496,N_15405);
nand U15748 (N_15748,N_15520,N_15521);
xor U15749 (N_15749,N_15525,N_15444);
nor U15750 (N_15750,N_15402,N_15448);
nand U15751 (N_15751,N_15583,N_15550);
nor U15752 (N_15752,N_15457,N_15414);
xor U15753 (N_15753,N_15594,N_15415);
or U15754 (N_15754,N_15414,N_15466);
nor U15755 (N_15755,N_15505,N_15432);
xor U15756 (N_15756,N_15498,N_15463);
or U15757 (N_15757,N_15447,N_15579);
or U15758 (N_15758,N_15554,N_15524);
and U15759 (N_15759,N_15454,N_15512);
or U15760 (N_15760,N_15546,N_15508);
or U15761 (N_15761,N_15596,N_15410);
and U15762 (N_15762,N_15561,N_15443);
xnor U15763 (N_15763,N_15414,N_15550);
nand U15764 (N_15764,N_15551,N_15581);
and U15765 (N_15765,N_15472,N_15566);
or U15766 (N_15766,N_15437,N_15461);
or U15767 (N_15767,N_15536,N_15407);
nor U15768 (N_15768,N_15479,N_15441);
xnor U15769 (N_15769,N_15488,N_15534);
and U15770 (N_15770,N_15527,N_15452);
nor U15771 (N_15771,N_15496,N_15501);
and U15772 (N_15772,N_15563,N_15570);
xnor U15773 (N_15773,N_15415,N_15464);
nor U15774 (N_15774,N_15520,N_15482);
nand U15775 (N_15775,N_15548,N_15474);
nor U15776 (N_15776,N_15479,N_15456);
and U15777 (N_15777,N_15536,N_15565);
nor U15778 (N_15778,N_15493,N_15472);
or U15779 (N_15779,N_15485,N_15460);
xor U15780 (N_15780,N_15521,N_15451);
xor U15781 (N_15781,N_15478,N_15521);
xnor U15782 (N_15782,N_15505,N_15441);
nor U15783 (N_15783,N_15518,N_15541);
xnor U15784 (N_15784,N_15455,N_15461);
nor U15785 (N_15785,N_15599,N_15476);
or U15786 (N_15786,N_15535,N_15571);
or U15787 (N_15787,N_15455,N_15587);
nand U15788 (N_15788,N_15567,N_15507);
nor U15789 (N_15789,N_15435,N_15494);
and U15790 (N_15790,N_15404,N_15570);
nor U15791 (N_15791,N_15431,N_15482);
or U15792 (N_15792,N_15577,N_15487);
nand U15793 (N_15793,N_15492,N_15586);
nand U15794 (N_15794,N_15494,N_15426);
and U15795 (N_15795,N_15535,N_15490);
and U15796 (N_15796,N_15565,N_15492);
or U15797 (N_15797,N_15497,N_15501);
nor U15798 (N_15798,N_15558,N_15475);
and U15799 (N_15799,N_15599,N_15528);
and U15800 (N_15800,N_15646,N_15711);
xor U15801 (N_15801,N_15753,N_15781);
nor U15802 (N_15802,N_15627,N_15709);
nand U15803 (N_15803,N_15616,N_15706);
and U15804 (N_15804,N_15644,N_15683);
nor U15805 (N_15805,N_15707,N_15654);
or U15806 (N_15806,N_15685,N_15780);
and U15807 (N_15807,N_15613,N_15757);
xnor U15808 (N_15808,N_15676,N_15673);
and U15809 (N_15809,N_15652,N_15731);
xor U15810 (N_15810,N_15720,N_15784);
or U15811 (N_15811,N_15642,N_15611);
xnor U15812 (N_15812,N_15689,N_15747);
or U15813 (N_15813,N_15733,N_15695);
or U15814 (N_15814,N_15632,N_15741);
xnor U15815 (N_15815,N_15788,N_15633);
or U15816 (N_15816,N_15620,N_15699);
nand U15817 (N_15817,N_15610,N_15766);
and U15818 (N_15818,N_15630,N_15797);
xor U15819 (N_15819,N_15617,N_15723);
or U15820 (N_15820,N_15771,N_15726);
nand U15821 (N_15821,N_15730,N_15792);
or U15822 (N_15822,N_15744,N_15649);
nand U15823 (N_15823,N_15715,N_15607);
or U15824 (N_15824,N_15614,N_15727);
and U15825 (N_15825,N_15653,N_15767);
and U15826 (N_15826,N_15629,N_15623);
xnor U15827 (N_15827,N_15664,N_15713);
and U15828 (N_15828,N_15751,N_15705);
nand U15829 (N_15829,N_15745,N_15693);
xnor U15830 (N_15830,N_15671,N_15722);
and U15831 (N_15831,N_15658,N_15645);
or U15832 (N_15832,N_15626,N_15735);
and U15833 (N_15833,N_15721,N_15691);
nor U15834 (N_15834,N_15750,N_15606);
nor U15835 (N_15835,N_15764,N_15748);
nand U15836 (N_15836,N_15643,N_15602);
nor U15837 (N_15837,N_15789,N_15637);
nor U15838 (N_15838,N_15687,N_15754);
nor U15839 (N_15839,N_15628,N_15675);
xor U15840 (N_15840,N_15700,N_15663);
or U15841 (N_15841,N_15682,N_15694);
nand U15842 (N_15842,N_15716,N_15679);
xnor U15843 (N_15843,N_15796,N_15625);
or U15844 (N_15844,N_15605,N_15634);
nor U15845 (N_15845,N_15657,N_15742);
and U15846 (N_15846,N_15774,N_15697);
nor U15847 (N_15847,N_15794,N_15677);
xor U15848 (N_15848,N_15698,N_15631);
or U15849 (N_15849,N_15684,N_15791);
or U15850 (N_15850,N_15725,N_15670);
or U15851 (N_15851,N_15786,N_15604);
nor U15852 (N_15852,N_15704,N_15612);
or U15853 (N_15853,N_15712,N_15656);
nand U15854 (N_15854,N_15667,N_15690);
nand U15855 (N_15855,N_15749,N_15708);
and U15856 (N_15856,N_15703,N_15669);
xor U15857 (N_15857,N_15680,N_15779);
and U15858 (N_15858,N_15717,N_15729);
or U15859 (N_15859,N_15692,N_15778);
nand U15860 (N_15860,N_15762,N_15795);
and U15861 (N_15861,N_15732,N_15724);
xnor U15862 (N_15862,N_15760,N_15743);
or U15863 (N_15863,N_15702,N_15769);
xor U15864 (N_15864,N_15672,N_15798);
and U15865 (N_15865,N_15661,N_15674);
nor U15866 (N_15866,N_15718,N_15752);
and U15867 (N_15867,N_15624,N_15609);
nand U15868 (N_15868,N_15768,N_15782);
nor U15869 (N_15869,N_15608,N_15701);
nand U15870 (N_15870,N_15619,N_15790);
nand U15871 (N_15871,N_15600,N_15777);
or U15872 (N_15872,N_15772,N_15775);
or U15873 (N_15873,N_15603,N_15696);
nand U15874 (N_15874,N_15662,N_15668);
or U15875 (N_15875,N_15755,N_15665);
nand U15876 (N_15876,N_15770,N_15785);
nand U15877 (N_15877,N_15601,N_15734);
or U15878 (N_15878,N_15678,N_15759);
or U15879 (N_15879,N_15641,N_15666);
nand U15880 (N_15880,N_15756,N_15776);
or U15881 (N_15881,N_15761,N_15615);
and U15882 (N_15882,N_15746,N_15622);
nand U15883 (N_15883,N_15648,N_15736);
xor U15884 (N_15884,N_15728,N_15650);
xor U15885 (N_15885,N_15660,N_15738);
or U15886 (N_15886,N_15618,N_15647);
nand U15887 (N_15887,N_15763,N_15655);
nor U15888 (N_15888,N_15635,N_15714);
nor U15889 (N_15889,N_15740,N_15710);
nand U15890 (N_15890,N_15659,N_15688);
or U15891 (N_15891,N_15765,N_15793);
nor U15892 (N_15892,N_15719,N_15799);
xnor U15893 (N_15893,N_15758,N_15621);
nor U15894 (N_15894,N_15773,N_15737);
xnor U15895 (N_15895,N_15640,N_15651);
and U15896 (N_15896,N_15783,N_15787);
nor U15897 (N_15897,N_15636,N_15739);
or U15898 (N_15898,N_15639,N_15686);
or U15899 (N_15899,N_15638,N_15681);
nor U15900 (N_15900,N_15708,N_15732);
xor U15901 (N_15901,N_15775,N_15623);
or U15902 (N_15902,N_15732,N_15687);
nor U15903 (N_15903,N_15604,N_15713);
nand U15904 (N_15904,N_15789,N_15695);
xor U15905 (N_15905,N_15728,N_15609);
nor U15906 (N_15906,N_15630,N_15736);
xnor U15907 (N_15907,N_15697,N_15744);
nor U15908 (N_15908,N_15621,N_15684);
nand U15909 (N_15909,N_15704,N_15747);
xor U15910 (N_15910,N_15650,N_15757);
nor U15911 (N_15911,N_15603,N_15654);
nor U15912 (N_15912,N_15738,N_15651);
nand U15913 (N_15913,N_15766,N_15741);
nor U15914 (N_15914,N_15686,N_15673);
nand U15915 (N_15915,N_15678,N_15633);
nor U15916 (N_15916,N_15650,N_15625);
xnor U15917 (N_15917,N_15680,N_15754);
nor U15918 (N_15918,N_15656,N_15666);
or U15919 (N_15919,N_15773,N_15612);
and U15920 (N_15920,N_15713,N_15667);
and U15921 (N_15921,N_15766,N_15773);
nor U15922 (N_15922,N_15604,N_15770);
and U15923 (N_15923,N_15692,N_15737);
xnor U15924 (N_15924,N_15603,N_15625);
nor U15925 (N_15925,N_15649,N_15799);
nand U15926 (N_15926,N_15647,N_15752);
and U15927 (N_15927,N_15773,N_15664);
xnor U15928 (N_15928,N_15719,N_15674);
or U15929 (N_15929,N_15671,N_15756);
or U15930 (N_15930,N_15761,N_15729);
xnor U15931 (N_15931,N_15746,N_15702);
or U15932 (N_15932,N_15740,N_15777);
xnor U15933 (N_15933,N_15690,N_15705);
nand U15934 (N_15934,N_15622,N_15741);
xnor U15935 (N_15935,N_15642,N_15637);
and U15936 (N_15936,N_15734,N_15772);
and U15937 (N_15937,N_15681,N_15662);
and U15938 (N_15938,N_15636,N_15658);
xor U15939 (N_15939,N_15632,N_15728);
nand U15940 (N_15940,N_15635,N_15615);
nor U15941 (N_15941,N_15620,N_15608);
nor U15942 (N_15942,N_15615,N_15725);
and U15943 (N_15943,N_15638,N_15702);
or U15944 (N_15944,N_15715,N_15681);
and U15945 (N_15945,N_15614,N_15743);
xnor U15946 (N_15946,N_15732,N_15753);
and U15947 (N_15947,N_15636,N_15784);
nand U15948 (N_15948,N_15628,N_15725);
nor U15949 (N_15949,N_15716,N_15754);
nand U15950 (N_15950,N_15769,N_15671);
nand U15951 (N_15951,N_15668,N_15601);
nand U15952 (N_15952,N_15724,N_15682);
nor U15953 (N_15953,N_15679,N_15618);
xnor U15954 (N_15954,N_15690,N_15798);
nor U15955 (N_15955,N_15713,N_15644);
or U15956 (N_15956,N_15743,N_15699);
nor U15957 (N_15957,N_15639,N_15625);
nand U15958 (N_15958,N_15665,N_15641);
and U15959 (N_15959,N_15604,N_15619);
or U15960 (N_15960,N_15655,N_15754);
xnor U15961 (N_15961,N_15651,N_15751);
or U15962 (N_15962,N_15753,N_15733);
nor U15963 (N_15963,N_15697,N_15640);
xnor U15964 (N_15964,N_15670,N_15626);
or U15965 (N_15965,N_15623,N_15622);
nand U15966 (N_15966,N_15776,N_15628);
or U15967 (N_15967,N_15740,N_15760);
nor U15968 (N_15968,N_15709,N_15740);
and U15969 (N_15969,N_15670,N_15780);
nand U15970 (N_15970,N_15656,N_15719);
xor U15971 (N_15971,N_15734,N_15643);
or U15972 (N_15972,N_15630,N_15794);
xnor U15973 (N_15973,N_15610,N_15773);
xor U15974 (N_15974,N_15655,N_15640);
xnor U15975 (N_15975,N_15773,N_15777);
nor U15976 (N_15976,N_15617,N_15648);
nand U15977 (N_15977,N_15680,N_15718);
and U15978 (N_15978,N_15691,N_15770);
and U15979 (N_15979,N_15652,N_15606);
and U15980 (N_15980,N_15720,N_15749);
nand U15981 (N_15981,N_15797,N_15736);
or U15982 (N_15982,N_15626,N_15744);
nor U15983 (N_15983,N_15692,N_15675);
nor U15984 (N_15984,N_15648,N_15768);
nand U15985 (N_15985,N_15649,N_15753);
or U15986 (N_15986,N_15618,N_15709);
or U15987 (N_15987,N_15710,N_15755);
and U15988 (N_15988,N_15612,N_15609);
nor U15989 (N_15989,N_15763,N_15686);
xnor U15990 (N_15990,N_15657,N_15683);
nor U15991 (N_15991,N_15633,N_15625);
or U15992 (N_15992,N_15731,N_15751);
and U15993 (N_15993,N_15796,N_15626);
and U15994 (N_15994,N_15749,N_15612);
nand U15995 (N_15995,N_15780,N_15773);
nor U15996 (N_15996,N_15784,N_15731);
or U15997 (N_15997,N_15745,N_15649);
and U15998 (N_15998,N_15747,N_15676);
and U15999 (N_15999,N_15730,N_15626);
and U16000 (N_16000,N_15800,N_15857);
nand U16001 (N_16001,N_15966,N_15894);
nand U16002 (N_16002,N_15917,N_15918);
and U16003 (N_16003,N_15981,N_15958);
or U16004 (N_16004,N_15906,N_15916);
and U16005 (N_16005,N_15880,N_15960);
or U16006 (N_16006,N_15867,N_15998);
xor U16007 (N_16007,N_15909,N_15869);
and U16008 (N_16008,N_15914,N_15812);
nor U16009 (N_16009,N_15984,N_15919);
nand U16010 (N_16010,N_15945,N_15961);
nand U16011 (N_16011,N_15992,N_15938);
and U16012 (N_16012,N_15892,N_15991);
xor U16013 (N_16013,N_15922,N_15833);
xnor U16014 (N_16014,N_15925,N_15935);
nand U16015 (N_16015,N_15969,N_15811);
xor U16016 (N_16016,N_15996,N_15801);
or U16017 (N_16017,N_15926,N_15878);
nor U16018 (N_16018,N_15974,N_15897);
or U16019 (N_16019,N_15825,N_15884);
nor U16020 (N_16020,N_15809,N_15879);
and U16021 (N_16021,N_15826,N_15828);
and U16022 (N_16022,N_15872,N_15893);
nor U16023 (N_16023,N_15865,N_15881);
nand U16024 (N_16024,N_15939,N_15837);
or U16025 (N_16025,N_15967,N_15844);
nand U16026 (N_16026,N_15882,N_15806);
nand U16027 (N_16027,N_15995,N_15810);
or U16028 (N_16028,N_15987,N_15861);
and U16029 (N_16029,N_15986,N_15920);
nor U16030 (N_16030,N_15823,N_15830);
nand U16031 (N_16031,N_15994,N_15968);
xor U16032 (N_16032,N_15942,N_15862);
nor U16033 (N_16033,N_15807,N_15817);
xnor U16034 (N_16034,N_15885,N_15999);
nand U16035 (N_16035,N_15965,N_15864);
nor U16036 (N_16036,N_15820,N_15927);
and U16037 (N_16037,N_15835,N_15886);
nand U16038 (N_16038,N_15977,N_15962);
and U16039 (N_16039,N_15841,N_15854);
nand U16040 (N_16040,N_15888,N_15921);
and U16041 (N_16041,N_15950,N_15815);
nand U16042 (N_16042,N_15976,N_15898);
nand U16043 (N_16043,N_15954,N_15838);
or U16044 (N_16044,N_15808,N_15863);
xor U16045 (N_16045,N_15870,N_15911);
xor U16046 (N_16046,N_15849,N_15816);
xnor U16047 (N_16047,N_15860,N_15840);
or U16048 (N_16048,N_15923,N_15947);
and U16049 (N_16049,N_15902,N_15813);
nor U16050 (N_16050,N_15877,N_15946);
or U16051 (N_16051,N_15876,N_15932);
nor U16052 (N_16052,N_15842,N_15929);
or U16053 (N_16053,N_15940,N_15943);
nand U16054 (N_16054,N_15871,N_15912);
nor U16055 (N_16055,N_15821,N_15874);
nand U16056 (N_16056,N_15802,N_15983);
and U16057 (N_16057,N_15953,N_15901);
xor U16058 (N_16058,N_15824,N_15819);
or U16059 (N_16059,N_15952,N_15889);
nand U16060 (N_16060,N_15964,N_15941);
and U16061 (N_16061,N_15899,N_15818);
nand U16062 (N_16062,N_15924,N_15890);
nor U16063 (N_16063,N_15937,N_15805);
xor U16064 (N_16064,N_15956,N_15915);
xnor U16065 (N_16065,N_15803,N_15848);
xor U16066 (N_16066,N_15887,N_15804);
and U16067 (N_16067,N_15907,N_15910);
or U16068 (N_16068,N_15936,N_15883);
nand U16069 (N_16069,N_15847,N_15970);
nor U16070 (N_16070,N_15829,N_15949);
nor U16071 (N_16071,N_15957,N_15948);
xnor U16072 (N_16072,N_15858,N_15856);
nand U16073 (N_16073,N_15839,N_15988);
xnor U16074 (N_16074,N_15827,N_15908);
or U16075 (N_16075,N_15982,N_15933);
xnor U16076 (N_16076,N_15875,N_15853);
nand U16077 (N_16077,N_15891,N_15980);
and U16078 (N_16078,N_15973,N_15903);
and U16079 (N_16079,N_15834,N_15866);
xor U16080 (N_16080,N_15997,N_15905);
and U16081 (N_16081,N_15993,N_15934);
xnor U16082 (N_16082,N_15895,N_15944);
nor U16083 (N_16083,N_15930,N_15843);
nor U16084 (N_16084,N_15959,N_15989);
xnor U16085 (N_16085,N_15836,N_15900);
nor U16086 (N_16086,N_15850,N_15928);
nor U16087 (N_16087,N_15978,N_15831);
or U16088 (N_16088,N_15955,N_15814);
xor U16089 (N_16089,N_15963,N_15985);
xnor U16090 (N_16090,N_15859,N_15868);
and U16091 (N_16091,N_15832,N_15855);
or U16092 (N_16092,N_15845,N_15822);
or U16093 (N_16093,N_15846,N_15851);
nor U16094 (N_16094,N_15896,N_15904);
nor U16095 (N_16095,N_15852,N_15913);
and U16096 (N_16096,N_15951,N_15979);
and U16097 (N_16097,N_15972,N_15931);
nand U16098 (N_16098,N_15975,N_15971);
and U16099 (N_16099,N_15990,N_15873);
xor U16100 (N_16100,N_15932,N_15840);
and U16101 (N_16101,N_15910,N_15952);
and U16102 (N_16102,N_15806,N_15819);
nand U16103 (N_16103,N_15940,N_15904);
nor U16104 (N_16104,N_15837,N_15817);
nand U16105 (N_16105,N_15883,N_15956);
and U16106 (N_16106,N_15974,N_15874);
nor U16107 (N_16107,N_15905,N_15844);
or U16108 (N_16108,N_15933,N_15973);
xor U16109 (N_16109,N_15882,N_15976);
nand U16110 (N_16110,N_15988,N_15853);
nand U16111 (N_16111,N_15800,N_15933);
or U16112 (N_16112,N_15875,N_15898);
and U16113 (N_16113,N_15810,N_15868);
nor U16114 (N_16114,N_15916,N_15861);
xnor U16115 (N_16115,N_15821,N_15985);
nand U16116 (N_16116,N_15884,N_15800);
and U16117 (N_16117,N_15875,N_15904);
and U16118 (N_16118,N_15864,N_15866);
xnor U16119 (N_16119,N_15988,N_15814);
xnor U16120 (N_16120,N_15984,N_15998);
nor U16121 (N_16121,N_15840,N_15952);
or U16122 (N_16122,N_15990,N_15994);
or U16123 (N_16123,N_15801,N_15831);
xor U16124 (N_16124,N_15821,N_15856);
xor U16125 (N_16125,N_15988,N_15911);
nand U16126 (N_16126,N_15801,N_15968);
xor U16127 (N_16127,N_15865,N_15908);
xor U16128 (N_16128,N_15825,N_15858);
nor U16129 (N_16129,N_15930,N_15934);
nand U16130 (N_16130,N_15953,N_15842);
xor U16131 (N_16131,N_15966,N_15809);
nand U16132 (N_16132,N_15889,N_15896);
nand U16133 (N_16133,N_15998,N_15877);
or U16134 (N_16134,N_15900,N_15807);
nor U16135 (N_16135,N_15842,N_15934);
xor U16136 (N_16136,N_15950,N_15820);
nor U16137 (N_16137,N_15972,N_15889);
nor U16138 (N_16138,N_15990,N_15894);
nand U16139 (N_16139,N_15989,N_15903);
xnor U16140 (N_16140,N_15898,N_15973);
nand U16141 (N_16141,N_15953,N_15829);
nor U16142 (N_16142,N_15976,N_15910);
or U16143 (N_16143,N_15913,N_15806);
nand U16144 (N_16144,N_15859,N_15912);
or U16145 (N_16145,N_15949,N_15989);
nand U16146 (N_16146,N_15936,N_15977);
nand U16147 (N_16147,N_15975,N_15834);
xor U16148 (N_16148,N_15823,N_15964);
nor U16149 (N_16149,N_15831,N_15901);
nand U16150 (N_16150,N_15937,N_15861);
and U16151 (N_16151,N_15955,N_15924);
or U16152 (N_16152,N_15935,N_15845);
nand U16153 (N_16153,N_15873,N_15931);
nor U16154 (N_16154,N_15995,N_15888);
nand U16155 (N_16155,N_15877,N_15848);
or U16156 (N_16156,N_15898,N_15887);
nor U16157 (N_16157,N_15915,N_15870);
nor U16158 (N_16158,N_15990,N_15844);
or U16159 (N_16159,N_15876,N_15822);
xor U16160 (N_16160,N_15982,N_15883);
and U16161 (N_16161,N_15956,N_15868);
nor U16162 (N_16162,N_15928,N_15899);
and U16163 (N_16163,N_15940,N_15822);
and U16164 (N_16164,N_15996,N_15979);
and U16165 (N_16165,N_15874,N_15851);
xnor U16166 (N_16166,N_15822,N_15886);
nor U16167 (N_16167,N_15919,N_15982);
or U16168 (N_16168,N_15961,N_15807);
and U16169 (N_16169,N_15901,N_15911);
nand U16170 (N_16170,N_15861,N_15830);
xnor U16171 (N_16171,N_15897,N_15930);
and U16172 (N_16172,N_15956,N_15866);
nand U16173 (N_16173,N_15841,N_15928);
and U16174 (N_16174,N_15829,N_15989);
or U16175 (N_16175,N_15934,N_15818);
and U16176 (N_16176,N_15916,N_15985);
and U16177 (N_16177,N_15967,N_15871);
and U16178 (N_16178,N_15935,N_15862);
xor U16179 (N_16179,N_15925,N_15996);
or U16180 (N_16180,N_15807,N_15878);
or U16181 (N_16181,N_15953,N_15997);
and U16182 (N_16182,N_15871,N_15937);
or U16183 (N_16183,N_15860,N_15900);
or U16184 (N_16184,N_15956,N_15923);
or U16185 (N_16185,N_15829,N_15864);
and U16186 (N_16186,N_15976,N_15964);
and U16187 (N_16187,N_15950,N_15933);
xor U16188 (N_16188,N_15870,N_15910);
xnor U16189 (N_16189,N_15885,N_15997);
nand U16190 (N_16190,N_15841,N_15941);
and U16191 (N_16191,N_15856,N_15908);
nand U16192 (N_16192,N_15964,N_15993);
nand U16193 (N_16193,N_15827,N_15880);
and U16194 (N_16194,N_15897,N_15978);
nor U16195 (N_16195,N_15955,N_15968);
nor U16196 (N_16196,N_15809,N_15943);
and U16197 (N_16197,N_15868,N_15836);
or U16198 (N_16198,N_15885,N_15899);
and U16199 (N_16199,N_15951,N_15925);
and U16200 (N_16200,N_16051,N_16150);
xor U16201 (N_16201,N_16019,N_16186);
xnor U16202 (N_16202,N_16118,N_16086);
and U16203 (N_16203,N_16030,N_16010);
xor U16204 (N_16204,N_16199,N_16114);
nor U16205 (N_16205,N_16140,N_16029);
nand U16206 (N_16206,N_16185,N_16097);
nor U16207 (N_16207,N_16164,N_16165);
or U16208 (N_16208,N_16149,N_16141);
xnor U16209 (N_16209,N_16128,N_16002);
or U16210 (N_16210,N_16139,N_16171);
xnor U16211 (N_16211,N_16194,N_16087);
xor U16212 (N_16212,N_16197,N_16060);
and U16213 (N_16213,N_16179,N_16028);
nor U16214 (N_16214,N_16110,N_16191);
xor U16215 (N_16215,N_16162,N_16154);
nand U16216 (N_16216,N_16063,N_16023);
xnor U16217 (N_16217,N_16046,N_16190);
nor U16218 (N_16218,N_16070,N_16104);
nor U16219 (N_16219,N_16142,N_16178);
and U16220 (N_16220,N_16092,N_16084);
xnor U16221 (N_16221,N_16182,N_16135);
or U16222 (N_16222,N_16069,N_16036);
xor U16223 (N_16223,N_16188,N_16033);
xnor U16224 (N_16224,N_16088,N_16056);
and U16225 (N_16225,N_16173,N_16172);
xor U16226 (N_16226,N_16168,N_16007);
nor U16227 (N_16227,N_16044,N_16055);
and U16228 (N_16228,N_16032,N_16038);
xor U16229 (N_16229,N_16027,N_16059);
or U16230 (N_16230,N_16057,N_16037);
nand U16231 (N_16231,N_16094,N_16120);
or U16232 (N_16232,N_16054,N_16126);
xor U16233 (N_16233,N_16123,N_16147);
xor U16234 (N_16234,N_16012,N_16052);
xnor U16235 (N_16235,N_16144,N_16025);
or U16236 (N_16236,N_16107,N_16176);
nor U16237 (N_16237,N_16050,N_16167);
xor U16238 (N_16238,N_16133,N_16064);
xor U16239 (N_16239,N_16014,N_16130);
or U16240 (N_16240,N_16075,N_16122);
or U16241 (N_16241,N_16161,N_16196);
and U16242 (N_16242,N_16192,N_16151);
nor U16243 (N_16243,N_16058,N_16145);
nor U16244 (N_16244,N_16006,N_16041);
xor U16245 (N_16245,N_16068,N_16066);
and U16246 (N_16246,N_16153,N_16187);
and U16247 (N_16247,N_16136,N_16105);
nor U16248 (N_16248,N_16170,N_16053);
or U16249 (N_16249,N_16001,N_16072);
nand U16250 (N_16250,N_16089,N_16106);
nand U16251 (N_16251,N_16184,N_16061);
or U16252 (N_16252,N_16183,N_16100);
and U16253 (N_16253,N_16174,N_16078);
and U16254 (N_16254,N_16049,N_16015);
nor U16255 (N_16255,N_16091,N_16022);
xor U16256 (N_16256,N_16040,N_16125);
xor U16257 (N_16257,N_16198,N_16143);
nor U16258 (N_16258,N_16166,N_16152);
and U16259 (N_16259,N_16035,N_16071);
xnor U16260 (N_16260,N_16129,N_16109);
or U16261 (N_16261,N_16117,N_16079);
or U16262 (N_16262,N_16031,N_16175);
xor U16263 (N_16263,N_16074,N_16156);
nor U16264 (N_16264,N_16034,N_16039);
xnor U16265 (N_16265,N_16138,N_16108);
or U16266 (N_16266,N_16062,N_16124);
or U16267 (N_16267,N_16111,N_16047);
and U16268 (N_16268,N_16065,N_16096);
nand U16269 (N_16269,N_16000,N_16017);
nor U16270 (N_16270,N_16116,N_16160);
nor U16271 (N_16271,N_16157,N_16132);
xnor U16272 (N_16272,N_16093,N_16146);
xnor U16273 (N_16273,N_16180,N_16021);
or U16274 (N_16274,N_16077,N_16181);
or U16275 (N_16275,N_16011,N_16131);
xor U16276 (N_16276,N_16102,N_16177);
or U16277 (N_16277,N_16013,N_16026);
nor U16278 (N_16278,N_16073,N_16134);
or U16279 (N_16279,N_16169,N_16195);
or U16280 (N_16280,N_16101,N_16018);
nor U16281 (N_16281,N_16043,N_16189);
or U16282 (N_16282,N_16005,N_16081);
xnor U16283 (N_16283,N_16083,N_16042);
xor U16284 (N_16284,N_16158,N_16137);
xnor U16285 (N_16285,N_16148,N_16085);
and U16286 (N_16286,N_16008,N_16113);
nand U16287 (N_16287,N_16067,N_16090);
or U16288 (N_16288,N_16016,N_16127);
nor U16289 (N_16289,N_16121,N_16004);
xor U16290 (N_16290,N_16076,N_16099);
nor U16291 (N_16291,N_16163,N_16119);
or U16292 (N_16292,N_16155,N_16082);
xnor U16293 (N_16293,N_16098,N_16024);
and U16294 (N_16294,N_16112,N_16045);
xor U16295 (N_16295,N_16193,N_16009);
or U16296 (N_16296,N_16095,N_16003);
xor U16297 (N_16297,N_16159,N_16048);
nand U16298 (N_16298,N_16020,N_16115);
or U16299 (N_16299,N_16103,N_16080);
xor U16300 (N_16300,N_16097,N_16107);
or U16301 (N_16301,N_16044,N_16130);
nand U16302 (N_16302,N_16017,N_16196);
or U16303 (N_16303,N_16081,N_16047);
nor U16304 (N_16304,N_16074,N_16188);
xor U16305 (N_16305,N_16049,N_16050);
nor U16306 (N_16306,N_16056,N_16024);
nand U16307 (N_16307,N_16001,N_16074);
xor U16308 (N_16308,N_16105,N_16038);
and U16309 (N_16309,N_16095,N_16178);
nor U16310 (N_16310,N_16025,N_16142);
xor U16311 (N_16311,N_16085,N_16033);
and U16312 (N_16312,N_16145,N_16106);
nand U16313 (N_16313,N_16133,N_16194);
xor U16314 (N_16314,N_16122,N_16004);
nand U16315 (N_16315,N_16033,N_16064);
and U16316 (N_16316,N_16147,N_16165);
or U16317 (N_16317,N_16109,N_16111);
nor U16318 (N_16318,N_16181,N_16019);
or U16319 (N_16319,N_16018,N_16181);
nand U16320 (N_16320,N_16079,N_16099);
or U16321 (N_16321,N_16109,N_16160);
or U16322 (N_16322,N_16139,N_16145);
nand U16323 (N_16323,N_16008,N_16172);
xnor U16324 (N_16324,N_16198,N_16040);
nor U16325 (N_16325,N_16075,N_16191);
xnor U16326 (N_16326,N_16169,N_16128);
xnor U16327 (N_16327,N_16076,N_16111);
and U16328 (N_16328,N_16050,N_16052);
or U16329 (N_16329,N_16099,N_16041);
nand U16330 (N_16330,N_16038,N_16179);
and U16331 (N_16331,N_16027,N_16072);
nand U16332 (N_16332,N_16073,N_16135);
xor U16333 (N_16333,N_16112,N_16004);
nand U16334 (N_16334,N_16028,N_16046);
nand U16335 (N_16335,N_16194,N_16184);
nand U16336 (N_16336,N_16035,N_16093);
or U16337 (N_16337,N_16189,N_16152);
xor U16338 (N_16338,N_16038,N_16187);
xor U16339 (N_16339,N_16035,N_16125);
or U16340 (N_16340,N_16020,N_16106);
or U16341 (N_16341,N_16098,N_16121);
nand U16342 (N_16342,N_16061,N_16104);
xor U16343 (N_16343,N_16100,N_16136);
xor U16344 (N_16344,N_16169,N_16072);
nor U16345 (N_16345,N_16041,N_16005);
or U16346 (N_16346,N_16191,N_16034);
or U16347 (N_16347,N_16019,N_16116);
or U16348 (N_16348,N_16120,N_16013);
xor U16349 (N_16349,N_16123,N_16161);
nand U16350 (N_16350,N_16073,N_16032);
and U16351 (N_16351,N_16126,N_16051);
and U16352 (N_16352,N_16015,N_16021);
xor U16353 (N_16353,N_16002,N_16059);
nor U16354 (N_16354,N_16094,N_16182);
nand U16355 (N_16355,N_16090,N_16194);
or U16356 (N_16356,N_16063,N_16001);
xor U16357 (N_16357,N_16044,N_16010);
xor U16358 (N_16358,N_16082,N_16099);
or U16359 (N_16359,N_16198,N_16086);
xnor U16360 (N_16360,N_16030,N_16196);
nor U16361 (N_16361,N_16194,N_16118);
xor U16362 (N_16362,N_16175,N_16121);
nand U16363 (N_16363,N_16151,N_16050);
nand U16364 (N_16364,N_16174,N_16083);
or U16365 (N_16365,N_16166,N_16126);
xor U16366 (N_16366,N_16129,N_16103);
and U16367 (N_16367,N_16115,N_16191);
nand U16368 (N_16368,N_16030,N_16142);
nor U16369 (N_16369,N_16002,N_16077);
xor U16370 (N_16370,N_16081,N_16044);
and U16371 (N_16371,N_16078,N_16088);
or U16372 (N_16372,N_16050,N_16105);
xor U16373 (N_16373,N_16111,N_16145);
and U16374 (N_16374,N_16085,N_16127);
and U16375 (N_16375,N_16137,N_16043);
and U16376 (N_16376,N_16107,N_16154);
and U16377 (N_16377,N_16104,N_16078);
nor U16378 (N_16378,N_16052,N_16009);
xnor U16379 (N_16379,N_16117,N_16133);
or U16380 (N_16380,N_16073,N_16008);
nand U16381 (N_16381,N_16156,N_16020);
nand U16382 (N_16382,N_16128,N_16031);
nand U16383 (N_16383,N_16000,N_16112);
or U16384 (N_16384,N_16093,N_16172);
nor U16385 (N_16385,N_16058,N_16075);
and U16386 (N_16386,N_16162,N_16012);
nor U16387 (N_16387,N_16193,N_16129);
nand U16388 (N_16388,N_16004,N_16052);
xor U16389 (N_16389,N_16160,N_16016);
nand U16390 (N_16390,N_16188,N_16122);
nor U16391 (N_16391,N_16063,N_16050);
nor U16392 (N_16392,N_16180,N_16072);
xor U16393 (N_16393,N_16167,N_16079);
or U16394 (N_16394,N_16167,N_16122);
and U16395 (N_16395,N_16152,N_16055);
nand U16396 (N_16396,N_16129,N_16043);
nor U16397 (N_16397,N_16072,N_16131);
xor U16398 (N_16398,N_16084,N_16094);
nor U16399 (N_16399,N_16140,N_16193);
nor U16400 (N_16400,N_16242,N_16248);
nor U16401 (N_16401,N_16228,N_16296);
or U16402 (N_16402,N_16222,N_16357);
nand U16403 (N_16403,N_16201,N_16306);
or U16404 (N_16404,N_16257,N_16331);
nor U16405 (N_16405,N_16313,N_16351);
and U16406 (N_16406,N_16226,N_16301);
and U16407 (N_16407,N_16227,N_16220);
and U16408 (N_16408,N_16346,N_16305);
nor U16409 (N_16409,N_16349,N_16369);
xnor U16410 (N_16410,N_16241,N_16310);
nor U16411 (N_16411,N_16332,N_16327);
nand U16412 (N_16412,N_16283,N_16221);
xnor U16413 (N_16413,N_16267,N_16224);
xor U16414 (N_16414,N_16352,N_16318);
nand U16415 (N_16415,N_16236,N_16270);
and U16416 (N_16416,N_16340,N_16384);
xor U16417 (N_16417,N_16280,N_16303);
and U16418 (N_16418,N_16254,N_16304);
nand U16419 (N_16419,N_16363,N_16311);
nand U16420 (N_16420,N_16354,N_16339);
xnor U16421 (N_16421,N_16381,N_16335);
or U16422 (N_16422,N_16288,N_16324);
nor U16423 (N_16423,N_16343,N_16292);
nand U16424 (N_16424,N_16252,N_16309);
or U16425 (N_16425,N_16266,N_16277);
and U16426 (N_16426,N_16230,N_16265);
or U16427 (N_16427,N_16203,N_16247);
xor U16428 (N_16428,N_16202,N_16263);
nor U16429 (N_16429,N_16359,N_16218);
nor U16430 (N_16430,N_16366,N_16232);
nand U16431 (N_16431,N_16214,N_16328);
nand U16432 (N_16432,N_16312,N_16205);
nor U16433 (N_16433,N_16209,N_16294);
and U16434 (N_16434,N_16361,N_16200);
nor U16435 (N_16435,N_16207,N_16269);
nor U16436 (N_16436,N_16317,N_16374);
xnor U16437 (N_16437,N_16278,N_16396);
nor U16438 (N_16438,N_16275,N_16212);
or U16439 (N_16439,N_16285,N_16326);
and U16440 (N_16440,N_16211,N_16382);
xnor U16441 (N_16441,N_16379,N_16219);
or U16442 (N_16442,N_16264,N_16344);
and U16443 (N_16443,N_16385,N_16245);
nand U16444 (N_16444,N_16253,N_16355);
nor U16445 (N_16445,N_16323,N_16386);
xor U16446 (N_16446,N_16330,N_16376);
and U16447 (N_16447,N_16213,N_16238);
or U16448 (N_16448,N_16320,N_16215);
or U16449 (N_16449,N_16286,N_16276);
nand U16450 (N_16450,N_16334,N_16290);
nand U16451 (N_16451,N_16373,N_16314);
xor U16452 (N_16452,N_16325,N_16341);
or U16453 (N_16453,N_16258,N_16279);
and U16454 (N_16454,N_16353,N_16239);
nor U16455 (N_16455,N_16260,N_16293);
nor U16456 (N_16456,N_16240,N_16393);
nor U16457 (N_16457,N_16235,N_16365);
or U16458 (N_16458,N_16300,N_16210);
xnor U16459 (N_16459,N_16298,N_16388);
and U16460 (N_16460,N_16255,N_16399);
xnor U16461 (N_16461,N_16249,N_16299);
and U16462 (N_16462,N_16234,N_16225);
nand U16463 (N_16463,N_16336,N_16380);
or U16464 (N_16464,N_16356,N_16295);
nand U16465 (N_16465,N_16217,N_16364);
nor U16466 (N_16466,N_16259,N_16329);
xnor U16467 (N_16467,N_16243,N_16395);
nor U16468 (N_16468,N_16272,N_16345);
xnor U16469 (N_16469,N_16397,N_16237);
xnor U16470 (N_16470,N_16370,N_16389);
or U16471 (N_16471,N_16291,N_16246);
or U16472 (N_16472,N_16244,N_16256);
xor U16473 (N_16473,N_16342,N_16204);
and U16474 (N_16474,N_16316,N_16321);
xor U16475 (N_16475,N_16289,N_16208);
nor U16476 (N_16476,N_16368,N_16375);
or U16477 (N_16477,N_16297,N_16231);
xor U16478 (N_16478,N_16308,N_16302);
nand U16479 (N_16479,N_16282,N_16372);
or U16480 (N_16480,N_16281,N_16333);
or U16481 (N_16481,N_16387,N_16315);
or U16482 (N_16482,N_16261,N_16391);
or U16483 (N_16483,N_16362,N_16268);
or U16484 (N_16484,N_16337,N_16358);
and U16485 (N_16485,N_16319,N_16371);
nor U16486 (N_16486,N_16274,N_16273);
nand U16487 (N_16487,N_16390,N_16347);
nand U16488 (N_16488,N_16350,N_16307);
xnor U16489 (N_16489,N_16392,N_16206);
and U16490 (N_16490,N_16377,N_16338);
and U16491 (N_16491,N_16322,N_16216);
and U16492 (N_16492,N_16287,N_16251);
xor U16493 (N_16493,N_16394,N_16233);
xnor U16494 (N_16494,N_16383,N_16398);
or U16495 (N_16495,N_16229,N_16367);
nand U16496 (N_16496,N_16378,N_16223);
xor U16497 (N_16497,N_16250,N_16271);
xnor U16498 (N_16498,N_16348,N_16284);
nor U16499 (N_16499,N_16360,N_16262);
xor U16500 (N_16500,N_16214,N_16277);
nand U16501 (N_16501,N_16236,N_16356);
nand U16502 (N_16502,N_16395,N_16389);
and U16503 (N_16503,N_16290,N_16305);
and U16504 (N_16504,N_16313,N_16250);
nand U16505 (N_16505,N_16257,N_16344);
and U16506 (N_16506,N_16204,N_16372);
or U16507 (N_16507,N_16371,N_16283);
and U16508 (N_16508,N_16374,N_16378);
xor U16509 (N_16509,N_16218,N_16312);
or U16510 (N_16510,N_16350,N_16397);
and U16511 (N_16511,N_16282,N_16272);
nand U16512 (N_16512,N_16292,N_16283);
nand U16513 (N_16513,N_16256,N_16336);
and U16514 (N_16514,N_16317,N_16216);
nor U16515 (N_16515,N_16368,N_16315);
nor U16516 (N_16516,N_16289,N_16398);
nor U16517 (N_16517,N_16212,N_16374);
nand U16518 (N_16518,N_16331,N_16259);
and U16519 (N_16519,N_16328,N_16394);
or U16520 (N_16520,N_16336,N_16371);
and U16521 (N_16521,N_16243,N_16269);
nand U16522 (N_16522,N_16271,N_16358);
xnor U16523 (N_16523,N_16217,N_16220);
nand U16524 (N_16524,N_16244,N_16286);
xnor U16525 (N_16525,N_16278,N_16266);
nor U16526 (N_16526,N_16316,N_16327);
and U16527 (N_16527,N_16303,N_16398);
nor U16528 (N_16528,N_16335,N_16283);
xnor U16529 (N_16529,N_16291,N_16224);
xor U16530 (N_16530,N_16367,N_16318);
or U16531 (N_16531,N_16285,N_16354);
nand U16532 (N_16532,N_16268,N_16363);
nor U16533 (N_16533,N_16330,N_16205);
xnor U16534 (N_16534,N_16387,N_16260);
nand U16535 (N_16535,N_16397,N_16289);
nand U16536 (N_16536,N_16325,N_16254);
or U16537 (N_16537,N_16394,N_16254);
nand U16538 (N_16538,N_16335,N_16234);
nand U16539 (N_16539,N_16288,N_16320);
and U16540 (N_16540,N_16397,N_16296);
and U16541 (N_16541,N_16360,N_16208);
nand U16542 (N_16542,N_16262,N_16286);
and U16543 (N_16543,N_16357,N_16261);
or U16544 (N_16544,N_16352,N_16365);
nor U16545 (N_16545,N_16228,N_16202);
xor U16546 (N_16546,N_16262,N_16355);
nand U16547 (N_16547,N_16212,N_16223);
and U16548 (N_16548,N_16351,N_16268);
or U16549 (N_16549,N_16291,N_16388);
nor U16550 (N_16550,N_16229,N_16391);
xor U16551 (N_16551,N_16331,N_16296);
nand U16552 (N_16552,N_16246,N_16255);
and U16553 (N_16553,N_16356,N_16371);
xnor U16554 (N_16554,N_16218,N_16308);
nand U16555 (N_16555,N_16228,N_16298);
or U16556 (N_16556,N_16264,N_16230);
and U16557 (N_16557,N_16248,N_16332);
and U16558 (N_16558,N_16210,N_16317);
xor U16559 (N_16559,N_16217,N_16355);
nor U16560 (N_16560,N_16344,N_16355);
nand U16561 (N_16561,N_16362,N_16298);
nor U16562 (N_16562,N_16350,N_16281);
nand U16563 (N_16563,N_16337,N_16367);
nor U16564 (N_16564,N_16208,N_16397);
xor U16565 (N_16565,N_16385,N_16333);
nand U16566 (N_16566,N_16330,N_16351);
and U16567 (N_16567,N_16301,N_16311);
nand U16568 (N_16568,N_16279,N_16241);
nor U16569 (N_16569,N_16207,N_16364);
and U16570 (N_16570,N_16244,N_16384);
xor U16571 (N_16571,N_16329,N_16231);
or U16572 (N_16572,N_16310,N_16352);
nand U16573 (N_16573,N_16288,N_16281);
xnor U16574 (N_16574,N_16225,N_16301);
xor U16575 (N_16575,N_16214,N_16307);
and U16576 (N_16576,N_16336,N_16247);
nor U16577 (N_16577,N_16236,N_16287);
and U16578 (N_16578,N_16291,N_16272);
nor U16579 (N_16579,N_16243,N_16350);
nor U16580 (N_16580,N_16267,N_16309);
nor U16581 (N_16581,N_16337,N_16226);
and U16582 (N_16582,N_16393,N_16300);
nor U16583 (N_16583,N_16226,N_16371);
nor U16584 (N_16584,N_16346,N_16289);
nand U16585 (N_16585,N_16228,N_16378);
xnor U16586 (N_16586,N_16305,N_16292);
nor U16587 (N_16587,N_16328,N_16288);
or U16588 (N_16588,N_16232,N_16225);
and U16589 (N_16589,N_16225,N_16380);
nor U16590 (N_16590,N_16254,N_16363);
or U16591 (N_16591,N_16338,N_16254);
or U16592 (N_16592,N_16222,N_16377);
or U16593 (N_16593,N_16207,N_16342);
and U16594 (N_16594,N_16263,N_16372);
xnor U16595 (N_16595,N_16285,N_16281);
nor U16596 (N_16596,N_16383,N_16270);
or U16597 (N_16597,N_16345,N_16294);
nand U16598 (N_16598,N_16232,N_16284);
or U16599 (N_16599,N_16344,N_16309);
xor U16600 (N_16600,N_16532,N_16490);
xnor U16601 (N_16601,N_16593,N_16411);
nor U16602 (N_16602,N_16450,N_16464);
nor U16603 (N_16603,N_16418,N_16576);
nor U16604 (N_16604,N_16572,N_16534);
and U16605 (N_16605,N_16446,N_16567);
or U16606 (N_16606,N_16432,N_16546);
and U16607 (N_16607,N_16560,N_16586);
nor U16608 (N_16608,N_16400,N_16582);
or U16609 (N_16609,N_16438,N_16448);
and U16610 (N_16610,N_16456,N_16497);
nand U16611 (N_16611,N_16443,N_16519);
nor U16612 (N_16612,N_16581,N_16498);
nand U16613 (N_16613,N_16554,N_16547);
nor U16614 (N_16614,N_16536,N_16422);
and U16615 (N_16615,N_16590,N_16525);
and U16616 (N_16616,N_16406,N_16454);
nor U16617 (N_16617,N_16500,N_16439);
xnor U16618 (N_16618,N_16542,N_16410);
nand U16619 (N_16619,N_16452,N_16592);
and U16620 (N_16620,N_16583,N_16539);
and U16621 (N_16621,N_16477,N_16544);
or U16622 (N_16622,N_16495,N_16436);
nor U16623 (N_16623,N_16496,N_16549);
and U16624 (N_16624,N_16565,N_16468);
or U16625 (N_16625,N_16573,N_16433);
nor U16626 (N_16626,N_16598,N_16595);
xor U16627 (N_16627,N_16533,N_16543);
nand U16628 (N_16628,N_16538,N_16413);
and U16629 (N_16629,N_16574,N_16481);
xnor U16630 (N_16630,N_16509,N_16514);
and U16631 (N_16631,N_16556,N_16467);
and U16632 (N_16632,N_16491,N_16435);
or U16633 (N_16633,N_16486,N_16506);
nand U16634 (N_16634,N_16451,N_16522);
and U16635 (N_16635,N_16568,N_16471);
nor U16636 (N_16636,N_16409,N_16499);
xnor U16637 (N_16637,N_16537,N_16501);
nand U16638 (N_16638,N_16473,N_16578);
xor U16639 (N_16639,N_16445,N_16575);
nand U16640 (N_16640,N_16561,N_16466);
xnor U16641 (N_16641,N_16510,N_16531);
nand U16642 (N_16642,N_16417,N_16484);
and U16643 (N_16643,N_16427,N_16570);
and U16644 (N_16644,N_16447,N_16442);
nand U16645 (N_16645,N_16597,N_16548);
or U16646 (N_16646,N_16557,N_16588);
and U16647 (N_16647,N_16403,N_16479);
and U16648 (N_16648,N_16485,N_16455);
nand U16649 (N_16649,N_16414,N_16416);
or U16650 (N_16650,N_16434,N_16492);
xor U16651 (N_16651,N_16523,N_16505);
nor U16652 (N_16652,N_16419,N_16569);
xor U16653 (N_16653,N_16579,N_16515);
or U16654 (N_16654,N_16552,N_16502);
nand U16655 (N_16655,N_16440,N_16553);
nand U16656 (N_16656,N_16429,N_16437);
or U16657 (N_16657,N_16520,N_16401);
or U16658 (N_16658,N_16483,N_16420);
or U16659 (N_16659,N_16530,N_16404);
or U16660 (N_16660,N_16441,N_16585);
nand U16661 (N_16661,N_16504,N_16587);
nor U16662 (N_16662,N_16405,N_16462);
nor U16663 (N_16663,N_16472,N_16529);
xor U16664 (N_16664,N_16541,N_16562);
nor U16665 (N_16665,N_16550,N_16558);
nand U16666 (N_16666,N_16566,N_16545);
or U16667 (N_16667,N_16535,N_16402);
nor U16668 (N_16668,N_16470,N_16453);
nand U16669 (N_16669,N_16571,N_16596);
or U16670 (N_16670,N_16407,N_16518);
xor U16671 (N_16671,N_16559,N_16508);
nor U16672 (N_16672,N_16521,N_16457);
and U16673 (N_16673,N_16589,N_16503);
xnor U16674 (N_16674,N_16423,N_16459);
nand U16675 (N_16675,N_16421,N_16474);
nand U16676 (N_16676,N_16431,N_16577);
xor U16677 (N_16677,N_16480,N_16584);
nand U16678 (N_16678,N_16412,N_16424);
xor U16679 (N_16679,N_16488,N_16580);
or U16680 (N_16680,N_16415,N_16563);
xor U16681 (N_16681,N_16527,N_16524);
nand U16682 (N_16682,N_16460,N_16444);
xnor U16683 (N_16683,N_16458,N_16594);
xor U16684 (N_16684,N_16591,N_16526);
nand U16685 (N_16685,N_16540,N_16469);
or U16686 (N_16686,N_16428,N_16461);
nand U16687 (N_16687,N_16489,N_16507);
xnor U16688 (N_16688,N_16408,N_16516);
and U16689 (N_16689,N_16478,N_16512);
and U16690 (N_16690,N_16528,N_16555);
nand U16691 (N_16691,N_16513,N_16463);
nor U16692 (N_16692,N_16449,N_16482);
xor U16693 (N_16693,N_16426,N_16599);
or U16694 (N_16694,N_16475,N_16494);
nand U16695 (N_16695,N_16425,N_16493);
or U16696 (N_16696,N_16517,N_16476);
or U16697 (N_16697,N_16551,N_16430);
xor U16698 (N_16698,N_16487,N_16511);
and U16699 (N_16699,N_16465,N_16564);
xor U16700 (N_16700,N_16433,N_16402);
and U16701 (N_16701,N_16566,N_16426);
nand U16702 (N_16702,N_16537,N_16476);
nor U16703 (N_16703,N_16401,N_16471);
nand U16704 (N_16704,N_16497,N_16538);
nor U16705 (N_16705,N_16554,N_16468);
nand U16706 (N_16706,N_16588,N_16527);
and U16707 (N_16707,N_16508,N_16428);
xnor U16708 (N_16708,N_16531,N_16414);
nor U16709 (N_16709,N_16595,N_16438);
xnor U16710 (N_16710,N_16507,N_16593);
nand U16711 (N_16711,N_16488,N_16463);
or U16712 (N_16712,N_16510,N_16586);
and U16713 (N_16713,N_16468,N_16556);
nor U16714 (N_16714,N_16559,N_16550);
or U16715 (N_16715,N_16484,N_16425);
and U16716 (N_16716,N_16433,N_16465);
and U16717 (N_16717,N_16519,N_16482);
xor U16718 (N_16718,N_16481,N_16422);
xnor U16719 (N_16719,N_16474,N_16436);
xor U16720 (N_16720,N_16500,N_16429);
and U16721 (N_16721,N_16541,N_16411);
nand U16722 (N_16722,N_16581,N_16551);
and U16723 (N_16723,N_16437,N_16563);
or U16724 (N_16724,N_16538,N_16463);
nor U16725 (N_16725,N_16525,N_16577);
and U16726 (N_16726,N_16400,N_16597);
nor U16727 (N_16727,N_16569,N_16592);
and U16728 (N_16728,N_16468,N_16580);
nor U16729 (N_16729,N_16568,N_16436);
and U16730 (N_16730,N_16527,N_16587);
xnor U16731 (N_16731,N_16463,N_16559);
nor U16732 (N_16732,N_16496,N_16401);
or U16733 (N_16733,N_16414,N_16403);
nand U16734 (N_16734,N_16484,N_16409);
nor U16735 (N_16735,N_16401,N_16528);
and U16736 (N_16736,N_16481,N_16480);
or U16737 (N_16737,N_16407,N_16557);
xnor U16738 (N_16738,N_16428,N_16437);
and U16739 (N_16739,N_16458,N_16529);
and U16740 (N_16740,N_16507,N_16569);
or U16741 (N_16741,N_16509,N_16581);
or U16742 (N_16742,N_16415,N_16584);
nand U16743 (N_16743,N_16495,N_16554);
and U16744 (N_16744,N_16587,N_16519);
or U16745 (N_16745,N_16574,N_16419);
nor U16746 (N_16746,N_16552,N_16466);
and U16747 (N_16747,N_16432,N_16438);
and U16748 (N_16748,N_16596,N_16570);
nor U16749 (N_16749,N_16455,N_16478);
and U16750 (N_16750,N_16457,N_16537);
and U16751 (N_16751,N_16402,N_16428);
nor U16752 (N_16752,N_16460,N_16530);
and U16753 (N_16753,N_16541,N_16427);
nand U16754 (N_16754,N_16567,N_16532);
or U16755 (N_16755,N_16570,N_16450);
and U16756 (N_16756,N_16596,N_16560);
xnor U16757 (N_16757,N_16403,N_16472);
nand U16758 (N_16758,N_16553,N_16542);
and U16759 (N_16759,N_16478,N_16541);
nand U16760 (N_16760,N_16581,N_16450);
xnor U16761 (N_16761,N_16554,N_16483);
or U16762 (N_16762,N_16528,N_16499);
xor U16763 (N_16763,N_16513,N_16517);
nand U16764 (N_16764,N_16485,N_16448);
nor U16765 (N_16765,N_16486,N_16518);
and U16766 (N_16766,N_16553,N_16497);
and U16767 (N_16767,N_16587,N_16406);
or U16768 (N_16768,N_16597,N_16500);
nand U16769 (N_16769,N_16529,N_16592);
or U16770 (N_16770,N_16411,N_16487);
or U16771 (N_16771,N_16596,N_16435);
xor U16772 (N_16772,N_16552,N_16542);
xor U16773 (N_16773,N_16554,N_16415);
and U16774 (N_16774,N_16400,N_16517);
nor U16775 (N_16775,N_16505,N_16476);
nand U16776 (N_16776,N_16402,N_16499);
nand U16777 (N_16777,N_16400,N_16411);
nor U16778 (N_16778,N_16540,N_16495);
nor U16779 (N_16779,N_16424,N_16567);
or U16780 (N_16780,N_16453,N_16515);
and U16781 (N_16781,N_16560,N_16570);
nor U16782 (N_16782,N_16531,N_16457);
xnor U16783 (N_16783,N_16556,N_16551);
xnor U16784 (N_16784,N_16553,N_16400);
nor U16785 (N_16785,N_16597,N_16576);
or U16786 (N_16786,N_16422,N_16521);
xor U16787 (N_16787,N_16453,N_16467);
xor U16788 (N_16788,N_16553,N_16461);
nor U16789 (N_16789,N_16539,N_16574);
and U16790 (N_16790,N_16568,N_16403);
nor U16791 (N_16791,N_16429,N_16556);
xnor U16792 (N_16792,N_16459,N_16557);
and U16793 (N_16793,N_16558,N_16526);
xnor U16794 (N_16794,N_16526,N_16537);
nor U16795 (N_16795,N_16438,N_16460);
nand U16796 (N_16796,N_16574,N_16500);
xnor U16797 (N_16797,N_16579,N_16439);
nand U16798 (N_16798,N_16470,N_16478);
nor U16799 (N_16799,N_16585,N_16400);
and U16800 (N_16800,N_16787,N_16662);
nand U16801 (N_16801,N_16743,N_16775);
or U16802 (N_16802,N_16695,N_16698);
xor U16803 (N_16803,N_16643,N_16674);
and U16804 (N_16804,N_16622,N_16704);
and U16805 (N_16805,N_16628,N_16679);
nor U16806 (N_16806,N_16609,N_16686);
xnor U16807 (N_16807,N_16641,N_16760);
or U16808 (N_16808,N_16715,N_16640);
or U16809 (N_16809,N_16677,N_16734);
nand U16810 (N_16810,N_16619,N_16736);
and U16811 (N_16811,N_16711,N_16762);
nand U16812 (N_16812,N_16645,N_16696);
nor U16813 (N_16813,N_16751,N_16650);
nand U16814 (N_16814,N_16769,N_16719);
nand U16815 (N_16815,N_16726,N_16685);
xnor U16816 (N_16816,N_16700,N_16788);
nor U16817 (N_16817,N_16768,N_16735);
xor U16818 (N_16818,N_16697,N_16668);
or U16819 (N_16819,N_16728,N_16730);
nand U16820 (N_16820,N_16667,N_16746);
and U16821 (N_16821,N_16601,N_16745);
or U16822 (N_16822,N_16659,N_16618);
and U16823 (N_16823,N_16636,N_16765);
xnor U16824 (N_16824,N_16613,N_16727);
nand U16825 (N_16825,N_16779,N_16753);
nor U16826 (N_16826,N_16632,N_16615);
nor U16827 (N_16827,N_16720,N_16770);
or U16828 (N_16828,N_16690,N_16729);
nand U16829 (N_16829,N_16651,N_16612);
nand U16830 (N_16830,N_16757,N_16795);
nor U16831 (N_16831,N_16611,N_16713);
or U16832 (N_16832,N_16664,N_16732);
xor U16833 (N_16833,N_16773,N_16605);
xnor U16834 (N_16834,N_16623,N_16600);
and U16835 (N_16835,N_16687,N_16656);
nor U16836 (N_16836,N_16692,N_16742);
nand U16837 (N_16837,N_16693,N_16797);
nand U16838 (N_16838,N_16639,N_16716);
and U16839 (N_16839,N_16680,N_16764);
nor U16840 (N_16840,N_16792,N_16767);
nand U16841 (N_16841,N_16660,N_16657);
and U16842 (N_16842,N_16725,N_16722);
or U16843 (N_16843,N_16635,N_16776);
or U16844 (N_16844,N_16782,N_16748);
and U16845 (N_16845,N_16625,N_16781);
xor U16846 (N_16846,N_16670,N_16647);
nand U16847 (N_16847,N_16718,N_16608);
nor U16848 (N_16848,N_16627,N_16629);
and U16849 (N_16849,N_16783,N_16733);
and U16850 (N_16850,N_16793,N_16638);
and U16851 (N_16851,N_16705,N_16663);
xor U16852 (N_16852,N_16666,N_16750);
nand U16853 (N_16853,N_16702,N_16772);
nand U16854 (N_16854,N_16684,N_16791);
or U16855 (N_16855,N_16724,N_16766);
or U16856 (N_16856,N_16784,N_16780);
nand U16857 (N_16857,N_16610,N_16691);
and U16858 (N_16858,N_16708,N_16634);
and U16859 (N_16859,N_16644,N_16790);
or U16860 (N_16860,N_16631,N_16794);
nand U16861 (N_16861,N_16675,N_16789);
or U16862 (N_16862,N_16761,N_16739);
nand U16863 (N_16863,N_16703,N_16665);
nand U16864 (N_16864,N_16723,N_16777);
nand U16865 (N_16865,N_16652,N_16785);
nor U16866 (N_16866,N_16653,N_16778);
nor U16867 (N_16867,N_16706,N_16774);
nand U16868 (N_16868,N_16759,N_16688);
and U16869 (N_16869,N_16633,N_16683);
or U16870 (N_16870,N_16689,N_16626);
or U16871 (N_16871,N_16649,N_16669);
nor U16872 (N_16872,N_16630,N_16799);
xnor U16873 (N_16873,N_16603,N_16714);
xor U16874 (N_16874,N_16709,N_16604);
and U16875 (N_16875,N_16710,N_16681);
and U16876 (N_16876,N_16646,N_16771);
nor U16877 (N_16877,N_16607,N_16763);
or U16878 (N_16878,N_16655,N_16672);
or U16879 (N_16879,N_16614,N_16741);
xnor U16880 (N_16880,N_16740,N_16658);
nor U16881 (N_16881,N_16621,N_16701);
and U16882 (N_16882,N_16678,N_16620);
nor U16883 (N_16883,N_16747,N_16744);
xnor U16884 (N_16884,N_16648,N_16661);
nand U16885 (N_16885,N_16738,N_16717);
and U16886 (N_16886,N_16637,N_16682);
and U16887 (N_16887,N_16731,N_16699);
nor U16888 (N_16888,N_16712,N_16673);
nor U16889 (N_16889,N_16756,N_16671);
nand U16890 (N_16890,N_16654,N_16754);
xnor U16891 (N_16891,N_16737,N_16694);
nand U16892 (N_16892,N_16707,N_16624);
nand U16893 (N_16893,N_16606,N_16642);
nand U16894 (N_16894,N_16617,N_16676);
xnor U16895 (N_16895,N_16798,N_16749);
nor U16896 (N_16896,N_16752,N_16602);
xnor U16897 (N_16897,N_16758,N_16796);
and U16898 (N_16898,N_16755,N_16786);
nor U16899 (N_16899,N_16721,N_16616);
or U16900 (N_16900,N_16604,N_16795);
xnor U16901 (N_16901,N_16635,N_16638);
xor U16902 (N_16902,N_16629,N_16771);
nand U16903 (N_16903,N_16600,N_16694);
or U16904 (N_16904,N_16777,N_16636);
nor U16905 (N_16905,N_16702,N_16691);
and U16906 (N_16906,N_16719,N_16717);
or U16907 (N_16907,N_16731,N_16711);
xnor U16908 (N_16908,N_16606,N_16687);
xor U16909 (N_16909,N_16722,N_16780);
or U16910 (N_16910,N_16641,N_16739);
nand U16911 (N_16911,N_16664,N_16773);
nor U16912 (N_16912,N_16711,N_16746);
or U16913 (N_16913,N_16646,N_16704);
xnor U16914 (N_16914,N_16651,N_16727);
nor U16915 (N_16915,N_16665,N_16648);
xor U16916 (N_16916,N_16753,N_16704);
nor U16917 (N_16917,N_16744,N_16645);
or U16918 (N_16918,N_16785,N_16757);
nand U16919 (N_16919,N_16627,N_16615);
xnor U16920 (N_16920,N_16739,N_16756);
nor U16921 (N_16921,N_16789,N_16674);
nand U16922 (N_16922,N_16790,N_16668);
nand U16923 (N_16923,N_16652,N_16657);
or U16924 (N_16924,N_16670,N_16766);
nand U16925 (N_16925,N_16652,N_16787);
nand U16926 (N_16926,N_16782,N_16662);
or U16927 (N_16927,N_16797,N_16672);
and U16928 (N_16928,N_16695,N_16688);
xor U16929 (N_16929,N_16744,N_16672);
or U16930 (N_16930,N_16793,N_16743);
or U16931 (N_16931,N_16709,N_16711);
nand U16932 (N_16932,N_16661,N_16714);
or U16933 (N_16933,N_16651,N_16656);
or U16934 (N_16934,N_16745,N_16642);
nand U16935 (N_16935,N_16687,N_16754);
and U16936 (N_16936,N_16645,N_16693);
xor U16937 (N_16937,N_16788,N_16745);
nand U16938 (N_16938,N_16719,N_16731);
xnor U16939 (N_16939,N_16682,N_16602);
or U16940 (N_16940,N_16672,N_16768);
and U16941 (N_16941,N_16605,N_16650);
and U16942 (N_16942,N_16614,N_16717);
xnor U16943 (N_16943,N_16614,N_16675);
and U16944 (N_16944,N_16674,N_16776);
nor U16945 (N_16945,N_16767,N_16689);
nand U16946 (N_16946,N_16674,N_16600);
nand U16947 (N_16947,N_16640,N_16673);
xor U16948 (N_16948,N_16784,N_16613);
and U16949 (N_16949,N_16744,N_16788);
or U16950 (N_16950,N_16772,N_16681);
nor U16951 (N_16951,N_16742,N_16731);
or U16952 (N_16952,N_16661,N_16726);
and U16953 (N_16953,N_16616,N_16766);
or U16954 (N_16954,N_16631,N_16614);
xor U16955 (N_16955,N_16791,N_16650);
nand U16956 (N_16956,N_16787,N_16613);
xnor U16957 (N_16957,N_16696,N_16682);
and U16958 (N_16958,N_16783,N_16738);
and U16959 (N_16959,N_16770,N_16611);
nor U16960 (N_16960,N_16763,N_16681);
nor U16961 (N_16961,N_16615,N_16685);
and U16962 (N_16962,N_16733,N_16671);
nand U16963 (N_16963,N_16759,N_16609);
or U16964 (N_16964,N_16741,N_16730);
nor U16965 (N_16965,N_16700,N_16741);
and U16966 (N_16966,N_16754,N_16782);
or U16967 (N_16967,N_16617,N_16732);
nor U16968 (N_16968,N_16746,N_16769);
nor U16969 (N_16969,N_16766,N_16790);
xor U16970 (N_16970,N_16725,N_16673);
nor U16971 (N_16971,N_16645,N_16789);
or U16972 (N_16972,N_16742,N_16606);
xor U16973 (N_16973,N_16630,N_16684);
and U16974 (N_16974,N_16761,N_16657);
xnor U16975 (N_16975,N_16708,N_16786);
or U16976 (N_16976,N_16735,N_16764);
nand U16977 (N_16977,N_16757,N_16729);
nor U16978 (N_16978,N_16719,N_16783);
and U16979 (N_16979,N_16636,N_16628);
or U16980 (N_16980,N_16643,N_16622);
and U16981 (N_16981,N_16707,N_16736);
nor U16982 (N_16982,N_16736,N_16797);
and U16983 (N_16983,N_16686,N_16633);
or U16984 (N_16984,N_16692,N_16637);
nor U16985 (N_16985,N_16789,N_16796);
or U16986 (N_16986,N_16629,N_16677);
nand U16987 (N_16987,N_16732,N_16727);
or U16988 (N_16988,N_16745,N_16645);
nor U16989 (N_16989,N_16766,N_16682);
or U16990 (N_16990,N_16678,N_16689);
and U16991 (N_16991,N_16679,N_16684);
nand U16992 (N_16992,N_16718,N_16691);
and U16993 (N_16993,N_16702,N_16655);
or U16994 (N_16994,N_16620,N_16656);
and U16995 (N_16995,N_16796,N_16767);
and U16996 (N_16996,N_16631,N_16767);
nand U16997 (N_16997,N_16629,N_16741);
or U16998 (N_16998,N_16786,N_16653);
xor U16999 (N_16999,N_16605,N_16670);
nand U17000 (N_17000,N_16882,N_16992);
xnor U17001 (N_17001,N_16890,N_16983);
and U17002 (N_17002,N_16815,N_16952);
nor U17003 (N_17003,N_16954,N_16941);
or U17004 (N_17004,N_16912,N_16802);
and U17005 (N_17005,N_16988,N_16861);
nor U17006 (N_17006,N_16873,N_16868);
nand U17007 (N_17007,N_16995,N_16929);
nor U17008 (N_17008,N_16851,N_16808);
nor U17009 (N_17009,N_16963,N_16888);
and U17010 (N_17010,N_16825,N_16836);
nand U17011 (N_17011,N_16845,N_16958);
nor U17012 (N_17012,N_16982,N_16820);
nor U17013 (N_17013,N_16897,N_16810);
or U17014 (N_17014,N_16998,N_16921);
or U17015 (N_17015,N_16872,N_16887);
xor U17016 (N_17016,N_16800,N_16804);
and U17017 (N_17017,N_16997,N_16817);
and U17018 (N_17018,N_16844,N_16940);
nand U17019 (N_17019,N_16919,N_16839);
or U17020 (N_17020,N_16848,N_16891);
or U17021 (N_17021,N_16937,N_16809);
xnor U17022 (N_17022,N_16870,N_16824);
nor U17023 (N_17023,N_16860,N_16904);
nand U17024 (N_17024,N_16920,N_16854);
and U17025 (N_17025,N_16812,N_16986);
xor U17026 (N_17026,N_16962,N_16840);
or U17027 (N_17027,N_16886,N_16857);
nor U17028 (N_17028,N_16990,N_16842);
nor U17029 (N_17029,N_16864,N_16834);
or U17030 (N_17030,N_16970,N_16907);
nor U17031 (N_17031,N_16884,N_16811);
nor U17032 (N_17032,N_16946,N_16908);
nand U17033 (N_17033,N_16866,N_16969);
nor U17034 (N_17034,N_16947,N_16837);
nand U17035 (N_17035,N_16913,N_16955);
xor U17036 (N_17036,N_16885,N_16926);
nor U17037 (N_17037,N_16938,N_16867);
nand U17038 (N_17038,N_16829,N_16917);
and U17039 (N_17039,N_16862,N_16974);
or U17040 (N_17040,N_16999,N_16852);
xor U17041 (N_17041,N_16827,N_16855);
or U17042 (N_17042,N_16977,N_16996);
and U17043 (N_17043,N_16879,N_16994);
xnor U17044 (N_17044,N_16874,N_16951);
xnor U17045 (N_17045,N_16973,N_16838);
nor U17046 (N_17046,N_16821,N_16899);
and U17047 (N_17047,N_16935,N_16987);
xor U17048 (N_17048,N_16918,N_16914);
nor U17049 (N_17049,N_16819,N_16949);
and U17050 (N_17050,N_16957,N_16883);
and U17051 (N_17051,N_16944,N_16847);
and U17052 (N_17052,N_16806,N_16959);
nand U17053 (N_17053,N_16985,N_16902);
and U17054 (N_17054,N_16801,N_16905);
nand U17055 (N_17055,N_16901,N_16953);
nand U17056 (N_17056,N_16943,N_16823);
and U17057 (N_17057,N_16871,N_16822);
xnor U17058 (N_17058,N_16828,N_16903);
nor U17059 (N_17059,N_16859,N_16939);
or U17060 (N_17060,N_16960,N_16975);
and U17061 (N_17061,N_16816,N_16928);
and U17062 (N_17062,N_16826,N_16923);
nor U17063 (N_17063,N_16813,N_16964);
nor U17064 (N_17064,N_16876,N_16832);
nor U17065 (N_17065,N_16835,N_16863);
nor U17066 (N_17066,N_16916,N_16865);
nor U17067 (N_17067,N_16878,N_16898);
and U17068 (N_17068,N_16980,N_16906);
nand U17069 (N_17069,N_16981,N_16893);
or U17070 (N_17070,N_16894,N_16895);
nor U17071 (N_17071,N_16841,N_16877);
nand U17072 (N_17072,N_16948,N_16850);
nor U17073 (N_17073,N_16933,N_16979);
or U17074 (N_17074,N_16831,N_16853);
or U17075 (N_17075,N_16910,N_16966);
nor U17076 (N_17076,N_16930,N_16950);
or U17077 (N_17077,N_16991,N_16961);
and U17078 (N_17078,N_16896,N_16932);
nor U17079 (N_17079,N_16849,N_16978);
or U17080 (N_17080,N_16843,N_16971);
xnor U17081 (N_17081,N_16846,N_16909);
xor U17082 (N_17082,N_16911,N_16984);
nand U17083 (N_17083,N_16875,N_16881);
nand U17084 (N_17084,N_16880,N_16972);
nor U17085 (N_17085,N_16869,N_16900);
nand U17086 (N_17086,N_16889,N_16931);
and U17087 (N_17087,N_16915,N_16967);
and U17088 (N_17088,N_16830,N_16993);
and U17089 (N_17089,N_16833,N_16856);
nand U17090 (N_17090,N_16922,N_16945);
and U17091 (N_17091,N_16818,N_16942);
xor U17092 (N_17092,N_16989,N_16968);
nor U17093 (N_17093,N_16924,N_16965);
or U17094 (N_17094,N_16927,N_16807);
or U17095 (N_17095,N_16858,N_16892);
nor U17096 (N_17096,N_16936,N_16925);
or U17097 (N_17097,N_16805,N_16934);
xnor U17098 (N_17098,N_16803,N_16814);
nand U17099 (N_17099,N_16976,N_16956);
and U17100 (N_17100,N_16961,N_16981);
and U17101 (N_17101,N_16816,N_16983);
nor U17102 (N_17102,N_16982,N_16898);
nand U17103 (N_17103,N_16894,N_16962);
and U17104 (N_17104,N_16876,N_16903);
nor U17105 (N_17105,N_16959,N_16820);
nand U17106 (N_17106,N_16900,N_16955);
nor U17107 (N_17107,N_16814,N_16996);
nor U17108 (N_17108,N_16903,N_16823);
or U17109 (N_17109,N_16838,N_16831);
nand U17110 (N_17110,N_16818,N_16931);
nand U17111 (N_17111,N_16887,N_16861);
or U17112 (N_17112,N_16824,N_16878);
nand U17113 (N_17113,N_16940,N_16908);
and U17114 (N_17114,N_16885,N_16924);
xnor U17115 (N_17115,N_16947,N_16972);
and U17116 (N_17116,N_16935,N_16905);
nor U17117 (N_17117,N_16986,N_16957);
nor U17118 (N_17118,N_16827,N_16992);
and U17119 (N_17119,N_16911,N_16851);
nor U17120 (N_17120,N_16943,N_16913);
xor U17121 (N_17121,N_16837,N_16817);
and U17122 (N_17122,N_16963,N_16920);
and U17123 (N_17123,N_16878,N_16980);
nor U17124 (N_17124,N_16847,N_16878);
nand U17125 (N_17125,N_16909,N_16901);
or U17126 (N_17126,N_16869,N_16951);
or U17127 (N_17127,N_16815,N_16964);
nor U17128 (N_17128,N_16836,N_16823);
or U17129 (N_17129,N_16837,N_16982);
nand U17130 (N_17130,N_16994,N_16988);
and U17131 (N_17131,N_16912,N_16997);
xor U17132 (N_17132,N_16816,N_16847);
nand U17133 (N_17133,N_16920,N_16979);
or U17134 (N_17134,N_16975,N_16983);
nand U17135 (N_17135,N_16915,N_16827);
xnor U17136 (N_17136,N_16843,N_16949);
nand U17137 (N_17137,N_16839,N_16801);
or U17138 (N_17138,N_16920,N_16928);
nand U17139 (N_17139,N_16992,N_16926);
and U17140 (N_17140,N_16967,N_16884);
xnor U17141 (N_17141,N_16800,N_16916);
nor U17142 (N_17142,N_16970,N_16948);
xor U17143 (N_17143,N_16995,N_16896);
or U17144 (N_17144,N_16844,N_16887);
nor U17145 (N_17145,N_16963,N_16853);
xnor U17146 (N_17146,N_16863,N_16814);
and U17147 (N_17147,N_16906,N_16879);
nand U17148 (N_17148,N_16921,N_16986);
xnor U17149 (N_17149,N_16892,N_16873);
nor U17150 (N_17150,N_16907,N_16897);
or U17151 (N_17151,N_16904,N_16982);
xor U17152 (N_17152,N_16856,N_16994);
or U17153 (N_17153,N_16991,N_16965);
and U17154 (N_17154,N_16986,N_16815);
xor U17155 (N_17155,N_16801,N_16900);
nor U17156 (N_17156,N_16854,N_16886);
nor U17157 (N_17157,N_16823,N_16806);
xnor U17158 (N_17158,N_16946,N_16884);
and U17159 (N_17159,N_16863,N_16891);
nor U17160 (N_17160,N_16927,N_16973);
nand U17161 (N_17161,N_16834,N_16942);
nor U17162 (N_17162,N_16936,N_16935);
xnor U17163 (N_17163,N_16858,N_16803);
or U17164 (N_17164,N_16815,N_16910);
or U17165 (N_17165,N_16800,N_16895);
xor U17166 (N_17166,N_16896,N_16912);
nor U17167 (N_17167,N_16808,N_16884);
nor U17168 (N_17168,N_16926,N_16925);
xor U17169 (N_17169,N_16985,N_16868);
and U17170 (N_17170,N_16879,N_16958);
xor U17171 (N_17171,N_16946,N_16990);
nand U17172 (N_17172,N_16803,N_16827);
nor U17173 (N_17173,N_16861,N_16853);
nand U17174 (N_17174,N_16838,N_16837);
nor U17175 (N_17175,N_16819,N_16920);
and U17176 (N_17176,N_16946,N_16850);
xor U17177 (N_17177,N_16943,N_16932);
and U17178 (N_17178,N_16804,N_16991);
nor U17179 (N_17179,N_16941,N_16935);
nand U17180 (N_17180,N_16996,N_16835);
or U17181 (N_17181,N_16899,N_16981);
xor U17182 (N_17182,N_16947,N_16941);
nand U17183 (N_17183,N_16960,N_16997);
xor U17184 (N_17184,N_16894,N_16969);
nand U17185 (N_17185,N_16876,N_16829);
and U17186 (N_17186,N_16912,N_16842);
nand U17187 (N_17187,N_16862,N_16934);
or U17188 (N_17188,N_16876,N_16972);
nor U17189 (N_17189,N_16890,N_16882);
xor U17190 (N_17190,N_16916,N_16972);
nand U17191 (N_17191,N_16908,N_16835);
and U17192 (N_17192,N_16961,N_16959);
or U17193 (N_17193,N_16866,N_16889);
xnor U17194 (N_17194,N_16871,N_16963);
nand U17195 (N_17195,N_16812,N_16898);
or U17196 (N_17196,N_16880,N_16870);
or U17197 (N_17197,N_16861,N_16978);
or U17198 (N_17198,N_16943,N_16936);
xnor U17199 (N_17199,N_16803,N_16967);
nand U17200 (N_17200,N_17105,N_17049);
nand U17201 (N_17201,N_17056,N_17077);
or U17202 (N_17202,N_17021,N_17175);
and U17203 (N_17203,N_17194,N_17071);
or U17204 (N_17204,N_17166,N_17060);
or U17205 (N_17205,N_17075,N_17184);
or U17206 (N_17206,N_17182,N_17180);
nand U17207 (N_17207,N_17000,N_17150);
or U17208 (N_17208,N_17098,N_17007);
or U17209 (N_17209,N_17011,N_17028);
and U17210 (N_17210,N_17043,N_17005);
and U17211 (N_17211,N_17193,N_17037);
xor U17212 (N_17212,N_17044,N_17106);
or U17213 (N_17213,N_17025,N_17055);
and U17214 (N_17214,N_17032,N_17008);
nor U17215 (N_17215,N_17086,N_17093);
nand U17216 (N_17216,N_17185,N_17165);
nand U17217 (N_17217,N_17127,N_17046);
and U17218 (N_17218,N_17178,N_17143);
nor U17219 (N_17219,N_17083,N_17097);
xor U17220 (N_17220,N_17048,N_17145);
or U17221 (N_17221,N_17036,N_17066);
nor U17222 (N_17222,N_17023,N_17009);
and U17223 (N_17223,N_17058,N_17074);
xor U17224 (N_17224,N_17198,N_17112);
nor U17225 (N_17225,N_17116,N_17039);
and U17226 (N_17226,N_17161,N_17001);
xnor U17227 (N_17227,N_17045,N_17092);
or U17228 (N_17228,N_17033,N_17133);
nand U17229 (N_17229,N_17014,N_17119);
or U17230 (N_17230,N_17131,N_17156);
xnor U17231 (N_17231,N_17004,N_17068);
nand U17232 (N_17232,N_17136,N_17129);
xor U17233 (N_17233,N_17163,N_17029);
and U17234 (N_17234,N_17095,N_17019);
or U17235 (N_17235,N_17190,N_17196);
and U17236 (N_17236,N_17110,N_17167);
or U17237 (N_17237,N_17067,N_17155);
or U17238 (N_17238,N_17016,N_17189);
nor U17239 (N_17239,N_17139,N_17038);
or U17240 (N_17240,N_17148,N_17051);
and U17241 (N_17241,N_17057,N_17158);
nand U17242 (N_17242,N_17177,N_17192);
nor U17243 (N_17243,N_17085,N_17128);
nor U17244 (N_17244,N_17146,N_17030);
nor U17245 (N_17245,N_17114,N_17174);
xnor U17246 (N_17246,N_17191,N_17135);
or U17247 (N_17247,N_17024,N_17186);
nor U17248 (N_17248,N_17078,N_17176);
nor U17249 (N_17249,N_17102,N_17173);
and U17250 (N_17250,N_17117,N_17113);
xor U17251 (N_17251,N_17153,N_17187);
and U17252 (N_17252,N_17100,N_17142);
or U17253 (N_17253,N_17080,N_17070);
and U17254 (N_17254,N_17052,N_17159);
xnor U17255 (N_17255,N_17027,N_17094);
and U17256 (N_17256,N_17041,N_17199);
nand U17257 (N_17257,N_17138,N_17101);
or U17258 (N_17258,N_17054,N_17061);
nand U17259 (N_17259,N_17144,N_17026);
or U17260 (N_17260,N_17157,N_17050);
nor U17261 (N_17261,N_17072,N_17076);
nand U17262 (N_17262,N_17126,N_17169);
and U17263 (N_17263,N_17034,N_17132);
and U17264 (N_17264,N_17195,N_17087);
or U17265 (N_17265,N_17121,N_17059);
nand U17266 (N_17266,N_17109,N_17134);
nand U17267 (N_17267,N_17149,N_17063);
nor U17268 (N_17268,N_17152,N_17179);
xnor U17269 (N_17269,N_17082,N_17012);
xnor U17270 (N_17270,N_17120,N_17140);
nand U17271 (N_17271,N_17010,N_17035);
or U17272 (N_17272,N_17002,N_17081);
and U17273 (N_17273,N_17141,N_17160);
nand U17274 (N_17274,N_17111,N_17123);
and U17275 (N_17275,N_17084,N_17088);
xnor U17276 (N_17276,N_17069,N_17107);
nor U17277 (N_17277,N_17183,N_17164);
nor U17278 (N_17278,N_17188,N_17096);
and U17279 (N_17279,N_17013,N_17047);
nand U17280 (N_17280,N_17003,N_17162);
nor U17281 (N_17281,N_17118,N_17031);
or U17282 (N_17282,N_17079,N_17089);
or U17283 (N_17283,N_17073,N_17064);
nand U17284 (N_17284,N_17099,N_17020);
nand U17285 (N_17285,N_17130,N_17015);
xnor U17286 (N_17286,N_17154,N_17197);
nor U17287 (N_17287,N_17042,N_17151);
nand U17288 (N_17288,N_17022,N_17170);
or U17289 (N_17289,N_17104,N_17115);
and U17290 (N_17290,N_17006,N_17122);
or U17291 (N_17291,N_17103,N_17018);
nor U17292 (N_17292,N_17172,N_17062);
xor U17293 (N_17293,N_17124,N_17168);
xor U17294 (N_17294,N_17147,N_17125);
and U17295 (N_17295,N_17181,N_17090);
xnor U17296 (N_17296,N_17040,N_17137);
nand U17297 (N_17297,N_17171,N_17017);
nand U17298 (N_17298,N_17065,N_17091);
and U17299 (N_17299,N_17053,N_17108);
and U17300 (N_17300,N_17144,N_17121);
and U17301 (N_17301,N_17035,N_17084);
and U17302 (N_17302,N_17009,N_17195);
and U17303 (N_17303,N_17025,N_17122);
nand U17304 (N_17304,N_17129,N_17100);
or U17305 (N_17305,N_17138,N_17018);
nand U17306 (N_17306,N_17102,N_17184);
or U17307 (N_17307,N_17059,N_17193);
nand U17308 (N_17308,N_17057,N_17094);
xnor U17309 (N_17309,N_17179,N_17018);
xnor U17310 (N_17310,N_17036,N_17027);
nor U17311 (N_17311,N_17007,N_17137);
and U17312 (N_17312,N_17097,N_17164);
nand U17313 (N_17313,N_17020,N_17167);
nor U17314 (N_17314,N_17155,N_17109);
and U17315 (N_17315,N_17158,N_17088);
or U17316 (N_17316,N_17162,N_17085);
xor U17317 (N_17317,N_17038,N_17067);
xnor U17318 (N_17318,N_17049,N_17111);
or U17319 (N_17319,N_17182,N_17092);
nand U17320 (N_17320,N_17003,N_17045);
and U17321 (N_17321,N_17090,N_17113);
or U17322 (N_17322,N_17030,N_17025);
or U17323 (N_17323,N_17125,N_17016);
or U17324 (N_17324,N_17192,N_17029);
and U17325 (N_17325,N_17002,N_17109);
and U17326 (N_17326,N_17182,N_17140);
and U17327 (N_17327,N_17097,N_17023);
and U17328 (N_17328,N_17003,N_17181);
nand U17329 (N_17329,N_17166,N_17130);
and U17330 (N_17330,N_17082,N_17145);
or U17331 (N_17331,N_17087,N_17033);
and U17332 (N_17332,N_17057,N_17153);
nor U17333 (N_17333,N_17033,N_17136);
and U17334 (N_17334,N_17196,N_17182);
nor U17335 (N_17335,N_17159,N_17019);
nand U17336 (N_17336,N_17113,N_17088);
xnor U17337 (N_17337,N_17194,N_17072);
and U17338 (N_17338,N_17167,N_17143);
nor U17339 (N_17339,N_17162,N_17053);
and U17340 (N_17340,N_17022,N_17043);
and U17341 (N_17341,N_17059,N_17060);
xor U17342 (N_17342,N_17089,N_17141);
or U17343 (N_17343,N_17182,N_17152);
and U17344 (N_17344,N_17006,N_17153);
and U17345 (N_17345,N_17162,N_17176);
nand U17346 (N_17346,N_17187,N_17099);
nand U17347 (N_17347,N_17178,N_17050);
or U17348 (N_17348,N_17115,N_17070);
xor U17349 (N_17349,N_17097,N_17114);
xnor U17350 (N_17350,N_17173,N_17088);
nor U17351 (N_17351,N_17160,N_17154);
nand U17352 (N_17352,N_17075,N_17048);
and U17353 (N_17353,N_17140,N_17164);
nor U17354 (N_17354,N_17081,N_17055);
nor U17355 (N_17355,N_17164,N_17075);
or U17356 (N_17356,N_17148,N_17120);
or U17357 (N_17357,N_17066,N_17163);
nor U17358 (N_17358,N_17166,N_17161);
nand U17359 (N_17359,N_17141,N_17192);
xor U17360 (N_17360,N_17190,N_17169);
or U17361 (N_17361,N_17023,N_17055);
nor U17362 (N_17362,N_17037,N_17005);
xnor U17363 (N_17363,N_17155,N_17068);
and U17364 (N_17364,N_17116,N_17087);
or U17365 (N_17365,N_17096,N_17179);
nand U17366 (N_17366,N_17106,N_17017);
nand U17367 (N_17367,N_17087,N_17076);
and U17368 (N_17368,N_17096,N_17037);
xnor U17369 (N_17369,N_17166,N_17198);
nand U17370 (N_17370,N_17039,N_17148);
xor U17371 (N_17371,N_17133,N_17142);
nand U17372 (N_17372,N_17001,N_17040);
and U17373 (N_17373,N_17087,N_17050);
and U17374 (N_17374,N_17160,N_17000);
xor U17375 (N_17375,N_17003,N_17173);
or U17376 (N_17376,N_17010,N_17129);
xnor U17377 (N_17377,N_17039,N_17008);
and U17378 (N_17378,N_17081,N_17198);
or U17379 (N_17379,N_17178,N_17117);
and U17380 (N_17380,N_17022,N_17081);
nand U17381 (N_17381,N_17108,N_17118);
nor U17382 (N_17382,N_17192,N_17108);
or U17383 (N_17383,N_17088,N_17002);
nand U17384 (N_17384,N_17115,N_17079);
xnor U17385 (N_17385,N_17136,N_17088);
nand U17386 (N_17386,N_17089,N_17025);
xnor U17387 (N_17387,N_17019,N_17188);
nor U17388 (N_17388,N_17042,N_17028);
nor U17389 (N_17389,N_17086,N_17198);
nand U17390 (N_17390,N_17101,N_17167);
nand U17391 (N_17391,N_17089,N_17162);
xor U17392 (N_17392,N_17056,N_17102);
nand U17393 (N_17393,N_17100,N_17056);
or U17394 (N_17394,N_17147,N_17167);
or U17395 (N_17395,N_17157,N_17161);
nand U17396 (N_17396,N_17050,N_17017);
nor U17397 (N_17397,N_17002,N_17196);
and U17398 (N_17398,N_17129,N_17152);
nand U17399 (N_17399,N_17031,N_17052);
and U17400 (N_17400,N_17392,N_17290);
nand U17401 (N_17401,N_17246,N_17225);
or U17402 (N_17402,N_17339,N_17322);
xor U17403 (N_17403,N_17226,N_17342);
and U17404 (N_17404,N_17311,N_17385);
or U17405 (N_17405,N_17352,N_17395);
xor U17406 (N_17406,N_17229,N_17285);
and U17407 (N_17407,N_17337,N_17308);
nor U17408 (N_17408,N_17353,N_17393);
nor U17409 (N_17409,N_17218,N_17275);
and U17410 (N_17410,N_17286,N_17384);
and U17411 (N_17411,N_17272,N_17224);
xnor U17412 (N_17412,N_17382,N_17294);
xor U17413 (N_17413,N_17377,N_17253);
nor U17414 (N_17414,N_17365,N_17251);
nor U17415 (N_17415,N_17212,N_17310);
nor U17416 (N_17416,N_17364,N_17330);
nand U17417 (N_17417,N_17305,N_17361);
and U17418 (N_17418,N_17367,N_17256);
nand U17419 (N_17419,N_17394,N_17213);
and U17420 (N_17420,N_17380,N_17201);
or U17421 (N_17421,N_17296,N_17379);
and U17422 (N_17422,N_17355,N_17237);
nor U17423 (N_17423,N_17345,N_17205);
xnor U17424 (N_17424,N_17265,N_17210);
nand U17425 (N_17425,N_17328,N_17239);
or U17426 (N_17426,N_17344,N_17232);
or U17427 (N_17427,N_17297,N_17207);
nor U17428 (N_17428,N_17397,N_17359);
nand U17429 (N_17429,N_17317,N_17289);
and U17430 (N_17430,N_17291,N_17278);
and U17431 (N_17431,N_17329,N_17302);
nand U17432 (N_17432,N_17321,N_17331);
nand U17433 (N_17433,N_17356,N_17368);
or U17434 (N_17434,N_17222,N_17348);
or U17435 (N_17435,N_17233,N_17371);
xor U17436 (N_17436,N_17252,N_17343);
and U17437 (N_17437,N_17214,N_17396);
xnor U17438 (N_17438,N_17314,N_17333);
xnor U17439 (N_17439,N_17363,N_17281);
nor U17440 (N_17440,N_17261,N_17273);
nor U17441 (N_17441,N_17318,N_17350);
and U17442 (N_17442,N_17200,N_17269);
and U17443 (N_17443,N_17284,N_17389);
nor U17444 (N_17444,N_17346,N_17262);
nor U17445 (N_17445,N_17301,N_17254);
xnor U17446 (N_17446,N_17245,N_17357);
or U17447 (N_17447,N_17387,N_17386);
xor U17448 (N_17448,N_17336,N_17341);
or U17449 (N_17449,N_17373,N_17258);
and U17450 (N_17450,N_17306,N_17366);
nand U17451 (N_17451,N_17255,N_17316);
or U17452 (N_17452,N_17347,N_17349);
xnor U17453 (N_17453,N_17282,N_17227);
nor U17454 (N_17454,N_17216,N_17325);
xor U17455 (N_17455,N_17388,N_17223);
xnor U17456 (N_17456,N_17264,N_17231);
nand U17457 (N_17457,N_17240,N_17219);
or U17458 (N_17458,N_17326,N_17370);
or U17459 (N_17459,N_17378,N_17241);
nand U17460 (N_17460,N_17259,N_17271);
nor U17461 (N_17461,N_17236,N_17335);
or U17462 (N_17462,N_17244,N_17369);
xor U17463 (N_17463,N_17228,N_17250);
nor U17464 (N_17464,N_17288,N_17332);
xnor U17465 (N_17465,N_17257,N_17360);
and U17466 (N_17466,N_17372,N_17238);
or U17467 (N_17467,N_17203,N_17381);
nor U17468 (N_17468,N_17260,N_17274);
and U17469 (N_17469,N_17234,N_17270);
xnor U17470 (N_17470,N_17221,N_17217);
xor U17471 (N_17471,N_17351,N_17279);
nor U17472 (N_17472,N_17398,N_17293);
or U17473 (N_17473,N_17263,N_17266);
nor U17474 (N_17474,N_17242,N_17340);
xor U17475 (N_17475,N_17206,N_17390);
xnor U17476 (N_17476,N_17299,N_17334);
xnor U17477 (N_17477,N_17208,N_17376);
or U17478 (N_17478,N_17309,N_17277);
nor U17479 (N_17479,N_17374,N_17383);
xnor U17480 (N_17480,N_17209,N_17338);
nor U17481 (N_17481,N_17313,N_17320);
and U17482 (N_17482,N_17375,N_17287);
xor U17483 (N_17483,N_17323,N_17399);
or U17484 (N_17484,N_17354,N_17319);
or U17485 (N_17485,N_17280,N_17202);
xor U17486 (N_17486,N_17327,N_17324);
xor U17487 (N_17487,N_17358,N_17243);
xor U17488 (N_17488,N_17283,N_17211);
nor U17489 (N_17489,N_17204,N_17230);
xnor U17490 (N_17490,N_17304,N_17215);
xor U17491 (N_17491,N_17220,N_17295);
nor U17492 (N_17492,N_17276,N_17249);
xnor U17493 (N_17493,N_17303,N_17307);
nand U17494 (N_17494,N_17235,N_17362);
xnor U17495 (N_17495,N_17300,N_17267);
and U17496 (N_17496,N_17247,N_17298);
nor U17497 (N_17497,N_17391,N_17312);
nand U17498 (N_17498,N_17315,N_17268);
or U17499 (N_17499,N_17292,N_17248);
or U17500 (N_17500,N_17214,N_17354);
or U17501 (N_17501,N_17327,N_17284);
and U17502 (N_17502,N_17314,N_17202);
or U17503 (N_17503,N_17363,N_17262);
xor U17504 (N_17504,N_17254,N_17344);
and U17505 (N_17505,N_17313,N_17373);
xor U17506 (N_17506,N_17251,N_17390);
and U17507 (N_17507,N_17205,N_17312);
xor U17508 (N_17508,N_17352,N_17295);
xor U17509 (N_17509,N_17297,N_17301);
nand U17510 (N_17510,N_17341,N_17253);
xnor U17511 (N_17511,N_17346,N_17277);
or U17512 (N_17512,N_17372,N_17257);
nand U17513 (N_17513,N_17297,N_17361);
nand U17514 (N_17514,N_17204,N_17245);
xor U17515 (N_17515,N_17383,N_17365);
and U17516 (N_17516,N_17212,N_17230);
and U17517 (N_17517,N_17297,N_17247);
and U17518 (N_17518,N_17222,N_17249);
nand U17519 (N_17519,N_17259,N_17326);
nand U17520 (N_17520,N_17344,N_17293);
nor U17521 (N_17521,N_17215,N_17218);
or U17522 (N_17522,N_17258,N_17243);
or U17523 (N_17523,N_17271,N_17230);
or U17524 (N_17524,N_17299,N_17261);
nand U17525 (N_17525,N_17238,N_17331);
xor U17526 (N_17526,N_17209,N_17273);
or U17527 (N_17527,N_17214,N_17276);
nor U17528 (N_17528,N_17384,N_17353);
nor U17529 (N_17529,N_17334,N_17344);
and U17530 (N_17530,N_17350,N_17295);
nand U17531 (N_17531,N_17274,N_17234);
nand U17532 (N_17532,N_17360,N_17256);
and U17533 (N_17533,N_17286,N_17383);
and U17534 (N_17534,N_17358,N_17357);
or U17535 (N_17535,N_17336,N_17205);
nand U17536 (N_17536,N_17321,N_17274);
nor U17537 (N_17537,N_17273,N_17298);
nor U17538 (N_17538,N_17293,N_17269);
xnor U17539 (N_17539,N_17242,N_17350);
nor U17540 (N_17540,N_17343,N_17270);
xnor U17541 (N_17541,N_17256,N_17217);
xnor U17542 (N_17542,N_17225,N_17281);
nor U17543 (N_17543,N_17293,N_17250);
or U17544 (N_17544,N_17395,N_17245);
xnor U17545 (N_17545,N_17321,N_17300);
and U17546 (N_17546,N_17332,N_17310);
or U17547 (N_17547,N_17263,N_17282);
nand U17548 (N_17548,N_17391,N_17303);
nor U17549 (N_17549,N_17281,N_17371);
or U17550 (N_17550,N_17213,N_17252);
nor U17551 (N_17551,N_17334,N_17250);
xor U17552 (N_17552,N_17267,N_17355);
and U17553 (N_17553,N_17368,N_17310);
and U17554 (N_17554,N_17351,N_17364);
and U17555 (N_17555,N_17311,N_17227);
and U17556 (N_17556,N_17376,N_17263);
and U17557 (N_17557,N_17252,N_17203);
nor U17558 (N_17558,N_17391,N_17343);
or U17559 (N_17559,N_17351,N_17370);
xnor U17560 (N_17560,N_17220,N_17302);
xor U17561 (N_17561,N_17233,N_17207);
xor U17562 (N_17562,N_17210,N_17268);
nor U17563 (N_17563,N_17207,N_17222);
and U17564 (N_17564,N_17223,N_17245);
nor U17565 (N_17565,N_17339,N_17208);
xor U17566 (N_17566,N_17252,N_17392);
nand U17567 (N_17567,N_17212,N_17229);
nand U17568 (N_17568,N_17245,N_17279);
nand U17569 (N_17569,N_17382,N_17309);
xnor U17570 (N_17570,N_17202,N_17228);
nor U17571 (N_17571,N_17251,N_17258);
xor U17572 (N_17572,N_17324,N_17315);
nand U17573 (N_17573,N_17260,N_17201);
and U17574 (N_17574,N_17274,N_17305);
or U17575 (N_17575,N_17204,N_17399);
and U17576 (N_17576,N_17338,N_17294);
nor U17577 (N_17577,N_17252,N_17310);
or U17578 (N_17578,N_17276,N_17257);
nand U17579 (N_17579,N_17385,N_17229);
xor U17580 (N_17580,N_17214,N_17372);
or U17581 (N_17581,N_17253,N_17217);
nor U17582 (N_17582,N_17307,N_17395);
xor U17583 (N_17583,N_17210,N_17385);
nor U17584 (N_17584,N_17298,N_17219);
nand U17585 (N_17585,N_17319,N_17279);
nand U17586 (N_17586,N_17220,N_17351);
and U17587 (N_17587,N_17335,N_17392);
nor U17588 (N_17588,N_17276,N_17305);
xor U17589 (N_17589,N_17350,N_17247);
xor U17590 (N_17590,N_17374,N_17223);
or U17591 (N_17591,N_17377,N_17371);
nand U17592 (N_17592,N_17287,N_17290);
and U17593 (N_17593,N_17204,N_17228);
nand U17594 (N_17594,N_17216,N_17276);
xnor U17595 (N_17595,N_17347,N_17368);
and U17596 (N_17596,N_17270,N_17221);
nor U17597 (N_17597,N_17298,N_17313);
nand U17598 (N_17598,N_17301,N_17353);
xor U17599 (N_17599,N_17361,N_17301);
or U17600 (N_17600,N_17558,N_17489);
and U17601 (N_17601,N_17465,N_17525);
nor U17602 (N_17602,N_17451,N_17504);
nand U17603 (N_17603,N_17548,N_17474);
xor U17604 (N_17604,N_17418,N_17562);
nor U17605 (N_17605,N_17446,N_17580);
xnor U17606 (N_17606,N_17579,N_17539);
and U17607 (N_17607,N_17431,N_17593);
nor U17608 (N_17608,N_17437,N_17488);
or U17609 (N_17609,N_17426,N_17427);
and U17610 (N_17610,N_17551,N_17450);
xor U17611 (N_17611,N_17498,N_17572);
or U17612 (N_17612,N_17567,N_17541);
nand U17613 (N_17613,N_17479,N_17573);
and U17614 (N_17614,N_17569,N_17520);
xor U17615 (N_17615,N_17590,N_17429);
nor U17616 (N_17616,N_17524,N_17534);
nor U17617 (N_17617,N_17405,N_17537);
and U17618 (N_17618,N_17597,N_17556);
or U17619 (N_17619,N_17436,N_17453);
xor U17620 (N_17620,N_17463,N_17420);
xor U17621 (N_17621,N_17528,N_17583);
and U17622 (N_17622,N_17598,N_17557);
or U17623 (N_17623,N_17447,N_17467);
xor U17624 (N_17624,N_17545,N_17501);
or U17625 (N_17625,N_17464,N_17403);
xor U17626 (N_17626,N_17515,N_17512);
or U17627 (N_17627,N_17589,N_17425);
xnor U17628 (N_17628,N_17540,N_17423);
nor U17629 (N_17629,N_17497,N_17484);
nand U17630 (N_17630,N_17435,N_17544);
xor U17631 (N_17631,N_17496,N_17588);
xnor U17632 (N_17632,N_17517,N_17411);
xor U17633 (N_17633,N_17454,N_17599);
and U17634 (N_17634,N_17442,N_17543);
xnor U17635 (N_17635,N_17581,N_17523);
xnor U17636 (N_17636,N_17417,N_17552);
or U17637 (N_17637,N_17519,N_17459);
and U17638 (N_17638,N_17486,N_17438);
nand U17639 (N_17639,N_17526,N_17502);
nor U17640 (N_17640,N_17550,N_17482);
and U17641 (N_17641,N_17565,N_17594);
and U17642 (N_17642,N_17509,N_17576);
nand U17643 (N_17643,N_17587,N_17505);
nor U17644 (N_17644,N_17582,N_17596);
and U17645 (N_17645,N_17412,N_17472);
or U17646 (N_17646,N_17428,N_17577);
or U17647 (N_17647,N_17564,N_17578);
nand U17648 (N_17648,N_17542,N_17460);
or U17649 (N_17649,N_17493,N_17470);
nand U17650 (N_17650,N_17455,N_17414);
nand U17651 (N_17651,N_17592,N_17401);
nand U17652 (N_17652,N_17494,N_17574);
xor U17653 (N_17653,N_17595,N_17457);
nor U17654 (N_17654,N_17575,N_17555);
xnor U17655 (N_17655,N_17406,N_17499);
nor U17656 (N_17656,N_17510,N_17409);
nor U17657 (N_17657,N_17476,N_17424);
nor U17658 (N_17658,N_17402,N_17585);
xnor U17659 (N_17659,N_17518,N_17553);
and U17660 (N_17660,N_17566,N_17570);
nand U17661 (N_17661,N_17527,N_17468);
xor U17662 (N_17662,N_17508,N_17485);
xnor U17663 (N_17663,N_17586,N_17487);
xnor U17664 (N_17664,N_17433,N_17445);
and U17665 (N_17665,N_17507,N_17419);
nor U17666 (N_17666,N_17416,N_17462);
xnor U17667 (N_17667,N_17404,N_17471);
and U17668 (N_17668,N_17535,N_17531);
nand U17669 (N_17669,N_17421,N_17461);
nor U17670 (N_17670,N_17521,N_17422);
or U17671 (N_17671,N_17452,N_17439);
or U17672 (N_17672,N_17483,N_17491);
nor U17673 (N_17673,N_17495,N_17481);
or U17674 (N_17674,N_17443,N_17530);
and U17675 (N_17675,N_17408,N_17532);
and U17676 (N_17676,N_17440,N_17563);
and U17677 (N_17677,N_17529,N_17473);
xor U17678 (N_17678,N_17536,N_17475);
nand U17679 (N_17679,N_17514,N_17533);
xnor U17680 (N_17680,N_17503,N_17466);
xor U17681 (N_17681,N_17559,N_17434);
nand U17682 (N_17682,N_17591,N_17546);
nand U17683 (N_17683,N_17477,N_17522);
or U17684 (N_17684,N_17432,N_17407);
and U17685 (N_17685,N_17584,N_17400);
or U17686 (N_17686,N_17415,N_17478);
nand U17687 (N_17687,N_17410,N_17441);
nor U17688 (N_17688,N_17480,N_17513);
nor U17689 (N_17689,N_17561,N_17547);
nor U17690 (N_17690,N_17456,N_17560);
xnor U17691 (N_17691,N_17492,N_17449);
xor U17692 (N_17692,N_17506,N_17444);
xor U17693 (N_17693,N_17511,N_17516);
nor U17694 (N_17694,N_17458,N_17549);
xnor U17695 (N_17695,N_17500,N_17448);
nor U17696 (N_17696,N_17568,N_17554);
or U17697 (N_17697,N_17430,N_17538);
nor U17698 (N_17698,N_17413,N_17490);
and U17699 (N_17699,N_17571,N_17469);
nor U17700 (N_17700,N_17403,N_17415);
xor U17701 (N_17701,N_17511,N_17555);
and U17702 (N_17702,N_17418,N_17411);
xor U17703 (N_17703,N_17581,N_17592);
xnor U17704 (N_17704,N_17529,N_17570);
nor U17705 (N_17705,N_17447,N_17574);
xnor U17706 (N_17706,N_17524,N_17432);
and U17707 (N_17707,N_17576,N_17471);
or U17708 (N_17708,N_17533,N_17471);
xnor U17709 (N_17709,N_17582,N_17412);
or U17710 (N_17710,N_17467,N_17586);
and U17711 (N_17711,N_17541,N_17488);
xnor U17712 (N_17712,N_17460,N_17582);
nor U17713 (N_17713,N_17470,N_17426);
or U17714 (N_17714,N_17511,N_17466);
or U17715 (N_17715,N_17582,N_17529);
or U17716 (N_17716,N_17596,N_17509);
or U17717 (N_17717,N_17451,N_17491);
or U17718 (N_17718,N_17425,N_17470);
nand U17719 (N_17719,N_17487,N_17552);
nand U17720 (N_17720,N_17533,N_17579);
or U17721 (N_17721,N_17536,N_17578);
nor U17722 (N_17722,N_17538,N_17435);
and U17723 (N_17723,N_17449,N_17518);
nor U17724 (N_17724,N_17453,N_17446);
nor U17725 (N_17725,N_17581,N_17521);
nand U17726 (N_17726,N_17594,N_17532);
nor U17727 (N_17727,N_17514,N_17459);
or U17728 (N_17728,N_17542,N_17421);
and U17729 (N_17729,N_17552,N_17580);
and U17730 (N_17730,N_17538,N_17464);
nor U17731 (N_17731,N_17553,N_17590);
and U17732 (N_17732,N_17518,N_17420);
xor U17733 (N_17733,N_17476,N_17516);
xnor U17734 (N_17734,N_17508,N_17554);
or U17735 (N_17735,N_17444,N_17504);
and U17736 (N_17736,N_17456,N_17545);
nand U17737 (N_17737,N_17548,N_17589);
or U17738 (N_17738,N_17470,N_17574);
xor U17739 (N_17739,N_17533,N_17406);
nor U17740 (N_17740,N_17489,N_17577);
nand U17741 (N_17741,N_17402,N_17546);
or U17742 (N_17742,N_17461,N_17407);
nor U17743 (N_17743,N_17513,N_17514);
nor U17744 (N_17744,N_17559,N_17407);
nor U17745 (N_17745,N_17463,N_17564);
nor U17746 (N_17746,N_17538,N_17490);
or U17747 (N_17747,N_17538,N_17424);
or U17748 (N_17748,N_17433,N_17453);
nor U17749 (N_17749,N_17543,N_17567);
xnor U17750 (N_17750,N_17423,N_17510);
and U17751 (N_17751,N_17476,N_17419);
nand U17752 (N_17752,N_17439,N_17453);
nor U17753 (N_17753,N_17452,N_17554);
and U17754 (N_17754,N_17450,N_17433);
nor U17755 (N_17755,N_17473,N_17463);
xor U17756 (N_17756,N_17485,N_17582);
nand U17757 (N_17757,N_17483,N_17523);
xor U17758 (N_17758,N_17459,N_17485);
or U17759 (N_17759,N_17446,N_17536);
nand U17760 (N_17760,N_17555,N_17513);
nor U17761 (N_17761,N_17412,N_17477);
and U17762 (N_17762,N_17415,N_17516);
nor U17763 (N_17763,N_17495,N_17424);
or U17764 (N_17764,N_17464,N_17499);
nor U17765 (N_17765,N_17559,N_17460);
and U17766 (N_17766,N_17533,N_17457);
xnor U17767 (N_17767,N_17491,N_17411);
or U17768 (N_17768,N_17408,N_17477);
xnor U17769 (N_17769,N_17532,N_17540);
nor U17770 (N_17770,N_17476,N_17474);
and U17771 (N_17771,N_17510,N_17598);
and U17772 (N_17772,N_17590,N_17409);
nor U17773 (N_17773,N_17516,N_17458);
xor U17774 (N_17774,N_17530,N_17489);
or U17775 (N_17775,N_17435,N_17452);
xnor U17776 (N_17776,N_17572,N_17549);
nand U17777 (N_17777,N_17442,N_17527);
xor U17778 (N_17778,N_17406,N_17540);
nor U17779 (N_17779,N_17569,N_17455);
xnor U17780 (N_17780,N_17418,N_17537);
nand U17781 (N_17781,N_17546,N_17553);
xor U17782 (N_17782,N_17590,N_17592);
nor U17783 (N_17783,N_17591,N_17538);
or U17784 (N_17784,N_17596,N_17561);
nand U17785 (N_17785,N_17452,N_17412);
nand U17786 (N_17786,N_17489,N_17428);
nor U17787 (N_17787,N_17510,N_17435);
nand U17788 (N_17788,N_17420,N_17556);
nor U17789 (N_17789,N_17501,N_17418);
or U17790 (N_17790,N_17438,N_17588);
or U17791 (N_17791,N_17534,N_17581);
xnor U17792 (N_17792,N_17513,N_17465);
and U17793 (N_17793,N_17556,N_17538);
xnor U17794 (N_17794,N_17499,N_17445);
nand U17795 (N_17795,N_17417,N_17502);
or U17796 (N_17796,N_17487,N_17472);
nand U17797 (N_17797,N_17550,N_17412);
nor U17798 (N_17798,N_17591,N_17464);
or U17799 (N_17799,N_17403,N_17507);
nand U17800 (N_17800,N_17745,N_17723);
nand U17801 (N_17801,N_17749,N_17759);
and U17802 (N_17802,N_17754,N_17651);
or U17803 (N_17803,N_17764,N_17696);
or U17804 (N_17804,N_17770,N_17683);
nand U17805 (N_17805,N_17733,N_17757);
nor U17806 (N_17806,N_17736,N_17741);
or U17807 (N_17807,N_17619,N_17701);
and U17808 (N_17808,N_17797,N_17767);
xnor U17809 (N_17809,N_17780,N_17628);
nand U17810 (N_17810,N_17667,N_17747);
nand U17811 (N_17811,N_17661,N_17671);
nand U17812 (N_17812,N_17756,N_17617);
xor U17813 (N_17813,N_17714,N_17607);
xor U17814 (N_17814,N_17717,N_17602);
nand U17815 (N_17815,N_17760,N_17758);
nor U17816 (N_17816,N_17703,N_17734);
or U17817 (N_17817,N_17687,N_17684);
nand U17818 (N_17818,N_17621,N_17689);
xnor U17819 (N_17819,N_17752,N_17640);
xor U17820 (N_17820,N_17601,N_17694);
nand U17821 (N_17821,N_17730,N_17707);
or U17822 (N_17822,N_17784,N_17670);
or U17823 (N_17823,N_17665,N_17704);
nand U17824 (N_17824,N_17765,N_17709);
nor U17825 (N_17825,N_17698,N_17654);
nor U17826 (N_17826,N_17750,N_17720);
nand U17827 (N_17827,N_17719,N_17708);
and U17828 (N_17828,N_17663,N_17630);
nand U17829 (N_17829,N_17695,N_17612);
nor U17830 (N_17830,N_17637,N_17716);
nor U17831 (N_17831,N_17674,N_17682);
or U17832 (N_17832,N_17715,N_17680);
or U17833 (N_17833,N_17693,N_17664);
xnor U17834 (N_17834,N_17632,N_17669);
nor U17835 (N_17835,N_17699,N_17657);
xor U17836 (N_17836,N_17610,N_17722);
nor U17837 (N_17837,N_17748,N_17614);
xnor U17838 (N_17838,N_17629,N_17773);
xor U17839 (N_17839,N_17761,N_17666);
xnor U17840 (N_17840,N_17660,N_17691);
xor U17841 (N_17841,N_17678,N_17799);
xor U17842 (N_17842,N_17721,N_17737);
and U17843 (N_17843,N_17606,N_17725);
and U17844 (N_17844,N_17774,N_17726);
xor U17845 (N_17845,N_17739,N_17755);
nand U17846 (N_17846,N_17727,N_17772);
or U17847 (N_17847,N_17681,N_17616);
xor U17848 (N_17848,N_17600,N_17627);
or U17849 (N_17849,N_17753,N_17624);
or U17850 (N_17850,N_17635,N_17743);
nor U17851 (N_17851,N_17643,N_17702);
nand U17852 (N_17852,N_17718,N_17650);
or U17853 (N_17853,N_17731,N_17705);
nand U17854 (N_17854,N_17613,N_17677);
or U17855 (N_17855,N_17762,N_17679);
nor U17856 (N_17856,N_17796,N_17798);
and U17857 (N_17857,N_17769,N_17639);
nand U17858 (N_17858,N_17644,N_17634);
or U17859 (N_17859,N_17655,N_17692);
nor U17860 (N_17860,N_17778,N_17633);
or U17861 (N_17861,N_17649,N_17668);
or U17862 (N_17862,N_17771,N_17700);
and U17863 (N_17863,N_17740,N_17648);
and U17864 (N_17864,N_17738,N_17656);
nor U17865 (N_17865,N_17751,N_17776);
and U17866 (N_17866,N_17779,N_17789);
nand U17867 (N_17867,N_17609,N_17673);
nor U17868 (N_17868,N_17615,N_17646);
xnor U17869 (N_17869,N_17729,N_17786);
nand U17870 (N_17870,N_17686,N_17685);
and U17871 (N_17871,N_17623,N_17712);
nor U17872 (N_17872,N_17653,N_17645);
nand U17873 (N_17873,N_17710,N_17782);
nand U17874 (N_17874,N_17631,N_17790);
nor U17875 (N_17875,N_17728,N_17794);
or U17876 (N_17876,N_17647,N_17697);
and U17877 (N_17877,N_17795,N_17706);
xor U17878 (N_17878,N_17688,N_17775);
nand U17879 (N_17879,N_17605,N_17611);
and U17880 (N_17880,N_17652,N_17724);
xnor U17881 (N_17881,N_17626,N_17787);
and U17882 (N_17882,N_17636,N_17608);
xnor U17883 (N_17883,N_17785,N_17659);
nor U17884 (N_17884,N_17622,N_17791);
and U17885 (N_17885,N_17711,N_17603);
and U17886 (N_17886,N_17690,N_17788);
xnor U17887 (N_17887,N_17777,N_17713);
and U17888 (N_17888,N_17618,N_17641);
or U17889 (N_17889,N_17742,N_17793);
or U17890 (N_17890,N_17604,N_17625);
nor U17891 (N_17891,N_17783,N_17675);
and U17892 (N_17892,N_17768,N_17662);
xnor U17893 (N_17893,N_17781,N_17642);
or U17894 (N_17894,N_17658,N_17676);
and U17895 (N_17895,N_17732,N_17735);
and U17896 (N_17896,N_17638,N_17620);
nor U17897 (N_17897,N_17744,N_17763);
or U17898 (N_17898,N_17792,N_17766);
xnor U17899 (N_17899,N_17672,N_17746);
nand U17900 (N_17900,N_17703,N_17756);
nand U17901 (N_17901,N_17652,N_17662);
nand U17902 (N_17902,N_17749,N_17636);
and U17903 (N_17903,N_17648,N_17774);
or U17904 (N_17904,N_17694,N_17604);
nand U17905 (N_17905,N_17600,N_17764);
nor U17906 (N_17906,N_17736,N_17728);
or U17907 (N_17907,N_17737,N_17657);
and U17908 (N_17908,N_17669,N_17737);
nand U17909 (N_17909,N_17633,N_17738);
xor U17910 (N_17910,N_17718,N_17766);
nand U17911 (N_17911,N_17690,N_17617);
nand U17912 (N_17912,N_17602,N_17715);
or U17913 (N_17913,N_17630,N_17612);
or U17914 (N_17914,N_17635,N_17628);
or U17915 (N_17915,N_17680,N_17690);
nand U17916 (N_17916,N_17622,N_17698);
xor U17917 (N_17917,N_17644,N_17775);
and U17918 (N_17918,N_17615,N_17683);
and U17919 (N_17919,N_17705,N_17651);
xor U17920 (N_17920,N_17778,N_17722);
nor U17921 (N_17921,N_17607,N_17674);
xnor U17922 (N_17922,N_17796,N_17626);
xnor U17923 (N_17923,N_17776,N_17794);
xor U17924 (N_17924,N_17636,N_17763);
nand U17925 (N_17925,N_17791,N_17686);
or U17926 (N_17926,N_17717,N_17651);
and U17927 (N_17927,N_17740,N_17634);
xnor U17928 (N_17928,N_17674,N_17738);
and U17929 (N_17929,N_17630,N_17620);
nand U17930 (N_17930,N_17655,N_17777);
and U17931 (N_17931,N_17741,N_17646);
xnor U17932 (N_17932,N_17763,N_17616);
nor U17933 (N_17933,N_17741,N_17694);
or U17934 (N_17934,N_17790,N_17748);
or U17935 (N_17935,N_17609,N_17662);
and U17936 (N_17936,N_17708,N_17664);
nand U17937 (N_17937,N_17637,N_17799);
and U17938 (N_17938,N_17667,N_17702);
nand U17939 (N_17939,N_17781,N_17790);
nand U17940 (N_17940,N_17749,N_17691);
nand U17941 (N_17941,N_17661,N_17616);
xnor U17942 (N_17942,N_17782,N_17692);
and U17943 (N_17943,N_17671,N_17726);
and U17944 (N_17944,N_17723,N_17683);
or U17945 (N_17945,N_17643,N_17704);
or U17946 (N_17946,N_17606,N_17668);
or U17947 (N_17947,N_17706,N_17649);
nor U17948 (N_17948,N_17766,N_17605);
xor U17949 (N_17949,N_17743,N_17758);
and U17950 (N_17950,N_17723,N_17601);
or U17951 (N_17951,N_17772,N_17685);
xnor U17952 (N_17952,N_17735,N_17631);
or U17953 (N_17953,N_17797,N_17753);
nand U17954 (N_17954,N_17727,N_17643);
or U17955 (N_17955,N_17775,N_17746);
or U17956 (N_17956,N_17692,N_17797);
or U17957 (N_17957,N_17705,N_17797);
and U17958 (N_17958,N_17711,N_17649);
xor U17959 (N_17959,N_17617,N_17759);
nand U17960 (N_17960,N_17741,N_17631);
nor U17961 (N_17961,N_17689,N_17696);
xnor U17962 (N_17962,N_17745,N_17715);
or U17963 (N_17963,N_17654,N_17704);
nand U17964 (N_17964,N_17658,N_17656);
and U17965 (N_17965,N_17629,N_17776);
and U17966 (N_17966,N_17751,N_17628);
or U17967 (N_17967,N_17780,N_17709);
and U17968 (N_17968,N_17718,N_17690);
nor U17969 (N_17969,N_17792,N_17725);
or U17970 (N_17970,N_17706,N_17671);
nor U17971 (N_17971,N_17658,N_17797);
xnor U17972 (N_17972,N_17790,N_17721);
xnor U17973 (N_17973,N_17742,N_17602);
and U17974 (N_17974,N_17723,N_17626);
xor U17975 (N_17975,N_17791,N_17741);
or U17976 (N_17976,N_17735,N_17610);
xnor U17977 (N_17977,N_17799,N_17729);
or U17978 (N_17978,N_17650,N_17686);
nor U17979 (N_17979,N_17605,N_17633);
nor U17980 (N_17980,N_17763,N_17707);
xor U17981 (N_17981,N_17633,N_17773);
nor U17982 (N_17982,N_17729,N_17780);
xor U17983 (N_17983,N_17627,N_17730);
nand U17984 (N_17984,N_17763,N_17635);
xor U17985 (N_17985,N_17671,N_17629);
or U17986 (N_17986,N_17689,N_17762);
nand U17987 (N_17987,N_17759,N_17766);
nor U17988 (N_17988,N_17608,N_17727);
or U17989 (N_17989,N_17778,N_17796);
nand U17990 (N_17990,N_17739,N_17747);
xnor U17991 (N_17991,N_17753,N_17615);
nand U17992 (N_17992,N_17746,N_17762);
nor U17993 (N_17993,N_17654,N_17793);
and U17994 (N_17994,N_17675,N_17651);
and U17995 (N_17995,N_17642,N_17761);
or U17996 (N_17996,N_17777,N_17616);
or U17997 (N_17997,N_17648,N_17689);
xnor U17998 (N_17998,N_17662,N_17709);
nor U17999 (N_17999,N_17722,N_17660);
and U18000 (N_18000,N_17958,N_17934);
nor U18001 (N_18001,N_17920,N_17843);
nand U18002 (N_18002,N_17944,N_17879);
nor U18003 (N_18003,N_17922,N_17907);
nand U18004 (N_18004,N_17827,N_17955);
and U18005 (N_18005,N_17924,N_17956);
or U18006 (N_18006,N_17926,N_17847);
nor U18007 (N_18007,N_17863,N_17960);
and U18008 (N_18008,N_17851,N_17901);
and U18009 (N_18009,N_17898,N_17892);
nand U18010 (N_18010,N_17835,N_17810);
and U18011 (N_18011,N_17981,N_17989);
nand U18012 (N_18012,N_17992,N_17900);
nor U18013 (N_18013,N_17919,N_17943);
or U18014 (N_18014,N_17839,N_17821);
or U18015 (N_18015,N_17980,N_17927);
or U18016 (N_18016,N_17914,N_17931);
or U18017 (N_18017,N_17826,N_17935);
or U18018 (N_18018,N_17825,N_17804);
nand U18019 (N_18019,N_17904,N_17991);
xnor U18020 (N_18020,N_17959,N_17890);
or U18021 (N_18021,N_17942,N_17868);
or U18022 (N_18022,N_17815,N_17972);
or U18023 (N_18023,N_17853,N_17856);
nand U18024 (N_18024,N_17897,N_17984);
xor U18025 (N_18025,N_17936,N_17928);
nor U18026 (N_18026,N_17995,N_17970);
nand U18027 (N_18027,N_17923,N_17805);
or U18028 (N_18028,N_17962,N_17882);
or U18029 (N_18029,N_17941,N_17896);
or U18030 (N_18030,N_17930,N_17834);
or U18031 (N_18031,N_17961,N_17964);
and U18032 (N_18032,N_17953,N_17945);
and U18033 (N_18033,N_17933,N_17862);
nor U18034 (N_18034,N_17824,N_17977);
nand U18035 (N_18035,N_17906,N_17891);
or U18036 (N_18036,N_17800,N_17967);
or U18037 (N_18037,N_17886,N_17908);
nor U18038 (N_18038,N_17986,N_17828);
nor U18039 (N_18039,N_17939,N_17838);
xnor U18040 (N_18040,N_17867,N_17850);
nand U18041 (N_18041,N_17811,N_17903);
or U18042 (N_18042,N_17966,N_17860);
nor U18043 (N_18043,N_17905,N_17997);
nor U18044 (N_18044,N_17858,N_17899);
and U18045 (N_18045,N_17916,N_17872);
nor U18046 (N_18046,N_17932,N_17951);
xnor U18047 (N_18047,N_17874,N_17988);
and U18048 (N_18048,N_17982,N_17957);
xnor U18049 (N_18049,N_17854,N_17887);
or U18050 (N_18050,N_17975,N_17921);
xor U18051 (N_18051,N_17844,N_17983);
and U18052 (N_18052,N_17833,N_17859);
xnor U18053 (N_18053,N_17809,N_17814);
nor U18054 (N_18054,N_17974,N_17865);
or U18055 (N_18055,N_17829,N_17870);
nor U18056 (N_18056,N_17902,N_17861);
xor U18057 (N_18057,N_17893,N_17820);
and U18058 (N_18058,N_17911,N_17946);
nor U18059 (N_18059,N_17841,N_17968);
and U18060 (N_18060,N_17880,N_17813);
nand U18061 (N_18061,N_17949,N_17915);
and U18062 (N_18062,N_17855,N_17876);
nand U18063 (N_18063,N_17837,N_17971);
nor U18064 (N_18064,N_17806,N_17913);
or U18065 (N_18065,N_17987,N_17895);
nor U18066 (N_18066,N_17998,N_17999);
xor U18067 (N_18067,N_17937,N_17849);
nor U18068 (N_18068,N_17917,N_17817);
nand U18069 (N_18069,N_17969,N_17963);
xor U18070 (N_18070,N_17846,N_17918);
nor U18071 (N_18071,N_17822,N_17994);
xor U18072 (N_18072,N_17993,N_17873);
nor U18073 (N_18073,N_17973,N_17877);
and U18074 (N_18074,N_17808,N_17801);
nor U18075 (N_18075,N_17938,N_17840);
nor U18076 (N_18076,N_17812,N_17889);
nor U18077 (N_18077,N_17848,N_17912);
or U18078 (N_18078,N_17864,N_17878);
xor U18079 (N_18079,N_17909,N_17954);
or U18080 (N_18080,N_17816,N_17881);
nand U18081 (N_18081,N_17869,N_17952);
nand U18082 (N_18082,N_17985,N_17996);
xnor U18083 (N_18083,N_17842,N_17925);
and U18084 (N_18084,N_17885,N_17866);
nand U18085 (N_18085,N_17802,N_17807);
xor U18086 (N_18086,N_17857,N_17910);
xnor U18087 (N_18087,N_17888,N_17832);
nor U18088 (N_18088,N_17883,N_17852);
and U18089 (N_18089,N_17803,N_17884);
nor U18090 (N_18090,N_17990,N_17947);
xnor U18091 (N_18091,N_17875,N_17830);
or U18092 (N_18092,N_17950,N_17976);
xnor U18093 (N_18093,N_17823,N_17894);
nor U18094 (N_18094,N_17831,N_17818);
nand U18095 (N_18095,N_17845,N_17940);
nor U18096 (N_18096,N_17819,N_17978);
or U18097 (N_18097,N_17871,N_17965);
nor U18098 (N_18098,N_17929,N_17979);
nor U18099 (N_18099,N_17948,N_17836);
nand U18100 (N_18100,N_17880,N_17906);
and U18101 (N_18101,N_17822,N_17957);
xnor U18102 (N_18102,N_17935,N_17801);
and U18103 (N_18103,N_17991,N_17943);
xnor U18104 (N_18104,N_17861,N_17809);
or U18105 (N_18105,N_17999,N_17816);
nand U18106 (N_18106,N_17874,N_17848);
and U18107 (N_18107,N_17962,N_17998);
nor U18108 (N_18108,N_17894,N_17913);
and U18109 (N_18109,N_17943,N_17822);
and U18110 (N_18110,N_17833,N_17986);
xnor U18111 (N_18111,N_17928,N_17850);
or U18112 (N_18112,N_17834,N_17814);
xor U18113 (N_18113,N_17808,N_17836);
or U18114 (N_18114,N_17826,N_17945);
nand U18115 (N_18115,N_17855,N_17922);
nor U18116 (N_18116,N_17889,N_17887);
or U18117 (N_18117,N_17830,N_17968);
and U18118 (N_18118,N_17948,N_17821);
xor U18119 (N_18119,N_17814,N_17989);
and U18120 (N_18120,N_17881,N_17800);
nor U18121 (N_18121,N_17869,N_17851);
nand U18122 (N_18122,N_17999,N_17928);
nor U18123 (N_18123,N_17808,N_17858);
nor U18124 (N_18124,N_17826,N_17862);
and U18125 (N_18125,N_17811,N_17921);
xor U18126 (N_18126,N_17897,N_17967);
and U18127 (N_18127,N_17946,N_17851);
nand U18128 (N_18128,N_17817,N_17968);
xor U18129 (N_18129,N_17933,N_17819);
or U18130 (N_18130,N_17923,N_17814);
nand U18131 (N_18131,N_17943,N_17873);
nor U18132 (N_18132,N_17990,N_17943);
and U18133 (N_18133,N_17857,N_17873);
and U18134 (N_18134,N_17957,N_17830);
xor U18135 (N_18135,N_17964,N_17870);
and U18136 (N_18136,N_17851,N_17879);
nor U18137 (N_18137,N_17980,N_17813);
xnor U18138 (N_18138,N_17920,N_17996);
and U18139 (N_18139,N_17829,N_17972);
and U18140 (N_18140,N_17856,N_17881);
xnor U18141 (N_18141,N_17839,N_17802);
nand U18142 (N_18142,N_17981,N_17826);
xnor U18143 (N_18143,N_17867,N_17993);
and U18144 (N_18144,N_17823,N_17849);
and U18145 (N_18145,N_17887,N_17904);
xor U18146 (N_18146,N_17855,N_17863);
nand U18147 (N_18147,N_17831,N_17842);
nor U18148 (N_18148,N_17900,N_17820);
nor U18149 (N_18149,N_17961,N_17802);
nor U18150 (N_18150,N_17891,N_17810);
and U18151 (N_18151,N_17925,N_17821);
or U18152 (N_18152,N_17802,N_17842);
or U18153 (N_18153,N_17990,N_17900);
xor U18154 (N_18154,N_17946,N_17919);
xor U18155 (N_18155,N_17898,N_17818);
nor U18156 (N_18156,N_17882,N_17900);
or U18157 (N_18157,N_17958,N_17853);
nand U18158 (N_18158,N_17982,N_17809);
xnor U18159 (N_18159,N_17969,N_17987);
xnor U18160 (N_18160,N_17908,N_17857);
and U18161 (N_18161,N_17863,N_17853);
nor U18162 (N_18162,N_17856,N_17948);
nand U18163 (N_18163,N_17981,N_17936);
nor U18164 (N_18164,N_17948,N_17958);
and U18165 (N_18165,N_17872,N_17800);
nor U18166 (N_18166,N_17874,N_17916);
and U18167 (N_18167,N_17814,N_17816);
xor U18168 (N_18168,N_17979,N_17927);
nand U18169 (N_18169,N_17882,N_17969);
xnor U18170 (N_18170,N_17885,N_17926);
xnor U18171 (N_18171,N_17937,N_17881);
nor U18172 (N_18172,N_17993,N_17954);
nor U18173 (N_18173,N_17841,N_17981);
nand U18174 (N_18174,N_17814,N_17935);
or U18175 (N_18175,N_17967,N_17824);
nand U18176 (N_18176,N_17952,N_17931);
or U18177 (N_18177,N_17889,N_17917);
and U18178 (N_18178,N_17933,N_17998);
nand U18179 (N_18179,N_17875,N_17859);
nor U18180 (N_18180,N_17899,N_17828);
nand U18181 (N_18181,N_17914,N_17902);
or U18182 (N_18182,N_17896,N_17808);
nand U18183 (N_18183,N_17817,N_17818);
nor U18184 (N_18184,N_17885,N_17939);
xnor U18185 (N_18185,N_17806,N_17832);
nor U18186 (N_18186,N_17811,N_17927);
or U18187 (N_18187,N_17801,N_17934);
nor U18188 (N_18188,N_17992,N_17999);
nor U18189 (N_18189,N_17892,N_17824);
nor U18190 (N_18190,N_17877,N_17981);
or U18191 (N_18191,N_17980,N_17979);
nand U18192 (N_18192,N_17990,N_17879);
or U18193 (N_18193,N_17831,N_17820);
nand U18194 (N_18194,N_17961,N_17853);
xnor U18195 (N_18195,N_17940,N_17918);
nand U18196 (N_18196,N_17997,N_17943);
xor U18197 (N_18197,N_17907,N_17920);
xnor U18198 (N_18198,N_17919,N_17979);
nor U18199 (N_18199,N_17885,N_17886);
nand U18200 (N_18200,N_18152,N_18024);
xnor U18201 (N_18201,N_18131,N_18060);
nor U18202 (N_18202,N_18017,N_18035);
or U18203 (N_18203,N_18002,N_18126);
xnor U18204 (N_18204,N_18049,N_18108);
nor U18205 (N_18205,N_18170,N_18096);
xnor U18206 (N_18206,N_18164,N_18184);
nor U18207 (N_18207,N_18168,N_18116);
and U18208 (N_18208,N_18023,N_18030);
and U18209 (N_18209,N_18136,N_18122);
nor U18210 (N_18210,N_18000,N_18032);
nand U18211 (N_18211,N_18065,N_18113);
and U18212 (N_18212,N_18103,N_18193);
xnor U18213 (N_18213,N_18021,N_18061);
nor U18214 (N_18214,N_18192,N_18094);
or U18215 (N_18215,N_18140,N_18132);
or U18216 (N_18216,N_18115,N_18182);
xnor U18217 (N_18217,N_18181,N_18078);
nand U18218 (N_18218,N_18147,N_18086);
nor U18219 (N_18219,N_18073,N_18111);
nand U18220 (N_18220,N_18051,N_18134);
or U18221 (N_18221,N_18015,N_18165);
and U18222 (N_18222,N_18011,N_18027);
or U18223 (N_18223,N_18055,N_18029);
or U18224 (N_18224,N_18180,N_18123);
xor U18225 (N_18225,N_18010,N_18092);
nor U18226 (N_18226,N_18036,N_18056);
nand U18227 (N_18227,N_18037,N_18095);
xnor U18228 (N_18228,N_18185,N_18007);
nor U18229 (N_18229,N_18106,N_18117);
nor U18230 (N_18230,N_18171,N_18133);
nor U18231 (N_18231,N_18158,N_18169);
nor U18232 (N_18232,N_18150,N_18098);
nor U18233 (N_18233,N_18105,N_18137);
or U18234 (N_18234,N_18082,N_18101);
xnor U18235 (N_18235,N_18160,N_18154);
xor U18236 (N_18236,N_18197,N_18173);
nand U18237 (N_18237,N_18198,N_18059);
and U18238 (N_18238,N_18179,N_18124);
nor U18239 (N_18239,N_18167,N_18139);
nand U18240 (N_18240,N_18144,N_18074);
or U18241 (N_18241,N_18058,N_18174);
nand U18242 (N_18242,N_18004,N_18039);
nor U18243 (N_18243,N_18044,N_18042);
nor U18244 (N_18244,N_18025,N_18149);
xnor U18245 (N_18245,N_18048,N_18166);
xor U18246 (N_18246,N_18083,N_18163);
nand U18247 (N_18247,N_18033,N_18156);
nand U18248 (N_18248,N_18148,N_18102);
or U18249 (N_18249,N_18142,N_18090);
nor U18250 (N_18250,N_18138,N_18091);
and U18251 (N_18251,N_18088,N_18031);
or U18252 (N_18252,N_18189,N_18014);
and U18253 (N_18253,N_18062,N_18008);
and U18254 (N_18254,N_18177,N_18112);
nand U18255 (N_18255,N_18079,N_18043);
or U18256 (N_18256,N_18087,N_18072);
xor U18257 (N_18257,N_18018,N_18012);
and U18258 (N_18258,N_18034,N_18199);
xnor U18259 (N_18259,N_18068,N_18127);
or U18260 (N_18260,N_18028,N_18041);
and U18261 (N_18261,N_18064,N_18069);
or U18262 (N_18262,N_18155,N_18130);
and U18263 (N_18263,N_18005,N_18070);
nor U18264 (N_18264,N_18019,N_18047);
nor U18265 (N_18265,N_18063,N_18040);
or U18266 (N_18266,N_18084,N_18097);
xnor U18267 (N_18267,N_18110,N_18120);
and U18268 (N_18268,N_18071,N_18172);
nor U18269 (N_18269,N_18178,N_18162);
xor U18270 (N_18270,N_18145,N_18186);
and U18271 (N_18271,N_18038,N_18175);
and U18272 (N_18272,N_18080,N_18066);
xnor U18273 (N_18273,N_18052,N_18057);
xor U18274 (N_18274,N_18075,N_18125);
nor U18275 (N_18275,N_18194,N_18129);
and U18276 (N_18276,N_18195,N_18081);
nor U18277 (N_18277,N_18104,N_18020);
nor U18278 (N_18278,N_18016,N_18067);
nor U18279 (N_18279,N_18159,N_18188);
nand U18280 (N_18280,N_18146,N_18006);
xnor U18281 (N_18281,N_18187,N_18157);
xor U18282 (N_18282,N_18076,N_18053);
and U18283 (N_18283,N_18128,N_18161);
nor U18284 (N_18284,N_18022,N_18013);
nor U18285 (N_18285,N_18143,N_18109);
nor U18286 (N_18286,N_18190,N_18100);
or U18287 (N_18287,N_18099,N_18141);
xor U18288 (N_18288,N_18114,N_18085);
or U18289 (N_18289,N_18191,N_18050);
xnor U18290 (N_18290,N_18077,N_18026);
nor U18291 (N_18291,N_18176,N_18093);
nand U18292 (N_18292,N_18045,N_18121);
nand U18293 (N_18293,N_18046,N_18001);
nand U18294 (N_18294,N_18135,N_18183);
xor U18295 (N_18295,N_18153,N_18107);
or U18296 (N_18296,N_18054,N_18196);
or U18297 (N_18297,N_18151,N_18003);
or U18298 (N_18298,N_18009,N_18089);
nand U18299 (N_18299,N_18119,N_18118);
nor U18300 (N_18300,N_18100,N_18181);
xor U18301 (N_18301,N_18100,N_18108);
xor U18302 (N_18302,N_18117,N_18169);
or U18303 (N_18303,N_18187,N_18038);
xor U18304 (N_18304,N_18137,N_18155);
xnor U18305 (N_18305,N_18153,N_18034);
nor U18306 (N_18306,N_18141,N_18038);
nor U18307 (N_18307,N_18189,N_18077);
xnor U18308 (N_18308,N_18175,N_18132);
or U18309 (N_18309,N_18059,N_18179);
and U18310 (N_18310,N_18140,N_18066);
nor U18311 (N_18311,N_18123,N_18195);
and U18312 (N_18312,N_18035,N_18082);
nor U18313 (N_18313,N_18132,N_18097);
nand U18314 (N_18314,N_18075,N_18032);
xnor U18315 (N_18315,N_18088,N_18029);
or U18316 (N_18316,N_18047,N_18093);
xor U18317 (N_18317,N_18033,N_18171);
nand U18318 (N_18318,N_18155,N_18182);
and U18319 (N_18319,N_18179,N_18041);
nand U18320 (N_18320,N_18112,N_18094);
and U18321 (N_18321,N_18159,N_18024);
or U18322 (N_18322,N_18041,N_18086);
and U18323 (N_18323,N_18181,N_18188);
nor U18324 (N_18324,N_18034,N_18163);
xnor U18325 (N_18325,N_18017,N_18175);
or U18326 (N_18326,N_18119,N_18007);
nand U18327 (N_18327,N_18056,N_18169);
xnor U18328 (N_18328,N_18168,N_18082);
nand U18329 (N_18329,N_18156,N_18187);
nand U18330 (N_18330,N_18078,N_18123);
or U18331 (N_18331,N_18042,N_18102);
nor U18332 (N_18332,N_18158,N_18013);
nand U18333 (N_18333,N_18167,N_18157);
or U18334 (N_18334,N_18039,N_18069);
or U18335 (N_18335,N_18112,N_18031);
or U18336 (N_18336,N_18030,N_18004);
nand U18337 (N_18337,N_18152,N_18187);
nand U18338 (N_18338,N_18197,N_18046);
nand U18339 (N_18339,N_18105,N_18071);
and U18340 (N_18340,N_18044,N_18129);
nand U18341 (N_18341,N_18079,N_18180);
and U18342 (N_18342,N_18115,N_18051);
nor U18343 (N_18343,N_18094,N_18062);
or U18344 (N_18344,N_18018,N_18081);
or U18345 (N_18345,N_18079,N_18002);
and U18346 (N_18346,N_18196,N_18088);
and U18347 (N_18347,N_18063,N_18140);
nand U18348 (N_18348,N_18066,N_18050);
xor U18349 (N_18349,N_18175,N_18005);
nand U18350 (N_18350,N_18088,N_18195);
xnor U18351 (N_18351,N_18168,N_18048);
nor U18352 (N_18352,N_18032,N_18113);
nand U18353 (N_18353,N_18053,N_18110);
and U18354 (N_18354,N_18044,N_18092);
nor U18355 (N_18355,N_18193,N_18025);
nor U18356 (N_18356,N_18089,N_18056);
nand U18357 (N_18357,N_18109,N_18151);
and U18358 (N_18358,N_18047,N_18045);
or U18359 (N_18359,N_18164,N_18013);
xnor U18360 (N_18360,N_18165,N_18055);
nand U18361 (N_18361,N_18045,N_18123);
nor U18362 (N_18362,N_18079,N_18118);
xnor U18363 (N_18363,N_18171,N_18194);
xor U18364 (N_18364,N_18191,N_18002);
nor U18365 (N_18365,N_18008,N_18032);
or U18366 (N_18366,N_18177,N_18101);
and U18367 (N_18367,N_18095,N_18169);
nand U18368 (N_18368,N_18023,N_18158);
nand U18369 (N_18369,N_18091,N_18095);
or U18370 (N_18370,N_18169,N_18130);
and U18371 (N_18371,N_18047,N_18143);
xor U18372 (N_18372,N_18055,N_18099);
nand U18373 (N_18373,N_18034,N_18166);
xor U18374 (N_18374,N_18001,N_18030);
nand U18375 (N_18375,N_18093,N_18114);
xnor U18376 (N_18376,N_18046,N_18177);
nor U18377 (N_18377,N_18156,N_18119);
nor U18378 (N_18378,N_18088,N_18120);
and U18379 (N_18379,N_18065,N_18074);
nand U18380 (N_18380,N_18138,N_18022);
nand U18381 (N_18381,N_18006,N_18085);
or U18382 (N_18382,N_18061,N_18039);
xnor U18383 (N_18383,N_18073,N_18035);
and U18384 (N_18384,N_18170,N_18016);
xnor U18385 (N_18385,N_18179,N_18184);
nand U18386 (N_18386,N_18099,N_18123);
nand U18387 (N_18387,N_18076,N_18001);
xor U18388 (N_18388,N_18131,N_18153);
or U18389 (N_18389,N_18102,N_18020);
or U18390 (N_18390,N_18181,N_18139);
nor U18391 (N_18391,N_18050,N_18160);
nor U18392 (N_18392,N_18022,N_18071);
nor U18393 (N_18393,N_18102,N_18087);
or U18394 (N_18394,N_18045,N_18122);
nand U18395 (N_18395,N_18135,N_18060);
xor U18396 (N_18396,N_18034,N_18132);
or U18397 (N_18397,N_18129,N_18199);
xor U18398 (N_18398,N_18161,N_18180);
xnor U18399 (N_18399,N_18040,N_18161);
xnor U18400 (N_18400,N_18237,N_18278);
nand U18401 (N_18401,N_18223,N_18352);
nor U18402 (N_18402,N_18357,N_18208);
nor U18403 (N_18403,N_18262,N_18320);
nand U18404 (N_18404,N_18318,N_18205);
and U18405 (N_18405,N_18319,N_18231);
xnor U18406 (N_18406,N_18292,N_18350);
nand U18407 (N_18407,N_18326,N_18203);
nor U18408 (N_18408,N_18244,N_18232);
nor U18409 (N_18409,N_18343,N_18202);
nor U18410 (N_18410,N_18282,N_18314);
or U18411 (N_18411,N_18209,N_18315);
nand U18412 (N_18412,N_18396,N_18340);
nand U18413 (N_18413,N_18269,N_18386);
and U18414 (N_18414,N_18291,N_18226);
and U18415 (N_18415,N_18236,N_18338);
nor U18416 (N_18416,N_18302,N_18275);
or U18417 (N_18417,N_18361,N_18222);
and U18418 (N_18418,N_18240,N_18309);
nand U18419 (N_18419,N_18200,N_18267);
and U18420 (N_18420,N_18329,N_18252);
nand U18421 (N_18421,N_18362,N_18331);
nor U18422 (N_18422,N_18288,N_18299);
and U18423 (N_18423,N_18294,N_18251);
and U18424 (N_18424,N_18347,N_18254);
nand U18425 (N_18425,N_18364,N_18349);
or U18426 (N_18426,N_18397,N_18284);
and U18427 (N_18427,N_18399,N_18368);
and U18428 (N_18428,N_18287,N_18286);
and U18429 (N_18429,N_18334,N_18253);
or U18430 (N_18430,N_18384,N_18298);
nor U18431 (N_18431,N_18215,N_18241);
nand U18432 (N_18432,N_18374,N_18395);
and U18433 (N_18433,N_18247,N_18392);
nand U18434 (N_18434,N_18276,N_18359);
or U18435 (N_18435,N_18367,N_18233);
nand U18436 (N_18436,N_18274,N_18266);
xor U18437 (N_18437,N_18207,N_18280);
or U18438 (N_18438,N_18210,N_18375);
nor U18439 (N_18439,N_18213,N_18295);
xor U18440 (N_18440,N_18256,N_18304);
xor U18441 (N_18441,N_18307,N_18211);
and U18442 (N_18442,N_18379,N_18279);
xnor U18443 (N_18443,N_18249,N_18393);
nand U18444 (N_18444,N_18370,N_18313);
nand U18445 (N_18445,N_18344,N_18355);
or U18446 (N_18446,N_18268,N_18212);
and U18447 (N_18447,N_18265,N_18325);
and U18448 (N_18448,N_18238,N_18248);
and U18449 (N_18449,N_18301,N_18218);
or U18450 (N_18450,N_18376,N_18380);
nand U18451 (N_18451,N_18354,N_18271);
and U18452 (N_18452,N_18214,N_18257);
and U18453 (N_18453,N_18259,N_18342);
xnor U18454 (N_18454,N_18303,N_18322);
and U18455 (N_18455,N_18391,N_18371);
or U18456 (N_18456,N_18270,N_18328);
and U18457 (N_18457,N_18337,N_18348);
xnor U18458 (N_18458,N_18378,N_18297);
nand U18459 (N_18459,N_18216,N_18220);
nand U18460 (N_18460,N_18281,N_18312);
nand U18461 (N_18461,N_18333,N_18332);
nand U18462 (N_18462,N_18385,N_18221);
or U18463 (N_18463,N_18227,N_18388);
and U18464 (N_18464,N_18234,N_18390);
or U18465 (N_18465,N_18243,N_18273);
nand U18466 (N_18466,N_18365,N_18263);
xnor U18467 (N_18467,N_18306,N_18296);
xor U18468 (N_18468,N_18356,N_18327);
or U18469 (N_18469,N_18235,N_18217);
nor U18470 (N_18470,N_18353,N_18289);
and U18471 (N_18471,N_18394,N_18339);
and U18472 (N_18472,N_18383,N_18311);
nand U18473 (N_18473,N_18317,N_18398);
nor U18474 (N_18474,N_18283,N_18246);
xnor U18475 (N_18475,N_18201,N_18285);
nand U18476 (N_18476,N_18366,N_18230);
nand U18477 (N_18477,N_18219,N_18377);
or U18478 (N_18478,N_18358,N_18372);
or U18479 (N_18479,N_18239,N_18321);
nand U18480 (N_18480,N_18228,N_18310);
nor U18481 (N_18481,N_18335,N_18324);
nor U18482 (N_18482,N_18389,N_18255);
or U18483 (N_18483,N_18204,N_18373);
and U18484 (N_18484,N_18225,N_18260);
nor U18485 (N_18485,N_18316,N_18261);
or U18486 (N_18486,N_18272,N_18250);
nand U18487 (N_18487,N_18229,N_18323);
xor U18488 (N_18488,N_18258,N_18346);
or U18489 (N_18489,N_18382,N_18242);
nand U18490 (N_18490,N_18245,N_18341);
xor U18491 (N_18491,N_18369,N_18264);
nand U18492 (N_18492,N_18363,N_18360);
nor U18493 (N_18493,N_18206,N_18351);
nand U18494 (N_18494,N_18308,N_18345);
nand U18495 (N_18495,N_18277,N_18224);
xnor U18496 (N_18496,N_18336,N_18330);
or U18497 (N_18497,N_18300,N_18305);
and U18498 (N_18498,N_18290,N_18293);
or U18499 (N_18499,N_18381,N_18387);
nor U18500 (N_18500,N_18297,N_18260);
nor U18501 (N_18501,N_18211,N_18306);
xnor U18502 (N_18502,N_18221,N_18235);
nand U18503 (N_18503,N_18356,N_18329);
nand U18504 (N_18504,N_18252,N_18392);
or U18505 (N_18505,N_18390,N_18284);
xor U18506 (N_18506,N_18275,N_18361);
nand U18507 (N_18507,N_18236,N_18298);
nand U18508 (N_18508,N_18341,N_18201);
or U18509 (N_18509,N_18310,N_18328);
nand U18510 (N_18510,N_18308,N_18370);
nor U18511 (N_18511,N_18326,N_18252);
and U18512 (N_18512,N_18223,N_18219);
nand U18513 (N_18513,N_18343,N_18385);
nor U18514 (N_18514,N_18274,N_18381);
nor U18515 (N_18515,N_18322,N_18317);
or U18516 (N_18516,N_18307,N_18236);
or U18517 (N_18517,N_18321,N_18277);
xnor U18518 (N_18518,N_18230,N_18212);
nor U18519 (N_18519,N_18383,N_18259);
xnor U18520 (N_18520,N_18302,N_18382);
or U18521 (N_18521,N_18372,N_18391);
and U18522 (N_18522,N_18351,N_18314);
or U18523 (N_18523,N_18333,N_18348);
nor U18524 (N_18524,N_18394,N_18271);
nand U18525 (N_18525,N_18380,N_18318);
nor U18526 (N_18526,N_18334,N_18381);
nor U18527 (N_18527,N_18396,N_18314);
nor U18528 (N_18528,N_18300,N_18342);
nand U18529 (N_18529,N_18360,N_18204);
xnor U18530 (N_18530,N_18343,N_18352);
and U18531 (N_18531,N_18320,N_18338);
xor U18532 (N_18532,N_18374,N_18292);
and U18533 (N_18533,N_18264,N_18257);
and U18534 (N_18534,N_18292,N_18391);
nor U18535 (N_18535,N_18358,N_18323);
or U18536 (N_18536,N_18227,N_18306);
or U18537 (N_18537,N_18263,N_18231);
or U18538 (N_18538,N_18368,N_18298);
nand U18539 (N_18539,N_18295,N_18385);
nand U18540 (N_18540,N_18234,N_18356);
and U18541 (N_18541,N_18387,N_18377);
nor U18542 (N_18542,N_18290,N_18218);
and U18543 (N_18543,N_18359,N_18252);
xnor U18544 (N_18544,N_18392,N_18346);
or U18545 (N_18545,N_18349,N_18209);
nand U18546 (N_18546,N_18357,N_18397);
or U18547 (N_18547,N_18208,N_18214);
and U18548 (N_18548,N_18257,N_18274);
xor U18549 (N_18549,N_18351,N_18245);
nor U18550 (N_18550,N_18270,N_18332);
or U18551 (N_18551,N_18224,N_18317);
xor U18552 (N_18552,N_18317,N_18298);
and U18553 (N_18553,N_18396,N_18262);
xnor U18554 (N_18554,N_18365,N_18399);
xnor U18555 (N_18555,N_18333,N_18340);
nor U18556 (N_18556,N_18333,N_18321);
nor U18557 (N_18557,N_18371,N_18289);
nand U18558 (N_18558,N_18355,N_18259);
nand U18559 (N_18559,N_18206,N_18220);
or U18560 (N_18560,N_18221,N_18373);
xor U18561 (N_18561,N_18253,N_18380);
nand U18562 (N_18562,N_18344,N_18361);
and U18563 (N_18563,N_18392,N_18334);
nor U18564 (N_18564,N_18242,N_18378);
or U18565 (N_18565,N_18298,N_18219);
nand U18566 (N_18566,N_18386,N_18352);
and U18567 (N_18567,N_18317,N_18399);
and U18568 (N_18568,N_18221,N_18200);
or U18569 (N_18569,N_18248,N_18351);
nor U18570 (N_18570,N_18370,N_18286);
or U18571 (N_18571,N_18285,N_18280);
nor U18572 (N_18572,N_18354,N_18363);
nand U18573 (N_18573,N_18374,N_18218);
nor U18574 (N_18574,N_18248,N_18232);
xor U18575 (N_18575,N_18297,N_18344);
or U18576 (N_18576,N_18214,N_18297);
or U18577 (N_18577,N_18304,N_18251);
xor U18578 (N_18578,N_18347,N_18251);
nand U18579 (N_18579,N_18397,N_18389);
xor U18580 (N_18580,N_18320,N_18301);
xor U18581 (N_18581,N_18212,N_18327);
nor U18582 (N_18582,N_18262,N_18249);
xnor U18583 (N_18583,N_18268,N_18216);
nor U18584 (N_18584,N_18369,N_18351);
xor U18585 (N_18585,N_18249,N_18260);
nor U18586 (N_18586,N_18312,N_18395);
and U18587 (N_18587,N_18345,N_18384);
xor U18588 (N_18588,N_18243,N_18350);
and U18589 (N_18589,N_18327,N_18217);
nor U18590 (N_18590,N_18353,N_18242);
xor U18591 (N_18591,N_18347,N_18273);
and U18592 (N_18592,N_18296,N_18293);
nor U18593 (N_18593,N_18303,N_18234);
and U18594 (N_18594,N_18396,N_18222);
nor U18595 (N_18595,N_18290,N_18204);
nand U18596 (N_18596,N_18233,N_18354);
nand U18597 (N_18597,N_18210,N_18336);
nor U18598 (N_18598,N_18259,N_18314);
or U18599 (N_18599,N_18209,N_18309);
or U18600 (N_18600,N_18466,N_18591);
nor U18601 (N_18601,N_18557,N_18577);
xor U18602 (N_18602,N_18400,N_18531);
xor U18603 (N_18603,N_18428,N_18496);
nand U18604 (N_18604,N_18538,N_18569);
nor U18605 (N_18605,N_18437,N_18404);
nand U18606 (N_18606,N_18424,N_18581);
nor U18607 (N_18607,N_18490,N_18588);
nor U18608 (N_18608,N_18590,N_18516);
xnor U18609 (N_18609,N_18498,N_18527);
xor U18610 (N_18610,N_18461,N_18559);
nand U18611 (N_18611,N_18578,N_18426);
or U18612 (N_18612,N_18505,N_18526);
nand U18613 (N_18613,N_18599,N_18440);
xor U18614 (N_18614,N_18471,N_18584);
xor U18615 (N_18615,N_18510,N_18512);
or U18616 (N_18616,N_18481,N_18525);
and U18617 (N_18617,N_18415,N_18451);
xnor U18618 (N_18618,N_18521,N_18450);
xnor U18619 (N_18619,N_18488,N_18585);
and U18620 (N_18620,N_18592,N_18519);
and U18621 (N_18621,N_18537,N_18432);
xor U18622 (N_18622,N_18473,N_18572);
nand U18623 (N_18623,N_18463,N_18555);
xor U18624 (N_18624,N_18552,N_18460);
xnor U18625 (N_18625,N_18542,N_18541);
xor U18626 (N_18626,N_18595,N_18467);
nor U18627 (N_18627,N_18545,N_18598);
or U18628 (N_18628,N_18554,N_18507);
nor U18629 (N_18629,N_18430,N_18586);
nand U18630 (N_18630,N_18532,N_18412);
nand U18631 (N_18631,N_18582,N_18539);
nand U18632 (N_18632,N_18534,N_18427);
or U18633 (N_18633,N_18580,N_18436);
nor U18634 (N_18634,N_18503,N_18423);
xnor U18635 (N_18635,N_18594,N_18402);
or U18636 (N_18636,N_18504,N_18449);
or U18637 (N_18637,N_18434,N_18459);
nor U18638 (N_18638,N_18597,N_18579);
xor U18639 (N_18639,N_18435,N_18566);
and U18640 (N_18640,N_18522,N_18462);
and U18641 (N_18641,N_18442,N_18421);
nor U18642 (N_18642,N_18484,N_18411);
nor U18643 (N_18643,N_18403,N_18487);
xor U18644 (N_18644,N_18414,N_18517);
and U18645 (N_18645,N_18506,N_18468);
xnor U18646 (N_18646,N_18509,N_18520);
nor U18647 (N_18647,N_18474,N_18448);
and U18648 (N_18648,N_18530,N_18493);
and U18649 (N_18649,N_18553,N_18438);
xor U18650 (N_18650,N_18413,N_18406);
or U18651 (N_18651,N_18514,N_18518);
and U18652 (N_18652,N_18533,N_18422);
xnor U18653 (N_18653,N_18429,N_18464);
or U18654 (N_18654,N_18575,N_18445);
xor U18655 (N_18655,N_18433,N_18556);
nor U18656 (N_18656,N_18513,N_18441);
nand U18657 (N_18657,N_18573,N_18465);
xor U18658 (N_18658,N_18478,N_18529);
nand U18659 (N_18659,N_18455,N_18407);
and U18660 (N_18660,N_18563,N_18535);
nand U18661 (N_18661,N_18476,N_18405);
nor U18662 (N_18662,N_18540,N_18502);
or U18663 (N_18663,N_18523,N_18494);
or U18664 (N_18664,N_18447,N_18486);
nor U18665 (N_18665,N_18475,N_18508);
nor U18666 (N_18666,N_18596,N_18470);
xnor U18667 (N_18667,N_18562,N_18408);
xor U18668 (N_18668,N_18558,N_18479);
or U18669 (N_18669,N_18564,N_18492);
nand U18670 (N_18670,N_18547,N_18551);
nor U18671 (N_18671,N_18458,N_18567);
xnor U18672 (N_18672,N_18528,N_18544);
nor U18673 (N_18673,N_18524,N_18401);
or U18674 (N_18674,N_18500,N_18477);
nor U18675 (N_18675,N_18560,N_18495);
xnor U18676 (N_18676,N_18420,N_18483);
nor U18677 (N_18677,N_18571,N_18565);
nor U18678 (N_18678,N_18431,N_18446);
nor U18679 (N_18679,N_18568,N_18469);
and U18680 (N_18680,N_18491,N_18444);
nand U18681 (N_18681,N_18417,N_18548);
and U18682 (N_18682,N_18418,N_18480);
xor U18683 (N_18683,N_18576,N_18589);
nand U18684 (N_18684,N_18515,N_18536);
nand U18685 (N_18685,N_18543,N_18416);
nand U18686 (N_18686,N_18425,N_18499);
nor U18687 (N_18687,N_18549,N_18419);
nor U18688 (N_18688,N_18570,N_18457);
or U18689 (N_18689,N_18443,N_18587);
nand U18690 (N_18690,N_18454,N_18583);
or U18691 (N_18691,N_18489,N_18550);
nor U18692 (N_18692,N_18497,N_18472);
or U18693 (N_18693,N_18593,N_18452);
nand U18694 (N_18694,N_18485,N_18561);
nor U18695 (N_18695,N_18456,N_18511);
nand U18696 (N_18696,N_18439,N_18482);
and U18697 (N_18697,N_18501,N_18546);
nand U18698 (N_18698,N_18410,N_18409);
nand U18699 (N_18699,N_18453,N_18574);
nor U18700 (N_18700,N_18455,N_18445);
and U18701 (N_18701,N_18429,N_18441);
nor U18702 (N_18702,N_18427,N_18576);
nand U18703 (N_18703,N_18523,N_18540);
and U18704 (N_18704,N_18457,N_18465);
nor U18705 (N_18705,N_18471,N_18494);
nand U18706 (N_18706,N_18459,N_18530);
and U18707 (N_18707,N_18445,N_18404);
or U18708 (N_18708,N_18489,N_18440);
or U18709 (N_18709,N_18450,N_18572);
nand U18710 (N_18710,N_18507,N_18559);
or U18711 (N_18711,N_18452,N_18574);
and U18712 (N_18712,N_18495,N_18504);
and U18713 (N_18713,N_18410,N_18447);
nor U18714 (N_18714,N_18400,N_18402);
nor U18715 (N_18715,N_18587,N_18519);
or U18716 (N_18716,N_18442,N_18581);
xnor U18717 (N_18717,N_18481,N_18571);
and U18718 (N_18718,N_18464,N_18407);
nand U18719 (N_18719,N_18459,N_18443);
and U18720 (N_18720,N_18546,N_18455);
or U18721 (N_18721,N_18557,N_18461);
nor U18722 (N_18722,N_18577,N_18527);
or U18723 (N_18723,N_18577,N_18589);
and U18724 (N_18724,N_18430,N_18440);
and U18725 (N_18725,N_18428,N_18475);
xnor U18726 (N_18726,N_18577,N_18455);
xnor U18727 (N_18727,N_18584,N_18449);
nand U18728 (N_18728,N_18419,N_18518);
nor U18729 (N_18729,N_18450,N_18411);
xnor U18730 (N_18730,N_18564,N_18550);
or U18731 (N_18731,N_18446,N_18417);
nand U18732 (N_18732,N_18495,N_18523);
nand U18733 (N_18733,N_18440,N_18593);
xnor U18734 (N_18734,N_18597,N_18465);
xnor U18735 (N_18735,N_18563,N_18515);
nand U18736 (N_18736,N_18518,N_18444);
or U18737 (N_18737,N_18426,N_18479);
nor U18738 (N_18738,N_18543,N_18462);
nand U18739 (N_18739,N_18515,N_18435);
nand U18740 (N_18740,N_18487,N_18578);
nor U18741 (N_18741,N_18527,N_18570);
and U18742 (N_18742,N_18563,N_18415);
xnor U18743 (N_18743,N_18431,N_18532);
xnor U18744 (N_18744,N_18405,N_18499);
or U18745 (N_18745,N_18543,N_18443);
nor U18746 (N_18746,N_18554,N_18456);
nand U18747 (N_18747,N_18464,N_18514);
nor U18748 (N_18748,N_18478,N_18517);
nor U18749 (N_18749,N_18535,N_18471);
or U18750 (N_18750,N_18486,N_18570);
and U18751 (N_18751,N_18597,N_18421);
and U18752 (N_18752,N_18446,N_18456);
and U18753 (N_18753,N_18416,N_18519);
or U18754 (N_18754,N_18416,N_18429);
nor U18755 (N_18755,N_18566,N_18535);
or U18756 (N_18756,N_18452,N_18456);
or U18757 (N_18757,N_18491,N_18461);
xnor U18758 (N_18758,N_18545,N_18445);
nand U18759 (N_18759,N_18536,N_18454);
or U18760 (N_18760,N_18423,N_18437);
or U18761 (N_18761,N_18405,N_18475);
or U18762 (N_18762,N_18407,N_18576);
nor U18763 (N_18763,N_18551,N_18440);
or U18764 (N_18764,N_18512,N_18459);
nor U18765 (N_18765,N_18461,N_18504);
nor U18766 (N_18766,N_18597,N_18517);
nand U18767 (N_18767,N_18518,N_18587);
and U18768 (N_18768,N_18506,N_18441);
and U18769 (N_18769,N_18422,N_18586);
nor U18770 (N_18770,N_18425,N_18512);
nor U18771 (N_18771,N_18591,N_18580);
nand U18772 (N_18772,N_18559,N_18489);
and U18773 (N_18773,N_18462,N_18577);
and U18774 (N_18774,N_18557,N_18429);
or U18775 (N_18775,N_18415,N_18582);
and U18776 (N_18776,N_18483,N_18545);
xnor U18777 (N_18777,N_18435,N_18443);
and U18778 (N_18778,N_18467,N_18548);
and U18779 (N_18779,N_18429,N_18467);
nor U18780 (N_18780,N_18506,N_18509);
or U18781 (N_18781,N_18528,N_18577);
nand U18782 (N_18782,N_18528,N_18476);
nor U18783 (N_18783,N_18444,N_18572);
xor U18784 (N_18784,N_18540,N_18524);
nor U18785 (N_18785,N_18414,N_18547);
nor U18786 (N_18786,N_18483,N_18588);
nor U18787 (N_18787,N_18530,N_18555);
nand U18788 (N_18788,N_18459,N_18494);
and U18789 (N_18789,N_18409,N_18477);
nand U18790 (N_18790,N_18482,N_18476);
xnor U18791 (N_18791,N_18589,N_18567);
nand U18792 (N_18792,N_18519,N_18500);
nand U18793 (N_18793,N_18572,N_18466);
nor U18794 (N_18794,N_18439,N_18528);
and U18795 (N_18795,N_18576,N_18450);
nor U18796 (N_18796,N_18417,N_18442);
nor U18797 (N_18797,N_18544,N_18445);
nand U18798 (N_18798,N_18580,N_18495);
or U18799 (N_18799,N_18557,N_18450);
or U18800 (N_18800,N_18755,N_18621);
nor U18801 (N_18801,N_18600,N_18625);
xnor U18802 (N_18802,N_18751,N_18614);
and U18803 (N_18803,N_18689,N_18602);
or U18804 (N_18804,N_18736,N_18762);
and U18805 (N_18805,N_18799,N_18604);
or U18806 (N_18806,N_18764,N_18745);
nand U18807 (N_18807,N_18617,N_18649);
nor U18808 (N_18808,N_18644,N_18633);
and U18809 (N_18809,N_18671,N_18746);
and U18810 (N_18810,N_18609,N_18712);
or U18811 (N_18811,N_18628,N_18668);
and U18812 (N_18812,N_18629,N_18687);
and U18813 (N_18813,N_18682,N_18646);
or U18814 (N_18814,N_18631,N_18678);
and U18815 (N_18815,N_18697,N_18605);
nand U18816 (N_18816,N_18722,N_18721);
or U18817 (N_18817,N_18684,N_18620);
and U18818 (N_18818,N_18793,N_18695);
and U18819 (N_18819,N_18707,N_18653);
nand U18820 (N_18820,N_18661,N_18703);
or U18821 (N_18821,N_18761,N_18640);
nor U18822 (N_18822,N_18723,N_18619);
and U18823 (N_18823,N_18692,N_18641);
or U18824 (N_18824,N_18654,N_18665);
nand U18825 (N_18825,N_18685,N_18622);
nor U18826 (N_18826,N_18716,N_18601);
nor U18827 (N_18827,N_18713,N_18709);
and U18828 (N_18828,N_18776,N_18710);
and U18829 (N_18829,N_18794,N_18626);
nor U18830 (N_18830,N_18650,N_18750);
nor U18831 (N_18831,N_18663,N_18708);
xnor U18832 (N_18832,N_18786,N_18611);
xnor U18833 (N_18833,N_18765,N_18769);
nand U18834 (N_18834,N_18796,N_18742);
nor U18835 (N_18835,N_18696,N_18766);
and U18836 (N_18836,N_18730,N_18787);
xor U18837 (N_18837,N_18676,N_18792);
or U18838 (N_18838,N_18795,N_18731);
nor U18839 (N_18839,N_18694,N_18674);
or U18840 (N_18840,N_18733,N_18760);
or U18841 (N_18841,N_18637,N_18777);
nor U18842 (N_18842,N_18771,N_18666);
nor U18843 (N_18843,N_18747,N_18789);
and U18844 (N_18844,N_18706,N_18607);
nand U18845 (N_18845,N_18748,N_18680);
nand U18846 (N_18846,N_18784,N_18632);
nor U18847 (N_18847,N_18691,N_18711);
xnor U18848 (N_18848,N_18701,N_18627);
xnor U18849 (N_18849,N_18624,N_18683);
nor U18850 (N_18850,N_18639,N_18659);
nor U18851 (N_18851,N_18774,N_18752);
nor U18852 (N_18852,N_18749,N_18727);
or U18853 (N_18853,N_18648,N_18744);
and U18854 (N_18854,N_18634,N_18688);
nand U18855 (N_18855,N_18705,N_18616);
nor U18856 (N_18856,N_18737,N_18642);
nor U18857 (N_18857,N_18728,N_18652);
nand U18858 (N_18858,N_18655,N_18606);
or U18859 (N_18859,N_18781,N_18779);
nor U18860 (N_18860,N_18636,N_18788);
nor U18861 (N_18861,N_18724,N_18719);
and U18862 (N_18862,N_18767,N_18657);
or U18863 (N_18863,N_18759,N_18756);
xor U18864 (N_18864,N_18690,N_18726);
and U18865 (N_18865,N_18613,N_18686);
xnor U18866 (N_18866,N_18673,N_18638);
nor U18867 (N_18867,N_18720,N_18772);
nand U18868 (N_18868,N_18718,N_18656);
nor U18869 (N_18869,N_18700,N_18635);
nand U18870 (N_18870,N_18735,N_18768);
and U18871 (N_18871,N_18757,N_18675);
and U18872 (N_18872,N_18739,N_18729);
nand U18873 (N_18873,N_18754,N_18725);
xor U18874 (N_18874,N_18603,N_18791);
or U18875 (N_18875,N_18658,N_18660);
nand U18876 (N_18876,N_18790,N_18797);
xor U18877 (N_18877,N_18782,N_18643);
xor U18878 (N_18878,N_18698,N_18669);
xnor U18879 (N_18879,N_18670,N_18679);
nor U18880 (N_18880,N_18667,N_18645);
nand U18881 (N_18881,N_18681,N_18647);
nor U18882 (N_18882,N_18783,N_18662);
or U18883 (N_18883,N_18741,N_18715);
nor U18884 (N_18884,N_18714,N_18610);
or U18885 (N_18885,N_18734,N_18758);
nor U18886 (N_18886,N_18798,N_18740);
nand U18887 (N_18887,N_18743,N_18763);
nor U18888 (N_18888,N_18732,N_18623);
or U18889 (N_18889,N_18699,N_18717);
nand U18890 (N_18890,N_18775,N_18608);
or U18891 (N_18891,N_18753,N_18704);
nand U18892 (N_18892,N_18693,N_18664);
xor U18893 (N_18893,N_18738,N_18702);
or U18894 (N_18894,N_18618,N_18773);
and U18895 (N_18895,N_18770,N_18615);
nor U18896 (N_18896,N_18651,N_18677);
or U18897 (N_18897,N_18785,N_18672);
nor U18898 (N_18898,N_18780,N_18630);
or U18899 (N_18899,N_18778,N_18612);
xor U18900 (N_18900,N_18687,N_18699);
and U18901 (N_18901,N_18786,N_18661);
or U18902 (N_18902,N_18656,N_18643);
and U18903 (N_18903,N_18673,N_18731);
nand U18904 (N_18904,N_18762,N_18613);
and U18905 (N_18905,N_18650,N_18667);
nand U18906 (N_18906,N_18776,N_18731);
xnor U18907 (N_18907,N_18725,N_18709);
nand U18908 (N_18908,N_18762,N_18653);
and U18909 (N_18909,N_18786,N_18798);
xor U18910 (N_18910,N_18774,N_18771);
nand U18911 (N_18911,N_18666,N_18684);
nand U18912 (N_18912,N_18740,N_18703);
xnor U18913 (N_18913,N_18745,N_18704);
and U18914 (N_18914,N_18660,N_18665);
xnor U18915 (N_18915,N_18608,N_18675);
and U18916 (N_18916,N_18632,N_18664);
nand U18917 (N_18917,N_18612,N_18667);
xor U18918 (N_18918,N_18799,N_18738);
nand U18919 (N_18919,N_18788,N_18777);
or U18920 (N_18920,N_18728,N_18761);
nor U18921 (N_18921,N_18703,N_18701);
or U18922 (N_18922,N_18735,N_18750);
xnor U18923 (N_18923,N_18667,N_18649);
nand U18924 (N_18924,N_18607,N_18695);
or U18925 (N_18925,N_18771,N_18785);
nor U18926 (N_18926,N_18779,N_18607);
nor U18927 (N_18927,N_18767,N_18685);
nand U18928 (N_18928,N_18785,N_18660);
nand U18929 (N_18929,N_18784,N_18749);
xnor U18930 (N_18930,N_18750,N_18709);
and U18931 (N_18931,N_18628,N_18736);
nor U18932 (N_18932,N_18628,N_18732);
nor U18933 (N_18933,N_18611,N_18631);
or U18934 (N_18934,N_18752,N_18787);
or U18935 (N_18935,N_18709,N_18759);
nor U18936 (N_18936,N_18613,N_18609);
and U18937 (N_18937,N_18797,N_18692);
or U18938 (N_18938,N_18775,N_18736);
nor U18939 (N_18939,N_18710,N_18674);
or U18940 (N_18940,N_18610,N_18793);
or U18941 (N_18941,N_18741,N_18794);
and U18942 (N_18942,N_18735,N_18740);
or U18943 (N_18943,N_18615,N_18714);
and U18944 (N_18944,N_18600,N_18626);
xor U18945 (N_18945,N_18733,N_18796);
xor U18946 (N_18946,N_18710,N_18635);
xor U18947 (N_18947,N_18713,N_18799);
nor U18948 (N_18948,N_18792,N_18693);
and U18949 (N_18949,N_18688,N_18786);
or U18950 (N_18950,N_18654,N_18628);
and U18951 (N_18951,N_18644,N_18773);
xor U18952 (N_18952,N_18768,N_18615);
nand U18953 (N_18953,N_18621,N_18747);
nor U18954 (N_18954,N_18629,N_18636);
nor U18955 (N_18955,N_18782,N_18758);
nor U18956 (N_18956,N_18743,N_18607);
nor U18957 (N_18957,N_18621,N_18785);
nor U18958 (N_18958,N_18757,N_18650);
and U18959 (N_18959,N_18701,N_18795);
xor U18960 (N_18960,N_18651,N_18619);
nor U18961 (N_18961,N_18762,N_18777);
or U18962 (N_18962,N_18769,N_18678);
or U18963 (N_18963,N_18707,N_18615);
and U18964 (N_18964,N_18677,N_18683);
nand U18965 (N_18965,N_18782,N_18673);
xor U18966 (N_18966,N_18773,N_18764);
or U18967 (N_18967,N_18682,N_18797);
nand U18968 (N_18968,N_18685,N_18613);
and U18969 (N_18969,N_18733,N_18750);
xor U18970 (N_18970,N_18647,N_18699);
or U18971 (N_18971,N_18762,N_18673);
and U18972 (N_18972,N_18739,N_18652);
nand U18973 (N_18973,N_18779,N_18745);
nand U18974 (N_18974,N_18604,N_18742);
or U18975 (N_18975,N_18693,N_18704);
nor U18976 (N_18976,N_18654,N_18726);
nor U18977 (N_18977,N_18692,N_18771);
or U18978 (N_18978,N_18731,N_18796);
or U18979 (N_18979,N_18744,N_18733);
xor U18980 (N_18980,N_18689,N_18694);
nand U18981 (N_18981,N_18796,N_18717);
nand U18982 (N_18982,N_18786,N_18765);
nor U18983 (N_18983,N_18679,N_18731);
nor U18984 (N_18984,N_18612,N_18729);
and U18985 (N_18985,N_18713,N_18662);
nand U18986 (N_18986,N_18734,N_18792);
xnor U18987 (N_18987,N_18671,N_18619);
or U18988 (N_18988,N_18781,N_18725);
and U18989 (N_18989,N_18796,N_18774);
and U18990 (N_18990,N_18738,N_18640);
and U18991 (N_18991,N_18784,N_18615);
nor U18992 (N_18992,N_18659,N_18634);
nor U18993 (N_18993,N_18726,N_18664);
and U18994 (N_18994,N_18675,N_18710);
nor U18995 (N_18995,N_18770,N_18731);
nor U18996 (N_18996,N_18765,N_18744);
nor U18997 (N_18997,N_18739,N_18709);
nor U18998 (N_18998,N_18617,N_18765);
nand U18999 (N_18999,N_18631,N_18616);
and U19000 (N_19000,N_18852,N_18897);
nor U19001 (N_19001,N_18913,N_18864);
nand U19002 (N_19002,N_18837,N_18804);
or U19003 (N_19003,N_18912,N_18896);
or U19004 (N_19004,N_18898,N_18857);
or U19005 (N_19005,N_18949,N_18978);
and U19006 (N_19006,N_18989,N_18809);
nand U19007 (N_19007,N_18942,N_18819);
or U19008 (N_19008,N_18840,N_18848);
and U19009 (N_19009,N_18824,N_18854);
nand U19010 (N_19010,N_18827,N_18881);
or U19011 (N_19011,N_18903,N_18810);
xor U19012 (N_19012,N_18836,N_18880);
xnor U19013 (N_19013,N_18966,N_18980);
or U19014 (N_19014,N_18862,N_18958);
nand U19015 (N_19015,N_18919,N_18917);
and U19016 (N_19016,N_18872,N_18944);
nand U19017 (N_19017,N_18952,N_18843);
nor U19018 (N_19018,N_18983,N_18877);
nand U19019 (N_19019,N_18911,N_18990);
and U19020 (N_19020,N_18988,N_18879);
and U19021 (N_19021,N_18977,N_18850);
or U19022 (N_19022,N_18930,N_18856);
or U19023 (N_19023,N_18891,N_18860);
and U19024 (N_19024,N_18950,N_18847);
and U19025 (N_19025,N_18982,N_18932);
xor U19026 (N_19026,N_18825,N_18866);
xnor U19027 (N_19027,N_18956,N_18985);
or U19028 (N_19028,N_18907,N_18961);
xor U19029 (N_19029,N_18914,N_18986);
or U19030 (N_19030,N_18935,N_18939);
and U19031 (N_19031,N_18931,N_18933);
nand U19032 (N_19032,N_18905,N_18899);
or U19033 (N_19033,N_18839,N_18938);
or U19034 (N_19034,N_18883,N_18865);
and U19035 (N_19035,N_18916,N_18926);
nand U19036 (N_19036,N_18820,N_18833);
xnor U19037 (N_19037,N_18909,N_18981);
nand U19038 (N_19038,N_18946,N_18993);
xnor U19039 (N_19039,N_18936,N_18940);
nand U19040 (N_19040,N_18995,N_18947);
or U19041 (N_19041,N_18889,N_18876);
nor U19042 (N_19042,N_18828,N_18984);
xnor U19043 (N_19043,N_18871,N_18967);
xnor U19044 (N_19044,N_18934,N_18972);
nor U19045 (N_19045,N_18953,N_18975);
or U19046 (N_19046,N_18813,N_18979);
and U19047 (N_19047,N_18875,N_18969);
or U19048 (N_19048,N_18849,N_18832);
and U19049 (N_19049,N_18888,N_18948);
nand U19050 (N_19050,N_18920,N_18838);
xor U19051 (N_19051,N_18830,N_18929);
or U19052 (N_19052,N_18844,N_18915);
nand U19053 (N_19053,N_18968,N_18823);
or U19054 (N_19054,N_18970,N_18957);
nand U19055 (N_19055,N_18811,N_18999);
nand U19056 (N_19056,N_18816,N_18894);
nor U19057 (N_19057,N_18800,N_18976);
nor U19058 (N_19058,N_18885,N_18951);
and U19059 (N_19059,N_18831,N_18812);
or U19060 (N_19060,N_18846,N_18807);
or U19061 (N_19061,N_18893,N_18895);
nor U19062 (N_19062,N_18806,N_18867);
xnor U19063 (N_19063,N_18863,N_18884);
and U19064 (N_19064,N_18964,N_18902);
nor U19065 (N_19065,N_18924,N_18887);
nor U19066 (N_19066,N_18861,N_18815);
or U19067 (N_19067,N_18996,N_18965);
nand U19068 (N_19068,N_18817,N_18808);
nand U19069 (N_19069,N_18925,N_18826);
nand U19070 (N_19070,N_18987,N_18900);
nor U19071 (N_19071,N_18959,N_18835);
nand U19072 (N_19072,N_18801,N_18998);
nor U19073 (N_19073,N_18921,N_18937);
nand U19074 (N_19074,N_18873,N_18878);
nor U19075 (N_19075,N_18906,N_18822);
xor U19076 (N_19076,N_18927,N_18997);
xor U19077 (N_19077,N_18992,N_18960);
nand U19078 (N_19078,N_18928,N_18802);
and U19079 (N_19079,N_18886,N_18974);
nor U19080 (N_19080,N_18834,N_18955);
and U19081 (N_19081,N_18901,N_18904);
xor U19082 (N_19082,N_18818,N_18910);
or U19083 (N_19083,N_18851,N_18954);
and U19084 (N_19084,N_18853,N_18962);
nand U19085 (N_19085,N_18973,N_18945);
and U19086 (N_19086,N_18814,N_18845);
nand U19087 (N_19087,N_18890,N_18918);
xor U19088 (N_19088,N_18923,N_18943);
or U19089 (N_19089,N_18941,N_18829);
nand U19090 (N_19090,N_18991,N_18922);
nand U19091 (N_19091,N_18971,N_18994);
nand U19092 (N_19092,N_18870,N_18805);
xnor U19093 (N_19093,N_18908,N_18874);
or U19094 (N_19094,N_18859,N_18869);
nor U19095 (N_19095,N_18821,N_18855);
nand U19096 (N_19096,N_18963,N_18841);
and U19097 (N_19097,N_18882,N_18892);
nor U19098 (N_19098,N_18858,N_18803);
nor U19099 (N_19099,N_18868,N_18842);
nand U19100 (N_19100,N_18919,N_18957);
nand U19101 (N_19101,N_18826,N_18850);
nor U19102 (N_19102,N_18878,N_18994);
nor U19103 (N_19103,N_18979,N_18984);
nand U19104 (N_19104,N_18830,N_18975);
xnor U19105 (N_19105,N_18961,N_18897);
nand U19106 (N_19106,N_18916,N_18869);
and U19107 (N_19107,N_18883,N_18977);
xor U19108 (N_19108,N_18903,N_18808);
nor U19109 (N_19109,N_18835,N_18841);
xnor U19110 (N_19110,N_18937,N_18862);
nand U19111 (N_19111,N_18891,N_18867);
nand U19112 (N_19112,N_18950,N_18806);
nand U19113 (N_19113,N_18949,N_18858);
nor U19114 (N_19114,N_18812,N_18863);
nand U19115 (N_19115,N_18899,N_18895);
and U19116 (N_19116,N_18811,N_18948);
nand U19117 (N_19117,N_18960,N_18857);
and U19118 (N_19118,N_18865,N_18845);
or U19119 (N_19119,N_18942,N_18900);
or U19120 (N_19120,N_18979,N_18930);
xor U19121 (N_19121,N_18895,N_18858);
nor U19122 (N_19122,N_18892,N_18933);
or U19123 (N_19123,N_18913,N_18870);
or U19124 (N_19124,N_18816,N_18965);
and U19125 (N_19125,N_18922,N_18872);
xnor U19126 (N_19126,N_18984,N_18834);
or U19127 (N_19127,N_18880,N_18982);
nand U19128 (N_19128,N_18809,N_18807);
nand U19129 (N_19129,N_18885,N_18803);
nand U19130 (N_19130,N_18954,N_18994);
nand U19131 (N_19131,N_18828,N_18903);
or U19132 (N_19132,N_18878,N_18995);
or U19133 (N_19133,N_18929,N_18934);
nor U19134 (N_19134,N_18869,N_18938);
xnor U19135 (N_19135,N_18823,N_18996);
or U19136 (N_19136,N_18906,N_18954);
xor U19137 (N_19137,N_18977,N_18888);
xor U19138 (N_19138,N_18861,N_18841);
nor U19139 (N_19139,N_18818,N_18977);
or U19140 (N_19140,N_18847,N_18944);
nor U19141 (N_19141,N_18880,N_18994);
nand U19142 (N_19142,N_18867,N_18972);
xnor U19143 (N_19143,N_18938,N_18996);
nor U19144 (N_19144,N_18844,N_18835);
and U19145 (N_19145,N_18958,N_18900);
or U19146 (N_19146,N_18895,N_18860);
and U19147 (N_19147,N_18889,N_18910);
nor U19148 (N_19148,N_18805,N_18888);
nor U19149 (N_19149,N_18843,N_18967);
xnor U19150 (N_19150,N_18803,N_18901);
xnor U19151 (N_19151,N_18876,N_18838);
nor U19152 (N_19152,N_18950,N_18944);
or U19153 (N_19153,N_18977,N_18894);
xnor U19154 (N_19154,N_18965,N_18896);
or U19155 (N_19155,N_18961,N_18899);
nand U19156 (N_19156,N_18842,N_18870);
nand U19157 (N_19157,N_18884,N_18841);
nand U19158 (N_19158,N_18877,N_18999);
or U19159 (N_19159,N_18949,N_18825);
and U19160 (N_19160,N_18977,N_18852);
and U19161 (N_19161,N_18970,N_18868);
nand U19162 (N_19162,N_18991,N_18999);
or U19163 (N_19163,N_18948,N_18946);
xnor U19164 (N_19164,N_18884,N_18808);
nor U19165 (N_19165,N_18818,N_18837);
or U19166 (N_19166,N_18965,N_18813);
nor U19167 (N_19167,N_18962,N_18873);
and U19168 (N_19168,N_18999,N_18887);
xnor U19169 (N_19169,N_18972,N_18940);
and U19170 (N_19170,N_18864,N_18862);
nor U19171 (N_19171,N_18945,N_18866);
nor U19172 (N_19172,N_18913,N_18938);
xnor U19173 (N_19173,N_18955,N_18900);
xor U19174 (N_19174,N_18928,N_18929);
nand U19175 (N_19175,N_18841,N_18810);
nand U19176 (N_19176,N_18852,N_18816);
and U19177 (N_19177,N_18960,N_18801);
and U19178 (N_19178,N_18980,N_18899);
and U19179 (N_19179,N_18942,N_18830);
nor U19180 (N_19180,N_18969,N_18937);
and U19181 (N_19181,N_18810,N_18974);
nor U19182 (N_19182,N_18952,N_18888);
and U19183 (N_19183,N_18985,N_18979);
or U19184 (N_19184,N_18858,N_18919);
xor U19185 (N_19185,N_18830,N_18815);
xnor U19186 (N_19186,N_18994,N_18822);
nor U19187 (N_19187,N_18914,N_18952);
or U19188 (N_19188,N_18864,N_18980);
nand U19189 (N_19189,N_18951,N_18849);
nor U19190 (N_19190,N_18941,N_18935);
xor U19191 (N_19191,N_18943,N_18969);
and U19192 (N_19192,N_18803,N_18868);
nand U19193 (N_19193,N_18981,N_18982);
nand U19194 (N_19194,N_18828,N_18908);
and U19195 (N_19195,N_18955,N_18847);
nor U19196 (N_19196,N_18834,N_18827);
nor U19197 (N_19197,N_18859,N_18865);
nor U19198 (N_19198,N_18878,N_18992);
and U19199 (N_19199,N_18929,N_18996);
xnor U19200 (N_19200,N_19041,N_19134);
or U19201 (N_19201,N_19170,N_19193);
or U19202 (N_19202,N_19045,N_19051);
nand U19203 (N_19203,N_19007,N_19077);
nand U19204 (N_19204,N_19130,N_19160);
nand U19205 (N_19205,N_19139,N_19164);
xnor U19206 (N_19206,N_19017,N_19064);
and U19207 (N_19207,N_19011,N_19083);
nand U19208 (N_19208,N_19123,N_19026);
and U19209 (N_19209,N_19122,N_19060);
xor U19210 (N_19210,N_19150,N_19132);
nand U19211 (N_19211,N_19096,N_19165);
or U19212 (N_19212,N_19102,N_19043);
xnor U19213 (N_19213,N_19162,N_19100);
nor U19214 (N_19214,N_19167,N_19035);
and U19215 (N_19215,N_19095,N_19014);
nand U19216 (N_19216,N_19019,N_19036);
or U19217 (N_19217,N_19144,N_19110);
xor U19218 (N_19218,N_19016,N_19173);
nand U19219 (N_19219,N_19010,N_19161);
and U19220 (N_19220,N_19079,N_19156);
or U19221 (N_19221,N_19091,N_19154);
and U19222 (N_19222,N_19056,N_19199);
nor U19223 (N_19223,N_19135,N_19053);
nand U19224 (N_19224,N_19190,N_19074);
xor U19225 (N_19225,N_19148,N_19000);
and U19226 (N_19226,N_19046,N_19128);
and U19227 (N_19227,N_19040,N_19001);
and U19228 (N_19228,N_19089,N_19068);
or U19229 (N_19229,N_19142,N_19039);
nand U19230 (N_19230,N_19143,N_19188);
nand U19231 (N_19231,N_19052,N_19197);
and U19232 (N_19232,N_19071,N_19157);
and U19233 (N_19233,N_19153,N_19012);
or U19234 (N_19234,N_19070,N_19159);
or U19235 (N_19235,N_19196,N_19112);
or U19236 (N_19236,N_19120,N_19126);
xnor U19237 (N_19237,N_19129,N_19048);
nor U19238 (N_19238,N_19082,N_19006);
nor U19239 (N_19239,N_19168,N_19054);
nand U19240 (N_19240,N_19088,N_19186);
nor U19241 (N_19241,N_19192,N_19030);
nand U19242 (N_19242,N_19034,N_19169);
nor U19243 (N_19243,N_19184,N_19166);
nand U19244 (N_19244,N_19015,N_19103);
or U19245 (N_19245,N_19076,N_19085);
or U19246 (N_19246,N_19124,N_19177);
nor U19247 (N_19247,N_19013,N_19158);
nand U19248 (N_19248,N_19063,N_19059);
and U19249 (N_19249,N_19055,N_19058);
or U19250 (N_19250,N_19018,N_19020);
or U19251 (N_19251,N_19118,N_19114);
xor U19252 (N_19252,N_19140,N_19025);
xor U19253 (N_19253,N_19176,N_19028);
nand U19254 (N_19254,N_19133,N_19042);
or U19255 (N_19255,N_19024,N_19141);
xnor U19256 (N_19256,N_19147,N_19104);
nor U19257 (N_19257,N_19065,N_19049);
or U19258 (N_19258,N_19174,N_19099);
nor U19259 (N_19259,N_19137,N_19131);
or U19260 (N_19260,N_19090,N_19163);
xnor U19261 (N_19261,N_19080,N_19119);
xor U19262 (N_19262,N_19037,N_19109);
nand U19263 (N_19263,N_19061,N_19097);
or U19264 (N_19264,N_19149,N_19022);
nor U19265 (N_19265,N_19194,N_19152);
nand U19266 (N_19266,N_19179,N_19044);
xnor U19267 (N_19267,N_19111,N_19138);
xnor U19268 (N_19268,N_19032,N_19023);
xnor U19269 (N_19269,N_19008,N_19182);
nor U19270 (N_19270,N_19066,N_19062);
nor U19271 (N_19271,N_19187,N_19106);
xor U19272 (N_19272,N_19004,N_19107);
nor U19273 (N_19273,N_19072,N_19151);
or U19274 (N_19274,N_19189,N_19191);
or U19275 (N_19275,N_19003,N_19092);
and U19276 (N_19276,N_19005,N_19108);
nand U19277 (N_19277,N_19069,N_19093);
or U19278 (N_19278,N_19021,N_19027);
nand U19279 (N_19279,N_19145,N_19031);
or U19280 (N_19280,N_19009,N_19101);
or U19281 (N_19281,N_19098,N_19127);
xnor U19282 (N_19282,N_19175,N_19075);
or U19283 (N_19283,N_19181,N_19002);
or U19284 (N_19284,N_19195,N_19105);
nand U19285 (N_19285,N_19050,N_19198);
nor U19286 (N_19286,N_19029,N_19185);
and U19287 (N_19287,N_19146,N_19094);
or U19288 (N_19288,N_19136,N_19121);
nand U19289 (N_19289,N_19172,N_19180);
and U19290 (N_19290,N_19057,N_19067);
nand U19291 (N_19291,N_19047,N_19087);
and U19292 (N_19292,N_19178,N_19033);
nand U19293 (N_19293,N_19116,N_19117);
or U19294 (N_19294,N_19113,N_19125);
or U19295 (N_19295,N_19155,N_19081);
xnor U19296 (N_19296,N_19078,N_19084);
and U19297 (N_19297,N_19038,N_19171);
nor U19298 (N_19298,N_19086,N_19183);
nor U19299 (N_19299,N_19073,N_19115);
nand U19300 (N_19300,N_19088,N_19003);
and U19301 (N_19301,N_19135,N_19190);
xnor U19302 (N_19302,N_19072,N_19168);
xnor U19303 (N_19303,N_19178,N_19199);
or U19304 (N_19304,N_19121,N_19070);
nor U19305 (N_19305,N_19084,N_19132);
and U19306 (N_19306,N_19131,N_19181);
nor U19307 (N_19307,N_19058,N_19195);
xnor U19308 (N_19308,N_19026,N_19138);
xor U19309 (N_19309,N_19015,N_19006);
or U19310 (N_19310,N_19164,N_19115);
nand U19311 (N_19311,N_19088,N_19064);
or U19312 (N_19312,N_19136,N_19005);
and U19313 (N_19313,N_19165,N_19052);
nand U19314 (N_19314,N_19006,N_19145);
or U19315 (N_19315,N_19142,N_19128);
and U19316 (N_19316,N_19018,N_19194);
nand U19317 (N_19317,N_19053,N_19098);
xnor U19318 (N_19318,N_19078,N_19171);
or U19319 (N_19319,N_19128,N_19179);
nor U19320 (N_19320,N_19169,N_19177);
xor U19321 (N_19321,N_19133,N_19062);
nand U19322 (N_19322,N_19009,N_19170);
or U19323 (N_19323,N_19038,N_19159);
nand U19324 (N_19324,N_19056,N_19154);
nor U19325 (N_19325,N_19163,N_19059);
nor U19326 (N_19326,N_19120,N_19053);
xor U19327 (N_19327,N_19192,N_19029);
xor U19328 (N_19328,N_19104,N_19012);
or U19329 (N_19329,N_19059,N_19085);
xor U19330 (N_19330,N_19102,N_19038);
and U19331 (N_19331,N_19011,N_19099);
nand U19332 (N_19332,N_19110,N_19035);
xor U19333 (N_19333,N_19146,N_19154);
and U19334 (N_19334,N_19158,N_19199);
or U19335 (N_19335,N_19118,N_19025);
or U19336 (N_19336,N_19082,N_19001);
and U19337 (N_19337,N_19085,N_19169);
or U19338 (N_19338,N_19086,N_19161);
xor U19339 (N_19339,N_19195,N_19049);
nand U19340 (N_19340,N_19092,N_19072);
and U19341 (N_19341,N_19084,N_19129);
nor U19342 (N_19342,N_19030,N_19070);
nor U19343 (N_19343,N_19010,N_19137);
and U19344 (N_19344,N_19059,N_19034);
nand U19345 (N_19345,N_19003,N_19035);
nor U19346 (N_19346,N_19006,N_19049);
nand U19347 (N_19347,N_19033,N_19052);
nand U19348 (N_19348,N_19172,N_19075);
and U19349 (N_19349,N_19128,N_19169);
or U19350 (N_19350,N_19136,N_19163);
or U19351 (N_19351,N_19024,N_19035);
or U19352 (N_19352,N_19140,N_19196);
and U19353 (N_19353,N_19007,N_19118);
nand U19354 (N_19354,N_19181,N_19059);
nor U19355 (N_19355,N_19093,N_19096);
xor U19356 (N_19356,N_19095,N_19111);
nor U19357 (N_19357,N_19076,N_19198);
and U19358 (N_19358,N_19050,N_19119);
or U19359 (N_19359,N_19113,N_19075);
and U19360 (N_19360,N_19011,N_19089);
and U19361 (N_19361,N_19190,N_19117);
and U19362 (N_19362,N_19003,N_19048);
and U19363 (N_19363,N_19128,N_19139);
nand U19364 (N_19364,N_19161,N_19152);
or U19365 (N_19365,N_19153,N_19090);
nor U19366 (N_19366,N_19101,N_19131);
xor U19367 (N_19367,N_19036,N_19113);
nor U19368 (N_19368,N_19189,N_19118);
nand U19369 (N_19369,N_19114,N_19091);
and U19370 (N_19370,N_19058,N_19183);
nor U19371 (N_19371,N_19161,N_19130);
nor U19372 (N_19372,N_19072,N_19170);
nand U19373 (N_19373,N_19058,N_19138);
nor U19374 (N_19374,N_19104,N_19181);
nor U19375 (N_19375,N_19134,N_19172);
or U19376 (N_19376,N_19154,N_19119);
nor U19377 (N_19377,N_19115,N_19179);
xnor U19378 (N_19378,N_19002,N_19068);
and U19379 (N_19379,N_19105,N_19059);
xnor U19380 (N_19380,N_19004,N_19161);
xnor U19381 (N_19381,N_19075,N_19146);
nor U19382 (N_19382,N_19066,N_19159);
nor U19383 (N_19383,N_19083,N_19106);
xor U19384 (N_19384,N_19165,N_19140);
nor U19385 (N_19385,N_19047,N_19095);
and U19386 (N_19386,N_19052,N_19132);
and U19387 (N_19387,N_19118,N_19129);
xor U19388 (N_19388,N_19161,N_19069);
and U19389 (N_19389,N_19184,N_19167);
or U19390 (N_19390,N_19195,N_19035);
and U19391 (N_19391,N_19109,N_19089);
or U19392 (N_19392,N_19177,N_19152);
xnor U19393 (N_19393,N_19195,N_19125);
nor U19394 (N_19394,N_19157,N_19116);
nor U19395 (N_19395,N_19060,N_19057);
or U19396 (N_19396,N_19148,N_19189);
or U19397 (N_19397,N_19154,N_19088);
xor U19398 (N_19398,N_19195,N_19072);
and U19399 (N_19399,N_19161,N_19158);
nor U19400 (N_19400,N_19374,N_19352);
or U19401 (N_19401,N_19387,N_19207);
nand U19402 (N_19402,N_19296,N_19355);
xor U19403 (N_19403,N_19278,N_19293);
nor U19404 (N_19404,N_19279,N_19329);
nor U19405 (N_19405,N_19258,N_19347);
nand U19406 (N_19406,N_19328,N_19336);
xnor U19407 (N_19407,N_19200,N_19262);
xnor U19408 (N_19408,N_19338,N_19227);
nand U19409 (N_19409,N_19234,N_19375);
nor U19410 (N_19410,N_19259,N_19340);
or U19411 (N_19411,N_19344,N_19333);
or U19412 (N_19412,N_19245,N_19252);
xnor U19413 (N_19413,N_19384,N_19261);
or U19414 (N_19414,N_19358,N_19208);
and U19415 (N_19415,N_19230,N_19270);
xor U19416 (N_19416,N_19289,N_19327);
nand U19417 (N_19417,N_19305,N_19390);
and U19418 (N_19418,N_19210,N_19345);
and U19419 (N_19419,N_19257,N_19382);
nand U19420 (N_19420,N_19370,N_19330);
xor U19421 (N_19421,N_19398,N_19343);
or U19422 (N_19422,N_19319,N_19211);
nand U19423 (N_19423,N_19348,N_19395);
nand U19424 (N_19424,N_19284,N_19315);
nor U19425 (N_19425,N_19251,N_19353);
and U19426 (N_19426,N_19307,N_19389);
nor U19427 (N_19427,N_19321,N_19372);
nand U19428 (N_19428,N_19268,N_19380);
or U19429 (N_19429,N_19265,N_19255);
nor U19430 (N_19430,N_19334,N_19264);
and U19431 (N_19431,N_19312,N_19383);
and U19432 (N_19432,N_19331,N_19341);
and U19433 (N_19433,N_19373,N_19256);
and U19434 (N_19434,N_19213,N_19297);
or U19435 (N_19435,N_19285,N_19359);
xor U19436 (N_19436,N_19295,N_19298);
nand U19437 (N_19437,N_19217,N_19274);
or U19438 (N_19438,N_19364,N_19287);
xor U19439 (N_19439,N_19392,N_19367);
nor U19440 (N_19440,N_19209,N_19394);
nand U19441 (N_19441,N_19281,N_19244);
or U19442 (N_19442,N_19228,N_19303);
nor U19443 (N_19443,N_19299,N_19231);
or U19444 (N_19444,N_19324,N_19369);
or U19445 (N_19445,N_19366,N_19306);
or U19446 (N_19446,N_19317,N_19335);
nor U19447 (N_19447,N_19277,N_19361);
or U19448 (N_19448,N_19325,N_19322);
xor U19449 (N_19449,N_19221,N_19246);
xor U19450 (N_19450,N_19357,N_19396);
nor U19451 (N_19451,N_19349,N_19204);
nand U19452 (N_19452,N_19350,N_19243);
xor U19453 (N_19453,N_19332,N_19381);
xor U19454 (N_19454,N_19313,N_19288);
or U19455 (N_19455,N_19360,N_19272);
and U19456 (N_19456,N_19388,N_19206);
nor U19457 (N_19457,N_19229,N_19290);
xnor U19458 (N_19458,N_19385,N_19393);
xor U19459 (N_19459,N_19283,N_19362);
nor U19460 (N_19460,N_19233,N_19275);
nor U19461 (N_19461,N_19269,N_19391);
xnor U19462 (N_19462,N_19236,N_19235);
nor U19463 (N_19463,N_19267,N_19376);
xnor U19464 (N_19464,N_19371,N_19240);
xnor U19465 (N_19465,N_19318,N_19316);
and U19466 (N_19466,N_19226,N_19308);
nand U19467 (N_19467,N_19377,N_19310);
or U19468 (N_19468,N_19280,N_19212);
nand U19469 (N_19469,N_19266,N_19368);
nor U19470 (N_19470,N_19271,N_19351);
nand U19471 (N_19471,N_19379,N_19238);
nand U19472 (N_19472,N_19309,N_19320);
or U19473 (N_19473,N_19237,N_19248);
or U19474 (N_19474,N_19304,N_19339);
xor U19475 (N_19475,N_19253,N_19249);
xnor U19476 (N_19476,N_19242,N_19314);
xnor U19477 (N_19477,N_19326,N_19223);
xnor U19478 (N_19478,N_19337,N_19386);
nor U19479 (N_19479,N_19276,N_19291);
or U19480 (N_19480,N_19250,N_19216);
or U19481 (N_19481,N_19202,N_19205);
and U19482 (N_19482,N_19346,N_19203);
nor U19483 (N_19483,N_19241,N_19363);
nor U19484 (N_19484,N_19219,N_19214);
nor U19485 (N_19485,N_19286,N_19292);
nand U19486 (N_19486,N_19378,N_19311);
nand U19487 (N_19487,N_19397,N_19273);
nand U19488 (N_19488,N_19302,N_19294);
nor U19489 (N_19489,N_19263,N_19224);
nand U19490 (N_19490,N_19239,N_19356);
and U19491 (N_19491,N_19323,N_19399);
nand U19492 (N_19492,N_19201,N_19254);
nand U19493 (N_19493,N_19220,N_19222);
and U19494 (N_19494,N_19342,N_19365);
or U19495 (N_19495,N_19301,N_19218);
or U19496 (N_19496,N_19232,N_19260);
xnor U19497 (N_19497,N_19247,N_19215);
and U19498 (N_19498,N_19354,N_19300);
nand U19499 (N_19499,N_19225,N_19282);
nand U19500 (N_19500,N_19342,N_19238);
nand U19501 (N_19501,N_19217,N_19315);
xor U19502 (N_19502,N_19372,N_19337);
xor U19503 (N_19503,N_19290,N_19351);
nor U19504 (N_19504,N_19371,N_19360);
or U19505 (N_19505,N_19357,N_19370);
and U19506 (N_19506,N_19305,N_19294);
nor U19507 (N_19507,N_19225,N_19384);
and U19508 (N_19508,N_19318,N_19202);
nand U19509 (N_19509,N_19311,N_19359);
nand U19510 (N_19510,N_19220,N_19273);
or U19511 (N_19511,N_19271,N_19326);
and U19512 (N_19512,N_19306,N_19263);
or U19513 (N_19513,N_19344,N_19280);
and U19514 (N_19514,N_19344,N_19346);
nand U19515 (N_19515,N_19382,N_19254);
nand U19516 (N_19516,N_19388,N_19348);
xor U19517 (N_19517,N_19276,N_19252);
or U19518 (N_19518,N_19201,N_19345);
and U19519 (N_19519,N_19231,N_19369);
nor U19520 (N_19520,N_19217,N_19316);
nand U19521 (N_19521,N_19310,N_19230);
and U19522 (N_19522,N_19281,N_19337);
nand U19523 (N_19523,N_19276,N_19280);
xor U19524 (N_19524,N_19313,N_19251);
or U19525 (N_19525,N_19353,N_19318);
xnor U19526 (N_19526,N_19330,N_19293);
nor U19527 (N_19527,N_19302,N_19396);
or U19528 (N_19528,N_19313,N_19341);
or U19529 (N_19529,N_19260,N_19395);
nand U19530 (N_19530,N_19347,N_19286);
nand U19531 (N_19531,N_19320,N_19351);
nand U19532 (N_19532,N_19272,N_19309);
and U19533 (N_19533,N_19387,N_19234);
and U19534 (N_19534,N_19261,N_19359);
nand U19535 (N_19535,N_19370,N_19251);
or U19536 (N_19536,N_19270,N_19302);
nor U19537 (N_19537,N_19253,N_19272);
or U19538 (N_19538,N_19347,N_19226);
nand U19539 (N_19539,N_19349,N_19387);
and U19540 (N_19540,N_19265,N_19215);
or U19541 (N_19541,N_19341,N_19269);
or U19542 (N_19542,N_19379,N_19389);
nand U19543 (N_19543,N_19343,N_19395);
nand U19544 (N_19544,N_19354,N_19371);
xor U19545 (N_19545,N_19321,N_19259);
nand U19546 (N_19546,N_19256,N_19272);
or U19547 (N_19547,N_19269,N_19305);
and U19548 (N_19548,N_19347,N_19266);
or U19549 (N_19549,N_19353,N_19283);
and U19550 (N_19550,N_19386,N_19370);
and U19551 (N_19551,N_19293,N_19303);
and U19552 (N_19552,N_19351,N_19384);
nor U19553 (N_19553,N_19267,N_19370);
xor U19554 (N_19554,N_19365,N_19374);
nor U19555 (N_19555,N_19344,N_19381);
nand U19556 (N_19556,N_19282,N_19246);
nand U19557 (N_19557,N_19310,N_19256);
nand U19558 (N_19558,N_19266,N_19205);
nor U19559 (N_19559,N_19275,N_19264);
or U19560 (N_19560,N_19386,N_19275);
xnor U19561 (N_19561,N_19283,N_19251);
and U19562 (N_19562,N_19299,N_19346);
and U19563 (N_19563,N_19249,N_19275);
nand U19564 (N_19564,N_19269,N_19219);
or U19565 (N_19565,N_19318,N_19395);
nand U19566 (N_19566,N_19341,N_19280);
and U19567 (N_19567,N_19368,N_19356);
nand U19568 (N_19568,N_19313,N_19225);
xnor U19569 (N_19569,N_19364,N_19279);
nor U19570 (N_19570,N_19244,N_19335);
or U19571 (N_19571,N_19342,N_19205);
nand U19572 (N_19572,N_19348,N_19303);
xnor U19573 (N_19573,N_19322,N_19265);
and U19574 (N_19574,N_19331,N_19241);
nand U19575 (N_19575,N_19383,N_19381);
xor U19576 (N_19576,N_19378,N_19296);
nor U19577 (N_19577,N_19371,N_19220);
nor U19578 (N_19578,N_19310,N_19354);
xor U19579 (N_19579,N_19224,N_19328);
and U19580 (N_19580,N_19302,N_19359);
or U19581 (N_19581,N_19340,N_19372);
and U19582 (N_19582,N_19322,N_19399);
xnor U19583 (N_19583,N_19314,N_19207);
xnor U19584 (N_19584,N_19338,N_19243);
nor U19585 (N_19585,N_19237,N_19249);
nor U19586 (N_19586,N_19355,N_19231);
xnor U19587 (N_19587,N_19270,N_19339);
or U19588 (N_19588,N_19360,N_19212);
nor U19589 (N_19589,N_19280,N_19215);
and U19590 (N_19590,N_19369,N_19367);
nor U19591 (N_19591,N_19220,N_19381);
or U19592 (N_19592,N_19390,N_19323);
and U19593 (N_19593,N_19220,N_19262);
xnor U19594 (N_19594,N_19216,N_19314);
xnor U19595 (N_19595,N_19238,N_19358);
or U19596 (N_19596,N_19376,N_19226);
nand U19597 (N_19597,N_19303,N_19385);
nand U19598 (N_19598,N_19250,N_19387);
and U19599 (N_19599,N_19222,N_19304);
xor U19600 (N_19600,N_19509,N_19428);
and U19601 (N_19601,N_19522,N_19514);
and U19602 (N_19602,N_19403,N_19532);
or U19603 (N_19603,N_19431,N_19411);
xnor U19604 (N_19604,N_19422,N_19478);
and U19605 (N_19605,N_19499,N_19437);
nor U19606 (N_19606,N_19423,N_19473);
and U19607 (N_19607,N_19495,N_19408);
and U19608 (N_19608,N_19545,N_19414);
or U19609 (N_19609,N_19407,N_19584);
or U19610 (N_19610,N_19511,N_19435);
nor U19611 (N_19611,N_19531,N_19488);
and U19612 (N_19612,N_19474,N_19560);
and U19613 (N_19613,N_19554,N_19452);
xor U19614 (N_19614,N_19525,N_19550);
and U19615 (N_19615,N_19445,N_19508);
nand U19616 (N_19616,N_19472,N_19464);
and U19617 (N_19617,N_19536,N_19589);
or U19618 (N_19618,N_19406,N_19461);
xor U19619 (N_19619,N_19573,N_19420);
nor U19620 (N_19620,N_19417,N_19564);
nor U19621 (N_19621,N_19555,N_19440);
nand U19622 (N_19622,N_19524,N_19418);
nor U19623 (N_19623,N_19505,N_19574);
nor U19624 (N_19624,N_19521,N_19503);
xnor U19625 (N_19625,N_19570,N_19439);
nand U19626 (N_19626,N_19492,N_19512);
nor U19627 (N_19627,N_19542,N_19463);
or U19628 (N_19628,N_19551,N_19527);
nor U19629 (N_19629,N_19426,N_19470);
or U19630 (N_19630,N_19544,N_19530);
or U19631 (N_19631,N_19599,N_19424);
and U19632 (N_19632,N_19547,N_19427);
nand U19633 (N_19633,N_19425,N_19562);
nand U19634 (N_19634,N_19490,N_19475);
or U19635 (N_19635,N_19563,N_19583);
nand U19636 (N_19636,N_19409,N_19523);
and U19637 (N_19637,N_19540,N_19448);
nand U19638 (N_19638,N_19400,N_19467);
nor U19639 (N_19639,N_19569,N_19405);
xnor U19640 (N_19640,N_19487,N_19526);
nand U19641 (N_19641,N_19486,N_19543);
xnor U19642 (N_19642,N_19450,N_19453);
and U19643 (N_19643,N_19535,N_19520);
xor U19644 (N_19644,N_19455,N_19594);
nand U19645 (N_19645,N_19410,N_19501);
xnor U19646 (N_19646,N_19558,N_19548);
or U19647 (N_19647,N_19586,N_19596);
nand U19648 (N_19648,N_19517,N_19592);
or U19649 (N_19649,N_19483,N_19556);
nor U19650 (N_19650,N_19581,N_19507);
and U19651 (N_19651,N_19539,N_19568);
nand U19652 (N_19652,N_19491,N_19485);
and U19653 (N_19653,N_19580,N_19438);
nor U19654 (N_19654,N_19595,N_19434);
or U19655 (N_19655,N_19585,N_19447);
and U19656 (N_19656,N_19582,N_19587);
xnor U19657 (N_19657,N_19515,N_19413);
or U19658 (N_19658,N_19458,N_19510);
xnor U19659 (N_19659,N_19518,N_19466);
nand U19660 (N_19660,N_19572,N_19469);
nor U19661 (N_19661,N_19482,N_19559);
nor U19662 (N_19662,N_19496,N_19541);
nand U19663 (N_19663,N_19549,N_19597);
nor U19664 (N_19664,N_19421,N_19567);
and U19665 (N_19665,N_19444,N_19449);
and U19666 (N_19666,N_19578,N_19519);
nand U19667 (N_19667,N_19529,N_19500);
and U19668 (N_19668,N_19591,N_19462);
xnor U19669 (N_19669,N_19576,N_19552);
nor U19670 (N_19670,N_19502,N_19489);
nand U19671 (N_19671,N_19534,N_19593);
nand U19672 (N_19672,N_19442,N_19415);
nor U19673 (N_19673,N_19471,N_19579);
and U19674 (N_19674,N_19430,N_19484);
and U19675 (N_19675,N_19504,N_19429);
or U19676 (N_19676,N_19433,N_19575);
or U19677 (N_19677,N_19533,N_19459);
xnor U19678 (N_19678,N_19506,N_19498);
or U19679 (N_19679,N_19598,N_19401);
nor U19680 (N_19680,N_19497,N_19553);
nand U19681 (N_19681,N_19476,N_19479);
and U19682 (N_19682,N_19561,N_19457);
or U19683 (N_19683,N_19432,N_19404);
xor U19684 (N_19684,N_19481,N_19454);
or U19685 (N_19685,N_19460,N_19565);
nor U19686 (N_19686,N_19516,N_19557);
nand U19687 (N_19687,N_19537,N_19546);
nor U19688 (N_19688,N_19477,N_19451);
xor U19689 (N_19689,N_19588,N_19456);
nor U19690 (N_19690,N_19566,N_19446);
xnor U19691 (N_19691,N_19468,N_19402);
xnor U19692 (N_19692,N_19571,N_19493);
or U19693 (N_19693,N_19480,N_19494);
xnor U19694 (N_19694,N_19528,N_19538);
or U19695 (N_19695,N_19513,N_19577);
nand U19696 (N_19696,N_19419,N_19443);
xnor U19697 (N_19697,N_19412,N_19441);
nand U19698 (N_19698,N_19590,N_19465);
or U19699 (N_19699,N_19416,N_19436);
xor U19700 (N_19700,N_19436,N_19555);
xor U19701 (N_19701,N_19591,N_19561);
nor U19702 (N_19702,N_19595,N_19573);
or U19703 (N_19703,N_19412,N_19541);
xnor U19704 (N_19704,N_19539,N_19563);
nand U19705 (N_19705,N_19491,N_19569);
nor U19706 (N_19706,N_19566,N_19407);
nand U19707 (N_19707,N_19425,N_19568);
and U19708 (N_19708,N_19437,N_19578);
or U19709 (N_19709,N_19522,N_19504);
or U19710 (N_19710,N_19407,N_19499);
nand U19711 (N_19711,N_19479,N_19484);
nor U19712 (N_19712,N_19578,N_19561);
nand U19713 (N_19713,N_19531,N_19573);
xnor U19714 (N_19714,N_19510,N_19560);
nor U19715 (N_19715,N_19455,N_19595);
nor U19716 (N_19716,N_19592,N_19501);
nor U19717 (N_19717,N_19515,N_19494);
nand U19718 (N_19718,N_19526,N_19594);
xor U19719 (N_19719,N_19422,N_19425);
nor U19720 (N_19720,N_19447,N_19559);
or U19721 (N_19721,N_19510,N_19528);
nand U19722 (N_19722,N_19556,N_19528);
nor U19723 (N_19723,N_19455,N_19515);
xor U19724 (N_19724,N_19424,N_19403);
nand U19725 (N_19725,N_19465,N_19447);
and U19726 (N_19726,N_19480,N_19579);
and U19727 (N_19727,N_19525,N_19459);
nand U19728 (N_19728,N_19540,N_19472);
or U19729 (N_19729,N_19504,N_19413);
xor U19730 (N_19730,N_19472,N_19521);
or U19731 (N_19731,N_19564,N_19500);
xor U19732 (N_19732,N_19490,N_19594);
and U19733 (N_19733,N_19515,N_19526);
nor U19734 (N_19734,N_19551,N_19462);
and U19735 (N_19735,N_19400,N_19437);
xnor U19736 (N_19736,N_19403,N_19490);
xnor U19737 (N_19737,N_19580,N_19553);
or U19738 (N_19738,N_19589,N_19588);
or U19739 (N_19739,N_19489,N_19412);
nand U19740 (N_19740,N_19441,N_19532);
or U19741 (N_19741,N_19526,N_19452);
or U19742 (N_19742,N_19550,N_19572);
or U19743 (N_19743,N_19443,N_19517);
or U19744 (N_19744,N_19428,N_19407);
xnor U19745 (N_19745,N_19460,N_19424);
or U19746 (N_19746,N_19428,N_19422);
or U19747 (N_19747,N_19555,N_19593);
nor U19748 (N_19748,N_19540,N_19572);
or U19749 (N_19749,N_19593,N_19536);
nor U19750 (N_19750,N_19476,N_19501);
xnor U19751 (N_19751,N_19468,N_19571);
or U19752 (N_19752,N_19513,N_19593);
xnor U19753 (N_19753,N_19515,N_19514);
xnor U19754 (N_19754,N_19584,N_19595);
nor U19755 (N_19755,N_19447,N_19581);
and U19756 (N_19756,N_19487,N_19535);
nand U19757 (N_19757,N_19542,N_19484);
nor U19758 (N_19758,N_19488,N_19466);
xnor U19759 (N_19759,N_19532,N_19420);
nand U19760 (N_19760,N_19428,N_19432);
and U19761 (N_19761,N_19559,N_19578);
nand U19762 (N_19762,N_19421,N_19517);
nor U19763 (N_19763,N_19443,N_19400);
xnor U19764 (N_19764,N_19562,N_19557);
or U19765 (N_19765,N_19460,N_19518);
or U19766 (N_19766,N_19538,N_19429);
nor U19767 (N_19767,N_19470,N_19588);
or U19768 (N_19768,N_19598,N_19527);
nor U19769 (N_19769,N_19446,N_19554);
and U19770 (N_19770,N_19558,N_19508);
xnor U19771 (N_19771,N_19516,N_19546);
or U19772 (N_19772,N_19552,N_19550);
or U19773 (N_19773,N_19534,N_19528);
nor U19774 (N_19774,N_19543,N_19588);
nand U19775 (N_19775,N_19534,N_19443);
xnor U19776 (N_19776,N_19569,N_19594);
nand U19777 (N_19777,N_19403,N_19421);
nand U19778 (N_19778,N_19438,N_19532);
and U19779 (N_19779,N_19541,N_19408);
or U19780 (N_19780,N_19404,N_19434);
nand U19781 (N_19781,N_19403,N_19546);
or U19782 (N_19782,N_19416,N_19550);
xnor U19783 (N_19783,N_19599,N_19480);
nand U19784 (N_19784,N_19439,N_19527);
and U19785 (N_19785,N_19503,N_19554);
and U19786 (N_19786,N_19506,N_19479);
or U19787 (N_19787,N_19586,N_19583);
and U19788 (N_19788,N_19438,N_19423);
and U19789 (N_19789,N_19513,N_19557);
or U19790 (N_19790,N_19598,N_19468);
or U19791 (N_19791,N_19456,N_19560);
xor U19792 (N_19792,N_19420,N_19554);
nor U19793 (N_19793,N_19484,N_19549);
nand U19794 (N_19794,N_19537,N_19488);
xor U19795 (N_19795,N_19447,N_19438);
xnor U19796 (N_19796,N_19490,N_19559);
and U19797 (N_19797,N_19424,N_19489);
and U19798 (N_19798,N_19473,N_19589);
or U19799 (N_19799,N_19540,N_19595);
and U19800 (N_19800,N_19669,N_19712);
xnor U19801 (N_19801,N_19608,N_19652);
nor U19802 (N_19802,N_19675,N_19695);
or U19803 (N_19803,N_19603,N_19690);
xor U19804 (N_19804,N_19676,N_19736);
xnor U19805 (N_19805,N_19672,N_19752);
or U19806 (N_19806,N_19708,N_19729);
and U19807 (N_19807,N_19659,N_19632);
or U19808 (N_19808,N_19778,N_19671);
or U19809 (N_19809,N_19693,N_19795);
nor U19810 (N_19810,N_19788,N_19770);
and U19811 (N_19811,N_19619,N_19750);
and U19812 (N_19812,N_19609,N_19747);
and U19813 (N_19813,N_19614,N_19699);
nand U19814 (N_19814,N_19776,N_19634);
nor U19815 (N_19815,N_19740,N_19687);
nand U19816 (N_19816,N_19626,N_19754);
nand U19817 (N_19817,N_19625,N_19683);
nand U19818 (N_19818,N_19719,N_19660);
nand U19819 (N_19819,N_19611,N_19725);
and U19820 (N_19820,N_19745,N_19735);
xor U19821 (N_19821,N_19791,N_19667);
nand U19822 (N_19822,N_19713,N_19756);
and U19823 (N_19823,N_19668,N_19673);
and U19824 (N_19824,N_19680,N_19782);
xor U19825 (N_19825,N_19615,N_19616);
or U19826 (N_19826,N_19704,N_19786);
or U19827 (N_19827,N_19710,N_19646);
and U19828 (N_19828,N_19686,N_19649);
and U19829 (N_19829,N_19732,N_19685);
xor U19830 (N_19830,N_19694,N_19650);
or U19831 (N_19831,N_19764,N_19620);
xnor U19832 (N_19832,N_19658,N_19692);
nor U19833 (N_19833,N_19792,N_19765);
and U19834 (N_19834,N_19697,N_19600);
and U19835 (N_19835,N_19709,N_19700);
and U19836 (N_19836,N_19630,N_19796);
and U19837 (N_19837,N_19767,N_19636);
and U19838 (N_19838,N_19731,N_19623);
xor U19839 (N_19839,N_19701,N_19703);
nor U19840 (N_19840,N_19793,N_19705);
xor U19841 (N_19841,N_19726,N_19737);
xnor U19842 (N_19842,N_19605,N_19761);
xor U19843 (N_19843,N_19717,N_19664);
and U19844 (N_19844,N_19768,N_19716);
nor U19845 (N_19845,N_19665,N_19787);
xor U19846 (N_19846,N_19612,N_19642);
xnor U19847 (N_19847,N_19784,N_19651);
xor U19848 (N_19848,N_19629,N_19627);
nand U19849 (N_19849,N_19728,N_19655);
and U19850 (N_19850,N_19621,N_19618);
nand U19851 (N_19851,N_19780,N_19774);
or U19852 (N_19852,N_19617,N_19633);
or U19853 (N_19853,N_19744,N_19763);
nor U19854 (N_19854,N_19643,N_19715);
and U19855 (N_19855,N_19679,N_19753);
and U19856 (N_19856,N_19734,N_19641);
or U19857 (N_19857,N_19730,N_19771);
nor U19858 (N_19858,N_19751,N_19727);
nand U19859 (N_19859,N_19714,N_19773);
nor U19860 (N_19860,N_19698,N_19769);
or U19861 (N_19861,N_19601,N_19631);
xnor U19862 (N_19862,N_19706,N_19762);
xor U19863 (N_19863,N_19613,N_19758);
nor U19864 (N_19864,N_19648,N_19647);
nand U19865 (N_19865,N_19640,N_19720);
and U19866 (N_19866,N_19749,N_19689);
nand U19867 (N_19867,N_19657,N_19742);
nor U19868 (N_19868,N_19653,N_19775);
or U19869 (N_19869,N_19739,N_19637);
nor U19870 (N_19870,N_19746,N_19661);
xnor U19871 (N_19871,N_19766,N_19602);
xor U19872 (N_19872,N_19798,N_19663);
xnor U19873 (N_19873,N_19738,N_19645);
nor U19874 (N_19874,N_19783,N_19723);
nor U19875 (N_19875,N_19794,N_19799);
nand U19876 (N_19876,N_19781,N_19722);
xnor U19877 (N_19877,N_19785,N_19654);
or U19878 (N_19878,N_19684,N_19748);
nor U19879 (N_19879,N_19662,N_19718);
and U19880 (N_19880,N_19702,N_19606);
xnor U19881 (N_19881,N_19635,N_19789);
and U19882 (N_19882,N_19682,N_19607);
nor U19883 (N_19883,N_19741,N_19755);
nand U19884 (N_19884,N_19707,N_19677);
or U19885 (N_19885,N_19644,N_19696);
nand U19886 (N_19886,N_19666,N_19674);
and U19887 (N_19887,N_19604,N_19656);
nand U19888 (N_19888,N_19688,N_19757);
or U19889 (N_19889,N_19733,N_19622);
nor U19890 (N_19890,N_19760,N_19790);
xor U19891 (N_19891,N_19678,N_19724);
xnor U19892 (N_19892,N_19638,N_19743);
or U19893 (N_19893,N_19639,N_19691);
nor U19894 (N_19894,N_19721,N_19759);
nor U19895 (N_19895,N_19624,N_19610);
xor U19896 (N_19896,N_19670,N_19777);
xor U19897 (N_19897,N_19779,N_19772);
and U19898 (N_19898,N_19797,N_19681);
nor U19899 (N_19899,N_19628,N_19711);
or U19900 (N_19900,N_19707,N_19690);
or U19901 (N_19901,N_19704,N_19735);
or U19902 (N_19902,N_19659,N_19755);
xor U19903 (N_19903,N_19685,N_19712);
or U19904 (N_19904,N_19700,N_19692);
xor U19905 (N_19905,N_19750,N_19799);
and U19906 (N_19906,N_19781,N_19644);
and U19907 (N_19907,N_19627,N_19769);
and U19908 (N_19908,N_19751,N_19775);
xnor U19909 (N_19909,N_19661,N_19604);
nand U19910 (N_19910,N_19733,N_19678);
xor U19911 (N_19911,N_19698,N_19644);
xnor U19912 (N_19912,N_19623,N_19622);
xor U19913 (N_19913,N_19699,N_19784);
nor U19914 (N_19914,N_19600,N_19641);
and U19915 (N_19915,N_19785,N_19773);
nor U19916 (N_19916,N_19609,N_19632);
xor U19917 (N_19917,N_19655,N_19698);
xnor U19918 (N_19918,N_19607,N_19672);
and U19919 (N_19919,N_19722,N_19715);
nand U19920 (N_19920,N_19674,N_19796);
or U19921 (N_19921,N_19757,N_19746);
nor U19922 (N_19922,N_19613,N_19699);
or U19923 (N_19923,N_19602,N_19715);
and U19924 (N_19924,N_19690,N_19664);
nand U19925 (N_19925,N_19602,N_19655);
xnor U19926 (N_19926,N_19672,N_19780);
or U19927 (N_19927,N_19793,N_19736);
and U19928 (N_19928,N_19727,N_19613);
nand U19929 (N_19929,N_19665,N_19653);
nor U19930 (N_19930,N_19746,N_19762);
nor U19931 (N_19931,N_19766,N_19714);
nor U19932 (N_19932,N_19623,N_19722);
or U19933 (N_19933,N_19714,N_19795);
and U19934 (N_19934,N_19707,N_19762);
nand U19935 (N_19935,N_19615,N_19710);
or U19936 (N_19936,N_19712,N_19766);
or U19937 (N_19937,N_19787,N_19678);
nand U19938 (N_19938,N_19691,N_19757);
xnor U19939 (N_19939,N_19638,N_19688);
nor U19940 (N_19940,N_19738,N_19695);
nand U19941 (N_19941,N_19619,N_19691);
and U19942 (N_19942,N_19791,N_19619);
and U19943 (N_19943,N_19631,N_19718);
or U19944 (N_19944,N_19719,N_19723);
nand U19945 (N_19945,N_19790,N_19674);
nand U19946 (N_19946,N_19704,N_19764);
xnor U19947 (N_19947,N_19610,N_19749);
xnor U19948 (N_19948,N_19652,N_19763);
nand U19949 (N_19949,N_19646,N_19732);
and U19950 (N_19950,N_19714,N_19605);
nor U19951 (N_19951,N_19641,N_19605);
nor U19952 (N_19952,N_19698,N_19637);
nor U19953 (N_19953,N_19620,N_19740);
or U19954 (N_19954,N_19776,N_19740);
xnor U19955 (N_19955,N_19770,N_19622);
nor U19956 (N_19956,N_19726,N_19796);
xnor U19957 (N_19957,N_19777,N_19606);
nand U19958 (N_19958,N_19728,N_19674);
nor U19959 (N_19959,N_19691,N_19697);
and U19960 (N_19960,N_19743,N_19629);
xnor U19961 (N_19961,N_19654,N_19770);
nor U19962 (N_19962,N_19728,N_19621);
or U19963 (N_19963,N_19704,N_19699);
and U19964 (N_19964,N_19644,N_19743);
and U19965 (N_19965,N_19618,N_19667);
xor U19966 (N_19966,N_19700,N_19710);
nand U19967 (N_19967,N_19768,N_19775);
xor U19968 (N_19968,N_19616,N_19632);
nor U19969 (N_19969,N_19659,N_19717);
xnor U19970 (N_19970,N_19670,N_19757);
nand U19971 (N_19971,N_19614,N_19780);
nor U19972 (N_19972,N_19776,N_19652);
nand U19973 (N_19973,N_19672,N_19745);
nand U19974 (N_19974,N_19611,N_19798);
and U19975 (N_19975,N_19725,N_19626);
and U19976 (N_19976,N_19732,N_19769);
nor U19977 (N_19977,N_19658,N_19729);
and U19978 (N_19978,N_19767,N_19694);
or U19979 (N_19979,N_19663,N_19740);
or U19980 (N_19980,N_19692,N_19606);
xor U19981 (N_19981,N_19749,N_19677);
xnor U19982 (N_19982,N_19693,N_19789);
and U19983 (N_19983,N_19664,N_19679);
or U19984 (N_19984,N_19655,N_19689);
nand U19985 (N_19985,N_19610,N_19746);
xor U19986 (N_19986,N_19744,N_19688);
or U19987 (N_19987,N_19717,N_19727);
nor U19988 (N_19988,N_19661,N_19750);
and U19989 (N_19989,N_19642,N_19693);
nand U19990 (N_19990,N_19601,N_19692);
nand U19991 (N_19991,N_19748,N_19642);
xor U19992 (N_19992,N_19771,N_19608);
nand U19993 (N_19993,N_19744,N_19669);
nand U19994 (N_19994,N_19692,N_19627);
and U19995 (N_19995,N_19633,N_19750);
xnor U19996 (N_19996,N_19798,N_19704);
nand U19997 (N_19997,N_19767,N_19639);
or U19998 (N_19998,N_19639,N_19765);
or U19999 (N_19999,N_19729,N_19692);
or UO_0 (O_0,N_19938,N_19994);
nand UO_1 (O_1,N_19879,N_19977);
nor UO_2 (O_2,N_19964,N_19970);
or UO_3 (O_3,N_19871,N_19881);
xor UO_4 (O_4,N_19842,N_19894);
or UO_5 (O_5,N_19914,N_19951);
and UO_6 (O_6,N_19957,N_19861);
and UO_7 (O_7,N_19857,N_19965);
xnor UO_8 (O_8,N_19876,N_19932);
nor UO_9 (O_9,N_19888,N_19893);
nand UO_10 (O_10,N_19972,N_19868);
nor UO_11 (O_11,N_19926,N_19940);
xnor UO_12 (O_12,N_19808,N_19802);
xor UO_13 (O_13,N_19824,N_19815);
nand UO_14 (O_14,N_19905,N_19930);
xnor UO_15 (O_15,N_19838,N_19955);
nand UO_16 (O_16,N_19903,N_19807);
nor UO_17 (O_17,N_19856,N_19919);
xor UO_18 (O_18,N_19963,N_19952);
and UO_19 (O_19,N_19939,N_19862);
and UO_20 (O_20,N_19877,N_19947);
nand UO_21 (O_21,N_19869,N_19835);
nand UO_22 (O_22,N_19916,N_19944);
or UO_23 (O_23,N_19969,N_19910);
and UO_24 (O_24,N_19827,N_19904);
xnor UO_25 (O_25,N_19925,N_19943);
and UO_26 (O_26,N_19899,N_19968);
nor UO_27 (O_27,N_19949,N_19883);
nand UO_28 (O_28,N_19967,N_19975);
nand UO_29 (O_29,N_19817,N_19870);
nor UO_30 (O_30,N_19836,N_19966);
xor UO_31 (O_31,N_19954,N_19821);
nand UO_32 (O_32,N_19831,N_19937);
xnor UO_33 (O_33,N_19995,N_19934);
nor UO_34 (O_34,N_19982,N_19875);
or UO_35 (O_35,N_19855,N_19991);
xnor UO_36 (O_36,N_19896,N_19889);
nor UO_37 (O_37,N_19872,N_19851);
or UO_38 (O_38,N_19895,N_19850);
nand UO_39 (O_39,N_19931,N_19958);
or UO_40 (O_40,N_19805,N_19946);
and UO_41 (O_41,N_19985,N_19843);
and UO_42 (O_42,N_19920,N_19941);
xor UO_43 (O_43,N_19839,N_19988);
nor UO_44 (O_44,N_19880,N_19921);
nand UO_45 (O_45,N_19810,N_19822);
xor UO_46 (O_46,N_19874,N_19885);
nor UO_47 (O_47,N_19993,N_19961);
xnor UO_48 (O_48,N_19986,N_19834);
nor UO_49 (O_49,N_19847,N_19812);
nand UO_50 (O_50,N_19829,N_19898);
nand UO_51 (O_51,N_19933,N_19927);
xnor UO_52 (O_52,N_19854,N_19953);
xnor UO_53 (O_53,N_19814,N_19803);
xor UO_54 (O_54,N_19917,N_19990);
nor UO_55 (O_55,N_19902,N_19859);
xnor UO_56 (O_56,N_19983,N_19820);
xor UO_57 (O_57,N_19992,N_19979);
xnor UO_58 (O_58,N_19973,N_19882);
nand UO_59 (O_59,N_19866,N_19924);
xnor UO_60 (O_60,N_19886,N_19962);
and UO_61 (O_61,N_19981,N_19813);
and UO_62 (O_62,N_19984,N_19950);
and UO_63 (O_63,N_19945,N_19897);
xnor UO_64 (O_64,N_19878,N_19922);
or UO_65 (O_65,N_19978,N_19907);
nor UO_66 (O_66,N_19833,N_19828);
nand UO_67 (O_67,N_19849,N_19852);
nand UO_68 (O_68,N_19891,N_19804);
nand UO_69 (O_69,N_19832,N_19935);
and UO_70 (O_70,N_19867,N_19809);
nor UO_71 (O_71,N_19976,N_19928);
nor UO_72 (O_72,N_19900,N_19890);
or UO_73 (O_73,N_19913,N_19818);
and UO_74 (O_74,N_19909,N_19929);
nand UO_75 (O_75,N_19942,N_19841);
nand UO_76 (O_76,N_19840,N_19918);
and UO_77 (O_77,N_19996,N_19860);
xor UO_78 (O_78,N_19892,N_19845);
xnor UO_79 (O_79,N_19956,N_19846);
nor UO_80 (O_80,N_19819,N_19873);
nor UO_81 (O_81,N_19936,N_19800);
or UO_82 (O_82,N_19884,N_19948);
or UO_83 (O_83,N_19823,N_19901);
nand UO_84 (O_84,N_19806,N_19911);
and UO_85 (O_85,N_19826,N_19997);
or UO_86 (O_86,N_19908,N_19960);
or UO_87 (O_87,N_19853,N_19864);
xor UO_88 (O_88,N_19844,N_19863);
xnor UO_89 (O_89,N_19974,N_19906);
or UO_90 (O_90,N_19825,N_19816);
nand UO_91 (O_91,N_19987,N_19971);
xnor UO_92 (O_92,N_19801,N_19989);
nand UO_93 (O_93,N_19998,N_19959);
and UO_94 (O_94,N_19865,N_19923);
and UO_95 (O_95,N_19837,N_19915);
or UO_96 (O_96,N_19980,N_19912);
xor UO_97 (O_97,N_19848,N_19887);
or UO_98 (O_98,N_19830,N_19811);
and UO_99 (O_99,N_19999,N_19858);
nor UO_100 (O_100,N_19859,N_19942);
or UO_101 (O_101,N_19889,N_19876);
nand UO_102 (O_102,N_19962,N_19814);
and UO_103 (O_103,N_19847,N_19988);
nand UO_104 (O_104,N_19977,N_19815);
nand UO_105 (O_105,N_19944,N_19950);
nor UO_106 (O_106,N_19889,N_19823);
or UO_107 (O_107,N_19860,N_19937);
or UO_108 (O_108,N_19887,N_19947);
and UO_109 (O_109,N_19979,N_19802);
nor UO_110 (O_110,N_19894,N_19809);
xor UO_111 (O_111,N_19840,N_19824);
nor UO_112 (O_112,N_19898,N_19945);
and UO_113 (O_113,N_19993,N_19836);
nor UO_114 (O_114,N_19919,N_19842);
and UO_115 (O_115,N_19815,N_19833);
nand UO_116 (O_116,N_19921,N_19991);
and UO_117 (O_117,N_19981,N_19844);
nand UO_118 (O_118,N_19978,N_19949);
nor UO_119 (O_119,N_19931,N_19913);
or UO_120 (O_120,N_19829,N_19990);
xor UO_121 (O_121,N_19966,N_19976);
nand UO_122 (O_122,N_19832,N_19870);
nand UO_123 (O_123,N_19953,N_19946);
and UO_124 (O_124,N_19858,N_19834);
nor UO_125 (O_125,N_19820,N_19951);
nand UO_126 (O_126,N_19819,N_19845);
xnor UO_127 (O_127,N_19805,N_19827);
or UO_128 (O_128,N_19922,N_19944);
xor UO_129 (O_129,N_19932,N_19860);
and UO_130 (O_130,N_19999,N_19832);
and UO_131 (O_131,N_19947,N_19898);
xor UO_132 (O_132,N_19819,N_19829);
xnor UO_133 (O_133,N_19851,N_19892);
nand UO_134 (O_134,N_19988,N_19865);
nor UO_135 (O_135,N_19971,N_19956);
or UO_136 (O_136,N_19851,N_19978);
and UO_137 (O_137,N_19876,N_19922);
xor UO_138 (O_138,N_19940,N_19942);
nor UO_139 (O_139,N_19863,N_19813);
or UO_140 (O_140,N_19949,N_19943);
or UO_141 (O_141,N_19868,N_19855);
nand UO_142 (O_142,N_19819,N_19965);
or UO_143 (O_143,N_19889,N_19884);
nor UO_144 (O_144,N_19976,N_19952);
or UO_145 (O_145,N_19805,N_19957);
and UO_146 (O_146,N_19829,N_19908);
and UO_147 (O_147,N_19858,N_19889);
or UO_148 (O_148,N_19825,N_19858);
and UO_149 (O_149,N_19939,N_19963);
nand UO_150 (O_150,N_19946,N_19836);
and UO_151 (O_151,N_19844,N_19807);
nor UO_152 (O_152,N_19943,N_19989);
and UO_153 (O_153,N_19831,N_19823);
and UO_154 (O_154,N_19899,N_19994);
xnor UO_155 (O_155,N_19810,N_19963);
or UO_156 (O_156,N_19963,N_19995);
nor UO_157 (O_157,N_19810,N_19988);
nor UO_158 (O_158,N_19976,N_19862);
or UO_159 (O_159,N_19856,N_19949);
xor UO_160 (O_160,N_19804,N_19956);
xor UO_161 (O_161,N_19966,N_19857);
nand UO_162 (O_162,N_19905,N_19900);
xor UO_163 (O_163,N_19983,N_19873);
xor UO_164 (O_164,N_19824,N_19947);
or UO_165 (O_165,N_19867,N_19900);
xnor UO_166 (O_166,N_19825,N_19899);
nor UO_167 (O_167,N_19876,N_19866);
nor UO_168 (O_168,N_19993,N_19877);
xnor UO_169 (O_169,N_19921,N_19884);
nand UO_170 (O_170,N_19852,N_19919);
nor UO_171 (O_171,N_19816,N_19951);
xnor UO_172 (O_172,N_19976,N_19817);
or UO_173 (O_173,N_19865,N_19864);
nand UO_174 (O_174,N_19866,N_19927);
and UO_175 (O_175,N_19869,N_19816);
nor UO_176 (O_176,N_19901,N_19894);
or UO_177 (O_177,N_19953,N_19915);
or UO_178 (O_178,N_19960,N_19923);
nor UO_179 (O_179,N_19950,N_19816);
xor UO_180 (O_180,N_19953,N_19810);
nor UO_181 (O_181,N_19931,N_19915);
nor UO_182 (O_182,N_19812,N_19813);
and UO_183 (O_183,N_19836,N_19923);
nor UO_184 (O_184,N_19956,N_19881);
xnor UO_185 (O_185,N_19811,N_19883);
xnor UO_186 (O_186,N_19875,N_19832);
nor UO_187 (O_187,N_19993,N_19913);
nand UO_188 (O_188,N_19857,N_19879);
nand UO_189 (O_189,N_19840,N_19825);
xor UO_190 (O_190,N_19984,N_19997);
and UO_191 (O_191,N_19966,N_19813);
nor UO_192 (O_192,N_19849,N_19916);
and UO_193 (O_193,N_19918,N_19905);
xor UO_194 (O_194,N_19996,N_19995);
nand UO_195 (O_195,N_19930,N_19845);
and UO_196 (O_196,N_19932,N_19898);
xnor UO_197 (O_197,N_19886,N_19943);
nand UO_198 (O_198,N_19967,N_19979);
or UO_199 (O_199,N_19875,N_19927);
nand UO_200 (O_200,N_19953,N_19950);
or UO_201 (O_201,N_19969,N_19841);
nor UO_202 (O_202,N_19801,N_19965);
nor UO_203 (O_203,N_19880,N_19978);
or UO_204 (O_204,N_19801,N_19802);
nor UO_205 (O_205,N_19837,N_19867);
nor UO_206 (O_206,N_19800,N_19981);
xor UO_207 (O_207,N_19892,N_19935);
or UO_208 (O_208,N_19970,N_19904);
and UO_209 (O_209,N_19982,N_19817);
nor UO_210 (O_210,N_19827,N_19929);
nor UO_211 (O_211,N_19924,N_19947);
nand UO_212 (O_212,N_19945,N_19907);
or UO_213 (O_213,N_19813,N_19874);
nor UO_214 (O_214,N_19814,N_19848);
nand UO_215 (O_215,N_19937,N_19854);
xnor UO_216 (O_216,N_19926,N_19800);
nand UO_217 (O_217,N_19963,N_19898);
or UO_218 (O_218,N_19810,N_19997);
nor UO_219 (O_219,N_19890,N_19897);
xor UO_220 (O_220,N_19838,N_19932);
nor UO_221 (O_221,N_19829,N_19925);
nand UO_222 (O_222,N_19957,N_19997);
xor UO_223 (O_223,N_19945,N_19832);
and UO_224 (O_224,N_19940,N_19801);
nand UO_225 (O_225,N_19918,N_19990);
nor UO_226 (O_226,N_19896,N_19985);
xor UO_227 (O_227,N_19806,N_19838);
nor UO_228 (O_228,N_19899,N_19829);
xnor UO_229 (O_229,N_19861,N_19830);
nand UO_230 (O_230,N_19895,N_19997);
nand UO_231 (O_231,N_19916,N_19812);
nand UO_232 (O_232,N_19864,N_19880);
xor UO_233 (O_233,N_19842,N_19930);
nand UO_234 (O_234,N_19852,N_19801);
nand UO_235 (O_235,N_19974,N_19818);
xor UO_236 (O_236,N_19833,N_19960);
or UO_237 (O_237,N_19944,N_19912);
nand UO_238 (O_238,N_19964,N_19918);
or UO_239 (O_239,N_19929,N_19990);
and UO_240 (O_240,N_19829,N_19927);
nor UO_241 (O_241,N_19880,N_19947);
xnor UO_242 (O_242,N_19981,N_19811);
nand UO_243 (O_243,N_19893,N_19828);
or UO_244 (O_244,N_19950,N_19995);
nor UO_245 (O_245,N_19954,N_19831);
and UO_246 (O_246,N_19893,N_19864);
xor UO_247 (O_247,N_19967,N_19870);
and UO_248 (O_248,N_19869,N_19839);
nor UO_249 (O_249,N_19943,N_19970);
nor UO_250 (O_250,N_19849,N_19902);
and UO_251 (O_251,N_19973,N_19919);
or UO_252 (O_252,N_19930,N_19932);
nor UO_253 (O_253,N_19976,N_19855);
nor UO_254 (O_254,N_19986,N_19989);
nor UO_255 (O_255,N_19849,N_19936);
or UO_256 (O_256,N_19983,N_19889);
nand UO_257 (O_257,N_19932,N_19903);
or UO_258 (O_258,N_19909,N_19910);
or UO_259 (O_259,N_19976,N_19838);
nor UO_260 (O_260,N_19940,N_19900);
xor UO_261 (O_261,N_19946,N_19856);
nor UO_262 (O_262,N_19868,N_19913);
nor UO_263 (O_263,N_19811,N_19813);
nor UO_264 (O_264,N_19969,N_19916);
xnor UO_265 (O_265,N_19867,N_19874);
and UO_266 (O_266,N_19872,N_19860);
nand UO_267 (O_267,N_19828,N_19923);
and UO_268 (O_268,N_19862,N_19872);
nor UO_269 (O_269,N_19897,N_19862);
and UO_270 (O_270,N_19928,N_19881);
xnor UO_271 (O_271,N_19873,N_19852);
and UO_272 (O_272,N_19857,N_19834);
or UO_273 (O_273,N_19870,N_19884);
nand UO_274 (O_274,N_19879,N_19893);
and UO_275 (O_275,N_19936,N_19846);
nand UO_276 (O_276,N_19843,N_19932);
nor UO_277 (O_277,N_19829,N_19980);
nor UO_278 (O_278,N_19881,N_19927);
xor UO_279 (O_279,N_19956,N_19890);
xor UO_280 (O_280,N_19839,N_19981);
xnor UO_281 (O_281,N_19853,N_19811);
or UO_282 (O_282,N_19892,N_19821);
xnor UO_283 (O_283,N_19891,N_19893);
or UO_284 (O_284,N_19901,N_19880);
or UO_285 (O_285,N_19934,N_19966);
or UO_286 (O_286,N_19802,N_19970);
nor UO_287 (O_287,N_19878,N_19945);
nand UO_288 (O_288,N_19811,N_19936);
xor UO_289 (O_289,N_19997,N_19855);
xor UO_290 (O_290,N_19943,N_19926);
nand UO_291 (O_291,N_19844,N_19871);
xnor UO_292 (O_292,N_19924,N_19814);
or UO_293 (O_293,N_19844,N_19984);
nand UO_294 (O_294,N_19892,N_19995);
nor UO_295 (O_295,N_19921,N_19900);
xor UO_296 (O_296,N_19868,N_19906);
or UO_297 (O_297,N_19870,N_19873);
nand UO_298 (O_298,N_19991,N_19913);
nor UO_299 (O_299,N_19905,N_19920);
or UO_300 (O_300,N_19909,N_19912);
nand UO_301 (O_301,N_19938,N_19897);
nor UO_302 (O_302,N_19983,N_19803);
nand UO_303 (O_303,N_19832,N_19857);
or UO_304 (O_304,N_19937,N_19964);
nor UO_305 (O_305,N_19950,N_19992);
nor UO_306 (O_306,N_19900,N_19902);
nor UO_307 (O_307,N_19870,N_19835);
xnor UO_308 (O_308,N_19823,N_19978);
nor UO_309 (O_309,N_19854,N_19843);
and UO_310 (O_310,N_19830,N_19909);
nand UO_311 (O_311,N_19931,N_19952);
or UO_312 (O_312,N_19980,N_19952);
nand UO_313 (O_313,N_19926,N_19990);
nand UO_314 (O_314,N_19907,N_19876);
nand UO_315 (O_315,N_19894,N_19823);
xnor UO_316 (O_316,N_19909,N_19853);
or UO_317 (O_317,N_19848,N_19946);
nand UO_318 (O_318,N_19829,N_19879);
xnor UO_319 (O_319,N_19893,N_19827);
nor UO_320 (O_320,N_19866,N_19881);
and UO_321 (O_321,N_19832,N_19930);
or UO_322 (O_322,N_19857,N_19800);
or UO_323 (O_323,N_19865,N_19905);
xor UO_324 (O_324,N_19942,N_19855);
or UO_325 (O_325,N_19921,N_19913);
and UO_326 (O_326,N_19839,N_19979);
xor UO_327 (O_327,N_19841,N_19819);
xor UO_328 (O_328,N_19827,N_19836);
nor UO_329 (O_329,N_19982,N_19837);
nor UO_330 (O_330,N_19808,N_19845);
xor UO_331 (O_331,N_19905,N_19968);
nor UO_332 (O_332,N_19997,N_19881);
and UO_333 (O_333,N_19818,N_19990);
nor UO_334 (O_334,N_19861,N_19985);
and UO_335 (O_335,N_19859,N_19917);
or UO_336 (O_336,N_19949,N_19952);
and UO_337 (O_337,N_19962,N_19949);
nand UO_338 (O_338,N_19991,N_19849);
nor UO_339 (O_339,N_19828,N_19882);
and UO_340 (O_340,N_19965,N_19917);
or UO_341 (O_341,N_19911,N_19974);
nor UO_342 (O_342,N_19999,N_19984);
xor UO_343 (O_343,N_19967,N_19807);
nor UO_344 (O_344,N_19990,N_19885);
nand UO_345 (O_345,N_19933,N_19802);
nor UO_346 (O_346,N_19847,N_19940);
xor UO_347 (O_347,N_19811,N_19905);
nand UO_348 (O_348,N_19832,N_19932);
nand UO_349 (O_349,N_19908,N_19933);
or UO_350 (O_350,N_19943,N_19947);
nor UO_351 (O_351,N_19877,N_19808);
and UO_352 (O_352,N_19882,N_19870);
and UO_353 (O_353,N_19827,N_19830);
and UO_354 (O_354,N_19898,N_19933);
nand UO_355 (O_355,N_19992,N_19872);
nor UO_356 (O_356,N_19900,N_19948);
or UO_357 (O_357,N_19925,N_19896);
xor UO_358 (O_358,N_19825,N_19866);
nand UO_359 (O_359,N_19965,N_19957);
nand UO_360 (O_360,N_19914,N_19807);
or UO_361 (O_361,N_19879,N_19915);
nand UO_362 (O_362,N_19840,N_19805);
xnor UO_363 (O_363,N_19860,N_19868);
nand UO_364 (O_364,N_19974,N_19840);
and UO_365 (O_365,N_19877,N_19926);
and UO_366 (O_366,N_19916,N_19907);
nor UO_367 (O_367,N_19939,N_19978);
nand UO_368 (O_368,N_19920,N_19865);
and UO_369 (O_369,N_19917,N_19985);
nor UO_370 (O_370,N_19912,N_19925);
nand UO_371 (O_371,N_19888,N_19949);
or UO_372 (O_372,N_19996,N_19857);
and UO_373 (O_373,N_19826,N_19994);
nor UO_374 (O_374,N_19806,N_19959);
nor UO_375 (O_375,N_19952,N_19907);
nor UO_376 (O_376,N_19841,N_19868);
and UO_377 (O_377,N_19998,N_19985);
and UO_378 (O_378,N_19948,N_19834);
xor UO_379 (O_379,N_19808,N_19826);
and UO_380 (O_380,N_19974,N_19912);
nand UO_381 (O_381,N_19962,N_19914);
or UO_382 (O_382,N_19923,N_19937);
or UO_383 (O_383,N_19833,N_19847);
or UO_384 (O_384,N_19816,N_19860);
xor UO_385 (O_385,N_19908,N_19840);
nand UO_386 (O_386,N_19937,N_19960);
or UO_387 (O_387,N_19915,N_19816);
or UO_388 (O_388,N_19949,N_19984);
nand UO_389 (O_389,N_19859,N_19946);
nand UO_390 (O_390,N_19938,N_19964);
xnor UO_391 (O_391,N_19972,N_19844);
nand UO_392 (O_392,N_19908,N_19964);
or UO_393 (O_393,N_19897,N_19803);
xor UO_394 (O_394,N_19943,N_19847);
and UO_395 (O_395,N_19891,N_19976);
or UO_396 (O_396,N_19869,N_19963);
or UO_397 (O_397,N_19841,N_19858);
or UO_398 (O_398,N_19902,N_19824);
and UO_399 (O_399,N_19925,N_19879);
nor UO_400 (O_400,N_19865,N_19845);
and UO_401 (O_401,N_19924,N_19912);
nand UO_402 (O_402,N_19912,N_19973);
nor UO_403 (O_403,N_19853,N_19874);
nor UO_404 (O_404,N_19987,N_19968);
nand UO_405 (O_405,N_19913,N_19992);
nand UO_406 (O_406,N_19932,N_19949);
xnor UO_407 (O_407,N_19861,N_19897);
and UO_408 (O_408,N_19801,N_19868);
and UO_409 (O_409,N_19801,N_19815);
nor UO_410 (O_410,N_19993,N_19940);
or UO_411 (O_411,N_19841,N_19811);
nand UO_412 (O_412,N_19991,N_19863);
xor UO_413 (O_413,N_19932,N_19888);
nand UO_414 (O_414,N_19864,N_19927);
nand UO_415 (O_415,N_19967,N_19989);
and UO_416 (O_416,N_19912,N_19840);
or UO_417 (O_417,N_19969,N_19975);
nor UO_418 (O_418,N_19886,N_19947);
nor UO_419 (O_419,N_19947,N_19981);
nor UO_420 (O_420,N_19949,N_19981);
nor UO_421 (O_421,N_19901,N_19918);
or UO_422 (O_422,N_19939,N_19958);
xnor UO_423 (O_423,N_19981,N_19991);
xnor UO_424 (O_424,N_19929,N_19835);
and UO_425 (O_425,N_19996,N_19892);
nand UO_426 (O_426,N_19982,N_19856);
and UO_427 (O_427,N_19888,N_19810);
nor UO_428 (O_428,N_19972,N_19914);
and UO_429 (O_429,N_19845,N_19969);
xor UO_430 (O_430,N_19921,N_19864);
nand UO_431 (O_431,N_19816,N_19813);
and UO_432 (O_432,N_19856,N_19801);
or UO_433 (O_433,N_19986,N_19835);
nor UO_434 (O_434,N_19944,N_19966);
nand UO_435 (O_435,N_19808,N_19838);
nor UO_436 (O_436,N_19853,N_19806);
and UO_437 (O_437,N_19942,N_19957);
or UO_438 (O_438,N_19917,N_19961);
nand UO_439 (O_439,N_19862,N_19990);
and UO_440 (O_440,N_19800,N_19875);
xor UO_441 (O_441,N_19930,N_19982);
nand UO_442 (O_442,N_19850,N_19954);
and UO_443 (O_443,N_19945,N_19900);
xnor UO_444 (O_444,N_19943,N_19884);
xor UO_445 (O_445,N_19902,N_19908);
xnor UO_446 (O_446,N_19830,N_19842);
nand UO_447 (O_447,N_19843,N_19818);
xor UO_448 (O_448,N_19948,N_19895);
nand UO_449 (O_449,N_19958,N_19969);
nand UO_450 (O_450,N_19935,N_19927);
or UO_451 (O_451,N_19852,N_19810);
nand UO_452 (O_452,N_19995,N_19873);
nand UO_453 (O_453,N_19805,N_19883);
nand UO_454 (O_454,N_19994,N_19995);
xnor UO_455 (O_455,N_19928,N_19871);
xnor UO_456 (O_456,N_19882,N_19925);
and UO_457 (O_457,N_19965,N_19817);
and UO_458 (O_458,N_19839,N_19843);
nand UO_459 (O_459,N_19977,N_19840);
xor UO_460 (O_460,N_19862,N_19910);
xnor UO_461 (O_461,N_19943,N_19897);
xnor UO_462 (O_462,N_19894,N_19929);
or UO_463 (O_463,N_19854,N_19864);
xor UO_464 (O_464,N_19902,N_19950);
nand UO_465 (O_465,N_19969,N_19838);
or UO_466 (O_466,N_19827,N_19930);
nand UO_467 (O_467,N_19900,N_19946);
nor UO_468 (O_468,N_19901,N_19968);
nand UO_469 (O_469,N_19968,N_19819);
nor UO_470 (O_470,N_19973,N_19891);
xnor UO_471 (O_471,N_19860,N_19982);
nor UO_472 (O_472,N_19860,N_19862);
or UO_473 (O_473,N_19835,N_19880);
nand UO_474 (O_474,N_19950,N_19933);
xnor UO_475 (O_475,N_19952,N_19921);
and UO_476 (O_476,N_19972,N_19931);
nand UO_477 (O_477,N_19875,N_19859);
xor UO_478 (O_478,N_19845,N_19959);
nor UO_479 (O_479,N_19897,N_19804);
nor UO_480 (O_480,N_19966,N_19868);
xnor UO_481 (O_481,N_19996,N_19898);
nor UO_482 (O_482,N_19889,N_19942);
nor UO_483 (O_483,N_19823,N_19817);
nor UO_484 (O_484,N_19869,N_19986);
nand UO_485 (O_485,N_19887,N_19997);
nor UO_486 (O_486,N_19911,N_19887);
and UO_487 (O_487,N_19963,N_19842);
nand UO_488 (O_488,N_19924,N_19807);
xor UO_489 (O_489,N_19828,N_19852);
nor UO_490 (O_490,N_19882,N_19872);
nor UO_491 (O_491,N_19895,N_19804);
or UO_492 (O_492,N_19810,N_19809);
nor UO_493 (O_493,N_19821,N_19921);
nand UO_494 (O_494,N_19870,N_19920);
or UO_495 (O_495,N_19824,N_19836);
or UO_496 (O_496,N_19991,N_19902);
and UO_497 (O_497,N_19896,N_19940);
nor UO_498 (O_498,N_19865,N_19830);
nor UO_499 (O_499,N_19882,N_19987);
nand UO_500 (O_500,N_19988,N_19844);
nor UO_501 (O_501,N_19931,N_19843);
or UO_502 (O_502,N_19978,N_19856);
or UO_503 (O_503,N_19845,N_19970);
nand UO_504 (O_504,N_19990,N_19837);
and UO_505 (O_505,N_19976,N_19982);
and UO_506 (O_506,N_19977,N_19874);
nor UO_507 (O_507,N_19871,N_19965);
nand UO_508 (O_508,N_19826,N_19963);
or UO_509 (O_509,N_19935,N_19828);
or UO_510 (O_510,N_19856,N_19840);
or UO_511 (O_511,N_19826,N_19833);
nand UO_512 (O_512,N_19801,N_19966);
and UO_513 (O_513,N_19805,N_19890);
nor UO_514 (O_514,N_19846,N_19818);
nor UO_515 (O_515,N_19938,N_19924);
and UO_516 (O_516,N_19903,N_19912);
and UO_517 (O_517,N_19957,N_19981);
xnor UO_518 (O_518,N_19840,N_19868);
xor UO_519 (O_519,N_19927,N_19943);
or UO_520 (O_520,N_19956,N_19965);
nand UO_521 (O_521,N_19987,N_19880);
nand UO_522 (O_522,N_19823,N_19855);
xnor UO_523 (O_523,N_19829,N_19921);
nor UO_524 (O_524,N_19839,N_19939);
nand UO_525 (O_525,N_19815,N_19976);
and UO_526 (O_526,N_19894,N_19895);
nand UO_527 (O_527,N_19845,N_19921);
nor UO_528 (O_528,N_19847,N_19890);
nor UO_529 (O_529,N_19906,N_19844);
nand UO_530 (O_530,N_19960,N_19928);
xnor UO_531 (O_531,N_19981,N_19911);
nand UO_532 (O_532,N_19996,N_19870);
or UO_533 (O_533,N_19850,N_19882);
nand UO_534 (O_534,N_19969,N_19982);
nand UO_535 (O_535,N_19845,N_19818);
and UO_536 (O_536,N_19940,N_19826);
nand UO_537 (O_537,N_19887,N_19916);
xnor UO_538 (O_538,N_19941,N_19804);
xor UO_539 (O_539,N_19870,N_19984);
and UO_540 (O_540,N_19937,N_19877);
or UO_541 (O_541,N_19817,N_19818);
xor UO_542 (O_542,N_19886,N_19805);
nand UO_543 (O_543,N_19814,N_19983);
and UO_544 (O_544,N_19877,N_19940);
xor UO_545 (O_545,N_19804,N_19978);
nor UO_546 (O_546,N_19939,N_19928);
or UO_547 (O_547,N_19954,N_19941);
and UO_548 (O_548,N_19951,N_19842);
nand UO_549 (O_549,N_19978,N_19999);
nand UO_550 (O_550,N_19936,N_19919);
nor UO_551 (O_551,N_19945,N_19809);
nor UO_552 (O_552,N_19915,N_19947);
xnor UO_553 (O_553,N_19866,N_19867);
nor UO_554 (O_554,N_19868,N_19884);
and UO_555 (O_555,N_19825,N_19994);
and UO_556 (O_556,N_19836,N_19808);
xnor UO_557 (O_557,N_19873,N_19835);
and UO_558 (O_558,N_19805,N_19998);
nor UO_559 (O_559,N_19949,N_19937);
or UO_560 (O_560,N_19892,N_19878);
or UO_561 (O_561,N_19858,N_19913);
and UO_562 (O_562,N_19847,N_19826);
nand UO_563 (O_563,N_19855,N_19928);
or UO_564 (O_564,N_19881,N_19987);
nand UO_565 (O_565,N_19812,N_19891);
nor UO_566 (O_566,N_19951,N_19940);
xnor UO_567 (O_567,N_19922,N_19869);
nor UO_568 (O_568,N_19930,N_19943);
xor UO_569 (O_569,N_19942,N_19980);
nor UO_570 (O_570,N_19802,N_19911);
nand UO_571 (O_571,N_19882,N_19912);
nor UO_572 (O_572,N_19945,N_19961);
nand UO_573 (O_573,N_19942,N_19915);
xor UO_574 (O_574,N_19989,N_19834);
nor UO_575 (O_575,N_19881,N_19892);
nand UO_576 (O_576,N_19802,N_19815);
xor UO_577 (O_577,N_19976,N_19961);
and UO_578 (O_578,N_19964,N_19808);
nand UO_579 (O_579,N_19963,N_19908);
and UO_580 (O_580,N_19979,N_19844);
and UO_581 (O_581,N_19801,N_19879);
and UO_582 (O_582,N_19997,N_19963);
nand UO_583 (O_583,N_19831,N_19889);
and UO_584 (O_584,N_19873,N_19821);
nor UO_585 (O_585,N_19910,N_19993);
xnor UO_586 (O_586,N_19802,N_19895);
and UO_587 (O_587,N_19890,N_19876);
and UO_588 (O_588,N_19841,N_19849);
nor UO_589 (O_589,N_19917,N_19934);
or UO_590 (O_590,N_19859,N_19987);
nand UO_591 (O_591,N_19847,N_19848);
xnor UO_592 (O_592,N_19910,N_19932);
nand UO_593 (O_593,N_19882,N_19806);
xnor UO_594 (O_594,N_19918,N_19942);
nor UO_595 (O_595,N_19950,N_19815);
xnor UO_596 (O_596,N_19822,N_19914);
nor UO_597 (O_597,N_19980,N_19802);
nor UO_598 (O_598,N_19840,N_19907);
nand UO_599 (O_599,N_19948,N_19917);
or UO_600 (O_600,N_19951,N_19807);
or UO_601 (O_601,N_19971,N_19829);
nor UO_602 (O_602,N_19902,N_19855);
nor UO_603 (O_603,N_19891,N_19875);
nand UO_604 (O_604,N_19893,N_19984);
nor UO_605 (O_605,N_19860,N_19988);
and UO_606 (O_606,N_19922,N_19887);
xor UO_607 (O_607,N_19860,N_19840);
and UO_608 (O_608,N_19917,N_19959);
or UO_609 (O_609,N_19852,N_19891);
nand UO_610 (O_610,N_19834,N_19830);
nand UO_611 (O_611,N_19898,N_19823);
or UO_612 (O_612,N_19882,N_19845);
nor UO_613 (O_613,N_19823,N_19929);
nor UO_614 (O_614,N_19976,N_19934);
nor UO_615 (O_615,N_19809,N_19937);
or UO_616 (O_616,N_19914,N_19975);
xor UO_617 (O_617,N_19971,N_19850);
nor UO_618 (O_618,N_19862,N_19955);
and UO_619 (O_619,N_19958,N_19844);
nand UO_620 (O_620,N_19978,N_19940);
nor UO_621 (O_621,N_19886,N_19861);
xnor UO_622 (O_622,N_19894,N_19843);
and UO_623 (O_623,N_19862,N_19820);
or UO_624 (O_624,N_19810,N_19970);
nor UO_625 (O_625,N_19842,N_19944);
or UO_626 (O_626,N_19872,N_19928);
nor UO_627 (O_627,N_19930,N_19867);
or UO_628 (O_628,N_19923,N_19893);
nand UO_629 (O_629,N_19953,N_19827);
nand UO_630 (O_630,N_19855,N_19984);
xnor UO_631 (O_631,N_19968,N_19988);
xnor UO_632 (O_632,N_19800,N_19979);
nand UO_633 (O_633,N_19864,N_19934);
nand UO_634 (O_634,N_19977,N_19942);
and UO_635 (O_635,N_19801,N_19928);
nand UO_636 (O_636,N_19844,N_19936);
xnor UO_637 (O_637,N_19847,N_19938);
and UO_638 (O_638,N_19948,N_19839);
nand UO_639 (O_639,N_19881,N_19964);
and UO_640 (O_640,N_19834,N_19803);
and UO_641 (O_641,N_19978,N_19925);
nor UO_642 (O_642,N_19806,N_19978);
nor UO_643 (O_643,N_19886,N_19825);
and UO_644 (O_644,N_19931,N_19850);
and UO_645 (O_645,N_19944,N_19936);
or UO_646 (O_646,N_19817,N_19871);
xnor UO_647 (O_647,N_19921,N_19983);
xnor UO_648 (O_648,N_19885,N_19986);
nand UO_649 (O_649,N_19807,N_19808);
nor UO_650 (O_650,N_19820,N_19852);
nand UO_651 (O_651,N_19929,N_19837);
xor UO_652 (O_652,N_19955,N_19923);
xor UO_653 (O_653,N_19888,N_19951);
or UO_654 (O_654,N_19880,N_19951);
or UO_655 (O_655,N_19849,N_19868);
or UO_656 (O_656,N_19949,N_19924);
or UO_657 (O_657,N_19888,N_19954);
or UO_658 (O_658,N_19807,N_19843);
or UO_659 (O_659,N_19815,N_19878);
nor UO_660 (O_660,N_19997,N_19952);
and UO_661 (O_661,N_19938,N_19834);
and UO_662 (O_662,N_19829,N_19876);
and UO_663 (O_663,N_19850,N_19990);
xor UO_664 (O_664,N_19935,N_19871);
and UO_665 (O_665,N_19963,N_19907);
xnor UO_666 (O_666,N_19960,N_19861);
nand UO_667 (O_667,N_19845,N_19968);
nand UO_668 (O_668,N_19940,N_19912);
or UO_669 (O_669,N_19896,N_19839);
and UO_670 (O_670,N_19815,N_19888);
and UO_671 (O_671,N_19978,N_19991);
nor UO_672 (O_672,N_19851,N_19898);
nor UO_673 (O_673,N_19843,N_19889);
xor UO_674 (O_674,N_19860,N_19839);
nor UO_675 (O_675,N_19900,N_19810);
or UO_676 (O_676,N_19873,N_19800);
nand UO_677 (O_677,N_19857,N_19827);
or UO_678 (O_678,N_19910,N_19884);
and UO_679 (O_679,N_19958,N_19830);
and UO_680 (O_680,N_19854,N_19959);
or UO_681 (O_681,N_19848,N_19854);
xnor UO_682 (O_682,N_19876,N_19912);
and UO_683 (O_683,N_19870,N_19811);
and UO_684 (O_684,N_19981,N_19831);
and UO_685 (O_685,N_19863,N_19909);
nor UO_686 (O_686,N_19852,N_19841);
xnor UO_687 (O_687,N_19940,N_19962);
and UO_688 (O_688,N_19984,N_19846);
nor UO_689 (O_689,N_19888,N_19990);
nand UO_690 (O_690,N_19812,N_19876);
xor UO_691 (O_691,N_19867,N_19984);
xor UO_692 (O_692,N_19923,N_19984);
and UO_693 (O_693,N_19860,N_19847);
and UO_694 (O_694,N_19955,N_19875);
nand UO_695 (O_695,N_19878,N_19828);
nand UO_696 (O_696,N_19919,N_19980);
xnor UO_697 (O_697,N_19996,N_19972);
xor UO_698 (O_698,N_19827,N_19878);
and UO_699 (O_699,N_19856,N_19921);
nor UO_700 (O_700,N_19914,N_19994);
nand UO_701 (O_701,N_19825,N_19896);
and UO_702 (O_702,N_19824,N_19813);
xnor UO_703 (O_703,N_19994,N_19816);
and UO_704 (O_704,N_19842,N_19887);
nand UO_705 (O_705,N_19828,N_19869);
and UO_706 (O_706,N_19944,N_19958);
nand UO_707 (O_707,N_19821,N_19866);
and UO_708 (O_708,N_19999,N_19887);
xor UO_709 (O_709,N_19986,N_19966);
nand UO_710 (O_710,N_19981,N_19961);
xor UO_711 (O_711,N_19940,N_19919);
nor UO_712 (O_712,N_19869,N_19843);
or UO_713 (O_713,N_19852,N_19937);
or UO_714 (O_714,N_19876,N_19994);
nand UO_715 (O_715,N_19866,N_19962);
or UO_716 (O_716,N_19869,N_19833);
or UO_717 (O_717,N_19828,N_19998);
nand UO_718 (O_718,N_19801,N_19872);
nand UO_719 (O_719,N_19879,N_19887);
or UO_720 (O_720,N_19921,N_19810);
or UO_721 (O_721,N_19830,N_19858);
and UO_722 (O_722,N_19967,N_19829);
and UO_723 (O_723,N_19925,N_19815);
or UO_724 (O_724,N_19912,N_19867);
or UO_725 (O_725,N_19947,N_19921);
and UO_726 (O_726,N_19870,N_19847);
and UO_727 (O_727,N_19878,N_19836);
nand UO_728 (O_728,N_19888,N_19931);
nor UO_729 (O_729,N_19885,N_19852);
xnor UO_730 (O_730,N_19800,N_19900);
or UO_731 (O_731,N_19801,N_19938);
nand UO_732 (O_732,N_19933,N_19892);
and UO_733 (O_733,N_19844,N_19963);
nor UO_734 (O_734,N_19844,N_19853);
xnor UO_735 (O_735,N_19848,N_19843);
xnor UO_736 (O_736,N_19990,N_19865);
or UO_737 (O_737,N_19818,N_19987);
and UO_738 (O_738,N_19820,N_19940);
and UO_739 (O_739,N_19958,N_19946);
and UO_740 (O_740,N_19868,N_19928);
nand UO_741 (O_741,N_19969,N_19816);
nand UO_742 (O_742,N_19979,N_19853);
nor UO_743 (O_743,N_19823,N_19853);
or UO_744 (O_744,N_19910,N_19824);
nor UO_745 (O_745,N_19955,N_19813);
xor UO_746 (O_746,N_19883,N_19801);
xor UO_747 (O_747,N_19852,N_19962);
nor UO_748 (O_748,N_19802,N_19937);
and UO_749 (O_749,N_19950,N_19974);
nand UO_750 (O_750,N_19925,N_19832);
nand UO_751 (O_751,N_19820,N_19909);
and UO_752 (O_752,N_19980,N_19924);
nand UO_753 (O_753,N_19996,N_19859);
nand UO_754 (O_754,N_19821,N_19845);
nand UO_755 (O_755,N_19846,N_19884);
and UO_756 (O_756,N_19843,N_19810);
and UO_757 (O_757,N_19989,N_19849);
xor UO_758 (O_758,N_19935,N_19880);
and UO_759 (O_759,N_19960,N_19899);
and UO_760 (O_760,N_19831,N_19956);
or UO_761 (O_761,N_19932,N_19879);
nand UO_762 (O_762,N_19863,N_19949);
nor UO_763 (O_763,N_19920,N_19957);
nor UO_764 (O_764,N_19912,N_19838);
nand UO_765 (O_765,N_19880,N_19957);
xor UO_766 (O_766,N_19900,N_19801);
xnor UO_767 (O_767,N_19956,N_19888);
xor UO_768 (O_768,N_19907,N_19893);
and UO_769 (O_769,N_19879,N_19843);
xnor UO_770 (O_770,N_19936,N_19921);
or UO_771 (O_771,N_19912,N_19815);
and UO_772 (O_772,N_19959,N_19840);
or UO_773 (O_773,N_19849,N_19977);
and UO_774 (O_774,N_19925,N_19977);
or UO_775 (O_775,N_19888,N_19860);
nand UO_776 (O_776,N_19929,N_19804);
xnor UO_777 (O_777,N_19861,N_19910);
nor UO_778 (O_778,N_19960,N_19821);
nand UO_779 (O_779,N_19868,N_19856);
nand UO_780 (O_780,N_19827,N_19844);
xor UO_781 (O_781,N_19985,N_19944);
nand UO_782 (O_782,N_19967,N_19910);
nand UO_783 (O_783,N_19995,N_19805);
xnor UO_784 (O_784,N_19942,N_19808);
or UO_785 (O_785,N_19963,N_19922);
and UO_786 (O_786,N_19907,N_19990);
or UO_787 (O_787,N_19851,N_19844);
xor UO_788 (O_788,N_19940,N_19976);
or UO_789 (O_789,N_19840,N_19810);
or UO_790 (O_790,N_19870,N_19802);
and UO_791 (O_791,N_19948,N_19904);
or UO_792 (O_792,N_19982,N_19869);
xnor UO_793 (O_793,N_19920,N_19923);
or UO_794 (O_794,N_19866,N_19806);
nand UO_795 (O_795,N_19866,N_19971);
or UO_796 (O_796,N_19951,N_19887);
nor UO_797 (O_797,N_19897,N_19838);
nor UO_798 (O_798,N_19879,N_19983);
nand UO_799 (O_799,N_19956,N_19822);
xnor UO_800 (O_800,N_19894,N_19988);
and UO_801 (O_801,N_19953,N_19976);
and UO_802 (O_802,N_19903,N_19962);
or UO_803 (O_803,N_19934,N_19971);
nor UO_804 (O_804,N_19956,N_19908);
nor UO_805 (O_805,N_19970,N_19863);
nand UO_806 (O_806,N_19882,N_19856);
or UO_807 (O_807,N_19943,N_19983);
xor UO_808 (O_808,N_19948,N_19903);
xnor UO_809 (O_809,N_19858,N_19992);
or UO_810 (O_810,N_19931,N_19960);
nor UO_811 (O_811,N_19960,N_19830);
and UO_812 (O_812,N_19896,N_19927);
or UO_813 (O_813,N_19998,N_19927);
xor UO_814 (O_814,N_19821,N_19888);
and UO_815 (O_815,N_19916,N_19909);
nand UO_816 (O_816,N_19912,N_19827);
nand UO_817 (O_817,N_19896,N_19818);
or UO_818 (O_818,N_19877,N_19928);
xnor UO_819 (O_819,N_19945,N_19838);
or UO_820 (O_820,N_19861,N_19965);
and UO_821 (O_821,N_19888,N_19856);
xor UO_822 (O_822,N_19948,N_19991);
and UO_823 (O_823,N_19881,N_19848);
nand UO_824 (O_824,N_19847,N_19946);
and UO_825 (O_825,N_19962,N_19980);
or UO_826 (O_826,N_19913,N_19841);
and UO_827 (O_827,N_19989,N_19853);
xor UO_828 (O_828,N_19993,N_19899);
nand UO_829 (O_829,N_19989,N_19905);
xnor UO_830 (O_830,N_19996,N_19918);
or UO_831 (O_831,N_19905,N_19802);
nor UO_832 (O_832,N_19997,N_19955);
or UO_833 (O_833,N_19845,N_19877);
nand UO_834 (O_834,N_19949,N_19955);
or UO_835 (O_835,N_19970,N_19830);
and UO_836 (O_836,N_19960,N_19945);
nor UO_837 (O_837,N_19827,N_19817);
and UO_838 (O_838,N_19994,N_19915);
and UO_839 (O_839,N_19871,N_19840);
nand UO_840 (O_840,N_19934,N_19935);
nand UO_841 (O_841,N_19951,N_19932);
nand UO_842 (O_842,N_19822,N_19981);
and UO_843 (O_843,N_19900,N_19832);
nor UO_844 (O_844,N_19846,N_19997);
xnor UO_845 (O_845,N_19862,N_19866);
nand UO_846 (O_846,N_19901,N_19931);
nor UO_847 (O_847,N_19958,N_19948);
nor UO_848 (O_848,N_19935,N_19836);
nand UO_849 (O_849,N_19993,N_19920);
and UO_850 (O_850,N_19925,N_19892);
nand UO_851 (O_851,N_19905,N_19999);
or UO_852 (O_852,N_19965,N_19888);
nor UO_853 (O_853,N_19959,N_19974);
xor UO_854 (O_854,N_19857,N_19805);
xnor UO_855 (O_855,N_19947,N_19807);
nand UO_856 (O_856,N_19838,N_19964);
nor UO_857 (O_857,N_19860,N_19965);
nor UO_858 (O_858,N_19846,N_19858);
nand UO_859 (O_859,N_19887,N_19958);
nand UO_860 (O_860,N_19983,N_19920);
nor UO_861 (O_861,N_19964,N_19916);
xnor UO_862 (O_862,N_19945,N_19844);
nor UO_863 (O_863,N_19849,N_19994);
or UO_864 (O_864,N_19898,N_19850);
or UO_865 (O_865,N_19889,N_19824);
nand UO_866 (O_866,N_19947,N_19867);
or UO_867 (O_867,N_19916,N_19917);
xnor UO_868 (O_868,N_19829,N_19919);
and UO_869 (O_869,N_19867,N_19918);
and UO_870 (O_870,N_19861,N_19813);
xor UO_871 (O_871,N_19885,N_19966);
xnor UO_872 (O_872,N_19987,N_19805);
xnor UO_873 (O_873,N_19935,N_19877);
or UO_874 (O_874,N_19809,N_19918);
nor UO_875 (O_875,N_19930,N_19969);
or UO_876 (O_876,N_19910,N_19890);
and UO_877 (O_877,N_19932,N_19858);
or UO_878 (O_878,N_19958,N_19897);
nor UO_879 (O_879,N_19950,N_19887);
or UO_880 (O_880,N_19879,N_19862);
and UO_881 (O_881,N_19931,N_19944);
xor UO_882 (O_882,N_19873,N_19816);
and UO_883 (O_883,N_19966,N_19812);
and UO_884 (O_884,N_19931,N_19824);
or UO_885 (O_885,N_19937,N_19904);
nand UO_886 (O_886,N_19866,N_19953);
nand UO_887 (O_887,N_19809,N_19935);
nor UO_888 (O_888,N_19954,N_19992);
and UO_889 (O_889,N_19892,N_19896);
or UO_890 (O_890,N_19834,N_19947);
and UO_891 (O_891,N_19846,N_19955);
nand UO_892 (O_892,N_19805,N_19869);
and UO_893 (O_893,N_19996,N_19845);
nand UO_894 (O_894,N_19859,N_19837);
and UO_895 (O_895,N_19909,N_19941);
xor UO_896 (O_896,N_19825,N_19984);
and UO_897 (O_897,N_19994,N_19968);
xor UO_898 (O_898,N_19914,N_19928);
or UO_899 (O_899,N_19962,N_19863);
nand UO_900 (O_900,N_19953,N_19845);
nand UO_901 (O_901,N_19830,N_19934);
xor UO_902 (O_902,N_19929,N_19953);
nand UO_903 (O_903,N_19975,N_19896);
nor UO_904 (O_904,N_19962,N_19994);
nor UO_905 (O_905,N_19898,N_19931);
nor UO_906 (O_906,N_19995,N_19847);
nand UO_907 (O_907,N_19871,N_19920);
nand UO_908 (O_908,N_19936,N_19880);
nor UO_909 (O_909,N_19839,N_19925);
xnor UO_910 (O_910,N_19836,N_19927);
nor UO_911 (O_911,N_19813,N_19962);
xnor UO_912 (O_912,N_19847,N_19883);
nor UO_913 (O_913,N_19883,N_19815);
or UO_914 (O_914,N_19821,N_19875);
nand UO_915 (O_915,N_19875,N_19978);
xor UO_916 (O_916,N_19873,N_19984);
nor UO_917 (O_917,N_19989,N_19840);
nand UO_918 (O_918,N_19861,N_19902);
nor UO_919 (O_919,N_19948,N_19952);
or UO_920 (O_920,N_19910,N_19908);
nand UO_921 (O_921,N_19854,N_19829);
nor UO_922 (O_922,N_19951,N_19835);
nor UO_923 (O_923,N_19804,N_19885);
and UO_924 (O_924,N_19841,N_19878);
or UO_925 (O_925,N_19910,N_19804);
and UO_926 (O_926,N_19973,N_19953);
nor UO_927 (O_927,N_19936,N_19821);
nand UO_928 (O_928,N_19861,N_19976);
or UO_929 (O_929,N_19920,N_19951);
xnor UO_930 (O_930,N_19954,N_19887);
xor UO_931 (O_931,N_19983,N_19952);
or UO_932 (O_932,N_19893,N_19802);
xor UO_933 (O_933,N_19810,N_19882);
xor UO_934 (O_934,N_19943,N_19838);
or UO_935 (O_935,N_19812,N_19887);
or UO_936 (O_936,N_19858,N_19843);
nor UO_937 (O_937,N_19838,N_19811);
xnor UO_938 (O_938,N_19975,N_19988);
xnor UO_939 (O_939,N_19982,N_19912);
nand UO_940 (O_940,N_19845,N_19913);
xor UO_941 (O_941,N_19819,N_19984);
xor UO_942 (O_942,N_19856,N_19886);
nor UO_943 (O_943,N_19809,N_19808);
xor UO_944 (O_944,N_19947,N_19951);
nor UO_945 (O_945,N_19906,N_19912);
xor UO_946 (O_946,N_19924,N_19842);
xor UO_947 (O_947,N_19842,N_19969);
nor UO_948 (O_948,N_19889,N_19960);
and UO_949 (O_949,N_19805,N_19925);
nand UO_950 (O_950,N_19900,N_19967);
or UO_951 (O_951,N_19970,N_19852);
nand UO_952 (O_952,N_19961,N_19925);
xnor UO_953 (O_953,N_19819,N_19885);
nand UO_954 (O_954,N_19830,N_19961);
and UO_955 (O_955,N_19834,N_19847);
or UO_956 (O_956,N_19829,N_19824);
or UO_957 (O_957,N_19890,N_19972);
nor UO_958 (O_958,N_19880,N_19942);
nor UO_959 (O_959,N_19943,N_19863);
nand UO_960 (O_960,N_19905,N_19810);
xnor UO_961 (O_961,N_19859,N_19977);
and UO_962 (O_962,N_19997,N_19947);
and UO_963 (O_963,N_19899,N_19815);
or UO_964 (O_964,N_19906,N_19833);
nor UO_965 (O_965,N_19829,N_19897);
and UO_966 (O_966,N_19827,N_19838);
xnor UO_967 (O_967,N_19899,N_19814);
and UO_968 (O_968,N_19930,N_19935);
nor UO_969 (O_969,N_19923,N_19885);
xor UO_970 (O_970,N_19914,N_19956);
nor UO_971 (O_971,N_19997,N_19896);
xor UO_972 (O_972,N_19815,N_19879);
xor UO_973 (O_973,N_19852,N_19925);
nand UO_974 (O_974,N_19925,N_19846);
nor UO_975 (O_975,N_19879,N_19950);
or UO_976 (O_976,N_19808,N_19865);
and UO_977 (O_977,N_19954,N_19959);
nor UO_978 (O_978,N_19888,N_19994);
nor UO_979 (O_979,N_19977,N_19950);
nor UO_980 (O_980,N_19899,N_19830);
nand UO_981 (O_981,N_19850,N_19800);
or UO_982 (O_982,N_19860,N_19817);
nor UO_983 (O_983,N_19977,N_19889);
or UO_984 (O_984,N_19907,N_19908);
and UO_985 (O_985,N_19864,N_19955);
nor UO_986 (O_986,N_19864,N_19843);
nor UO_987 (O_987,N_19935,N_19888);
nand UO_988 (O_988,N_19975,N_19891);
nor UO_989 (O_989,N_19824,N_19991);
or UO_990 (O_990,N_19909,N_19937);
nor UO_991 (O_991,N_19955,N_19933);
and UO_992 (O_992,N_19945,N_19919);
and UO_993 (O_993,N_19908,N_19878);
and UO_994 (O_994,N_19811,N_19932);
or UO_995 (O_995,N_19981,N_19840);
or UO_996 (O_996,N_19870,N_19901);
and UO_997 (O_997,N_19804,N_19879);
and UO_998 (O_998,N_19881,N_19991);
and UO_999 (O_999,N_19892,N_19919);
xnor UO_1000 (O_1000,N_19809,N_19876);
and UO_1001 (O_1001,N_19800,N_19945);
or UO_1002 (O_1002,N_19939,N_19920);
xnor UO_1003 (O_1003,N_19880,N_19894);
and UO_1004 (O_1004,N_19967,N_19803);
and UO_1005 (O_1005,N_19879,N_19994);
or UO_1006 (O_1006,N_19808,N_19895);
and UO_1007 (O_1007,N_19882,N_19989);
or UO_1008 (O_1008,N_19877,N_19859);
xnor UO_1009 (O_1009,N_19981,N_19936);
or UO_1010 (O_1010,N_19930,N_19830);
nor UO_1011 (O_1011,N_19888,N_19993);
and UO_1012 (O_1012,N_19885,N_19948);
nor UO_1013 (O_1013,N_19849,N_19866);
xor UO_1014 (O_1014,N_19912,N_19926);
xor UO_1015 (O_1015,N_19830,N_19878);
or UO_1016 (O_1016,N_19971,N_19926);
xnor UO_1017 (O_1017,N_19952,N_19946);
nand UO_1018 (O_1018,N_19980,N_19902);
xor UO_1019 (O_1019,N_19812,N_19987);
nor UO_1020 (O_1020,N_19829,N_19902);
and UO_1021 (O_1021,N_19920,N_19832);
nand UO_1022 (O_1022,N_19854,N_19833);
xor UO_1023 (O_1023,N_19922,N_19845);
nor UO_1024 (O_1024,N_19939,N_19987);
nor UO_1025 (O_1025,N_19988,N_19826);
and UO_1026 (O_1026,N_19895,N_19933);
nor UO_1027 (O_1027,N_19957,N_19969);
and UO_1028 (O_1028,N_19867,N_19974);
and UO_1029 (O_1029,N_19918,N_19977);
xnor UO_1030 (O_1030,N_19802,N_19925);
nand UO_1031 (O_1031,N_19855,N_19888);
nor UO_1032 (O_1032,N_19841,N_19999);
nor UO_1033 (O_1033,N_19924,N_19932);
or UO_1034 (O_1034,N_19933,N_19858);
xnor UO_1035 (O_1035,N_19849,N_19869);
and UO_1036 (O_1036,N_19873,N_19871);
nor UO_1037 (O_1037,N_19928,N_19953);
nand UO_1038 (O_1038,N_19916,N_19869);
nand UO_1039 (O_1039,N_19890,N_19946);
and UO_1040 (O_1040,N_19811,N_19960);
nor UO_1041 (O_1041,N_19952,N_19951);
nor UO_1042 (O_1042,N_19923,N_19978);
or UO_1043 (O_1043,N_19877,N_19876);
xor UO_1044 (O_1044,N_19904,N_19971);
and UO_1045 (O_1045,N_19872,N_19972);
xnor UO_1046 (O_1046,N_19925,N_19969);
nor UO_1047 (O_1047,N_19829,N_19861);
and UO_1048 (O_1048,N_19972,N_19983);
xnor UO_1049 (O_1049,N_19839,N_19950);
nand UO_1050 (O_1050,N_19974,N_19996);
nand UO_1051 (O_1051,N_19984,N_19955);
nand UO_1052 (O_1052,N_19964,N_19933);
xor UO_1053 (O_1053,N_19824,N_19857);
nor UO_1054 (O_1054,N_19817,N_19840);
nand UO_1055 (O_1055,N_19945,N_19908);
or UO_1056 (O_1056,N_19893,N_19979);
nor UO_1057 (O_1057,N_19950,N_19934);
xor UO_1058 (O_1058,N_19903,N_19817);
nand UO_1059 (O_1059,N_19898,N_19995);
nand UO_1060 (O_1060,N_19867,N_19869);
and UO_1061 (O_1061,N_19858,N_19956);
or UO_1062 (O_1062,N_19863,N_19921);
xor UO_1063 (O_1063,N_19978,N_19902);
or UO_1064 (O_1064,N_19964,N_19960);
or UO_1065 (O_1065,N_19964,N_19997);
nor UO_1066 (O_1066,N_19971,N_19855);
nor UO_1067 (O_1067,N_19987,N_19986);
nor UO_1068 (O_1068,N_19890,N_19891);
and UO_1069 (O_1069,N_19857,N_19985);
and UO_1070 (O_1070,N_19968,N_19829);
and UO_1071 (O_1071,N_19856,N_19824);
nor UO_1072 (O_1072,N_19961,N_19978);
xor UO_1073 (O_1073,N_19818,N_19873);
and UO_1074 (O_1074,N_19812,N_19968);
nor UO_1075 (O_1075,N_19842,N_19978);
xor UO_1076 (O_1076,N_19940,N_19986);
nand UO_1077 (O_1077,N_19967,N_19991);
nand UO_1078 (O_1078,N_19876,N_19867);
and UO_1079 (O_1079,N_19857,N_19994);
nor UO_1080 (O_1080,N_19979,N_19981);
and UO_1081 (O_1081,N_19904,N_19859);
nand UO_1082 (O_1082,N_19971,N_19878);
or UO_1083 (O_1083,N_19802,N_19810);
nand UO_1084 (O_1084,N_19961,N_19865);
xor UO_1085 (O_1085,N_19989,N_19852);
xnor UO_1086 (O_1086,N_19848,N_19972);
or UO_1087 (O_1087,N_19968,N_19951);
or UO_1088 (O_1088,N_19886,N_19874);
nor UO_1089 (O_1089,N_19836,N_19942);
nand UO_1090 (O_1090,N_19941,N_19823);
and UO_1091 (O_1091,N_19893,N_19885);
and UO_1092 (O_1092,N_19872,N_19904);
nand UO_1093 (O_1093,N_19883,N_19800);
nand UO_1094 (O_1094,N_19998,N_19834);
xor UO_1095 (O_1095,N_19870,N_19939);
nor UO_1096 (O_1096,N_19984,N_19868);
xor UO_1097 (O_1097,N_19955,N_19887);
nand UO_1098 (O_1098,N_19854,N_19855);
xor UO_1099 (O_1099,N_19818,N_19884);
nand UO_1100 (O_1100,N_19947,N_19826);
or UO_1101 (O_1101,N_19916,N_19834);
and UO_1102 (O_1102,N_19870,N_19863);
nor UO_1103 (O_1103,N_19997,N_19878);
nand UO_1104 (O_1104,N_19985,N_19975);
and UO_1105 (O_1105,N_19955,N_19954);
nor UO_1106 (O_1106,N_19968,N_19838);
or UO_1107 (O_1107,N_19829,N_19803);
nor UO_1108 (O_1108,N_19861,N_19866);
nand UO_1109 (O_1109,N_19829,N_19882);
and UO_1110 (O_1110,N_19931,N_19879);
nand UO_1111 (O_1111,N_19981,N_19910);
or UO_1112 (O_1112,N_19947,N_19833);
or UO_1113 (O_1113,N_19968,N_19945);
nor UO_1114 (O_1114,N_19975,N_19817);
xor UO_1115 (O_1115,N_19812,N_19857);
and UO_1116 (O_1116,N_19800,N_19983);
nor UO_1117 (O_1117,N_19926,N_19909);
or UO_1118 (O_1118,N_19948,N_19817);
nor UO_1119 (O_1119,N_19947,N_19800);
xnor UO_1120 (O_1120,N_19854,N_19912);
or UO_1121 (O_1121,N_19900,N_19941);
and UO_1122 (O_1122,N_19918,N_19826);
nand UO_1123 (O_1123,N_19950,N_19867);
and UO_1124 (O_1124,N_19965,N_19855);
or UO_1125 (O_1125,N_19984,N_19962);
and UO_1126 (O_1126,N_19832,N_19846);
nor UO_1127 (O_1127,N_19957,N_19868);
xor UO_1128 (O_1128,N_19972,N_19984);
or UO_1129 (O_1129,N_19888,N_19845);
nor UO_1130 (O_1130,N_19814,N_19845);
xor UO_1131 (O_1131,N_19884,N_19920);
and UO_1132 (O_1132,N_19826,N_19949);
nand UO_1133 (O_1133,N_19896,N_19894);
xnor UO_1134 (O_1134,N_19800,N_19815);
nand UO_1135 (O_1135,N_19860,N_19866);
xnor UO_1136 (O_1136,N_19847,N_19891);
and UO_1137 (O_1137,N_19896,N_19871);
xor UO_1138 (O_1138,N_19962,N_19910);
or UO_1139 (O_1139,N_19978,N_19977);
nor UO_1140 (O_1140,N_19993,N_19964);
xor UO_1141 (O_1141,N_19959,N_19810);
nand UO_1142 (O_1142,N_19908,N_19930);
xor UO_1143 (O_1143,N_19860,N_19878);
or UO_1144 (O_1144,N_19941,N_19910);
nand UO_1145 (O_1145,N_19881,N_19875);
nand UO_1146 (O_1146,N_19947,N_19852);
nand UO_1147 (O_1147,N_19974,N_19864);
nor UO_1148 (O_1148,N_19844,N_19850);
nor UO_1149 (O_1149,N_19932,N_19973);
nor UO_1150 (O_1150,N_19957,N_19935);
or UO_1151 (O_1151,N_19903,N_19875);
and UO_1152 (O_1152,N_19990,N_19832);
xor UO_1153 (O_1153,N_19800,N_19986);
or UO_1154 (O_1154,N_19928,N_19915);
or UO_1155 (O_1155,N_19853,N_19972);
and UO_1156 (O_1156,N_19901,N_19888);
xor UO_1157 (O_1157,N_19963,N_19879);
xor UO_1158 (O_1158,N_19810,N_19830);
or UO_1159 (O_1159,N_19906,N_19911);
nand UO_1160 (O_1160,N_19876,N_19906);
or UO_1161 (O_1161,N_19872,N_19844);
xor UO_1162 (O_1162,N_19952,N_19929);
nand UO_1163 (O_1163,N_19808,N_19989);
xor UO_1164 (O_1164,N_19985,N_19829);
nor UO_1165 (O_1165,N_19949,N_19982);
nand UO_1166 (O_1166,N_19881,N_19833);
and UO_1167 (O_1167,N_19909,N_19813);
and UO_1168 (O_1168,N_19838,N_19909);
or UO_1169 (O_1169,N_19839,N_19840);
or UO_1170 (O_1170,N_19901,N_19929);
nor UO_1171 (O_1171,N_19901,N_19848);
or UO_1172 (O_1172,N_19859,N_19972);
nor UO_1173 (O_1173,N_19812,N_19934);
or UO_1174 (O_1174,N_19995,N_19914);
nand UO_1175 (O_1175,N_19850,N_19929);
or UO_1176 (O_1176,N_19806,N_19900);
nor UO_1177 (O_1177,N_19811,N_19850);
xnor UO_1178 (O_1178,N_19940,N_19804);
nand UO_1179 (O_1179,N_19822,N_19943);
xnor UO_1180 (O_1180,N_19960,N_19900);
or UO_1181 (O_1181,N_19871,N_19836);
and UO_1182 (O_1182,N_19954,N_19811);
nor UO_1183 (O_1183,N_19876,N_19963);
and UO_1184 (O_1184,N_19868,N_19878);
and UO_1185 (O_1185,N_19961,N_19942);
nor UO_1186 (O_1186,N_19845,N_19898);
xnor UO_1187 (O_1187,N_19963,N_19803);
and UO_1188 (O_1188,N_19839,N_19845);
or UO_1189 (O_1189,N_19848,N_19857);
nor UO_1190 (O_1190,N_19993,N_19943);
or UO_1191 (O_1191,N_19838,N_19977);
xor UO_1192 (O_1192,N_19972,N_19916);
nand UO_1193 (O_1193,N_19853,N_19923);
xor UO_1194 (O_1194,N_19905,N_19925);
nand UO_1195 (O_1195,N_19804,N_19981);
nand UO_1196 (O_1196,N_19920,N_19940);
nand UO_1197 (O_1197,N_19926,N_19897);
nor UO_1198 (O_1198,N_19906,N_19882);
xnor UO_1199 (O_1199,N_19862,N_19837);
xnor UO_1200 (O_1200,N_19814,N_19878);
or UO_1201 (O_1201,N_19870,N_19941);
nor UO_1202 (O_1202,N_19918,N_19893);
nand UO_1203 (O_1203,N_19811,N_19985);
and UO_1204 (O_1204,N_19944,N_19997);
and UO_1205 (O_1205,N_19942,N_19866);
or UO_1206 (O_1206,N_19949,N_19872);
xnor UO_1207 (O_1207,N_19886,N_19871);
xor UO_1208 (O_1208,N_19800,N_19831);
nor UO_1209 (O_1209,N_19913,N_19932);
nor UO_1210 (O_1210,N_19996,N_19882);
nor UO_1211 (O_1211,N_19864,N_19950);
xor UO_1212 (O_1212,N_19815,N_19934);
xor UO_1213 (O_1213,N_19930,N_19891);
nand UO_1214 (O_1214,N_19901,N_19861);
and UO_1215 (O_1215,N_19911,N_19869);
nand UO_1216 (O_1216,N_19905,N_19913);
xor UO_1217 (O_1217,N_19968,N_19975);
and UO_1218 (O_1218,N_19959,N_19914);
xor UO_1219 (O_1219,N_19859,N_19973);
and UO_1220 (O_1220,N_19927,N_19912);
xnor UO_1221 (O_1221,N_19876,N_19851);
nand UO_1222 (O_1222,N_19869,N_19893);
nor UO_1223 (O_1223,N_19824,N_19916);
or UO_1224 (O_1224,N_19836,N_19978);
and UO_1225 (O_1225,N_19916,N_19999);
xnor UO_1226 (O_1226,N_19929,N_19865);
nand UO_1227 (O_1227,N_19999,N_19920);
or UO_1228 (O_1228,N_19875,N_19842);
xnor UO_1229 (O_1229,N_19973,N_19821);
or UO_1230 (O_1230,N_19872,N_19805);
xor UO_1231 (O_1231,N_19927,N_19986);
and UO_1232 (O_1232,N_19921,N_19865);
xor UO_1233 (O_1233,N_19974,N_19837);
and UO_1234 (O_1234,N_19801,N_19987);
xnor UO_1235 (O_1235,N_19897,N_19915);
nor UO_1236 (O_1236,N_19891,N_19954);
xnor UO_1237 (O_1237,N_19931,N_19981);
and UO_1238 (O_1238,N_19944,N_19802);
or UO_1239 (O_1239,N_19871,N_19860);
nor UO_1240 (O_1240,N_19879,N_19896);
and UO_1241 (O_1241,N_19956,N_19941);
xnor UO_1242 (O_1242,N_19932,N_19968);
nand UO_1243 (O_1243,N_19855,N_19809);
or UO_1244 (O_1244,N_19857,N_19865);
and UO_1245 (O_1245,N_19818,N_19902);
or UO_1246 (O_1246,N_19839,N_19970);
and UO_1247 (O_1247,N_19875,N_19958);
or UO_1248 (O_1248,N_19972,N_19942);
and UO_1249 (O_1249,N_19934,N_19901);
and UO_1250 (O_1250,N_19904,N_19819);
xor UO_1251 (O_1251,N_19891,N_19833);
or UO_1252 (O_1252,N_19949,N_19881);
xnor UO_1253 (O_1253,N_19824,N_19963);
and UO_1254 (O_1254,N_19865,N_19997);
nor UO_1255 (O_1255,N_19849,N_19933);
nand UO_1256 (O_1256,N_19849,N_19818);
or UO_1257 (O_1257,N_19954,N_19999);
or UO_1258 (O_1258,N_19941,N_19819);
nor UO_1259 (O_1259,N_19949,N_19929);
nor UO_1260 (O_1260,N_19877,N_19901);
nand UO_1261 (O_1261,N_19808,N_19831);
nand UO_1262 (O_1262,N_19990,N_19807);
nand UO_1263 (O_1263,N_19888,N_19950);
nor UO_1264 (O_1264,N_19823,N_19842);
or UO_1265 (O_1265,N_19884,N_19843);
or UO_1266 (O_1266,N_19979,N_19971);
xnor UO_1267 (O_1267,N_19847,N_19971);
nand UO_1268 (O_1268,N_19896,N_19809);
or UO_1269 (O_1269,N_19950,N_19975);
nor UO_1270 (O_1270,N_19907,N_19838);
xor UO_1271 (O_1271,N_19893,N_19832);
or UO_1272 (O_1272,N_19920,N_19839);
and UO_1273 (O_1273,N_19845,N_19858);
nor UO_1274 (O_1274,N_19960,N_19869);
nand UO_1275 (O_1275,N_19994,N_19841);
nor UO_1276 (O_1276,N_19901,N_19987);
and UO_1277 (O_1277,N_19800,N_19923);
or UO_1278 (O_1278,N_19977,N_19832);
nor UO_1279 (O_1279,N_19935,N_19996);
xor UO_1280 (O_1280,N_19899,N_19910);
or UO_1281 (O_1281,N_19982,N_19963);
nor UO_1282 (O_1282,N_19840,N_19904);
nor UO_1283 (O_1283,N_19926,N_19884);
and UO_1284 (O_1284,N_19893,N_19961);
xnor UO_1285 (O_1285,N_19930,N_19906);
xnor UO_1286 (O_1286,N_19937,N_19813);
nand UO_1287 (O_1287,N_19931,N_19833);
or UO_1288 (O_1288,N_19911,N_19933);
or UO_1289 (O_1289,N_19901,N_19914);
and UO_1290 (O_1290,N_19887,N_19888);
xor UO_1291 (O_1291,N_19935,N_19844);
nor UO_1292 (O_1292,N_19855,N_19921);
or UO_1293 (O_1293,N_19929,N_19866);
nand UO_1294 (O_1294,N_19956,N_19894);
and UO_1295 (O_1295,N_19995,N_19801);
nand UO_1296 (O_1296,N_19993,N_19952);
nand UO_1297 (O_1297,N_19803,N_19886);
nand UO_1298 (O_1298,N_19950,N_19927);
or UO_1299 (O_1299,N_19854,N_19991);
xnor UO_1300 (O_1300,N_19886,N_19995);
or UO_1301 (O_1301,N_19810,N_19878);
nor UO_1302 (O_1302,N_19832,N_19922);
and UO_1303 (O_1303,N_19856,N_19838);
or UO_1304 (O_1304,N_19894,N_19945);
nand UO_1305 (O_1305,N_19926,N_19981);
nand UO_1306 (O_1306,N_19882,N_19986);
xor UO_1307 (O_1307,N_19863,N_19896);
xnor UO_1308 (O_1308,N_19892,N_19953);
xor UO_1309 (O_1309,N_19805,N_19836);
and UO_1310 (O_1310,N_19803,N_19959);
and UO_1311 (O_1311,N_19900,N_19870);
xnor UO_1312 (O_1312,N_19825,N_19900);
or UO_1313 (O_1313,N_19978,N_19998);
or UO_1314 (O_1314,N_19959,N_19915);
xor UO_1315 (O_1315,N_19988,N_19837);
and UO_1316 (O_1316,N_19949,N_19845);
or UO_1317 (O_1317,N_19887,N_19880);
nand UO_1318 (O_1318,N_19844,N_19909);
xor UO_1319 (O_1319,N_19845,N_19937);
nand UO_1320 (O_1320,N_19905,N_19857);
or UO_1321 (O_1321,N_19973,N_19986);
nor UO_1322 (O_1322,N_19978,N_19868);
xnor UO_1323 (O_1323,N_19928,N_19811);
and UO_1324 (O_1324,N_19915,N_19961);
nor UO_1325 (O_1325,N_19835,N_19908);
or UO_1326 (O_1326,N_19974,N_19925);
and UO_1327 (O_1327,N_19950,N_19895);
and UO_1328 (O_1328,N_19952,N_19902);
and UO_1329 (O_1329,N_19946,N_19990);
or UO_1330 (O_1330,N_19861,N_19867);
or UO_1331 (O_1331,N_19872,N_19947);
or UO_1332 (O_1332,N_19916,N_19816);
xnor UO_1333 (O_1333,N_19957,N_19874);
or UO_1334 (O_1334,N_19857,N_19822);
and UO_1335 (O_1335,N_19953,N_19844);
or UO_1336 (O_1336,N_19873,N_19929);
nand UO_1337 (O_1337,N_19913,N_19816);
or UO_1338 (O_1338,N_19897,N_19946);
or UO_1339 (O_1339,N_19975,N_19971);
nand UO_1340 (O_1340,N_19949,N_19987);
or UO_1341 (O_1341,N_19849,N_19809);
or UO_1342 (O_1342,N_19970,N_19874);
and UO_1343 (O_1343,N_19965,N_19987);
or UO_1344 (O_1344,N_19856,N_19943);
nor UO_1345 (O_1345,N_19919,N_19951);
or UO_1346 (O_1346,N_19879,N_19832);
and UO_1347 (O_1347,N_19970,N_19956);
and UO_1348 (O_1348,N_19806,N_19800);
nor UO_1349 (O_1349,N_19918,N_19902);
and UO_1350 (O_1350,N_19881,N_19933);
nor UO_1351 (O_1351,N_19836,N_19901);
nor UO_1352 (O_1352,N_19876,N_19968);
and UO_1353 (O_1353,N_19899,N_19842);
and UO_1354 (O_1354,N_19862,N_19833);
xor UO_1355 (O_1355,N_19898,N_19953);
nand UO_1356 (O_1356,N_19824,N_19955);
and UO_1357 (O_1357,N_19904,N_19994);
nand UO_1358 (O_1358,N_19875,N_19974);
and UO_1359 (O_1359,N_19942,N_19964);
nor UO_1360 (O_1360,N_19925,N_19993);
and UO_1361 (O_1361,N_19841,N_19910);
xnor UO_1362 (O_1362,N_19847,N_19985);
and UO_1363 (O_1363,N_19898,N_19812);
nand UO_1364 (O_1364,N_19914,N_19814);
and UO_1365 (O_1365,N_19854,N_19908);
nand UO_1366 (O_1366,N_19986,N_19863);
and UO_1367 (O_1367,N_19883,N_19846);
nand UO_1368 (O_1368,N_19862,N_19858);
and UO_1369 (O_1369,N_19826,N_19980);
xor UO_1370 (O_1370,N_19946,N_19875);
and UO_1371 (O_1371,N_19966,N_19858);
or UO_1372 (O_1372,N_19886,N_19917);
or UO_1373 (O_1373,N_19842,N_19935);
and UO_1374 (O_1374,N_19884,N_19869);
nand UO_1375 (O_1375,N_19947,N_19806);
xnor UO_1376 (O_1376,N_19983,N_19996);
nand UO_1377 (O_1377,N_19967,N_19930);
or UO_1378 (O_1378,N_19836,N_19848);
and UO_1379 (O_1379,N_19872,N_19951);
nor UO_1380 (O_1380,N_19859,N_19960);
xor UO_1381 (O_1381,N_19961,N_19918);
xnor UO_1382 (O_1382,N_19824,N_19844);
and UO_1383 (O_1383,N_19969,N_19834);
nor UO_1384 (O_1384,N_19859,N_19823);
or UO_1385 (O_1385,N_19917,N_19904);
xnor UO_1386 (O_1386,N_19940,N_19819);
nor UO_1387 (O_1387,N_19853,N_19952);
nand UO_1388 (O_1388,N_19880,N_19879);
nor UO_1389 (O_1389,N_19949,N_19850);
or UO_1390 (O_1390,N_19863,N_19886);
or UO_1391 (O_1391,N_19825,N_19959);
xor UO_1392 (O_1392,N_19838,N_19915);
xnor UO_1393 (O_1393,N_19912,N_19878);
nand UO_1394 (O_1394,N_19891,N_19805);
and UO_1395 (O_1395,N_19969,N_19898);
or UO_1396 (O_1396,N_19908,N_19920);
and UO_1397 (O_1397,N_19826,N_19925);
nor UO_1398 (O_1398,N_19818,N_19991);
or UO_1399 (O_1399,N_19880,N_19892);
nand UO_1400 (O_1400,N_19893,N_19857);
nand UO_1401 (O_1401,N_19949,N_19961);
and UO_1402 (O_1402,N_19839,N_19854);
nand UO_1403 (O_1403,N_19832,N_19885);
xor UO_1404 (O_1404,N_19855,N_19802);
and UO_1405 (O_1405,N_19874,N_19908);
and UO_1406 (O_1406,N_19964,N_19982);
or UO_1407 (O_1407,N_19908,N_19941);
xnor UO_1408 (O_1408,N_19988,N_19843);
nor UO_1409 (O_1409,N_19943,N_19921);
xor UO_1410 (O_1410,N_19951,N_19900);
nor UO_1411 (O_1411,N_19833,N_19936);
nand UO_1412 (O_1412,N_19835,N_19970);
xnor UO_1413 (O_1413,N_19949,N_19871);
and UO_1414 (O_1414,N_19900,N_19947);
and UO_1415 (O_1415,N_19844,N_19969);
nand UO_1416 (O_1416,N_19830,N_19837);
xnor UO_1417 (O_1417,N_19953,N_19901);
nand UO_1418 (O_1418,N_19985,N_19820);
nor UO_1419 (O_1419,N_19992,N_19944);
and UO_1420 (O_1420,N_19821,N_19978);
or UO_1421 (O_1421,N_19947,N_19902);
nor UO_1422 (O_1422,N_19948,N_19893);
nor UO_1423 (O_1423,N_19842,N_19827);
xnor UO_1424 (O_1424,N_19916,N_19929);
nor UO_1425 (O_1425,N_19859,N_19879);
nand UO_1426 (O_1426,N_19920,N_19955);
or UO_1427 (O_1427,N_19812,N_19975);
and UO_1428 (O_1428,N_19982,N_19866);
nand UO_1429 (O_1429,N_19942,N_19844);
nor UO_1430 (O_1430,N_19848,N_19981);
or UO_1431 (O_1431,N_19989,N_19835);
nor UO_1432 (O_1432,N_19849,N_19967);
and UO_1433 (O_1433,N_19803,N_19880);
nand UO_1434 (O_1434,N_19810,N_19850);
nand UO_1435 (O_1435,N_19891,N_19914);
or UO_1436 (O_1436,N_19818,N_19802);
xor UO_1437 (O_1437,N_19896,N_19904);
nor UO_1438 (O_1438,N_19923,N_19823);
or UO_1439 (O_1439,N_19827,N_19921);
nand UO_1440 (O_1440,N_19902,N_19983);
xor UO_1441 (O_1441,N_19922,N_19850);
nor UO_1442 (O_1442,N_19923,N_19857);
nand UO_1443 (O_1443,N_19974,N_19955);
or UO_1444 (O_1444,N_19848,N_19942);
or UO_1445 (O_1445,N_19802,N_19847);
and UO_1446 (O_1446,N_19829,N_19983);
or UO_1447 (O_1447,N_19833,N_19840);
nor UO_1448 (O_1448,N_19863,N_19872);
xnor UO_1449 (O_1449,N_19931,N_19845);
or UO_1450 (O_1450,N_19920,N_19984);
and UO_1451 (O_1451,N_19848,N_19863);
nand UO_1452 (O_1452,N_19904,N_19817);
and UO_1453 (O_1453,N_19897,N_19900);
nand UO_1454 (O_1454,N_19889,N_19841);
and UO_1455 (O_1455,N_19886,N_19924);
or UO_1456 (O_1456,N_19815,N_19914);
nand UO_1457 (O_1457,N_19968,N_19957);
xor UO_1458 (O_1458,N_19807,N_19977);
nand UO_1459 (O_1459,N_19885,N_19950);
xnor UO_1460 (O_1460,N_19924,N_19877);
nand UO_1461 (O_1461,N_19936,N_19949);
and UO_1462 (O_1462,N_19987,N_19819);
and UO_1463 (O_1463,N_19862,N_19850);
and UO_1464 (O_1464,N_19978,N_19943);
nor UO_1465 (O_1465,N_19857,N_19888);
and UO_1466 (O_1466,N_19913,N_19823);
and UO_1467 (O_1467,N_19983,N_19843);
and UO_1468 (O_1468,N_19889,N_19965);
xnor UO_1469 (O_1469,N_19879,N_19863);
nor UO_1470 (O_1470,N_19996,N_19941);
or UO_1471 (O_1471,N_19890,N_19922);
xor UO_1472 (O_1472,N_19972,N_19897);
and UO_1473 (O_1473,N_19894,N_19890);
nor UO_1474 (O_1474,N_19811,N_19800);
or UO_1475 (O_1475,N_19829,N_19915);
or UO_1476 (O_1476,N_19981,N_19986);
xor UO_1477 (O_1477,N_19801,N_19950);
nand UO_1478 (O_1478,N_19944,N_19867);
nor UO_1479 (O_1479,N_19993,N_19931);
or UO_1480 (O_1480,N_19842,N_19976);
or UO_1481 (O_1481,N_19876,N_19857);
or UO_1482 (O_1482,N_19860,N_19909);
or UO_1483 (O_1483,N_19956,N_19901);
xor UO_1484 (O_1484,N_19946,N_19868);
or UO_1485 (O_1485,N_19979,N_19821);
nand UO_1486 (O_1486,N_19977,N_19971);
and UO_1487 (O_1487,N_19927,N_19957);
and UO_1488 (O_1488,N_19974,N_19819);
xor UO_1489 (O_1489,N_19870,N_19950);
nand UO_1490 (O_1490,N_19877,N_19888);
nor UO_1491 (O_1491,N_19955,N_19903);
xor UO_1492 (O_1492,N_19921,N_19933);
nand UO_1493 (O_1493,N_19850,N_19867);
nor UO_1494 (O_1494,N_19872,N_19808);
xnor UO_1495 (O_1495,N_19900,N_19935);
or UO_1496 (O_1496,N_19817,N_19924);
and UO_1497 (O_1497,N_19807,N_19859);
nor UO_1498 (O_1498,N_19972,N_19936);
and UO_1499 (O_1499,N_19840,N_19902);
nand UO_1500 (O_1500,N_19955,N_19843);
nor UO_1501 (O_1501,N_19944,N_19980);
nand UO_1502 (O_1502,N_19823,N_19996);
or UO_1503 (O_1503,N_19873,N_19928);
and UO_1504 (O_1504,N_19800,N_19847);
nor UO_1505 (O_1505,N_19972,N_19950);
nand UO_1506 (O_1506,N_19969,N_19835);
and UO_1507 (O_1507,N_19920,N_19902);
xor UO_1508 (O_1508,N_19863,N_19802);
xor UO_1509 (O_1509,N_19892,N_19963);
and UO_1510 (O_1510,N_19946,N_19882);
nand UO_1511 (O_1511,N_19812,N_19863);
or UO_1512 (O_1512,N_19937,N_19934);
nor UO_1513 (O_1513,N_19968,N_19921);
and UO_1514 (O_1514,N_19928,N_19985);
or UO_1515 (O_1515,N_19936,N_19897);
xnor UO_1516 (O_1516,N_19937,N_19978);
nor UO_1517 (O_1517,N_19983,N_19907);
and UO_1518 (O_1518,N_19912,N_19953);
and UO_1519 (O_1519,N_19854,N_19888);
xnor UO_1520 (O_1520,N_19894,N_19973);
and UO_1521 (O_1521,N_19802,N_19996);
xnor UO_1522 (O_1522,N_19971,N_19890);
nand UO_1523 (O_1523,N_19810,N_19889);
nand UO_1524 (O_1524,N_19987,N_19950);
xnor UO_1525 (O_1525,N_19852,N_19867);
nand UO_1526 (O_1526,N_19912,N_19962);
nand UO_1527 (O_1527,N_19919,N_19825);
nand UO_1528 (O_1528,N_19832,N_19858);
and UO_1529 (O_1529,N_19947,N_19876);
and UO_1530 (O_1530,N_19989,N_19913);
xor UO_1531 (O_1531,N_19892,N_19987);
and UO_1532 (O_1532,N_19924,N_19812);
nor UO_1533 (O_1533,N_19874,N_19969);
nand UO_1534 (O_1534,N_19877,N_19884);
xor UO_1535 (O_1535,N_19918,N_19907);
nor UO_1536 (O_1536,N_19982,N_19848);
or UO_1537 (O_1537,N_19955,N_19821);
nand UO_1538 (O_1538,N_19844,N_19920);
nor UO_1539 (O_1539,N_19853,N_19850);
nor UO_1540 (O_1540,N_19971,N_19951);
nand UO_1541 (O_1541,N_19817,N_19831);
or UO_1542 (O_1542,N_19942,N_19992);
and UO_1543 (O_1543,N_19833,N_19853);
nand UO_1544 (O_1544,N_19864,N_19943);
and UO_1545 (O_1545,N_19804,N_19801);
or UO_1546 (O_1546,N_19995,N_19872);
and UO_1547 (O_1547,N_19854,N_19921);
nand UO_1548 (O_1548,N_19902,N_19926);
nand UO_1549 (O_1549,N_19827,N_19800);
or UO_1550 (O_1550,N_19810,N_19922);
nor UO_1551 (O_1551,N_19984,N_19935);
or UO_1552 (O_1552,N_19865,N_19947);
or UO_1553 (O_1553,N_19975,N_19842);
or UO_1554 (O_1554,N_19942,N_19893);
nand UO_1555 (O_1555,N_19896,N_19969);
nand UO_1556 (O_1556,N_19946,N_19887);
xor UO_1557 (O_1557,N_19912,N_19947);
and UO_1558 (O_1558,N_19954,N_19915);
or UO_1559 (O_1559,N_19985,N_19923);
nand UO_1560 (O_1560,N_19916,N_19994);
nor UO_1561 (O_1561,N_19921,N_19832);
or UO_1562 (O_1562,N_19800,N_19924);
and UO_1563 (O_1563,N_19912,N_19822);
and UO_1564 (O_1564,N_19906,N_19917);
xnor UO_1565 (O_1565,N_19860,N_19990);
xor UO_1566 (O_1566,N_19874,N_19918);
and UO_1567 (O_1567,N_19907,N_19954);
nor UO_1568 (O_1568,N_19881,N_19951);
and UO_1569 (O_1569,N_19900,N_19861);
nand UO_1570 (O_1570,N_19888,N_19838);
nand UO_1571 (O_1571,N_19993,N_19978);
nor UO_1572 (O_1572,N_19982,N_19877);
and UO_1573 (O_1573,N_19983,N_19975);
nor UO_1574 (O_1574,N_19874,N_19875);
and UO_1575 (O_1575,N_19935,N_19879);
nor UO_1576 (O_1576,N_19831,N_19896);
and UO_1577 (O_1577,N_19877,N_19853);
nand UO_1578 (O_1578,N_19906,N_19855);
or UO_1579 (O_1579,N_19969,N_19973);
nor UO_1580 (O_1580,N_19994,N_19941);
nand UO_1581 (O_1581,N_19976,N_19824);
nor UO_1582 (O_1582,N_19822,N_19974);
nor UO_1583 (O_1583,N_19953,N_19978);
nand UO_1584 (O_1584,N_19871,N_19834);
xnor UO_1585 (O_1585,N_19882,N_19812);
nor UO_1586 (O_1586,N_19987,N_19904);
xnor UO_1587 (O_1587,N_19897,N_19937);
xor UO_1588 (O_1588,N_19892,N_19810);
and UO_1589 (O_1589,N_19981,N_19874);
nand UO_1590 (O_1590,N_19923,N_19832);
nand UO_1591 (O_1591,N_19966,N_19845);
and UO_1592 (O_1592,N_19871,N_19847);
nand UO_1593 (O_1593,N_19966,N_19830);
nand UO_1594 (O_1594,N_19995,N_19944);
or UO_1595 (O_1595,N_19881,N_19831);
xnor UO_1596 (O_1596,N_19946,N_19919);
nand UO_1597 (O_1597,N_19940,N_19886);
nor UO_1598 (O_1598,N_19986,N_19962);
nand UO_1599 (O_1599,N_19882,N_19950);
nor UO_1600 (O_1600,N_19894,N_19835);
xnor UO_1601 (O_1601,N_19882,N_19867);
or UO_1602 (O_1602,N_19947,N_19906);
or UO_1603 (O_1603,N_19901,N_19863);
nor UO_1604 (O_1604,N_19915,N_19810);
nor UO_1605 (O_1605,N_19920,N_19900);
and UO_1606 (O_1606,N_19820,N_19808);
nand UO_1607 (O_1607,N_19910,N_19898);
nor UO_1608 (O_1608,N_19882,N_19877);
and UO_1609 (O_1609,N_19935,N_19874);
or UO_1610 (O_1610,N_19991,N_19899);
and UO_1611 (O_1611,N_19867,N_19816);
xor UO_1612 (O_1612,N_19891,N_19837);
or UO_1613 (O_1613,N_19966,N_19834);
xor UO_1614 (O_1614,N_19856,N_19853);
nand UO_1615 (O_1615,N_19835,N_19834);
nor UO_1616 (O_1616,N_19917,N_19846);
nor UO_1617 (O_1617,N_19904,N_19855);
and UO_1618 (O_1618,N_19959,N_19987);
nor UO_1619 (O_1619,N_19947,N_19894);
and UO_1620 (O_1620,N_19917,N_19982);
nor UO_1621 (O_1621,N_19879,N_19851);
nand UO_1622 (O_1622,N_19803,N_19947);
nor UO_1623 (O_1623,N_19989,N_19859);
xor UO_1624 (O_1624,N_19814,N_19917);
or UO_1625 (O_1625,N_19823,N_19949);
or UO_1626 (O_1626,N_19896,N_19847);
xnor UO_1627 (O_1627,N_19935,N_19805);
nor UO_1628 (O_1628,N_19897,N_19962);
nor UO_1629 (O_1629,N_19816,N_19981);
xor UO_1630 (O_1630,N_19881,N_19970);
nor UO_1631 (O_1631,N_19817,N_19839);
and UO_1632 (O_1632,N_19929,N_19998);
nor UO_1633 (O_1633,N_19822,N_19992);
nand UO_1634 (O_1634,N_19869,N_19864);
nor UO_1635 (O_1635,N_19952,N_19874);
xnor UO_1636 (O_1636,N_19998,N_19873);
nand UO_1637 (O_1637,N_19875,N_19965);
nand UO_1638 (O_1638,N_19872,N_19817);
xnor UO_1639 (O_1639,N_19955,N_19980);
or UO_1640 (O_1640,N_19835,N_19899);
and UO_1641 (O_1641,N_19897,N_19923);
or UO_1642 (O_1642,N_19988,N_19808);
or UO_1643 (O_1643,N_19809,N_19834);
and UO_1644 (O_1644,N_19809,N_19804);
and UO_1645 (O_1645,N_19901,N_19917);
nor UO_1646 (O_1646,N_19884,N_19996);
nand UO_1647 (O_1647,N_19964,N_19988);
nand UO_1648 (O_1648,N_19812,N_19969);
nand UO_1649 (O_1649,N_19892,N_19936);
xnor UO_1650 (O_1650,N_19879,N_19842);
nor UO_1651 (O_1651,N_19961,N_19848);
or UO_1652 (O_1652,N_19821,N_19847);
nor UO_1653 (O_1653,N_19875,N_19811);
or UO_1654 (O_1654,N_19917,N_19973);
or UO_1655 (O_1655,N_19916,N_19838);
or UO_1656 (O_1656,N_19893,N_19985);
nand UO_1657 (O_1657,N_19875,N_19948);
or UO_1658 (O_1658,N_19939,N_19872);
nand UO_1659 (O_1659,N_19880,N_19976);
nor UO_1660 (O_1660,N_19923,N_19847);
nand UO_1661 (O_1661,N_19972,N_19911);
or UO_1662 (O_1662,N_19890,N_19966);
xor UO_1663 (O_1663,N_19832,N_19826);
nand UO_1664 (O_1664,N_19852,N_19822);
xnor UO_1665 (O_1665,N_19978,N_19819);
or UO_1666 (O_1666,N_19903,N_19820);
nand UO_1667 (O_1667,N_19923,N_19980);
nand UO_1668 (O_1668,N_19818,N_19812);
or UO_1669 (O_1669,N_19816,N_19943);
xor UO_1670 (O_1670,N_19814,N_19909);
nand UO_1671 (O_1671,N_19818,N_19923);
nor UO_1672 (O_1672,N_19922,N_19801);
or UO_1673 (O_1673,N_19940,N_19901);
nor UO_1674 (O_1674,N_19978,N_19870);
and UO_1675 (O_1675,N_19881,N_19914);
and UO_1676 (O_1676,N_19826,N_19856);
xnor UO_1677 (O_1677,N_19943,N_19965);
xor UO_1678 (O_1678,N_19988,N_19827);
nand UO_1679 (O_1679,N_19925,N_19996);
xnor UO_1680 (O_1680,N_19965,N_19994);
and UO_1681 (O_1681,N_19812,N_19973);
nor UO_1682 (O_1682,N_19955,N_19804);
and UO_1683 (O_1683,N_19919,N_19964);
nand UO_1684 (O_1684,N_19807,N_19888);
nor UO_1685 (O_1685,N_19813,N_19834);
and UO_1686 (O_1686,N_19858,N_19824);
xor UO_1687 (O_1687,N_19958,N_19804);
nor UO_1688 (O_1688,N_19812,N_19943);
nor UO_1689 (O_1689,N_19813,N_19904);
nor UO_1690 (O_1690,N_19972,N_19842);
nand UO_1691 (O_1691,N_19991,N_19800);
or UO_1692 (O_1692,N_19932,N_19957);
or UO_1693 (O_1693,N_19904,N_19963);
nor UO_1694 (O_1694,N_19902,N_19810);
nand UO_1695 (O_1695,N_19994,N_19804);
or UO_1696 (O_1696,N_19812,N_19890);
or UO_1697 (O_1697,N_19863,N_19989);
nand UO_1698 (O_1698,N_19844,N_19952);
xor UO_1699 (O_1699,N_19859,N_19864);
nor UO_1700 (O_1700,N_19886,N_19811);
or UO_1701 (O_1701,N_19831,N_19996);
xor UO_1702 (O_1702,N_19801,N_19888);
xnor UO_1703 (O_1703,N_19948,N_19876);
nor UO_1704 (O_1704,N_19889,N_19958);
nand UO_1705 (O_1705,N_19876,N_19822);
or UO_1706 (O_1706,N_19917,N_19810);
nor UO_1707 (O_1707,N_19988,N_19882);
nor UO_1708 (O_1708,N_19995,N_19951);
nand UO_1709 (O_1709,N_19938,N_19899);
and UO_1710 (O_1710,N_19988,N_19935);
or UO_1711 (O_1711,N_19868,N_19973);
or UO_1712 (O_1712,N_19889,N_19871);
xor UO_1713 (O_1713,N_19966,N_19906);
or UO_1714 (O_1714,N_19962,N_19958);
and UO_1715 (O_1715,N_19908,N_19919);
nor UO_1716 (O_1716,N_19936,N_19969);
xor UO_1717 (O_1717,N_19977,N_19886);
nor UO_1718 (O_1718,N_19829,N_19905);
nor UO_1719 (O_1719,N_19931,N_19934);
nor UO_1720 (O_1720,N_19872,N_19879);
and UO_1721 (O_1721,N_19927,N_19941);
nor UO_1722 (O_1722,N_19812,N_19902);
and UO_1723 (O_1723,N_19819,N_19976);
nand UO_1724 (O_1724,N_19949,N_19874);
or UO_1725 (O_1725,N_19861,N_19883);
or UO_1726 (O_1726,N_19917,N_19940);
nand UO_1727 (O_1727,N_19926,N_19863);
or UO_1728 (O_1728,N_19902,N_19816);
nor UO_1729 (O_1729,N_19996,N_19878);
xor UO_1730 (O_1730,N_19800,N_19834);
nand UO_1731 (O_1731,N_19972,N_19908);
xnor UO_1732 (O_1732,N_19805,N_19994);
or UO_1733 (O_1733,N_19887,N_19840);
nor UO_1734 (O_1734,N_19917,N_19971);
nor UO_1735 (O_1735,N_19997,N_19886);
nand UO_1736 (O_1736,N_19808,N_19975);
or UO_1737 (O_1737,N_19922,N_19965);
xnor UO_1738 (O_1738,N_19996,N_19891);
and UO_1739 (O_1739,N_19938,N_19869);
xor UO_1740 (O_1740,N_19857,N_19942);
nand UO_1741 (O_1741,N_19826,N_19870);
nand UO_1742 (O_1742,N_19969,N_19903);
nor UO_1743 (O_1743,N_19970,N_19993);
or UO_1744 (O_1744,N_19913,N_19937);
nor UO_1745 (O_1745,N_19903,N_19907);
xor UO_1746 (O_1746,N_19904,N_19905);
or UO_1747 (O_1747,N_19940,N_19842);
and UO_1748 (O_1748,N_19817,N_19979);
nand UO_1749 (O_1749,N_19870,N_19819);
nor UO_1750 (O_1750,N_19863,N_19969);
nor UO_1751 (O_1751,N_19821,N_19972);
or UO_1752 (O_1752,N_19907,N_19955);
or UO_1753 (O_1753,N_19825,N_19863);
or UO_1754 (O_1754,N_19925,N_19924);
or UO_1755 (O_1755,N_19861,N_19931);
nand UO_1756 (O_1756,N_19819,N_19880);
or UO_1757 (O_1757,N_19865,N_19911);
nor UO_1758 (O_1758,N_19831,N_19968);
nand UO_1759 (O_1759,N_19914,N_19900);
and UO_1760 (O_1760,N_19831,N_19982);
or UO_1761 (O_1761,N_19874,N_19844);
nor UO_1762 (O_1762,N_19866,N_19940);
or UO_1763 (O_1763,N_19996,N_19840);
nand UO_1764 (O_1764,N_19857,N_19930);
or UO_1765 (O_1765,N_19999,N_19888);
and UO_1766 (O_1766,N_19956,N_19973);
or UO_1767 (O_1767,N_19939,N_19968);
nor UO_1768 (O_1768,N_19923,N_19876);
or UO_1769 (O_1769,N_19983,N_19934);
nor UO_1770 (O_1770,N_19818,N_19955);
nand UO_1771 (O_1771,N_19880,N_19911);
nor UO_1772 (O_1772,N_19966,N_19832);
or UO_1773 (O_1773,N_19917,N_19893);
nand UO_1774 (O_1774,N_19916,N_19981);
and UO_1775 (O_1775,N_19930,N_19898);
nor UO_1776 (O_1776,N_19842,N_19991);
xnor UO_1777 (O_1777,N_19894,N_19887);
nor UO_1778 (O_1778,N_19964,N_19967);
xor UO_1779 (O_1779,N_19942,N_19966);
nor UO_1780 (O_1780,N_19824,N_19932);
and UO_1781 (O_1781,N_19884,N_19956);
xor UO_1782 (O_1782,N_19879,N_19839);
nand UO_1783 (O_1783,N_19870,N_19994);
nor UO_1784 (O_1784,N_19878,N_19906);
and UO_1785 (O_1785,N_19806,N_19938);
xnor UO_1786 (O_1786,N_19877,N_19932);
xnor UO_1787 (O_1787,N_19849,N_19932);
nand UO_1788 (O_1788,N_19875,N_19980);
xor UO_1789 (O_1789,N_19934,N_19841);
or UO_1790 (O_1790,N_19901,N_19908);
and UO_1791 (O_1791,N_19825,N_19946);
or UO_1792 (O_1792,N_19859,N_19999);
and UO_1793 (O_1793,N_19951,N_19962);
xnor UO_1794 (O_1794,N_19941,N_19854);
or UO_1795 (O_1795,N_19864,N_19851);
or UO_1796 (O_1796,N_19852,N_19830);
xnor UO_1797 (O_1797,N_19910,N_19991);
and UO_1798 (O_1798,N_19995,N_19962);
xor UO_1799 (O_1799,N_19889,N_19950);
nand UO_1800 (O_1800,N_19867,N_19935);
nor UO_1801 (O_1801,N_19955,N_19871);
nand UO_1802 (O_1802,N_19946,N_19916);
or UO_1803 (O_1803,N_19807,N_19994);
xnor UO_1804 (O_1804,N_19948,N_19823);
xor UO_1805 (O_1805,N_19848,N_19958);
and UO_1806 (O_1806,N_19844,N_19896);
and UO_1807 (O_1807,N_19963,N_19859);
or UO_1808 (O_1808,N_19838,N_19995);
nor UO_1809 (O_1809,N_19939,N_19898);
xnor UO_1810 (O_1810,N_19995,N_19812);
nor UO_1811 (O_1811,N_19859,N_19980);
xnor UO_1812 (O_1812,N_19980,N_19950);
or UO_1813 (O_1813,N_19994,N_19837);
and UO_1814 (O_1814,N_19861,N_19926);
or UO_1815 (O_1815,N_19846,N_19981);
nand UO_1816 (O_1816,N_19947,N_19960);
or UO_1817 (O_1817,N_19866,N_19891);
and UO_1818 (O_1818,N_19850,N_19840);
or UO_1819 (O_1819,N_19872,N_19926);
and UO_1820 (O_1820,N_19973,N_19944);
or UO_1821 (O_1821,N_19803,N_19932);
or UO_1822 (O_1822,N_19873,N_19950);
and UO_1823 (O_1823,N_19852,N_19847);
or UO_1824 (O_1824,N_19960,N_19924);
nand UO_1825 (O_1825,N_19931,N_19862);
or UO_1826 (O_1826,N_19975,N_19851);
or UO_1827 (O_1827,N_19815,N_19890);
xnor UO_1828 (O_1828,N_19946,N_19941);
and UO_1829 (O_1829,N_19970,N_19824);
xor UO_1830 (O_1830,N_19826,N_19992);
nand UO_1831 (O_1831,N_19945,N_19937);
nor UO_1832 (O_1832,N_19984,N_19804);
and UO_1833 (O_1833,N_19879,N_19966);
nand UO_1834 (O_1834,N_19957,N_19977);
nor UO_1835 (O_1835,N_19994,N_19877);
or UO_1836 (O_1836,N_19871,N_19829);
nand UO_1837 (O_1837,N_19811,N_19942);
and UO_1838 (O_1838,N_19942,N_19882);
nor UO_1839 (O_1839,N_19800,N_19888);
xnor UO_1840 (O_1840,N_19971,N_19802);
and UO_1841 (O_1841,N_19936,N_19864);
or UO_1842 (O_1842,N_19813,N_19917);
and UO_1843 (O_1843,N_19956,N_19845);
xnor UO_1844 (O_1844,N_19957,N_19851);
xnor UO_1845 (O_1845,N_19908,N_19831);
and UO_1846 (O_1846,N_19882,N_19939);
or UO_1847 (O_1847,N_19821,N_19939);
nor UO_1848 (O_1848,N_19892,N_19877);
or UO_1849 (O_1849,N_19858,N_19820);
xor UO_1850 (O_1850,N_19886,N_19850);
xnor UO_1851 (O_1851,N_19906,N_19957);
xnor UO_1852 (O_1852,N_19889,N_19816);
and UO_1853 (O_1853,N_19916,N_19868);
nand UO_1854 (O_1854,N_19949,N_19885);
and UO_1855 (O_1855,N_19812,N_19927);
nor UO_1856 (O_1856,N_19953,N_19995);
or UO_1857 (O_1857,N_19807,N_19931);
nor UO_1858 (O_1858,N_19919,N_19872);
or UO_1859 (O_1859,N_19962,N_19867);
xor UO_1860 (O_1860,N_19906,N_19973);
and UO_1861 (O_1861,N_19846,N_19970);
nand UO_1862 (O_1862,N_19893,N_19972);
and UO_1863 (O_1863,N_19951,N_19877);
nand UO_1864 (O_1864,N_19934,N_19818);
xor UO_1865 (O_1865,N_19901,N_19989);
or UO_1866 (O_1866,N_19982,N_19815);
nor UO_1867 (O_1867,N_19819,N_19912);
nand UO_1868 (O_1868,N_19840,N_19818);
nor UO_1869 (O_1869,N_19947,N_19891);
or UO_1870 (O_1870,N_19818,N_19984);
nand UO_1871 (O_1871,N_19954,N_19976);
and UO_1872 (O_1872,N_19994,N_19981);
nand UO_1873 (O_1873,N_19802,N_19872);
xor UO_1874 (O_1874,N_19871,N_19868);
or UO_1875 (O_1875,N_19899,N_19869);
or UO_1876 (O_1876,N_19890,N_19849);
nor UO_1877 (O_1877,N_19900,N_19865);
nand UO_1878 (O_1878,N_19866,N_19822);
nand UO_1879 (O_1879,N_19910,N_19916);
and UO_1880 (O_1880,N_19877,N_19942);
nor UO_1881 (O_1881,N_19904,N_19995);
xor UO_1882 (O_1882,N_19886,N_19879);
nand UO_1883 (O_1883,N_19814,N_19998);
and UO_1884 (O_1884,N_19901,N_19838);
nand UO_1885 (O_1885,N_19877,N_19855);
and UO_1886 (O_1886,N_19807,N_19926);
nor UO_1887 (O_1887,N_19872,N_19897);
xnor UO_1888 (O_1888,N_19857,N_19950);
xor UO_1889 (O_1889,N_19852,N_19988);
or UO_1890 (O_1890,N_19846,N_19983);
or UO_1891 (O_1891,N_19804,N_19906);
xnor UO_1892 (O_1892,N_19917,N_19935);
xor UO_1893 (O_1893,N_19858,N_19850);
xor UO_1894 (O_1894,N_19858,N_19994);
or UO_1895 (O_1895,N_19861,N_19842);
and UO_1896 (O_1896,N_19905,N_19895);
nand UO_1897 (O_1897,N_19973,N_19820);
xnor UO_1898 (O_1898,N_19962,N_19916);
nor UO_1899 (O_1899,N_19964,N_19882);
xor UO_1900 (O_1900,N_19911,N_19943);
xnor UO_1901 (O_1901,N_19968,N_19863);
or UO_1902 (O_1902,N_19860,N_19952);
and UO_1903 (O_1903,N_19826,N_19930);
xnor UO_1904 (O_1904,N_19955,N_19989);
or UO_1905 (O_1905,N_19929,N_19995);
and UO_1906 (O_1906,N_19999,N_19925);
nor UO_1907 (O_1907,N_19915,N_19845);
or UO_1908 (O_1908,N_19838,N_19991);
nor UO_1909 (O_1909,N_19997,N_19854);
or UO_1910 (O_1910,N_19846,N_19986);
nand UO_1911 (O_1911,N_19882,N_19927);
and UO_1912 (O_1912,N_19900,N_19874);
xor UO_1913 (O_1913,N_19925,N_19872);
xor UO_1914 (O_1914,N_19837,N_19920);
nand UO_1915 (O_1915,N_19818,N_19860);
nand UO_1916 (O_1916,N_19872,N_19920);
and UO_1917 (O_1917,N_19999,N_19889);
or UO_1918 (O_1918,N_19904,N_19833);
nand UO_1919 (O_1919,N_19900,N_19849);
and UO_1920 (O_1920,N_19868,N_19992);
nor UO_1921 (O_1921,N_19891,N_19941);
or UO_1922 (O_1922,N_19943,N_19979);
or UO_1923 (O_1923,N_19931,N_19943);
or UO_1924 (O_1924,N_19985,N_19887);
or UO_1925 (O_1925,N_19808,N_19885);
and UO_1926 (O_1926,N_19986,N_19960);
nand UO_1927 (O_1927,N_19834,N_19882);
or UO_1928 (O_1928,N_19976,N_19995);
nand UO_1929 (O_1929,N_19835,N_19975);
xor UO_1930 (O_1930,N_19849,N_19889);
nor UO_1931 (O_1931,N_19873,N_19982);
or UO_1932 (O_1932,N_19912,N_19825);
and UO_1933 (O_1933,N_19961,N_19975);
nand UO_1934 (O_1934,N_19976,N_19895);
xnor UO_1935 (O_1935,N_19970,N_19815);
nand UO_1936 (O_1936,N_19873,N_19952);
nand UO_1937 (O_1937,N_19939,N_19873);
nand UO_1938 (O_1938,N_19855,N_19925);
nand UO_1939 (O_1939,N_19945,N_19934);
or UO_1940 (O_1940,N_19825,N_19993);
and UO_1941 (O_1941,N_19979,N_19924);
xnor UO_1942 (O_1942,N_19883,N_19842);
nand UO_1943 (O_1943,N_19948,N_19901);
xor UO_1944 (O_1944,N_19955,N_19962);
nand UO_1945 (O_1945,N_19956,N_19824);
or UO_1946 (O_1946,N_19919,N_19978);
and UO_1947 (O_1947,N_19913,N_19959);
xor UO_1948 (O_1948,N_19807,N_19987);
nand UO_1949 (O_1949,N_19809,N_19893);
xnor UO_1950 (O_1950,N_19909,N_19827);
nor UO_1951 (O_1951,N_19980,N_19920);
xor UO_1952 (O_1952,N_19982,N_19859);
or UO_1953 (O_1953,N_19803,N_19841);
or UO_1954 (O_1954,N_19975,N_19904);
xnor UO_1955 (O_1955,N_19975,N_19807);
and UO_1956 (O_1956,N_19899,N_19908);
and UO_1957 (O_1957,N_19893,N_19876);
or UO_1958 (O_1958,N_19869,N_19815);
nand UO_1959 (O_1959,N_19898,N_19954);
nor UO_1960 (O_1960,N_19863,N_19990);
nor UO_1961 (O_1961,N_19841,N_19921);
xor UO_1962 (O_1962,N_19892,N_19903);
and UO_1963 (O_1963,N_19889,N_19986);
nand UO_1964 (O_1964,N_19867,N_19802);
xor UO_1965 (O_1965,N_19960,N_19806);
or UO_1966 (O_1966,N_19886,N_19836);
or UO_1967 (O_1967,N_19825,N_19849);
or UO_1968 (O_1968,N_19956,N_19892);
or UO_1969 (O_1969,N_19997,N_19972);
nor UO_1970 (O_1970,N_19819,N_19900);
xor UO_1971 (O_1971,N_19931,N_19910);
nor UO_1972 (O_1972,N_19926,N_19854);
xnor UO_1973 (O_1973,N_19813,N_19972);
and UO_1974 (O_1974,N_19881,N_19864);
nand UO_1975 (O_1975,N_19958,N_19908);
or UO_1976 (O_1976,N_19979,N_19938);
xnor UO_1977 (O_1977,N_19916,N_19928);
xor UO_1978 (O_1978,N_19905,N_19803);
or UO_1979 (O_1979,N_19920,N_19833);
xor UO_1980 (O_1980,N_19977,N_19882);
or UO_1981 (O_1981,N_19955,N_19805);
nand UO_1982 (O_1982,N_19861,N_19906);
nor UO_1983 (O_1983,N_19905,N_19902);
xnor UO_1984 (O_1984,N_19905,N_19969);
or UO_1985 (O_1985,N_19831,N_19927);
nor UO_1986 (O_1986,N_19915,N_19849);
nor UO_1987 (O_1987,N_19898,N_19839);
and UO_1988 (O_1988,N_19894,N_19980);
nor UO_1989 (O_1989,N_19905,N_19937);
nor UO_1990 (O_1990,N_19817,N_19967);
and UO_1991 (O_1991,N_19823,N_19938);
xor UO_1992 (O_1992,N_19889,N_19913);
nand UO_1993 (O_1993,N_19837,N_19842);
nand UO_1994 (O_1994,N_19969,N_19867);
xnor UO_1995 (O_1995,N_19876,N_19940);
and UO_1996 (O_1996,N_19964,N_19974);
nor UO_1997 (O_1997,N_19981,N_19894);
and UO_1998 (O_1998,N_19953,N_19812);
and UO_1999 (O_1999,N_19882,N_19975);
or UO_2000 (O_2000,N_19816,N_19979);
and UO_2001 (O_2001,N_19864,N_19822);
and UO_2002 (O_2002,N_19827,N_19936);
xor UO_2003 (O_2003,N_19944,N_19866);
or UO_2004 (O_2004,N_19871,N_19947);
and UO_2005 (O_2005,N_19986,N_19860);
nor UO_2006 (O_2006,N_19952,N_19839);
nor UO_2007 (O_2007,N_19942,N_19821);
nand UO_2008 (O_2008,N_19954,N_19977);
nand UO_2009 (O_2009,N_19862,N_19933);
nand UO_2010 (O_2010,N_19835,N_19985);
nor UO_2011 (O_2011,N_19848,N_19898);
nor UO_2012 (O_2012,N_19909,N_19899);
or UO_2013 (O_2013,N_19859,N_19968);
and UO_2014 (O_2014,N_19853,N_19838);
nand UO_2015 (O_2015,N_19917,N_19969);
and UO_2016 (O_2016,N_19956,N_19833);
or UO_2017 (O_2017,N_19925,N_19899);
nand UO_2018 (O_2018,N_19837,N_19996);
nor UO_2019 (O_2019,N_19820,N_19824);
nor UO_2020 (O_2020,N_19872,N_19963);
and UO_2021 (O_2021,N_19833,N_19875);
nor UO_2022 (O_2022,N_19892,N_19984);
and UO_2023 (O_2023,N_19899,N_19937);
nor UO_2024 (O_2024,N_19962,N_19800);
and UO_2025 (O_2025,N_19923,N_19962);
and UO_2026 (O_2026,N_19917,N_19995);
nor UO_2027 (O_2027,N_19936,N_19922);
or UO_2028 (O_2028,N_19965,N_19961);
nor UO_2029 (O_2029,N_19856,N_19809);
or UO_2030 (O_2030,N_19966,N_19835);
xor UO_2031 (O_2031,N_19950,N_19877);
and UO_2032 (O_2032,N_19928,N_19874);
or UO_2033 (O_2033,N_19980,N_19800);
and UO_2034 (O_2034,N_19821,N_19961);
nand UO_2035 (O_2035,N_19861,N_19890);
nand UO_2036 (O_2036,N_19967,N_19981);
xor UO_2037 (O_2037,N_19878,N_19934);
or UO_2038 (O_2038,N_19954,N_19960);
and UO_2039 (O_2039,N_19866,N_19850);
nand UO_2040 (O_2040,N_19975,N_19846);
nor UO_2041 (O_2041,N_19909,N_19936);
or UO_2042 (O_2042,N_19956,N_19930);
nand UO_2043 (O_2043,N_19932,N_19942);
or UO_2044 (O_2044,N_19871,N_19819);
nor UO_2045 (O_2045,N_19965,N_19829);
xor UO_2046 (O_2046,N_19822,N_19869);
or UO_2047 (O_2047,N_19958,N_19910);
nand UO_2048 (O_2048,N_19947,N_19953);
xnor UO_2049 (O_2049,N_19950,N_19829);
nand UO_2050 (O_2050,N_19866,N_19856);
nor UO_2051 (O_2051,N_19933,N_19882);
nor UO_2052 (O_2052,N_19859,N_19858);
xnor UO_2053 (O_2053,N_19997,N_19872);
or UO_2054 (O_2054,N_19842,N_19871);
nor UO_2055 (O_2055,N_19964,N_19874);
or UO_2056 (O_2056,N_19927,N_19817);
xnor UO_2057 (O_2057,N_19877,N_19805);
nand UO_2058 (O_2058,N_19912,N_19986);
or UO_2059 (O_2059,N_19941,N_19841);
nor UO_2060 (O_2060,N_19975,N_19929);
xor UO_2061 (O_2061,N_19917,N_19945);
and UO_2062 (O_2062,N_19884,N_19965);
and UO_2063 (O_2063,N_19833,N_19894);
nor UO_2064 (O_2064,N_19929,N_19985);
and UO_2065 (O_2065,N_19839,N_19943);
xnor UO_2066 (O_2066,N_19901,N_19859);
nand UO_2067 (O_2067,N_19896,N_19880);
nand UO_2068 (O_2068,N_19840,N_19988);
and UO_2069 (O_2069,N_19927,N_19884);
xnor UO_2070 (O_2070,N_19834,N_19894);
or UO_2071 (O_2071,N_19812,N_19895);
and UO_2072 (O_2072,N_19838,N_19835);
and UO_2073 (O_2073,N_19907,N_19806);
nand UO_2074 (O_2074,N_19935,N_19876);
nand UO_2075 (O_2075,N_19888,N_19930);
nor UO_2076 (O_2076,N_19902,N_19949);
nor UO_2077 (O_2077,N_19929,N_19855);
or UO_2078 (O_2078,N_19943,N_19883);
nand UO_2079 (O_2079,N_19957,N_19870);
nor UO_2080 (O_2080,N_19944,N_19862);
or UO_2081 (O_2081,N_19826,N_19905);
xor UO_2082 (O_2082,N_19886,N_19854);
and UO_2083 (O_2083,N_19846,N_19833);
nand UO_2084 (O_2084,N_19973,N_19908);
nor UO_2085 (O_2085,N_19839,N_19876);
nand UO_2086 (O_2086,N_19815,N_19983);
and UO_2087 (O_2087,N_19963,N_19825);
xnor UO_2088 (O_2088,N_19911,N_19853);
and UO_2089 (O_2089,N_19879,N_19985);
or UO_2090 (O_2090,N_19852,N_19934);
and UO_2091 (O_2091,N_19883,N_19927);
and UO_2092 (O_2092,N_19914,N_19838);
nor UO_2093 (O_2093,N_19888,N_19927);
nand UO_2094 (O_2094,N_19885,N_19998);
and UO_2095 (O_2095,N_19811,N_19914);
nand UO_2096 (O_2096,N_19907,N_19935);
and UO_2097 (O_2097,N_19920,N_19994);
and UO_2098 (O_2098,N_19988,N_19841);
nand UO_2099 (O_2099,N_19986,N_19990);
nand UO_2100 (O_2100,N_19817,N_19933);
nand UO_2101 (O_2101,N_19838,N_19804);
or UO_2102 (O_2102,N_19969,N_19839);
nor UO_2103 (O_2103,N_19970,N_19817);
xor UO_2104 (O_2104,N_19916,N_19821);
nand UO_2105 (O_2105,N_19844,N_19922);
nand UO_2106 (O_2106,N_19884,N_19845);
xor UO_2107 (O_2107,N_19823,N_19914);
xor UO_2108 (O_2108,N_19942,N_19908);
nand UO_2109 (O_2109,N_19800,N_19860);
xnor UO_2110 (O_2110,N_19834,N_19845);
nor UO_2111 (O_2111,N_19935,N_19956);
or UO_2112 (O_2112,N_19989,N_19927);
nand UO_2113 (O_2113,N_19902,N_19841);
nand UO_2114 (O_2114,N_19841,N_19964);
xor UO_2115 (O_2115,N_19838,N_19869);
nand UO_2116 (O_2116,N_19915,N_19988);
nor UO_2117 (O_2117,N_19932,N_19992);
nor UO_2118 (O_2118,N_19880,N_19845);
and UO_2119 (O_2119,N_19873,N_19825);
xnor UO_2120 (O_2120,N_19807,N_19836);
nor UO_2121 (O_2121,N_19979,N_19915);
or UO_2122 (O_2122,N_19837,N_19983);
nor UO_2123 (O_2123,N_19949,N_19957);
or UO_2124 (O_2124,N_19966,N_19840);
nand UO_2125 (O_2125,N_19966,N_19994);
and UO_2126 (O_2126,N_19960,N_19879);
and UO_2127 (O_2127,N_19819,N_19872);
nand UO_2128 (O_2128,N_19872,N_19836);
xnor UO_2129 (O_2129,N_19835,N_19968);
or UO_2130 (O_2130,N_19830,N_19851);
or UO_2131 (O_2131,N_19977,N_19904);
xor UO_2132 (O_2132,N_19932,N_19946);
and UO_2133 (O_2133,N_19888,N_19973);
xor UO_2134 (O_2134,N_19951,N_19861);
or UO_2135 (O_2135,N_19920,N_19979);
and UO_2136 (O_2136,N_19884,N_19828);
nand UO_2137 (O_2137,N_19999,N_19839);
xnor UO_2138 (O_2138,N_19995,N_19991);
nand UO_2139 (O_2139,N_19967,N_19815);
or UO_2140 (O_2140,N_19874,N_19838);
nand UO_2141 (O_2141,N_19870,N_19845);
nand UO_2142 (O_2142,N_19953,N_19811);
nand UO_2143 (O_2143,N_19947,N_19832);
and UO_2144 (O_2144,N_19848,N_19912);
nand UO_2145 (O_2145,N_19965,N_19958);
and UO_2146 (O_2146,N_19968,N_19824);
nor UO_2147 (O_2147,N_19926,N_19987);
nand UO_2148 (O_2148,N_19863,N_19842);
xnor UO_2149 (O_2149,N_19802,N_19820);
or UO_2150 (O_2150,N_19985,N_19960);
or UO_2151 (O_2151,N_19966,N_19863);
xor UO_2152 (O_2152,N_19951,N_19869);
or UO_2153 (O_2153,N_19952,N_19885);
and UO_2154 (O_2154,N_19917,N_19989);
nor UO_2155 (O_2155,N_19918,N_19885);
or UO_2156 (O_2156,N_19829,N_19945);
or UO_2157 (O_2157,N_19987,N_19911);
nor UO_2158 (O_2158,N_19944,N_19859);
nand UO_2159 (O_2159,N_19806,N_19834);
nor UO_2160 (O_2160,N_19959,N_19927);
xnor UO_2161 (O_2161,N_19814,N_19801);
or UO_2162 (O_2162,N_19924,N_19884);
xor UO_2163 (O_2163,N_19879,N_19924);
and UO_2164 (O_2164,N_19813,N_19853);
nor UO_2165 (O_2165,N_19988,N_19884);
xor UO_2166 (O_2166,N_19824,N_19943);
nand UO_2167 (O_2167,N_19928,N_19866);
nor UO_2168 (O_2168,N_19891,N_19998);
nor UO_2169 (O_2169,N_19832,N_19800);
and UO_2170 (O_2170,N_19923,N_19957);
xor UO_2171 (O_2171,N_19806,N_19944);
nor UO_2172 (O_2172,N_19836,N_19928);
or UO_2173 (O_2173,N_19924,N_19851);
or UO_2174 (O_2174,N_19809,N_19954);
nand UO_2175 (O_2175,N_19940,N_19879);
or UO_2176 (O_2176,N_19853,N_19984);
nor UO_2177 (O_2177,N_19887,N_19876);
xor UO_2178 (O_2178,N_19919,N_19971);
or UO_2179 (O_2179,N_19891,N_19911);
and UO_2180 (O_2180,N_19891,N_19979);
xor UO_2181 (O_2181,N_19965,N_19806);
and UO_2182 (O_2182,N_19820,N_19827);
and UO_2183 (O_2183,N_19984,N_19936);
nand UO_2184 (O_2184,N_19872,N_19885);
nand UO_2185 (O_2185,N_19989,N_19979);
nand UO_2186 (O_2186,N_19975,N_19836);
and UO_2187 (O_2187,N_19951,N_19994);
nand UO_2188 (O_2188,N_19876,N_19816);
or UO_2189 (O_2189,N_19912,N_19866);
or UO_2190 (O_2190,N_19814,N_19830);
and UO_2191 (O_2191,N_19994,N_19847);
and UO_2192 (O_2192,N_19819,N_19932);
nor UO_2193 (O_2193,N_19973,N_19920);
xnor UO_2194 (O_2194,N_19839,N_19924);
or UO_2195 (O_2195,N_19900,N_19999);
and UO_2196 (O_2196,N_19862,N_19874);
and UO_2197 (O_2197,N_19973,N_19895);
nand UO_2198 (O_2198,N_19910,N_19950);
xor UO_2199 (O_2199,N_19892,N_19951);
xnor UO_2200 (O_2200,N_19984,N_19959);
or UO_2201 (O_2201,N_19901,N_19951);
nor UO_2202 (O_2202,N_19834,N_19942);
nor UO_2203 (O_2203,N_19957,N_19871);
nor UO_2204 (O_2204,N_19864,N_19807);
nor UO_2205 (O_2205,N_19892,N_19832);
or UO_2206 (O_2206,N_19837,N_19889);
or UO_2207 (O_2207,N_19818,N_19899);
xor UO_2208 (O_2208,N_19950,N_19959);
nand UO_2209 (O_2209,N_19922,N_19967);
nand UO_2210 (O_2210,N_19911,N_19825);
or UO_2211 (O_2211,N_19940,N_19881);
or UO_2212 (O_2212,N_19816,N_19896);
nor UO_2213 (O_2213,N_19898,N_19915);
or UO_2214 (O_2214,N_19964,N_19941);
and UO_2215 (O_2215,N_19826,N_19974);
nor UO_2216 (O_2216,N_19843,N_19979);
nor UO_2217 (O_2217,N_19915,N_19891);
or UO_2218 (O_2218,N_19930,N_19927);
nand UO_2219 (O_2219,N_19819,N_19875);
nor UO_2220 (O_2220,N_19989,N_19962);
and UO_2221 (O_2221,N_19977,N_19966);
xnor UO_2222 (O_2222,N_19882,N_19951);
and UO_2223 (O_2223,N_19846,N_19831);
or UO_2224 (O_2224,N_19825,N_19859);
and UO_2225 (O_2225,N_19899,N_19801);
or UO_2226 (O_2226,N_19934,N_19890);
and UO_2227 (O_2227,N_19873,N_19860);
and UO_2228 (O_2228,N_19977,N_19963);
nor UO_2229 (O_2229,N_19924,N_19935);
or UO_2230 (O_2230,N_19821,N_19835);
xor UO_2231 (O_2231,N_19878,N_19829);
nor UO_2232 (O_2232,N_19807,N_19849);
and UO_2233 (O_2233,N_19989,N_19941);
or UO_2234 (O_2234,N_19815,N_19843);
xor UO_2235 (O_2235,N_19929,N_19913);
nor UO_2236 (O_2236,N_19916,N_19806);
nand UO_2237 (O_2237,N_19904,N_19831);
nand UO_2238 (O_2238,N_19956,N_19859);
nor UO_2239 (O_2239,N_19895,N_19838);
xor UO_2240 (O_2240,N_19924,N_19801);
nand UO_2241 (O_2241,N_19920,N_19986);
or UO_2242 (O_2242,N_19871,N_19855);
nand UO_2243 (O_2243,N_19932,N_19887);
or UO_2244 (O_2244,N_19910,N_19827);
xor UO_2245 (O_2245,N_19924,N_19936);
or UO_2246 (O_2246,N_19993,N_19844);
and UO_2247 (O_2247,N_19896,N_19952);
or UO_2248 (O_2248,N_19859,N_19838);
nand UO_2249 (O_2249,N_19987,N_19997);
or UO_2250 (O_2250,N_19800,N_19973);
nor UO_2251 (O_2251,N_19851,N_19943);
nand UO_2252 (O_2252,N_19813,N_19900);
or UO_2253 (O_2253,N_19966,N_19892);
nor UO_2254 (O_2254,N_19815,N_19818);
xor UO_2255 (O_2255,N_19976,N_19843);
and UO_2256 (O_2256,N_19808,N_19843);
nor UO_2257 (O_2257,N_19841,N_19872);
nand UO_2258 (O_2258,N_19958,N_19920);
and UO_2259 (O_2259,N_19864,N_19906);
nor UO_2260 (O_2260,N_19875,N_19977);
xnor UO_2261 (O_2261,N_19924,N_19835);
xor UO_2262 (O_2262,N_19808,N_19973);
or UO_2263 (O_2263,N_19975,N_19936);
and UO_2264 (O_2264,N_19919,N_19960);
or UO_2265 (O_2265,N_19875,N_19914);
nor UO_2266 (O_2266,N_19924,N_19926);
or UO_2267 (O_2267,N_19995,N_19910);
nor UO_2268 (O_2268,N_19924,N_19808);
and UO_2269 (O_2269,N_19904,N_19862);
and UO_2270 (O_2270,N_19866,N_19816);
nand UO_2271 (O_2271,N_19995,N_19920);
or UO_2272 (O_2272,N_19843,N_19825);
xor UO_2273 (O_2273,N_19954,N_19938);
or UO_2274 (O_2274,N_19881,N_19867);
or UO_2275 (O_2275,N_19808,N_19853);
xnor UO_2276 (O_2276,N_19967,N_19812);
or UO_2277 (O_2277,N_19909,N_19867);
nand UO_2278 (O_2278,N_19880,N_19863);
xor UO_2279 (O_2279,N_19922,N_19886);
or UO_2280 (O_2280,N_19898,N_19919);
nor UO_2281 (O_2281,N_19837,N_19928);
and UO_2282 (O_2282,N_19878,N_19845);
nand UO_2283 (O_2283,N_19897,N_19905);
xor UO_2284 (O_2284,N_19945,N_19978);
nand UO_2285 (O_2285,N_19937,N_19865);
nor UO_2286 (O_2286,N_19929,N_19947);
and UO_2287 (O_2287,N_19905,N_19953);
nand UO_2288 (O_2288,N_19890,N_19800);
xnor UO_2289 (O_2289,N_19993,N_19817);
nand UO_2290 (O_2290,N_19899,N_19952);
and UO_2291 (O_2291,N_19865,N_19969);
nand UO_2292 (O_2292,N_19907,N_19970);
nand UO_2293 (O_2293,N_19874,N_19833);
or UO_2294 (O_2294,N_19997,N_19802);
or UO_2295 (O_2295,N_19867,N_19875);
xnor UO_2296 (O_2296,N_19818,N_19875);
nor UO_2297 (O_2297,N_19895,N_19826);
nor UO_2298 (O_2298,N_19917,N_19932);
or UO_2299 (O_2299,N_19892,N_19994);
nor UO_2300 (O_2300,N_19879,N_19954);
xor UO_2301 (O_2301,N_19926,N_19953);
nor UO_2302 (O_2302,N_19846,N_19899);
nand UO_2303 (O_2303,N_19824,N_19874);
or UO_2304 (O_2304,N_19956,N_19826);
nand UO_2305 (O_2305,N_19942,N_19955);
nand UO_2306 (O_2306,N_19926,N_19803);
or UO_2307 (O_2307,N_19889,N_19856);
and UO_2308 (O_2308,N_19909,N_19857);
or UO_2309 (O_2309,N_19935,N_19986);
nor UO_2310 (O_2310,N_19853,N_19954);
nand UO_2311 (O_2311,N_19958,N_19914);
nor UO_2312 (O_2312,N_19885,N_19981);
xor UO_2313 (O_2313,N_19889,N_19834);
and UO_2314 (O_2314,N_19978,N_19928);
or UO_2315 (O_2315,N_19855,N_19887);
nand UO_2316 (O_2316,N_19827,N_19850);
nor UO_2317 (O_2317,N_19935,N_19810);
and UO_2318 (O_2318,N_19848,N_19930);
nand UO_2319 (O_2319,N_19920,N_19985);
nor UO_2320 (O_2320,N_19833,N_19897);
nor UO_2321 (O_2321,N_19827,N_19816);
xor UO_2322 (O_2322,N_19952,N_19898);
or UO_2323 (O_2323,N_19924,N_19904);
or UO_2324 (O_2324,N_19946,N_19970);
xnor UO_2325 (O_2325,N_19841,N_19850);
and UO_2326 (O_2326,N_19808,N_19932);
and UO_2327 (O_2327,N_19913,N_19870);
or UO_2328 (O_2328,N_19859,N_19936);
or UO_2329 (O_2329,N_19915,N_19913);
and UO_2330 (O_2330,N_19844,N_19892);
nand UO_2331 (O_2331,N_19978,N_19926);
nor UO_2332 (O_2332,N_19829,N_19933);
xnor UO_2333 (O_2333,N_19879,N_19848);
xnor UO_2334 (O_2334,N_19991,N_19972);
nand UO_2335 (O_2335,N_19841,N_19924);
or UO_2336 (O_2336,N_19899,N_19886);
xnor UO_2337 (O_2337,N_19878,N_19855);
and UO_2338 (O_2338,N_19965,N_19877);
and UO_2339 (O_2339,N_19880,N_19983);
nand UO_2340 (O_2340,N_19886,N_19972);
nand UO_2341 (O_2341,N_19830,N_19863);
or UO_2342 (O_2342,N_19943,N_19842);
nand UO_2343 (O_2343,N_19966,N_19993);
or UO_2344 (O_2344,N_19820,N_19914);
xor UO_2345 (O_2345,N_19989,N_19825);
nand UO_2346 (O_2346,N_19963,N_19889);
xnor UO_2347 (O_2347,N_19920,N_19953);
nor UO_2348 (O_2348,N_19835,N_19918);
nor UO_2349 (O_2349,N_19832,N_19851);
xnor UO_2350 (O_2350,N_19876,N_19837);
nor UO_2351 (O_2351,N_19886,N_19964);
xor UO_2352 (O_2352,N_19838,N_19896);
or UO_2353 (O_2353,N_19823,N_19821);
or UO_2354 (O_2354,N_19965,N_19896);
xnor UO_2355 (O_2355,N_19893,N_19937);
and UO_2356 (O_2356,N_19959,N_19831);
or UO_2357 (O_2357,N_19881,N_19921);
nand UO_2358 (O_2358,N_19868,N_19809);
and UO_2359 (O_2359,N_19867,N_19895);
xnor UO_2360 (O_2360,N_19971,N_19938);
nand UO_2361 (O_2361,N_19952,N_19919);
nor UO_2362 (O_2362,N_19864,N_19998);
and UO_2363 (O_2363,N_19855,N_19813);
xnor UO_2364 (O_2364,N_19832,N_19864);
nand UO_2365 (O_2365,N_19839,N_19931);
nand UO_2366 (O_2366,N_19977,N_19921);
or UO_2367 (O_2367,N_19962,N_19895);
xor UO_2368 (O_2368,N_19985,N_19828);
and UO_2369 (O_2369,N_19952,N_19909);
xnor UO_2370 (O_2370,N_19885,N_19890);
xnor UO_2371 (O_2371,N_19960,N_19996);
xnor UO_2372 (O_2372,N_19862,N_19811);
or UO_2373 (O_2373,N_19934,N_19822);
xnor UO_2374 (O_2374,N_19999,N_19845);
nand UO_2375 (O_2375,N_19803,N_19822);
and UO_2376 (O_2376,N_19928,N_19834);
or UO_2377 (O_2377,N_19986,N_19813);
xor UO_2378 (O_2378,N_19888,N_19953);
and UO_2379 (O_2379,N_19881,N_19954);
xor UO_2380 (O_2380,N_19834,N_19818);
and UO_2381 (O_2381,N_19986,N_19871);
or UO_2382 (O_2382,N_19804,N_19944);
xor UO_2383 (O_2383,N_19921,N_19861);
nand UO_2384 (O_2384,N_19841,N_19838);
xor UO_2385 (O_2385,N_19882,N_19943);
or UO_2386 (O_2386,N_19997,N_19852);
or UO_2387 (O_2387,N_19812,N_19926);
nor UO_2388 (O_2388,N_19914,N_19974);
nand UO_2389 (O_2389,N_19982,N_19994);
nand UO_2390 (O_2390,N_19948,N_19972);
nand UO_2391 (O_2391,N_19848,N_19938);
and UO_2392 (O_2392,N_19815,N_19892);
or UO_2393 (O_2393,N_19908,N_19800);
and UO_2394 (O_2394,N_19974,N_19916);
or UO_2395 (O_2395,N_19820,N_19916);
or UO_2396 (O_2396,N_19806,N_19951);
nand UO_2397 (O_2397,N_19862,N_19969);
and UO_2398 (O_2398,N_19903,N_19842);
or UO_2399 (O_2399,N_19855,N_19950);
and UO_2400 (O_2400,N_19807,N_19800);
or UO_2401 (O_2401,N_19947,N_19816);
xor UO_2402 (O_2402,N_19871,N_19833);
nor UO_2403 (O_2403,N_19949,N_19989);
nor UO_2404 (O_2404,N_19800,N_19812);
and UO_2405 (O_2405,N_19919,N_19882);
nand UO_2406 (O_2406,N_19933,N_19841);
and UO_2407 (O_2407,N_19842,N_19997);
nor UO_2408 (O_2408,N_19802,N_19811);
and UO_2409 (O_2409,N_19863,N_19815);
nand UO_2410 (O_2410,N_19957,N_19959);
nor UO_2411 (O_2411,N_19841,N_19861);
nor UO_2412 (O_2412,N_19933,N_19923);
nand UO_2413 (O_2413,N_19931,N_19806);
and UO_2414 (O_2414,N_19910,N_19845);
xor UO_2415 (O_2415,N_19931,N_19941);
xor UO_2416 (O_2416,N_19829,N_19942);
nor UO_2417 (O_2417,N_19954,N_19833);
or UO_2418 (O_2418,N_19868,N_19845);
xor UO_2419 (O_2419,N_19829,N_19881);
xnor UO_2420 (O_2420,N_19855,N_19831);
or UO_2421 (O_2421,N_19846,N_19863);
and UO_2422 (O_2422,N_19922,N_19897);
or UO_2423 (O_2423,N_19926,N_19962);
nor UO_2424 (O_2424,N_19884,N_19858);
and UO_2425 (O_2425,N_19885,N_19896);
nand UO_2426 (O_2426,N_19812,N_19805);
or UO_2427 (O_2427,N_19994,N_19925);
or UO_2428 (O_2428,N_19819,N_19890);
xor UO_2429 (O_2429,N_19887,N_19993);
nand UO_2430 (O_2430,N_19921,N_19858);
and UO_2431 (O_2431,N_19837,N_19954);
nand UO_2432 (O_2432,N_19997,N_19834);
and UO_2433 (O_2433,N_19993,N_19996);
or UO_2434 (O_2434,N_19910,N_19837);
or UO_2435 (O_2435,N_19932,N_19934);
or UO_2436 (O_2436,N_19800,N_19877);
nand UO_2437 (O_2437,N_19937,N_19804);
nand UO_2438 (O_2438,N_19906,N_19807);
nor UO_2439 (O_2439,N_19838,N_19846);
or UO_2440 (O_2440,N_19910,N_19858);
nand UO_2441 (O_2441,N_19804,N_19886);
nand UO_2442 (O_2442,N_19906,N_19801);
xnor UO_2443 (O_2443,N_19840,N_19883);
xnor UO_2444 (O_2444,N_19987,N_19825);
or UO_2445 (O_2445,N_19921,N_19870);
and UO_2446 (O_2446,N_19816,N_19957);
or UO_2447 (O_2447,N_19813,N_19857);
nand UO_2448 (O_2448,N_19845,N_19875);
xnor UO_2449 (O_2449,N_19976,N_19810);
or UO_2450 (O_2450,N_19854,N_19930);
nor UO_2451 (O_2451,N_19821,N_19982);
nor UO_2452 (O_2452,N_19994,N_19822);
xnor UO_2453 (O_2453,N_19838,N_19836);
nor UO_2454 (O_2454,N_19880,N_19912);
nand UO_2455 (O_2455,N_19823,N_19902);
or UO_2456 (O_2456,N_19911,N_19897);
xor UO_2457 (O_2457,N_19977,N_19853);
nand UO_2458 (O_2458,N_19973,N_19987);
or UO_2459 (O_2459,N_19889,N_19873);
and UO_2460 (O_2460,N_19806,N_19908);
xor UO_2461 (O_2461,N_19829,N_19844);
xnor UO_2462 (O_2462,N_19970,N_19813);
or UO_2463 (O_2463,N_19953,N_19998);
nor UO_2464 (O_2464,N_19979,N_19805);
nor UO_2465 (O_2465,N_19827,N_19992);
xnor UO_2466 (O_2466,N_19978,N_19976);
nand UO_2467 (O_2467,N_19942,N_19990);
and UO_2468 (O_2468,N_19962,N_19879);
nand UO_2469 (O_2469,N_19801,N_19920);
nand UO_2470 (O_2470,N_19820,N_19976);
or UO_2471 (O_2471,N_19811,N_19935);
or UO_2472 (O_2472,N_19999,N_19963);
nand UO_2473 (O_2473,N_19933,N_19976);
and UO_2474 (O_2474,N_19956,N_19857);
nor UO_2475 (O_2475,N_19911,N_19960);
nand UO_2476 (O_2476,N_19951,N_19852);
or UO_2477 (O_2477,N_19804,N_19935);
nand UO_2478 (O_2478,N_19962,N_19967);
or UO_2479 (O_2479,N_19998,N_19899);
nand UO_2480 (O_2480,N_19896,N_19949);
nor UO_2481 (O_2481,N_19820,N_19908);
nand UO_2482 (O_2482,N_19996,N_19872);
and UO_2483 (O_2483,N_19918,N_19997);
nor UO_2484 (O_2484,N_19806,N_19928);
and UO_2485 (O_2485,N_19991,N_19836);
nand UO_2486 (O_2486,N_19909,N_19870);
and UO_2487 (O_2487,N_19920,N_19901);
or UO_2488 (O_2488,N_19874,N_19835);
nor UO_2489 (O_2489,N_19981,N_19888);
and UO_2490 (O_2490,N_19935,N_19913);
and UO_2491 (O_2491,N_19856,N_19942);
and UO_2492 (O_2492,N_19934,N_19858);
and UO_2493 (O_2493,N_19802,N_19991);
xnor UO_2494 (O_2494,N_19825,N_19992);
nand UO_2495 (O_2495,N_19823,N_19878);
or UO_2496 (O_2496,N_19904,N_19878);
or UO_2497 (O_2497,N_19965,N_19926);
nor UO_2498 (O_2498,N_19863,N_19878);
nand UO_2499 (O_2499,N_19866,N_19810);
endmodule