module basic_3000_30000_3500_150_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
and U0 (N_0,In_205,In_2992);
nand U1 (N_1,In_192,In_2485);
or U2 (N_2,In_888,In_2802);
nor U3 (N_3,In_991,In_2411);
nor U4 (N_4,In_1497,In_943);
xor U5 (N_5,In_2666,In_1196);
xor U6 (N_6,In_180,In_2255);
xnor U7 (N_7,In_2360,In_237);
xnor U8 (N_8,In_1019,In_2664);
xor U9 (N_9,In_1121,In_2810);
xor U10 (N_10,In_770,In_2791);
nor U11 (N_11,In_2168,In_2310);
or U12 (N_12,In_158,In_2646);
xnor U13 (N_13,In_465,In_663);
nor U14 (N_14,In_1869,In_141);
nand U15 (N_15,In_1775,In_329);
or U16 (N_16,In_594,In_681);
nor U17 (N_17,In_1906,In_1919);
xor U18 (N_18,In_394,In_1052);
and U19 (N_19,In_1447,In_214);
and U20 (N_20,In_2916,In_1727);
or U21 (N_21,In_246,In_643);
nor U22 (N_22,In_1818,In_2221);
nor U23 (N_23,In_1256,In_79);
and U24 (N_24,In_2288,In_2275);
and U25 (N_25,In_1507,In_646);
nand U26 (N_26,In_1281,In_1228);
or U27 (N_27,In_2227,In_190);
or U28 (N_28,In_2548,In_426);
and U29 (N_29,In_880,In_2053);
xnor U30 (N_30,In_1086,In_1306);
nand U31 (N_31,In_1672,In_863);
nor U32 (N_32,In_587,In_2052);
xor U33 (N_33,In_1479,In_1174);
xor U34 (N_34,In_658,In_1324);
nor U35 (N_35,In_199,In_605);
nor U36 (N_36,In_1848,In_2070);
and U37 (N_37,In_771,In_2497);
xnor U38 (N_38,In_659,In_2378);
and U39 (N_39,In_371,In_172);
or U40 (N_40,In_1406,In_2060);
and U41 (N_41,In_1565,In_1269);
or U42 (N_42,In_2491,In_2072);
nand U43 (N_43,In_2804,In_2469);
and U44 (N_44,In_19,In_1071);
and U45 (N_45,In_2960,In_431);
or U46 (N_46,In_2343,In_2772);
xnor U47 (N_47,In_1193,In_1960);
and U48 (N_48,In_1018,In_1874);
nand U49 (N_49,In_1203,In_2092);
nand U50 (N_50,In_151,In_1561);
nor U51 (N_51,In_1474,In_621);
or U52 (N_52,In_1751,In_2235);
or U53 (N_53,In_1393,In_2761);
nand U54 (N_54,In_1369,In_1850);
or U55 (N_55,In_344,In_1084);
nand U56 (N_56,In_1961,In_2321);
or U57 (N_57,In_869,In_853);
and U58 (N_58,In_2678,In_2393);
or U59 (N_59,In_1682,In_357);
xnor U60 (N_60,In_5,In_1711);
nand U61 (N_61,In_2619,In_2532);
xor U62 (N_62,In_1648,In_130);
nand U63 (N_63,In_2935,In_2312);
and U64 (N_64,In_2910,In_731);
and U65 (N_65,In_43,In_1326);
nor U66 (N_66,In_2345,In_2823);
nand U67 (N_67,In_2254,In_2387);
nand U68 (N_68,In_2408,In_2170);
or U69 (N_69,In_1245,In_241);
and U70 (N_70,In_2568,In_1097);
nand U71 (N_71,In_704,In_1255);
or U72 (N_72,In_528,In_2549);
nor U73 (N_73,In_496,In_2199);
xor U74 (N_74,In_562,In_359);
or U75 (N_75,In_2702,In_70);
and U76 (N_76,In_1892,In_2332);
nand U77 (N_77,In_2692,In_2529);
nor U78 (N_78,In_2507,In_2969);
nor U79 (N_79,In_97,In_657);
nand U80 (N_80,In_1580,In_1272);
nand U81 (N_81,In_1233,In_2596);
xor U82 (N_82,In_234,In_2657);
and U83 (N_83,In_1237,In_1585);
or U84 (N_84,In_1146,In_764);
nor U85 (N_85,In_2103,In_1885);
xnor U86 (N_86,In_1043,In_2371);
or U87 (N_87,In_872,In_381);
xnor U88 (N_88,In_1724,In_1540);
nand U89 (N_89,In_1800,In_150);
nand U90 (N_90,In_538,In_1622);
or U91 (N_91,In_1236,In_2020);
and U92 (N_92,In_873,In_446);
xor U93 (N_93,In_610,In_1931);
xor U94 (N_94,In_1488,In_2899);
nand U95 (N_95,In_2137,In_352);
nand U96 (N_96,In_1697,In_2127);
and U97 (N_97,In_466,In_1487);
or U98 (N_98,In_1504,In_469);
nand U99 (N_99,In_418,In_2089);
nand U100 (N_100,In_1472,In_1963);
and U101 (N_101,In_2731,In_523);
xnor U102 (N_102,In_1460,In_48);
xor U103 (N_103,In_2465,In_2264);
nor U104 (N_104,In_1061,In_1400);
nor U105 (N_105,In_2400,In_2155);
nand U106 (N_106,In_2233,In_2659);
nand U107 (N_107,In_1415,In_890);
or U108 (N_108,In_2977,In_2021);
or U109 (N_109,In_2237,In_1403);
and U110 (N_110,In_1574,In_938);
nor U111 (N_111,In_1897,In_1559);
and U112 (N_112,In_1187,In_1912);
and U113 (N_113,In_987,In_1270);
nor U114 (N_114,In_1787,In_2669);
or U115 (N_115,In_277,In_833);
nand U116 (N_116,In_174,In_1277);
nand U117 (N_117,In_617,In_2708);
nand U118 (N_118,In_1597,In_198);
nand U119 (N_119,In_2816,In_498);
or U120 (N_120,In_837,In_1240);
xnor U121 (N_121,In_1340,In_2487);
and U122 (N_122,In_2427,In_1160);
or U123 (N_123,In_2163,In_2908);
nor U124 (N_124,In_2434,In_564);
xor U125 (N_125,In_328,In_456);
or U126 (N_126,In_188,In_239);
xor U127 (N_127,In_817,In_2043);
nand U128 (N_128,In_815,In_2689);
nand U129 (N_129,In_2138,In_149);
or U130 (N_130,In_2156,In_143);
or U131 (N_131,In_1327,In_145);
nor U132 (N_132,In_103,In_399);
xnor U133 (N_133,In_666,In_1982);
nor U134 (N_134,In_1986,In_631);
and U135 (N_135,In_1420,In_1035);
nor U136 (N_136,In_2388,In_2962);
nor U137 (N_137,In_2871,In_950);
xnor U138 (N_138,In_2697,In_979);
and U139 (N_139,In_1038,In_374);
nor U140 (N_140,In_1396,In_2311);
xor U141 (N_141,In_2826,In_2431);
and U142 (N_142,In_2190,In_1341);
and U143 (N_143,In_376,In_1127);
and U144 (N_144,In_2281,In_1323);
and U145 (N_145,In_2304,In_812);
nor U146 (N_146,In_1490,In_292);
nand U147 (N_147,In_2048,In_2894);
and U148 (N_148,In_2918,In_1463);
or U149 (N_149,In_1795,In_509);
xor U150 (N_150,In_1915,In_1829);
or U151 (N_151,In_1894,In_1675);
and U152 (N_152,In_1158,In_2209);
nor U153 (N_153,In_2954,In_1070);
nand U154 (N_154,In_40,In_1657);
nand U155 (N_155,In_64,In_2001);
or U156 (N_156,In_1527,In_651);
or U157 (N_157,In_2970,In_2982);
nor U158 (N_158,In_1455,In_692);
or U159 (N_159,In_721,In_2153);
and U160 (N_160,In_1016,In_1512);
and U161 (N_161,In_2890,In_1405);
nor U162 (N_162,In_2699,In_449);
nor U163 (N_163,In_2464,In_316);
and U164 (N_164,In_2779,In_2618);
nor U165 (N_165,In_1433,In_2205);
xnor U166 (N_166,In_744,In_856);
or U167 (N_167,In_1826,In_897);
xor U168 (N_168,In_2,In_436);
or U169 (N_169,In_1048,In_209);
or U170 (N_170,In_536,In_1688);
nor U171 (N_171,In_1589,In_1284);
nand U172 (N_172,In_1558,In_1769);
and U173 (N_173,In_1099,In_1810);
nor U174 (N_174,In_1092,In_1744);
nor U175 (N_175,In_726,In_53);
nor U176 (N_176,In_361,In_848);
nand U177 (N_177,In_1654,In_1047);
and U178 (N_178,In_2905,In_1737);
or U179 (N_179,In_261,In_541);
xnor U180 (N_180,In_1950,In_322);
nand U181 (N_181,In_1571,In_849);
and U182 (N_182,In_1861,In_690);
xor U183 (N_183,In_1582,In_122);
nand U184 (N_184,In_2746,In_558);
nand U185 (N_185,In_1592,In_2315);
or U186 (N_186,In_1481,In_2513);
xnor U187 (N_187,In_1884,In_1870);
or U188 (N_188,In_2650,In_2914);
nor U189 (N_189,In_2883,In_2284);
and U190 (N_190,In_257,In_989);
nor U191 (N_191,In_1660,In_1204);
and U192 (N_192,In_506,In_1350);
nor U193 (N_193,In_1685,In_2068);
or U194 (N_194,In_1937,In_2055);
nor U195 (N_195,In_1087,In_1090);
or U196 (N_196,In_2616,In_1318);
or U197 (N_197,In_655,In_1927);
nand U198 (N_198,In_423,In_1473);
and U199 (N_199,In_2269,In_1839);
nand U200 (N_200,In_458,In_1069);
and U201 (N_201,In_1772,N_89);
nor U202 (N_202,In_2476,In_569);
nor U203 (N_203,In_638,In_1480);
xnor U204 (N_204,N_53,In_2161);
xor U205 (N_205,In_696,In_1109);
and U206 (N_206,In_922,In_823);
xnor U207 (N_207,In_232,In_1469);
or U208 (N_208,In_1786,N_130);
or U209 (N_209,In_2189,In_2850);
nor U210 (N_210,In_262,In_228);
and U211 (N_211,In_264,In_1254);
nand U212 (N_212,In_337,In_1542);
nor U213 (N_213,In_566,In_1432);
or U214 (N_214,In_2733,In_8);
xor U215 (N_215,In_1185,In_2014);
nand U216 (N_216,In_1820,In_334);
and U217 (N_217,In_902,In_2830);
nor U218 (N_218,N_43,In_2869);
nor U219 (N_219,In_1312,In_1696);
nor U220 (N_220,In_580,In_850);
nor U221 (N_221,In_1649,In_1266);
xnor U222 (N_222,In_1450,In_2739);
nand U223 (N_223,In_1532,In_414);
nor U224 (N_224,In_2024,In_2492);
or U225 (N_225,In_2817,In_1719);
nand U226 (N_226,In_2394,In_2088);
or U227 (N_227,In_2564,N_135);
xnor U228 (N_228,In_2653,In_1032);
nor U229 (N_229,In_947,In_1921);
nor U230 (N_230,In_2012,In_2122);
nand U231 (N_231,In_2645,In_369);
nand U232 (N_232,In_1599,In_1855);
xor U233 (N_233,In_37,In_1259);
and U234 (N_234,In_219,In_1928);
nand U235 (N_235,N_83,In_2167);
nand U236 (N_236,In_2061,In_2824);
xnor U237 (N_237,N_105,N_154);
or U238 (N_238,In_2546,In_1638);
and U239 (N_239,In_2740,In_2098);
nand U240 (N_240,In_94,In_1107);
and U241 (N_241,In_1389,In_975);
and U242 (N_242,In_518,In_2035);
and U243 (N_243,In_2204,In_2778);
xnor U244 (N_244,In_516,In_137);
xnor U245 (N_245,In_1524,In_1890);
or U246 (N_246,In_2114,In_2803);
and U247 (N_247,In_1129,N_142);
nand U248 (N_248,In_1082,In_2839);
nand U249 (N_249,In_2142,In_495);
nand U250 (N_250,In_2323,In_18);
or U251 (N_251,In_2065,In_1947);
and U252 (N_252,In_311,In_886);
or U253 (N_253,In_2860,In_912);
nand U254 (N_254,In_248,In_27);
and U255 (N_255,In_2352,In_388);
nand U256 (N_256,In_2196,In_2051);
nand U257 (N_257,N_75,In_274);
nand U258 (N_258,In_308,N_4);
and U259 (N_259,In_2732,In_949);
and U260 (N_260,In_2843,In_1801);
nor U261 (N_261,In_2931,In_1922);
nor U262 (N_262,In_1679,In_1546);
nor U263 (N_263,In_2078,In_1948);
nand U264 (N_264,In_756,In_1550);
xor U265 (N_265,In_884,In_1208);
nand U266 (N_266,In_1872,In_1741);
or U267 (N_267,In_755,In_772);
nor U268 (N_268,In_1011,In_1918);
and U269 (N_269,In_951,In_283);
nand U270 (N_270,In_2223,In_624);
nand U271 (N_271,In_2978,In_2928);
nand U272 (N_272,In_2643,In_404);
xnor U273 (N_273,In_2895,N_178);
xor U274 (N_274,In_2289,In_2423);
nand U275 (N_275,In_1513,In_427);
nor U276 (N_276,In_207,In_2220);
nand U277 (N_277,In_2555,N_31);
and U278 (N_278,In_2923,In_99);
nor U279 (N_279,In_769,In_2414);
nor U280 (N_280,In_1669,In_2228);
nor U281 (N_281,In_708,In_2855);
nor U282 (N_282,In_1276,In_2131);
nor U283 (N_283,In_1118,In_1262);
xnor U284 (N_284,In_2822,In_342);
nand U285 (N_285,In_1799,In_16);
nor U286 (N_286,N_169,In_602);
nand U287 (N_287,In_2663,In_223);
xor U288 (N_288,In_1845,In_284);
or U289 (N_289,In_1505,In_2744);
nand U290 (N_290,In_1548,In_2759);
xnor U291 (N_291,In_1837,In_1362);
nor U292 (N_292,In_1722,In_782);
nand U293 (N_293,In_967,In_1162);
or U294 (N_294,In_2239,N_137);
or U295 (N_295,In_953,In_1503);
nand U296 (N_296,In_2166,In_941);
xor U297 (N_297,In_1287,In_2903);
xor U298 (N_298,In_410,In_2107);
or U299 (N_299,In_472,In_2187);
xor U300 (N_300,In_2374,N_58);
nor U301 (N_301,In_1085,In_2880);
xnor U302 (N_302,In_570,In_1111);
xor U303 (N_303,In_2533,In_164);
and U304 (N_304,In_306,In_1310);
and U305 (N_305,In_87,In_1014);
xor U306 (N_306,In_703,In_1625);
xor U307 (N_307,N_174,In_459);
nand U308 (N_308,In_350,In_1893);
xor U309 (N_309,In_1040,In_2994);
or U310 (N_310,In_182,In_727);
or U311 (N_311,N_85,In_12);
or U312 (N_312,In_1367,In_2133);
nor U313 (N_313,In_2652,In_1611);
nor U314 (N_314,In_2683,In_996);
or U315 (N_315,In_1384,In_400);
nor U316 (N_316,In_2921,In_1847);
nand U317 (N_317,In_607,In_1764);
nand U318 (N_318,In_358,In_196);
or U319 (N_319,In_2398,In_993);
xnor U320 (N_320,In_1655,In_642);
and U321 (N_321,In_2490,In_1910);
nand U322 (N_322,In_1316,In_1157);
or U323 (N_323,In_2842,In_2277);
xor U324 (N_324,In_2541,In_2242);
and U325 (N_325,In_1267,In_2225);
nand U326 (N_326,N_132,In_299);
xnor U327 (N_327,In_2436,In_1429);
nand U328 (N_328,In_356,In_2536);
xor U329 (N_329,In_2481,In_76);
nand U330 (N_330,In_1049,In_111);
nand U331 (N_331,In_2306,In_2213);
nand U332 (N_332,In_741,In_2044);
or U333 (N_333,In_448,In_2856);
or U334 (N_334,In_482,In_2134);
nand U335 (N_335,In_1138,In_2256);
nor U336 (N_336,In_2219,In_476);
nor U337 (N_337,In_224,In_1002);
nor U338 (N_338,In_1357,In_120);
nor U339 (N_339,In_416,In_2537);
and U340 (N_340,In_233,In_442);
xnor U341 (N_341,In_2795,In_181);
nand U342 (N_342,In_905,In_489);
nand U343 (N_343,In_2105,In_1286);
nand U344 (N_344,N_74,N_57);
nor U345 (N_345,N_160,In_827);
nand U346 (N_346,In_811,In_924);
or U347 (N_347,N_171,In_2317);
xnor U348 (N_348,In_2101,In_2151);
nand U349 (N_349,In_1135,In_927);
nand U350 (N_350,In_242,In_445);
xnor U351 (N_351,In_461,In_2948);
nor U352 (N_352,In_1687,In_2725);
or U353 (N_353,In_2140,In_2927);
or U354 (N_354,In_2756,In_2493);
xor U355 (N_355,In_2463,In_152);
nor U356 (N_356,In_47,In_1545);
and U357 (N_357,In_1934,In_1621);
or U358 (N_358,In_675,N_109);
and U359 (N_359,In_2297,In_255);
xnor U360 (N_360,In_1006,In_2113);
and U361 (N_361,In_2974,In_603);
xor U362 (N_362,In_2967,In_1533);
and U363 (N_363,In_1788,In_1511);
or U364 (N_364,In_2447,In_2329);
nand U365 (N_365,In_2334,In_718);
nand U366 (N_366,In_1975,N_50);
nor U367 (N_367,In_355,In_2303);
or U368 (N_368,In_2520,In_1924);
xnor U369 (N_369,In_2644,In_2571);
or U370 (N_370,In_1656,In_742);
xnor U371 (N_371,In_1944,In_629);
and U372 (N_372,In_453,In_543);
nand U373 (N_373,In_1761,In_29);
or U374 (N_374,In_170,N_12);
and U375 (N_375,N_80,In_2988);
nor U376 (N_376,In_2963,In_619);
and U377 (N_377,In_1750,In_1232);
or U378 (N_378,In_1202,In_2123);
and U379 (N_379,In_2715,In_834);
and U380 (N_380,In_1067,In_1541);
nand U381 (N_381,In_1017,In_1796);
or U382 (N_382,N_46,In_1205);
and U383 (N_383,In_49,In_26);
and U384 (N_384,In_66,In_857);
nand U385 (N_385,N_60,In_2724);
nand U386 (N_386,In_438,In_450);
nand U387 (N_387,In_2353,In_2483);
and U388 (N_388,N_124,N_44);
xnor U389 (N_389,In_1123,In_1417);
and U390 (N_390,In_1154,In_2718);
xnor U391 (N_391,In_1275,In_2557);
or U392 (N_392,In_434,N_64);
xor U393 (N_393,In_2039,In_377);
and U394 (N_394,In_1115,In_1189);
nand U395 (N_395,In_980,In_866);
nor U396 (N_396,In_317,In_2471);
and U397 (N_397,In_1021,In_1965);
nor U398 (N_398,In_678,In_432);
or U399 (N_399,In_1206,In_2747);
and U400 (N_400,N_294,In_1386);
xor U401 (N_401,N_383,In_2207);
xnor U402 (N_402,In_1673,In_1586);
nor U403 (N_403,In_2745,In_2835);
nand U404 (N_404,In_707,In_669);
xnor U405 (N_405,In_2419,N_213);
and U406 (N_406,In_1242,In_2703);
or U407 (N_407,In_2631,In_294);
xnor U408 (N_408,In_2682,In_1435);
and U409 (N_409,In_36,In_1449);
nor U410 (N_410,In_2130,In_61);
or U411 (N_411,In_1112,In_325);
nand U412 (N_412,In_2143,In_945);
xnor U413 (N_413,In_1445,In_830);
xor U414 (N_414,In_2511,In_2265);
xnor U415 (N_415,In_1785,In_184);
xnor U416 (N_416,In_1819,In_1853);
or U417 (N_417,In_958,In_1025);
and U418 (N_418,In_1590,N_317);
and U419 (N_419,N_251,In_499);
nor U420 (N_420,In_1780,In_333);
and U421 (N_421,In_917,In_2152);
nor U422 (N_422,N_6,N_81);
nor U423 (N_423,In_2047,N_259);
and U424 (N_424,In_2628,In_168);
nand U425 (N_425,In_2449,N_293);
or U426 (N_426,N_241,In_2552);
xor U427 (N_427,In_112,N_236);
and U428 (N_428,In_1343,N_147);
nand U429 (N_429,In_2050,In_1430);
nor U430 (N_430,N_289,N_226);
or U431 (N_431,N_8,N_387);
or U432 (N_432,In_2980,In_1570);
nor U433 (N_433,In_2093,In_1066);
nand U434 (N_434,N_98,In_1078);
and U435 (N_435,N_398,In_1282);
nor U436 (N_436,In_2837,In_1062);
and U437 (N_437,In_1584,N_66);
or U438 (N_438,In_1954,In_2307);
nand U439 (N_439,In_403,In_1168);
or U440 (N_440,N_248,In_2293);
and U441 (N_441,N_108,N_276);
nor U442 (N_442,In_1846,In_90);
nor U443 (N_443,N_245,In_1939);
and U444 (N_444,In_719,In_2097);
nor U445 (N_445,N_35,In_1268);
nand U446 (N_446,In_252,In_503);
nor U447 (N_447,In_487,In_2981);
xor U448 (N_448,In_165,In_1483);
nand U449 (N_449,N_390,In_2911);
and U450 (N_450,In_2128,In_1502);
or U451 (N_451,N_188,In_2809);
or U452 (N_452,In_354,In_253);
nor U453 (N_453,In_1331,In_1662);
and U454 (N_454,In_128,In_2925);
or U455 (N_455,In_2836,In_829);
and U456 (N_456,In_1218,In_1891);
xnor U457 (N_457,In_665,In_123);
or U458 (N_458,In_1972,In_1989);
nand U459 (N_459,In_684,In_673);
and U460 (N_460,In_2399,In_963);
nor U461 (N_461,In_183,In_2587);
or U462 (N_462,N_393,In_2146);
nand U463 (N_463,In_1770,In_2893);
or U464 (N_464,N_201,In_117);
nor U465 (N_465,N_21,In_1875);
nand U466 (N_466,N_219,In_2096);
nand U467 (N_467,In_2726,In_1949);
and U468 (N_468,In_2762,In_353);
xnor U469 (N_469,In_1349,In_1383);
xor U470 (N_470,In_2503,N_113);
nor U471 (N_471,N_388,In_2523);
or U472 (N_472,In_940,In_1905);
and U473 (N_473,In_1783,In_822);
nand U474 (N_474,N_76,In_2441);
and U475 (N_475,N_318,In_2569);
nand U476 (N_476,In_2456,In_2391);
or U477 (N_477,In_2117,In_1163);
nand U478 (N_478,In_2593,In_383);
or U479 (N_479,In_2665,In_272);
or U480 (N_480,In_1103,In_173);
nor U481 (N_481,In_2287,In_1752);
nand U482 (N_482,In_2116,N_26);
xor U483 (N_483,In_1251,In_714);
and U484 (N_484,In_1791,In_746);
nand U485 (N_485,In_2016,In_615);
xnor U486 (N_486,In_1454,In_961);
xnor U487 (N_487,In_1210,In_1740);
nor U488 (N_488,In_1227,In_2578);
xor U489 (N_489,In_1178,In_722);
xnor U490 (N_490,In_1661,In_1832);
or U491 (N_491,In_421,N_90);
nand U492 (N_492,In_74,N_344);
nor U493 (N_493,In_1581,In_1694);
nand U494 (N_494,In_2775,In_1217);
and U495 (N_495,In_1626,In_2976);
xor U496 (N_496,In_2807,In_240);
xor U497 (N_497,In_923,In_625);
xor U498 (N_498,In_2252,In_2685);
and U499 (N_499,In_793,In_2506);
and U500 (N_500,In_1354,In_1302);
xor U501 (N_501,In_1703,In_1140);
and U502 (N_502,In_1765,In_415);
xor U503 (N_503,In_1091,In_2862);
or U504 (N_504,In_1075,In_2815);
nor U505 (N_505,In_2877,In_2208);
nand U506 (N_506,In_127,In_490);
and U507 (N_507,In_2728,In_1666);
xnor U508 (N_508,N_300,In_2714);
or U509 (N_509,In_100,In_1739);
nand U510 (N_510,In_2933,In_1992);
nand U511 (N_511,In_125,In_1346);
nor U512 (N_512,In_542,In_676);
or U513 (N_513,In_1055,In_2349);
and U514 (N_514,N_197,In_845);
and U515 (N_515,In_1184,In_1640);
or U516 (N_516,In_131,In_1865);
or U517 (N_517,In_368,In_1706);
and U518 (N_518,In_844,In_2308);
nor U519 (N_519,In_2185,N_378);
xnor U520 (N_520,In_1636,In_1036);
xnor U521 (N_521,N_55,In_2084);
and U522 (N_522,In_1738,In_781);
and U523 (N_523,In_60,In_2214);
nand U524 (N_524,N_273,In_375);
and U525 (N_525,In_832,In_904);
or U526 (N_526,In_2338,In_2291);
or U527 (N_527,In_2621,In_1246);
xnor U528 (N_528,In_1882,In_501);
xor U529 (N_529,In_2104,In_2385);
nor U530 (N_530,In_338,In_1946);
xor U531 (N_531,In_2147,In_1176);
xnor U532 (N_532,In_2690,In_2328);
nand U533 (N_533,In_2301,In_1977);
xor U534 (N_534,In_613,In_780);
and U535 (N_535,N_167,In_2961);
nor U536 (N_536,In_493,In_1619);
xor U537 (N_537,N_72,In_124);
nor U538 (N_538,In_2958,In_2290);
nor U539 (N_539,In_2783,In_1811);
nand U540 (N_540,N_330,In_1003);
nor U541 (N_541,In_2342,In_2482);
nand U542 (N_542,In_505,In_2386);
nand U543 (N_543,In_1593,In_988);
nor U544 (N_544,In_671,In_437);
or U545 (N_545,In_485,In_1000);
nor U546 (N_546,In_2845,N_112);
or U547 (N_547,In_507,N_222);
nor U548 (N_548,In_1495,In_2340);
nor U549 (N_549,In_2430,In_2995);
nand U550 (N_550,N_96,In_2821);
nor U551 (N_551,N_184,In_1577);
nor U552 (N_552,In_1807,In_1475);
and U553 (N_553,In_2135,In_1864);
nand U554 (N_554,In_601,In_2554);
xnor U555 (N_555,In_1419,N_281);
or U556 (N_556,In_1743,In_2331);
and U557 (N_557,In_2531,In_1414);
xor U558 (N_558,In_310,In_579);
or U559 (N_559,In_1757,In_1710);
xnor U560 (N_560,In_2466,In_1311);
nand U561 (N_561,N_68,In_537);
or U562 (N_562,In_1222,N_380);
nand U563 (N_563,In_38,In_2852);
and U564 (N_564,In_2499,In_674);
or U565 (N_565,In_2647,In_2322);
nand U566 (N_566,In_492,In_2853);
nor U567 (N_567,In_2276,In_2542);
or U568 (N_568,In_2267,In_502);
nand U569 (N_569,In_725,In_439);
xnor U570 (N_570,In_1817,In_583);
or U571 (N_571,In_2629,In_2550);
nand U572 (N_572,In_1113,In_592);
xor U573 (N_573,In_2013,In_1155);
or U574 (N_574,In_1792,In_1351);
nor U575 (N_575,In_384,In_2884);
nor U576 (N_576,In_2486,In_1149);
nand U577 (N_577,In_1332,In_2222);
nor U578 (N_578,In_1423,In_2741);
xnor U579 (N_579,In_876,In_2410);
xnor U580 (N_580,In_1628,In_2661);
and U581 (N_581,In_799,In_195);
xor U582 (N_582,In_1911,In_1364);
or U583 (N_583,In_390,In_309);
nor U584 (N_584,In_2118,In_2944);
or U585 (N_585,In_743,In_2194);
nor U586 (N_586,In_1776,In_1427);
nand U587 (N_587,In_101,N_231);
and U588 (N_588,In_712,In_1781);
nand U589 (N_589,In_555,In_2253);
nand U590 (N_590,In_451,In_1691);
or U591 (N_591,In_556,In_1179);
nor U592 (N_592,In_1314,N_296);
xor U593 (N_593,N_302,In_441);
nor U594 (N_594,In_2169,In_2900);
and U595 (N_595,In_1841,In_295);
xnor U596 (N_596,In_1418,In_959);
or U597 (N_597,N_223,In_21);
nor U598 (N_598,N_33,In_296);
nand U599 (N_599,In_2319,In_1809);
xor U600 (N_600,N_298,In_2341);
xor U601 (N_601,In_870,N_290);
xor U602 (N_602,N_180,In_1623);
nand U603 (N_603,In_389,In_852);
nor U604 (N_604,In_1150,In_565);
nor U605 (N_605,In_2811,In_560);
nor U606 (N_606,In_2162,In_1665);
nor U607 (N_607,N_478,In_2259);
nor U608 (N_608,In_1583,N_490);
nor U609 (N_609,In_662,In_1436);
or U610 (N_610,In_153,In_1642);
nor U611 (N_611,N_368,In_80);
or U612 (N_612,In_1380,In_2673);
xor U613 (N_613,In_1526,In_710);
nor U614 (N_614,N_177,In_69);
or U615 (N_615,In_1098,N_111);
and U616 (N_616,In_4,In_794);
or U617 (N_617,In_545,In_1096);
xnor U618 (N_618,In_1936,In_760);
xor U619 (N_619,In_1220,N_527);
nor U620 (N_620,In_307,In_1325);
or U621 (N_621,N_110,In_1453);
nand U622 (N_622,In_2608,N_551);
nand U623 (N_623,In_1195,N_377);
nand U624 (N_624,In_977,In_1684);
and U625 (N_625,N_165,In_530);
and U626 (N_626,In_1725,N_181);
xnor U627 (N_627,In_2723,In_1244);
or U628 (N_628,In_2054,In_831);
and U629 (N_629,In_1736,In_738);
nor U630 (N_630,In_1401,In_2909);
xor U631 (N_631,In_2413,In_2675);
nand U632 (N_632,In_1605,In_2882);
and U633 (N_633,In_2734,N_539);
or U634 (N_634,In_634,In_96);
xnor U635 (N_635,In_1289,In_1437);
xor U636 (N_636,N_595,N_484);
xnor U637 (N_637,In_2330,N_13);
nand U638 (N_638,In_406,In_1057);
or U639 (N_639,In_654,N_559);
xnor U640 (N_640,N_435,In_649);
and U641 (N_641,In_1955,N_23);
and U642 (N_642,In_2261,In_2108);
or U643 (N_643,In_1122,In_2782);
and U644 (N_644,In_2881,In_1054);
nand U645 (N_645,N_136,In_1440);
nand U646 (N_646,N_565,N_345);
xor U647 (N_647,N_593,In_2100);
and U648 (N_648,In_121,In_1298);
and U649 (N_649,In_1482,N_534);
nand U650 (N_650,In_1397,In_2316);
or U651 (N_651,N_292,In_324);
and U652 (N_652,In_970,In_42);
or U653 (N_653,In_340,In_1767);
xor U654 (N_654,In_2710,In_1439);
or U655 (N_655,In_2292,In_2272);
nand U656 (N_656,N_91,In_1699);
and U657 (N_657,In_1632,In_2069);
and U658 (N_658,In_1899,In_2580);
and U659 (N_659,N_185,N_410);
xor U660 (N_660,In_1613,N_30);
and U661 (N_661,In_2864,In_1603);
and U662 (N_662,In_1288,In_2038);
xnor U663 (N_663,In_1042,In_1079);
and U664 (N_664,In_2736,In_636);
or U665 (N_665,In_1307,N_205);
xnor U666 (N_666,N_2,In_862);
nor U667 (N_667,N_562,In_2891);
and U668 (N_668,In_2245,In_1973);
xor U669 (N_669,In_2937,In_1979);
or U670 (N_670,In_939,In_1615);
xnor U671 (N_671,In_2594,In_2757);
nor U672 (N_672,In_1330,In_1372);
nor U673 (N_673,In_2444,In_997);
nor U674 (N_674,In_1895,N_326);
nand U675 (N_675,In_2501,In_2416);
nand U676 (N_676,N_24,In_2848);
nand U677 (N_677,In_1537,N_238);
or U678 (N_678,In_1838,In_2355);
or U679 (N_679,N_253,In_1538);
xnor U680 (N_680,In_1539,In_473);
nor U681 (N_681,N_578,In_6);
nand U682 (N_682,In_2144,In_1514);
and U683 (N_683,In_1072,In_2354);
nor U684 (N_684,In_139,In_2597);
and U685 (N_685,In_2073,In_1285);
xor U686 (N_686,N_99,In_2525);
nand U687 (N_687,In_1468,In_1012);
nor U688 (N_688,In_2781,In_650);
and U689 (N_689,N_40,In_142);
xnor U690 (N_690,N_414,In_1768);
nor U691 (N_691,In_648,In_2365);
and U692 (N_692,In_1608,In_312);
and U693 (N_693,In_1260,In_529);
or U694 (N_694,In_2879,N_524);
nand U695 (N_695,In_1650,In_2787);
xor U696 (N_696,N_584,In_900);
nand U697 (N_697,In_1523,In_1089);
nor U698 (N_698,N_427,In_935);
xor U699 (N_699,N_379,N_339);
nor U700 (N_700,In_728,In_2799);
nor U701 (N_701,In_1144,In_1366);
and U702 (N_702,In_305,N_324);
or U703 (N_703,In_2359,In_1602);
nor U704 (N_704,In_2515,In_1471);
nor U705 (N_705,In_2868,In_2602);
or U706 (N_706,In_300,In_1001);
xor U707 (N_707,In_2579,In_211);
nand U708 (N_708,In_2679,In_1145);
nand U709 (N_709,In_478,In_179);
or U710 (N_710,In_1104,In_568);
or U711 (N_711,N_592,In_1224);
xnor U712 (N_712,In_1843,N_331);
or U713 (N_713,N_284,In_600);
xnor U714 (N_714,In_2717,In_2585);
nor U715 (N_715,In_2825,In_753);
or U716 (N_716,In_82,In_1171);
xnor U717 (N_717,In_2812,N_469);
nand U718 (N_718,In_1379,In_2514);
nand U719 (N_719,In_35,In_942);
and U720 (N_720,N_221,N_510);
and U721 (N_721,N_515,In_954);
and U722 (N_722,N_202,In_798);
xor U723 (N_723,In_639,In_2929);
nor U724 (N_724,In_628,In_1368);
or U725 (N_725,N_364,In_1797);
nand U726 (N_726,N_509,In_894);
nand U727 (N_727,In_1653,In_2907);
or U728 (N_728,In_1422,In_1568);
nand U729 (N_729,In_366,In_2033);
or U730 (N_730,In_1974,In_1443);
and U731 (N_731,N_84,In_1130);
nand U732 (N_732,In_887,N_283);
nand U733 (N_733,In_835,N_338);
nor U734 (N_734,In_1375,N_311);
nand U735 (N_735,In_2164,In_1394);
or U736 (N_736,N_369,In_1390);
nand U737 (N_737,In_889,In_775);
or U738 (N_738,In_1529,In_641);
xnor U739 (N_739,In_2160,In_803);
nor U740 (N_740,In_2898,In_1177);
and U741 (N_741,N_573,In_1470);
or U742 (N_742,N_417,In_2528);
xor U743 (N_743,In_1243,N_428);
nor U744 (N_744,In_2649,In_2369);
xnor U745 (N_745,In_470,In_1569);
or U746 (N_746,In_2119,In_321);
nand U747 (N_747,N_454,In_2247);
or U748 (N_748,N_352,In_2432);
nor U749 (N_749,In_2770,N_119);
or U750 (N_750,In_1296,N_419);
xor U751 (N_751,In_2612,In_2007);
xor U752 (N_752,In_2010,In_1943);
or U753 (N_753,In_2902,In_1695);
or U754 (N_754,N_247,In_788);
nand U755 (N_755,N_360,In_2986);
nand U756 (N_756,N_228,In_1466);
nor U757 (N_757,In_1486,In_2681);
and U758 (N_758,In_711,In_2889);
or U759 (N_759,In_2614,In_413);
xor U760 (N_760,In_106,N_246);
or U761 (N_761,N_25,In_1438);
or U762 (N_762,N_3,In_2833);
or U763 (N_763,N_586,N_122);
xnor U764 (N_764,N_82,In_1456);
nand U765 (N_765,In_185,N_497);
or U766 (N_766,In_1223,In_393);
xor U767 (N_767,N_94,In_222);
nand U768 (N_768,In_471,In_715);
or U769 (N_769,N_441,N_240);
nor U770 (N_770,In_138,N_9);
nor U771 (N_771,In_2171,In_2324);
nand U772 (N_772,In_2111,N_459);
nor U773 (N_773,In_41,In_2081);
nand U774 (N_774,In_893,In_1416);
nor U775 (N_775,In_2186,In_774);
or U776 (N_776,In_2372,In_2755);
nand U777 (N_777,In_1026,In_2640);
and U778 (N_778,In_259,N_395);
and U779 (N_779,In_1360,In_379);
or U780 (N_780,In_609,In_2278);
nand U781 (N_781,In_298,N_268);
or U782 (N_782,In_899,In_1141);
nor U783 (N_783,In_526,N_521);
xor U784 (N_784,In_2892,N_305);
or U785 (N_785,In_1659,In_1452);
nor U786 (N_786,N_512,In_2455);
xor U787 (N_787,In_2454,N_483);
or U788 (N_788,In_2934,In_786);
xor U789 (N_789,In_2638,In_1183);
and U790 (N_790,In_2197,N_408);
and U791 (N_791,In_460,In_1257);
nor U792 (N_792,In_851,In_946);
or U793 (N_793,In_2712,In_1644);
nor U794 (N_794,N_541,In_210);
xor U795 (N_795,N_431,In_1081);
or U796 (N_796,In_1771,In_1729);
xor U797 (N_797,N_152,In_51);
and U798 (N_798,In_2438,In_488);
or U799 (N_799,In_2922,In_1595);
nor U800 (N_800,In_454,In_2535);
or U801 (N_801,In_1983,N_366);
nand U802 (N_802,N_216,In_532);
xnor U803 (N_803,N_336,In_962);
and U804 (N_804,In_2721,In_2786);
or U805 (N_805,In_903,In_2581);
xnor U806 (N_806,N_372,N_570);
nor U807 (N_807,In_623,In_1013);
or U808 (N_808,In_2610,In_1631);
nor U809 (N_809,In_572,In_46);
and U810 (N_810,In_1723,N_218);
or U811 (N_811,In_1898,In_1134);
xnor U812 (N_812,N_703,In_2145);
nand U813 (N_813,In_1498,In_964);
nor U814 (N_814,N_321,In_1731);
or U815 (N_815,In_2015,In_2806);
nand U816 (N_816,In_1990,In_396);
and U817 (N_817,In_2192,N_745);
nor U818 (N_818,In_2403,N_162);
xnor U819 (N_819,In_2840,N_176);
and U820 (N_820,In_281,In_2538);
nor U821 (N_821,In_578,In_191);
nor U822 (N_822,In_2609,In_1693);
nand U823 (N_823,In_2178,In_582);
and U824 (N_824,In_2458,In_1945);
or U825 (N_825,In_2818,N_642);
xnor U826 (N_826,N_106,N_545);
nand U827 (N_827,In_1039,In_2313);
xnor U828 (N_828,In_346,In_2773);
xor U829 (N_829,In_2872,In_1248);
or U830 (N_830,In_2534,N_536);
nor U831 (N_831,N_335,In_475);
and U832 (N_832,N_151,In_1301);
xor U833 (N_833,In_243,N_161);
xnor U834 (N_834,N_635,In_573);
nand U835 (N_835,In_2518,N_59);
nor U836 (N_836,N_118,In_2271);
nand U837 (N_837,In_1303,In_2987);
nor U838 (N_838,In_1076,In_896);
or U839 (N_839,In_11,In_2442);
xor U840 (N_840,N_115,N_457);
nand U841 (N_841,In_2124,N_420);
nor U842 (N_842,N_288,In_1690);
nor U843 (N_843,In_1674,In_1261);
and U844 (N_844,In_2562,In_2379);
nand U845 (N_845,In_1434,In_126);
xnor U846 (N_846,In_883,In_679);
xnor U847 (N_847,N_341,In_23);
and U848 (N_848,In_982,N_173);
or U849 (N_849,In_2606,In_2184);
nand U850 (N_850,In_218,In_2827);
xnor U851 (N_851,N_793,In_2279);
nand U852 (N_852,In_1247,In_1278);
nand U853 (N_853,In_2658,In_1755);
and U854 (N_854,In_1620,In_2510);
and U855 (N_855,In_575,In_1198);
and U856 (N_856,In_1216,In_428);
nand U857 (N_857,In_1059,In_705);
nand U858 (N_858,In_276,In_59);
and U859 (N_859,In_1197,In_95);
xor U860 (N_860,In_1033,In_1824);
nor U861 (N_861,N_437,In_392);
or U862 (N_862,N_705,In_86);
xor U863 (N_863,In_552,In_2000);
nand U864 (N_864,N_511,N_448);
xor U865 (N_865,N_45,In_1297);
and U866 (N_866,N_694,In_217);
and U867 (N_867,In_206,N_444);
nor U868 (N_868,In_1517,In_349);
or U869 (N_869,N_28,In_2768);
xnor U870 (N_870,In_263,In_2023);
xnor U871 (N_871,In_2504,In_1860);
xor U872 (N_872,N_492,In_2985);
or U873 (N_873,In_1388,In_2350);
and U874 (N_874,In_802,N_7);
xnor U875 (N_875,In_467,In_1344);
xor U876 (N_876,In_2173,In_2368);
or U877 (N_877,In_1215,In_15);
and U878 (N_878,In_1428,In_1053);
and U879 (N_879,In_2796,In_1652);
and U880 (N_880,N_482,In_2095);
or U881 (N_881,In_2639,In_2849);
or U882 (N_882,N_456,In_1271);
nand U883 (N_883,In_167,In_1101);
nand U884 (N_884,In_2769,In_1572);
or U885 (N_885,N_287,N_714);
xor U886 (N_886,N_148,In_2654);
or U887 (N_887,In_1790,In_2695);
and U888 (N_888,In_193,In_653);
nand U889 (N_889,In_1143,N_797);
nor U890 (N_890,In_776,In_189);
nand U891 (N_891,In_314,In_397);
nand U892 (N_892,In_640,In_2502);
nor U893 (N_893,In_1063,In_1214);
nor U894 (N_894,N_279,In_1280);
xnor U895 (N_895,In_1212,N_107);
xor U896 (N_896,In_2588,N_309);
or U897 (N_897,In_56,In_2865);
or U898 (N_898,N_737,N_750);
nand U899 (N_899,N_86,N_190);
and U900 (N_900,In_1766,N_720);
and U901 (N_901,In_1816,In_279);
xnor U902 (N_902,In_405,N_525);
nand U903 (N_903,In_735,In_435);
xor U904 (N_904,In_2945,N_477);
xor U905 (N_905,In_1951,N_631);
nor U906 (N_906,In_1762,In_1213);
or U907 (N_907,N_409,In_2059);
or U908 (N_908,In_119,In_2605);
nand U909 (N_909,In_254,In_1426);
or U910 (N_910,In_1962,In_2011);
xor U911 (N_911,In_135,In_1987);
xor U912 (N_912,N_687,In_2136);
nor U913 (N_913,In_611,N_206);
nor U914 (N_914,In_2694,In_2320);
xnor U915 (N_915,In_2709,In_2409);
or U916 (N_916,In_1534,In_986);
nand U917 (N_917,N_229,In_737);
nand U918 (N_918,In_2286,In_1747);
nand U919 (N_919,In_2424,In_1980);
xor U920 (N_920,N_572,In_550);
xnor U921 (N_921,In_670,In_1929);
xor U922 (N_922,In_2716,In_226);
or U923 (N_923,N_333,In_1477);
or U924 (N_924,In_1718,In_1676);
nand U925 (N_925,In_1333,N_755);
nand U926 (N_926,In_2077,In_2595);
nor U927 (N_927,In_75,In_2380);
nor U928 (N_928,In_2129,In_2066);
or U929 (N_929,N_523,In_819);
or U930 (N_930,In_2688,N_485);
nor U931 (N_931,In_1034,In_2120);
nand U932 (N_932,N_170,In_468);
nand U933 (N_933,In_1120,N_591);
nand U934 (N_934,In_944,In_203);
or U935 (N_935,N_239,In_1252);
nand U936 (N_936,In_2576,In_2217);
nand U937 (N_937,N_653,In_2950);
nand U938 (N_938,In_2484,In_2866);
nand U939 (N_939,N_52,N_698);
and U940 (N_940,In_2561,In_39);
xnor U941 (N_941,In_479,In_1748);
nor U942 (N_942,In_2071,In_966);
xnor U943 (N_943,In_1573,In_2032);
or U944 (N_944,In_687,N_346);
nand U945 (N_945,In_508,In_71);
or U946 (N_946,In_2874,N_365);
xor U947 (N_947,In_1392,In_2392);
nor U948 (N_948,In_163,In_574);
nor U949 (N_949,N_645,In_2148);
and U950 (N_950,In_2049,In_2997);
or U951 (N_951,In_2959,In_2159);
nor U952 (N_952,In_1190,In_1683);
or U953 (N_953,In_1064,In_1805);
nand U954 (N_954,In_1391,In_2941);
nor U955 (N_955,In_1606,In_391);
nor U956 (N_956,In_140,In_1320);
nor U957 (N_957,In_2999,In_1553);
nand U958 (N_958,In_1956,In_1803);
nor U959 (N_959,In_1907,In_236);
nand U960 (N_960,N_358,In_1667);
xnor U961 (N_961,In_2819,In_2457);
or U962 (N_962,N_325,N_322);
nand U963 (N_963,N_465,N_489);
xnor U964 (N_964,In_2335,In_25);
nand U965 (N_965,N_633,In_664);
and U966 (N_966,In_477,In_881);
nor U967 (N_967,In_2034,In_2382);
nor U968 (N_968,N_638,In_1041);
nor U969 (N_969,In_859,In_1338);
or U970 (N_970,In_2648,N_712);
nand U971 (N_971,In_2083,In_1821);
and U972 (N_972,In_227,In_2526);
or U973 (N_973,In_250,N_531);
or U974 (N_974,In_736,N_618);
nor U975 (N_975,N_747,In_419);
xor U976 (N_976,In_2964,In_1578);
or U977 (N_977,In_1866,In_2704);
nand U978 (N_978,In_430,In_1170);
nand U979 (N_979,In_1735,In_2838);
nor U980 (N_980,In_1500,In_55);
xor U981 (N_981,In_2031,N_783);
nor U982 (N_982,In_2611,In_1159);
nand U983 (N_983,N_606,In_906);
nand U984 (N_984,In_2446,N_744);
nor U985 (N_985,In_230,In_2302);
xor U986 (N_986,N_233,In_2415);
or U987 (N_987,In_1131,N_274);
xnor U988 (N_988,In_107,In_412);
or U989 (N_989,N_587,In_2383);
xnor U990 (N_990,In_287,In_2373);
or U991 (N_991,In_2973,In_1065);
or U992 (N_992,In_2461,In_72);
nand U993 (N_993,In_115,N_319);
xor U994 (N_994,In_411,N_449);
or U995 (N_995,In_7,In_2210);
or U996 (N_996,In_1709,N_356);
nor U997 (N_997,N_316,In_1749);
and U998 (N_998,In_1856,In_2468);
or U999 (N_999,In_1153,In_1562);
nand U1000 (N_1000,In_1376,In_864);
nor U1001 (N_1001,In_200,In_455);
xor U1002 (N_1002,In_315,N_227);
nand U1003 (N_1003,In_765,N_569);
nand U1004 (N_1004,N_911,N_577);
and U1005 (N_1005,In_757,N_314);
or U1006 (N_1006,In_524,N_262);
or U1007 (N_1007,In_50,In_2943);
nor U1008 (N_1008,In_2296,N_450);
xnor U1009 (N_1009,In_2662,In_425);
or U1010 (N_1010,N_935,In_520);
xor U1011 (N_1011,In_2042,In_2417);
xnor U1012 (N_1012,In_1971,N_22);
and U1013 (N_1013,In_1201,In_57);
and U1014 (N_1014,In_1175,N_467);
nand U1015 (N_1015,N_386,In_2099);
or U1016 (N_1016,In_335,In_108);
nand U1017 (N_1017,In_2401,N_832);
or U1018 (N_1018,N_590,In_1172);
and U1019 (N_1019,In_2700,In_1802);
and U1020 (N_1020,In_178,N_664);
nor U1021 (N_1021,N_114,In_148);
and U1022 (N_1022,In_2767,In_622);
and U1023 (N_1023,N_726,In_956);
nand U1024 (N_1024,N_736,In_166);
or U1025 (N_1025,In_2676,In_2076);
and U1026 (N_1026,In_796,In_2157);
nand U1027 (N_1027,N_146,In_2358);
and U1028 (N_1028,In_2112,In_213);
and U1029 (N_1029,N_824,In_1630);
nand U1030 (N_1030,In_1361,In_2854);
and U1031 (N_1031,In_1139,In_2336);
or U1032 (N_1032,N_285,N_158);
xor U1033 (N_1033,In_2738,In_2750);
or U1034 (N_1034,N_941,In_1528);
nor U1035 (N_1035,In_2236,In_1756);
or U1036 (N_1036,In_2730,N_873);
or U1037 (N_1037,In_1782,In_1510);
xnor U1038 (N_1038,N_991,In_1300);
nor U1039 (N_1039,N_297,In_58);
and U1040 (N_1040,In_2574,N_632);
nor U1041 (N_1041,N_667,N_889);
xnor U1042 (N_1042,N_998,In_825);
or U1043 (N_1043,In_871,In_373);
nand U1044 (N_1044,In_596,In_1322);
and U1045 (N_1045,In_2957,N_780);
nand U1046 (N_1046,In_1840,In_1188);
nor U1047 (N_1047,N_626,N_451);
or U1048 (N_1048,In_1823,In_931);
xor U1049 (N_1049,In_1871,In_2777);
and U1050 (N_1050,In_875,In_362);
and U1051 (N_1051,In_2087,In_2851);
nor U1052 (N_1052,N_850,In_1813);
and U1053 (N_1053,N_254,In_2670);
nor U1054 (N_1054,N_79,N_355);
and U1055 (N_1055,In_2405,In_212);
nand U1056 (N_1056,N_910,In_504);
nand U1057 (N_1057,N_867,In_595);
nand U1058 (N_1058,N_649,N_447);
xor U1059 (N_1059,In_1457,In_2121);
xor U1060 (N_1060,In_688,N_840);
xor U1061 (N_1061,N_960,N_438);
xor U1062 (N_1062,In_301,In_1941);
nor U1063 (N_1063,In_1377,In_1421);
nor U1064 (N_1064,In_1506,In_895);
nor U1065 (N_1065,N_351,In_2180);
nor U1066 (N_1066,In_265,In_1745);
or U1067 (N_1067,N_243,In_2636);
and U1068 (N_1068,In_1116,In_668);
and U1069 (N_1069,N_502,In_593);
or U1070 (N_1070,N_674,In_13);
or U1071 (N_1071,In_2231,In_402);
nor U1072 (N_1072,N_877,In_2743);
nor U1073 (N_1073,In_1485,N_563);
nor U1074 (N_1074,N_430,N_400);
nor U1075 (N_1075,In_1913,In_2870);
nand U1076 (N_1076,N_814,In_549);
nor U1077 (N_1077,In_2058,N_820);
or U1078 (N_1078,N_462,In_2599);
and U1079 (N_1079,In_2539,In_2005);
and U1080 (N_1080,In_1253,In_2508);
xnor U1081 (N_1081,In_937,In_1981);
nor U1082 (N_1082,N_602,In_633);
xor U1083 (N_1083,In_2283,In_2930);
nor U1084 (N_1084,N_537,In_820);
or U1085 (N_1085,In_2126,N_903);
or U1086 (N_1086,In_2412,In_1348);
and U1087 (N_1087,In_1442,N_163);
and U1088 (N_1088,In_1953,N_735);
and U1089 (N_1089,In_1617,In_1588);
or U1090 (N_1090,In_2627,In_1173);
and U1091 (N_1091,In_515,In_395);
or U1092 (N_1092,N_717,In_2046);
nand U1093 (N_1093,In_1024,In_652);
or U1094 (N_1094,In_2624,In_285);
nand U1095 (N_1095,In_928,In_1412);
and U1096 (N_1096,In_1408,In_1876);
or U1097 (N_1097,In_2498,In_1137);
and U1098 (N_1098,N_842,In_2752);
nor U1099 (N_1099,N_871,In_2200);
nand U1100 (N_1100,In_855,N_678);
xnor U1101 (N_1101,In_1133,N_813);
and U1102 (N_1102,In_161,In_635);
xnor U1103 (N_1103,In_878,N_320);
nor U1104 (N_1104,In_531,In_867);
xor U1105 (N_1105,N_748,In_1575);
xnor U1106 (N_1106,N_203,In_1920);
nand U1107 (N_1107,N_925,In_1598);
nand U1108 (N_1108,In_2737,In_32);
nor U1109 (N_1109,In_2592,N_772);
nand U1110 (N_1110,In_63,N_19);
and U1111 (N_1111,In_171,In_1646);
xnor U1112 (N_1112,N_558,N_957);
or U1113 (N_1113,N_597,In_2489);
and U1114 (N_1114,In_1604,N_224);
xnor U1115 (N_1115,In_1935,In_251);
and U1116 (N_1116,In_919,N_412);
or U1117 (N_1117,In_484,In_319);
and U1118 (N_1118,In_1543,N_433);
nand U1119 (N_1119,N_376,N_829);
xnor U1120 (N_1120,N_948,In_2615);
nor U1121 (N_1121,In_1136,In_1754);
nor U1122 (N_1122,In_2150,N_37);
and U1123 (N_1123,In_994,N_609);
and U1124 (N_1124,In_891,In_2829);
and U1125 (N_1125,In_1496,In_1713);
nor U1126 (N_1126,In_1023,In_1484);
xnor U1127 (N_1127,In_2979,N_733);
and U1128 (N_1128,N_822,In_220);
nand U1129 (N_1129,N_884,In_510);
and U1130 (N_1130,In_114,N_965);
nor U1131 (N_1131,N_392,In_1878);
or U1132 (N_1132,In_407,In_282);
or U1133 (N_1133,In_983,N_834);
xor U1134 (N_1134,In_667,In_447);
and U1135 (N_1135,N_354,In_1371);
xnor U1136 (N_1136,In_1378,N_133);
or U1137 (N_1137,In_2859,N_686);
nand U1138 (N_1138,In_2257,In_1125);
nor U1139 (N_1139,In_2655,In_2651);
nand U1140 (N_1140,N_608,In_2687);
or U1141 (N_1141,In_1704,N_835);
xnor U1142 (N_1142,In_2325,In_1556);
and U1143 (N_1143,In_323,In_547);
and U1144 (N_1144,In_156,In_146);
nor U1145 (N_1145,In_926,N_913);
nor U1146 (N_1146,In_1462,N_257);
nand U1147 (N_1147,N_138,In_177);
nand U1148 (N_1148,N_70,In_604);
nand U1149 (N_1149,In_10,N_230);
nor U1150 (N_1150,In_2952,In_1917);
or U1151 (N_1151,N_102,In_1901);
nor U1152 (N_1152,N_466,N_476);
nand U1153 (N_1153,In_948,In_273);
nor U1154 (N_1154,In_1806,In_720);
xnor U1155 (N_1155,In_1591,N_746);
nor U1156 (N_1156,In_976,In_1629);
nor U1157 (N_1157,N_275,In_591);
nand U1158 (N_1158,In_1579,In_2932);
and U1159 (N_1159,In_2635,In_2165);
and U1160 (N_1160,N_423,N_455);
nor U1161 (N_1161,In_2470,In_313);
and U1162 (N_1162,In_1909,In_2800);
and U1163 (N_1163,N_361,N_370);
nor U1164 (N_1164,In_1702,In_1707);
nor U1165 (N_1165,In_93,In_934);
and U1166 (N_1166,In_554,In_2080);
xnor U1167 (N_1167,N_574,N_915);
nand U1168 (N_1168,In_1535,N_337);
nor U1169 (N_1169,In_861,In_443);
xnor U1170 (N_1170,N_743,N_272);
xnor U1171 (N_1171,In_2395,In_2789);
and U1172 (N_1172,N_661,N_210);
and U1173 (N_1173,In_1881,In_2025);
or U1174 (N_1174,N_855,N_860);
nand U1175 (N_1175,N_504,N_266);
nand U1176 (N_1176,In_341,In_985);
or U1177 (N_1177,In_2620,In_1319);
and U1178 (N_1178,In_540,N_199);
or U1179 (N_1179,In_695,In_2203);
and U1180 (N_1180,In_706,N_561);
nor U1181 (N_1181,In_877,In_2425);
and U1182 (N_1182,In_270,In_2763);
nand U1183 (N_1183,In_2057,In_1902);
and U1184 (N_1184,N_373,In_1549);
or U1185 (N_1185,In_1194,In_995);
nand U1186 (N_1186,N_198,N_671);
and U1187 (N_1187,In_1209,N_406);
nand U1188 (N_1188,In_2437,In_2248);
nor U1189 (N_1189,In_2861,N_384);
nor U1190 (N_1190,In_288,N_721);
nor U1191 (N_1191,In_984,N_891);
nand U1192 (N_1192,N_519,N_825);
and U1193 (N_1193,In_801,In_1425);
nor U1194 (N_1194,In_620,N_668);
xnor U1195 (N_1195,N_751,N_643);
nand U1196 (N_1196,N_347,In_1293);
nor U1197 (N_1197,N_615,In_1999);
nand U1198 (N_1198,In_2766,In_1088);
and U1199 (N_1199,N_978,In_915);
and U1200 (N_1200,N_458,N_628);
nor U1201 (N_1201,In_34,In_1814);
xnor U1202 (N_1202,In_1292,In_2793);
and U1203 (N_1203,N_1030,In_2022);
xnor U1204 (N_1204,N_947,In_2295);
and U1205 (N_1205,N_851,N_175);
or U1206 (N_1206,N_896,In_2575);
nand U1207 (N_1207,In_616,In_1413);
xor U1208 (N_1208,N_49,N_191);
or U1209 (N_1209,In_92,In_1102);
nand U1210 (N_1210,N_1045,N_1044);
xor U1211 (N_1211,In_247,In_1651);
xnor U1212 (N_1212,N_549,N_520);
and U1213 (N_1213,N_1001,In_491);
xnor U1214 (N_1214,In_1923,In_2522);
nor U1215 (N_1215,N_768,In_2240);
or U1216 (N_1216,In_1889,In_201);
nor U1217 (N_1217,N_1174,In_409);
or U1218 (N_1218,N_964,In_2363);
xnor U1219 (N_1219,In_2660,N_962);
nand U1220 (N_1220,N_984,In_134);
xor U1221 (N_1221,In_517,In_767);
and U1222 (N_1222,In_1353,In_1461);
and U1223 (N_1223,In_1742,In_1060);
and U1224 (N_1224,In_1555,In_1365);
nand U1225 (N_1225,In_2857,N_654);
or U1226 (N_1226,N_619,In_865);
nand U1227 (N_1227,In_440,N_402);
and U1228 (N_1228,N_987,In_1492);
nor U1229 (N_1229,In_1836,In_1273);
xnor U1230 (N_1230,N_186,In_2754);
and U1231 (N_1231,In_1027,In_1995);
nor U1232 (N_1232,N_71,In_1046);
nand U1233 (N_1233,In_2521,N_495);
xor U1234 (N_1234,N_700,N_580);
and U1235 (N_1235,In_1004,N_73);
xor U1236 (N_1236,N_1011,N_641);
and U1237 (N_1237,N_603,N_1075);
nor U1238 (N_1238,N_415,In_1329);
nor U1239 (N_1239,N_468,N_892);
nand U1240 (N_1240,N_836,In_1015);
or U1241 (N_1241,In_1645,N_1195);
xor U1242 (N_1242,In_1250,In_2226);
nand U1243 (N_1243,N_1114,In_494);
and U1244 (N_1244,In_1641,N_685);
and U1245 (N_1245,In_271,N_1068);
or U1246 (N_1246,In_320,In_157);
or U1247 (N_1247,N_676,In_1831);
and U1248 (N_1248,N_919,N_658);
nand U1249 (N_1249,In_2067,In_1700);
xor U1250 (N_1250,N_688,In_2418);
xnor U1251 (N_1251,In_2079,In_444);
nor U1252 (N_1252,N_101,N_652);
nor U1253 (N_1253,In_2586,N_357);
and U1254 (N_1254,In_2115,In_929);
xnor U1255 (N_1255,In_1411,In_221);
or U1256 (N_1256,In_2433,In_2713);
nor U1257 (N_1257,In_385,In_408);
nand U1258 (N_1258,In_1464,In_2193);
nand U1259 (N_1259,In_2939,In_925);
and U1260 (N_1260,N_445,In_2947);
and U1261 (N_1261,N_1166,N_890);
and U1262 (N_1262,In_2396,N_1173);
and U1263 (N_1263,In_647,N_1094);
and U1264 (N_1264,N_809,In_1156);
and U1265 (N_1265,N_134,In_33);
nor U1266 (N_1266,In_2090,In_1596);
nor U1267 (N_1267,N_1163,N_1164);
nand U1268 (N_1268,In_1093,N_362);
and U1269 (N_1269,In_2495,N_1092);
nand U1270 (N_1270,In_551,In_2547);
or U1271 (N_1271,In_1967,N_557);
nor U1272 (N_1272,N_985,N_385);
xnor U1273 (N_1273,N_225,In_828);
xor U1274 (N_1274,N_662,In_1363);
xor U1275 (N_1275,N_513,N_852);
xnor U1276 (N_1276,N_334,In_1265);
nor U1277 (N_1277,N_1115,In_2820);
xor U1278 (N_1278,In_2630,In_2711);
nor U1279 (N_1279,In_577,In_1627);
and U1280 (N_1280,In_1926,In_1778);
nor U1281 (N_1281,N_728,In_1835);
and U1282 (N_1282,N_900,N_1101);
xnor U1283 (N_1283,N_529,N_403);
xor U1284 (N_1284,In_2591,In_1759);
or U1285 (N_1285,N_1067,N_1054);
and U1286 (N_1286,In_778,N_605);
nor U1287 (N_1287,N_986,N_1187);
nor U1288 (N_1288,In_1900,In_1494);
xnor U1289 (N_1289,In_2938,N_255);
and U1290 (N_1290,N_731,In_1794);
xor U1291 (N_1291,N_887,In_2390);
nand U1292 (N_1292,In_2106,In_1342);
nor U1293 (N_1293,In_1726,In_2748);
nand U1294 (N_1294,N_480,In_238);
nor U1295 (N_1295,N_1197,N_501);
and U1296 (N_1296,In_1701,In_2584);
xor U1297 (N_1297,N_232,N_888);
and U1298 (N_1298,N_1063,In_2407);
nor U1299 (N_1299,In_1521,In_1382);
xor U1300 (N_1300,N_234,In_2188);
nor U1301 (N_1301,N_722,In_826);
nor U1302 (N_1302,N_673,N_1077);
nand U1303 (N_1303,In_1407,N_486);
nor U1304 (N_1304,In_1808,N_1029);
nand U1305 (N_1305,N_217,N_1168);
or U1306 (N_1306,In_2426,N_1132);
nor U1307 (N_1307,In_972,In_700);
or U1308 (N_1308,N_681,In_2479);
nand U1309 (N_1309,In_463,In_813);
and U1310 (N_1310,N_709,N_994);
nand U1311 (N_1311,In_2218,In_548);
nand U1312 (N_1312,In_1932,N_648);
nand U1313 (N_1313,In_67,In_2241);
or U1314 (N_1314,In_1106,In_2553);
xnor U1315 (N_1315,N_1123,N_785);
nand U1316 (N_1316,N_1082,N_754);
or U1317 (N_1317,In_2625,In_1714);
or U1318 (N_1318,N_1014,N_878);
xor U1319 (N_1319,In_680,N_41);
and U1320 (N_1320,In_2348,N_1193);
nor U1321 (N_1321,N_946,N_528);
and U1322 (N_1322,In_2788,In_2765);
nor U1323 (N_1323,N_299,In_2366);
nor U1324 (N_1324,In_1515,In_77);
or U1325 (N_1325,In_1373,N_200);
and U1326 (N_1326,N_116,In_836);
nand U1327 (N_1327,N_323,N_640);
xnor U1328 (N_1328,In_598,In_1020);
and U1329 (N_1329,N_967,In_2834);
xor U1330 (N_1330,In_1308,N_1182);
xnor U1331 (N_1331,In_474,In_1235);
or U1332 (N_1332,In_2473,In_1518);
xnor U1333 (N_1333,In_630,In_1225);
and U1334 (N_1334,In_2132,N_993);
or U1335 (N_1335,In_89,N_1023);
nor U1336 (N_1336,N_411,N_439);
and U1337 (N_1337,In_1180,In_278);
nand U1338 (N_1338,N_522,N_882);
nor U1339 (N_1339,In_1940,N_304);
xor U1340 (N_1340,N_552,In_2459);
nand U1341 (N_1341,In_1402,N_540);
nor U1342 (N_1342,In_2966,N_970);
nor U1343 (N_1343,In_806,In_2965);
nor U1344 (N_1344,In_2004,In_783);
nand U1345 (N_1345,N_263,In_2913);
nand U1346 (N_1346,In_661,In_2701);
and U1347 (N_1347,In_1191,N_846);
and U1348 (N_1348,In_2008,In_689);
nand U1349 (N_1349,In_576,N_0);
and U1350 (N_1350,N_1145,In_1857);
nand U1351 (N_1351,In_1124,In_1531);
xnor U1352 (N_1352,N_249,N_164);
xor U1353 (N_1353,N_1005,In_1499);
and U1354 (N_1354,In_588,In_1637);
nor U1355 (N_1355,In_2246,In_1686);
and U1356 (N_1356,In_2149,N_934);
nand U1357 (N_1357,In_2559,N_908);
or U1358 (N_1358,In_2305,In_1896);
nand U1359 (N_1359,In_1600,N_327);
nor U1360 (N_1360,N_893,In_1844);
and U1361 (N_1361,In_2377,N_1037);
xor U1362 (N_1362,In_879,N_278);
xnor U1363 (N_1363,N_1119,N_1093);
or U1364 (N_1364,N_1026,In_2367);
xor U1365 (N_1365,In_2477,In_998);
nor U1366 (N_1366,In_2904,In_289);
nand U1367 (N_1367,In_1663,N_742);
nand U1368 (N_1368,N_461,In_1867);
nor U1369 (N_1369,N_599,N_1041);
xor U1370 (N_1370,In_1717,In_1789);
nand U1371 (N_1371,N_498,N_749);
xor U1372 (N_1372,In_2583,N_242);
or U1373 (N_1373,In_2698,In_2216);
or U1374 (N_1374,In_1618,In_1080);
xnor U1375 (N_1375,N_267,N_928);
nor U1376 (N_1376,In_2742,In_457);
xor U1377 (N_1377,In_2064,N_258);
xnor U1378 (N_1378,N_727,In_838);
xor U1379 (N_1379,N_585,In_1263);
nor U1380 (N_1380,In_2280,In_290);
nand U1381 (N_1381,N_799,N_350);
nand U1382 (N_1382,In_2814,In_360);
or U1383 (N_1383,In_1291,In_2632);
xnor U1384 (N_1384,In_1733,In_808);
and U1385 (N_1385,In_2832,In_2260);
nor U1386 (N_1386,N_487,In_2500);
or U1387 (N_1387,In_2337,In_2243);
xor U1388 (N_1388,N_801,In_44);
xor U1389 (N_1389,In_1880,In_1458);
nor U1390 (N_1390,N_1150,In_398);
nand U1391 (N_1391,N_625,N_936);
nand U1392 (N_1392,In_585,In_2448);
nor U1393 (N_1393,In_821,In_486);
nor U1394 (N_1394,N_1117,In_1959);
and U1395 (N_1395,In_2572,In_1304);
nor U1396 (N_1396,N_1007,N_1060);
nor U1397 (N_1397,N_1190,In_1045);
or U1398 (N_1398,In_1777,In_216);
and U1399 (N_1399,N_214,In_1886);
xor U1400 (N_1400,N_1142,N_128);
and U1401 (N_1401,In_109,N_215);
and U1402 (N_1402,N_1088,In_2249);
nor U1403 (N_1403,N_1089,In_1887);
or U1404 (N_1404,In_2224,N_1381);
or U1405 (N_1405,In_2951,N_792);
xor U1406 (N_1406,In_2917,In_761);
nor U1407 (N_1407,In_1825,N_1249);
xnor U1408 (N_1408,In_2244,In_2551);
nor U1409 (N_1409,N_650,N_1396);
or U1410 (N_1410,In_724,N_930);
or U1411 (N_1411,N_100,N_844);
xnor U1412 (N_1412,N_1313,In_533);
and U1413 (N_1413,In_525,In_1863);
nor U1414 (N_1414,In_2450,In_2362);
and U1415 (N_1415,N_396,In_2475);
nor U1416 (N_1416,N_481,In_345);
xnor U1417 (N_1417,N_1189,In_2445);
or U1418 (N_1418,N_303,In_2567);
and U1419 (N_1419,In_608,N_976);
or U1420 (N_1420,N_1278,N_756);
xor U1421 (N_1421,N_308,In_1166);
nand U1422 (N_1422,In_88,N_464);
nand U1423 (N_1423,N_491,N_636);
nor U1424 (N_1424,In_797,N_706);
nor U1425 (N_1425,In_387,N_1218);
nor U1426 (N_1426,N_1212,N_29);
nand U1427 (N_1427,N_1346,N_973);
nand U1428 (N_1428,N_759,N_1289);
xnor U1429 (N_1429,In_1664,N_774);
or U1430 (N_1430,N_1216,N_975);
nand U1431 (N_1431,In_2886,In_14);
or U1432 (N_1432,N_581,In_54);
nand U1433 (N_1433,In_2613,N_1253);
nor U1434 (N_1434,N_1245,In_1567);
xor U1435 (N_1435,In_1192,N_196);
and U1436 (N_1436,In_0,N_1273);
nor U1437 (N_1437,In_116,In_567);
nand U1438 (N_1438,N_87,In_2603);
nor U1439 (N_1439,N_69,N_505);
nor U1440 (N_1440,In_2524,In_932);
or U1441 (N_1441,In_1647,N_696);
and U1442 (N_1442,In_1720,In_586);
nor U1443 (N_1443,N_270,In_2509);
xnor U1444 (N_1444,N_943,In_1100);
and U1445 (N_1445,N_295,In_2440);
nor U1446 (N_1446,In_1358,In_2706);
or U1447 (N_1447,N_499,N_194);
xor U1448 (N_1448,In_2182,N_264);
or U1449 (N_1449,In_372,N_1387);
or U1450 (N_1450,In_2975,N_621);
xnor U1451 (N_1451,In_2875,In_534);
or U1452 (N_1452,In_1721,N_1131);
or U1453 (N_1453,N_1285,N_1034);
and U1454 (N_1454,In_544,In_1200);
nand U1455 (N_1455,In_1516,In_1522);
xor U1456 (N_1456,N_371,In_2460);
nand U1457 (N_1457,N_624,In_2936);
xnor U1458 (N_1458,In_2563,N_707);
nor U1459 (N_1459,N_1084,In_2846);
nor U1460 (N_1460,In_535,N_1390);
or U1461 (N_1461,N_594,N_831);
or U1462 (N_1462,In_1773,In_779);
or U1463 (N_1463,N_1327,N_634);
and U1464 (N_1464,N_1181,In_1404);
or U1465 (N_1465,N_1250,N_1279);
nor U1466 (N_1466,In_2751,In_1339);
nor U1467 (N_1467,In_2177,In_2339);
or U1468 (N_1468,N_1307,In_3);
or U1469 (N_1469,In_144,In_1446);
nand U1470 (N_1470,N_1363,N_1252);
nor U1471 (N_1471,In_751,N_1019);
nand U1472 (N_1472,N_1036,In_327);
nor U1473 (N_1473,In_208,N_1204);
nand U1474 (N_1474,N_1233,In_22);
nand U1475 (N_1475,In_1074,N_1107);
nand U1476 (N_1476,N_1340,N_1172);
and U1477 (N_1477,N_1116,In_981);
nor U1478 (N_1478,In_2462,In_1110);
nand U1479 (N_1479,In_370,N_1240);
nand U1480 (N_1480,In_1812,In_1639);
and U1481 (N_1481,N_1090,In_2030);
and U1482 (N_1482,In_1668,N_544);
nor U1483 (N_1483,N_1299,N_1065);
and U1484 (N_1484,N_938,In_1299);
nor U1485 (N_1485,In_1938,In_1313);
or U1486 (N_1486,In_363,N_858);
and U1487 (N_1487,N_729,In_155);
xnor U1488 (N_1488,N_826,N_168);
or U1489 (N_1489,N_1316,In_1985);
and U1490 (N_1490,In_1309,In_2774);
xor U1491 (N_1491,In_1169,N_1003);
xnor U1492 (N_1492,In_2623,N_1122);
xnor U1493 (N_1493,N_969,In_2274);
or U1494 (N_1494,In_2601,In_1705);
and U1495 (N_1495,N_838,In_1774);
nor U1496 (N_1496,In_2085,In_717);
or U1497 (N_1497,In_2873,N_1269);
or U1498 (N_1498,N_1322,In_2347);
or U1499 (N_1499,N_1179,In_2478);
or U1500 (N_1500,N_1392,In_336);
xnor U1501 (N_1501,N_1207,In_1833);
nor U1502 (N_1502,In_2238,N_1006);
xor U1503 (N_1503,N_1024,N_980);
nand U1504 (N_1504,N_770,N_752);
and U1505 (N_1505,N_679,In_102);
or U1506 (N_1506,N_567,In_302);
and U1507 (N_1507,N_764,N_261);
nor U1508 (N_1508,N_1356,In_1993);
or U1509 (N_1509,N_952,In_2607);
nor U1510 (N_1510,N_1033,N_918);
xnor U1511 (N_1511,In_777,N_77);
nor U1512 (N_1512,N_95,In_800);
xnor U1513 (N_1513,N_1056,In_571);
xnor U1514 (N_1514,N_508,N_237);
nand U1515 (N_1515,In_1186,N_995);
and U1516 (N_1516,In_2467,N_1010);
and U1517 (N_1517,In_957,N_1399);
xor U1518 (N_1518,N_518,In_1862);
and U1519 (N_1519,In_1347,In_1976);
or U1520 (N_1520,In_841,N_39);
nor U1521 (N_1521,In_1552,N_157);
or U1522 (N_1522,In_677,N_1383);
and U1523 (N_1523,In_1151,In_1732);
or U1524 (N_1524,In_699,N_389);
nand U1525 (N_1525,In_2212,In_1164);
or U1526 (N_1526,In_1030,In_758);
or U1527 (N_1527,N_924,N_1329);
nand U1528 (N_1528,N_131,N_1379);
and U1529 (N_1529,In_260,In_745);
nor U1530 (N_1530,N_1022,In_2983);
and U1531 (N_1531,In_2494,N_394);
or U1532 (N_1532,In_2110,In_1029);
or U1533 (N_1533,N_604,In_2764);
nor U1534 (N_1534,In_965,N_546);
nor U1535 (N_1535,In_2808,N_811);
xor U1536 (N_1536,In_563,In_2672);
xnor U1537 (N_1537,In_2828,In_245);
xnor U1538 (N_1538,N_208,In_759);
or U1539 (N_1539,N_1248,N_500);
or U1540 (N_1540,N_328,N_36);
nor U1541 (N_1541,In_1547,In_2327);
or U1542 (N_1542,In_1077,In_901);
and U1543 (N_1543,N_1357,N_786);
xnor U1544 (N_1544,N_803,In_249);
and U1545 (N_1545,N_442,In_1028);
xor U1546 (N_1546,N_869,In_1715);
xor U1547 (N_1547,In_702,N_1342);
or U1548 (N_1548,N_1028,N_1059);
or U1549 (N_1549,N_1157,In_1851);
nand U1550 (N_1550,N_956,N_156);
nand U1551 (N_1551,In_1904,N_63);
nor U1552 (N_1552,In_787,In_367);
and U1553 (N_1553,N_503,N_143);
nand U1554 (N_1554,N_1221,N_1306);
nor U1555 (N_1555,In_2229,In_1914);
and U1556 (N_1556,N_514,In_2268);
nor U1557 (N_1557,In_557,N_1319);
nor U1558 (N_1558,In_231,N_1228);
nand U1559 (N_1559,N_901,In_73);
xor U1560 (N_1560,In_2642,N_88);
nand U1561 (N_1561,In_2439,N_1276);
nand U1562 (N_1562,N_269,In_330);
nand U1563 (N_1563,N_397,In_686);
nand U1564 (N_1564,In_1258,N_981);
nand U1565 (N_1565,N_872,N_150);
nor U1566 (N_1566,N_1018,In_748);
or U1567 (N_1567,In_2792,In_30);
or U1568 (N_1568,N_1149,N_879);
nand U1569 (N_1569,N_1137,In_514);
nor U1570 (N_1570,N_715,In_1610);
xnor U1571 (N_1571,In_854,In_365);
or U1572 (N_1572,In_2406,N_1328);
or U1573 (N_1573,N_1105,N_1311);
and U1574 (N_1574,In_62,N_516);
nor U1575 (N_1575,In_2831,N_1049);
and U1576 (N_1576,N_1154,N_904);
xnor U1577 (N_1577,N_1310,N_791);
or U1578 (N_1578,N_1219,In_2971);
or U1579 (N_1579,In_2989,N_193);
xnor U1580 (N_1580,In_1073,N_1);
or U1581 (N_1581,N_1275,In_1356);
and U1582 (N_1582,In_1830,N_1009);
xor U1583 (N_1583,N_1027,N_470);
xor U1584 (N_1584,N_1042,N_1295);
and U1585 (N_1585,In_1908,In_1614);
or U1586 (N_1586,In_584,N_1158);
nor U1587 (N_1587,N_1135,In_118);
or U1588 (N_1588,N_1246,In_332);
nor U1589 (N_1589,N_183,N_422);
nand U1590 (N_1590,N_1264,N_1083);
nor U1591 (N_1591,In_347,N_425);
or U1592 (N_1592,In_2344,In_1991);
nand U1593 (N_1593,In_974,N_778);
nor U1594 (N_1594,N_828,In_612);
nand U1595 (N_1595,In_2674,In_1448);
nor U1596 (N_1596,In_1671,In_204);
and U1597 (N_1597,In_1355,N_827);
nor U1598 (N_1598,In_2109,N_1143);
nand U1599 (N_1599,N_895,In_1525);
or U1600 (N_1600,In_202,In_2364);
nand U1601 (N_1601,In_2102,In_839);
xnor U1602 (N_1602,N_1087,In_1784);
or U1603 (N_1603,N_141,N_1466);
and U1604 (N_1604,In_2634,N_1473);
nor U1605 (N_1605,N_1236,In_909);
xnor U1606 (N_1606,In_1010,N_982);
xnor U1607 (N_1607,In_297,In_1395);
xor U1608 (N_1608,N_849,In_709);
nand U1609 (N_1609,N_732,N_909);
or U1610 (N_1610,In_1283,N_1434);
and U1611 (N_1611,In_1566,N_139);
nand U1612 (N_1612,In_1601,N_833);
or U1613 (N_1613,In_644,In_2517);
nor U1614 (N_1614,N_1568,N_145);
or U1615 (N_1615,In_2867,In_1734);
nor U1616 (N_1616,In_2179,In_1670);
nor U1617 (N_1617,In_1978,N_367);
nor U1618 (N_1618,N_1368,In_1681);
or U1619 (N_1619,N_1589,In_1410);
and U1620 (N_1620,In_1199,N_738);
nand U1621 (N_1621,N_883,N_929);
nand U1622 (N_1622,N_62,In_1321);
and U1623 (N_1623,In_1489,N_166);
nand U1624 (N_1624,In_293,N_1479);
xnor U1625 (N_1625,N_1177,N_1530);
nand U1626 (N_1626,N_808,N_699);
nand U1627 (N_1627,N_1331,N_684);
nand U1628 (N_1628,N_1120,In_2002);
xor U1629 (N_1629,N_657,N_1572);
nor U1630 (N_1630,In_2040,N_1533);
nand U1631 (N_1631,In_2617,In_1451);
xnor U1632 (N_1632,In_874,N_856);
xnor U1633 (N_1633,N_1039,In_2805);
xor U1634 (N_1634,N_1208,In_618);
nand U1635 (N_1635,N_1433,N_1152);
xnor U1636 (N_1636,In_1716,In_1576);
nor U1637 (N_1637,In_1877,N_620);
xnor U1638 (N_1638,In_698,In_2273);
or U1639 (N_1639,N_868,N_1508);
and U1640 (N_1640,N_1526,N_907);
or U1641 (N_1641,N_1543,N_1004);
xor U1642 (N_1642,N_958,N_1557);
and U1643 (N_1643,In_2684,N_1282);
nand U1644 (N_1644,N_1231,N_1575);
and U1645 (N_1645,In_480,In_1635);
xnor U1646 (N_1646,In_2357,In_2181);
and U1647 (N_1647,N_1170,In_1114);
and U1648 (N_1648,In_2953,In_2298);
or U1649 (N_1649,In_614,In_2680);
nor U1650 (N_1650,In_9,In_1167);
nand U1651 (N_1651,In_1352,In_1231);
and U1652 (N_1652,In_1008,N_375);
xor U1653 (N_1653,In_1044,In_1031);
nand U1654 (N_1654,N_1214,In_2026);
or U1655 (N_1655,N_1565,N_926);
or U1656 (N_1656,N_125,In_81);
xnor U1657 (N_1657,In_2519,In_672);
xnor U1658 (N_1658,In_85,N_1244);
or U1659 (N_1659,N_753,N_1382);
nor U1660 (N_1660,In_2472,N_479);
nand U1661 (N_1661,In_933,N_1418);
nand U1662 (N_1662,In_1658,In_590);
nand U1663 (N_1663,N_1496,In_197);
or U1664 (N_1664,N_506,In_626);
nand U1665 (N_1665,In_2887,In_920);
nor U1666 (N_1666,N_1021,In_637);
and U1667 (N_1667,N_391,N_1303);
or U1668 (N_1668,In_2949,N_1456);
nand U1669 (N_1669,N_1393,In_318);
xnor U1670 (N_1670,N_1354,N_723);
or U1671 (N_1671,N_187,In_2888);
xnor U1672 (N_1672,N_1472,In_2794);
or U1673 (N_1673,In_244,In_2361);
or U1674 (N_1674,In_527,In_860);
and U1675 (N_1675,N_1171,N_159);
nor U1676 (N_1676,In_2158,N_179);
nor U1677 (N_1677,N_1203,In_2633);
or U1678 (N_1678,In_1798,In_1399);
nand U1679 (N_1679,In_1998,In_734);
nor U1680 (N_1680,N_1450,In_773);
xnor U1681 (N_1681,N_1153,N_656);
or U1682 (N_1682,N_905,N_761);
or U1683 (N_1683,In_2018,In_2876);
nand U1684 (N_1684,N_968,In_754);
nor U1685 (N_1685,N_67,In_2094);
nand U1686 (N_1686,In_2560,N_556);
nor U1687 (N_1687,N_1258,N_1238);
and U1688 (N_1688,In_1238,In_2566);
and U1689 (N_1689,N_1465,In_2801);
xor U1690 (N_1690,In_1264,In_511);
xor U1691 (N_1691,N_1071,In_2590);
and U1692 (N_1692,N_1389,N_1370);
and U1693 (N_1693,N_1224,N_1569);
nor U1694 (N_1694,N_859,N_1523);
and U1695 (N_1695,N_1000,N_1391);
or U1696 (N_1696,N_812,N_1320);
xor U1697 (N_1697,N_1527,N_843);
nor U1698 (N_1698,In_1229,In_401);
nor U1699 (N_1699,N_1415,N_1337);
nor U1700 (N_1700,In_701,In_1147);
nor U1701 (N_1701,In_1234,In_2314);
nand U1702 (N_1702,In_2813,In_2729);
xor U1703 (N_1703,N_1542,N_1043);
nor U1704 (N_1704,N_1175,N_922);
or U1705 (N_1705,N_1262,In_186);
nor U1706 (N_1706,N_989,In_104);
xnor U1707 (N_1707,N_207,N_1375);
xor U1708 (N_1708,In_2422,N_1429);
xnor U1709 (N_1709,N_1191,N_1482);
and U1710 (N_1710,In_2637,N_1257);
nand U1711 (N_1711,N_598,In_539);
and U1712 (N_1712,In_842,N_777);
or U1713 (N_1713,N_11,In_24);
and U1714 (N_1714,N_1057,N_1499);
xor U1715 (N_1715,In_154,In_280);
nand U1716 (N_1716,N_1593,N_575);
or U1717 (N_1717,N_708,In_162);
nor U1718 (N_1718,N_1165,In_2919);
or U1719 (N_1719,N_1511,In_129);
nand U1720 (N_1720,N_313,N_1096);
xor U1721 (N_1721,N_560,In_452);
or U1722 (N_1722,N_399,In_1117);
nand U1723 (N_1723,In_65,N_1442);
and U1724 (N_1724,N_1560,N_1571);
or U1725 (N_1725,In_936,N_127);
nand U1726 (N_1726,N_1529,In_1854);
and U1727 (N_1727,In_2201,In_1295);
nor U1728 (N_1728,N_1545,In_918);
nor U1729 (N_1729,N_1330,N_959);
or U1730 (N_1730,In_2530,N_349);
nand U1731 (N_1731,N_1247,N_921);
and U1732 (N_1732,N_711,In_2056);
nand U1733 (N_1733,N_806,N_961);
nor U1734 (N_1734,N_1167,In_483);
or U1735 (N_1735,In_2720,N_1076);
xnor U1736 (N_1736,N_1104,N_1078);
xnor U1737 (N_1737,In_1827,In_2858);
nor U1738 (N_1738,In_816,N_1349);
or U1739 (N_1739,N_1326,In_2622);
nor U1740 (N_1740,N_381,N_1226);
nor U1741 (N_1741,N_1437,N_265);
and U1742 (N_1742,N_1124,N_773);
nor U1743 (N_1743,In_522,N_951);
nor U1744 (N_1744,In_968,N_475);
xnor U1745 (N_1745,In_723,N_1317);
xnor U1746 (N_1746,In_999,N_1180);
and U1747 (N_1747,N_853,In_805);
and U1748 (N_1748,In_2082,N_1294);
or U1749 (N_1749,N_34,In_2589);
xor U1750 (N_1750,N_1485,In_2318);
or U1751 (N_1751,N_38,In_589);
or U1752 (N_1752,N_473,In_2356);
and U1753 (N_1753,N_568,N_472);
xor U1754 (N_1754,N_1352,In_656);
or U1755 (N_1755,In_2202,N_579);
nand U1756 (N_1756,N_1364,N_1520);
xnor U1757 (N_1757,N_307,In_2749);
or U1758 (N_1758,In_2677,N_1314);
nand U1759 (N_1759,N_655,N_1424);
or U1760 (N_1760,N_1386,N_460);
or U1761 (N_1761,N_129,N_20);
nand U1762 (N_1762,N_1491,N_691);
nor U1763 (N_1763,N_32,N_1136);
or U1764 (N_1764,N_854,In_810);
or U1765 (N_1765,In_660,N_613);
nor U1766 (N_1766,In_858,In_2139);
and U1767 (N_1767,In_1530,N_1409);
xnor U1768 (N_1768,In_2878,In_1609);
nor U1769 (N_1769,In_17,In_2488);
xnor U1770 (N_1770,N_1256,N_1467);
and U1771 (N_1771,N_1483,N_1209);
or U1772 (N_1772,N_1332,N_1596);
or U1773 (N_1773,In_132,N_1270);
and U1774 (N_1774,In_2027,N_693);
or U1775 (N_1775,N_610,N_1528);
and U1776 (N_1776,In_348,In_1970);
nand U1777 (N_1777,In_2421,N_212);
xnor U1778 (N_1778,In_91,N_923);
or U1779 (N_1779,N_1595,N_1344);
nor U1780 (N_1780,In_235,N_1298);
nor U1781 (N_1781,N_1373,N_983);
xnor U1782 (N_1782,N_47,N_1064);
and U1783 (N_1783,N_963,In_1022);
nand U1784 (N_1784,In_2251,In_911);
and U1785 (N_1785,N_937,N_1015);
and U1786 (N_1786,In_2154,In_1554);
or U1787 (N_1787,N_914,N_939);
xor U1788 (N_1788,N_413,N_353);
or U1789 (N_1789,N_1532,In_1132);
nand U1790 (N_1790,N_1414,N_1497);
and U1791 (N_1791,N_690,In_1984);
or U1792 (N_1792,N_1050,N_493);
and U1793 (N_1793,In_2722,In_2641);
nand U1794 (N_1794,In_1249,In_364);
xor U1795 (N_1795,N_894,In_1852);
xnor U1796 (N_1796,In_1444,N_282);
xnor U1797 (N_1797,In_2956,N_1052);
or U1798 (N_1798,N_429,N_1498);
nand U1799 (N_1799,N_564,N_418);
nand U1800 (N_1800,N_1619,N_702);
nand U1801 (N_1801,N_1770,In_785);
xor U1802 (N_1802,In_1335,N_1582);
nand U1803 (N_1803,In_2582,N_1397);
and U1804 (N_1804,N_1345,In_2125);
and U1805 (N_1805,In_266,N_1435);
or U1806 (N_1806,In_1988,N_1121);
nor U1807 (N_1807,N_1035,N_566);
xnor U1808 (N_1808,In_2435,N_1795);
xor U1809 (N_1809,In_1677,N_1098);
or U1810 (N_1810,N_1731,In_175);
or U1811 (N_1811,N_1645,N_1425);
nor U1812 (N_1812,N_942,N_974);
nand U1813 (N_1813,In_1207,N_1446);
xnor U1814 (N_1814,In_2920,In_2183);
xor U1815 (N_1815,In_1148,N_1367);
xor U1816 (N_1816,N_1051,N_1601);
nand U1817 (N_1817,N_999,N_1685);
nor U1818 (N_1818,N_1797,In_326);
xor U1819 (N_1819,N_97,N_496);
nor U1820 (N_1820,In_1868,N_1405);
nand U1821 (N_1821,N_1427,In_2705);
xnor U1822 (N_1822,N_1506,N_1355);
or U1823 (N_1823,In_1007,In_2402);
xor U1824 (N_1824,N_823,N_120);
xor U1825 (N_1825,In_382,N_1680);
nor U1826 (N_1826,N_1524,In_2062);
nor U1827 (N_1827,N_1099,N_1111);
or U1828 (N_1828,N_663,In_916);
or U1829 (N_1829,In_2258,In_380);
xor U1830 (N_1830,In_978,N_1505);
or U1831 (N_1831,In_2003,N_211);
or U1832 (N_1832,In_2915,N_48);
and U1833 (N_1833,N_800,In_2797);
or U1834 (N_1834,N_713,N_1283);
and U1835 (N_1835,N_1759,In_256);
nor U1836 (N_1836,N_312,N_972);
and U1837 (N_1837,N_1070,N_885);
nor U1838 (N_1838,In_176,N_1302);
xnor U1839 (N_1839,In_351,In_546);
nor U1840 (N_1840,N_1564,In_1633);
nand U1841 (N_1841,N_1449,In_2389);
or U1842 (N_1842,N_1750,N_1790);
xor U1843 (N_1843,In_481,N_1159);
nand U1844 (N_1844,N_725,N_1438);
or U1845 (N_1845,In_68,N_343);
nand U1846 (N_1846,N_1678,In_133);
xor U1847 (N_1847,N_1764,N_760);
and U1848 (N_1848,N_1535,In_2901);
nor U1849 (N_1849,In_187,In_2758);
xor U1850 (N_1850,In_2017,N_1100);
nand U1851 (N_1851,N_1741,N_730);
nor U1852 (N_1852,In_1274,N_1614);
nor U1853 (N_1853,In_1930,N_1640);
nand U1854 (N_1854,In_1519,N_359);
xor U1855 (N_1855,N_1488,N_1672);
or U1856 (N_1856,In_907,N_1586);
xnor U1857 (N_1857,In_898,N_1176);
or U1858 (N_1858,N_781,N_329);
nor U1859 (N_1859,In_2577,N_1551);
or U1860 (N_1860,N_865,N_1610);
xor U1861 (N_1861,N_1268,N_1369);
or U1862 (N_1862,In_2282,In_1804);
nor U1863 (N_1863,N_977,N_1155);
nand U1864 (N_1864,N_1468,In_1491);
nor U1865 (N_1865,In_740,N_906);
nand U1866 (N_1866,In_2381,N_306);
nand U1867 (N_1867,N_15,N_1760);
and U1868 (N_1868,N_1738,N_1724);
xor U1869 (N_1869,N_1492,N_436);
nand U1870 (N_1870,N_17,In_2543);
and U1871 (N_1871,N_1730,In_1241);
nor U1872 (N_1872,N_1507,In_2656);
or U1873 (N_1873,N_1786,In_1828);
and U1874 (N_1874,N_1066,N_1277);
xnor U1875 (N_1875,N_1200,In_713);
or U1876 (N_1876,N_1243,N_1623);
nor U1877 (N_1877,N_1689,In_519);
nand U1878 (N_1878,N_291,N_1215);
nand U1879 (N_1879,In_2346,In_1142);
xnor U1880 (N_1880,N_1732,N_1146);
xor U1881 (N_1881,N_1301,N_189);
and U1882 (N_1882,In_2512,N_1509);
nand U1883 (N_1883,N_740,N_1148);
xor U1884 (N_1884,In_1563,N_1350);
xor U1885 (N_1885,In_1317,In_2036);
nor U1886 (N_1886,N_630,N_1737);
and U1887 (N_1887,N_453,In_386);
xor U1888 (N_1888,N_195,N_1549);
or U1889 (N_1889,N_644,N_757);
nand U1890 (N_1890,In_1478,In_1508);
xor U1891 (N_1891,N_1341,In_2558);
and U1892 (N_1892,N_1799,N_1254);
and U1893 (N_1893,In_1345,N_1792);
xor U1894 (N_1894,In_2428,N_1630);
nand U1895 (N_1895,In_1692,N_1108);
nand U1896 (N_1896,In_1128,In_2262);
nor U1897 (N_1897,N_1227,N_1727);
nand U1898 (N_1898,In_2294,N_1380);
xor U1899 (N_1899,N_526,N_798);
xor U1900 (N_1900,In_1624,In_2544);
nor U1901 (N_1901,In_581,N_862);
nand U1902 (N_1902,In_2540,In_194);
and U1903 (N_1903,In_1290,N_1398);
and U1904 (N_1904,N_600,N_1156);
xor U1905 (N_1905,In_512,In_1424);
xnor U1906 (N_1906,N_1550,In_1037);
xnor U1907 (N_1907,In_2176,N_1462);
nand U1908 (N_1908,N_1413,In_417);
or U1909 (N_1909,In_1564,N_1522);
and U1910 (N_1910,In_136,N_614);
or U1911 (N_1911,N_1649,N_1734);
nor U1912 (N_1912,N_1284,N_790);
and U1913 (N_1913,N_1774,In_792);
and U1914 (N_1914,N_1772,N_1681);
nand U1915 (N_1915,N_1280,N_1217);
xnor U1916 (N_1916,N_784,N_1016);
or U1917 (N_1917,N_65,N_955);
nor U1918 (N_1918,N_1079,N_1494);
nor U1919 (N_1919,N_1744,N_1255);
nor U1920 (N_1920,In_847,In_795);
xnor U1921 (N_1921,In_807,N_1073);
or U1922 (N_1922,In_2309,N_821);
nor U1923 (N_1923,In_2370,N_665);
xnor U1924 (N_1924,N_533,N_719);
or U1925 (N_1925,In_1964,In_2019);
xor U1926 (N_1926,N_1476,In_28);
xnor U1927 (N_1927,N_554,N_1272);
and U1928 (N_1928,N_1118,N_701);
nor U1929 (N_1929,N_1133,N_1223);
and U1930 (N_1930,In_992,In_1879);
xnor U1931 (N_1931,N_807,In_160);
nand U1932 (N_1932,In_2074,N_1430);
xnor U1933 (N_1933,In_2029,N_659);
and U1934 (N_1934,N_1080,In_2480);
and U1935 (N_1935,N_1404,N_1703);
and U1936 (N_1936,N_1038,In_2443);
or U1937 (N_1937,In_682,N_1141);
and U1938 (N_1938,N_1017,In_2333);
and U1939 (N_1939,In_1903,In_2006);
nand U1940 (N_1940,N_1686,N_1635);
and U1941 (N_1941,In_1958,N_1721);
nor U1942 (N_1942,In_1315,N_446);
nor U1943 (N_1943,N_1745,In_269);
nor U1944 (N_1944,N_582,N_1102);
or U1945 (N_1945,N_1241,N_1714);
and U1946 (N_1946,N_1220,In_762);
xnor U1947 (N_1947,N_1235,N_1725);
xnor U1948 (N_1948,N_1371,N_1647);
nor U1949 (N_1949,N_1566,In_291);
xor U1950 (N_1950,N_1534,N_1766);
or U1951 (N_1951,In_2285,In_809);
xor U1952 (N_1952,N_1583,In_229);
nand U1953 (N_1953,N_1361,In_1969);
nor U1954 (N_1954,In_1883,In_885);
nor U1955 (N_1955,N_675,In_716);
or U1956 (N_1956,N_1715,N_1334);
and U1957 (N_1957,In_697,N_1338);
nand U1958 (N_1958,In_52,N_1682);
nor U1959 (N_1959,In_2141,In_2234);
xor U1960 (N_1960,In_1239,In_1942);
nand U1961 (N_1961,N_348,N_1581);
nor U1962 (N_1962,N_1785,In_693);
nand U1963 (N_1963,N_881,In_1680);
xor U1964 (N_1964,N_1463,N_18);
xnor U1965 (N_1965,In_497,N_27);
nand U1966 (N_1966,In_645,N_1698);
and U1967 (N_1967,N_1723,In_1119);
or U1968 (N_1968,N_1567,N_1325);
or U1969 (N_1969,N_443,N_1490);
xor U1970 (N_1970,In_1763,N_54);
and U1971 (N_1971,N_1756,N_1659);
or U1972 (N_1972,N_1454,N_1128);
and U1973 (N_1973,N_1705,N_1426);
xor U1974 (N_1974,In_2527,N_1587);
and U1975 (N_1975,N_795,N_1336);
nand U1976 (N_1976,N_235,N_1169);
or U1977 (N_1977,N_1662,N_452);
nor U1978 (N_1978,N_1777,In_2270);
xnor U1979 (N_1979,N_1525,In_500);
or U1980 (N_1980,In_2998,In_1957);
nand U1981 (N_1981,N_1638,N_204);
and U1982 (N_1982,N_103,N_1109);
nand U1983 (N_1983,In_632,N_182);
xnor U1984 (N_1984,In_1925,In_2780);
nor U1985 (N_1985,N_121,In_749);
or U1986 (N_1986,N_1561,N_1608);
nand U1987 (N_1987,N_1787,N_1002);
and U1988 (N_1988,N_596,N_763);
nor U1989 (N_1989,N_1627,In_2351);
nand U1990 (N_1990,N_1144,In_20);
nand U1991 (N_1991,In_2250,N_1713);
nor U1992 (N_1992,N_1451,N_848);
nand U1993 (N_1993,N_1707,In_973);
and U1994 (N_1994,N_1376,In_846);
nor U1995 (N_1995,N_1666,N_992);
and U1996 (N_1996,In_521,N_5);
xnor U1997 (N_1997,N_1594,N_1213);
or U1998 (N_1998,In_2175,N_51);
nand U1999 (N_1999,N_144,In_2760);
nor U2000 (N_2000,In_2009,N_1694);
or U2001 (N_2001,In_2686,In_1181);
xnor U2002 (N_2002,N_1964,N_1198);
xor U2003 (N_2003,N_1824,N_1445);
or U2004 (N_2004,N_1973,N_1539);
and U2005 (N_2005,In_789,N_1834);
or U2006 (N_2006,N_1471,N_1151);
xor U2007 (N_2007,In_2600,N_927);
and U2008 (N_2008,N_1267,N_1970);
nand U2009 (N_2009,In_1560,N_1374);
and U2010 (N_2010,N_779,N_1884);
or U2011 (N_2011,N_1259,N_1706);
or U2012 (N_2012,N_1504,In_597);
nand U2013 (N_2013,N_1394,N_841);
nor U2014 (N_2014,N_1953,N_1646);
and U2015 (N_2015,N_1554,N_1654);
xnor U2016 (N_2016,In_2968,N_342);
or U2017 (N_2017,N_1576,In_2940);
and U2018 (N_2018,N_117,N_1606);
nor U2019 (N_2019,N_1675,In_1849);
and U2020 (N_2020,N_1072,N_1905);
and U2021 (N_2021,N_787,N_818);
xor U2022 (N_2022,N_588,N_471);
nand U2023 (N_2023,N_1684,In_424);
xor U2024 (N_2024,In_1551,N_1962);
nand U2025 (N_2025,N_1989,In_1161);
xnor U2026 (N_2026,N_1924,In_2626);
nor U2027 (N_2027,N_920,N_1263);
and U2028 (N_2028,In_2556,N_1712);
xor U2029 (N_2029,N_716,N_870);
or U2030 (N_2030,In_908,N_1271);
nor U2031 (N_2031,In_1712,N_1829);
nor U2032 (N_2032,N_875,N_123);
xnor U2033 (N_2033,N_1733,N_1802);
nand U2034 (N_2034,N_880,N_1260);
nand U2035 (N_2035,N_1883,N_1911);
nand U2036 (N_2036,In_331,In_1441);
nor U2037 (N_2037,N_692,In_429);
or U2038 (N_2038,N_1881,N_1086);
nor U2039 (N_2039,In_553,N_155);
nand U2040 (N_2040,In_2990,N_1676);
nand U2041 (N_2041,N_1600,In_2326);
and U2042 (N_2042,N_1147,In_462);
nand U2043 (N_2043,N_250,In_1334);
nand U2044 (N_2044,In_1279,In_804);
nor U2045 (N_2045,N_576,In_691);
nand U2046 (N_2046,N_1867,In_1431);
and U2047 (N_2047,N_616,In_2496);
or U2048 (N_2048,N_1847,N_1958);
nand U2049 (N_2049,N_1826,In_2075);
or U2050 (N_2050,N_1673,N_1910);
and U2051 (N_2051,N_1455,N_1997);
nor U2052 (N_2052,N_830,In_304);
nor U2053 (N_2053,N_1232,In_2790);
and U2054 (N_2054,In_1230,N_804);
nand U2055 (N_2055,N_666,N_1555);
nand U2056 (N_2056,N_220,In_2863);
xor U2057 (N_2057,In_2991,N_1679);
nand U2058 (N_2058,In_971,In_2451);
nor U2059 (N_2059,N_1487,In_2573);
xnor U2060 (N_2060,N_724,N_1613);
and U2061 (N_2061,N_1584,In_1779);
or U2062 (N_2062,N_1692,N_507);
nor U2063 (N_2063,N_775,N_1993);
and U2064 (N_2064,In_2604,N_612);
xor U2065 (N_2065,In_2420,N_1819);
xor U2066 (N_2066,In_739,In_1634);
nor U2067 (N_2067,N_1184,N_1878);
nand U2068 (N_2068,N_1791,In_2086);
nor U2069 (N_2069,N_1751,In_1105);
xnor U2070 (N_2070,N_1814,N_1753);
and U2071 (N_2071,N_1667,N_1605);
nor U2072 (N_2072,N_553,N_1968);
or U2073 (N_2073,In_1337,In_1501);
or U2074 (N_2074,In_2771,N_1178);
or U2075 (N_2075,N_1477,In_843);
xor U2076 (N_2076,N_1835,N_1932);
nand U2077 (N_2077,N_1995,N_1663);
or U2078 (N_2078,N_1967,N_1362);
nand U2079 (N_2079,N_1453,N_1720);
nand U2080 (N_2080,N_1873,In_1108);
nor U2081 (N_2081,N_1406,N_104);
or U2082 (N_2082,N_1832,N_1950);
nand U2083 (N_2083,N_1852,In_2897);
or U2084 (N_2084,N_1321,N_1384);
and U2085 (N_2085,N_1502,N_1578);
and U2086 (N_2086,N_1440,N_1830);
xnor U2087 (N_2087,N_1652,N_837);
nor U2088 (N_2088,N_1211,N_1046);
and U2089 (N_2089,N_1460,N_1655);
and U2090 (N_2090,N_1927,In_1336);
xor U2091 (N_2091,N_1711,N_1854);
nor U2092 (N_2092,N_886,In_2906);
xor U2093 (N_2093,N_1746,In_268);
xnor U2094 (N_2094,N_1335,N_1305);
and U2095 (N_2095,N_1125,N_1519);
and U2096 (N_2096,N_933,N_1866);
or U2097 (N_2097,In_2753,N_1771);
nand U2098 (N_2098,In_1815,N_1933);
nor U2099 (N_2099,N_149,N_1622);
or U2100 (N_2100,In_882,N_1518);
and U2101 (N_2101,In_730,In_1858);
and U2102 (N_2102,N_1312,N_301);
xnor U2103 (N_2103,N_1461,N_1318);
nor U2104 (N_2104,N_1935,N_1222);
nor U2105 (N_2105,In_2993,N_1906);
and U2106 (N_2106,In_2784,N_1385);
or U2107 (N_2107,N_1653,N_767);
or U2108 (N_2108,N_782,N_1025);
xor U2109 (N_2109,In_2565,N_543);
nor U2110 (N_2110,N_1769,N_1230);
or U2111 (N_2111,N_1012,N_1815);
nand U2112 (N_2112,N_898,N_1683);
nand U2113 (N_2113,In_606,In_1058);
nand U2114 (N_2114,In_45,In_559);
xnor U2115 (N_2115,In_1509,N_1982);
nand U2116 (N_2116,N_1417,N_280);
xor U2117 (N_2117,N_538,In_1493);
nor U2118 (N_2118,N_1763,N_950);
and U2119 (N_2119,N_1800,N_1266);
xor U2120 (N_2120,N_1923,N_1718);
or U2121 (N_2121,N_1823,In_339);
xor U2122 (N_2122,In_790,N_1674);
or U2123 (N_2123,N_845,In_2942);
nand U2124 (N_2124,N_1537,In_1385);
xor U2125 (N_2125,In_1966,In_1834);
or U2126 (N_2126,N_1201,N_1609);
or U2127 (N_2127,N_1892,N_140);
and U2128 (N_2128,N_1748,N_1514);
or U2129 (N_2129,N_1287,N_252);
or U2130 (N_2130,N_1474,In_105);
xor U2131 (N_2131,N_1296,In_1009);
nand U2132 (N_2132,In_840,N_627);
xor U2133 (N_2133,N_771,N_1677);
nand U2134 (N_2134,N_1856,N_1900);
and U2135 (N_2135,In_1997,N_1687);
or U2136 (N_2136,N_695,N_1281);
nand U2137 (N_2137,N_1671,N_1898);
nor U2138 (N_2138,N_1951,In_159);
nand U2139 (N_2139,N_463,N_1288);
nor U2140 (N_2140,N_1861,N_1972);
and U2141 (N_2141,N_689,N_1495);
nand U2142 (N_2142,N_1915,N_1458);
nor U2143 (N_2143,N_1952,N_1742);
or U2144 (N_2144,In_303,N_1510);
xnor U2145 (N_2145,N_1735,N_1801);
xor U2146 (N_2146,N_401,N_1928);
xnor U2147 (N_2147,N_340,N_1286);
or U2148 (N_2148,N_1916,In_1793);
and U2149 (N_2149,In_2671,N_1743);
and U2150 (N_2150,N_1620,N_940);
nand U2151 (N_2151,N_1804,N_945);
or U2152 (N_2152,N_1293,N_1930);
and U2153 (N_2153,N_1469,In_2996);
or U2154 (N_2154,N_1055,N_1548);
nand U2155 (N_2155,N_1979,N_1047);
xor U2156 (N_2156,N_1940,N_405);
and U2157 (N_2157,N_954,N_1934);
xnor U2158 (N_2158,N_1942,N_1196);
nor U2159 (N_2159,N_1809,N_1323);
xor U2160 (N_2160,N_996,In_1536);
nand U2161 (N_2161,N_1949,In_930);
and U2162 (N_2162,N_1343,N_1980);
nand U2163 (N_2163,N_1848,N_1500);
and U2164 (N_2164,N_1470,N_1110);
xor U2165 (N_2165,N_209,N_1650);
nor U2166 (N_2166,N_1740,N_1945);
or U2167 (N_2167,N_583,N_1206);
or U2168 (N_2168,N_1192,N_1719);
xor U2169 (N_2169,N_1831,N_1621);
xor U2170 (N_2170,N_1531,N_1709);
and U2171 (N_2171,In_1612,N_1868);
and U2172 (N_2172,N_1013,N_1855);
xor U2173 (N_2173,In_910,N_874);
xnor U2174 (N_2174,In_2570,In_2946);
or U2175 (N_2175,N_847,N_1747);
or U2176 (N_2176,N_1726,N_789);
and U2177 (N_2177,N_1309,N_876);
or U2178 (N_2178,N_1896,In_1888);
xnor U2179 (N_2179,N_1444,N_1782);
xor U2180 (N_2180,In_147,N_1985);
and U2181 (N_2181,N_1697,In_2955);
nand U2182 (N_2182,N_555,N_1941);
or U2183 (N_2183,N_1597,N_1113);
nand U2184 (N_2184,N_404,In_1095);
or U2185 (N_2185,N_1818,In_258);
and U2186 (N_2186,N_1634,N_1372);
and U2187 (N_2187,N_1890,N_796);
and U2188 (N_2188,In_343,N_912);
nand U2189 (N_2189,N_440,N_1996);
and U2190 (N_2190,In_1594,In_824);
nand U2191 (N_2191,N_1710,N_1889);
nor U2192 (N_2192,In_1698,N_256);
xnor U2193 (N_2193,In_2598,In_98);
and U2194 (N_2194,N_1907,N_1882);
or U2195 (N_2195,N_1562,In_2037);
or U2196 (N_2196,N_1728,N_1696);
nor U2197 (N_2197,In_2232,N_1657);
nor U2198 (N_2198,N_864,In_2397);
xnor U2199 (N_2199,N_1339,N_1843);
or U2200 (N_2200,In_1678,N_1358);
nand U2201 (N_2201,N_1783,N_2158);
xor U2202 (N_2202,N_2058,N_494);
or U2203 (N_2203,In_1746,In_1996);
nand U2204 (N_2204,In_1968,In_1056);
or U2205 (N_2205,N_1407,N_971);
xnor U2206 (N_2206,N_1501,N_2167);
or U2207 (N_2207,N_1765,In_729);
nand U2208 (N_2208,N_682,N_1242);
xnor U2209 (N_2209,N_1447,N_1912);
and U2210 (N_2210,N_1629,N_1186);
or U2211 (N_2211,N_2060,N_2025);
nand U2212 (N_2212,N_2186,N_1704);
nand U2213 (N_2213,In_275,N_1624);
or U2214 (N_2214,In_1211,In_1467);
and U2215 (N_2215,N_2181,N_1773);
xnor U2216 (N_2216,N_1820,N_1833);
xor U2217 (N_2217,N_629,N_1761);
nand U2218 (N_2218,In_2667,N_1130);
xor U2219 (N_2219,N_1439,N_1512);
and U2220 (N_2220,N_1229,N_1484);
and U2221 (N_2221,In_2198,N_1865);
nor U2222 (N_2222,N_1961,N_1938);
nand U2223 (N_2223,N_1990,N_1604);
nor U2224 (N_2224,N_277,N_1475);
xor U2225 (N_2225,N_1822,N_1842);
xor U2226 (N_2226,In_1758,N_1922);
or U2227 (N_2227,In_2452,N_1902);
or U2228 (N_2228,In_784,In_1933);
nand U2229 (N_2229,In_83,N_2185);
or U2230 (N_2230,N_1946,In_2668);
or U2231 (N_2231,N_1716,N_2106);
nand U2232 (N_2232,N_1897,N_1965);
nor U2233 (N_2233,N_2049,N_1577);
nor U2234 (N_2234,N_2030,N_639);
and U2235 (N_2235,N_2097,N_1886);
or U2236 (N_2236,In_1520,In_1068);
nor U2237 (N_2237,N_1805,N_1811);
xnor U2238 (N_2238,N_1552,In_1994);
xor U2239 (N_2239,N_1333,N_2110);
nor U2240 (N_2240,N_2055,N_1420);
xor U2241 (N_2241,N_2059,N_2015);
nand U2242 (N_2242,N_932,In_2847);
nand U2243 (N_2243,N_1633,In_750);
and U2244 (N_2244,N_1513,N_1775);
or U2245 (N_2245,N_902,N_1251);
or U2246 (N_2246,N_2048,N_2169);
nand U2247 (N_2247,N_2117,N_2040);
or U2248 (N_2248,N_1091,In_1152);
nor U2249 (N_2249,N_861,N_1948);
nand U2250 (N_2250,N_2126,N_1161);
nand U2251 (N_2251,In_747,N_1377);
nand U2252 (N_2252,N_2197,N_2011);
nor U2253 (N_2253,N_1788,In_2841);
and U2254 (N_2254,N_1300,N_1378);
xnor U2255 (N_2255,N_2033,N_1691);
nor U2256 (N_2256,N_2184,N_1977);
and U2257 (N_2257,N_1846,N_794);
nand U2258 (N_2258,N_1441,N_1290);
nor U2259 (N_2259,N_1860,N_1858);
and U2260 (N_2260,N_1062,N_1776);
nand U2261 (N_2261,N_1423,N_2115);
xnor U2262 (N_2262,N_1069,N_2071);
or U2263 (N_2263,N_14,N_2037);
nand U2264 (N_2264,N_1739,N_1538);
xor U2265 (N_2265,N_1862,N_2136);
xnor U2266 (N_2266,N_2148,N_2176);
nor U2267 (N_2267,N_734,In_2735);
nand U2268 (N_2268,In_1753,N_1436);
nand U2269 (N_2269,In_752,N_2138);
or U2270 (N_2270,N_2026,N_1664);
nor U2271 (N_2271,N_1755,N_1708);
nor U2272 (N_2272,N_1827,N_2123);
and U2273 (N_2273,N_2020,N_1616);
and U2274 (N_2274,N_2160,N_1825);
xnor U2275 (N_2275,N_1401,N_2111);
xor U2276 (N_2276,N_426,N_1590);
nor U2277 (N_2277,N_2008,N_1939);
or U2278 (N_2278,In_766,N_819);
nand U2279 (N_2279,N_2116,In_1643);
xnor U2280 (N_2280,N_1917,N_1901);
nor U2281 (N_2281,N_2014,N_1095);
and U2282 (N_2282,N_1779,In_420);
nand U2283 (N_2283,N_2162,N_672);
or U2284 (N_2284,N_1481,N_2113);
or U2285 (N_2285,N_1891,N_718);
nand U2286 (N_2286,N_607,N_2093);
xor U2287 (N_2287,N_1205,N_1403);
nand U2288 (N_2288,N_1541,N_2129);
xor U2289 (N_2289,N_1877,N_2121);
nand U2290 (N_2290,N_1573,N_2046);
and U2291 (N_2291,N_2021,N_1690);
nor U2292 (N_2292,In_683,N_2109);
nand U2293 (N_2293,N_1598,N_2177);
nand U2294 (N_2294,N_535,In_1328);
xor U2295 (N_2295,N_2170,N_1908);
xnor U2296 (N_2296,N_1736,N_153);
and U2297 (N_2297,N_710,N_2188);
or U2298 (N_2298,N_1348,In_1607);
nand U2299 (N_2299,N_1366,N_2174);
nor U2300 (N_2300,N_2163,N_1032);
and U2301 (N_2301,In_2691,N_1899);
nand U2302 (N_2302,N_1853,N_2127);
or U2303 (N_2303,N_1626,N_2198);
nand U2304 (N_2304,N_2178,N_1489);
and U2305 (N_2305,N_1591,N_1558);
nand U2306 (N_2306,In_2384,N_680);
and U2307 (N_2307,N_622,N_1936);
xor U2308 (N_2308,N_1670,N_1134);
or U2309 (N_2309,N_2057,In_1476);
or U2310 (N_2310,N_2050,N_1202);
nor U2311 (N_2311,N_517,N_1957);
xnor U2312 (N_2312,In_2798,N_56);
nor U2313 (N_2313,N_1885,N_1020);
nor U2314 (N_2314,N_1943,In_694);
xor U2315 (N_2315,N_1658,N_2006);
or U2316 (N_2316,N_1994,N_1074);
and U2317 (N_2317,In_286,N_1956);
or U2318 (N_2318,N_2104,In_2912);
and U2319 (N_2319,N_1602,In_169);
nand U2320 (N_2320,N_1794,N_1040);
and U2321 (N_2321,N_2054,N_2146);
nor U2322 (N_2322,N_434,N_1234);
nand U2323 (N_2323,N_2149,N_1480);
or U2324 (N_2324,N_260,N_2105);
xnor U2325 (N_2325,N_2141,N_2094);
and U2326 (N_2326,N_2195,N_1611);
nand U2327 (N_2327,N_2134,N_1798);
nor U2328 (N_2328,N_1579,In_2174);
and U2329 (N_2329,N_2073,N_1837);
xnor U2330 (N_2330,N_1894,N_1839);
or U2331 (N_2331,N_944,N_897);
or U2332 (N_2332,N_966,N_765);
xor U2333 (N_2333,N_1412,In_1557);
and U2334 (N_2334,N_1808,N_2112);
xor U2335 (N_2335,N_1871,N_2091);
nand U2336 (N_2336,In_1587,N_2157);
nand U2337 (N_2337,N_1126,N_1304);
and U2338 (N_2338,N_1103,N_571);
nand U2339 (N_2339,N_1588,N_2102);
nor U2340 (N_2340,N_1517,In_791);
or U2341 (N_2341,N_2150,N_2084);
or U2342 (N_2342,N_1918,N_2007);
and U2343 (N_2343,N_2077,N_530);
or U2344 (N_2344,N_1422,N_547);
nand U2345 (N_2345,N_1291,N_2063);
xor U2346 (N_2346,N_1806,N_1400);
and U2347 (N_2347,In_1005,N_2128);
or U2348 (N_2348,N_1813,N_532);
nor U2349 (N_2349,N_1669,In_1051);
and U2350 (N_2350,N_1324,N_2190);
nor U2351 (N_2351,N_1955,N_683);
nor U2352 (N_2352,In_378,N_2018);
nor U2353 (N_2353,N_1612,N_1493);
nor U2354 (N_2354,N_2156,N_1292);
xor U2355 (N_2355,N_2124,N_1947);
nor U2356 (N_2356,N_1411,N_1974);
nor U2357 (N_2357,In_955,N_1651);
xor U2358 (N_2358,N_2151,N_1580);
nand U2359 (N_2359,In_1359,N_488);
or U2360 (N_2360,N_2081,N_1625);
nor U2361 (N_2361,N_988,In_2230);
and U2362 (N_2362,N_1631,N_1983);
or U2363 (N_2363,In_2505,N_2032);
or U2364 (N_2364,N_1999,N_1225);
or U2365 (N_2365,N_1789,N_2119);
xor U2366 (N_2366,N_310,N_2165);
nand U2367 (N_2367,N_1857,In_2696);
and U2368 (N_2368,N_2088,N_1636);
xnor U2369 (N_2369,N_1503,N_1784);
xnor U2370 (N_2370,N_2196,In_921);
or U2371 (N_2371,N_550,N_758);
nand U2372 (N_2372,N_432,In_2263);
xnor U2373 (N_2373,N_1976,In_1226);
or U2374 (N_2374,In_110,N_1536);
nand U2375 (N_2375,N_1875,N_1642);
and U2376 (N_2376,In_561,In_1387);
or U2377 (N_2377,N_1486,N_1544);
or U2378 (N_2378,N_1926,N_1297);
or U2379 (N_2379,N_2016,N_1851);
and U2380 (N_2380,N_899,N_2024);
xor U2381 (N_2381,In_1873,N_1408);
nor U2382 (N_2382,In_1544,In_464);
or U2383 (N_2383,In_225,N_1920);
and U2384 (N_2384,N_1160,N_2182);
xor U2385 (N_2385,N_1478,N_2166);
nor U2386 (N_2386,N_766,N_1464);
nor U2387 (N_2387,In_2045,N_1641);
nand U2388 (N_2388,N_1559,In_2516);
and U2389 (N_2389,In_215,N_2133);
nor U2390 (N_2390,N_1365,N_1998);
nand U2391 (N_2391,N_1880,N_1821);
or U2392 (N_2392,In_768,N_1984);
and U2393 (N_2393,N_61,N_2183);
xnor U2394 (N_2394,N_2140,N_2155);
or U2395 (N_2395,In_1916,N_1803);
or U2396 (N_2396,N_1981,In_1381);
and U2397 (N_2397,N_1637,N_1864);
nor U2398 (N_2398,N_1978,N_2034);
and U2399 (N_2399,N_1971,In_1305);
nand U2400 (N_2400,N_1540,N_2363);
nor U2401 (N_2401,In_2375,N_1700);
nand U2402 (N_2402,N_2272,N_16);
xor U2403 (N_2403,N_2259,N_363);
and U2404 (N_2404,N_2053,N_244);
xnor U2405 (N_2405,N_2090,N_2137);
or U2406 (N_2406,N_2396,N_817);
nand U2407 (N_2407,N_2374,N_2179);
nand U2408 (N_2408,N_2070,N_2268);
nand U2409 (N_2409,N_271,N_2216);
nor U2410 (N_2410,N_949,N_424);
xor U2411 (N_2411,N_2282,N_2144);
and U2412 (N_2412,N_78,N_2202);
or U2413 (N_2413,N_1841,N_1656);
xor U2414 (N_2414,N_2293,In_422);
nand U2415 (N_2415,N_1695,N_2304);
or U2416 (N_2416,N_2079,N_2366);
nor U2417 (N_2417,N_2271,N_617);
and U2418 (N_2418,N_2211,N_2281);
nand U2419 (N_2419,N_2227,In_513);
or U2420 (N_2420,N_1828,N_2107);
and U2421 (N_2421,N_2336,N_2219);
nor U2422 (N_2422,N_2122,N_548);
nand U2423 (N_2423,N_2191,N_2239);
nand U2424 (N_2424,N_42,N_1929);
nand U2425 (N_2425,N_2321,N_637);
xnor U2426 (N_2426,N_2319,N_2237);
nor U2427 (N_2427,N_1419,N_704);
nor U2428 (N_2428,N_1648,In_814);
nand U2429 (N_2429,N_2047,N_2382);
nor U2430 (N_2430,N_2348,N_1183);
xnor U2431 (N_2431,N_1353,In_969);
and U2432 (N_2432,N_2118,N_931);
nand U2433 (N_2433,N_2233,N_2353);
xnor U2434 (N_2434,N_1428,N_2279);
and U2435 (N_2435,N_2242,N_2296);
nand U2436 (N_2436,N_1053,N_2043);
nor U2437 (N_2437,N_1758,N_2042);
xnor U2438 (N_2438,N_2315,N_1553);
xnor U2439 (N_2439,In_599,N_2012);
xor U2440 (N_2440,N_1909,N_1431);
and U2441 (N_2441,In_84,N_1793);
nand U2442 (N_2442,N_2300,N_2347);
xor U2443 (N_2443,N_623,N_2052);
xor U2444 (N_2444,N_802,N_2385);
nand U2445 (N_2445,N_2292,In_2896);
and U2446 (N_2446,N_2225,In_1094);
nor U2447 (N_2447,N_1812,N_2354);
and U2448 (N_2448,N_1570,In_2972);
nand U2449 (N_2449,N_2082,N_2171);
or U2450 (N_2450,N_1603,N_2028);
or U2451 (N_2451,N_2313,N_2301);
xor U2452 (N_2452,N_1239,N_2311);
nor U2453 (N_2453,N_670,N_2383);
and U2454 (N_2454,N_2263,N_2332);
xor U2455 (N_2455,N_2051,N_2373);
nor U2456 (N_2456,In_113,N_816);
nor U2457 (N_2457,In_1,In_2300);
and U2458 (N_2458,In_2453,N_2131);
or U2459 (N_2459,N_2253,N_2302);
and U2460 (N_2460,N_1585,N_1546);
or U2461 (N_2461,N_1963,N_2255);
nor U2462 (N_2462,In_763,N_2343);
xor U2463 (N_2463,N_1960,N_1416);
or U2464 (N_2464,N_2265,N_1660);
and U2465 (N_2465,N_2261,N_1058);
and U2466 (N_2466,N_2305,N_2205);
xnor U2467 (N_2467,In_952,N_1188);
xnor U2468 (N_2468,N_2377,N_2080);
nand U2469 (N_2469,In_2429,In_31);
nor U2470 (N_2470,N_739,N_697);
and U2471 (N_2471,N_776,N_1315);
xor U2472 (N_2472,N_2287,N_1850);
xor U2473 (N_2473,N_2023,N_407);
xnor U2474 (N_2474,N_2273,N_1757);
nor U2475 (N_2475,N_1816,N_1031);
nand U2476 (N_2476,N_1991,N_589);
and U2477 (N_2477,N_2004,N_2266);
xnor U2478 (N_2478,N_1893,N_2284);
and U2479 (N_2479,In_1370,N_2114);
nand U2480 (N_2480,In_2926,N_2194);
xor U2481 (N_2481,In_892,N_1688);
nand U2482 (N_2482,In_2885,N_2230);
nand U2483 (N_2483,N_2218,N_2340);
xnor U2484 (N_2484,In_1616,N_2379);
nor U2485 (N_2485,N_2326,N_1081);
or U2486 (N_2486,N_2365,N_2002);
or U2487 (N_2487,N_2000,N_2089);
nand U2488 (N_2488,N_2217,N_1754);
xnor U2489 (N_2489,In_818,N_2370);
xor U2490 (N_2490,N_2278,N_126);
and U2491 (N_2491,N_2378,N_1665);
nor U2492 (N_2492,N_2041,N_2264);
or U2493 (N_2493,In_1730,In_2266);
or U2494 (N_2494,N_1921,N_1351);
nand U2495 (N_2495,In_1465,N_1904);
xnor U2496 (N_2496,N_1944,N_2339);
nand U2497 (N_2497,N_788,N_2371);
xor U2498 (N_2498,N_1265,N_1975);
xnor U2499 (N_2499,N_2223,N_1308);
xnor U2500 (N_2500,N_2294,N_382);
nand U2501 (N_2501,N_1874,N_1762);
nand U2502 (N_2502,N_2251,N_2369);
or U2503 (N_2503,In_1822,N_2044);
or U2504 (N_2504,N_2350,N_2276);
or U2505 (N_2505,N_2323,N_93);
nand U2506 (N_2506,In_2693,N_2390);
nor U2507 (N_2507,N_2360,N_2221);
xor U2508 (N_2508,In_2063,N_1838);
nor U2509 (N_2509,In_1219,N_2289);
or U2510 (N_2510,N_1644,N_1574);
xnor U2511 (N_2511,N_1872,N_2260);
nand U2512 (N_2512,N_2153,N_2100);
xor U2513 (N_2513,N_2389,In_2474);
or U2514 (N_2514,N_1138,N_1421);
or U2515 (N_2515,N_2243,N_2240);
xor U2516 (N_2516,N_2215,In_2299);
xnor U2517 (N_2517,N_1888,N_2393);
nand U2518 (N_2518,N_1859,N_2291);
or U2519 (N_2519,N_2331,N_1402);
nand U2520 (N_2520,N_2388,In_2211);
and U2521 (N_2521,N_286,N_2035);
xor U2522 (N_2522,N_2038,N_805);
nand U2523 (N_2523,N_10,N_1237);
and U2524 (N_2524,N_2290,N_2248);
or U2525 (N_2525,N_2208,N_2065);
nor U2526 (N_2526,N_1106,N_1448);
nand U2527 (N_2527,N_1903,N_374);
or U2528 (N_2528,N_1140,In_1689);
nor U2529 (N_2529,N_1592,N_2309);
and U2530 (N_2530,N_2220,N_2394);
and U2531 (N_2531,N_1768,N_1722);
nor U2532 (N_2532,N_1194,N_1112);
nor U2533 (N_2533,N_2245,In_1221);
nor U2534 (N_2534,N_1556,N_2192);
xor U2535 (N_2535,N_2335,N_2384);
and U2536 (N_2536,N_2173,N_741);
nand U2537 (N_2537,N_1701,In_868);
or U2538 (N_2538,N_2013,N_2397);
or U2539 (N_2539,In_1398,N_2325);
and U2540 (N_2540,N_2187,N_2213);
or U2541 (N_2541,N_1639,N_2303);
xnor U2542 (N_2542,In_2215,N_1443);
and U2543 (N_2543,N_1876,In_2719);
nor U2544 (N_2544,N_2346,N_866);
nor U2545 (N_2545,N_2236,N_1778);
xor U2546 (N_2546,N_2045,N_2380);
and U2547 (N_2547,N_172,N_1969);
xor U2548 (N_2548,N_2099,N_2022);
nand U2549 (N_2549,N_2375,N_2238);
nor U2550 (N_2550,N_2145,N_416);
xnor U2551 (N_2551,N_2154,N_1185);
nand U2552 (N_2552,N_2334,N_2103);
and U2553 (N_2553,N_2308,N_1274);
or U2554 (N_2554,N_1432,N_2241);
and U2555 (N_2555,In_990,N_2372);
xor U2556 (N_2556,N_1618,N_2076);
and U2557 (N_2557,N_2246,N_2256);
xnor U2558 (N_2558,In_2191,N_2226);
or U2559 (N_2559,N_2395,N_1693);
or U2560 (N_2560,In_2404,N_1347);
or U2561 (N_2561,N_2086,N_1729);
nand U2562 (N_2562,N_1615,N_2142);
nand U2563 (N_2563,N_611,N_2322);
nor U2564 (N_2564,N_2201,N_2306);
and U2565 (N_2565,In_732,N_1931);
or U2566 (N_2566,N_2207,N_192);
nand U2567 (N_2567,N_2376,In_627);
xnor U2568 (N_2568,N_1127,N_2288);
xor U2569 (N_2569,N_2074,N_2039);
and U2570 (N_2570,N_332,N_2078);
or U2571 (N_2571,In_1459,N_2338);
and U2572 (N_2572,In_1842,N_2244);
and U2573 (N_2573,N_2027,N_1599);
nor U2574 (N_2574,N_762,N_1987);
or U2575 (N_2575,N_2399,N_2139);
xor U2576 (N_2576,N_1162,N_2232);
xor U2577 (N_2577,In_914,N_2199);
nor U2578 (N_2578,N_1937,N_1359);
nor U2579 (N_2579,N_2337,N_2361);
nand U2580 (N_2580,N_2387,N_2168);
and U2581 (N_2581,N_1261,N_1913);
or U2582 (N_2582,In_2924,N_651);
or U2583 (N_2583,N_2392,N_2095);
nor U2584 (N_2584,N_2064,N_2307);
nor U2585 (N_2585,N_2327,In_685);
nand U2586 (N_2586,N_1869,N_2355);
and U2587 (N_2587,N_1780,N_1632);
or U2588 (N_2588,N_2200,N_2083);
and U2589 (N_2589,N_2019,N_2224);
or U2590 (N_2590,N_1643,N_2258);
or U2591 (N_2591,N_1129,N_1360);
xor U2592 (N_2592,N_917,N_2061);
nand U2593 (N_2593,In_1294,N_2029);
nand U2594 (N_2594,N_2359,In_2206);
and U2595 (N_2595,N_1986,N_1702);
and U2596 (N_2596,In_2844,N_1457);
nand U2597 (N_2597,N_2231,N_2228);
or U2598 (N_2598,N_474,N_990);
nor U2599 (N_2599,N_2252,N_2344);
and U2600 (N_2600,N_2445,N_2555);
nand U2601 (N_2601,N_997,N_2212);
nand U2602 (N_2602,N_2562,N_1139);
nand U2603 (N_2603,N_2010,N_2521);
or U2604 (N_2604,N_1914,N_2534);
xnor U2605 (N_2605,N_2443,N_2330);
xnor U2606 (N_2606,N_2554,N_1870);
xor U2607 (N_2607,N_2092,N_1563);
nor U2608 (N_2608,N_2556,N_2531);
nand U2609 (N_2609,N_2062,N_2275);
or U2610 (N_2610,N_2509,N_2430);
nand U2611 (N_2611,N_2193,N_2535);
nor U2612 (N_2612,N_810,N_2532);
and U2613 (N_2613,N_2257,N_1210);
nand U2614 (N_2614,N_2479,N_2143);
xnor U2615 (N_2615,N_2437,In_1952);
nor U2616 (N_2616,In_1374,N_2596);
and U2617 (N_2617,N_2530,N_2180);
nor U2618 (N_2618,N_2574,In_2727);
or U2619 (N_2619,N_2464,N_2503);
xor U2620 (N_2620,N_2585,N_2249);
or U2621 (N_2621,N_2565,N_2410);
nand U2622 (N_2622,N_2564,N_2405);
or U2623 (N_2623,N_542,N_2458);
xor U2624 (N_2624,N_2506,N_2483);
nor U2625 (N_2625,N_2481,N_2547);
nand U2626 (N_2626,N_2130,N_2203);
nor U2627 (N_2627,N_2001,N_2423);
nand U2628 (N_2628,N_2072,N_2206);
xnor U2629 (N_2629,N_2567,N_646);
nand U2630 (N_2630,N_2277,N_2132);
and U2631 (N_2631,N_2222,N_2229);
xor U2632 (N_2632,N_647,N_2578);
and U2633 (N_2633,N_2404,N_2560);
and U2634 (N_2634,N_2283,N_2175);
nor U2635 (N_2635,N_2408,N_2468);
and U2636 (N_2636,N_2362,N_2594);
and U2637 (N_2637,N_1817,In_733);
or U2638 (N_2638,N_2514,N_2501);
nor U2639 (N_2639,N_2269,N_2511);
nor U2640 (N_2640,N_863,N_1887);
or U2641 (N_2641,In_2776,In_433);
nand U2642 (N_2642,N_2096,N_2566);
and U2643 (N_2643,N_2570,N_1547);
nand U2644 (N_2644,N_1661,N_2391);
or U2645 (N_2645,N_2583,N_1628);
or U2646 (N_2646,N_2415,N_2235);
nand U2647 (N_2647,N_2444,N_2407);
xnor U2648 (N_2648,N_1767,N_2416);
or U2649 (N_2649,N_2490,N_2411);
nor U2650 (N_2650,N_2418,N_2398);
nand U2651 (N_2651,N_2358,N_2247);
nand U2652 (N_2652,N_2270,N_2250);
or U2653 (N_2653,N_1919,N_2066);
nor U2654 (N_2654,In_2376,N_2469);
xnor U2655 (N_2655,N_2285,N_2572);
nor U2656 (N_2656,N_2496,N_2493);
and U2657 (N_2657,N_2492,In_2028);
or U2658 (N_2658,N_916,N_2455);
xor U2659 (N_2659,N_2502,N_2381);
xnor U2660 (N_2660,N_2526,N_2428);
nand U2661 (N_2661,N_1668,In_1728);
and U2662 (N_2662,N_2573,N_2352);
and U2663 (N_2663,N_2459,N_2403);
nand U2664 (N_2664,N_2460,N_1845);
nor U2665 (N_2665,N_1863,N_2009);
nor U2666 (N_2666,In_913,N_2429);
and U2667 (N_2667,N_1849,N_2274);
or U2668 (N_2668,N_2449,N_2262);
xor U2669 (N_2669,N_2056,In_2195);
and U2670 (N_2670,N_2210,N_2448);
or U2671 (N_2671,N_2489,N_2523);
or U2672 (N_2672,N_2351,N_2364);
and U2673 (N_2673,N_2579,N_2474);
nand U2674 (N_2674,N_2482,N_2172);
xnor U2675 (N_2675,N_2451,N_2552);
and U2676 (N_2676,N_2558,In_1126);
and U2677 (N_2677,N_2505,In_1083);
and U2678 (N_2678,N_1008,N_1607);
nor U2679 (N_2679,N_2582,N_2568);
nand U2680 (N_2680,N_2541,N_2368);
or U2681 (N_2681,N_857,N_2591);
or U2682 (N_2682,N_1844,N_2527);
xnor U2683 (N_2683,N_421,In_267);
and U2684 (N_2684,N_2546,N_2462);
nand U2685 (N_2685,N_2441,N_2345);
nor U2686 (N_2686,In_1050,N_2414);
nand U2687 (N_2687,N_2328,N_1749);
and U2688 (N_2688,N_2597,N_1895);
xnor U2689 (N_2689,N_2475,N_2500);
nor U2690 (N_2690,N_2473,N_2520);
nand U2691 (N_2691,N_2067,N_2525);
xnor U2692 (N_2692,N_2539,N_2519);
or U2693 (N_2693,N_2401,N_769);
nor U2694 (N_2694,N_2320,N_2152);
and U2695 (N_2695,N_2497,N_1959);
nand U2696 (N_2696,In_1708,N_1521);
nand U2697 (N_2697,N_1836,N_2518);
nor U2698 (N_2698,N_1781,N_2433);
xnor U2699 (N_2699,N_2280,In_1859);
nor U2700 (N_2700,N_2588,N_2386);
nor U2701 (N_2701,N_1388,N_2420);
nand U2702 (N_2702,N_601,N_2517);
nor U2703 (N_2703,N_1699,N_2478);
nand U2704 (N_2704,N_2593,N_2333);
nor U2705 (N_2705,N_1752,N_2467);
and U2706 (N_2706,N_2314,N_1061);
nor U2707 (N_2707,N_2159,N_2349);
xor U2708 (N_2708,N_2412,N_2559);
and U2709 (N_2709,N_2550,N_2341);
nor U2710 (N_2710,N_2569,N_2499);
nor U2711 (N_2711,N_2453,N_2135);
nand U2712 (N_2712,N_2254,N_2424);
or U2713 (N_2713,N_2164,N_2427);
xor U2714 (N_2714,N_2598,N_2356);
nor U2715 (N_2715,N_1966,N_2480);
xor U2716 (N_2716,N_2298,N_2161);
nand U2717 (N_2717,N_2471,N_2486);
or U2718 (N_2718,N_2297,N_2592);
or U2719 (N_2719,N_2295,N_1395);
and U2720 (N_2720,N_2540,N_1459);
xor U2721 (N_2721,N_2576,N_2317);
or U2722 (N_2722,N_2204,N_677);
xnor U2723 (N_2723,N_2507,N_1410);
xor U2724 (N_2724,In_1409,In_2984);
or U2725 (N_2725,N_2584,N_839);
xor U2726 (N_2726,N_2108,N_2465);
nand U2727 (N_2727,N_2561,N_1807);
or U2728 (N_2728,N_1515,N_2545);
nor U2729 (N_2729,N_1516,N_2442);
or U2730 (N_2730,N_2438,N_2557);
nor U2731 (N_2731,N_2495,N_2512);
or U2732 (N_2732,N_2447,N_2456);
xnor U2733 (N_2733,In_2091,N_2536);
nand U2734 (N_2734,N_2528,N_2425);
and U2735 (N_2735,N_2426,N_2577);
nor U2736 (N_2736,N_1097,N_2068);
nand U2737 (N_2737,N_2586,N_979);
or U2738 (N_2738,N_2085,N_2440);
nor U2739 (N_2739,N_1840,N_2413);
nor U2740 (N_2740,N_2087,N_1954);
xnor U2741 (N_2741,N_2548,N_2533);
xor U2742 (N_2742,N_1992,In_2545);
nor U2743 (N_2743,N_660,N_2357);
or U2744 (N_2744,N_2452,N_2421);
xnor U2745 (N_2745,In_960,N_1925);
and U2746 (N_2746,N_2147,In_2041);
and U2747 (N_2747,N_2120,N_2436);
nand U2748 (N_2748,N_2286,N_2036);
or U2749 (N_2749,N_2101,N_1717);
nor U2750 (N_2750,N_2402,N_2522);
and U2751 (N_2751,N_2516,N_2422);
nor U2752 (N_2752,N_2457,N_2267);
xor U2753 (N_2753,N_2214,N_2510);
nand U2754 (N_2754,N_2069,N_2537);
or U2755 (N_2755,N_2553,N_315);
nor U2756 (N_2756,N_2316,N_2590);
nand U2757 (N_2757,N_2406,N_2551);
nand U2758 (N_2758,N_2312,N_2544);
nor U2759 (N_2759,N_2342,N_2450);
or U2760 (N_2760,N_2581,N_2542);
nand U2761 (N_2761,N_2329,N_2589);
nand U2762 (N_2762,N_2461,N_1048);
nor U2763 (N_2763,N_2435,N_2538);
nand U2764 (N_2764,N_815,N_2487);
nor U2765 (N_2765,N_2367,N_2324);
nand U2766 (N_2766,N_2466,N_2234);
nor U2767 (N_2767,N_2599,N_669);
nand U2768 (N_2768,N_2549,N_1879);
and U2769 (N_2769,N_2299,N_2431);
or U2770 (N_2770,N_2580,N_2515);
nand U2771 (N_2771,In_1760,N_2494);
nand U2772 (N_2772,N_2470,N_1452);
nand U2773 (N_2773,In_1165,N_2595);
nor U2774 (N_2774,N_2031,In_78);
or U2775 (N_2775,N_2563,N_2472);
and U2776 (N_2776,N_2571,N_2543);
xor U2777 (N_2777,N_2318,N_1085);
or U2778 (N_2778,N_1617,N_2463);
nor U2779 (N_2779,In_2785,N_1199);
nor U2780 (N_2780,N_1796,N_2513);
or U2781 (N_2781,N_2005,N_2524);
nor U2782 (N_2782,N_2446,N_2075);
and U2783 (N_2783,N_2504,N_1810);
and U2784 (N_2784,N_2529,N_2400);
nor U2785 (N_2785,N_2209,N_2125);
xor U2786 (N_2786,N_2477,N_2432);
nand U2787 (N_2787,N_2409,N_2488);
nor U2788 (N_2788,N_2587,N_2498);
xnor U2789 (N_2789,N_2419,N_2098);
and U2790 (N_2790,N_2189,N_1988);
nand U2791 (N_2791,N_953,N_2003);
and U2792 (N_2792,N_2508,N_2017);
and U2793 (N_2793,In_2172,N_2417);
xnor U2794 (N_2794,N_2484,N_2491);
and U2795 (N_2795,N_2454,N_2310);
and U2796 (N_2796,N_2476,In_1182);
nand U2797 (N_2797,N_2439,N_2575);
xor U2798 (N_2798,N_2485,In_2707);
nor U2799 (N_2799,N_2434,N_92);
and U2800 (N_2800,N_2605,N_2727);
nor U2801 (N_2801,N_2721,N_2682);
xnor U2802 (N_2802,N_2645,N_2704);
or U2803 (N_2803,N_2603,N_2644);
xor U2804 (N_2804,N_2623,N_2696);
nor U2805 (N_2805,N_2638,N_2674);
nand U2806 (N_2806,N_2720,N_2730);
nand U2807 (N_2807,N_2765,N_2627);
and U2808 (N_2808,N_2745,N_2626);
and U2809 (N_2809,N_2617,N_2635);
xor U2810 (N_2810,N_2772,N_2607);
or U2811 (N_2811,N_2742,N_2622);
or U2812 (N_2812,N_2641,N_2652);
nor U2813 (N_2813,N_2666,N_2744);
and U2814 (N_2814,N_2633,N_2631);
and U2815 (N_2815,N_2698,N_2783);
and U2816 (N_2816,N_2781,N_2695);
nor U2817 (N_2817,N_2612,N_2752);
xor U2818 (N_2818,N_2675,N_2618);
nor U2819 (N_2819,N_2750,N_2782);
nor U2820 (N_2820,N_2705,N_2743);
xnor U2821 (N_2821,N_2667,N_2653);
and U2822 (N_2822,N_2699,N_2639);
and U2823 (N_2823,N_2620,N_2774);
nand U2824 (N_2824,N_2646,N_2606);
nand U2825 (N_2825,N_2658,N_2724);
and U2826 (N_2826,N_2685,N_2797);
nand U2827 (N_2827,N_2679,N_2648);
nand U2828 (N_2828,N_2647,N_2790);
nand U2829 (N_2829,N_2740,N_2616);
xnor U2830 (N_2830,N_2661,N_2792);
or U2831 (N_2831,N_2747,N_2655);
or U2832 (N_2832,N_2650,N_2628);
or U2833 (N_2833,N_2716,N_2656);
nor U2834 (N_2834,N_2643,N_2692);
nand U2835 (N_2835,N_2689,N_2799);
nor U2836 (N_2836,N_2725,N_2755);
or U2837 (N_2837,N_2654,N_2634);
nor U2838 (N_2838,N_2714,N_2708);
nor U2839 (N_2839,N_2604,N_2768);
nor U2840 (N_2840,N_2673,N_2707);
and U2841 (N_2841,N_2751,N_2660);
or U2842 (N_2842,N_2736,N_2702);
nand U2843 (N_2843,N_2624,N_2786);
nand U2844 (N_2844,N_2659,N_2798);
xor U2845 (N_2845,N_2629,N_2757);
or U2846 (N_2846,N_2741,N_2601);
or U2847 (N_2847,N_2722,N_2737);
and U2848 (N_2848,N_2614,N_2684);
and U2849 (N_2849,N_2677,N_2780);
and U2850 (N_2850,N_2651,N_2632);
or U2851 (N_2851,N_2715,N_2610);
xor U2852 (N_2852,N_2678,N_2733);
nand U2853 (N_2853,N_2795,N_2630);
xor U2854 (N_2854,N_2680,N_2686);
nor U2855 (N_2855,N_2770,N_2749);
nor U2856 (N_2856,N_2760,N_2717);
or U2857 (N_2857,N_2636,N_2611);
nor U2858 (N_2858,N_2694,N_2762);
or U2859 (N_2859,N_2640,N_2602);
nor U2860 (N_2860,N_2642,N_2621);
nand U2861 (N_2861,N_2681,N_2787);
xnor U2862 (N_2862,N_2738,N_2663);
nor U2863 (N_2863,N_2687,N_2697);
and U2864 (N_2864,N_2665,N_2711);
nor U2865 (N_2865,N_2637,N_2764);
or U2866 (N_2866,N_2784,N_2701);
or U2867 (N_2867,N_2718,N_2615);
or U2868 (N_2868,N_2761,N_2734);
nor U2869 (N_2869,N_2777,N_2723);
xnor U2870 (N_2870,N_2671,N_2703);
nor U2871 (N_2871,N_2662,N_2769);
nor U2872 (N_2872,N_2785,N_2608);
nand U2873 (N_2873,N_2683,N_2773);
or U2874 (N_2874,N_2791,N_2710);
nand U2875 (N_2875,N_2657,N_2719);
nand U2876 (N_2876,N_2753,N_2691);
xnor U2877 (N_2877,N_2731,N_2771);
nand U2878 (N_2878,N_2759,N_2739);
and U2879 (N_2879,N_2778,N_2735);
nand U2880 (N_2880,N_2775,N_2609);
and U2881 (N_2881,N_2713,N_2709);
nand U2882 (N_2882,N_2712,N_2726);
nor U2883 (N_2883,N_2670,N_2788);
and U2884 (N_2884,N_2728,N_2796);
or U2885 (N_2885,N_2690,N_2668);
xor U2886 (N_2886,N_2688,N_2763);
xor U2887 (N_2887,N_2625,N_2732);
nand U2888 (N_2888,N_2729,N_2706);
nor U2889 (N_2889,N_2754,N_2779);
or U2890 (N_2890,N_2776,N_2766);
or U2891 (N_2891,N_2758,N_2793);
nor U2892 (N_2892,N_2672,N_2756);
or U2893 (N_2893,N_2619,N_2676);
xnor U2894 (N_2894,N_2746,N_2767);
nor U2895 (N_2895,N_2748,N_2700);
xnor U2896 (N_2896,N_2794,N_2600);
xor U2897 (N_2897,N_2693,N_2613);
or U2898 (N_2898,N_2669,N_2789);
xnor U2899 (N_2899,N_2649,N_2664);
nor U2900 (N_2900,N_2718,N_2689);
xor U2901 (N_2901,N_2703,N_2716);
and U2902 (N_2902,N_2723,N_2661);
and U2903 (N_2903,N_2605,N_2668);
nand U2904 (N_2904,N_2615,N_2653);
or U2905 (N_2905,N_2612,N_2771);
nor U2906 (N_2906,N_2774,N_2729);
nor U2907 (N_2907,N_2600,N_2629);
and U2908 (N_2908,N_2601,N_2762);
nand U2909 (N_2909,N_2782,N_2761);
nor U2910 (N_2910,N_2760,N_2761);
or U2911 (N_2911,N_2789,N_2790);
xnor U2912 (N_2912,N_2678,N_2766);
nand U2913 (N_2913,N_2656,N_2788);
or U2914 (N_2914,N_2615,N_2612);
xnor U2915 (N_2915,N_2771,N_2770);
xor U2916 (N_2916,N_2648,N_2607);
xor U2917 (N_2917,N_2679,N_2700);
nor U2918 (N_2918,N_2775,N_2778);
and U2919 (N_2919,N_2658,N_2691);
nand U2920 (N_2920,N_2715,N_2686);
nand U2921 (N_2921,N_2786,N_2698);
and U2922 (N_2922,N_2750,N_2739);
or U2923 (N_2923,N_2738,N_2696);
and U2924 (N_2924,N_2682,N_2722);
nor U2925 (N_2925,N_2791,N_2796);
nor U2926 (N_2926,N_2635,N_2783);
nor U2927 (N_2927,N_2746,N_2673);
and U2928 (N_2928,N_2681,N_2613);
nand U2929 (N_2929,N_2620,N_2637);
nand U2930 (N_2930,N_2789,N_2626);
or U2931 (N_2931,N_2620,N_2757);
or U2932 (N_2932,N_2788,N_2782);
nor U2933 (N_2933,N_2609,N_2787);
nor U2934 (N_2934,N_2717,N_2742);
or U2935 (N_2935,N_2601,N_2655);
xor U2936 (N_2936,N_2607,N_2793);
or U2937 (N_2937,N_2709,N_2706);
nand U2938 (N_2938,N_2667,N_2698);
or U2939 (N_2939,N_2651,N_2734);
nor U2940 (N_2940,N_2653,N_2787);
xnor U2941 (N_2941,N_2639,N_2683);
or U2942 (N_2942,N_2727,N_2632);
nor U2943 (N_2943,N_2679,N_2615);
nor U2944 (N_2944,N_2696,N_2790);
or U2945 (N_2945,N_2649,N_2669);
nand U2946 (N_2946,N_2739,N_2623);
nor U2947 (N_2947,N_2603,N_2642);
nor U2948 (N_2948,N_2601,N_2646);
nand U2949 (N_2949,N_2747,N_2674);
or U2950 (N_2950,N_2657,N_2771);
nand U2951 (N_2951,N_2640,N_2752);
and U2952 (N_2952,N_2696,N_2683);
and U2953 (N_2953,N_2748,N_2697);
nand U2954 (N_2954,N_2787,N_2638);
or U2955 (N_2955,N_2684,N_2739);
nand U2956 (N_2956,N_2649,N_2705);
nand U2957 (N_2957,N_2704,N_2724);
nor U2958 (N_2958,N_2689,N_2760);
or U2959 (N_2959,N_2724,N_2631);
and U2960 (N_2960,N_2789,N_2695);
nand U2961 (N_2961,N_2647,N_2693);
nand U2962 (N_2962,N_2602,N_2644);
nor U2963 (N_2963,N_2612,N_2623);
xnor U2964 (N_2964,N_2680,N_2752);
nand U2965 (N_2965,N_2798,N_2679);
nand U2966 (N_2966,N_2627,N_2754);
xor U2967 (N_2967,N_2793,N_2634);
and U2968 (N_2968,N_2730,N_2617);
xor U2969 (N_2969,N_2716,N_2782);
nand U2970 (N_2970,N_2701,N_2655);
and U2971 (N_2971,N_2677,N_2619);
nand U2972 (N_2972,N_2772,N_2755);
xnor U2973 (N_2973,N_2763,N_2656);
nor U2974 (N_2974,N_2705,N_2774);
nor U2975 (N_2975,N_2668,N_2609);
nor U2976 (N_2976,N_2680,N_2638);
nor U2977 (N_2977,N_2762,N_2708);
and U2978 (N_2978,N_2716,N_2772);
nor U2979 (N_2979,N_2777,N_2747);
and U2980 (N_2980,N_2653,N_2793);
xnor U2981 (N_2981,N_2603,N_2660);
nand U2982 (N_2982,N_2656,N_2705);
xor U2983 (N_2983,N_2698,N_2668);
nand U2984 (N_2984,N_2737,N_2676);
nor U2985 (N_2985,N_2796,N_2798);
xor U2986 (N_2986,N_2638,N_2773);
nor U2987 (N_2987,N_2652,N_2660);
or U2988 (N_2988,N_2787,N_2783);
nor U2989 (N_2989,N_2686,N_2641);
or U2990 (N_2990,N_2791,N_2688);
or U2991 (N_2991,N_2724,N_2634);
or U2992 (N_2992,N_2737,N_2760);
xor U2993 (N_2993,N_2671,N_2773);
and U2994 (N_2994,N_2753,N_2757);
nand U2995 (N_2995,N_2760,N_2695);
and U2996 (N_2996,N_2733,N_2729);
nand U2997 (N_2997,N_2666,N_2672);
nor U2998 (N_2998,N_2759,N_2624);
nor U2999 (N_2999,N_2758,N_2759);
xnor U3000 (N_3000,N_2958,N_2982);
nand U3001 (N_3001,N_2924,N_2996);
and U3002 (N_3002,N_2963,N_2940);
nor U3003 (N_3003,N_2992,N_2935);
nor U3004 (N_3004,N_2960,N_2879);
or U3005 (N_3005,N_2939,N_2878);
or U3006 (N_3006,N_2834,N_2814);
nand U3007 (N_3007,N_2829,N_2852);
nor U3008 (N_3008,N_2919,N_2951);
or U3009 (N_3009,N_2943,N_2946);
and U3010 (N_3010,N_2848,N_2941);
and U3011 (N_3011,N_2962,N_2923);
or U3012 (N_3012,N_2983,N_2858);
and U3013 (N_3013,N_2802,N_2945);
and U3014 (N_3014,N_2804,N_2977);
or U3015 (N_3015,N_2920,N_2808);
nand U3016 (N_3016,N_2965,N_2849);
or U3017 (N_3017,N_2926,N_2894);
or U3018 (N_3018,N_2971,N_2961);
and U3019 (N_3019,N_2856,N_2954);
xnor U3020 (N_3020,N_2861,N_2973);
xor U3021 (N_3021,N_2978,N_2869);
xor U3022 (N_3022,N_2981,N_2985);
or U3023 (N_3023,N_2832,N_2929);
or U3024 (N_3024,N_2831,N_2901);
xnor U3025 (N_3025,N_2807,N_2937);
nor U3026 (N_3026,N_2957,N_2905);
xnor U3027 (N_3027,N_2847,N_2893);
nand U3028 (N_3028,N_2842,N_2944);
nor U3029 (N_3029,N_2864,N_2956);
and U3030 (N_3030,N_2874,N_2866);
or U3031 (N_3031,N_2953,N_2865);
xnor U3032 (N_3032,N_2896,N_2863);
xor U3033 (N_3033,N_2969,N_2948);
nand U3034 (N_3034,N_2815,N_2855);
nor U3035 (N_3035,N_2952,N_2881);
or U3036 (N_3036,N_2833,N_2989);
xor U3037 (N_3037,N_2936,N_2843);
and U3038 (N_3038,N_2922,N_2892);
nand U3039 (N_3039,N_2931,N_2818);
xor U3040 (N_3040,N_2925,N_2942);
or U3041 (N_3041,N_2914,N_2980);
or U3042 (N_3042,N_2909,N_2912);
xnor U3043 (N_3043,N_2972,N_2876);
nor U3044 (N_3044,N_2964,N_2853);
or U3045 (N_3045,N_2838,N_2836);
nor U3046 (N_3046,N_2870,N_2900);
nand U3047 (N_3047,N_2993,N_2850);
and U3048 (N_3048,N_2970,N_2805);
and U3049 (N_3049,N_2888,N_2809);
or U3050 (N_3050,N_2932,N_2860);
xnor U3051 (N_3051,N_2800,N_2979);
nand U3052 (N_3052,N_2955,N_2872);
and U3053 (N_3053,N_2908,N_2950);
nand U3054 (N_3054,N_2810,N_2975);
xnor U3055 (N_3055,N_2806,N_2895);
or U3056 (N_3056,N_2835,N_2968);
or U3057 (N_3057,N_2873,N_2928);
xor U3058 (N_3058,N_2885,N_2917);
or U3059 (N_3059,N_2839,N_2986);
or U3060 (N_3060,N_2907,N_2841);
nand U3061 (N_3061,N_2903,N_2898);
or U3062 (N_3062,N_2817,N_2840);
xor U3063 (N_3063,N_2915,N_2974);
or U3064 (N_3064,N_2882,N_2813);
xor U3065 (N_3065,N_2811,N_2824);
nand U3066 (N_3066,N_2837,N_2823);
nor U3067 (N_3067,N_2845,N_2877);
nand U3068 (N_3068,N_2934,N_2987);
xor U3069 (N_3069,N_2868,N_2906);
nor U3070 (N_3070,N_2889,N_2820);
and U3071 (N_3071,N_2984,N_2854);
or U3072 (N_3072,N_2887,N_2918);
xor U3073 (N_3073,N_2844,N_2827);
nand U3074 (N_3074,N_2990,N_2812);
or U3075 (N_3075,N_2826,N_2947);
or U3076 (N_3076,N_2959,N_2891);
nor U3077 (N_3077,N_2988,N_2995);
nand U3078 (N_3078,N_2933,N_2949);
and U3079 (N_3079,N_2830,N_2902);
nand U3080 (N_3080,N_2857,N_2897);
xor U3081 (N_3081,N_2910,N_2999);
and U3082 (N_3082,N_2927,N_2938);
or U3083 (N_3083,N_2967,N_2913);
nand U3084 (N_3084,N_2880,N_2821);
nor U3085 (N_3085,N_2801,N_2871);
or U3086 (N_3086,N_2991,N_2930);
and U3087 (N_3087,N_2884,N_2846);
nor U3088 (N_3088,N_2828,N_2899);
nand U3089 (N_3089,N_2998,N_2822);
nand U3090 (N_3090,N_2883,N_2976);
nor U3091 (N_3091,N_2890,N_2875);
xor U3092 (N_3092,N_2911,N_2916);
nand U3093 (N_3093,N_2904,N_2859);
nor U3094 (N_3094,N_2867,N_2851);
or U3095 (N_3095,N_2862,N_2921);
xor U3096 (N_3096,N_2825,N_2997);
nand U3097 (N_3097,N_2886,N_2816);
nand U3098 (N_3098,N_2803,N_2994);
xor U3099 (N_3099,N_2819,N_2966);
xor U3100 (N_3100,N_2938,N_2910);
and U3101 (N_3101,N_2928,N_2857);
nand U3102 (N_3102,N_2907,N_2868);
nand U3103 (N_3103,N_2942,N_2853);
and U3104 (N_3104,N_2921,N_2930);
xnor U3105 (N_3105,N_2848,N_2832);
xor U3106 (N_3106,N_2880,N_2887);
nor U3107 (N_3107,N_2888,N_2911);
and U3108 (N_3108,N_2881,N_2872);
nor U3109 (N_3109,N_2915,N_2984);
xor U3110 (N_3110,N_2962,N_2886);
nand U3111 (N_3111,N_2931,N_2830);
nand U3112 (N_3112,N_2858,N_2924);
or U3113 (N_3113,N_2857,N_2806);
xnor U3114 (N_3114,N_2892,N_2913);
or U3115 (N_3115,N_2910,N_2834);
and U3116 (N_3116,N_2875,N_2800);
and U3117 (N_3117,N_2939,N_2868);
nor U3118 (N_3118,N_2810,N_2969);
or U3119 (N_3119,N_2961,N_2830);
or U3120 (N_3120,N_2943,N_2800);
nand U3121 (N_3121,N_2993,N_2803);
nor U3122 (N_3122,N_2842,N_2942);
or U3123 (N_3123,N_2838,N_2988);
and U3124 (N_3124,N_2933,N_2919);
and U3125 (N_3125,N_2898,N_2808);
nand U3126 (N_3126,N_2813,N_2902);
nand U3127 (N_3127,N_2827,N_2832);
nand U3128 (N_3128,N_2871,N_2816);
and U3129 (N_3129,N_2970,N_2934);
and U3130 (N_3130,N_2911,N_2870);
or U3131 (N_3131,N_2862,N_2946);
nand U3132 (N_3132,N_2846,N_2972);
and U3133 (N_3133,N_2996,N_2879);
and U3134 (N_3134,N_2918,N_2965);
nor U3135 (N_3135,N_2847,N_2967);
nor U3136 (N_3136,N_2923,N_2934);
or U3137 (N_3137,N_2814,N_2911);
xor U3138 (N_3138,N_2808,N_2974);
nor U3139 (N_3139,N_2883,N_2813);
xnor U3140 (N_3140,N_2818,N_2853);
nor U3141 (N_3141,N_2818,N_2938);
and U3142 (N_3142,N_2923,N_2822);
nor U3143 (N_3143,N_2917,N_2992);
nand U3144 (N_3144,N_2862,N_2972);
and U3145 (N_3145,N_2916,N_2844);
and U3146 (N_3146,N_2936,N_2983);
or U3147 (N_3147,N_2896,N_2844);
nand U3148 (N_3148,N_2931,N_2855);
nor U3149 (N_3149,N_2909,N_2827);
and U3150 (N_3150,N_2877,N_2964);
nand U3151 (N_3151,N_2813,N_2858);
nand U3152 (N_3152,N_2885,N_2877);
nand U3153 (N_3153,N_2893,N_2918);
nand U3154 (N_3154,N_2820,N_2964);
nand U3155 (N_3155,N_2867,N_2922);
nor U3156 (N_3156,N_2891,N_2827);
and U3157 (N_3157,N_2876,N_2906);
and U3158 (N_3158,N_2927,N_2943);
nand U3159 (N_3159,N_2909,N_2800);
nand U3160 (N_3160,N_2810,N_2861);
or U3161 (N_3161,N_2913,N_2836);
or U3162 (N_3162,N_2944,N_2826);
nor U3163 (N_3163,N_2985,N_2800);
nor U3164 (N_3164,N_2992,N_2874);
xor U3165 (N_3165,N_2967,N_2810);
and U3166 (N_3166,N_2830,N_2932);
xnor U3167 (N_3167,N_2835,N_2853);
nor U3168 (N_3168,N_2868,N_2803);
and U3169 (N_3169,N_2958,N_2806);
or U3170 (N_3170,N_2885,N_2950);
xor U3171 (N_3171,N_2809,N_2841);
nand U3172 (N_3172,N_2828,N_2907);
nor U3173 (N_3173,N_2953,N_2801);
and U3174 (N_3174,N_2827,N_2871);
and U3175 (N_3175,N_2859,N_2824);
and U3176 (N_3176,N_2824,N_2973);
nor U3177 (N_3177,N_2915,N_2859);
or U3178 (N_3178,N_2983,N_2922);
or U3179 (N_3179,N_2879,N_2918);
and U3180 (N_3180,N_2807,N_2983);
or U3181 (N_3181,N_2837,N_2865);
and U3182 (N_3182,N_2810,N_2805);
and U3183 (N_3183,N_2982,N_2837);
xor U3184 (N_3184,N_2964,N_2902);
xnor U3185 (N_3185,N_2974,N_2900);
xor U3186 (N_3186,N_2960,N_2975);
xor U3187 (N_3187,N_2925,N_2958);
and U3188 (N_3188,N_2925,N_2948);
nand U3189 (N_3189,N_2870,N_2847);
nand U3190 (N_3190,N_2822,N_2813);
xor U3191 (N_3191,N_2852,N_2969);
xor U3192 (N_3192,N_2828,N_2930);
nand U3193 (N_3193,N_2826,N_2829);
nor U3194 (N_3194,N_2857,N_2985);
nand U3195 (N_3195,N_2924,N_2912);
nor U3196 (N_3196,N_2829,N_2825);
nand U3197 (N_3197,N_2909,N_2868);
and U3198 (N_3198,N_2943,N_2807);
xnor U3199 (N_3199,N_2887,N_2940);
nand U3200 (N_3200,N_3081,N_3003);
nor U3201 (N_3201,N_3133,N_3039);
xnor U3202 (N_3202,N_3014,N_3076);
nor U3203 (N_3203,N_3082,N_3012);
and U3204 (N_3204,N_3096,N_3086);
nor U3205 (N_3205,N_3038,N_3103);
or U3206 (N_3206,N_3106,N_3060);
or U3207 (N_3207,N_3063,N_3089);
nor U3208 (N_3208,N_3011,N_3113);
nor U3209 (N_3209,N_3020,N_3144);
nor U3210 (N_3210,N_3079,N_3136);
nor U3211 (N_3211,N_3173,N_3025);
xnor U3212 (N_3212,N_3016,N_3049);
xor U3213 (N_3213,N_3057,N_3167);
xor U3214 (N_3214,N_3178,N_3157);
or U3215 (N_3215,N_3108,N_3116);
xor U3216 (N_3216,N_3091,N_3110);
xnor U3217 (N_3217,N_3028,N_3188);
and U3218 (N_3218,N_3042,N_3018);
nand U3219 (N_3219,N_3143,N_3168);
xor U3220 (N_3220,N_3004,N_3111);
nand U3221 (N_3221,N_3069,N_3169);
nor U3222 (N_3222,N_3187,N_3029);
nor U3223 (N_3223,N_3000,N_3033);
and U3224 (N_3224,N_3052,N_3162);
or U3225 (N_3225,N_3185,N_3040);
or U3226 (N_3226,N_3022,N_3154);
or U3227 (N_3227,N_3146,N_3164);
nand U3228 (N_3228,N_3182,N_3026);
and U3229 (N_3229,N_3195,N_3140);
or U3230 (N_3230,N_3002,N_3165);
nor U3231 (N_3231,N_3074,N_3075);
xor U3232 (N_3232,N_3067,N_3114);
nor U3233 (N_3233,N_3083,N_3071);
xor U3234 (N_3234,N_3104,N_3017);
nand U3235 (N_3235,N_3007,N_3027);
nor U3236 (N_3236,N_3019,N_3117);
and U3237 (N_3237,N_3112,N_3088);
xnor U3238 (N_3238,N_3031,N_3070);
nand U3239 (N_3239,N_3066,N_3134);
xnor U3240 (N_3240,N_3189,N_3190);
nor U3241 (N_3241,N_3062,N_3090);
and U3242 (N_3242,N_3056,N_3186);
nand U3243 (N_3243,N_3199,N_3142);
or U3244 (N_3244,N_3045,N_3092);
and U3245 (N_3245,N_3183,N_3051);
and U3246 (N_3246,N_3087,N_3149);
or U3247 (N_3247,N_3135,N_3175);
nand U3248 (N_3248,N_3046,N_3158);
nor U3249 (N_3249,N_3184,N_3148);
nand U3250 (N_3250,N_3196,N_3121);
xnor U3251 (N_3251,N_3137,N_3155);
nor U3252 (N_3252,N_3156,N_3159);
nor U3253 (N_3253,N_3170,N_3115);
and U3254 (N_3254,N_3145,N_3053);
or U3255 (N_3255,N_3109,N_3043);
nor U3256 (N_3256,N_3166,N_3101);
nor U3257 (N_3257,N_3085,N_3153);
nand U3258 (N_3258,N_3160,N_3191);
nor U3259 (N_3259,N_3006,N_3107);
nor U3260 (N_3260,N_3102,N_3163);
nand U3261 (N_3261,N_3094,N_3118);
and U3262 (N_3262,N_3047,N_3098);
xnor U3263 (N_3263,N_3124,N_3129);
and U3264 (N_3264,N_3032,N_3192);
and U3265 (N_3265,N_3127,N_3130);
nand U3266 (N_3266,N_3036,N_3035);
xor U3267 (N_3267,N_3010,N_3198);
xnor U3268 (N_3268,N_3015,N_3123);
or U3269 (N_3269,N_3197,N_3044);
xor U3270 (N_3270,N_3050,N_3030);
or U3271 (N_3271,N_3065,N_3179);
nor U3272 (N_3272,N_3013,N_3024);
nand U3273 (N_3273,N_3001,N_3095);
xor U3274 (N_3274,N_3194,N_3008);
nand U3275 (N_3275,N_3005,N_3084);
or U3276 (N_3276,N_3152,N_3141);
nand U3277 (N_3277,N_3171,N_3105);
xnor U3278 (N_3278,N_3055,N_3122);
xnor U3279 (N_3279,N_3072,N_3119);
or U3280 (N_3280,N_3061,N_3068);
nand U3281 (N_3281,N_3093,N_3037);
or U3282 (N_3282,N_3120,N_3100);
or U3283 (N_3283,N_3150,N_3174);
xnor U3284 (N_3284,N_3126,N_3128);
or U3285 (N_3285,N_3147,N_3161);
and U3286 (N_3286,N_3009,N_3041);
or U3287 (N_3287,N_3097,N_3048);
nand U3288 (N_3288,N_3172,N_3193);
nand U3289 (N_3289,N_3058,N_3080);
xor U3290 (N_3290,N_3021,N_3034);
xnor U3291 (N_3291,N_3099,N_3073);
nand U3292 (N_3292,N_3054,N_3078);
or U3293 (N_3293,N_3131,N_3125);
xor U3294 (N_3294,N_3064,N_3176);
and U3295 (N_3295,N_3151,N_3059);
and U3296 (N_3296,N_3181,N_3023);
xnor U3297 (N_3297,N_3077,N_3138);
xor U3298 (N_3298,N_3139,N_3177);
and U3299 (N_3299,N_3180,N_3132);
nor U3300 (N_3300,N_3039,N_3071);
and U3301 (N_3301,N_3114,N_3021);
nand U3302 (N_3302,N_3168,N_3060);
nand U3303 (N_3303,N_3105,N_3113);
or U3304 (N_3304,N_3161,N_3032);
and U3305 (N_3305,N_3060,N_3019);
xor U3306 (N_3306,N_3169,N_3053);
nand U3307 (N_3307,N_3140,N_3078);
or U3308 (N_3308,N_3017,N_3032);
and U3309 (N_3309,N_3137,N_3177);
and U3310 (N_3310,N_3042,N_3192);
nand U3311 (N_3311,N_3098,N_3029);
or U3312 (N_3312,N_3058,N_3084);
and U3313 (N_3313,N_3096,N_3190);
xor U3314 (N_3314,N_3051,N_3060);
or U3315 (N_3315,N_3176,N_3019);
or U3316 (N_3316,N_3036,N_3015);
nand U3317 (N_3317,N_3082,N_3134);
and U3318 (N_3318,N_3031,N_3037);
xnor U3319 (N_3319,N_3024,N_3127);
xnor U3320 (N_3320,N_3009,N_3095);
or U3321 (N_3321,N_3006,N_3047);
and U3322 (N_3322,N_3111,N_3128);
nor U3323 (N_3323,N_3011,N_3033);
and U3324 (N_3324,N_3135,N_3088);
and U3325 (N_3325,N_3000,N_3071);
nand U3326 (N_3326,N_3121,N_3151);
or U3327 (N_3327,N_3059,N_3092);
xor U3328 (N_3328,N_3129,N_3194);
nor U3329 (N_3329,N_3032,N_3039);
nor U3330 (N_3330,N_3139,N_3082);
nand U3331 (N_3331,N_3097,N_3002);
and U3332 (N_3332,N_3136,N_3167);
nand U3333 (N_3333,N_3084,N_3025);
xnor U3334 (N_3334,N_3080,N_3037);
xor U3335 (N_3335,N_3150,N_3181);
nand U3336 (N_3336,N_3129,N_3030);
xor U3337 (N_3337,N_3006,N_3179);
nand U3338 (N_3338,N_3156,N_3083);
xnor U3339 (N_3339,N_3064,N_3148);
nand U3340 (N_3340,N_3121,N_3079);
nor U3341 (N_3341,N_3161,N_3146);
or U3342 (N_3342,N_3021,N_3092);
and U3343 (N_3343,N_3087,N_3190);
nor U3344 (N_3344,N_3062,N_3129);
and U3345 (N_3345,N_3111,N_3114);
nand U3346 (N_3346,N_3151,N_3072);
nand U3347 (N_3347,N_3064,N_3007);
and U3348 (N_3348,N_3130,N_3124);
and U3349 (N_3349,N_3071,N_3031);
nor U3350 (N_3350,N_3173,N_3093);
nand U3351 (N_3351,N_3083,N_3016);
nand U3352 (N_3352,N_3198,N_3083);
xnor U3353 (N_3353,N_3155,N_3003);
nand U3354 (N_3354,N_3085,N_3195);
nand U3355 (N_3355,N_3147,N_3039);
nor U3356 (N_3356,N_3098,N_3074);
and U3357 (N_3357,N_3009,N_3066);
and U3358 (N_3358,N_3009,N_3177);
nand U3359 (N_3359,N_3115,N_3049);
nand U3360 (N_3360,N_3194,N_3155);
nor U3361 (N_3361,N_3003,N_3158);
and U3362 (N_3362,N_3112,N_3086);
or U3363 (N_3363,N_3090,N_3118);
xor U3364 (N_3364,N_3131,N_3169);
nand U3365 (N_3365,N_3079,N_3147);
or U3366 (N_3366,N_3161,N_3014);
or U3367 (N_3367,N_3104,N_3175);
nand U3368 (N_3368,N_3094,N_3014);
or U3369 (N_3369,N_3189,N_3000);
nor U3370 (N_3370,N_3034,N_3089);
nand U3371 (N_3371,N_3191,N_3093);
xnor U3372 (N_3372,N_3011,N_3082);
nor U3373 (N_3373,N_3154,N_3171);
or U3374 (N_3374,N_3176,N_3186);
xor U3375 (N_3375,N_3047,N_3126);
nand U3376 (N_3376,N_3141,N_3092);
xor U3377 (N_3377,N_3119,N_3022);
or U3378 (N_3378,N_3028,N_3126);
and U3379 (N_3379,N_3125,N_3018);
nor U3380 (N_3380,N_3050,N_3022);
nand U3381 (N_3381,N_3010,N_3024);
xnor U3382 (N_3382,N_3194,N_3158);
or U3383 (N_3383,N_3042,N_3051);
xor U3384 (N_3384,N_3093,N_3147);
and U3385 (N_3385,N_3016,N_3105);
or U3386 (N_3386,N_3158,N_3099);
nor U3387 (N_3387,N_3151,N_3031);
or U3388 (N_3388,N_3092,N_3043);
and U3389 (N_3389,N_3035,N_3094);
nand U3390 (N_3390,N_3044,N_3036);
xor U3391 (N_3391,N_3027,N_3180);
xnor U3392 (N_3392,N_3188,N_3128);
nor U3393 (N_3393,N_3120,N_3093);
nand U3394 (N_3394,N_3094,N_3182);
nor U3395 (N_3395,N_3121,N_3193);
or U3396 (N_3396,N_3027,N_3135);
nand U3397 (N_3397,N_3018,N_3116);
and U3398 (N_3398,N_3100,N_3193);
nor U3399 (N_3399,N_3145,N_3153);
and U3400 (N_3400,N_3312,N_3287);
or U3401 (N_3401,N_3202,N_3272);
or U3402 (N_3402,N_3271,N_3256);
and U3403 (N_3403,N_3374,N_3263);
and U3404 (N_3404,N_3297,N_3356);
or U3405 (N_3405,N_3361,N_3336);
or U3406 (N_3406,N_3252,N_3317);
nand U3407 (N_3407,N_3338,N_3227);
nand U3408 (N_3408,N_3396,N_3214);
and U3409 (N_3409,N_3388,N_3352);
xor U3410 (N_3410,N_3372,N_3373);
or U3411 (N_3411,N_3275,N_3264);
nor U3412 (N_3412,N_3237,N_3207);
or U3413 (N_3413,N_3344,N_3323);
and U3414 (N_3414,N_3333,N_3395);
or U3415 (N_3415,N_3345,N_3258);
nor U3416 (N_3416,N_3239,N_3268);
and U3417 (N_3417,N_3234,N_3328);
nor U3418 (N_3418,N_3203,N_3254);
nand U3419 (N_3419,N_3353,N_3224);
xnor U3420 (N_3420,N_3211,N_3267);
xor U3421 (N_3421,N_3209,N_3307);
xnor U3422 (N_3422,N_3376,N_3285);
and U3423 (N_3423,N_3265,N_3358);
nand U3424 (N_3424,N_3380,N_3223);
nand U3425 (N_3425,N_3289,N_3226);
xor U3426 (N_3426,N_3398,N_3300);
nor U3427 (N_3427,N_3269,N_3213);
or U3428 (N_3428,N_3340,N_3343);
nand U3429 (N_3429,N_3377,N_3246);
xnor U3430 (N_3430,N_3393,N_3219);
nor U3431 (N_3431,N_3248,N_3277);
nand U3432 (N_3432,N_3389,N_3257);
or U3433 (N_3433,N_3278,N_3316);
or U3434 (N_3434,N_3337,N_3291);
and U3435 (N_3435,N_3390,N_3384);
and U3436 (N_3436,N_3200,N_3362);
or U3437 (N_3437,N_3304,N_3230);
nand U3438 (N_3438,N_3310,N_3319);
xnor U3439 (N_3439,N_3397,N_3235);
or U3440 (N_3440,N_3279,N_3220);
nand U3441 (N_3441,N_3222,N_3311);
xnor U3442 (N_3442,N_3244,N_3309);
nand U3443 (N_3443,N_3386,N_3321);
or U3444 (N_3444,N_3332,N_3243);
xor U3445 (N_3445,N_3253,N_3331);
xnor U3446 (N_3446,N_3349,N_3280);
and U3447 (N_3447,N_3341,N_3357);
nor U3448 (N_3448,N_3329,N_3273);
nor U3449 (N_3449,N_3205,N_3301);
or U3450 (N_3450,N_3387,N_3232);
xnor U3451 (N_3451,N_3318,N_3313);
nor U3452 (N_3452,N_3355,N_3382);
nand U3453 (N_3453,N_3201,N_3363);
nor U3454 (N_3454,N_3378,N_3283);
and U3455 (N_3455,N_3351,N_3281);
or U3456 (N_3456,N_3262,N_3231);
or U3457 (N_3457,N_3294,N_3322);
or U3458 (N_3458,N_3293,N_3216);
and U3459 (N_3459,N_3247,N_3303);
and U3460 (N_3460,N_3290,N_3369);
and U3461 (N_3461,N_3210,N_3391);
nand U3462 (N_3462,N_3324,N_3367);
nand U3463 (N_3463,N_3233,N_3326);
nor U3464 (N_3464,N_3302,N_3276);
and U3465 (N_3465,N_3347,N_3270);
or U3466 (N_3466,N_3298,N_3330);
nor U3467 (N_3467,N_3334,N_3348);
nand U3468 (N_3468,N_3305,N_3241);
nand U3469 (N_3469,N_3259,N_3274);
nand U3470 (N_3470,N_3217,N_3370);
xor U3471 (N_3471,N_3229,N_3260);
or U3472 (N_3472,N_3365,N_3394);
xor U3473 (N_3473,N_3206,N_3250);
xor U3474 (N_3474,N_3299,N_3315);
and U3475 (N_3475,N_3245,N_3379);
nor U3476 (N_3476,N_3335,N_3339);
nor U3477 (N_3477,N_3251,N_3212);
xnor U3478 (N_3478,N_3366,N_3383);
and U3479 (N_3479,N_3266,N_3359);
and U3480 (N_3480,N_3236,N_3385);
and U3481 (N_3481,N_3399,N_3306);
nand U3482 (N_3482,N_3371,N_3346);
and U3483 (N_3483,N_3238,N_3288);
nand U3484 (N_3484,N_3221,N_3296);
or U3485 (N_3485,N_3295,N_3225);
nor U3486 (N_3486,N_3392,N_3215);
xor U3487 (N_3487,N_3375,N_3350);
nand U3488 (N_3488,N_3354,N_3240);
xor U3489 (N_3489,N_3292,N_3368);
or U3490 (N_3490,N_3325,N_3282);
xor U3491 (N_3491,N_3342,N_3249);
or U3492 (N_3492,N_3286,N_3218);
nand U3493 (N_3493,N_3284,N_3327);
or U3494 (N_3494,N_3320,N_3261);
nand U3495 (N_3495,N_3255,N_3228);
and U3496 (N_3496,N_3208,N_3314);
nand U3497 (N_3497,N_3364,N_3242);
xor U3498 (N_3498,N_3308,N_3204);
nor U3499 (N_3499,N_3381,N_3360);
nor U3500 (N_3500,N_3356,N_3339);
nor U3501 (N_3501,N_3264,N_3397);
nand U3502 (N_3502,N_3325,N_3224);
nor U3503 (N_3503,N_3393,N_3256);
nand U3504 (N_3504,N_3278,N_3214);
and U3505 (N_3505,N_3215,N_3324);
or U3506 (N_3506,N_3378,N_3272);
and U3507 (N_3507,N_3312,N_3210);
nor U3508 (N_3508,N_3245,N_3244);
nor U3509 (N_3509,N_3216,N_3214);
nor U3510 (N_3510,N_3382,N_3364);
or U3511 (N_3511,N_3268,N_3371);
nand U3512 (N_3512,N_3313,N_3391);
nor U3513 (N_3513,N_3200,N_3209);
and U3514 (N_3514,N_3375,N_3259);
nand U3515 (N_3515,N_3304,N_3233);
nand U3516 (N_3516,N_3383,N_3292);
or U3517 (N_3517,N_3241,N_3266);
or U3518 (N_3518,N_3292,N_3359);
xor U3519 (N_3519,N_3280,N_3376);
nor U3520 (N_3520,N_3253,N_3286);
nand U3521 (N_3521,N_3394,N_3393);
nor U3522 (N_3522,N_3328,N_3305);
or U3523 (N_3523,N_3282,N_3378);
xnor U3524 (N_3524,N_3229,N_3290);
xor U3525 (N_3525,N_3264,N_3308);
xor U3526 (N_3526,N_3304,N_3297);
and U3527 (N_3527,N_3215,N_3250);
or U3528 (N_3528,N_3334,N_3226);
xnor U3529 (N_3529,N_3316,N_3227);
and U3530 (N_3530,N_3252,N_3366);
and U3531 (N_3531,N_3379,N_3263);
nand U3532 (N_3532,N_3304,N_3339);
xnor U3533 (N_3533,N_3241,N_3301);
xor U3534 (N_3534,N_3236,N_3255);
xnor U3535 (N_3535,N_3250,N_3217);
and U3536 (N_3536,N_3281,N_3337);
and U3537 (N_3537,N_3208,N_3362);
nand U3538 (N_3538,N_3270,N_3326);
nand U3539 (N_3539,N_3352,N_3272);
and U3540 (N_3540,N_3384,N_3327);
xnor U3541 (N_3541,N_3282,N_3309);
and U3542 (N_3542,N_3208,N_3289);
and U3543 (N_3543,N_3371,N_3261);
nand U3544 (N_3544,N_3374,N_3334);
or U3545 (N_3545,N_3275,N_3257);
and U3546 (N_3546,N_3336,N_3283);
or U3547 (N_3547,N_3253,N_3327);
nand U3548 (N_3548,N_3325,N_3395);
and U3549 (N_3549,N_3389,N_3376);
nor U3550 (N_3550,N_3284,N_3238);
nand U3551 (N_3551,N_3287,N_3329);
and U3552 (N_3552,N_3334,N_3376);
or U3553 (N_3553,N_3320,N_3235);
and U3554 (N_3554,N_3264,N_3343);
and U3555 (N_3555,N_3291,N_3213);
and U3556 (N_3556,N_3279,N_3326);
nand U3557 (N_3557,N_3355,N_3296);
nand U3558 (N_3558,N_3358,N_3293);
and U3559 (N_3559,N_3203,N_3397);
and U3560 (N_3560,N_3375,N_3271);
nor U3561 (N_3561,N_3274,N_3366);
xor U3562 (N_3562,N_3319,N_3216);
and U3563 (N_3563,N_3338,N_3263);
nand U3564 (N_3564,N_3354,N_3324);
and U3565 (N_3565,N_3362,N_3375);
or U3566 (N_3566,N_3350,N_3347);
and U3567 (N_3567,N_3274,N_3260);
nand U3568 (N_3568,N_3268,N_3396);
and U3569 (N_3569,N_3257,N_3224);
xor U3570 (N_3570,N_3216,N_3317);
and U3571 (N_3571,N_3254,N_3211);
xor U3572 (N_3572,N_3376,N_3384);
or U3573 (N_3573,N_3350,N_3367);
nand U3574 (N_3574,N_3308,N_3223);
or U3575 (N_3575,N_3249,N_3228);
nand U3576 (N_3576,N_3202,N_3338);
xnor U3577 (N_3577,N_3349,N_3246);
nor U3578 (N_3578,N_3382,N_3396);
and U3579 (N_3579,N_3315,N_3246);
and U3580 (N_3580,N_3231,N_3324);
or U3581 (N_3581,N_3302,N_3297);
nand U3582 (N_3582,N_3377,N_3233);
or U3583 (N_3583,N_3383,N_3356);
nand U3584 (N_3584,N_3293,N_3340);
or U3585 (N_3585,N_3346,N_3298);
nand U3586 (N_3586,N_3261,N_3326);
nor U3587 (N_3587,N_3315,N_3215);
nand U3588 (N_3588,N_3206,N_3246);
nand U3589 (N_3589,N_3251,N_3290);
xnor U3590 (N_3590,N_3240,N_3244);
xor U3591 (N_3591,N_3384,N_3301);
nand U3592 (N_3592,N_3257,N_3246);
xnor U3593 (N_3593,N_3284,N_3260);
nand U3594 (N_3594,N_3317,N_3267);
and U3595 (N_3595,N_3373,N_3202);
nand U3596 (N_3596,N_3342,N_3285);
or U3597 (N_3597,N_3235,N_3386);
xnor U3598 (N_3598,N_3225,N_3203);
or U3599 (N_3599,N_3335,N_3366);
nor U3600 (N_3600,N_3517,N_3415);
xor U3601 (N_3601,N_3524,N_3430);
nand U3602 (N_3602,N_3449,N_3538);
nand U3603 (N_3603,N_3539,N_3411);
xnor U3604 (N_3604,N_3454,N_3514);
nand U3605 (N_3605,N_3552,N_3495);
xor U3606 (N_3606,N_3402,N_3545);
nand U3607 (N_3607,N_3522,N_3544);
nand U3608 (N_3608,N_3547,N_3442);
nor U3609 (N_3609,N_3407,N_3473);
xor U3610 (N_3610,N_3497,N_3464);
or U3611 (N_3611,N_3462,N_3597);
or U3612 (N_3612,N_3559,N_3551);
nor U3613 (N_3613,N_3558,N_3416);
nand U3614 (N_3614,N_3577,N_3422);
xor U3615 (N_3615,N_3479,N_3516);
nor U3616 (N_3616,N_3492,N_3521);
and U3617 (N_3617,N_3489,N_3465);
nand U3618 (N_3618,N_3532,N_3571);
nand U3619 (N_3619,N_3595,N_3427);
and U3620 (N_3620,N_3406,N_3490);
or U3621 (N_3621,N_3588,N_3506);
and U3622 (N_3622,N_3400,N_3535);
xnor U3623 (N_3623,N_3596,N_3556);
nand U3624 (N_3624,N_3537,N_3515);
xnor U3625 (N_3625,N_3429,N_3513);
and U3626 (N_3626,N_3459,N_3484);
nor U3627 (N_3627,N_3448,N_3441);
or U3628 (N_3628,N_3564,N_3580);
nor U3629 (N_3629,N_3549,N_3413);
or U3630 (N_3630,N_3414,N_3557);
and U3631 (N_3631,N_3421,N_3566);
or U3632 (N_3632,N_3498,N_3599);
or U3633 (N_3633,N_3472,N_3423);
and U3634 (N_3634,N_3589,N_3584);
and U3635 (N_3635,N_3534,N_3579);
nor U3636 (N_3636,N_3582,N_3512);
nand U3637 (N_3637,N_3541,N_3494);
or U3638 (N_3638,N_3468,N_3563);
or U3639 (N_3639,N_3426,N_3530);
nor U3640 (N_3640,N_3403,N_3425);
nand U3641 (N_3641,N_3446,N_3405);
xor U3642 (N_3642,N_3573,N_3554);
or U3643 (N_3643,N_3543,N_3508);
and U3644 (N_3644,N_3594,N_3493);
nand U3645 (N_3645,N_3451,N_3452);
nor U3646 (N_3646,N_3504,N_3592);
xor U3647 (N_3647,N_3478,N_3457);
or U3648 (N_3648,N_3540,N_3439);
or U3649 (N_3649,N_3455,N_3433);
nand U3650 (N_3650,N_3434,N_3436);
and U3651 (N_3651,N_3410,N_3401);
xnor U3652 (N_3652,N_3466,N_3431);
xnor U3653 (N_3653,N_3503,N_3420);
nand U3654 (N_3654,N_3550,N_3458);
xnor U3655 (N_3655,N_3586,N_3435);
and U3656 (N_3656,N_3443,N_3419);
nand U3657 (N_3657,N_3553,N_3501);
or U3658 (N_3658,N_3502,N_3590);
nor U3659 (N_3659,N_3569,N_3483);
nor U3660 (N_3660,N_3536,N_3475);
nor U3661 (N_3661,N_3499,N_3424);
nor U3662 (N_3662,N_3477,N_3404);
xor U3663 (N_3663,N_3505,N_3519);
nand U3664 (N_3664,N_3531,N_3445);
or U3665 (N_3665,N_3507,N_3518);
xor U3666 (N_3666,N_3574,N_3591);
nand U3667 (N_3667,N_3418,N_3438);
or U3668 (N_3668,N_3480,N_3523);
xor U3669 (N_3669,N_3461,N_3528);
nor U3670 (N_3670,N_3510,N_3412);
nand U3671 (N_3671,N_3575,N_3437);
nor U3672 (N_3672,N_3585,N_3565);
and U3673 (N_3673,N_3496,N_3444);
and U3674 (N_3674,N_3568,N_3511);
nand U3675 (N_3675,N_3560,N_3525);
nand U3676 (N_3676,N_3587,N_3481);
xnor U3677 (N_3677,N_3527,N_3428);
and U3678 (N_3678,N_3409,N_3476);
or U3679 (N_3679,N_3533,N_3487);
xor U3680 (N_3680,N_3432,N_3485);
nand U3681 (N_3681,N_3598,N_3546);
and U3682 (N_3682,N_3520,N_3562);
xnor U3683 (N_3683,N_3576,N_3500);
nand U3684 (N_3684,N_3488,N_3471);
and U3685 (N_3685,N_3529,N_3456);
and U3686 (N_3686,N_3572,N_3470);
or U3687 (N_3687,N_3570,N_3482);
and U3688 (N_3688,N_3509,N_3453);
nor U3689 (N_3689,N_3578,N_3491);
nand U3690 (N_3690,N_3474,N_3467);
xnor U3691 (N_3691,N_3450,N_3581);
xnor U3692 (N_3692,N_3561,N_3417);
and U3693 (N_3693,N_3567,N_3447);
nand U3694 (N_3694,N_3486,N_3542);
or U3695 (N_3695,N_3593,N_3469);
nor U3696 (N_3696,N_3463,N_3583);
or U3697 (N_3697,N_3555,N_3548);
nand U3698 (N_3698,N_3440,N_3460);
nor U3699 (N_3699,N_3408,N_3526);
nor U3700 (N_3700,N_3551,N_3449);
and U3701 (N_3701,N_3418,N_3511);
nand U3702 (N_3702,N_3558,N_3421);
and U3703 (N_3703,N_3479,N_3519);
nand U3704 (N_3704,N_3450,N_3454);
or U3705 (N_3705,N_3423,N_3587);
nor U3706 (N_3706,N_3450,N_3548);
or U3707 (N_3707,N_3557,N_3579);
and U3708 (N_3708,N_3543,N_3475);
nand U3709 (N_3709,N_3415,N_3483);
and U3710 (N_3710,N_3537,N_3560);
nor U3711 (N_3711,N_3513,N_3445);
and U3712 (N_3712,N_3439,N_3417);
nand U3713 (N_3713,N_3468,N_3597);
nand U3714 (N_3714,N_3537,N_3506);
or U3715 (N_3715,N_3572,N_3479);
nand U3716 (N_3716,N_3559,N_3566);
nand U3717 (N_3717,N_3520,N_3428);
xor U3718 (N_3718,N_3582,N_3547);
or U3719 (N_3719,N_3529,N_3552);
and U3720 (N_3720,N_3459,N_3429);
nand U3721 (N_3721,N_3591,N_3511);
xnor U3722 (N_3722,N_3595,N_3540);
or U3723 (N_3723,N_3560,N_3576);
nand U3724 (N_3724,N_3464,N_3573);
nand U3725 (N_3725,N_3531,N_3529);
xor U3726 (N_3726,N_3551,N_3436);
nand U3727 (N_3727,N_3546,N_3495);
nor U3728 (N_3728,N_3554,N_3471);
and U3729 (N_3729,N_3533,N_3588);
or U3730 (N_3730,N_3521,N_3448);
nand U3731 (N_3731,N_3549,N_3457);
xnor U3732 (N_3732,N_3445,N_3518);
xnor U3733 (N_3733,N_3479,N_3501);
nor U3734 (N_3734,N_3563,N_3494);
nand U3735 (N_3735,N_3558,N_3533);
nor U3736 (N_3736,N_3597,N_3449);
and U3737 (N_3737,N_3527,N_3471);
and U3738 (N_3738,N_3416,N_3577);
or U3739 (N_3739,N_3487,N_3485);
xor U3740 (N_3740,N_3536,N_3559);
and U3741 (N_3741,N_3451,N_3529);
nor U3742 (N_3742,N_3592,N_3530);
nor U3743 (N_3743,N_3513,N_3424);
or U3744 (N_3744,N_3593,N_3505);
nor U3745 (N_3745,N_3463,N_3558);
or U3746 (N_3746,N_3453,N_3553);
xnor U3747 (N_3747,N_3529,N_3491);
nor U3748 (N_3748,N_3437,N_3492);
and U3749 (N_3749,N_3546,N_3571);
xor U3750 (N_3750,N_3458,N_3563);
xnor U3751 (N_3751,N_3456,N_3515);
or U3752 (N_3752,N_3515,N_3433);
nor U3753 (N_3753,N_3548,N_3466);
and U3754 (N_3754,N_3499,N_3553);
nor U3755 (N_3755,N_3593,N_3590);
xor U3756 (N_3756,N_3448,N_3487);
nor U3757 (N_3757,N_3418,N_3538);
and U3758 (N_3758,N_3507,N_3596);
or U3759 (N_3759,N_3535,N_3528);
or U3760 (N_3760,N_3536,N_3439);
nand U3761 (N_3761,N_3595,N_3413);
and U3762 (N_3762,N_3548,N_3585);
or U3763 (N_3763,N_3428,N_3523);
nand U3764 (N_3764,N_3520,N_3589);
nor U3765 (N_3765,N_3485,N_3511);
and U3766 (N_3766,N_3436,N_3547);
nand U3767 (N_3767,N_3560,N_3400);
or U3768 (N_3768,N_3578,N_3596);
and U3769 (N_3769,N_3417,N_3544);
nor U3770 (N_3770,N_3564,N_3422);
and U3771 (N_3771,N_3554,N_3432);
xnor U3772 (N_3772,N_3475,N_3407);
nor U3773 (N_3773,N_3511,N_3446);
nand U3774 (N_3774,N_3582,N_3474);
or U3775 (N_3775,N_3473,N_3520);
xnor U3776 (N_3776,N_3437,N_3547);
nand U3777 (N_3777,N_3493,N_3513);
nand U3778 (N_3778,N_3443,N_3553);
xnor U3779 (N_3779,N_3416,N_3569);
nand U3780 (N_3780,N_3522,N_3540);
nor U3781 (N_3781,N_3500,N_3527);
nor U3782 (N_3782,N_3567,N_3507);
or U3783 (N_3783,N_3442,N_3421);
xnor U3784 (N_3784,N_3447,N_3532);
nand U3785 (N_3785,N_3465,N_3557);
and U3786 (N_3786,N_3599,N_3403);
nor U3787 (N_3787,N_3596,N_3592);
and U3788 (N_3788,N_3523,N_3467);
and U3789 (N_3789,N_3458,N_3444);
or U3790 (N_3790,N_3510,N_3467);
or U3791 (N_3791,N_3438,N_3494);
or U3792 (N_3792,N_3577,N_3572);
and U3793 (N_3793,N_3526,N_3488);
xor U3794 (N_3794,N_3505,N_3559);
xor U3795 (N_3795,N_3559,N_3596);
and U3796 (N_3796,N_3522,N_3473);
or U3797 (N_3797,N_3549,N_3412);
or U3798 (N_3798,N_3457,N_3414);
xnor U3799 (N_3799,N_3567,N_3453);
nor U3800 (N_3800,N_3612,N_3652);
and U3801 (N_3801,N_3759,N_3797);
nor U3802 (N_3802,N_3795,N_3656);
nand U3803 (N_3803,N_3735,N_3604);
nor U3804 (N_3804,N_3637,N_3617);
nor U3805 (N_3805,N_3746,N_3635);
or U3806 (N_3806,N_3703,N_3672);
xnor U3807 (N_3807,N_3794,N_3654);
or U3808 (N_3808,N_3718,N_3695);
or U3809 (N_3809,N_3751,N_3753);
and U3810 (N_3810,N_3742,N_3616);
nor U3811 (N_3811,N_3680,N_3688);
nor U3812 (N_3812,N_3793,N_3778);
nor U3813 (N_3813,N_3646,N_3723);
and U3814 (N_3814,N_3770,N_3701);
nor U3815 (N_3815,N_3705,N_3775);
and U3816 (N_3816,N_3752,N_3730);
nor U3817 (N_3817,N_3645,N_3769);
or U3818 (N_3818,N_3639,N_3766);
nand U3819 (N_3819,N_3749,N_3613);
nor U3820 (N_3820,N_3761,N_3748);
and U3821 (N_3821,N_3606,N_3659);
xor U3822 (N_3822,N_3707,N_3643);
or U3823 (N_3823,N_3649,N_3763);
or U3824 (N_3824,N_3711,N_3663);
nand U3825 (N_3825,N_3762,N_3768);
nand U3826 (N_3826,N_3697,N_3605);
nand U3827 (N_3827,N_3736,N_3626);
and U3828 (N_3828,N_3683,N_3782);
nand U3829 (N_3829,N_3758,N_3765);
nor U3830 (N_3830,N_3733,N_3610);
nand U3831 (N_3831,N_3726,N_3615);
and U3832 (N_3832,N_3764,N_3727);
or U3833 (N_3833,N_3690,N_3771);
nand U3834 (N_3834,N_3757,N_3774);
nand U3835 (N_3835,N_3756,N_3798);
and U3836 (N_3836,N_3673,N_3648);
or U3837 (N_3837,N_3719,N_3618);
nand U3838 (N_3838,N_3651,N_3712);
or U3839 (N_3839,N_3738,N_3647);
or U3840 (N_3840,N_3787,N_3745);
nand U3841 (N_3841,N_3729,N_3603);
nand U3842 (N_3842,N_3731,N_3661);
xor U3843 (N_3843,N_3725,N_3772);
and U3844 (N_3844,N_3668,N_3693);
or U3845 (N_3845,N_3796,N_3644);
xor U3846 (N_3846,N_3621,N_3678);
nand U3847 (N_3847,N_3722,N_3706);
and U3848 (N_3848,N_3653,N_3658);
and U3849 (N_3849,N_3676,N_3602);
nor U3850 (N_3850,N_3627,N_3620);
xnor U3851 (N_3851,N_3657,N_3691);
nand U3852 (N_3852,N_3767,N_3669);
or U3853 (N_3853,N_3721,N_3624);
xor U3854 (N_3854,N_3664,N_3720);
nand U3855 (N_3855,N_3694,N_3609);
xor U3856 (N_3856,N_3785,N_3783);
xor U3857 (N_3857,N_3716,N_3781);
nand U3858 (N_3858,N_3760,N_3717);
xnor U3859 (N_3859,N_3641,N_3777);
or U3860 (N_3860,N_3619,N_3743);
nand U3861 (N_3861,N_3611,N_3724);
or U3862 (N_3862,N_3642,N_3786);
xnor U3863 (N_3863,N_3773,N_3715);
nor U3864 (N_3864,N_3698,N_3709);
xor U3865 (N_3865,N_3686,N_3629);
and U3866 (N_3866,N_3739,N_3702);
or U3867 (N_3867,N_3754,N_3666);
nand U3868 (N_3868,N_3684,N_3789);
xor U3869 (N_3869,N_3671,N_3640);
or U3870 (N_3870,N_3700,N_3708);
xnor U3871 (N_3871,N_3655,N_3631);
or U3872 (N_3872,N_3681,N_3674);
nand U3873 (N_3873,N_3662,N_3670);
nor U3874 (N_3874,N_3734,N_3638);
xor U3875 (N_3875,N_3792,N_3632);
and U3876 (N_3876,N_3732,N_3685);
and U3877 (N_3877,N_3665,N_3625);
nor U3878 (N_3878,N_3636,N_3623);
nor U3879 (N_3879,N_3714,N_3601);
nor U3880 (N_3880,N_3784,N_3689);
or U3881 (N_3881,N_3750,N_3704);
xor U3882 (N_3882,N_3744,N_3628);
nand U3883 (N_3883,N_3692,N_3740);
xnor U3884 (N_3884,N_3622,N_3713);
nor U3885 (N_3885,N_3675,N_3607);
or U3886 (N_3886,N_3699,N_3696);
and U3887 (N_3887,N_3776,N_3650);
or U3888 (N_3888,N_3788,N_3679);
nor U3889 (N_3889,N_3600,N_3633);
and U3890 (N_3890,N_3737,N_3634);
nand U3891 (N_3891,N_3790,N_3660);
and U3892 (N_3892,N_3614,N_3608);
nor U3893 (N_3893,N_3667,N_3677);
xor U3894 (N_3894,N_3710,N_3630);
nor U3895 (N_3895,N_3747,N_3728);
nand U3896 (N_3896,N_3741,N_3682);
nand U3897 (N_3897,N_3779,N_3755);
and U3898 (N_3898,N_3799,N_3791);
xor U3899 (N_3899,N_3687,N_3780);
nor U3900 (N_3900,N_3642,N_3794);
and U3901 (N_3901,N_3796,N_3791);
xnor U3902 (N_3902,N_3710,N_3691);
nand U3903 (N_3903,N_3670,N_3619);
or U3904 (N_3904,N_3720,N_3698);
or U3905 (N_3905,N_3665,N_3601);
xnor U3906 (N_3906,N_3776,N_3721);
nor U3907 (N_3907,N_3774,N_3645);
xnor U3908 (N_3908,N_3703,N_3601);
nor U3909 (N_3909,N_3780,N_3775);
and U3910 (N_3910,N_3675,N_3672);
nor U3911 (N_3911,N_3793,N_3682);
xor U3912 (N_3912,N_3661,N_3708);
and U3913 (N_3913,N_3750,N_3644);
xor U3914 (N_3914,N_3764,N_3690);
nor U3915 (N_3915,N_3753,N_3613);
xnor U3916 (N_3916,N_3650,N_3648);
xnor U3917 (N_3917,N_3680,N_3630);
or U3918 (N_3918,N_3693,N_3756);
nand U3919 (N_3919,N_3686,N_3753);
or U3920 (N_3920,N_3670,N_3724);
nand U3921 (N_3921,N_3712,N_3697);
nand U3922 (N_3922,N_3694,N_3674);
and U3923 (N_3923,N_3712,N_3654);
xor U3924 (N_3924,N_3697,N_3668);
nand U3925 (N_3925,N_3793,N_3701);
nor U3926 (N_3926,N_3702,N_3638);
nand U3927 (N_3927,N_3698,N_3604);
xnor U3928 (N_3928,N_3796,N_3776);
nor U3929 (N_3929,N_3781,N_3731);
xnor U3930 (N_3930,N_3674,N_3710);
nor U3931 (N_3931,N_3792,N_3691);
nand U3932 (N_3932,N_3671,N_3719);
and U3933 (N_3933,N_3629,N_3684);
nor U3934 (N_3934,N_3749,N_3724);
and U3935 (N_3935,N_3725,N_3651);
xnor U3936 (N_3936,N_3692,N_3715);
xor U3937 (N_3937,N_3691,N_3752);
and U3938 (N_3938,N_3794,N_3694);
nor U3939 (N_3939,N_3614,N_3697);
nand U3940 (N_3940,N_3771,N_3699);
xnor U3941 (N_3941,N_3667,N_3665);
or U3942 (N_3942,N_3669,N_3716);
or U3943 (N_3943,N_3611,N_3602);
xnor U3944 (N_3944,N_3667,N_3649);
nand U3945 (N_3945,N_3683,N_3670);
or U3946 (N_3946,N_3604,N_3660);
nor U3947 (N_3947,N_3746,N_3628);
or U3948 (N_3948,N_3686,N_3759);
or U3949 (N_3949,N_3787,N_3784);
and U3950 (N_3950,N_3664,N_3648);
xor U3951 (N_3951,N_3601,N_3771);
nand U3952 (N_3952,N_3735,N_3700);
or U3953 (N_3953,N_3671,N_3626);
nor U3954 (N_3954,N_3651,N_3683);
nand U3955 (N_3955,N_3666,N_3683);
nor U3956 (N_3956,N_3671,N_3690);
and U3957 (N_3957,N_3710,N_3724);
xor U3958 (N_3958,N_3729,N_3623);
nand U3959 (N_3959,N_3621,N_3797);
nand U3960 (N_3960,N_3685,N_3770);
and U3961 (N_3961,N_3638,N_3754);
nand U3962 (N_3962,N_3777,N_3632);
nor U3963 (N_3963,N_3624,N_3617);
xnor U3964 (N_3964,N_3655,N_3650);
and U3965 (N_3965,N_3688,N_3700);
nor U3966 (N_3966,N_3663,N_3635);
nor U3967 (N_3967,N_3659,N_3680);
xnor U3968 (N_3968,N_3676,N_3660);
and U3969 (N_3969,N_3783,N_3763);
nand U3970 (N_3970,N_3666,N_3737);
or U3971 (N_3971,N_3631,N_3754);
nand U3972 (N_3972,N_3602,N_3722);
or U3973 (N_3973,N_3673,N_3678);
and U3974 (N_3974,N_3681,N_3613);
xnor U3975 (N_3975,N_3644,N_3777);
and U3976 (N_3976,N_3765,N_3786);
xor U3977 (N_3977,N_3764,N_3677);
nand U3978 (N_3978,N_3726,N_3757);
or U3979 (N_3979,N_3632,N_3620);
or U3980 (N_3980,N_3778,N_3759);
xor U3981 (N_3981,N_3739,N_3616);
nor U3982 (N_3982,N_3752,N_3733);
nand U3983 (N_3983,N_3728,N_3777);
or U3984 (N_3984,N_3612,N_3643);
and U3985 (N_3985,N_3655,N_3749);
xnor U3986 (N_3986,N_3657,N_3653);
and U3987 (N_3987,N_3623,N_3797);
or U3988 (N_3988,N_3736,N_3723);
and U3989 (N_3989,N_3640,N_3697);
nand U3990 (N_3990,N_3605,N_3709);
and U3991 (N_3991,N_3783,N_3703);
xor U3992 (N_3992,N_3644,N_3707);
nor U3993 (N_3993,N_3708,N_3782);
nand U3994 (N_3994,N_3635,N_3782);
or U3995 (N_3995,N_3765,N_3669);
xnor U3996 (N_3996,N_3721,N_3760);
and U3997 (N_3997,N_3614,N_3623);
nor U3998 (N_3998,N_3774,N_3771);
nand U3999 (N_3999,N_3707,N_3733);
nor U4000 (N_4000,N_3949,N_3805);
xor U4001 (N_4001,N_3939,N_3897);
nand U4002 (N_4002,N_3832,N_3906);
nor U4003 (N_4003,N_3820,N_3872);
xnor U4004 (N_4004,N_3887,N_3888);
and U4005 (N_4005,N_3837,N_3978);
xnor U4006 (N_4006,N_3833,N_3974);
nor U4007 (N_4007,N_3952,N_3899);
nand U4008 (N_4008,N_3990,N_3986);
and U4009 (N_4009,N_3890,N_3854);
nand U4010 (N_4010,N_3848,N_3898);
and U4011 (N_4011,N_3896,N_3958);
or U4012 (N_4012,N_3876,N_3992);
xor U4013 (N_4013,N_3807,N_3856);
nor U4014 (N_4014,N_3991,N_3847);
and U4015 (N_4015,N_3983,N_3968);
xnor U4016 (N_4016,N_3989,N_3932);
xnor U4017 (N_4017,N_3829,N_3886);
xnor U4018 (N_4018,N_3919,N_3916);
and U4019 (N_4019,N_3971,N_3944);
and U4020 (N_4020,N_3937,N_3948);
and U4021 (N_4021,N_3933,N_3843);
xnor U4022 (N_4022,N_3950,N_3883);
and U4023 (N_4023,N_3809,N_3825);
and U4024 (N_4024,N_3976,N_3925);
and U4025 (N_4025,N_3884,N_3965);
nor U4026 (N_4026,N_3838,N_3815);
xor U4027 (N_4027,N_3900,N_3977);
xnor U4028 (N_4028,N_3816,N_3980);
xnor U4029 (N_4029,N_3979,N_3935);
nor U4030 (N_4030,N_3960,N_3982);
nor U4031 (N_4031,N_3889,N_3885);
xor U4032 (N_4032,N_3943,N_3803);
nand U4033 (N_4033,N_3844,N_3894);
and U4034 (N_4034,N_3857,N_3951);
nor U4035 (N_4035,N_3909,N_3873);
or U4036 (N_4036,N_3967,N_3914);
or U4037 (N_4037,N_3969,N_3869);
or U4038 (N_4038,N_3938,N_3924);
nand U4039 (N_4039,N_3830,N_3877);
and U4040 (N_4040,N_3998,N_3975);
or U4041 (N_4041,N_3845,N_3834);
nand U4042 (N_4042,N_3811,N_3963);
nand U4043 (N_4043,N_3831,N_3859);
xnor U4044 (N_4044,N_3840,N_3855);
nor U4045 (N_4045,N_3984,N_3861);
nand U4046 (N_4046,N_3964,N_3867);
and U4047 (N_4047,N_3863,N_3945);
or U4048 (N_4048,N_3920,N_3871);
and U4049 (N_4049,N_3814,N_3961);
and U4050 (N_4050,N_3801,N_3865);
xnor U4051 (N_4051,N_3878,N_3875);
xor U4052 (N_4052,N_3817,N_3839);
nor U4053 (N_4053,N_3996,N_3849);
nand U4054 (N_4054,N_3930,N_3926);
nand U4055 (N_4055,N_3842,N_3866);
and U4056 (N_4056,N_3846,N_3882);
and U4057 (N_4057,N_3918,N_3800);
nor U4058 (N_4058,N_3962,N_3841);
and U4059 (N_4059,N_3852,N_3880);
xnor U4060 (N_4060,N_3804,N_3895);
and U4061 (N_4061,N_3911,N_3850);
nand U4062 (N_4062,N_3826,N_3901);
nor U4063 (N_4063,N_3910,N_3928);
or U4064 (N_4064,N_3987,N_3905);
nand U4065 (N_4065,N_3959,N_3947);
and U4066 (N_4066,N_3828,N_3908);
and U4067 (N_4067,N_3808,N_3981);
nand U4068 (N_4068,N_3966,N_3940);
xnor U4069 (N_4069,N_3922,N_3891);
xor U4070 (N_4070,N_3864,N_3912);
nand U4071 (N_4071,N_3993,N_3999);
nand U4072 (N_4072,N_3902,N_3936);
nor U4073 (N_4073,N_3915,N_3874);
nor U4074 (N_4074,N_3819,N_3812);
or U4075 (N_4075,N_3836,N_3818);
nor U4076 (N_4076,N_3917,N_3879);
nand U4077 (N_4077,N_3913,N_3985);
and U4078 (N_4078,N_3927,N_3941);
or U4079 (N_4079,N_3827,N_3921);
nor U4080 (N_4080,N_3823,N_3892);
or U4081 (N_4081,N_3853,N_3954);
or U4082 (N_4082,N_3810,N_3997);
nand U4083 (N_4083,N_3953,N_3806);
or U4084 (N_4084,N_3881,N_3868);
nor U4085 (N_4085,N_3907,N_3821);
xor U4086 (N_4086,N_3851,N_3860);
or U4087 (N_4087,N_3929,N_3957);
nor U4088 (N_4088,N_3994,N_3870);
and U4089 (N_4089,N_3835,N_3995);
nand U4090 (N_4090,N_3813,N_3956);
or U4091 (N_4091,N_3931,N_3822);
nand U4092 (N_4092,N_3972,N_3862);
nand U4093 (N_4093,N_3934,N_3903);
nor U4094 (N_4094,N_3946,N_3973);
nand U4095 (N_4095,N_3988,N_3858);
or U4096 (N_4096,N_3802,N_3824);
nand U4097 (N_4097,N_3955,N_3893);
nand U4098 (N_4098,N_3904,N_3970);
nor U4099 (N_4099,N_3923,N_3942);
or U4100 (N_4100,N_3926,N_3900);
or U4101 (N_4101,N_3850,N_3903);
xor U4102 (N_4102,N_3872,N_3997);
nand U4103 (N_4103,N_3943,N_3907);
nand U4104 (N_4104,N_3904,N_3943);
and U4105 (N_4105,N_3930,N_3946);
and U4106 (N_4106,N_3949,N_3913);
xnor U4107 (N_4107,N_3949,N_3882);
and U4108 (N_4108,N_3821,N_3810);
xor U4109 (N_4109,N_3902,N_3989);
nand U4110 (N_4110,N_3842,N_3893);
or U4111 (N_4111,N_3895,N_3968);
or U4112 (N_4112,N_3890,N_3989);
nor U4113 (N_4113,N_3981,N_3965);
or U4114 (N_4114,N_3995,N_3807);
or U4115 (N_4115,N_3962,N_3898);
and U4116 (N_4116,N_3929,N_3862);
nor U4117 (N_4117,N_3849,N_3883);
xnor U4118 (N_4118,N_3919,N_3966);
and U4119 (N_4119,N_3944,N_3936);
xnor U4120 (N_4120,N_3822,N_3833);
nand U4121 (N_4121,N_3993,N_3822);
nand U4122 (N_4122,N_3846,N_3820);
nand U4123 (N_4123,N_3839,N_3841);
nor U4124 (N_4124,N_3903,N_3932);
xnor U4125 (N_4125,N_3820,N_3884);
or U4126 (N_4126,N_3848,N_3947);
xor U4127 (N_4127,N_3815,N_3851);
nand U4128 (N_4128,N_3817,N_3829);
and U4129 (N_4129,N_3802,N_3972);
nor U4130 (N_4130,N_3976,N_3868);
or U4131 (N_4131,N_3826,N_3892);
nor U4132 (N_4132,N_3979,N_3973);
nand U4133 (N_4133,N_3870,N_3840);
nor U4134 (N_4134,N_3914,N_3862);
or U4135 (N_4135,N_3872,N_3946);
or U4136 (N_4136,N_3849,N_3928);
or U4137 (N_4137,N_3925,N_3872);
nand U4138 (N_4138,N_3888,N_3816);
nand U4139 (N_4139,N_3880,N_3928);
xnor U4140 (N_4140,N_3815,N_3924);
xor U4141 (N_4141,N_3992,N_3872);
or U4142 (N_4142,N_3807,N_3921);
and U4143 (N_4143,N_3823,N_3806);
or U4144 (N_4144,N_3832,N_3985);
xor U4145 (N_4145,N_3930,N_3832);
nor U4146 (N_4146,N_3902,N_3892);
nor U4147 (N_4147,N_3862,N_3892);
or U4148 (N_4148,N_3902,N_3826);
nor U4149 (N_4149,N_3834,N_3901);
or U4150 (N_4150,N_3948,N_3851);
and U4151 (N_4151,N_3931,N_3836);
nor U4152 (N_4152,N_3988,N_3931);
nand U4153 (N_4153,N_3884,N_3870);
xor U4154 (N_4154,N_3977,N_3810);
nand U4155 (N_4155,N_3966,N_3971);
and U4156 (N_4156,N_3905,N_3975);
and U4157 (N_4157,N_3893,N_3911);
and U4158 (N_4158,N_3961,N_3842);
and U4159 (N_4159,N_3817,N_3889);
xor U4160 (N_4160,N_3921,N_3987);
or U4161 (N_4161,N_3826,N_3875);
and U4162 (N_4162,N_3983,N_3867);
nand U4163 (N_4163,N_3966,N_3922);
and U4164 (N_4164,N_3853,N_3811);
or U4165 (N_4165,N_3821,N_3898);
nand U4166 (N_4166,N_3805,N_3954);
xor U4167 (N_4167,N_3992,N_3987);
nand U4168 (N_4168,N_3805,N_3865);
and U4169 (N_4169,N_3857,N_3890);
nor U4170 (N_4170,N_3872,N_3918);
nand U4171 (N_4171,N_3956,N_3957);
xor U4172 (N_4172,N_3939,N_3813);
nor U4173 (N_4173,N_3990,N_3959);
nor U4174 (N_4174,N_3846,N_3934);
xor U4175 (N_4175,N_3940,N_3848);
or U4176 (N_4176,N_3834,N_3800);
and U4177 (N_4177,N_3862,N_3881);
nand U4178 (N_4178,N_3997,N_3913);
nand U4179 (N_4179,N_3905,N_3921);
xnor U4180 (N_4180,N_3847,N_3800);
nand U4181 (N_4181,N_3814,N_3866);
nand U4182 (N_4182,N_3992,N_3900);
or U4183 (N_4183,N_3903,N_3920);
nand U4184 (N_4184,N_3910,N_3941);
or U4185 (N_4185,N_3867,N_3961);
xor U4186 (N_4186,N_3835,N_3837);
xor U4187 (N_4187,N_3996,N_3827);
and U4188 (N_4188,N_3910,N_3944);
xnor U4189 (N_4189,N_3890,N_3804);
or U4190 (N_4190,N_3955,N_3862);
xor U4191 (N_4191,N_3931,N_3968);
nand U4192 (N_4192,N_3909,N_3811);
nand U4193 (N_4193,N_3915,N_3919);
and U4194 (N_4194,N_3993,N_3989);
nand U4195 (N_4195,N_3905,N_3871);
or U4196 (N_4196,N_3941,N_3935);
and U4197 (N_4197,N_3952,N_3869);
or U4198 (N_4198,N_3962,N_3953);
nand U4199 (N_4199,N_3970,N_3991);
nand U4200 (N_4200,N_4183,N_4105);
and U4201 (N_4201,N_4008,N_4065);
nor U4202 (N_4202,N_4102,N_4019);
and U4203 (N_4203,N_4029,N_4042);
and U4204 (N_4204,N_4161,N_4158);
nor U4205 (N_4205,N_4049,N_4088);
nand U4206 (N_4206,N_4156,N_4140);
nor U4207 (N_4207,N_4083,N_4166);
and U4208 (N_4208,N_4092,N_4177);
and U4209 (N_4209,N_4135,N_4068);
nor U4210 (N_4210,N_4142,N_4016);
nand U4211 (N_4211,N_4101,N_4027);
and U4212 (N_4212,N_4072,N_4132);
and U4213 (N_4213,N_4084,N_4117);
nor U4214 (N_4214,N_4162,N_4089);
and U4215 (N_4215,N_4178,N_4009);
nand U4216 (N_4216,N_4044,N_4024);
xor U4217 (N_4217,N_4122,N_4022);
xnor U4218 (N_4218,N_4062,N_4059);
nor U4219 (N_4219,N_4074,N_4136);
or U4220 (N_4220,N_4041,N_4104);
nor U4221 (N_4221,N_4113,N_4037);
nand U4222 (N_4222,N_4121,N_4096);
nor U4223 (N_4223,N_4118,N_4171);
and U4224 (N_4224,N_4036,N_4130);
and U4225 (N_4225,N_4047,N_4091);
and U4226 (N_4226,N_4197,N_4126);
nor U4227 (N_4227,N_4198,N_4189);
nand U4228 (N_4228,N_4040,N_4128);
nand U4229 (N_4229,N_4039,N_4034);
and U4230 (N_4230,N_4075,N_4160);
nand U4231 (N_4231,N_4149,N_4120);
xnor U4232 (N_4232,N_4069,N_4058);
or U4233 (N_4233,N_4098,N_4015);
nand U4234 (N_4234,N_4119,N_4152);
and U4235 (N_4235,N_4137,N_4107);
or U4236 (N_4236,N_4014,N_4030);
and U4237 (N_4237,N_4176,N_4153);
or U4238 (N_4238,N_4077,N_4060);
or U4239 (N_4239,N_4129,N_4080);
nand U4240 (N_4240,N_4070,N_4038);
nor U4241 (N_4241,N_4085,N_4017);
xor U4242 (N_4242,N_4081,N_4163);
or U4243 (N_4243,N_4146,N_4103);
xor U4244 (N_4244,N_4054,N_4064);
and U4245 (N_4245,N_4108,N_4097);
and U4246 (N_4246,N_4031,N_4006);
nor U4247 (N_4247,N_4011,N_4199);
and U4248 (N_4248,N_4071,N_4168);
nand U4249 (N_4249,N_4051,N_4001);
nor U4250 (N_4250,N_4182,N_4195);
nand U4251 (N_4251,N_4180,N_4141);
nor U4252 (N_4252,N_4112,N_4094);
nor U4253 (N_4253,N_4086,N_4013);
or U4254 (N_4254,N_4133,N_4110);
xnor U4255 (N_4255,N_4061,N_4190);
and U4256 (N_4256,N_4063,N_4123);
and U4257 (N_4257,N_4193,N_4045);
and U4258 (N_4258,N_4115,N_4002);
or U4259 (N_4259,N_4020,N_4018);
nor U4260 (N_4260,N_4100,N_4185);
or U4261 (N_4261,N_4157,N_4090);
or U4262 (N_4262,N_4124,N_4078);
nor U4263 (N_4263,N_4188,N_4150);
nand U4264 (N_4264,N_4032,N_4134);
or U4265 (N_4265,N_4007,N_4154);
nand U4266 (N_4266,N_4026,N_4170);
nand U4267 (N_4267,N_4093,N_4046);
or U4268 (N_4268,N_4165,N_4173);
nor U4269 (N_4269,N_4151,N_4194);
and U4270 (N_4270,N_4184,N_4053);
nand U4271 (N_4271,N_4196,N_4004);
nor U4272 (N_4272,N_4192,N_4079);
and U4273 (N_4273,N_4159,N_4010);
nor U4274 (N_4274,N_4067,N_4003);
xor U4275 (N_4275,N_4138,N_4033);
nand U4276 (N_4276,N_4076,N_4035);
and U4277 (N_4277,N_4021,N_4175);
and U4278 (N_4278,N_4169,N_4174);
and U4279 (N_4279,N_4111,N_4172);
xnor U4280 (N_4280,N_4147,N_4082);
nand U4281 (N_4281,N_4028,N_4116);
nand U4282 (N_4282,N_4114,N_4164);
and U4283 (N_4283,N_4073,N_4145);
nor U4284 (N_4284,N_4052,N_4005);
nor U4285 (N_4285,N_4179,N_4109);
and U4286 (N_4286,N_4095,N_4087);
and U4287 (N_4287,N_4055,N_4143);
xnor U4288 (N_4288,N_4186,N_4099);
nand U4289 (N_4289,N_4023,N_4125);
or U4290 (N_4290,N_4043,N_4066);
or U4291 (N_4291,N_4057,N_4148);
nand U4292 (N_4292,N_4131,N_4191);
xnor U4293 (N_4293,N_4181,N_4139);
nand U4294 (N_4294,N_4106,N_4048);
xor U4295 (N_4295,N_4155,N_4187);
and U4296 (N_4296,N_4127,N_4144);
and U4297 (N_4297,N_4050,N_4012);
xnor U4298 (N_4298,N_4056,N_4000);
or U4299 (N_4299,N_4167,N_4025);
and U4300 (N_4300,N_4002,N_4091);
nor U4301 (N_4301,N_4155,N_4056);
nand U4302 (N_4302,N_4148,N_4001);
or U4303 (N_4303,N_4141,N_4002);
xor U4304 (N_4304,N_4006,N_4137);
nand U4305 (N_4305,N_4105,N_4161);
nand U4306 (N_4306,N_4106,N_4054);
nand U4307 (N_4307,N_4124,N_4180);
and U4308 (N_4308,N_4170,N_4147);
and U4309 (N_4309,N_4022,N_4000);
or U4310 (N_4310,N_4163,N_4067);
and U4311 (N_4311,N_4119,N_4148);
nand U4312 (N_4312,N_4169,N_4075);
nand U4313 (N_4313,N_4166,N_4122);
and U4314 (N_4314,N_4091,N_4133);
or U4315 (N_4315,N_4135,N_4102);
or U4316 (N_4316,N_4120,N_4039);
or U4317 (N_4317,N_4185,N_4020);
and U4318 (N_4318,N_4193,N_4059);
nand U4319 (N_4319,N_4078,N_4055);
nor U4320 (N_4320,N_4098,N_4007);
or U4321 (N_4321,N_4094,N_4110);
and U4322 (N_4322,N_4004,N_4018);
and U4323 (N_4323,N_4009,N_4095);
xnor U4324 (N_4324,N_4125,N_4097);
nor U4325 (N_4325,N_4113,N_4127);
or U4326 (N_4326,N_4167,N_4024);
xor U4327 (N_4327,N_4028,N_4097);
or U4328 (N_4328,N_4030,N_4085);
or U4329 (N_4329,N_4072,N_4047);
and U4330 (N_4330,N_4074,N_4058);
and U4331 (N_4331,N_4119,N_4150);
xnor U4332 (N_4332,N_4024,N_4036);
xor U4333 (N_4333,N_4106,N_4131);
or U4334 (N_4334,N_4102,N_4054);
nand U4335 (N_4335,N_4120,N_4115);
nor U4336 (N_4336,N_4013,N_4043);
nor U4337 (N_4337,N_4022,N_4183);
and U4338 (N_4338,N_4096,N_4067);
xnor U4339 (N_4339,N_4145,N_4120);
nor U4340 (N_4340,N_4177,N_4034);
and U4341 (N_4341,N_4183,N_4033);
nor U4342 (N_4342,N_4087,N_4062);
nor U4343 (N_4343,N_4126,N_4082);
and U4344 (N_4344,N_4128,N_4063);
nand U4345 (N_4345,N_4168,N_4183);
and U4346 (N_4346,N_4145,N_4198);
xor U4347 (N_4347,N_4121,N_4054);
nor U4348 (N_4348,N_4126,N_4015);
nor U4349 (N_4349,N_4067,N_4071);
and U4350 (N_4350,N_4198,N_4006);
and U4351 (N_4351,N_4112,N_4068);
or U4352 (N_4352,N_4192,N_4016);
xnor U4353 (N_4353,N_4060,N_4170);
nor U4354 (N_4354,N_4171,N_4043);
xor U4355 (N_4355,N_4116,N_4072);
or U4356 (N_4356,N_4017,N_4003);
nand U4357 (N_4357,N_4074,N_4146);
or U4358 (N_4358,N_4067,N_4196);
nor U4359 (N_4359,N_4123,N_4034);
and U4360 (N_4360,N_4130,N_4081);
and U4361 (N_4361,N_4013,N_4049);
and U4362 (N_4362,N_4052,N_4163);
nand U4363 (N_4363,N_4074,N_4109);
nand U4364 (N_4364,N_4175,N_4131);
xor U4365 (N_4365,N_4117,N_4106);
nand U4366 (N_4366,N_4056,N_4145);
or U4367 (N_4367,N_4008,N_4051);
or U4368 (N_4368,N_4056,N_4094);
nor U4369 (N_4369,N_4029,N_4197);
nor U4370 (N_4370,N_4008,N_4178);
nand U4371 (N_4371,N_4152,N_4093);
xor U4372 (N_4372,N_4139,N_4131);
nand U4373 (N_4373,N_4192,N_4082);
xnor U4374 (N_4374,N_4131,N_4019);
xnor U4375 (N_4375,N_4061,N_4157);
xor U4376 (N_4376,N_4125,N_4079);
or U4377 (N_4377,N_4113,N_4074);
nand U4378 (N_4378,N_4047,N_4156);
nor U4379 (N_4379,N_4134,N_4147);
or U4380 (N_4380,N_4076,N_4043);
nand U4381 (N_4381,N_4046,N_4107);
and U4382 (N_4382,N_4051,N_4150);
nor U4383 (N_4383,N_4033,N_4148);
xnor U4384 (N_4384,N_4190,N_4157);
and U4385 (N_4385,N_4146,N_4038);
nand U4386 (N_4386,N_4118,N_4129);
and U4387 (N_4387,N_4030,N_4189);
nand U4388 (N_4388,N_4196,N_4049);
nor U4389 (N_4389,N_4045,N_4070);
nand U4390 (N_4390,N_4080,N_4005);
nand U4391 (N_4391,N_4005,N_4143);
nand U4392 (N_4392,N_4055,N_4131);
nand U4393 (N_4393,N_4071,N_4149);
nand U4394 (N_4394,N_4184,N_4034);
and U4395 (N_4395,N_4076,N_4154);
nor U4396 (N_4396,N_4101,N_4054);
or U4397 (N_4397,N_4080,N_4058);
and U4398 (N_4398,N_4042,N_4057);
nand U4399 (N_4399,N_4109,N_4166);
or U4400 (N_4400,N_4291,N_4316);
nand U4401 (N_4401,N_4230,N_4365);
or U4402 (N_4402,N_4278,N_4341);
nand U4403 (N_4403,N_4363,N_4358);
and U4404 (N_4404,N_4205,N_4368);
nor U4405 (N_4405,N_4269,N_4227);
and U4406 (N_4406,N_4236,N_4399);
nor U4407 (N_4407,N_4301,N_4279);
xor U4408 (N_4408,N_4287,N_4307);
nand U4409 (N_4409,N_4334,N_4203);
xnor U4410 (N_4410,N_4394,N_4296);
nor U4411 (N_4411,N_4367,N_4293);
nand U4412 (N_4412,N_4209,N_4309);
nand U4413 (N_4413,N_4322,N_4201);
and U4414 (N_4414,N_4229,N_4328);
nand U4415 (N_4415,N_4366,N_4225);
xor U4416 (N_4416,N_4349,N_4338);
nor U4417 (N_4417,N_4221,N_4352);
or U4418 (N_4418,N_4331,N_4396);
xnor U4419 (N_4419,N_4387,N_4350);
nand U4420 (N_4420,N_4343,N_4323);
nand U4421 (N_4421,N_4379,N_4335);
xor U4422 (N_4422,N_4284,N_4295);
xnor U4423 (N_4423,N_4255,N_4235);
nand U4424 (N_4424,N_4391,N_4330);
nand U4425 (N_4425,N_4377,N_4243);
or U4426 (N_4426,N_4212,N_4257);
nand U4427 (N_4427,N_4305,N_4283);
nand U4428 (N_4428,N_4364,N_4310);
nand U4429 (N_4429,N_4226,N_4324);
or U4430 (N_4430,N_4300,N_4206);
or U4431 (N_4431,N_4228,N_4261);
nand U4432 (N_4432,N_4329,N_4355);
and U4433 (N_4433,N_4250,N_4319);
nand U4434 (N_4434,N_4266,N_4360);
xnor U4435 (N_4435,N_4382,N_4248);
or U4436 (N_4436,N_4288,N_4372);
or U4437 (N_4437,N_4302,N_4265);
xnor U4438 (N_4438,N_4327,N_4304);
nor U4439 (N_4439,N_4217,N_4274);
or U4440 (N_4440,N_4380,N_4325);
nand U4441 (N_4441,N_4306,N_4345);
nand U4442 (N_4442,N_4247,N_4245);
or U4443 (N_4443,N_4240,N_4336);
nand U4444 (N_4444,N_4390,N_4200);
nand U4445 (N_4445,N_4219,N_4220);
nand U4446 (N_4446,N_4348,N_4214);
nand U4447 (N_4447,N_4210,N_4342);
nor U4448 (N_4448,N_4373,N_4246);
nand U4449 (N_4449,N_4359,N_4356);
or U4450 (N_4450,N_4260,N_4393);
nand U4451 (N_4451,N_4320,N_4285);
and U4452 (N_4452,N_4299,N_4292);
nor U4453 (N_4453,N_4369,N_4276);
or U4454 (N_4454,N_4262,N_4244);
and U4455 (N_4455,N_4381,N_4361);
nand U4456 (N_4456,N_4384,N_4242);
nor U4457 (N_4457,N_4339,N_4234);
nand U4458 (N_4458,N_4268,N_4254);
nand U4459 (N_4459,N_4233,N_4282);
and U4460 (N_4460,N_4264,N_4267);
nor U4461 (N_4461,N_4202,N_4375);
nand U4462 (N_4462,N_4371,N_4232);
xnor U4463 (N_4463,N_4303,N_4340);
or U4464 (N_4464,N_4223,N_4294);
xor U4465 (N_4465,N_4318,N_4256);
nand U4466 (N_4466,N_4351,N_4277);
or U4467 (N_4467,N_4290,N_4337);
or U4468 (N_4468,N_4353,N_4374);
xnor U4469 (N_4469,N_4392,N_4272);
nor U4470 (N_4470,N_4326,N_4241);
nand U4471 (N_4471,N_4204,N_4386);
and U4472 (N_4472,N_4286,N_4270);
and U4473 (N_4473,N_4346,N_4252);
xnor U4474 (N_4474,N_4333,N_4280);
nor U4475 (N_4475,N_4208,N_4397);
or U4476 (N_4476,N_4395,N_4357);
nand U4477 (N_4477,N_4213,N_4224);
xor U4478 (N_4478,N_4311,N_4332);
and U4479 (N_4479,N_4275,N_4238);
and U4480 (N_4480,N_4385,N_4388);
nand U4481 (N_4481,N_4258,N_4347);
or U4482 (N_4482,N_4315,N_4211);
nand U4483 (N_4483,N_4362,N_4271);
xnor U4484 (N_4484,N_4289,N_4259);
nand U4485 (N_4485,N_4222,N_4249);
and U4486 (N_4486,N_4207,N_4383);
nand U4487 (N_4487,N_4370,N_4321);
xor U4488 (N_4488,N_4297,N_4398);
nor U4489 (N_4489,N_4239,N_4215);
nand U4490 (N_4490,N_4298,N_4313);
nand U4491 (N_4491,N_4376,N_4253);
and U4492 (N_4492,N_4314,N_4237);
and U4493 (N_4493,N_4281,N_4273);
nand U4494 (N_4494,N_4389,N_4231);
nand U4495 (N_4495,N_4344,N_4216);
nand U4496 (N_4496,N_4312,N_4308);
and U4497 (N_4497,N_4218,N_4354);
nand U4498 (N_4498,N_4251,N_4378);
xnor U4499 (N_4499,N_4317,N_4263);
nor U4500 (N_4500,N_4204,N_4264);
and U4501 (N_4501,N_4284,N_4298);
nor U4502 (N_4502,N_4345,N_4399);
xor U4503 (N_4503,N_4214,N_4368);
xnor U4504 (N_4504,N_4381,N_4352);
nand U4505 (N_4505,N_4224,N_4327);
and U4506 (N_4506,N_4201,N_4280);
xor U4507 (N_4507,N_4239,N_4399);
and U4508 (N_4508,N_4232,N_4356);
nand U4509 (N_4509,N_4213,N_4274);
nor U4510 (N_4510,N_4388,N_4380);
or U4511 (N_4511,N_4323,N_4213);
nor U4512 (N_4512,N_4263,N_4278);
nor U4513 (N_4513,N_4398,N_4253);
xnor U4514 (N_4514,N_4251,N_4283);
xor U4515 (N_4515,N_4273,N_4251);
nand U4516 (N_4516,N_4361,N_4326);
or U4517 (N_4517,N_4311,N_4276);
xnor U4518 (N_4518,N_4383,N_4387);
xnor U4519 (N_4519,N_4388,N_4313);
nor U4520 (N_4520,N_4347,N_4208);
nor U4521 (N_4521,N_4267,N_4339);
xor U4522 (N_4522,N_4359,N_4332);
nand U4523 (N_4523,N_4294,N_4278);
nor U4524 (N_4524,N_4328,N_4204);
nand U4525 (N_4525,N_4317,N_4200);
or U4526 (N_4526,N_4259,N_4363);
nor U4527 (N_4527,N_4326,N_4296);
nand U4528 (N_4528,N_4308,N_4294);
nor U4529 (N_4529,N_4314,N_4260);
nor U4530 (N_4530,N_4204,N_4380);
xor U4531 (N_4531,N_4298,N_4373);
and U4532 (N_4532,N_4261,N_4207);
nor U4533 (N_4533,N_4390,N_4241);
nand U4534 (N_4534,N_4324,N_4234);
nor U4535 (N_4535,N_4267,N_4273);
or U4536 (N_4536,N_4333,N_4367);
nor U4537 (N_4537,N_4355,N_4381);
or U4538 (N_4538,N_4252,N_4272);
or U4539 (N_4539,N_4356,N_4222);
nand U4540 (N_4540,N_4246,N_4297);
nor U4541 (N_4541,N_4348,N_4351);
nor U4542 (N_4542,N_4234,N_4210);
and U4543 (N_4543,N_4369,N_4213);
or U4544 (N_4544,N_4221,N_4339);
xor U4545 (N_4545,N_4257,N_4273);
xor U4546 (N_4546,N_4261,N_4265);
nor U4547 (N_4547,N_4267,N_4305);
or U4548 (N_4548,N_4309,N_4296);
nand U4549 (N_4549,N_4269,N_4211);
nor U4550 (N_4550,N_4257,N_4326);
and U4551 (N_4551,N_4334,N_4227);
and U4552 (N_4552,N_4218,N_4387);
nor U4553 (N_4553,N_4274,N_4209);
nor U4554 (N_4554,N_4323,N_4206);
nand U4555 (N_4555,N_4310,N_4339);
xnor U4556 (N_4556,N_4345,N_4286);
and U4557 (N_4557,N_4207,N_4279);
nand U4558 (N_4558,N_4284,N_4291);
nor U4559 (N_4559,N_4357,N_4378);
nand U4560 (N_4560,N_4243,N_4281);
nor U4561 (N_4561,N_4361,N_4207);
and U4562 (N_4562,N_4336,N_4304);
nand U4563 (N_4563,N_4383,N_4258);
nand U4564 (N_4564,N_4228,N_4225);
nor U4565 (N_4565,N_4316,N_4383);
xnor U4566 (N_4566,N_4398,N_4317);
nand U4567 (N_4567,N_4220,N_4265);
nand U4568 (N_4568,N_4273,N_4208);
and U4569 (N_4569,N_4296,N_4365);
or U4570 (N_4570,N_4233,N_4315);
and U4571 (N_4571,N_4369,N_4321);
and U4572 (N_4572,N_4371,N_4261);
xnor U4573 (N_4573,N_4376,N_4252);
xnor U4574 (N_4574,N_4343,N_4221);
xnor U4575 (N_4575,N_4347,N_4308);
nand U4576 (N_4576,N_4375,N_4281);
nor U4577 (N_4577,N_4225,N_4399);
xor U4578 (N_4578,N_4382,N_4201);
nor U4579 (N_4579,N_4394,N_4330);
nand U4580 (N_4580,N_4234,N_4341);
xnor U4581 (N_4581,N_4200,N_4311);
nand U4582 (N_4582,N_4248,N_4268);
nor U4583 (N_4583,N_4350,N_4389);
or U4584 (N_4584,N_4347,N_4273);
or U4585 (N_4585,N_4367,N_4290);
and U4586 (N_4586,N_4256,N_4210);
and U4587 (N_4587,N_4273,N_4234);
or U4588 (N_4588,N_4387,N_4271);
xnor U4589 (N_4589,N_4267,N_4376);
and U4590 (N_4590,N_4227,N_4354);
nand U4591 (N_4591,N_4242,N_4320);
xor U4592 (N_4592,N_4339,N_4270);
xnor U4593 (N_4593,N_4393,N_4293);
nor U4594 (N_4594,N_4371,N_4272);
or U4595 (N_4595,N_4200,N_4315);
nand U4596 (N_4596,N_4261,N_4210);
xor U4597 (N_4597,N_4381,N_4262);
nand U4598 (N_4598,N_4238,N_4202);
or U4599 (N_4599,N_4219,N_4332);
or U4600 (N_4600,N_4508,N_4455);
and U4601 (N_4601,N_4478,N_4504);
or U4602 (N_4602,N_4497,N_4511);
nor U4603 (N_4603,N_4551,N_4586);
nor U4604 (N_4604,N_4408,N_4481);
or U4605 (N_4605,N_4470,N_4419);
or U4606 (N_4606,N_4598,N_4593);
nor U4607 (N_4607,N_4479,N_4487);
and U4608 (N_4608,N_4403,N_4447);
and U4609 (N_4609,N_4444,N_4473);
nand U4610 (N_4610,N_4416,N_4463);
nand U4611 (N_4611,N_4579,N_4472);
or U4612 (N_4612,N_4407,N_4568);
nor U4613 (N_4613,N_4558,N_4476);
xor U4614 (N_4614,N_4599,N_4486);
nand U4615 (N_4615,N_4522,N_4505);
and U4616 (N_4616,N_4450,N_4523);
xnor U4617 (N_4617,N_4437,N_4510);
and U4618 (N_4618,N_4443,N_4424);
or U4619 (N_4619,N_4496,N_4545);
and U4620 (N_4620,N_4432,N_4411);
and U4621 (N_4621,N_4596,N_4552);
xor U4622 (N_4622,N_4571,N_4536);
nand U4623 (N_4623,N_4595,N_4493);
nor U4624 (N_4624,N_4445,N_4557);
or U4625 (N_4625,N_4588,N_4454);
nand U4626 (N_4626,N_4576,N_4560);
and U4627 (N_4627,N_4495,N_4405);
nand U4628 (N_4628,N_4442,N_4460);
or U4629 (N_4629,N_4426,N_4499);
nor U4630 (N_4630,N_4529,N_4439);
nand U4631 (N_4631,N_4452,N_4448);
or U4632 (N_4632,N_4457,N_4489);
xnor U4633 (N_4633,N_4500,N_4467);
nand U4634 (N_4634,N_4412,N_4513);
nor U4635 (N_4635,N_4570,N_4514);
nand U4636 (N_4636,N_4532,N_4546);
nor U4637 (N_4637,N_4469,N_4485);
and U4638 (N_4638,N_4429,N_4582);
nor U4639 (N_4639,N_4440,N_4520);
xor U4640 (N_4640,N_4578,N_4526);
and U4641 (N_4641,N_4466,N_4528);
xor U4642 (N_4642,N_4561,N_4451);
nor U4643 (N_4643,N_4559,N_4482);
and U4644 (N_4644,N_4527,N_4550);
nand U4645 (N_4645,N_4516,N_4406);
nor U4646 (N_4646,N_4543,N_4572);
nor U4647 (N_4647,N_4471,N_4542);
and U4648 (N_4648,N_4584,N_4464);
and U4649 (N_4649,N_4427,N_4446);
and U4650 (N_4650,N_4512,N_4556);
xor U4651 (N_4651,N_4502,N_4468);
xnor U4652 (N_4652,N_4539,N_4554);
nor U4653 (N_4653,N_4400,N_4569);
and U4654 (N_4654,N_4541,N_4458);
and U4655 (N_4655,N_4515,N_4538);
or U4656 (N_4656,N_4567,N_4591);
or U4657 (N_4657,N_4453,N_4535);
nand U4658 (N_4658,N_4435,N_4404);
nand U4659 (N_4659,N_4597,N_4413);
xnor U4660 (N_4660,N_4492,N_4540);
and U4661 (N_4661,N_4480,N_4438);
and U4662 (N_4662,N_4401,N_4580);
nor U4663 (N_4663,N_4488,N_4533);
and U4664 (N_4664,N_4420,N_4402);
or U4665 (N_4665,N_4433,N_4577);
xnor U4666 (N_4666,N_4421,N_4575);
nor U4667 (N_4667,N_4415,N_4537);
nor U4668 (N_4668,N_4410,N_4428);
nor U4669 (N_4669,N_4507,N_4518);
nor U4670 (N_4670,N_4549,N_4587);
nand U4671 (N_4671,N_4491,N_4498);
nand U4672 (N_4672,N_4553,N_4494);
nor U4673 (N_4673,N_4521,N_4436);
or U4674 (N_4674,N_4434,N_4563);
nand U4675 (N_4675,N_4585,N_4484);
nor U4676 (N_4676,N_4509,N_4565);
nand U4677 (N_4677,N_4564,N_4462);
nand U4678 (N_4678,N_4501,N_4506);
nor U4679 (N_4679,N_4566,N_4459);
and U4680 (N_4680,N_4441,N_4519);
nor U4681 (N_4681,N_4456,N_4423);
or U4682 (N_4682,N_4525,N_4461);
nor U4683 (N_4683,N_4581,N_4594);
nor U4684 (N_4684,N_4490,N_4418);
nand U4685 (N_4685,N_4555,N_4562);
and U4686 (N_4686,N_4465,N_4548);
or U4687 (N_4687,N_4449,N_4573);
or U4688 (N_4688,N_4544,N_4590);
nor U4689 (N_4689,N_4574,N_4414);
nor U4690 (N_4690,N_4534,N_4592);
nor U4691 (N_4691,N_4417,N_4583);
or U4692 (N_4692,N_4474,N_4517);
or U4693 (N_4693,N_4409,N_4589);
or U4694 (N_4694,N_4477,N_4483);
xnor U4695 (N_4695,N_4547,N_4431);
xor U4696 (N_4696,N_4422,N_4531);
nor U4697 (N_4697,N_4503,N_4430);
or U4698 (N_4698,N_4475,N_4524);
and U4699 (N_4699,N_4530,N_4425);
nand U4700 (N_4700,N_4510,N_4454);
xor U4701 (N_4701,N_4412,N_4598);
nor U4702 (N_4702,N_4479,N_4491);
or U4703 (N_4703,N_4413,N_4523);
and U4704 (N_4704,N_4428,N_4407);
or U4705 (N_4705,N_4495,N_4419);
and U4706 (N_4706,N_4482,N_4424);
or U4707 (N_4707,N_4595,N_4407);
or U4708 (N_4708,N_4495,N_4408);
nor U4709 (N_4709,N_4561,N_4567);
nor U4710 (N_4710,N_4530,N_4477);
or U4711 (N_4711,N_4598,N_4462);
nor U4712 (N_4712,N_4541,N_4402);
or U4713 (N_4713,N_4490,N_4458);
and U4714 (N_4714,N_4491,N_4567);
nor U4715 (N_4715,N_4589,N_4441);
xor U4716 (N_4716,N_4574,N_4425);
xnor U4717 (N_4717,N_4440,N_4498);
xnor U4718 (N_4718,N_4574,N_4534);
or U4719 (N_4719,N_4404,N_4594);
or U4720 (N_4720,N_4401,N_4533);
or U4721 (N_4721,N_4430,N_4438);
nor U4722 (N_4722,N_4598,N_4449);
xnor U4723 (N_4723,N_4423,N_4448);
or U4724 (N_4724,N_4414,N_4433);
xnor U4725 (N_4725,N_4466,N_4536);
nor U4726 (N_4726,N_4489,N_4596);
nor U4727 (N_4727,N_4437,N_4467);
or U4728 (N_4728,N_4574,N_4508);
and U4729 (N_4729,N_4589,N_4508);
xor U4730 (N_4730,N_4418,N_4454);
or U4731 (N_4731,N_4458,N_4590);
xor U4732 (N_4732,N_4528,N_4456);
nand U4733 (N_4733,N_4435,N_4580);
nand U4734 (N_4734,N_4560,N_4566);
nor U4735 (N_4735,N_4472,N_4573);
or U4736 (N_4736,N_4505,N_4516);
and U4737 (N_4737,N_4412,N_4481);
nor U4738 (N_4738,N_4475,N_4468);
nor U4739 (N_4739,N_4574,N_4457);
nand U4740 (N_4740,N_4457,N_4444);
or U4741 (N_4741,N_4437,N_4503);
nor U4742 (N_4742,N_4513,N_4536);
and U4743 (N_4743,N_4538,N_4483);
nor U4744 (N_4744,N_4563,N_4475);
nor U4745 (N_4745,N_4596,N_4590);
nand U4746 (N_4746,N_4466,N_4488);
or U4747 (N_4747,N_4559,N_4562);
or U4748 (N_4748,N_4503,N_4553);
nand U4749 (N_4749,N_4574,N_4579);
or U4750 (N_4750,N_4437,N_4562);
xor U4751 (N_4751,N_4476,N_4522);
nor U4752 (N_4752,N_4544,N_4503);
nand U4753 (N_4753,N_4467,N_4596);
xor U4754 (N_4754,N_4527,N_4400);
xnor U4755 (N_4755,N_4481,N_4585);
and U4756 (N_4756,N_4504,N_4526);
nand U4757 (N_4757,N_4422,N_4467);
xor U4758 (N_4758,N_4534,N_4484);
nand U4759 (N_4759,N_4442,N_4578);
nand U4760 (N_4760,N_4508,N_4483);
xnor U4761 (N_4761,N_4468,N_4408);
or U4762 (N_4762,N_4544,N_4555);
nand U4763 (N_4763,N_4525,N_4427);
nand U4764 (N_4764,N_4489,N_4458);
nor U4765 (N_4765,N_4404,N_4419);
nor U4766 (N_4766,N_4578,N_4418);
nand U4767 (N_4767,N_4446,N_4426);
xnor U4768 (N_4768,N_4537,N_4571);
and U4769 (N_4769,N_4432,N_4554);
nand U4770 (N_4770,N_4563,N_4449);
or U4771 (N_4771,N_4541,N_4573);
nand U4772 (N_4772,N_4562,N_4445);
xor U4773 (N_4773,N_4561,N_4464);
nor U4774 (N_4774,N_4565,N_4581);
xnor U4775 (N_4775,N_4565,N_4556);
or U4776 (N_4776,N_4529,N_4411);
xnor U4777 (N_4777,N_4466,N_4527);
xnor U4778 (N_4778,N_4453,N_4503);
xnor U4779 (N_4779,N_4560,N_4411);
xnor U4780 (N_4780,N_4484,N_4569);
nor U4781 (N_4781,N_4466,N_4496);
nand U4782 (N_4782,N_4520,N_4542);
nand U4783 (N_4783,N_4498,N_4444);
nor U4784 (N_4784,N_4590,N_4465);
or U4785 (N_4785,N_4427,N_4487);
or U4786 (N_4786,N_4535,N_4523);
xnor U4787 (N_4787,N_4418,N_4453);
xnor U4788 (N_4788,N_4537,N_4568);
or U4789 (N_4789,N_4574,N_4442);
xor U4790 (N_4790,N_4429,N_4514);
xor U4791 (N_4791,N_4462,N_4482);
or U4792 (N_4792,N_4426,N_4506);
nand U4793 (N_4793,N_4442,N_4414);
xnor U4794 (N_4794,N_4492,N_4487);
nand U4795 (N_4795,N_4571,N_4544);
nor U4796 (N_4796,N_4470,N_4547);
nor U4797 (N_4797,N_4523,N_4568);
or U4798 (N_4798,N_4435,N_4590);
and U4799 (N_4799,N_4425,N_4583);
nor U4800 (N_4800,N_4637,N_4709);
nand U4801 (N_4801,N_4766,N_4729);
nor U4802 (N_4802,N_4621,N_4797);
nor U4803 (N_4803,N_4792,N_4755);
and U4804 (N_4804,N_4635,N_4751);
or U4805 (N_4805,N_4644,N_4604);
nor U4806 (N_4806,N_4638,N_4676);
xor U4807 (N_4807,N_4671,N_4752);
and U4808 (N_4808,N_4688,N_4723);
nand U4809 (N_4809,N_4682,N_4666);
and U4810 (N_4810,N_4720,N_4603);
or U4811 (N_4811,N_4663,N_4767);
nand U4812 (N_4812,N_4626,N_4754);
nor U4813 (N_4813,N_4707,N_4774);
xnor U4814 (N_4814,N_4669,N_4656);
and U4815 (N_4815,N_4794,N_4736);
nand U4816 (N_4816,N_4672,N_4629);
or U4817 (N_4817,N_4654,N_4619);
nand U4818 (N_4818,N_4616,N_4703);
nor U4819 (N_4819,N_4612,N_4643);
nand U4820 (N_4820,N_4717,N_4658);
nor U4821 (N_4821,N_4650,N_4674);
xor U4822 (N_4822,N_4789,N_4726);
and U4823 (N_4823,N_4750,N_4628);
nor U4824 (N_4824,N_4799,N_4613);
and U4825 (N_4825,N_4744,N_4689);
nor U4826 (N_4826,N_4795,N_4694);
and U4827 (N_4827,N_4732,N_4623);
nor U4828 (N_4828,N_4741,N_4790);
or U4829 (N_4829,N_4695,N_4714);
xor U4830 (N_4830,N_4692,N_4618);
and U4831 (N_4831,N_4735,N_4609);
xor U4832 (N_4832,N_4696,N_4710);
or U4833 (N_4833,N_4749,N_4759);
and U4834 (N_4834,N_4639,N_4733);
nand U4835 (N_4835,N_4611,N_4620);
nand U4836 (N_4836,N_4675,N_4781);
nor U4837 (N_4837,N_4697,N_4768);
nor U4838 (N_4838,N_4648,N_4719);
or U4839 (N_4839,N_4716,N_4779);
nor U4840 (N_4840,N_4763,N_4640);
nor U4841 (N_4841,N_4748,N_4783);
nand U4842 (N_4842,N_4702,N_4602);
nand U4843 (N_4843,N_4764,N_4739);
or U4844 (N_4844,N_4728,N_4785);
and U4845 (N_4845,N_4681,N_4634);
xnor U4846 (N_4846,N_4691,N_4686);
or U4847 (N_4847,N_4601,N_4765);
or U4848 (N_4848,N_4718,N_4683);
or U4849 (N_4849,N_4659,N_4679);
or U4850 (N_4850,N_4678,N_4798);
and U4851 (N_4851,N_4606,N_4778);
and U4852 (N_4852,N_4771,N_4665);
xnor U4853 (N_4853,N_4622,N_4756);
or U4854 (N_4854,N_4704,N_4746);
and U4855 (N_4855,N_4610,N_4647);
or U4856 (N_4856,N_4657,N_4630);
nand U4857 (N_4857,N_4670,N_4605);
nand U4858 (N_4858,N_4615,N_4760);
nand U4859 (N_4859,N_4633,N_4753);
nand U4860 (N_4860,N_4793,N_4770);
nor U4861 (N_4861,N_4780,N_4711);
or U4862 (N_4862,N_4787,N_4699);
nor U4863 (N_4863,N_4667,N_4715);
and U4864 (N_4864,N_4705,N_4734);
nand U4865 (N_4865,N_4776,N_4645);
xor U4866 (N_4866,N_4617,N_4607);
and U4867 (N_4867,N_4742,N_4796);
nor U4868 (N_4868,N_4773,N_4641);
nand U4869 (N_4869,N_4700,N_4632);
nand U4870 (N_4870,N_4725,N_4646);
xnor U4871 (N_4871,N_4677,N_4724);
nand U4872 (N_4872,N_4745,N_4786);
nor U4873 (N_4873,N_4687,N_4747);
and U4874 (N_4874,N_4758,N_4791);
nor U4875 (N_4875,N_4631,N_4730);
xor U4876 (N_4876,N_4668,N_4706);
or U4877 (N_4877,N_4651,N_4738);
nand U4878 (N_4878,N_4762,N_4661);
xor U4879 (N_4879,N_4673,N_4772);
nor U4880 (N_4880,N_4698,N_4624);
nor U4881 (N_4881,N_4690,N_4684);
or U4882 (N_4882,N_4775,N_4731);
and U4883 (N_4883,N_4777,N_4761);
xnor U4884 (N_4884,N_4757,N_4693);
and U4885 (N_4885,N_4784,N_4788);
and U4886 (N_4886,N_4664,N_4722);
or U4887 (N_4887,N_4608,N_4660);
xor U4888 (N_4888,N_4655,N_4713);
nor U4889 (N_4889,N_4727,N_4712);
and U4890 (N_4890,N_4701,N_4642);
xnor U4891 (N_4891,N_4662,N_4708);
nor U4892 (N_4892,N_4625,N_4782);
or U4893 (N_4893,N_4740,N_4600);
nor U4894 (N_4894,N_4652,N_4627);
and U4895 (N_4895,N_4769,N_4636);
or U4896 (N_4896,N_4653,N_4737);
nand U4897 (N_4897,N_4614,N_4743);
nor U4898 (N_4898,N_4685,N_4680);
and U4899 (N_4899,N_4649,N_4721);
or U4900 (N_4900,N_4623,N_4781);
or U4901 (N_4901,N_4600,N_4653);
xnor U4902 (N_4902,N_4699,N_4774);
nand U4903 (N_4903,N_4728,N_4641);
nor U4904 (N_4904,N_4705,N_4618);
nand U4905 (N_4905,N_4646,N_4685);
nand U4906 (N_4906,N_4718,N_4669);
xnor U4907 (N_4907,N_4790,N_4788);
nand U4908 (N_4908,N_4600,N_4781);
nand U4909 (N_4909,N_4613,N_4674);
nand U4910 (N_4910,N_4775,N_4772);
nand U4911 (N_4911,N_4768,N_4702);
nand U4912 (N_4912,N_4792,N_4665);
nand U4913 (N_4913,N_4608,N_4659);
xor U4914 (N_4914,N_4605,N_4705);
nor U4915 (N_4915,N_4611,N_4702);
xor U4916 (N_4916,N_4756,N_4794);
nand U4917 (N_4917,N_4771,N_4798);
nor U4918 (N_4918,N_4693,N_4738);
nor U4919 (N_4919,N_4647,N_4709);
nand U4920 (N_4920,N_4612,N_4722);
or U4921 (N_4921,N_4688,N_4771);
and U4922 (N_4922,N_4771,N_4657);
nor U4923 (N_4923,N_4655,N_4641);
xor U4924 (N_4924,N_4708,N_4679);
xor U4925 (N_4925,N_4643,N_4741);
nor U4926 (N_4926,N_4658,N_4728);
nor U4927 (N_4927,N_4673,N_4612);
or U4928 (N_4928,N_4711,N_4645);
xor U4929 (N_4929,N_4773,N_4760);
nor U4930 (N_4930,N_4726,N_4785);
and U4931 (N_4931,N_4704,N_4739);
nand U4932 (N_4932,N_4611,N_4694);
or U4933 (N_4933,N_4609,N_4761);
xor U4934 (N_4934,N_4694,N_4603);
nand U4935 (N_4935,N_4695,N_4618);
xor U4936 (N_4936,N_4638,N_4758);
xnor U4937 (N_4937,N_4723,N_4643);
or U4938 (N_4938,N_4621,N_4684);
nand U4939 (N_4939,N_4706,N_4691);
xor U4940 (N_4940,N_4673,N_4759);
and U4941 (N_4941,N_4759,N_4734);
nor U4942 (N_4942,N_4758,N_4653);
or U4943 (N_4943,N_4612,N_4795);
or U4944 (N_4944,N_4712,N_4708);
or U4945 (N_4945,N_4721,N_4706);
xnor U4946 (N_4946,N_4706,N_4669);
or U4947 (N_4947,N_4736,N_4764);
and U4948 (N_4948,N_4609,N_4779);
xnor U4949 (N_4949,N_4626,N_4789);
and U4950 (N_4950,N_4634,N_4679);
nor U4951 (N_4951,N_4692,N_4659);
nand U4952 (N_4952,N_4679,N_4722);
nand U4953 (N_4953,N_4702,N_4676);
or U4954 (N_4954,N_4683,N_4715);
or U4955 (N_4955,N_4742,N_4647);
and U4956 (N_4956,N_4788,N_4629);
nor U4957 (N_4957,N_4725,N_4611);
or U4958 (N_4958,N_4796,N_4627);
nor U4959 (N_4959,N_4745,N_4778);
or U4960 (N_4960,N_4736,N_4647);
nand U4961 (N_4961,N_4659,N_4616);
or U4962 (N_4962,N_4614,N_4769);
and U4963 (N_4963,N_4669,N_4670);
xnor U4964 (N_4964,N_4743,N_4733);
or U4965 (N_4965,N_4732,N_4758);
and U4966 (N_4966,N_4765,N_4701);
or U4967 (N_4967,N_4714,N_4799);
nor U4968 (N_4968,N_4610,N_4746);
and U4969 (N_4969,N_4716,N_4721);
xor U4970 (N_4970,N_4674,N_4737);
nor U4971 (N_4971,N_4657,N_4693);
and U4972 (N_4972,N_4749,N_4799);
nor U4973 (N_4973,N_4661,N_4681);
nand U4974 (N_4974,N_4766,N_4654);
or U4975 (N_4975,N_4637,N_4646);
xnor U4976 (N_4976,N_4773,N_4610);
and U4977 (N_4977,N_4719,N_4654);
and U4978 (N_4978,N_4656,N_4676);
nor U4979 (N_4979,N_4757,N_4600);
and U4980 (N_4980,N_4671,N_4775);
nand U4981 (N_4981,N_4749,N_4668);
nand U4982 (N_4982,N_4603,N_4750);
xnor U4983 (N_4983,N_4654,N_4602);
and U4984 (N_4984,N_4608,N_4710);
and U4985 (N_4985,N_4791,N_4771);
nand U4986 (N_4986,N_4690,N_4730);
and U4987 (N_4987,N_4611,N_4726);
nor U4988 (N_4988,N_4713,N_4743);
nand U4989 (N_4989,N_4764,N_4734);
xor U4990 (N_4990,N_4742,N_4683);
xor U4991 (N_4991,N_4701,N_4682);
nor U4992 (N_4992,N_4640,N_4637);
nor U4993 (N_4993,N_4621,N_4680);
nand U4994 (N_4994,N_4790,N_4775);
xnor U4995 (N_4995,N_4784,N_4748);
nand U4996 (N_4996,N_4712,N_4782);
or U4997 (N_4997,N_4774,N_4737);
or U4998 (N_4998,N_4786,N_4642);
nand U4999 (N_4999,N_4690,N_4735);
or U5000 (N_5000,N_4915,N_4998);
nor U5001 (N_5001,N_4982,N_4885);
or U5002 (N_5002,N_4892,N_4948);
xnor U5003 (N_5003,N_4831,N_4932);
xnor U5004 (N_5004,N_4891,N_4873);
and U5005 (N_5005,N_4909,N_4936);
nand U5006 (N_5006,N_4843,N_4957);
and U5007 (N_5007,N_4938,N_4889);
nor U5008 (N_5008,N_4821,N_4958);
or U5009 (N_5009,N_4806,N_4952);
xnor U5010 (N_5010,N_4974,N_4816);
and U5011 (N_5011,N_4906,N_4835);
xnor U5012 (N_5012,N_4839,N_4870);
nand U5013 (N_5013,N_4829,N_4971);
xnor U5014 (N_5014,N_4973,N_4987);
and U5015 (N_5015,N_4991,N_4939);
or U5016 (N_5016,N_4819,N_4813);
nand U5017 (N_5017,N_4913,N_4901);
xor U5018 (N_5018,N_4921,N_4807);
nand U5019 (N_5019,N_4812,N_4865);
or U5020 (N_5020,N_4853,N_4801);
or U5021 (N_5021,N_4844,N_4988);
and U5022 (N_5022,N_4896,N_4852);
and U5023 (N_5023,N_4818,N_4809);
xor U5024 (N_5024,N_4934,N_4800);
nand U5025 (N_5025,N_4872,N_4840);
or U5026 (N_5026,N_4895,N_4900);
nor U5027 (N_5027,N_4834,N_4908);
xnor U5028 (N_5028,N_4856,N_4826);
xor U5029 (N_5029,N_4959,N_4850);
nand U5030 (N_5030,N_4965,N_4960);
xnor U5031 (N_5031,N_4802,N_4868);
or U5032 (N_5032,N_4810,N_4851);
or U5033 (N_5033,N_4949,N_4880);
or U5034 (N_5034,N_4846,N_4966);
nand U5035 (N_5035,N_4878,N_4942);
or U5036 (N_5036,N_4922,N_4953);
or U5037 (N_5037,N_4997,N_4989);
and U5038 (N_5038,N_4863,N_4832);
nor U5039 (N_5039,N_4907,N_4984);
xnor U5040 (N_5040,N_4916,N_4947);
nor U5041 (N_5041,N_4904,N_4980);
xor U5042 (N_5042,N_4940,N_4817);
nand U5043 (N_5043,N_4968,N_4924);
and U5044 (N_5044,N_4910,N_4943);
nand U5045 (N_5045,N_4955,N_4867);
xor U5046 (N_5046,N_4864,N_4847);
or U5047 (N_5047,N_4841,N_4963);
and U5048 (N_5048,N_4927,N_4905);
xnor U5049 (N_5049,N_4866,N_4979);
and U5050 (N_5050,N_4962,N_4879);
or U5051 (N_5051,N_4956,N_4838);
nor U5052 (N_5052,N_4887,N_4890);
nor U5053 (N_5053,N_4862,N_4860);
nor U5054 (N_5054,N_4950,N_4861);
xor U5055 (N_5055,N_4914,N_4898);
or U5056 (N_5056,N_4981,N_4875);
nor U5057 (N_5057,N_4894,N_4937);
and U5058 (N_5058,N_4995,N_4928);
or U5059 (N_5059,N_4899,N_4897);
nand U5060 (N_5060,N_4911,N_4884);
or U5061 (N_5061,N_4808,N_4869);
and U5062 (N_5062,N_4944,N_4859);
and U5063 (N_5063,N_4820,N_4985);
nor U5064 (N_5064,N_4970,N_4804);
xnor U5065 (N_5065,N_4920,N_4814);
and U5066 (N_5066,N_4992,N_4977);
nand U5067 (N_5067,N_4976,N_4803);
or U5068 (N_5068,N_4815,N_4858);
xor U5069 (N_5069,N_4929,N_4828);
xnor U5070 (N_5070,N_4871,N_4877);
nand U5071 (N_5071,N_4972,N_4999);
xor U5072 (N_5072,N_4886,N_4811);
xnor U5073 (N_5073,N_4912,N_4983);
nand U5074 (N_5074,N_4964,N_4931);
xnor U5075 (N_5075,N_4893,N_4946);
and U5076 (N_5076,N_4993,N_4805);
or U5077 (N_5077,N_4926,N_4941);
nor U5078 (N_5078,N_4823,N_4935);
nand U5079 (N_5079,N_4903,N_4978);
nand U5080 (N_5080,N_4822,N_4990);
or U5081 (N_5081,N_4967,N_4881);
or U5082 (N_5082,N_4825,N_4888);
or U5083 (N_5083,N_4994,N_4857);
and U5084 (N_5084,N_4975,N_4933);
nor U5085 (N_5085,N_4882,N_4951);
xor U5086 (N_5086,N_4925,N_4837);
and U5087 (N_5087,N_4855,N_4836);
nand U5088 (N_5088,N_4954,N_4849);
xor U5089 (N_5089,N_4883,N_4874);
and U5090 (N_5090,N_4848,N_4961);
nor U5091 (N_5091,N_4902,N_4923);
nand U5092 (N_5092,N_4845,N_4986);
nor U5093 (N_5093,N_4996,N_4830);
xnor U5094 (N_5094,N_4945,N_4827);
and U5095 (N_5095,N_4854,N_4842);
or U5096 (N_5096,N_4824,N_4930);
nand U5097 (N_5097,N_4969,N_4917);
nand U5098 (N_5098,N_4918,N_4919);
nor U5099 (N_5099,N_4833,N_4876);
xor U5100 (N_5100,N_4816,N_4883);
nand U5101 (N_5101,N_4867,N_4841);
nand U5102 (N_5102,N_4925,N_4876);
nand U5103 (N_5103,N_4811,N_4937);
or U5104 (N_5104,N_4881,N_4849);
and U5105 (N_5105,N_4844,N_4860);
xor U5106 (N_5106,N_4919,N_4859);
nand U5107 (N_5107,N_4873,N_4947);
and U5108 (N_5108,N_4999,N_4880);
or U5109 (N_5109,N_4903,N_4860);
nand U5110 (N_5110,N_4871,N_4907);
nor U5111 (N_5111,N_4936,N_4969);
and U5112 (N_5112,N_4823,N_4820);
or U5113 (N_5113,N_4843,N_4865);
nand U5114 (N_5114,N_4906,N_4936);
and U5115 (N_5115,N_4896,N_4897);
nand U5116 (N_5116,N_4839,N_4990);
nor U5117 (N_5117,N_4952,N_4897);
or U5118 (N_5118,N_4931,N_4873);
xor U5119 (N_5119,N_4995,N_4903);
nand U5120 (N_5120,N_4984,N_4888);
or U5121 (N_5121,N_4961,N_4949);
xor U5122 (N_5122,N_4894,N_4802);
nor U5123 (N_5123,N_4903,N_4823);
or U5124 (N_5124,N_4934,N_4815);
nand U5125 (N_5125,N_4868,N_4891);
and U5126 (N_5126,N_4854,N_4991);
and U5127 (N_5127,N_4821,N_4805);
nor U5128 (N_5128,N_4927,N_4860);
xnor U5129 (N_5129,N_4803,N_4809);
and U5130 (N_5130,N_4905,N_4843);
nand U5131 (N_5131,N_4856,N_4900);
nor U5132 (N_5132,N_4889,N_4870);
nand U5133 (N_5133,N_4813,N_4861);
nand U5134 (N_5134,N_4988,N_4856);
xnor U5135 (N_5135,N_4816,N_4833);
nor U5136 (N_5136,N_4897,N_4911);
and U5137 (N_5137,N_4888,N_4923);
nor U5138 (N_5138,N_4912,N_4988);
xnor U5139 (N_5139,N_4810,N_4917);
and U5140 (N_5140,N_4958,N_4875);
and U5141 (N_5141,N_4904,N_4999);
nor U5142 (N_5142,N_4809,N_4828);
xor U5143 (N_5143,N_4931,N_4989);
nand U5144 (N_5144,N_4913,N_4923);
nor U5145 (N_5145,N_4917,N_4937);
nor U5146 (N_5146,N_4933,N_4876);
and U5147 (N_5147,N_4991,N_4952);
nor U5148 (N_5148,N_4930,N_4842);
and U5149 (N_5149,N_4890,N_4986);
xor U5150 (N_5150,N_4831,N_4878);
nor U5151 (N_5151,N_4951,N_4885);
or U5152 (N_5152,N_4955,N_4921);
or U5153 (N_5153,N_4946,N_4914);
nand U5154 (N_5154,N_4818,N_4878);
or U5155 (N_5155,N_4909,N_4869);
and U5156 (N_5156,N_4809,N_4874);
nor U5157 (N_5157,N_4840,N_4947);
nor U5158 (N_5158,N_4939,N_4890);
or U5159 (N_5159,N_4885,N_4857);
nand U5160 (N_5160,N_4920,N_4839);
and U5161 (N_5161,N_4993,N_4987);
or U5162 (N_5162,N_4876,N_4884);
and U5163 (N_5163,N_4848,N_4884);
nand U5164 (N_5164,N_4829,N_4922);
and U5165 (N_5165,N_4815,N_4830);
nor U5166 (N_5166,N_4979,N_4996);
nand U5167 (N_5167,N_4907,N_4966);
xor U5168 (N_5168,N_4944,N_4853);
nor U5169 (N_5169,N_4854,N_4807);
nand U5170 (N_5170,N_4851,N_4910);
or U5171 (N_5171,N_4994,N_4829);
nand U5172 (N_5172,N_4922,N_4993);
xor U5173 (N_5173,N_4921,N_4833);
xor U5174 (N_5174,N_4893,N_4924);
nand U5175 (N_5175,N_4805,N_4802);
nand U5176 (N_5176,N_4853,N_4978);
nor U5177 (N_5177,N_4980,N_4803);
nor U5178 (N_5178,N_4873,N_4859);
xor U5179 (N_5179,N_4846,N_4912);
nand U5180 (N_5180,N_4843,N_4857);
nand U5181 (N_5181,N_4989,N_4864);
nor U5182 (N_5182,N_4921,N_4823);
or U5183 (N_5183,N_4881,N_4922);
nand U5184 (N_5184,N_4829,N_4929);
or U5185 (N_5185,N_4912,N_4806);
and U5186 (N_5186,N_4918,N_4809);
nor U5187 (N_5187,N_4954,N_4845);
nor U5188 (N_5188,N_4972,N_4842);
nand U5189 (N_5189,N_4881,N_4932);
xnor U5190 (N_5190,N_4996,N_4833);
or U5191 (N_5191,N_4992,N_4980);
or U5192 (N_5192,N_4854,N_4867);
or U5193 (N_5193,N_4923,N_4889);
xor U5194 (N_5194,N_4890,N_4863);
or U5195 (N_5195,N_4869,N_4812);
or U5196 (N_5196,N_4842,N_4962);
xnor U5197 (N_5197,N_4969,N_4945);
or U5198 (N_5198,N_4988,N_4960);
nand U5199 (N_5199,N_4896,N_4959);
and U5200 (N_5200,N_5154,N_5147);
nand U5201 (N_5201,N_5090,N_5112);
nor U5202 (N_5202,N_5063,N_5084);
and U5203 (N_5203,N_5070,N_5135);
nand U5204 (N_5204,N_5197,N_5015);
nor U5205 (N_5205,N_5034,N_5176);
nor U5206 (N_5206,N_5083,N_5156);
nor U5207 (N_5207,N_5093,N_5194);
xor U5208 (N_5208,N_5172,N_5150);
or U5209 (N_5209,N_5097,N_5199);
xor U5210 (N_5210,N_5082,N_5024);
nor U5211 (N_5211,N_5125,N_5107);
and U5212 (N_5212,N_5177,N_5038);
xor U5213 (N_5213,N_5127,N_5058);
nor U5214 (N_5214,N_5163,N_5062);
and U5215 (N_5215,N_5168,N_5109);
nor U5216 (N_5216,N_5078,N_5030);
nor U5217 (N_5217,N_5146,N_5032);
xor U5218 (N_5218,N_5026,N_5033);
nand U5219 (N_5219,N_5045,N_5118);
nor U5220 (N_5220,N_5020,N_5041);
nor U5221 (N_5221,N_5017,N_5099);
and U5222 (N_5222,N_5077,N_5061);
nor U5223 (N_5223,N_5133,N_5193);
nand U5224 (N_5224,N_5046,N_5003);
xnor U5225 (N_5225,N_5065,N_5067);
xnor U5226 (N_5226,N_5101,N_5142);
nor U5227 (N_5227,N_5126,N_5183);
or U5228 (N_5228,N_5191,N_5117);
nand U5229 (N_5229,N_5068,N_5031);
xor U5230 (N_5230,N_5180,N_5042);
or U5231 (N_5231,N_5123,N_5014);
and U5232 (N_5232,N_5013,N_5010);
xor U5233 (N_5233,N_5087,N_5174);
xnor U5234 (N_5234,N_5007,N_5162);
or U5235 (N_5235,N_5073,N_5171);
nor U5236 (N_5236,N_5170,N_5064);
nand U5237 (N_5237,N_5102,N_5182);
nor U5238 (N_5238,N_5119,N_5044);
or U5239 (N_5239,N_5186,N_5116);
xnor U5240 (N_5240,N_5100,N_5009);
or U5241 (N_5241,N_5029,N_5179);
and U5242 (N_5242,N_5155,N_5021);
nand U5243 (N_5243,N_5166,N_5131);
nor U5244 (N_5244,N_5108,N_5055);
xor U5245 (N_5245,N_5103,N_5027);
nor U5246 (N_5246,N_5023,N_5066);
and U5247 (N_5247,N_5105,N_5006);
xnor U5248 (N_5248,N_5114,N_5001);
and U5249 (N_5249,N_5169,N_5074);
nor U5250 (N_5250,N_5022,N_5059);
or U5251 (N_5251,N_5151,N_5095);
nor U5252 (N_5252,N_5075,N_5128);
nor U5253 (N_5253,N_5129,N_5040);
or U5254 (N_5254,N_5122,N_5164);
or U5255 (N_5255,N_5173,N_5195);
nand U5256 (N_5256,N_5005,N_5057);
nor U5257 (N_5257,N_5184,N_5048);
xnor U5258 (N_5258,N_5158,N_5165);
xnor U5259 (N_5259,N_5091,N_5196);
and U5260 (N_5260,N_5019,N_5137);
xor U5261 (N_5261,N_5076,N_5036);
or U5262 (N_5262,N_5069,N_5120);
nand U5263 (N_5263,N_5145,N_5160);
or U5264 (N_5264,N_5111,N_5192);
or U5265 (N_5265,N_5016,N_5043);
and U5266 (N_5266,N_5035,N_5051);
nand U5267 (N_5267,N_5148,N_5079);
or U5268 (N_5268,N_5106,N_5025);
and U5269 (N_5269,N_5188,N_5088);
xor U5270 (N_5270,N_5139,N_5152);
and U5271 (N_5271,N_5081,N_5161);
nor U5272 (N_5272,N_5187,N_5190);
nor U5273 (N_5273,N_5096,N_5086);
nor U5274 (N_5274,N_5167,N_5011);
and U5275 (N_5275,N_5149,N_5159);
xnor U5276 (N_5276,N_5056,N_5141);
xnor U5277 (N_5277,N_5175,N_5000);
xor U5278 (N_5278,N_5028,N_5002);
xor U5279 (N_5279,N_5130,N_5085);
nand U5280 (N_5280,N_5050,N_5132);
and U5281 (N_5281,N_5018,N_5110);
nand U5282 (N_5282,N_5039,N_5181);
nand U5283 (N_5283,N_5189,N_5094);
and U5284 (N_5284,N_5124,N_5134);
and U5285 (N_5285,N_5157,N_5072);
nand U5286 (N_5286,N_5037,N_5004);
xor U5287 (N_5287,N_5047,N_5080);
nand U5288 (N_5288,N_5115,N_5121);
xnor U5289 (N_5289,N_5071,N_5178);
or U5290 (N_5290,N_5185,N_5089);
nand U5291 (N_5291,N_5012,N_5138);
and U5292 (N_5292,N_5144,N_5143);
nor U5293 (N_5293,N_5113,N_5053);
nand U5294 (N_5294,N_5049,N_5136);
nand U5295 (N_5295,N_5153,N_5092);
xnor U5296 (N_5296,N_5098,N_5060);
xor U5297 (N_5297,N_5052,N_5104);
nand U5298 (N_5298,N_5198,N_5140);
nor U5299 (N_5299,N_5054,N_5008);
or U5300 (N_5300,N_5061,N_5096);
or U5301 (N_5301,N_5018,N_5006);
xor U5302 (N_5302,N_5035,N_5137);
xor U5303 (N_5303,N_5093,N_5110);
nor U5304 (N_5304,N_5063,N_5098);
xnor U5305 (N_5305,N_5074,N_5190);
nor U5306 (N_5306,N_5037,N_5088);
or U5307 (N_5307,N_5013,N_5106);
xnor U5308 (N_5308,N_5155,N_5114);
xnor U5309 (N_5309,N_5081,N_5077);
xnor U5310 (N_5310,N_5164,N_5141);
or U5311 (N_5311,N_5046,N_5088);
and U5312 (N_5312,N_5133,N_5040);
and U5313 (N_5313,N_5161,N_5091);
or U5314 (N_5314,N_5044,N_5162);
xor U5315 (N_5315,N_5055,N_5186);
nand U5316 (N_5316,N_5068,N_5175);
nor U5317 (N_5317,N_5085,N_5102);
xnor U5318 (N_5318,N_5149,N_5177);
and U5319 (N_5319,N_5121,N_5143);
or U5320 (N_5320,N_5076,N_5115);
and U5321 (N_5321,N_5172,N_5153);
nand U5322 (N_5322,N_5006,N_5030);
or U5323 (N_5323,N_5040,N_5058);
xnor U5324 (N_5324,N_5028,N_5014);
nor U5325 (N_5325,N_5146,N_5096);
nor U5326 (N_5326,N_5163,N_5074);
nand U5327 (N_5327,N_5041,N_5143);
nand U5328 (N_5328,N_5096,N_5025);
xor U5329 (N_5329,N_5139,N_5005);
or U5330 (N_5330,N_5129,N_5046);
nor U5331 (N_5331,N_5116,N_5054);
xor U5332 (N_5332,N_5160,N_5033);
xor U5333 (N_5333,N_5060,N_5064);
nor U5334 (N_5334,N_5124,N_5002);
nor U5335 (N_5335,N_5161,N_5000);
xnor U5336 (N_5336,N_5046,N_5049);
or U5337 (N_5337,N_5018,N_5086);
xnor U5338 (N_5338,N_5110,N_5031);
nor U5339 (N_5339,N_5169,N_5091);
nand U5340 (N_5340,N_5161,N_5164);
nand U5341 (N_5341,N_5058,N_5004);
nand U5342 (N_5342,N_5101,N_5080);
nand U5343 (N_5343,N_5163,N_5048);
or U5344 (N_5344,N_5109,N_5047);
xor U5345 (N_5345,N_5183,N_5062);
nor U5346 (N_5346,N_5192,N_5009);
and U5347 (N_5347,N_5081,N_5080);
nand U5348 (N_5348,N_5015,N_5054);
nor U5349 (N_5349,N_5142,N_5179);
nand U5350 (N_5350,N_5048,N_5106);
nor U5351 (N_5351,N_5100,N_5122);
and U5352 (N_5352,N_5047,N_5055);
nor U5353 (N_5353,N_5098,N_5120);
nand U5354 (N_5354,N_5131,N_5025);
or U5355 (N_5355,N_5152,N_5161);
and U5356 (N_5356,N_5150,N_5093);
xnor U5357 (N_5357,N_5198,N_5066);
and U5358 (N_5358,N_5090,N_5070);
and U5359 (N_5359,N_5102,N_5184);
and U5360 (N_5360,N_5016,N_5078);
nor U5361 (N_5361,N_5100,N_5181);
nand U5362 (N_5362,N_5009,N_5183);
or U5363 (N_5363,N_5124,N_5116);
nand U5364 (N_5364,N_5079,N_5190);
nand U5365 (N_5365,N_5136,N_5119);
and U5366 (N_5366,N_5040,N_5119);
xnor U5367 (N_5367,N_5064,N_5009);
and U5368 (N_5368,N_5132,N_5080);
or U5369 (N_5369,N_5150,N_5029);
or U5370 (N_5370,N_5157,N_5106);
nor U5371 (N_5371,N_5060,N_5138);
nor U5372 (N_5372,N_5171,N_5149);
xnor U5373 (N_5373,N_5199,N_5070);
nor U5374 (N_5374,N_5097,N_5175);
nand U5375 (N_5375,N_5068,N_5010);
xor U5376 (N_5376,N_5119,N_5197);
nand U5377 (N_5377,N_5045,N_5019);
or U5378 (N_5378,N_5006,N_5087);
nor U5379 (N_5379,N_5042,N_5007);
and U5380 (N_5380,N_5129,N_5054);
nand U5381 (N_5381,N_5072,N_5047);
or U5382 (N_5382,N_5095,N_5074);
nor U5383 (N_5383,N_5158,N_5051);
or U5384 (N_5384,N_5173,N_5131);
nor U5385 (N_5385,N_5168,N_5039);
xor U5386 (N_5386,N_5162,N_5182);
nand U5387 (N_5387,N_5011,N_5036);
xor U5388 (N_5388,N_5033,N_5002);
and U5389 (N_5389,N_5144,N_5152);
or U5390 (N_5390,N_5016,N_5001);
xnor U5391 (N_5391,N_5128,N_5066);
or U5392 (N_5392,N_5137,N_5068);
nand U5393 (N_5393,N_5024,N_5173);
nor U5394 (N_5394,N_5033,N_5117);
nand U5395 (N_5395,N_5053,N_5191);
nand U5396 (N_5396,N_5094,N_5053);
nor U5397 (N_5397,N_5125,N_5081);
nand U5398 (N_5398,N_5056,N_5033);
xnor U5399 (N_5399,N_5007,N_5000);
and U5400 (N_5400,N_5238,N_5323);
xor U5401 (N_5401,N_5206,N_5259);
nor U5402 (N_5402,N_5264,N_5336);
and U5403 (N_5403,N_5309,N_5283);
nor U5404 (N_5404,N_5210,N_5222);
nor U5405 (N_5405,N_5288,N_5330);
nor U5406 (N_5406,N_5253,N_5341);
nand U5407 (N_5407,N_5287,N_5257);
nand U5408 (N_5408,N_5396,N_5362);
nand U5409 (N_5409,N_5338,N_5386);
nand U5410 (N_5410,N_5232,N_5250);
xor U5411 (N_5411,N_5270,N_5337);
nor U5412 (N_5412,N_5392,N_5350);
or U5413 (N_5413,N_5344,N_5312);
and U5414 (N_5414,N_5237,N_5282);
nand U5415 (N_5415,N_5248,N_5387);
nand U5416 (N_5416,N_5200,N_5243);
and U5417 (N_5417,N_5390,N_5202);
nor U5418 (N_5418,N_5296,N_5249);
xnor U5419 (N_5419,N_5244,N_5346);
nor U5420 (N_5420,N_5213,N_5315);
xor U5421 (N_5421,N_5385,N_5240);
xnor U5422 (N_5422,N_5217,N_5317);
xor U5423 (N_5423,N_5394,N_5384);
nor U5424 (N_5424,N_5355,N_5221);
or U5425 (N_5425,N_5310,N_5335);
or U5426 (N_5426,N_5377,N_5354);
and U5427 (N_5427,N_5290,N_5300);
xnor U5428 (N_5428,N_5308,N_5298);
or U5429 (N_5429,N_5383,N_5280);
or U5430 (N_5430,N_5381,N_5365);
or U5431 (N_5431,N_5228,N_5242);
or U5432 (N_5432,N_5361,N_5379);
nor U5433 (N_5433,N_5297,N_5372);
nor U5434 (N_5434,N_5271,N_5274);
nor U5435 (N_5435,N_5316,N_5291);
xnor U5436 (N_5436,N_5299,N_5320);
nor U5437 (N_5437,N_5364,N_5289);
nand U5438 (N_5438,N_5371,N_5329);
or U5439 (N_5439,N_5233,N_5333);
nand U5440 (N_5440,N_5351,N_5269);
or U5441 (N_5441,N_5395,N_5214);
nor U5442 (N_5442,N_5295,N_5245);
or U5443 (N_5443,N_5332,N_5281);
and U5444 (N_5444,N_5260,N_5305);
nor U5445 (N_5445,N_5363,N_5227);
xnor U5446 (N_5446,N_5375,N_5339);
and U5447 (N_5447,N_5321,N_5302);
nor U5448 (N_5448,N_5314,N_5359);
and U5449 (N_5449,N_5224,N_5223);
and U5450 (N_5450,N_5307,N_5277);
and U5451 (N_5451,N_5360,N_5311);
xor U5452 (N_5452,N_5211,N_5328);
xnor U5453 (N_5453,N_5231,N_5239);
and U5454 (N_5454,N_5391,N_5398);
nand U5455 (N_5455,N_5201,N_5345);
nor U5456 (N_5456,N_5258,N_5215);
xor U5457 (N_5457,N_5216,N_5380);
nor U5458 (N_5458,N_5342,N_5207);
xor U5459 (N_5459,N_5251,N_5292);
xnor U5460 (N_5460,N_5236,N_5278);
nor U5461 (N_5461,N_5263,N_5225);
nand U5462 (N_5462,N_5266,N_5349);
nor U5463 (N_5463,N_5294,N_5261);
or U5464 (N_5464,N_5370,N_5252);
nor U5465 (N_5465,N_5268,N_5397);
and U5466 (N_5466,N_5319,N_5352);
nor U5467 (N_5467,N_5325,N_5208);
nand U5468 (N_5468,N_5322,N_5255);
and U5469 (N_5469,N_5357,N_5348);
nand U5470 (N_5470,N_5284,N_5212);
nor U5471 (N_5471,N_5306,N_5301);
and U5472 (N_5472,N_5367,N_5229);
nor U5473 (N_5473,N_5303,N_5209);
and U5474 (N_5474,N_5389,N_5234);
xor U5475 (N_5475,N_5230,N_5254);
xor U5476 (N_5476,N_5246,N_5399);
or U5477 (N_5477,N_5279,N_5376);
nor U5478 (N_5478,N_5369,N_5334);
and U5479 (N_5479,N_5358,N_5219);
xnor U5480 (N_5480,N_5313,N_5275);
or U5481 (N_5481,N_5327,N_5293);
nand U5482 (N_5482,N_5347,N_5286);
nand U5483 (N_5483,N_5204,N_5318);
and U5484 (N_5484,N_5326,N_5220);
or U5485 (N_5485,N_5247,N_5356);
nor U5486 (N_5486,N_5343,N_5304);
and U5487 (N_5487,N_5273,N_5374);
xor U5488 (N_5488,N_5331,N_5340);
nor U5489 (N_5489,N_5285,N_5256);
and U5490 (N_5490,N_5393,N_5235);
nand U5491 (N_5491,N_5218,N_5324);
and U5492 (N_5492,N_5241,N_5388);
xnor U5493 (N_5493,N_5226,N_5373);
nand U5494 (N_5494,N_5267,N_5382);
nand U5495 (N_5495,N_5366,N_5265);
nor U5496 (N_5496,N_5203,N_5272);
xor U5497 (N_5497,N_5276,N_5262);
nand U5498 (N_5498,N_5205,N_5368);
nand U5499 (N_5499,N_5353,N_5378);
nand U5500 (N_5500,N_5357,N_5251);
or U5501 (N_5501,N_5200,N_5371);
nor U5502 (N_5502,N_5347,N_5209);
nand U5503 (N_5503,N_5356,N_5387);
nor U5504 (N_5504,N_5389,N_5209);
and U5505 (N_5505,N_5215,N_5381);
xnor U5506 (N_5506,N_5284,N_5323);
and U5507 (N_5507,N_5272,N_5342);
nand U5508 (N_5508,N_5286,N_5203);
or U5509 (N_5509,N_5317,N_5374);
and U5510 (N_5510,N_5229,N_5299);
nand U5511 (N_5511,N_5347,N_5350);
or U5512 (N_5512,N_5348,N_5337);
and U5513 (N_5513,N_5210,N_5372);
and U5514 (N_5514,N_5369,N_5229);
xnor U5515 (N_5515,N_5211,N_5262);
xnor U5516 (N_5516,N_5209,N_5292);
xnor U5517 (N_5517,N_5261,N_5315);
nor U5518 (N_5518,N_5303,N_5359);
nand U5519 (N_5519,N_5318,N_5289);
xor U5520 (N_5520,N_5335,N_5390);
xor U5521 (N_5521,N_5231,N_5284);
and U5522 (N_5522,N_5350,N_5209);
or U5523 (N_5523,N_5295,N_5261);
nand U5524 (N_5524,N_5329,N_5261);
nor U5525 (N_5525,N_5335,N_5301);
nand U5526 (N_5526,N_5343,N_5370);
nand U5527 (N_5527,N_5356,N_5232);
nor U5528 (N_5528,N_5347,N_5394);
and U5529 (N_5529,N_5245,N_5240);
nand U5530 (N_5530,N_5383,N_5288);
or U5531 (N_5531,N_5256,N_5260);
nor U5532 (N_5532,N_5261,N_5300);
xor U5533 (N_5533,N_5302,N_5396);
or U5534 (N_5534,N_5351,N_5392);
nor U5535 (N_5535,N_5378,N_5359);
nor U5536 (N_5536,N_5223,N_5350);
or U5537 (N_5537,N_5395,N_5272);
nor U5538 (N_5538,N_5324,N_5302);
xor U5539 (N_5539,N_5271,N_5341);
xor U5540 (N_5540,N_5367,N_5218);
and U5541 (N_5541,N_5285,N_5292);
nor U5542 (N_5542,N_5216,N_5236);
or U5543 (N_5543,N_5392,N_5396);
or U5544 (N_5544,N_5308,N_5378);
nand U5545 (N_5545,N_5226,N_5325);
nand U5546 (N_5546,N_5319,N_5219);
nand U5547 (N_5547,N_5208,N_5298);
xnor U5548 (N_5548,N_5361,N_5350);
and U5549 (N_5549,N_5326,N_5203);
xnor U5550 (N_5550,N_5293,N_5369);
and U5551 (N_5551,N_5346,N_5285);
and U5552 (N_5552,N_5312,N_5386);
or U5553 (N_5553,N_5289,N_5250);
nand U5554 (N_5554,N_5224,N_5219);
or U5555 (N_5555,N_5366,N_5260);
xnor U5556 (N_5556,N_5350,N_5340);
or U5557 (N_5557,N_5374,N_5230);
or U5558 (N_5558,N_5379,N_5348);
and U5559 (N_5559,N_5263,N_5223);
and U5560 (N_5560,N_5329,N_5256);
and U5561 (N_5561,N_5286,N_5243);
and U5562 (N_5562,N_5366,N_5318);
xor U5563 (N_5563,N_5283,N_5236);
or U5564 (N_5564,N_5293,N_5300);
xor U5565 (N_5565,N_5200,N_5257);
or U5566 (N_5566,N_5312,N_5255);
nand U5567 (N_5567,N_5263,N_5329);
nand U5568 (N_5568,N_5343,N_5273);
nand U5569 (N_5569,N_5340,N_5330);
and U5570 (N_5570,N_5215,N_5263);
or U5571 (N_5571,N_5243,N_5394);
nand U5572 (N_5572,N_5209,N_5253);
or U5573 (N_5573,N_5358,N_5275);
or U5574 (N_5574,N_5228,N_5375);
nand U5575 (N_5575,N_5391,N_5314);
nor U5576 (N_5576,N_5335,N_5340);
or U5577 (N_5577,N_5207,N_5256);
xnor U5578 (N_5578,N_5268,N_5266);
nand U5579 (N_5579,N_5277,N_5217);
nand U5580 (N_5580,N_5272,N_5287);
nor U5581 (N_5581,N_5214,N_5292);
or U5582 (N_5582,N_5203,N_5219);
nand U5583 (N_5583,N_5353,N_5256);
nand U5584 (N_5584,N_5201,N_5306);
xnor U5585 (N_5585,N_5203,N_5287);
nor U5586 (N_5586,N_5315,N_5205);
nor U5587 (N_5587,N_5399,N_5326);
nand U5588 (N_5588,N_5343,N_5219);
or U5589 (N_5589,N_5387,N_5256);
or U5590 (N_5590,N_5206,N_5325);
or U5591 (N_5591,N_5397,N_5243);
xnor U5592 (N_5592,N_5271,N_5202);
nor U5593 (N_5593,N_5353,N_5360);
nand U5594 (N_5594,N_5311,N_5320);
xnor U5595 (N_5595,N_5212,N_5255);
nor U5596 (N_5596,N_5351,N_5204);
nand U5597 (N_5597,N_5235,N_5326);
xnor U5598 (N_5598,N_5203,N_5213);
nor U5599 (N_5599,N_5340,N_5381);
xnor U5600 (N_5600,N_5555,N_5505);
and U5601 (N_5601,N_5460,N_5583);
nor U5602 (N_5602,N_5418,N_5480);
nor U5603 (N_5603,N_5552,N_5519);
xor U5604 (N_5604,N_5446,N_5501);
and U5605 (N_5605,N_5550,N_5454);
or U5606 (N_5606,N_5523,N_5544);
or U5607 (N_5607,N_5512,N_5477);
nor U5608 (N_5608,N_5518,N_5577);
and U5609 (N_5609,N_5411,N_5504);
nor U5610 (N_5610,N_5484,N_5497);
xnor U5611 (N_5611,N_5511,N_5543);
nor U5612 (N_5612,N_5459,N_5409);
or U5613 (N_5613,N_5462,N_5469);
and U5614 (N_5614,N_5472,N_5467);
nand U5615 (N_5615,N_5545,N_5572);
or U5616 (N_5616,N_5553,N_5458);
nor U5617 (N_5617,N_5468,N_5506);
and U5618 (N_5618,N_5440,N_5529);
and U5619 (N_5619,N_5508,N_5428);
nand U5620 (N_5620,N_5489,N_5490);
or U5621 (N_5621,N_5502,N_5499);
nand U5622 (N_5622,N_5455,N_5481);
xnor U5623 (N_5623,N_5548,N_5558);
nor U5624 (N_5624,N_5566,N_5561);
or U5625 (N_5625,N_5534,N_5461);
or U5626 (N_5626,N_5444,N_5495);
or U5627 (N_5627,N_5582,N_5594);
or U5628 (N_5628,N_5406,N_5524);
xor U5629 (N_5629,N_5551,N_5403);
and U5630 (N_5630,N_5588,N_5598);
and U5631 (N_5631,N_5465,N_5479);
nand U5632 (N_5632,N_5562,N_5414);
or U5633 (N_5633,N_5424,N_5421);
nor U5634 (N_5634,N_5537,N_5590);
nor U5635 (N_5635,N_5532,N_5464);
or U5636 (N_5636,N_5563,N_5533);
nor U5637 (N_5637,N_5522,N_5434);
or U5638 (N_5638,N_5536,N_5457);
and U5639 (N_5639,N_5515,N_5585);
or U5640 (N_5640,N_5436,N_5422);
or U5641 (N_5641,N_5596,N_5581);
xnor U5642 (N_5642,N_5439,N_5416);
nor U5643 (N_5643,N_5575,N_5541);
nor U5644 (N_5644,N_5516,N_5432);
nor U5645 (N_5645,N_5520,N_5576);
xnor U5646 (N_5646,N_5456,N_5503);
nor U5647 (N_5647,N_5531,N_5586);
xnor U5648 (N_5648,N_5571,N_5540);
and U5649 (N_5649,N_5412,N_5452);
nor U5650 (N_5650,N_5592,N_5538);
nor U5651 (N_5651,N_5599,N_5494);
nand U5652 (N_5652,N_5500,N_5400);
or U5653 (N_5653,N_5591,N_5405);
or U5654 (N_5654,N_5569,N_5466);
or U5655 (N_5655,N_5483,N_5478);
nand U5656 (N_5656,N_5574,N_5413);
and U5657 (N_5657,N_5450,N_5514);
and U5658 (N_5658,N_5485,N_5560);
and U5659 (N_5659,N_5493,N_5567);
and U5660 (N_5660,N_5535,N_5445);
xnor U5661 (N_5661,N_5539,N_5476);
and U5662 (N_5662,N_5438,N_5573);
xor U5663 (N_5663,N_5557,N_5530);
or U5664 (N_5664,N_5463,N_5587);
and U5665 (N_5665,N_5473,N_5447);
nor U5666 (N_5666,N_5407,N_5488);
nor U5667 (N_5667,N_5401,N_5580);
or U5668 (N_5668,N_5408,N_5417);
xor U5669 (N_5669,N_5584,N_5420);
xnor U5670 (N_5670,N_5559,N_5443);
or U5671 (N_5671,N_5429,N_5509);
and U5672 (N_5672,N_5542,N_5433);
xnor U5673 (N_5673,N_5423,N_5517);
or U5674 (N_5674,N_5482,N_5597);
or U5675 (N_5675,N_5507,N_5496);
xnor U5676 (N_5676,N_5510,N_5492);
nand U5677 (N_5677,N_5431,N_5570);
and U5678 (N_5678,N_5528,N_5449);
nor U5679 (N_5679,N_5498,N_5593);
nand U5680 (N_5680,N_5521,N_5474);
nand U5681 (N_5681,N_5410,N_5426);
nor U5682 (N_5682,N_5442,N_5453);
and U5683 (N_5683,N_5475,N_5487);
xor U5684 (N_5684,N_5549,N_5564);
nand U5685 (N_5685,N_5595,N_5427);
or U5686 (N_5686,N_5513,N_5402);
xnor U5687 (N_5687,N_5486,N_5554);
or U5688 (N_5688,N_5404,N_5578);
xor U5689 (N_5689,N_5430,N_5419);
xor U5690 (N_5690,N_5546,N_5526);
xor U5691 (N_5691,N_5441,N_5435);
nand U5692 (N_5692,N_5425,N_5451);
or U5693 (N_5693,N_5527,N_5547);
nand U5694 (N_5694,N_5556,N_5579);
and U5695 (N_5695,N_5470,N_5491);
xor U5696 (N_5696,N_5565,N_5448);
and U5697 (N_5697,N_5589,N_5568);
or U5698 (N_5698,N_5471,N_5525);
xnor U5699 (N_5699,N_5437,N_5415);
nand U5700 (N_5700,N_5543,N_5578);
or U5701 (N_5701,N_5423,N_5569);
nand U5702 (N_5702,N_5579,N_5557);
nor U5703 (N_5703,N_5413,N_5568);
nor U5704 (N_5704,N_5485,N_5418);
xnor U5705 (N_5705,N_5581,N_5521);
nand U5706 (N_5706,N_5410,N_5492);
xor U5707 (N_5707,N_5406,N_5494);
and U5708 (N_5708,N_5569,N_5541);
nand U5709 (N_5709,N_5430,N_5444);
or U5710 (N_5710,N_5478,N_5468);
and U5711 (N_5711,N_5594,N_5541);
xnor U5712 (N_5712,N_5533,N_5461);
xor U5713 (N_5713,N_5526,N_5434);
or U5714 (N_5714,N_5450,N_5470);
nand U5715 (N_5715,N_5543,N_5529);
nor U5716 (N_5716,N_5456,N_5545);
or U5717 (N_5717,N_5497,N_5530);
nand U5718 (N_5718,N_5548,N_5492);
nor U5719 (N_5719,N_5596,N_5488);
nor U5720 (N_5720,N_5409,N_5527);
xor U5721 (N_5721,N_5502,N_5512);
nand U5722 (N_5722,N_5500,N_5519);
xnor U5723 (N_5723,N_5513,N_5541);
or U5724 (N_5724,N_5466,N_5581);
and U5725 (N_5725,N_5488,N_5412);
and U5726 (N_5726,N_5527,N_5566);
or U5727 (N_5727,N_5447,N_5523);
nand U5728 (N_5728,N_5501,N_5485);
or U5729 (N_5729,N_5421,N_5432);
and U5730 (N_5730,N_5454,N_5557);
or U5731 (N_5731,N_5468,N_5438);
and U5732 (N_5732,N_5599,N_5443);
xnor U5733 (N_5733,N_5557,N_5559);
and U5734 (N_5734,N_5407,N_5497);
xnor U5735 (N_5735,N_5448,N_5481);
and U5736 (N_5736,N_5504,N_5470);
nand U5737 (N_5737,N_5585,N_5430);
and U5738 (N_5738,N_5562,N_5426);
and U5739 (N_5739,N_5531,N_5490);
nand U5740 (N_5740,N_5416,N_5573);
or U5741 (N_5741,N_5533,N_5428);
xor U5742 (N_5742,N_5543,N_5502);
nand U5743 (N_5743,N_5471,N_5494);
or U5744 (N_5744,N_5578,N_5410);
or U5745 (N_5745,N_5570,N_5481);
or U5746 (N_5746,N_5523,N_5599);
and U5747 (N_5747,N_5519,N_5547);
nor U5748 (N_5748,N_5503,N_5553);
nor U5749 (N_5749,N_5524,N_5456);
nand U5750 (N_5750,N_5587,N_5450);
or U5751 (N_5751,N_5527,N_5453);
or U5752 (N_5752,N_5470,N_5505);
and U5753 (N_5753,N_5511,N_5524);
or U5754 (N_5754,N_5479,N_5464);
nand U5755 (N_5755,N_5442,N_5562);
and U5756 (N_5756,N_5501,N_5490);
nand U5757 (N_5757,N_5593,N_5426);
nand U5758 (N_5758,N_5567,N_5410);
nand U5759 (N_5759,N_5459,N_5515);
xor U5760 (N_5760,N_5583,N_5406);
nand U5761 (N_5761,N_5416,N_5428);
nor U5762 (N_5762,N_5498,N_5538);
xnor U5763 (N_5763,N_5451,N_5597);
nor U5764 (N_5764,N_5536,N_5413);
and U5765 (N_5765,N_5488,N_5566);
and U5766 (N_5766,N_5550,N_5429);
nand U5767 (N_5767,N_5464,N_5531);
or U5768 (N_5768,N_5499,N_5460);
or U5769 (N_5769,N_5436,N_5469);
and U5770 (N_5770,N_5430,N_5455);
xnor U5771 (N_5771,N_5479,N_5406);
or U5772 (N_5772,N_5541,N_5411);
nor U5773 (N_5773,N_5544,N_5498);
nor U5774 (N_5774,N_5526,N_5485);
nand U5775 (N_5775,N_5552,N_5459);
xor U5776 (N_5776,N_5512,N_5535);
nor U5777 (N_5777,N_5583,N_5491);
nor U5778 (N_5778,N_5472,N_5486);
nor U5779 (N_5779,N_5562,N_5558);
nor U5780 (N_5780,N_5582,N_5473);
nand U5781 (N_5781,N_5593,N_5583);
or U5782 (N_5782,N_5451,N_5591);
or U5783 (N_5783,N_5580,N_5439);
or U5784 (N_5784,N_5575,N_5478);
and U5785 (N_5785,N_5496,N_5495);
xnor U5786 (N_5786,N_5502,N_5566);
nor U5787 (N_5787,N_5513,N_5597);
and U5788 (N_5788,N_5546,N_5466);
xnor U5789 (N_5789,N_5510,N_5435);
nor U5790 (N_5790,N_5466,N_5597);
nor U5791 (N_5791,N_5583,N_5550);
xnor U5792 (N_5792,N_5493,N_5434);
nand U5793 (N_5793,N_5410,N_5505);
xnor U5794 (N_5794,N_5551,N_5435);
xnor U5795 (N_5795,N_5430,N_5530);
and U5796 (N_5796,N_5511,N_5484);
nand U5797 (N_5797,N_5570,N_5534);
nand U5798 (N_5798,N_5539,N_5465);
or U5799 (N_5799,N_5423,N_5558);
xor U5800 (N_5800,N_5780,N_5746);
xor U5801 (N_5801,N_5618,N_5745);
nand U5802 (N_5802,N_5647,N_5695);
nand U5803 (N_5803,N_5787,N_5794);
xor U5804 (N_5804,N_5681,N_5732);
nor U5805 (N_5805,N_5636,N_5737);
and U5806 (N_5806,N_5799,N_5699);
nor U5807 (N_5807,N_5782,N_5710);
nor U5808 (N_5808,N_5676,N_5701);
nor U5809 (N_5809,N_5649,N_5735);
nand U5810 (N_5810,N_5715,N_5606);
nor U5811 (N_5811,N_5684,N_5631);
or U5812 (N_5812,N_5702,N_5633);
nor U5813 (N_5813,N_5602,N_5688);
nor U5814 (N_5814,N_5690,N_5734);
nand U5815 (N_5815,N_5640,N_5784);
or U5816 (N_5816,N_5739,N_5608);
and U5817 (N_5817,N_5652,N_5668);
nand U5818 (N_5818,N_5788,N_5726);
nor U5819 (N_5819,N_5617,N_5660);
nand U5820 (N_5820,N_5654,N_5667);
nand U5821 (N_5821,N_5741,N_5712);
nand U5822 (N_5822,N_5758,N_5722);
or U5823 (N_5823,N_5718,N_5653);
nand U5824 (N_5824,N_5719,N_5616);
xnor U5825 (N_5825,N_5641,N_5709);
nor U5826 (N_5826,N_5796,N_5656);
nor U5827 (N_5827,N_5723,N_5630);
and U5828 (N_5828,N_5779,N_5672);
or U5829 (N_5829,N_5757,N_5603);
xor U5830 (N_5830,N_5687,N_5748);
or U5831 (N_5831,N_5786,N_5717);
xor U5832 (N_5832,N_5626,N_5771);
and U5833 (N_5833,N_5697,N_5772);
and U5834 (N_5834,N_5624,N_5670);
or U5835 (N_5835,N_5696,N_5728);
xnor U5836 (N_5836,N_5713,N_5655);
or U5837 (N_5837,N_5673,N_5763);
nand U5838 (N_5838,N_5762,N_5691);
or U5839 (N_5839,N_5604,N_5749);
xnor U5840 (N_5840,N_5611,N_5642);
and U5841 (N_5841,N_5623,N_5674);
and U5842 (N_5842,N_5694,N_5774);
and U5843 (N_5843,N_5738,N_5760);
nor U5844 (N_5844,N_5704,N_5679);
nand U5845 (N_5845,N_5620,N_5650);
nor U5846 (N_5846,N_5662,N_5659);
xnor U5847 (N_5847,N_5683,N_5638);
nor U5848 (N_5848,N_5761,N_5783);
xnor U5849 (N_5849,N_5797,N_5751);
or U5850 (N_5850,N_5756,N_5613);
xnor U5851 (N_5851,N_5768,N_5663);
nor U5852 (N_5852,N_5629,N_5635);
nor U5853 (N_5853,N_5675,N_5628);
or U5854 (N_5854,N_5736,N_5773);
and U5855 (N_5855,N_5750,N_5610);
or U5856 (N_5856,N_5625,N_5680);
xnor U5857 (N_5857,N_5619,N_5733);
xor U5858 (N_5858,N_5791,N_5744);
and U5859 (N_5859,N_5708,N_5765);
or U5860 (N_5860,N_5692,N_5648);
nor U5861 (N_5861,N_5781,N_5764);
or U5862 (N_5862,N_5789,N_5689);
nor U5863 (N_5863,N_5790,N_5643);
and U5864 (N_5864,N_5686,N_5615);
nand U5865 (N_5865,N_5767,N_5705);
xor U5866 (N_5866,N_5612,N_5727);
or U5867 (N_5867,N_5622,N_5716);
nand U5868 (N_5868,N_5698,N_5775);
xnor U5869 (N_5869,N_5682,N_5747);
or U5870 (N_5870,N_5706,N_5777);
nor U5871 (N_5871,N_5766,N_5651);
nor U5872 (N_5872,N_5645,N_5609);
nor U5873 (N_5873,N_5671,N_5785);
xor U5874 (N_5874,N_5795,N_5637);
nand U5875 (N_5875,N_5605,N_5634);
xnor U5876 (N_5876,N_5644,N_5664);
and U5877 (N_5877,N_5601,N_5769);
and U5878 (N_5878,N_5770,N_5752);
and U5879 (N_5879,N_5731,N_5753);
or U5880 (N_5880,N_5776,N_5798);
or U5881 (N_5881,N_5661,N_5632);
or U5882 (N_5882,N_5754,N_5729);
xor U5883 (N_5883,N_5600,N_5730);
nand U5884 (N_5884,N_5721,N_5685);
xnor U5885 (N_5885,N_5725,N_5703);
nand U5886 (N_5886,N_5627,N_5759);
nor U5887 (N_5887,N_5714,N_5700);
nand U5888 (N_5888,N_5639,N_5724);
nand U5889 (N_5889,N_5742,N_5665);
nor U5890 (N_5890,N_5711,N_5621);
and U5891 (N_5891,N_5666,N_5793);
nor U5892 (N_5892,N_5607,N_5707);
or U5893 (N_5893,N_5658,N_5677);
nand U5894 (N_5894,N_5693,N_5778);
xnor U5895 (N_5895,N_5720,N_5792);
nor U5896 (N_5896,N_5678,N_5669);
and U5897 (N_5897,N_5646,N_5740);
and U5898 (N_5898,N_5657,N_5614);
or U5899 (N_5899,N_5755,N_5743);
or U5900 (N_5900,N_5643,N_5746);
nor U5901 (N_5901,N_5782,N_5643);
nand U5902 (N_5902,N_5663,N_5682);
nand U5903 (N_5903,N_5656,N_5652);
xor U5904 (N_5904,N_5702,N_5729);
and U5905 (N_5905,N_5686,N_5794);
and U5906 (N_5906,N_5724,N_5780);
or U5907 (N_5907,N_5790,N_5724);
and U5908 (N_5908,N_5792,N_5649);
xor U5909 (N_5909,N_5647,N_5752);
or U5910 (N_5910,N_5688,N_5727);
nand U5911 (N_5911,N_5651,N_5714);
or U5912 (N_5912,N_5774,N_5685);
and U5913 (N_5913,N_5778,N_5690);
xor U5914 (N_5914,N_5696,N_5638);
nand U5915 (N_5915,N_5773,N_5622);
nand U5916 (N_5916,N_5663,N_5694);
or U5917 (N_5917,N_5641,N_5606);
or U5918 (N_5918,N_5689,N_5704);
nor U5919 (N_5919,N_5745,N_5779);
nor U5920 (N_5920,N_5787,N_5641);
nand U5921 (N_5921,N_5613,N_5615);
nand U5922 (N_5922,N_5775,N_5696);
or U5923 (N_5923,N_5772,N_5775);
nor U5924 (N_5924,N_5705,N_5738);
or U5925 (N_5925,N_5792,N_5622);
or U5926 (N_5926,N_5621,N_5623);
or U5927 (N_5927,N_5632,N_5656);
or U5928 (N_5928,N_5745,N_5794);
nand U5929 (N_5929,N_5650,N_5681);
and U5930 (N_5930,N_5703,N_5696);
and U5931 (N_5931,N_5684,N_5640);
nand U5932 (N_5932,N_5606,N_5720);
nand U5933 (N_5933,N_5734,N_5692);
xor U5934 (N_5934,N_5635,N_5776);
and U5935 (N_5935,N_5689,N_5611);
and U5936 (N_5936,N_5677,N_5615);
nand U5937 (N_5937,N_5652,N_5613);
nor U5938 (N_5938,N_5627,N_5760);
xor U5939 (N_5939,N_5650,N_5667);
and U5940 (N_5940,N_5795,N_5787);
nand U5941 (N_5941,N_5783,N_5644);
or U5942 (N_5942,N_5771,N_5709);
and U5943 (N_5943,N_5640,N_5783);
and U5944 (N_5944,N_5763,N_5733);
nand U5945 (N_5945,N_5601,N_5759);
xnor U5946 (N_5946,N_5753,N_5767);
and U5947 (N_5947,N_5673,N_5649);
xnor U5948 (N_5948,N_5719,N_5686);
and U5949 (N_5949,N_5780,N_5791);
and U5950 (N_5950,N_5669,N_5657);
xor U5951 (N_5951,N_5601,N_5626);
nand U5952 (N_5952,N_5673,N_5658);
or U5953 (N_5953,N_5669,N_5652);
and U5954 (N_5954,N_5687,N_5738);
xor U5955 (N_5955,N_5635,N_5630);
nor U5956 (N_5956,N_5608,N_5694);
nor U5957 (N_5957,N_5695,N_5762);
xnor U5958 (N_5958,N_5693,N_5620);
and U5959 (N_5959,N_5708,N_5794);
nor U5960 (N_5960,N_5684,N_5783);
nor U5961 (N_5961,N_5628,N_5760);
xnor U5962 (N_5962,N_5724,N_5743);
nand U5963 (N_5963,N_5715,N_5745);
and U5964 (N_5964,N_5746,N_5676);
and U5965 (N_5965,N_5722,N_5639);
nor U5966 (N_5966,N_5678,N_5697);
nand U5967 (N_5967,N_5701,N_5782);
nor U5968 (N_5968,N_5678,N_5712);
nand U5969 (N_5969,N_5700,N_5710);
nor U5970 (N_5970,N_5798,N_5792);
xnor U5971 (N_5971,N_5736,N_5656);
nor U5972 (N_5972,N_5700,N_5797);
or U5973 (N_5973,N_5731,N_5777);
or U5974 (N_5974,N_5606,N_5690);
xor U5975 (N_5975,N_5667,N_5629);
or U5976 (N_5976,N_5765,N_5611);
and U5977 (N_5977,N_5647,N_5634);
nor U5978 (N_5978,N_5690,N_5684);
and U5979 (N_5979,N_5698,N_5705);
nand U5980 (N_5980,N_5709,N_5644);
xor U5981 (N_5981,N_5698,N_5759);
or U5982 (N_5982,N_5603,N_5663);
xnor U5983 (N_5983,N_5612,N_5788);
xor U5984 (N_5984,N_5675,N_5622);
nand U5985 (N_5985,N_5714,N_5799);
or U5986 (N_5986,N_5756,N_5754);
and U5987 (N_5987,N_5641,N_5689);
or U5988 (N_5988,N_5681,N_5625);
xnor U5989 (N_5989,N_5627,N_5689);
nand U5990 (N_5990,N_5627,N_5633);
or U5991 (N_5991,N_5753,N_5626);
xnor U5992 (N_5992,N_5631,N_5725);
or U5993 (N_5993,N_5612,N_5741);
nand U5994 (N_5994,N_5623,N_5642);
or U5995 (N_5995,N_5645,N_5713);
nand U5996 (N_5996,N_5610,N_5764);
or U5997 (N_5997,N_5728,N_5722);
or U5998 (N_5998,N_5629,N_5779);
or U5999 (N_5999,N_5679,N_5632);
and U6000 (N_6000,N_5916,N_5880);
xor U6001 (N_6001,N_5985,N_5894);
nor U6002 (N_6002,N_5874,N_5929);
and U6003 (N_6003,N_5865,N_5914);
and U6004 (N_6004,N_5942,N_5906);
and U6005 (N_6005,N_5863,N_5861);
nand U6006 (N_6006,N_5869,N_5912);
nand U6007 (N_6007,N_5956,N_5901);
nand U6008 (N_6008,N_5803,N_5954);
xor U6009 (N_6009,N_5802,N_5815);
nand U6010 (N_6010,N_5896,N_5948);
nor U6011 (N_6011,N_5936,N_5826);
or U6012 (N_6012,N_5975,N_5873);
xnor U6013 (N_6013,N_5945,N_5836);
nor U6014 (N_6014,N_5862,N_5959);
nor U6015 (N_6015,N_5932,N_5966);
nand U6016 (N_6016,N_5980,N_5918);
nor U6017 (N_6017,N_5951,N_5893);
nand U6018 (N_6018,N_5997,N_5976);
xnor U6019 (N_6019,N_5859,N_5995);
nor U6020 (N_6020,N_5983,N_5847);
nand U6021 (N_6021,N_5941,N_5950);
or U6022 (N_6022,N_5907,N_5828);
and U6023 (N_6023,N_5899,N_5852);
nand U6024 (N_6024,N_5813,N_5905);
xnor U6025 (N_6025,N_5903,N_5943);
or U6026 (N_6026,N_5807,N_5969);
xor U6027 (N_6027,N_5931,N_5804);
nand U6028 (N_6028,N_5871,N_5811);
nand U6029 (N_6029,N_5844,N_5938);
nand U6030 (N_6030,N_5827,N_5808);
nand U6031 (N_6031,N_5935,N_5934);
xnor U6032 (N_6032,N_5940,N_5961);
nor U6033 (N_6033,N_5921,N_5825);
xor U6034 (N_6034,N_5977,N_5832);
nor U6035 (N_6035,N_5973,N_5917);
nor U6036 (N_6036,N_5879,N_5947);
or U6037 (N_6037,N_5970,N_5854);
nor U6038 (N_6038,N_5992,N_5930);
nor U6039 (N_6039,N_5988,N_5843);
nor U6040 (N_6040,N_5989,N_5994);
or U6041 (N_6041,N_5814,N_5974);
or U6042 (N_6042,N_5849,N_5913);
nor U6043 (N_6043,N_5923,N_5864);
nand U6044 (N_6044,N_5919,N_5888);
and U6045 (N_6045,N_5810,N_5845);
xnor U6046 (N_6046,N_5805,N_5897);
xnor U6047 (N_6047,N_5927,N_5818);
nand U6048 (N_6048,N_5908,N_5915);
nor U6049 (N_6049,N_5999,N_5860);
and U6050 (N_6050,N_5993,N_5881);
or U6051 (N_6051,N_5911,N_5822);
nor U6052 (N_6052,N_5851,N_5839);
or U6053 (N_6053,N_5886,N_5925);
nand U6054 (N_6054,N_5955,N_5960);
or U6055 (N_6055,N_5830,N_5885);
and U6056 (N_6056,N_5867,N_5957);
or U6057 (N_6057,N_5823,N_5816);
nor U6058 (N_6058,N_5904,N_5853);
or U6059 (N_6059,N_5909,N_5834);
or U6060 (N_6060,N_5987,N_5882);
nor U6061 (N_6061,N_5926,N_5883);
and U6062 (N_6062,N_5986,N_5878);
xnor U6063 (N_6063,N_5842,N_5900);
xor U6064 (N_6064,N_5809,N_5922);
or U6065 (N_6065,N_5981,N_5962);
xor U6066 (N_6066,N_5996,N_5949);
and U6067 (N_6067,N_5857,N_5991);
nor U6068 (N_6068,N_5990,N_5856);
xnor U6069 (N_6069,N_5846,N_5806);
and U6070 (N_6070,N_5958,N_5963);
and U6071 (N_6071,N_5819,N_5801);
and U6072 (N_6072,N_5829,N_5920);
nor U6073 (N_6073,N_5939,N_5875);
nand U6074 (N_6074,N_5946,N_5964);
nand U6075 (N_6075,N_5850,N_5812);
or U6076 (N_6076,N_5820,N_5877);
nor U6077 (N_6077,N_5933,N_5835);
nor U6078 (N_6078,N_5876,N_5984);
xnor U6079 (N_6079,N_5891,N_5872);
nor U6080 (N_6080,N_5892,N_5972);
and U6081 (N_6081,N_5821,N_5887);
xor U6082 (N_6082,N_5910,N_5944);
or U6083 (N_6083,N_5841,N_5979);
nand U6084 (N_6084,N_5833,N_5965);
nand U6085 (N_6085,N_5800,N_5868);
nor U6086 (N_6086,N_5928,N_5952);
xnor U6087 (N_6087,N_5895,N_5870);
xor U6088 (N_6088,N_5998,N_5890);
and U6089 (N_6089,N_5968,N_5837);
nand U6090 (N_6090,N_5840,N_5937);
xnor U6091 (N_6091,N_5924,N_5855);
or U6092 (N_6092,N_5967,N_5889);
or U6093 (N_6093,N_5858,N_5902);
nor U6094 (N_6094,N_5866,N_5978);
or U6095 (N_6095,N_5848,N_5817);
xor U6096 (N_6096,N_5953,N_5884);
and U6097 (N_6097,N_5824,N_5982);
and U6098 (N_6098,N_5898,N_5831);
and U6099 (N_6099,N_5971,N_5838);
xnor U6100 (N_6100,N_5826,N_5914);
nor U6101 (N_6101,N_5890,N_5922);
or U6102 (N_6102,N_5849,N_5959);
nand U6103 (N_6103,N_5846,N_5982);
and U6104 (N_6104,N_5880,N_5890);
nor U6105 (N_6105,N_5917,N_5963);
and U6106 (N_6106,N_5900,N_5958);
or U6107 (N_6107,N_5831,N_5982);
or U6108 (N_6108,N_5819,N_5836);
and U6109 (N_6109,N_5989,N_5953);
nor U6110 (N_6110,N_5809,N_5884);
and U6111 (N_6111,N_5964,N_5941);
nand U6112 (N_6112,N_5964,N_5816);
nor U6113 (N_6113,N_5913,N_5802);
nand U6114 (N_6114,N_5966,N_5845);
and U6115 (N_6115,N_5945,N_5891);
xor U6116 (N_6116,N_5859,N_5873);
and U6117 (N_6117,N_5995,N_5853);
nor U6118 (N_6118,N_5851,N_5834);
nor U6119 (N_6119,N_5929,N_5985);
xor U6120 (N_6120,N_5841,N_5910);
nor U6121 (N_6121,N_5952,N_5832);
xor U6122 (N_6122,N_5838,N_5815);
nand U6123 (N_6123,N_5998,N_5881);
xor U6124 (N_6124,N_5875,N_5842);
nand U6125 (N_6125,N_5809,N_5956);
nor U6126 (N_6126,N_5833,N_5908);
xnor U6127 (N_6127,N_5959,N_5814);
nor U6128 (N_6128,N_5839,N_5865);
and U6129 (N_6129,N_5902,N_5941);
and U6130 (N_6130,N_5801,N_5905);
nor U6131 (N_6131,N_5824,N_5878);
and U6132 (N_6132,N_5831,N_5820);
xor U6133 (N_6133,N_5953,N_5919);
and U6134 (N_6134,N_5807,N_5846);
nor U6135 (N_6135,N_5989,N_5885);
or U6136 (N_6136,N_5809,N_5902);
and U6137 (N_6137,N_5968,N_5955);
xor U6138 (N_6138,N_5851,N_5916);
nor U6139 (N_6139,N_5800,N_5929);
nand U6140 (N_6140,N_5989,N_5810);
and U6141 (N_6141,N_5864,N_5964);
xor U6142 (N_6142,N_5973,N_5887);
nor U6143 (N_6143,N_5911,N_5828);
nor U6144 (N_6144,N_5952,N_5956);
nor U6145 (N_6145,N_5913,N_5985);
xor U6146 (N_6146,N_5946,N_5838);
and U6147 (N_6147,N_5932,N_5918);
or U6148 (N_6148,N_5992,N_5859);
nand U6149 (N_6149,N_5937,N_5886);
xnor U6150 (N_6150,N_5934,N_5835);
xnor U6151 (N_6151,N_5905,N_5916);
and U6152 (N_6152,N_5906,N_5894);
or U6153 (N_6153,N_5982,N_5966);
nor U6154 (N_6154,N_5918,N_5869);
or U6155 (N_6155,N_5819,N_5948);
and U6156 (N_6156,N_5863,N_5866);
and U6157 (N_6157,N_5848,N_5860);
or U6158 (N_6158,N_5841,N_5880);
or U6159 (N_6159,N_5809,N_5906);
and U6160 (N_6160,N_5888,N_5871);
or U6161 (N_6161,N_5849,N_5950);
xnor U6162 (N_6162,N_5867,N_5803);
nor U6163 (N_6163,N_5980,N_5990);
xor U6164 (N_6164,N_5909,N_5844);
nor U6165 (N_6165,N_5894,N_5807);
and U6166 (N_6166,N_5917,N_5866);
nor U6167 (N_6167,N_5963,N_5889);
and U6168 (N_6168,N_5858,N_5833);
nand U6169 (N_6169,N_5941,N_5960);
nor U6170 (N_6170,N_5953,N_5846);
nor U6171 (N_6171,N_5817,N_5850);
nand U6172 (N_6172,N_5895,N_5910);
or U6173 (N_6173,N_5920,N_5838);
nor U6174 (N_6174,N_5930,N_5965);
xor U6175 (N_6175,N_5887,N_5926);
or U6176 (N_6176,N_5956,N_5857);
and U6177 (N_6177,N_5838,N_5988);
nor U6178 (N_6178,N_5989,N_5903);
or U6179 (N_6179,N_5936,N_5918);
nand U6180 (N_6180,N_5908,N_5830);
or U6181 (N_6181,N_5878,N_5929);
and U6182 (N_6182,N_5988,N_5980);
nand U6183 (N_6183,N_5997,N_5851);
nand U6184 (N_6184,N_5898,N_5844);
or U6185 (N_6185,N_5831,N_5827);
xnor U6186 (N_6186,N_5949,N_5885);
xnor U6187 (N_6187,N_5928,N_5947);
nor U6188 (N_6188,N_5842,N_5869);
or U6189 (N_6189,N_5823,N_5998);
and U6190 (N_6190,N_5884,N_5817);
xor U6191 (N_6191,N_5942,N_5980);
xor U6192 (N_6192,N_5812,N_5891);
or U6193 (N_6193,N_5897,N_5816);
xnor U6194 (N_6194,N_5914,N_5841);
and U6195 (N_6195,N_5800,N_5807);
nor U6196 (N_6196,N_5887,N_5968);
or U6197 (N_6197,N_5818,N_5900);
nor U6198 (N_6198,N_5835,N_5983);
nor U6199 (N_6199,N_5809,N_5936);
or U6200 (N_6200,N_6170,N_6024);
and U6201 (N_6201,N_6192,N_6076);
nor U6202 (N_6202,N_6087,N_6162);
xor U6203 (N_6203,N_6010,N_6189);
nand U6204 (N_6204,N_6169,N_6048);
xnor U6205 (N_6205,N_6075,N_6098);
and U6206 (N_6206,N_6091,N_6196);
and U6207 (N_6207,N_6119,N_6140);
xnor U6208 (N_6208,N_6051,N_6017);
and U6209 (N_6209,N_6052,N_6164);
or U6210 (N_6210,N_6131,N_6155);
xnor U6211 (N_6211,N_6022,N_6159);
nor U6212 (N_6212,N_6197,N_6148);
or U6213 (N_6213,N_6013,N_6103);
or U6214 (N_6214,N_6102,N_6107);
or U6215 (N_6215,N_6109,N_6199);
xor U6216 (N_6216,N_6007,N_6030);
nand U6217 (N_6217,N_6080,N_6019);
xor U6218 (N_6218,N_6021,N_6161);
nor U6219 (N_6219,N_6183,N_6151);
nand U6220 (N_6220,N_6032,N_6039);
and U6221 (N_6221,N_6049,N_6128);
or U6222 (N_6222,N_6000,N_6187);
and U6223 (N_6223,N_6168,N_6094);
nand U6224 (N_6224,N_6176,N_6029);
nor U6225 (N_6225,N_6079,N_6110);
or U6226 (N_6226,N_6043,N_6115);
xnor U6227 (N_6227,N_6071,N_6020);
and U6228 (N_6228,N_6114,N_6191);
xnor U6229 (N_6229,N_6068,N_6121);
and U6230 (N_6230,N_6085,N_6108);
xnor U6231 (N_6231,N_6088,N_6046);
xnor U6232 (N_6232,N_6179,N_6171);
or U6233 (N_6233,N_6070,N_6012);
nor U6234 (N_6234,N_6047,N_6064);
or U6235 (N_6235,N_6058,N_6113);
nand U6236 (N_6236,N_6129,N_6074);
xnor U6237 (N_6237,N_6042,N_6056);
nand U6238 (N_6238,N_6180,N_6090);
xor U6239 (N_6239,N_6186,N_6037);
xnor U6240 (N_6240,N_6116,N_6157);
nand U6241 (N_6241,N_6057,N_6027);
nand U6242 (N_6242,N_6003,N_6072);
or U6243 (N_6243,N_6040,N_6005);
nor U6244 (N_6244,N_6073,N_6190);
xor U6245 (N_6245,N_6106,N_6004);
and U6246 (N_6246,N_6077,N_6055);
and U6247 (N_6247,N_6099,N_6104);
or U6248 (N_6248,N_6036,N_6025);
nor U6249 (N_6249,N_6001,N_6044);
xor U6250 (N_6250,N_6084,N_6124);
nor U6251 (N_6251,N_6153,N_6078);
nor U6252 (N_6252,N_6002,N_6134);
or U6253 (N_6253,N_6093,N_6137);
nand U6254 (N_6254,N_6156,N_6172);
nand U6255 (N_6255,N_6143,N_6060);
nor U6256 (N_6256,N_6092,N_6066);
xor U6257 (N_6257,N_6086,N_6011);
or U6258 (N_6258,N_6163,N_6125);
xnor U6259 (N_6259,N_6152,N_6033);
nand U6260 (N_6260,N_6178,N_6082);
xnor U6261 (N_6261,N_6041,N_6081);
nor U6262 (N_6262,N_6132,N_6194);
xnor U6263 (N_6263,N_6038,N_6138);
or U6264 (N_6264,N_6141,N_6136);
or U6265 (N_6265,N_6028,N_6018);
xor U6266 (N_6266,N_6133,N_6184);
and U6267 (N_6267,N_6101,N_6089);
and U6268 (N_6268,N_6195,N_6142);
xnor U6269 (N_6269,N_6146,N_6139);
and U6270 (N_6270,N_6185,N_6009);
and U6271 (N_6271,N_6160,N_6045);
nor U6272 (N_6272,N_6198,N_6135);
xnor U6273 (N_6273,N_6126,N_6026);
nand U6274 (N_6274,N_6150,N_6112);
or U6275 (N_6275,N_6120,N_6167);
and U6276 (N_6276,N_6158,N_6117);
nand U6277 (N_6277,N_6069,N_6065);
xor U6278 (N_6278,N_6123,N_6034);
nand U6279 (N_6279,N_6111,N_6054);
xnor U6280 (N_6280,N_6177,N_6118);
and U6281 (N_6281,N_6062,N_6127);
xnor U6282 (N_6282,N_6015,N_6061);
or U6283 (N_6283,N_6014,N_6097);
or U6284 (N_6284,N_6130,N_6188);
or U6285 (N_6285,N_6100,N_6006);
nor U6286 (N_6286,N_6059,N_6174);
nand U6287 (N_6287,N_6147,N_6031);
xnor U6288 (N_6288,N_6181,N_6145);
nand U6289 (N_6289,N_6096,N_6175);
xnor U6290 (N_6290,N_6193,N_6067);
nand U6291 (N_6291,N_6154,N_6023);
nor U6292 (N_6292,N_6166,N_6149);
nor U6293 (N_6293,N_6144,N_6095);
and U6294 (N_6294,N_6165,N_6182);
nor U6295 (N_6295,N_6105,N_6122);
xnor U6296 (N_6296,N_6008,N_6050);
nand U6297 (N_6297,N_6053,N_6035);
and U6298 (N_6298,N_6063,N_6173);
xnor U6299 (N_6299,N_6016,N_6083);
nand U6300 (N_6300,N_6156,N_6007);
nand U6301 (N_6301,N_6116,N_6040);
xor U6302 (N_6302,N_6150,N_6171);
or U6303 (N_6303,N_6194,N_6153);
and U6304 (N_6304,N_6071,N_6037);
xnor U6305 (N_6305,N_6091,N_6186);
and U6306 (N_6306,N_6012,N_6160);
and U6307 (N_6307,N_6198,N_6099);
and U6308 (N_6308,N_6100,N_6158);
nor U6309 (N_6309,N_6112,N_6019);
nor U6310 (N_6310,N_6144,N_6082);
nor U6311 (N_6311,N_6119,N_6181);
nor U6312 (N_6312,N_6184,N_6178);
and U6313 (N_6313,N_6176,N_6123);
xor U6314 (N_6314,N_6033,N_6059);
nor U6315 (N_6315,N_6189,N_6159);
xnor U6316 (N_6316,N_6197,N_6130);
and U6317 (N_6317,N_6100,N_6067);
or U6318 (N_6318,N_6155,N_6044);
nand U6319 (N_6319,N_6184,N_6029);
and U6320 (N_6320,N_6048,N_6120);
or U6321 (N_6321,N_6074,N_6113);
and U6322 (N_6322,N_6059,N_6005);
nand U6323 (N_6323,N_6045,N_6098);
nor U6324 (N_6324,N_6161,N_6084);
xnor U6325 (N_6325,N_6061,N_6097);
and U6326 (N_6326,N_6130,N_6105);
nand U6327 (N_6327,N_6022,N_6015);
and U6328 (N_6328,N_6084,N_6032);
xnor U6329 (N_6329,N_6077,N_6134);
xor U6330 (N_6330,N_6120,N_6139);
and U6331 (N_6331,N_6003,N_6176);
nor U6332 (N_6332,N_6144,N_6059);
or U6333 (N_6333,N_6036,N_6049);
nor U6334 (N_6334,N_6057,N_6015);
and U6335 (N_6335,N_6096,N_6157);
xor U6336 (N_6336,N_6161,N_6191);
or U6337 (N_6337,N_6074,N_6102);
nor U6338 (N_6338,N_6142,N_6055);
nor U6339 (N_6339,N_6075,N_6073);
and U6340 (N_6340,N_6128,N_6152);
nand U6341 (N_6341,N_6188,N_6022);
nor U6342 (N_6342,N_6105,N_6087);
xnor U6343 (N_6343,N_6065,N_6030);
nor U6344 (N_6344,N_6078,N_6124);
nor U6345 (N_6345,N_6124,N_6179);
nand U6346 (N_6346,N_6042,N_6128);
xor U6347 (N_6347,N_6026,N_6007);
nand U6348 (N_6348,N_6029,N_6057);
or U6349 (N_6349,N_6124,N_6132);
or U6350 (N_6350,N_6165,N_6156);
and U6351 (N_6351,N_6133,N_6073);
or U6352 (N_6352,N_6183,N_6110);
xor U6353 (N_6353,N_6072,N_6175);
nand U6354 (N_6354,N_6166,N_6199);
nor U6355 (N_6355,N_6097,N_6106);
nand U6356 (N_6356,N_6174,N_6089);
xnor U6357 (N_6357,N_6063,N_6022);
and U6358 (N_6358,N_6040,N_6101);
nand U6359 (N_6359,N_6099,N_6082);
or U6360 (N_6360,N_6185,N_6071);
and U6361 (N_6361,N_6079,N_6124);
or U6362 (N_6362,N_6119,N_6065);
nand U6363 (N_6363,N_6017,N_6128);
nand U6364 (N_6364,N_6142,N_6138);
xor U6365 (N_6365,N_6071,N_6103);
xor U6366 (N_6366,N_6019,N_6017);
or U6367 (N_6367,N_6164,N_6056);
nand U6368 (N_6368,N_6034,N_6170);
nor U6369 (N_6369,N_6009,N_6006);
nand U6370 (N_6370,N_6049,N_6013);
nand U6371 (N_6371,N_6018,N_6190);
nor U6372 (N_6372,N_6130,N_6190);
and U6373 (N_6373,N_6035,N_6146);
nor U6374 (N_6374,N_6181,N_6027);
xnor U6375 (N_6375,N_6169,N_6054);
xor U6376 (N_6376,N_6091,N_6004);
and U6377 (N_6377,N_6026,N_6185);
and U6378 (N_6378,N_6134,N_6011);
or U6379 (N_6379,N_6000,N_6149);
nor U6380 (N_6380,N_6059,N_6162);
xor U6381 (N_6381,N_6004,N_6077);
or U6382 (N_6382,N_6118,N_6191);
nand U6383 (N_6383,N_6167,N_6170);
nand U6384 (N_6384,N_6166,N_6106);
nor U6385 (N_6385,N_6093,N_6002);
and U6386 (N_6386,N_6049,N_6199);
xnor U6387 (N_6387,N_6162,N_6136);
or U6388 (N_6388,N_6056,N_6012);
or U6389 (N_6389,N_6051,N_6062);
nor U6390 (N_6390,N_6029,N_6074);
or U6391 (N_6391,N_6060,N_6017);
xnor U6392 (N_6392,N_6018,N_6068);
and U6393 (N_6393,N_6029,N_6086);
or U6394 (N_6394,N_6191,N_6141);
and U6395 (N_6395,N_6121,N_6038);
or U6396 (N_6396,N_6176,N_6109);
or U6397 (N_6397,N_6083,N_6025);
or U6398 (N_6398,N_6073,N_6188);
nor U6399 (N_6399,N_6156,N_6068);
xnor U6400 (N_6400,N_6244,N_6268);
and U6401 (N_6401,N_6397,N_6352);
nand U6402 (N_6402,N_6277,N_6335);
xor U6403 (N_6403,N_6217,N_6325);
or U6404 (N_6404,N_6236,N_6247);
and U6405 (N_6405,N_6326,N_6355);
xnor U6406 (N_6406,N_6253,N_6350);
xnor U6407 (N_6407,N_6299,N_6390);
nand U6408 (N_6408,N_6233,N_6235);
nor U6409 (N_6409,N_6317,N_6227);
or U6410 (N_6410,N_6209,N_6257);
or U6411 (N_6411,N_6238,N_6384);
nand U6412 (N_6412,N_6279,N_6290);
xnor U6413 (N_6413,N_6309,N_6369);
xnor U6414 (N_6414,N_6376,N_6319);
nand U6415 (N_6415,N_6315,N_6220);
nand U6416 (N_6416,N_6379,N_6380);
and U6417 (N_6417,N_6264,N_6362);
and U6418 (N_6418,N_6243,N_6222);
xor U6419 (N_6419,N_6221,N_6381);
nand U6420 (N_6420,N_6385,N_6337);
nor U6421 (N_6421,N_6311,N_6274);
nand U6422 (N_6422,N_6214,N_6330);
and U6423 (N_6423,N_6202,N_6305);
and U6424 (N_6424,N_6373,N_6344);
nand U6425 (N_6425,N_6357,N_6327);
nor U6426 (N_6426,N_6377,N_6246);
or U6427 (N_6427,N_6275,N_6256);
nor U6428 (N_6428,N_6356,N_6241);
xor U6429 (N_6429,N_6292,N_6307);
and U6430 (N_6430,N_6278,N_6273);
nor U6431 (N_6431,N_6231,N_6333);
nand U6432 (N_6432,N_6225,N_6254);
xor U6433 (N_6433,N_6383,N_6210);
nand U6434 (N_6434,N_6271,N_6258);
nor U6435 (N_6435,N_6282,N_6249);
or U6436 (N_6436,N_6321,N_6294);
nor U6437 (N_6437,N_6239,N_6353);
nor U6438 (N_6438,N_6331,N_6371);
nor U6439 (N_6439,N_6200,N_6375);
and U6440 (N_6440,N_6252,N_6389);
nand U6441 (N_6441,N_6208,N_6363);
and U6442 (N_6442,N_6266,N_6285);
nand U6443 (N_6443,N_6374,N_6270);
nor U6444 (N_6444,N_6391,N_6295);
nor U6445 (N_6445,N_6250,N_6365);
nor U6446 (N_6446,N_6395,N_6284);
xnor U6447 (N_6447,N_6320,N_6338);
xnor U6448 (N_6448,N_6367,N_6240);
nor U6449 (N_6449,N_6394,N_6261);
or U6450 (N_6450,N_6229,N_6280);
nand U6451 (N_6451,N_6201,N_6289);
and U6452 (N_6452,N_6354,N_6205);
or U6453 (N_6453,N_6312,N_6297);
nand U6454 (N_6454,N_6260,N_6328);
and U6455 (N_6455,N_6263,N_6393);
nor U6456 (N_6456,N_6334,N_6219);
or U6457 (N_6457,N_6303,N_6358);
nand U6458 (N_6458,N_6316,N_6207);
nor U6459 (N_6459,N_6230,N_6370);
xor U6460 (N_6460,N_6286,N_6346);
xnor U6461 (N_6461,N_6242,N_6206);
xnor U6462 (N_6462,N_6388,N_6361);
and U6463 (N_6463,N_6378,N_6298);
or U6464 (N_6464,N_6399,N_6226);
or U6465 (N_6465,N_6396,N_6324);
nand U6466 (N_6466,N_6234,N_6215);
xnor U6467 (N_6467,N_6359,N_6204);
nand U6468 (N_6468,N_6287,N_6213);
and U6469 (N_6469,N_6329,N_6313);
nor U6470 (N_6470,N_6341,N_6339);
and U6471 (N_6471,N_6281,N_6237);
nor U6472 (N_6472,N_6387,N_6343);
nor U6473 (N_6473,N_6348,N_6364);
and U6474 (N_6474,N_6216,N_6288);
or U6475 (N_6475,N_6302,N_6347);
xnor U6476 (N_6476,N_6228,N_6269);
xor U6477 (N_6477,N_6310,N_6308);
nor U6478 (N_6478,N_6336,N_6224);
nor U6479 (N_6479,N_6265,N_6322);
xnor U6480 (N_6480,N_6276,N_6245);
and U6481 (N_6481,N_6349,N_6267);
and U6482 (N_6482,N_6300,N_6291);
or U6483 (N_6483,N_6345,N_6259);
nand U6484 (N_6484,N_6314,N_6323);
nor U6485 (N_6485,N_6293,N_6392);
xor U6486 (N_6486,N_6255,N_6368);
and U6487 (N_6487,N_6262,N_6212);
xor U6488 (N_6488,N_6283,N_6366);
and U6489 (N_6489,N_6223,N_6398);
or U6490 (N_6490,N_6232,N_6203);
and U6491 (N_6491,N_6318,N_6211);
or U6492 (N_6492,N_6251,N_6332);
or U6493 (N_6493,N_6301,N_6296);
nor U6494 (N_6494,N_6218,N_6272);
nand U6495 (N_6495,N_6248,N_6372);
xnor U6496 (N_6496,N_6351,N_6342);
and U6497 (N_6497,N_6306,N_6382);
and U6498 (N_6498,N_6340,N_6360);
nor U6499 (N_6499,N_6304,N_6386);
nor U6500 (N_6500,N_6282,N_6251);
xnor U6501 (N_6501,N_6205,N_6377);
nor U6502 (N_6502,N_6242,N_6240);
and U6503 (N_6503,N_6297,N_6315);
nand U6504 (N_6504,N_6356,N_6323);
nor U6505 (N_6505,N_6214,N_6302);
and U6506 (N_6506,N_6252,N_6336);
xnor U6507 (N_6507,N_6302,N_6263);
or U6508 (N_6508,N_6216,N_6322);
nor U6509 (N_6509,N_6363,N_6268);
or U6510 (N_6510,N_6287,N_6242);
and U6511 (N_6511,N_6292,N_6397);
xor U6512 (N_6512,N_6258,N_6321);
and U6513 (N_6513,N_6212,N_6365);
nand U6514 (N_6514,N_6252,N_6253);
nor U6515 (N_6515,N_6383,N_6251);
nand U6516 (N_6516,N_6260,N_6312);
xor U6517 (N_6517,N_6319,N_6274);
nand U6518 (N_6518,N_6303,N_6356);
or U6519 (N_6519,N_6201,N_6333);
nor U6520 (N_6520,N_6336,N_6289);
nor U6521 (N_6521,N_6222,N_6375);
nor U6522 (N_6522,N_6277,N_6368);
nand U6523 (N_6523,N_6267,N_6235);
xor U6524 (N_6524,N_6337,N_6335);
and U6525 (N_6525,N_6366,N_6264);
nor U6526 (N_6526,N_6379,N_6213);
or U6527 (N_6527,N_6312,N_6268);
nor U6528 (N_6528,N_6263,N_6352);
and U6529 (N_6529,N_6224,N_6313);
nor U6530 (N_6530,N_6223,N_6338);
nand U6531 (N_6531,N_6316,N_6204);
nand U6532 (N_6532,N_6389,N_6359);
xnor U6533 (N_6533,N_6389,N_6371);
nor U6534 (N_6534,N_6268,N_6348);
nand U6535 (N_6535,N_6385,N_6214);
and U6536 (N_6536,N_6343,N_6359);
or U6537 (N_6537,N_6322,N_6392);
or U6538 (N_6538,N_6266,N_6209);
nand U6539 (N_6539,N_6368,N_6396);
or U6540 (N_6540,N_6276,N_6293);
nor U6541 (N_6541,N_6223,N_6218);
xnor U6542 (N_6542,N_6202,N_6327);
nor U6543 (N_6543,N_6228,N_6371);
nand U6544 (N_6544,N_6310,N_6397);
xnor U6545 (N_6545,N_6340,N_6281);
and U6546 (N_6546,N_6388,N_6230);
nor U6547 (N_6547,N_6235,N_6269);
nor U6548 (N_6548,N_6333,N_6316);
and U6549 (N_6549,N_6304,N_6355);
nand U6550 (N_6550,N_6253,N_6347);
and U6551 (N_6551,N_6327,N_6311);
or U6552 (N_6552,N_6382,N_6215);
nand U6553 (N_6553,N_6232,N_6227);
and U6554 (N_6554,N_6331,N_6377);
nor U6555 (N_6555,N_6318,N_6364);
nand U6556 (N_6556,N_6307,N_6334);
xnor U6557 (N_6557,N_6241,N_6217);
or U6558 (N_6558,N_6320,N_6279);
or U6559 (N_6559,N_6229,N_6265);
xor U6560 (N_6560,N_6229,N_6206);
nand U6561 (N_6561,N_6331,N_6251);
nand U6562 (N_6562,N_6334,N_6279);
nor U6563 (N_6563,N_6313,N_6335);
or U6564 (N_6564,N_6258,N_6254);
nor U6565 (N_6565,N_6266,N_6223);
nand U6566 (N_6566,N_6376,N_6351);
or U6567 (N_6567,N_6319,N_6360);
nand U6568 (N_6568,N_6324,N_6377);
and U6569 (N_6569,N_6376,N_6386);
or U6570 (N_6570,N_6292,N_6245);
or U6571 (N_6571,N_6376,N_6234);
or U6572 (N_6572,N_6330,N_6327);
or U6573 (N_6573,N_6329,N_6206);
nor U6574 (N_6574,N_6341,N_6211);
nor U6575 (N_6575,N_6372,N_6331);
xor U6576 (N_6576,N_6229,N_6385);
nor U6577 (N_6577,N_6271,N_6322);
xor U6578 (N_6578,N_6344,N_6333);
and U6579 (N_6579,N_6368,N_6331);
or U6580 (N_6580,N_6302,N_6320);
nor U6581 (N_6581,N_6270,N_6204);
nor U6582 (N_6582,N_6338,N_6392);
and U6583 (N_6583,N_6273,N_6397);
nor U6584 (N_6584,N_6257,N_6260);
xnor U6585 (N_6585,N_6298,N_6308);
xor U6586 (N_6586,N_6205,N_6330);
and U6587 (N_6587,N_6224,N_6231);
xor U6588 (N_6588,N_6341,N_6220);
nor U6589 (N_6589,N_6219,N_6290);
and U6590 (N_6590,N_6212,N_6374);
nor U6591 (N_6591,N_6361,N_6261);
or U6592 (N_6592,N_6252,N_6317);
and U6593 (N_6593,N_6275,N_6349);
or U6594 (N_6594,N_6395,N_6256);
and U6595 (N_6595,N_6272,N_6383);
nand U6596 (N_6596,N_6334,N_6255);
nor U6597 (N_6597,N_6262,N_6267);
and U6598 (N_6598,N_6215,N_6225);
or U6599 (N_6599,N_6334,N_6352);
or U6600 (N_6600,N_6539,N_6465);
and U6601 (N_6601,N_6444,N_6557);
or U6602 (N_6602,N_6563,N_6541);
or U6603 (N_6603,N_6499,N_6418);
nor U6604 (N_6604,N_6427,N_6508);
and U6605 (N_6605,N_6515,N_6533);
or U6606 (N_6606,N_6431,N_6560);
xor U6607 (N_6607,N_6435,N_6459);
nand U6608 (N_6608,N_6480,N_6489);
or U6609 (N_6609,N_6577,N_6407);
and U6610 (N_6610,N_6487,N_6502);
xor U6611 (N_6611,N_6512,N_6482);
and U6612 (N_6612,N_6597,N_6583);
xor U6613 (N_6613,N_6421,N_6440);
and U6614 (N_6614,N_6599,N_6478);
and U6615 (N_6615,N_6536,N_6438);
xor U6616 (N_6616,N_6494,N_6552);
nand U6617 (N_6617,N_6424,N_6432);
nand U6618 (N_6618,N_6486,N_6446);
or U6619 (N_6619,N_6522,N_6400);
or U6620 (N_6620,N_6544,N_6466);
nor U6621 (N_6621,N_6419,N_6517);
nor U6622 (N_6622,N_6523,N_6568);
xnor U6623 (N_6623,N_6509,N_6469);
nor U6624 (N_6624,N_6475,N_6524);
and U6625 (N_6625,N_6507,N_6437);
nor U6626 (N_6626,N_6518,N_6485);
and U6627 (N_6627,N_6406,N_6417);
nor U6628 (N_6628,N_6570,N_6575);
nor U6629 (N_6629,N_6450,N_6497);
or U6630 (N_6630,N_6455,N_6590);
and U6631 (N_6631,N_6554,N_6545);
or U6632 (N_6632,N_6439,N_6445);
or U6633 (N_6633,N_6596,N_6551);
nor U6634 (N_6634,N_6409,N_6495);
or U6635 (N_6635,N_6503,N_6537);
nand U6636 (N_6636,N_6525,N_6462);
or U6637 (N_6637,N_6553,N_6423);
nand U6638 (N_6638,N_6404,N_6413);
and U6639 (N_6639,N_6416,N_6488);
and U6640 (N_6640,N_6578,N_6441);
and U6641 (N_6641,N_6569,N_6405);
nand U6642 (N_6642,N_6479,N_6505);
nand U6643 (N_6643,N_6456,N_6550);
or U6644 (N_6644,N_6592,N_6476);
nor U6645 (N_6645,N_6588,N_6579);
or U6646 (N_6646,N_6510,N_6521);
and U6647 (N_6647,N_6585,N_6561);
xnor U6648 (N_6648,N_6567,N_6460);
nor U6649 (N_6649,N_6410,N_6565);
nor U6650 (N_6650,N_6470,N_6457);
xor U6651 (N_6651,N_6540,N_6464);
nand U6652 (N_6652,N_6402,N_6415);
xnor U6653 (N_6653,N_6582,N_6527);
nand U6654 (N_6654,N_6436,N_6449);
nor U6655 (N_6655,N_6474,N_6443);
or U6656 (N_6656,N_6555,N_6411);
or U6657 (N_6657,N_6534,N_6549);
nor U6658 (N_6658,N_6492,N_6453);
or U6659 (N_6659,N_6587,N_6403);
nand U6660 (N_6660,N_6401,N_6467);
and U6661 (N_6661,N_6463,N_6498);
and U6662 (N_6662,N_6589,N_6434);
and U6663 (N_6663,N_6574,N_6538);
or U6664 (N_6664,N_6501,N_6581);
or U6665 (N_6665,N_6426,N_6520);
or U6666 (N_6666,N_6556,N_6483);
or U6667 (N_6667,N_6513,N_6530);
xor U6668 (N_6668,N_6473,N_6429);
and U6669 (N_6669,N_6535,N_6430);
xnor U6670 (N_6670,N_6448,N_6566);
nor U6671 (N_6671,N_6526,N_6580);
or U6672 (N_6672,N_6591,N_6594);
nand U6673 (N_6673,N_6472,N_6595);
and U6674 (N_6674,N_6425,N_6451);
nand U6675 (N_6675,N_6543,N_6433);
nor U6676 (N_6676,N_6461,N_6516);
nand U6677 (N_6677,N_6452,N_6458);
and U6678 (N_6678,N_6428,N_6414);
nand U6679 (N_6679,N_6447,N_6573);
nand U6680 (N_6680,N_6420,N_6559);
nand U6681 (N_6681,N_6572,N_6471);
or U6682 (N_6682,N_6547,N_6442);
nand U6683 (N_6683,N_6412,N_6564);
xnor U6684 (N_6684,N_6511,N_6506);
xor U6685 (N_6685,N_6542,N_6558);
or U6686 (N_6686,N_6593,N_6422);
or U6687 (N_6687,N_6484,N_6519);
nand U6688 (N_6688,N_6548,N_6571);
or U6689 (N_6689,N_6491,N_6468);
or U6690 (N_6690,N_6584,N_6576);
xnor U6691 (N_6691,N_6529,N_6598);
or U6692 (N_6692,N_6490,N_6496);
nor U6693 (N_6693,N_6514,N_6562);
and U6694 (N_6694,N_6493,N_6528);
nand U6695 (N_6695,N_6454,N_6531);
xor U6696 (N_6696,N_6586,N_6504);
nor U6697 (N_6697,N_6500,N_6546);
and U6698 (N_6698,N_6481,N_6477);
or U6699 (N_6699,N_6532,N_6408);
and U6700 (N_6700,N_6551,N_6500);
and U6701 (N_6701,N_6516,N_6467);
nor U6702 (N_6702,N_6438,N_6403);
xor U6703 (N_6703,N_6501,N_6518);
nor U6704 (N_6704,N_6559,N_6438);
or U6705 (N_6705,N_6553,N_6562);
xnor U6706 (N_6706,N_6417,N_6456);
xnor U6707 (N_6707,N_6504,N_6483);
or U6708 (N_6708,N_6471,N_6424);
or U6709 (N_6709,N_6568,N_6413);
nand U6710 (N_6710,N_6432,N_6440);
or U6711 (N_6711,N_6597,N_6430);
or U6712 (N_6712,N_6551,N_6408);
and U6713 (N_6713,N_6444,N_6433);
nor U6714 (N_6714,N_6500,N_6427);
xnor U6715 (N_6715,N_6489,N_6496);
and U6716 (N_6716,N_6482,N_6502);
xor U6717 (N_6717,N_6494,N_6544);
nor U6718 (N_6718,N_6435,N_6453);
nand U6719 (N_6719,N_6544,N_6560);
nor U6720 (N_6720,N_6419,N_6404);
or U6721 (N_6721,N_6465,N_6556);
and U6722 (N_6722,N_6556,N_6562);
and U6723 (N_6723,N_6555,N_6444);
nand U6724 (N_6724,N_6474,N_6541);
xor U6725 (N_6725,N_6525,N_6517);
nand U6726 (N_6726,N_6441,N_6571);
nor U6727 (N_6727,N_6449,N_6561);
nor U6728 (N_6728,N_6404,N_6472);
nor U6729 (N_6729,N_6411,N_6494);
xor U6730 (N_6730,N_6523,N_6532);
nand U6731 (N_6731,N_6507,N_6591);
nand U6732 (N_6732,N_6432,N_6454);
or U6733 (N_6733,N_6444,N_6400);
and U6734 (N_6734,N_6498,N_6421);
or U6735 (N_6735,N_6463,N_6580);
or U6736 (N_6736,N_6434,N_6407);
or U6737 (N_6737,N_6542,N_6597);
nor U6738 (N_6738,N_6412,N_6466);
nand U6739 (N_6739,N_6443,N_6468);
or U6740 (N_6740,N_6553,N_6493);
xor U6741 (N_6741,N_6522,N_6403);
nand U6742 (N_6742,N_6475,N_6411);
or U6743 (N_6743,N_6547,N_6566);
nand U6744 (N_6744,N_6480,N_6431);
nor U6745 (N_6745,N_6557,N_6555);
and U6746 (N_6746,N_6583,N_6466);
nor U6747 (N_6747,N_6475,N_6538);
or U6748 (N_6748,N_6414,N_6400);
or U6749 (N_6749,N_6571,N_6435);
xnor U6750 (N_6750,N_6400,N_6508);
nand U6751 (N_6751,N_6420,N_6565);
xor U6752 (N_6752,N_6574,N_6550);
or U6753 (N_6753,N_6575,N_6434);
or U6754 (N_6754,N_6512,N_6402);
nand U6755 (N_6755,N_6510,N_6542);
nor U6756 (N_6756,N_6437,N_6452);
nand U6757 (N_6757,N_6529,N_6586);
xor U6758 (N_6758,N_6433,N_6501);
or U6759 (N_6759,N_6470,N_6443);
nor U6760 (N_6760,N_6596,N_6564);
and U6761 (N_6761,N_6508,N_6503);
and U6762 (N_6762,N_6425,N_6589);
nor U6763 (N_6763,N_6437,N_6471);
or U6764 (N_6764,N_6511,N_6596);
and U6765 (N_6765,N_6540,N_6521);
or U6766 (N_6766,N_6581,N_6580);
or U6767 (N_6767,N_6455,N_6511);
xor U6768 (N_6768,N_6530,N_6592);
nor U6769 (N_6769,N_6544,N_6446);
nor U6770 (N_6770,N_6482,N_6423);
and U6771 (N_6771,N_6454,N_6541);
xor U6772 (N_6772,N_6407,N_6421);
xor U6773 (N_6773,N_6529,N_6572);
xor U6774 (N_6774,N_6429,N_6548);
or U6775 (N_6775,N_6550,N_6561);
nand U6776 (N_6776,N_6569,N_6538);
nand U6777 (N_6777,N_6584,N_6532);
xor U6778 (N_6778,N_6592,N_6454);
and U6779 (N_6779,N_6429,N_6438);
nor U6780 (N_6780,N_6504,N_6562);
or U6781 (N_6781,N_6594,N_6431);
xnor U6782 (N_6782,N_6492,N_6412);
xor U6783 (N_6783,N_6454,N_6416);
or U6784 (N_6784,N_6514,N_6556);
and U6785 (N_6785,N_6524,N_6545);
and U6786 (N_6786,N_6578,N_6532);
nor U6787 (N_6787,N_6427,N_6408);
or U6788 (N_6788,N_6549,N_6542);
xnor U6789 (N_6789,N_6439,N_6423);
nand U6790 (N_6790,N_6430,N_6454);
and U6791 (N_6791,N_6559,N_6501);
xor U6792 (N_6792,N_6516,N_6518);
nor U6793 (N_6793,N_6528,N_6524);
nand U6794 (N_6794,N_6516,N_6508);
and U6795 (N_6795,N_6556,N_6498);
xor U6796 (N_6796,N_6539,N_6438);
xor U6797 (N_6797,N_6478,N_6438);
and U6798 (N_6798,N_6460,N_6540);
or U6799 (N_6799,N_6411,N_6405);
xor U6800 (N_6800,N_6723,N_6726);
and U6801 (N_6801,N_6799,N_6622);
nand U6802 (N_6802,N_6651,N_6797);
and U6803 (N_6803,N_6618,N_6719);
nand U6804 (N_6804,N_6738,N_6714);
or U6805 (N_6805,N_6696,N_6706);
or U6806 (N_6806,N_6683,N_6785);
nor U6807 (N_6807,N_6774,N_6659);
and U6808 (N_6808,N_6675,N_6689);
xor U6809 (N_6809,N_6676,N_6761);
xor U6810 (N_6810,N_6750,N_6656);
nand U6811 (N_6811,N_6624,N_6710);
nor U6812 (N_6812,N_6602,N_6769);
nand U6813 (N_6813,N_6627,N_6679);
or U6814 (N_6814,N_6791,N_6678);
xor U6815 (N_6815,N_6768,N_6783);
xor U6816 (N_6816,N_6708,N_6741);
or U6817 (N_6817,N_6619,N_6691);
and U6818 (N_6818,N_6648,N_6729);
nor U6819 (N_6819,N_6647,N_6749);
nand U6820 (N_6820,N_6787,N_6636);
xnor U6821 (N_6821,N_6615,N_6788);
xnor U6822 (N_6822,N_6620,N_6645);
or U6823 (N_6823,N_6740,N_6649);
nand U6824 (N_6824,N_6668,N_6680);
or U6825 (N_6825,N_6767,N_6611);
nand U6826 (N_6826,N_6658,N_6784);
xor U6827 (N_6827,N_6746,N_6792);
xnor U6828 (N_6828,N_6600,N_6638);
or U6829 (N_6829,N_6661,N_6654);
nor U6830 (N_6830,N_6616,N_6662);
nand U6831 (N_6831,N_6730,N_6798);
and U6832 (N_6832,N_6709,N_6786);
nand U6833 (N_6833,N_6629,N_6663);
or U6834 (N_6834,N_6763,N_6694);
nand U6835 (N_6835,N_6736,N_6666);
or U6836 (N_6836,N_6695,N_6715);
or U6837 (N_6837,N_6707,N_6644);
or U6838 (N_6838,N_6742,N_6657);
nand U6839 (N_6839,N_6609,N_6630);
nand U6840 (N_6840,N_6725,N_6607);
xnor U6841 (N_6841,N_6720,N_6766);
xnor U6842 (N_6842,N_6665,N_6628);
nor U6843 (N_6843,N_6605,N_6664);
or U6844 (N_6844,N_6732,N_6617);
nand U6845 (N_6845,N_6603,N_6782);
nor U6846 (N_6846,N_6660,N_6608);
nor U6847 (N_6847,N_6751,N_6756);
xnor U6848 (N_6848,N_6671,N_6765);
or U6849 (N_6849,N_6634,N_6612);
and U6850 (N_6850,N_6743,N_6639);
xnor U6851 (N_6851,N_6686,N_6698);
xor U6852 (N_6852,N_6670,N_6745);
nand U6853 (N_6853,N_6739,N_6727);
and U6854 (N_6854,N_6758,N_6734);
or U6855 (N_6855,N_6684,N_6781);
or U6856 (N_6856,N_6633,N_6673);
xor U6857 (N_6857,N_6757,N_6753);
nand U6858 (N_6858,N_6655,N_6701);
nand U6859 (N_6859,N_6748,N_6712);
nor U6860 (N_6860,N_6772,N_6637);
or U6861 (N_6861,N_6704,N_6646);
and U6862 (N_6862,N_6718,N_6692);
and U6863 (N_6863,N_6631,N_6604);
nand U6864 (N_6864,N_6790,N_6737);
xor U6865 (N_6865,N_6653,N_6780);
nor U6866 (N_6866,N_6724,N_6735);
nand U6867 (N_6867,N_6764,N_6721);
nand U6868 (N_6868,N_6697,N_6793);
and U6869 (N_6869,N_6690,N_6652);
nor U6870 (N_6870,N_6667,N_6744);
or U6871 (N_6871,N_6601,N_6755);
or U6872 (N_6872,N_6747,N_6635);
xor U6873 (N_6873,N_6771,N_6632);
nand U6874 (N_6874,N_6703,N_6682);
and U6875 (N_6875,N_6794,N_6777);
xor U6876 (N_6876,N_6672,N_6669);
nor U6877 (N_6877,N_6702,N_6716);
nor U6878 (N_6878,N_6693,N_6681);
and U6879 (N_6879,N_6711,N_6687);
nand U6880 (N_6880,N_6640,N_6677);
xor U6881 (N_6881,N_6625,N_6779);
and U6882 (N_6882,N_6775,N_6795);
or U6883 (N_6883,N_6713,N_6643);
and U6884 (N_6884,N_6688,N_6759);
xor U6885 (N_6885,N_6778,N_6650);
nor U6886 (N_6886,N_6623,N_6610);
or U6887 (N_6887,N_6642,N_6728);
nand U6888 (N_6888,N_6776,N_6614);
nand U6889 (N_6889,N_6626,N_6731);
nor U6890 (N_6890,N_6641,N_6717);
or U6891 (N_6891,N_6699,N_6705);
xnor U6892 (N_6892,N_6796,N_6621);
and U6893 (N_6893,N_6674,N_6700);
or U6894 (N_6894,N_6752,N_6773);
xnor U6895 (N_6895,N_6760,N_6770);
xor U6896 (N_6896,N_6606,N_6789);
xor U6897 (N_6897,N_6613,N_6762);
and U6898 (N_6898,N_6685,N_6722);
nor U6899 (N_6899,N_6733,N_6754);
nand U6900 (N_6900,N_6712,N_6702);
nand U6901 (N_6901,N_6630,N_6673);
or U6902 (N_6902,N_6751,N_6719);
xnor U6903 (N_6903,N_6698,N_6706);
nand U6904 (N_6904,N_6787,N_6644);
nor U6905 (N_6905,N_6637,N_6679);
nand U6906 (N_6906,N_6713,N_6723);
and U6907 (N_6907,N_6678,N_6662);
and U6908 (N_6908,N_6777,N_6751);
xnor U6909 (N_6909,N_6784,N_6747);
nand U6910 (N_6910,N_6629,N_6748);
nor U6911 (N_6911,N_6629,N_6650);
or U6912 (N_6912,N_6663,N_6706);
nor U6913 (N_6913,N_6651,N_6787);
or U6914 (N_6914,N_6726,N_6790);
nor U6915 (N_6915,N_6615,N_6743);
nand U6916 (N_6916,N_6692,N_6653);
nand U6917 (N_6917,N_6677,N_6724);
and U6918 (N_6918,N_6653,N_6796);
or U6919 (N_6919,N_6681,N_6723);
or U6920 (N_6920,N_6638,N_6653);
xor U6921 (N_6921,N_6681,N_6668);
and U6922 (N_6922,N_6679,N_6691);
nor U6923 (N_6923,N_6631,N_6695);
xnor U6924 (N_6924,N_6675,N_6657);
xor U6925 (N_6925,N_6621,N_6614);
nand U6926 (N_6926,N_6666,N_6763);
xnor U6927 (N_6927,N_6712,N_6744);
or U6928 (N_6928,N_6645,N_6771);
xnor U6929 (N_6929,N_6743,N_6793);
or U6930 (N_6930,N_6644,N_6672);
or U6931 (N_6931,N_6699,N_6629);
nand U6932 (N_6932,N_6647,N_6698);
nor U6933 (N_6933,N_6644,N_6637);
nand U6934 (N_6934,N_6773,N_6797);
or U6935 (N_6935,N_6653,N_6783);
xnor U6936 (N_6936,N_6663,N_6739);
or U6937 (N_6937,N_6701,N_6642);
nand U6938 (N_6938,N_6787,N_6721);
xor U6939 (N_6939,N_6710,N_6679);
nor U6940 (N_6940,N_6768,N_6619);
xnor U6941 (N_6941,N_6682,N_6619);
nor U6942 (N_6942,N_6666,N_6672);
and U6943 (N_6943,N_6773,N_6763);
and U6944 (N_6944,N_6782,N_6713);
or U6945 (N_6945,N_6689,N_6661);
nor U6946 (N_6946,N_6688,N_6656);
or U6947 (N_6947,N_6693,N_6611);
nand U6948 (N_6948,N_6797,N_6603);
or U6949 (N_6949,N_6638,N_6711);
and U6950 (N_6950,N_6645,N_6790);
and U6951 (N_6951,N_6797,N_6770);
nand U6952 (N_6952,N_6686,N_6756);
or U6953 (N_6953,N_6673,N_6784);
and U6954 (N_6954,N_6753,N_6765);
xor U6955 (N_6955,N_6670,N_6774);
nand U6956 (N_6956,N_6758,N_6746);
and U6957 (N_6957,N_6775,N_6617);
nand U6958 (N_6958,N_6621,N_6667);
and U6959 (N_6959,N_6747,N_6621);
nand U6960 (N_6960,N_6663,N_6746);
xnor U6961 (N_6961,N_6722,N_6782);
and U6962 (N_6962,N_6626,N_6732);
nor U6963 (N_6963,N_6675,N_6679);
and U6964 (N_6964,N_6640,N_6780);
and U6965 (N_6965,N_6677,N_6636);
xnor U6966 (N_6966,N_6639,N_6669);
or U6967 (N_6967,N_6702,N_6658);
nor U6968 (N_6968,N_6718,N_6768);
and U6969 (N_6969,N_6780,N_6786);
or U6970 (N_6970,N_6767,N_6781);
nand U6971 (N_6971,N_6794,N_6747);
nor U6972 (N_6972,N_6709,N_6730);
nand U6973 (N_6973,N_6714,N_6656);
xor U6974 (N_6974,N_6768,N_6763);
nor U6975 (N_6975,N_6657,N_6654);
nor U6976 (N_6976,N_6603,N_6724);
nor U6977 (N_6977,N_6775,N_6735);
and U6978 (N_6978,N_6684,N_6735);
nand U6979 (N_6979,N_6785,N_6786);
and U6980 (N_6980,N_6653,N_6642);
or U6981 (N_6981,N_6606,N_6652);
nand U6982 (N_6982,N_6671,N_6700);
nor U6983 (N_6983,N_6698,N_6601);
nor U6984 (N_6984,N_6769,N_6615);
nor U6985 (N_6985,N_6604,N_6651);
xnor U6986 (N_6986,N_6697,N_6784);
xnor U6987 (N_6987,N_6625,N_6743);
or U6988 (N_6988,N_6642,N_6698);
or U6989 (N_6989,N_6628,N_6688);
and U6990 (N_6990,N_6766,N_6699);
xor U6991 (N_6991,N_6791,N_6668);
nor U6992 (N_6992,N_6602,N_6660);
nand U6993 (N_6993,N_6627,N_6701);
nor U6994 (N_6994,N_6627,N_6751);
nor U6995 (N_6995,N_6633,N_6776);
nand U6996 (N_6996,N_6777,N_6681);
nor U6997 (N_6997,N_6708,N_6632);
nand U6998 (N_6998,N_6672,N_6638);
nand U6999 (N_6999,N_6712,N_6650);
nor U7000 (N_7000,N_6920,N_6835);
and U7001 (N_7001,N_6857,N_6867);
nand U7002 (N_7002,N_6912,N_6845);
or U7003 (N_7003,N_6931,N_6900);
and U7004 (N_7004,N_6877,N_6975);
nor U7005 (N_7005,N_6914,N_6910);
nand U7006 (N_7006,N_6947,N_6919);
nor U7007 (N_7007,N_6979,N_6959);
or U7008 (N_7008,N_6834,N_6872);
and U7009 (N_7009,N_6941,N_6879);
xor U7010 (N_7010,N_6952,N_6842);
nor U7011 (N_7011,N_6820,N_6862);
nand U7012 (N_7012,N_6921,N_6812);
nand U7013 (N_7013,N_6936,N_6897);
and U7014 (N_7014,N_6996,N_6930);
nand U7015 (N_7015,N_6839,N_6894);
and U7016 (N_7016,N_6837,N_6932);
nor U7017 (N_7017,N_6859,N_6871);
and U7018 (N_7018,N_6822,N_6965);
or U7019 (N_7019,N_6966,N_6805);
xor U7020 (N_7020,N_6808,N_6810);
xnor U7021 (N_7021,N_6831,N_6978);
nand U7022 (N_7022,N_6998,N_6824);
nand U7023 (N_7023,N_6861,N_6850);
and U7024 (N_7024,N_6991,N_6823);
xnor U7025 (N_7025,N_6875,N_6880);
nand U7026 (N_7026,N_6816,N_6899);
xor U7027 (N_7027,N_6818,N_6889);
nand U7028 (N_7028,N_6866,N_6939);
nand U7029 (N_7029,N_6985,N_6876);
xor U7030 (N_7030,N_6874,N_6892);
or U7031 (N_7031,N_6945,N_6869);
nand U7032 (N_7032,N_6934,N_6854);
and U7033 (N_7033,N_6986,N_6827);
xor U7034 (N_7034,N_6988,N_6977);
xnor U7035 (N_7035,N_6815,N_6883);
nor U7036 (N_7036,N_6951,N_6956);
and U7037 (N_7037,N_6911,N_6813);
or U7038 (N_7038,N_6963,N_6992);
and U7039 (N_7039,N_6830,N_6851);
and U7040 (N_7040,N_6961,N_6846);
nor U7041 (N_7041,N_6925,N_6873);
nor U7042 (N_7042,N_6960,N_6974);
nand U7043 (N_7043,N_6888,N_6980);
nand U7044 (N_7044,N_6895,N_6848);
nand U7045 (N_7045,N_6942,N_6968);
or U7046 (N_7046,N_6949,N_6967);
xor U7047 (N_7047,N_6887,N_6800);
nand U7048 (N_7048,N_6863,N_6946);
nor U7049 (N_7049,N_6817,N_6964);
xor U7050 (N_7050,N_6806,N_6804);
nor U7051 (N_7051,N_6913,N_6994);
or U7052 (N_7052,N_6836,N_6864);
nand U7053 (N_7053,N_6807,N_6896);
nand U7054 (N_7054,N_6999,N_6907);
nand U7055 (N_7055,N_6915,N_6844);
nor U7056 (N_7056,N_6937,N_6981);
nand U7057 (N_7057,N_6924,N_6971);
or U7058 (N_7058,N_6860,N_6840);
xnor U7059 (N_7059,N_6908,N_6833);
or U7060 (N_7060,N_6909,N_6809);
nand U7061 (N_7061,N_6898,N_6893);
xor U7062 (N_7062,N_6922,N_6841);
nor U7063 (N_7063,N_6995,N_6878);
or U7064 (N_7064,N_6955,N_6825);
nor U7065 (N_7065,N_6917,N_6870);
or U7066 (N_7066,N_6828,N_6987);
nand U7067 (N_7067,N_6928,N_6997);
nor U7068 (N_7068,N_6856,N_6940);
xnor U7069 (N_7069,N_6927,N_6802);
nor U7070 (N_7070,N_6935,N_6847);
nand U7071 (N_7071,N_6826,N_6821);
or U7072 (N_7072,N_6906,N_6918);
nand U7073 (N_7073,N_6904,N_6972);
nor U7074 (N_7074,N_6969,N_6948);
nor U7075 (N_7075,N_6916,N_6853);
xor U7076 (N_7076,N_6957,N_6953);
or U7077 (N_7077,N_6838,N_6881);
nand U7078 (N_7078,N_6882,N_6929);
nand U7079 (N_7079,N_6885,N_6843);
and U7080 (N_7080,N_6868,N_6970);
and U7081 (N_7081,N_6829,N_6886);
nor U7082 (N_7082,N_6944,N_6819);
or U7083 (N_7083,N_6903,N_6950);
xnor U7084 (N_7084,N_6855,N_6990);
xnor U7085 (N_7085,N_6938,N_6803);
and U7086 (N_7086,N_6962,N_6958);
or U7087 (N_7087,N_6943,N_6905);
nand U7088 (N_7088,N_6801,N_6926);
xor U7089 (N_7089,N_6954,N_6993);
and U7090 (N_7090,N_6852,N_6976);
and U7091 (N_7091,N_6811,N_6849);
and U7092 (N_7092,N_6858,N_6865);
nand U7093 (N_7093,N_6814,N_6901);
and U7094 (N_7094,N_6933,N_6989);
or U7095 (N_7095,N_6983,N_6984);
or U7096 (N_7096,N_6923,N_6902);
nor U7097 (N_7097,N_6973,N_6891);
nor U7098 (N_7098,N_6890,N_6832);
nor U7099 (N_7099,N_6982,N_6884);
xnor U7100 (N_7100,N_6991,N_6928);
nand U7101 (N_7101,N_6927,N_6949);
nand U7102 (N_7102,N_6808,N_6950);
nor U7103 (N_7103,N_6824,N_6883);
and U7104 (N_7104,N_6908,N_6869);
nor U7105 (N_7105,N_6847,N_6844);
and U7106 (N_7106,N_6978,N_6918);
nor U7107 (N_7107,N_6881,N_6872);
nand U7108 (N_7108,N_6967,N_6922);
nand U7109 (N_7109,N_6995,N_6874);
xnor U7110 (N_7110,N_6941,N_6901);
or U7111 (N_7111,N_6884,N_6886);
and U7112 (N_7112,N_6896,N_6965);
and U7113 (N_7113,N_6949,N_6920);
and U7114 (N_7114,N_6803,N_6996);
nor U7115 (N_7115,N_6830,N_6876);
xnor U7116 (N_7116,N_6973,N_6806);
nand U7117 (N_7117,N_6972,N_6873);
nand U7118 (N_7118,N_6947,N_6977);
and U7119 (N_7119,N_6870,N_6810);
nand U7120 (N_7120,N_6824,N_6982);
nor U7121 (N_7121,N_6812,N_6965);
and U7122 (N_7122,N_6879,N_6910);
xor U7123 (N_7123,N_6851,N_6958);
nand U7124 (N_7124,N_6803,N_6944);
nor U7125 (N_7125,N_6847,N_6866);
xnor U7126 (N_7126,N_6886,N_6985);
nor U7127 (N_7127,N_6955,N_6904);
nor U7128 (N_7128,N_6825,N_6849);
or U7129 (N_7129,N_6815,N_6948);
or U7130 (N_7130,N_6903,N_6913);
nand U7131 (N_7131,N_6989,N_6955);
or U7132 (N_7132,N_6941,N_6884);
or U7133 (N_7133,N_6983,N_6860);
nor U7134 (N_7134,N_6967,N_6849);
or U7135 (N_7135,N_6833,N_6958);
nor U7136 (N_7136,N_6957,N_6917);
nor U7137 (N_7137,N_6930,N_6920);
or U7138 (N_7138,N_6970,N_6801);
xor U7139 (N_7139,N_6906,N_6915);
nor U7140 (N_7140,N_6899,N_6852);
nand U7141 (N_7141,N_6844,N_6973);
or U7142 (N_7142,N_6997,N_6986);
or U7143 (N_7143,N_6918,N_6887);
xnor U7144 (N_7144,N_6958,N_6809);
xnor U7145 (N_7145,N_6839,N_6996);
xnor U7146 (N_7146,N_6955,N_6874);
nand U7147 (N_7147,N_6830,N_6948);
and U7148 (N_7148,N_6986,N_6862);
xnor U7149 (N_7149,N_6818,N_6867);
xor U7150 (N_7150,N_6942,N_6868);
and U7151 (N_7151,N_6853,N_6910);
and U7152 (N_7152,N_6937,N_6841);
xnor U7153 (N_7153,N_6898,N_6824);
or U7154 (N_7154,N_6873,N_6896);
xnor U7155 (N_7155,N_6811,N_6890);
xnor U7156 (N_7156,N_6904,N_6806);
xor U7157 (N_7157,N_6986,N_6970);
and U7158 (N_7158,N_6915,N_6837);
nand U7159 (N_7159,N_6963,N_6888);
and U7160 (N_7160,N_6920,N_6817);
and U7161 (N_7161,N_6997,N_6876);
nor U7162 (N_7162,N_6908,N_6921);
and U7163 (N_7163,N_6973,N_6830);
or U7164 (N_7164,N_6968,N_6932);
or U7165 (N_7165,N_6986,N_6907);
and U7166 (N_7166,N_6809,N_6974);
xor U7167 (N_7167,N_6853,N_6822);
or U7168 (N_7168,N_6803,N_6820);
nand U7169 (N_7169,N_6961,N_6874);
xnor U7170 (N_7170,N_6878,N_6968);
or U7171 (N_7171,N_6829,N_6872);
xor U7172 (N_7172,N_6813,N_6930);
xnor U7173 (N_7173,N_6966,N_6922);
xnor U7174 (N_7174,N_6979,N_6952);
or U7175 (N_7175,N_6908,N_6889);
and U7176 (N_7176,N_6847,N_6934);
xor U7177 (N_7177,N_6817,N_6879);
and U7178 (N_7178,N_6934,N_6999);
xnor U7179 (N_7179,N_6844,N_6800);
nor U7180 (N_7180,N_6968,N_6970);
and U7181 (N_7181,N_6974,N_6979);
nor U7182 (N_7182,N_6956,N_6816);
and U7183 (N_7183,N_6861,N_6928);
and U7184 (N_7184,N_6957,N_6819);
xnor U7185 (N_7185,N_6987,N_6892);
xnor U7186 (N_7186,N_6981,N_6956);
or U7187 (N_7187,N_6881,N_6837);
and U7188 (N_7188,N_6923,N_6919);
or U7189 (N_7189,N_6902,N_6854);
xnor U7190 (N_7190,N_6948,N_6881);
and U7191 (N_7191,N_6833,N_6801);
xnor U7192 (N_7192,N_6876,N_6877);
or U7193 (N_7193,N_6874,N_6993);
xor U7194 (N_7194,N_6840,N_6832);
nor U7195 (N_7195,N_6981,N_6869);
and U7196 (N_7196,N_6917,N_6923);
and U7197 (N_7197,N_6920,N_6868);
or U7198 (N_7198,N_6922,N_6837);
xnor U7199 (N_7199,N_6898,N_6909);
nor U7200 (N_7200,N_7173,N_7162);
and U7201 (N_7201,N_7095,N_7174);
and U7202 (N_7202,N_7104,N_7100);
and U7203 (N_7203,N_7134,N_7029);
nor U7204 (N_7204,N_7068,N_7098);
or U7205 (N_7205,N_7198,N_7096);
xor U7206 (N_7206,N_7151,N_7181);
nor U7207 (N_7207,N_7054,N_7111);
nand U7208 (N_7208,N_7031,N_7081);
xor U7209 (N_7209,N_7113,N_7086);
nor U7210 (N_7210,N_7088,N_7193);
or U7211 (N_7211,N_7144,N_7172);
and U7212 (N_7212,N_7101,N_7016);
xor U7213 (N_7213,N_7147,N_7012);
and U7214 (N_7214,N_7002,N_7003);
xnor U7215 (N_7215,N_7176,N_7056);
nor U7216 (N_7216,N_7126,N_7057);
xnor U7217 (N_7217,N_7155,N_7121);
and U7218 (N_7218,N_7059,N_7131);
nor U7219 (N_7219,N_7011,N_7123);
and U7220 (N_7220,N_7133,N_7149);
and U7221 (N_7221,N_7199,N_7037);
and U7222 (N_7222,N_7022,N_7175);
nand U7223 (N_7223,N_7132,N_7180);
xnor U7224 (N_7224,N_7072,N_7141);
nand U7225 (N_7225,N_7076,N_7116);
or U7226 (N_7226,N_7182,N_7156);
nand U7227 (N_7227,N_7046,N_7035);
nand U7228 (N_7228,N_7196,N_7118);
nor U7229 (N_7229,N_7148,N_7130);
xnor U7230 (N_7230,N_7032,N_7060);
and U7231 (N_7231,N_7167,N_7197);
nor U7232 (N_7232,N_7083,N_7119);
xor U7233 (N_7233,N_7129,N_7103);
or U7234 (N_7234,N_7023,N_7062);
xor U7235 (N_7235,N_7170,N_7106);
xor U7236 (N_7236,N_7179,N_7145);
xor U7237 (N_7237,N_7157,N_7138);
nand U7238 (N_7238,N_7108,N_7004);
nor U7239 (N_7239,N_7066,N_7027);
nand U7240 (N_7240,N_7073,N_7099);
or U7241 (N_7241,N_7093,N_7109);
nand U7242 (N_7242,N_7183,N_7028);
nor U7243 (N_7243,N_7077,N_7064);
or U7244 (N_7244,N_7114,N_7184);
xnor U7245 (N_7245,N_7122,N_7102);
and U7246 (N_7246,N_7191,N_7137);
xor U7247 (N_7247,N_7052,N_7140);
xnor U7248 (N_7248,N_7018,N_7110);
nor U7249 (N_7249,N_7007,N_7153);
xor U7250 (N_7250,N_7079,N_7047);
nand U7251 (N_7251,N_7034,N_7026);
nand U7252 (N_7252,N_7020,N_7120);
and U7253 (N_7253,N_7009,N_7014);
xnor U7254 (N_7254,N_7082,N_7069);
nand U7255 (N_7255,N_7165,N_7067);
xnor U7256 (N_7256,N_7041,N_7000);
and U7257 (N_7257,N_7063,N_7042);
nor U7258 (N_7258,N_7117,N_7136);
or U7259 (N_7259,N_7049,N_7158);
or U7260 (N_7260,N_7070,N_7115);
xor U7261 (N_7261,N_7127,N_7139);
nor U7262 (N_7262,N_7163,N_7024);
xnor U7263 (N_7263,N_7017,N_7154);
or U7264 (N_7264,N_7015,N_7159);
or U7265 (N_7265,N_7021,N_7005);
or U7266 (N_7266,N_7161,N_7089);
nor U7267 (N_7267,N_7178,N_7013);
xor U7268 (N_7268,N_7177,N_7045);
or U7269 (N_7269,N_7128,N_7053);
or U7270 (N_7270,N_7025,N_7010);
nand U7271 (N_7271,N_7164,N_7055);
nor U7272 (N_7272,N_7065,N_7074);
nor U7273 (N_7273,N_7087,N_7048);
nand U7274 (N_7274,N_7008,N_7143);
nand U7275 (N_7275,N_7125,N_7166);
nor U7276 (N_7276,N_7006,N_7186);
xnor U7277 (N_7277,N_7171,N_7189);
nand U7278 (N_7278,N_7192,N_7061);
and U7279 (N_7279,N_7080,N_7085);
nor U7280 (N_7280,N_7150,N_7188);
xnor U7281 (N_7281,N_7038,N_7160);
and U7282 (N_7282,N_7058,N_7040);
or U7283 (N_7283,N_7078,N_7043);
and U7284 (N_7284,N_7195,N_7124);
or U7285 (N_7285,N_7091,N_7097);
and U7286 (N_7286,N_7142,N_7135);
or U7287 (N_7287,N_7094,N_7107);
xor U7288 (N_7288,N_7185,N_7090);
xnor U7289 (N_7289,N_7033,N_7030);
xnor U7290 (N_7290,N_7169,N_7044);
nor U7291 (N_7291,N_7152,N_7019);
or U7292 (N_7292,N_7190,N_7001);
nor U7293 (N_7293,N_7039,N_7075);
and U7294 (N_7294,N_7112,N_7187);
and U7295 (N_7295,N_7084,N_7146);
or U7296 (N_7296,N_7050,N_7168);
nand U7297 (N_7297,N_7036,N_7071);
and U7298 (N_7298,N_7194,N_7051);
or U7299 (N_7299,N_7092,N_7105);
nand U7300 (N_7300,N_7080,N_7193);
nor U7301 (N_7301,N_7000,N_7155);
xnor U7302 (N_7302,N_7129,N_7033);
nor U7303 (N_7303,N_7058,N_7085);
and U7304 (N_7304,N_7186,N_7059);
xnor U7305 (N_7305,N_7190,N_7127);
nand U7306 (N_7306,N_7047,N_7196);
and U7307 (N_7307,N_7188,N_7111);
nor U7308 (N_7308,N_7092,N_7068);
nand U7309 (N_7309,N_7002,N_7137);
nand U7310 (N_7310,N_7064,N_7048);
xor U7311 (N_7311,N_7180,N_7043);
or U7312 (N_7312,N_7032,N_7075);
nor U7313 (N_7313,N_7090,N_7096);
xnor U7314 (N_7314,N_7020,N_7135);
or U7315 (N_7315,N_7049,N_7028);
or U7316 (N_7316,N_7000,N_7085);
and U7317 (N_7317,N_7195,N_7006);
nand U7318 (N_7318,N_7162,N_7064);
nor U7319 (N_7319,N_7166,N_7120);
xor U7320 (N_7320,N_7102,N_7160);
xor U7321 (N_7321,N_7061,N_7137);
and U7322 (N_7322,N_7007,N_7004);
or U7323 (N_7323,N_7037,N_7057);
nand U7324 (N_7324,N_7184,N_7174);
or U7325 (N_7325,N_7097,N_7123);
or U7326 (N_7326,N_7044,N_7113);
xnor U7327 (N_7327,N_7191,N_7174);
nor U7328 (N_7328,N_7191,N_7138);
nor U7329 (N_7329,N_7138,N_7137);
and U7330 (N_7330,N_7136,N_7006);
nor U7331 (N_7331,N_7126,N_7119);
and U7332 (N_7332,N_7152,N_7009);
xnor U7333 (N_7333,N_7043,N_7026);
xnor U7334 (N_7334,N_7144,N_7041);
nor U7335 (N_7335,N_7074,N_7161);
or U7336 (N_7336,N_7066,N_7004);
or U7337 (N_7337,N_7080,N_7189);
and U7338 (N_7338,N_7160,N_7039);
or U7339 (N_7339,N_7152,N_7094);
or U7340 (N_7340,N_7077,N_7101);
or U7341 (N_7341,N_7027,N_7188);
nor U7342 (N_7342,N_7101,N_7129);
and U7343 (N_7343,N_7135,N_7012);
nand U7344 (N_7344,N_7058,N_7019);
or U7345 (N_7345,N_7005,N_7013);
nand U7346 (N_7346,N_7056,N_7103);
nand U7347 (N_7347,N_7176,N_7034);
xnor U7348 (N_7348,N_7056,N_7140);
and U7349 (N_7349,N_7119,N_7104);
xnor U7350 (N_7350,N_7171,N_7030);
xor U7351 (N_7351,N_7169,N_7128);
nand U7352 (N_7352,N_7165,N_7130);
and U7353 (N_7353,N_7199,N_7183);
and U7354 (N_7354,N_7155,N_7159);
and U7355 (N_7355,N_7044,N_7069);
nand U7356 (N_7356,N_7172,N_7195);
and U7357 (N_7357,N_7100,N_7135);
xor U7358 (N_7358,N_7062,N_7154);
xnor U7359 (N_7359,N_7011,N_7147);
xor U7360 (N_7360,N_7054,N_7099);
or U7361 (N_7361,N_7163,N_7100);
nand U7362 (N_7362,N_7147,N_7104);
nand U7363 (N_7363,N_7134,N_7022);
and U7364 (N_7364,N_7154,N_7043);
nand U7365 (N_7365,N_7162,N_7063);
nand U7366 (N_7366,N_7000,N_7186);
or U7367 (N_7367,N_7066,N_7021);
and U7368 (N_7368,N_7166,N_7092);
xnor U7369 (N_7369,N_7125,N_7009);
nor U7370 (N_7370,N_7055,N_7016);
and U7371 (N_7371,N_7102,N_7045);
and U7372 (N_7372,N_7130,N_7069);
xnor U7373 (N_7373,N_7101,N_7085);
and U7374 (N_7374,N_7052,N_7038);
and U7375 (N_7375,N_7122,N_7049);
and U7376 (N_7376,N_7041,N_7069);
nor U7377 (N_7377,N_7092,N_7110);
nor U7378 (N_7378,N_7116,N_7059);
xor U7379 (N_7379,N_7114,N_7055);
or U7380 (N_7380,N_7015,N_7022);
nand U7381 (N_7381,N_7068,N_7152);
nand U7382 (N_7382,N_7100,N_7015);
xor U7383 (N_7383,N_7165,N_7045);
or U7384 (N_7384,N_7161,N_7050);
nand U7385 (N_7385,N_7163,N_7113);
nand U7386 (N_7386,N_7103,N_7105);
nor U7387 (N_7387,N_7013,N_7105);
or U7388 (N_7388,N_7048,N_7103);
nand U7389 (N_7389,N_7068,N_7168);
xnor U7390 (N_7390,N_7036,N_7171);
nor U7391 (N_7391,N_7047,N_7048);
xnor U7392 (N_7392,N_7090,N_7117);
nor U7393 (N_7393,N_7109,N_7139);
nor U7394 (N_7394,N_7134,N_7069);
nor U7395 (N_7395,N_7151,N_7052);
xor U7396 (N_7396,N_7143,N_7004);
or U7397 (N_7397,N_7087,N_7187);
and U7398 (N_7398,N_7013,N_7048);
or U7399 (N_7399,N_7066,N_7069);
nand U7400 (N_7400,N_7230,N_7334);
nor U7401 (N_7401,N_7381,N_7300);
and U7402 (N_7402,N_7345,N_7255);
nand U7403 (N_7403,N_7353,N_7214);
xnor U7404 (N_7404,N_7307,N_7327);
xor U7405 (N_7405,N_7321,N_7217);
nand U7406 (N_7406,N_7212,N_7236);
nor U7407 (N_7407,N_7383,N_7318);
or U7408 (N_7408,N_7280,N_7365);
or U7409 (N_7409,N_7283,N_7380);
xnor U7410 (N_7410,N_7223,N_7256);
xnor U7411 (N_7411,N_7225,N_7397);
or U7412 (N_7412,N_7257,N_7332);
or U7413 (N_7413,N_7314,N_7267);
nand U7414 (N_7414,N_7388,N_7316);
or U7415 (N_7415,N_7277,N_7398);
nor U7416 (N_7416,N_7363,N_7385);
or U7417 (N_7417,N_7343,N_7295);
or U7418 (N_7418,N_7200,N_7292);
nand U7419 (N_7419,N_7320,N_7370);
or U7420 (N_7420,N_7352,N_7358);
nand U7421 (N_7421,N_7306,N_7279);
and U7422 (N_7422,N_7243,N_7245);
nand U7423 (N_7423,N_7325,N_7261);
nand U7424 (N_7424,N_7297,N_7204);
nor U7425 (N_7425,N_7241,N_7342);
or U7426 (N_7426,N_7284,N_7310);
nand U7427 (N_7427,N_7260,N_7235);
and U7428 (N_7428,N_7369,N_7250);
xor U7429 (N_7429,N_7382,N_7226);
and U7430 (N_7430,N_7244,N_7216);
xor U7431 (N_7431,N_7289,N_7364);
nor U7432 (N_7432,N_7251,N_7351);
nor U7433 (N_7433,N_7268,N_7228);
nand U7434 (N_7434,N_7312,N_7207);
or U7435 (N_7435,N_7227,N_7340);
and U7436 (N_7436,N_7341,N_7220);
nor U7437 (N_7437,N_7391,N_7390);
or U7438 (N_7438,N_7324,N_7311);
xnor U7439 (N_7439,N_7273,N_7329);
nand U7440 (N_7440,N_7309,N_7288);
nand U7441 (N_7441,N_7269,N_7221);
nand U7442 (N_7442,N_7252,N_7202);
nor U7443 (N_7443,N_7265,N_7215);
and U7444 (N_7444,N_7330,N_7258);
xor U7445 (N_7445,N_7360,N_7234);
xor U7446 (N_7446,N_7337,N_7387);
xor U7447 (N_7447,N_7331,N_7304);
or U7448 (N_7448,N_7237,N_7264);
nand U7449 (N_7449,N_7394,N_7285);
or U7450 (N_7450,N_7368,N_7246);
nor U7451 (N_7451,N_7208,N_7378);
nand U7452 (N_7452,N_7308,N_7272);
xor U7453 (N_7453,N_7287,N_7354);
or U7454 (N_7454,N_7373,N_7395);
or U7455 (N_7455,N_7282,N_7286);
or U7456 (N_7456,N_7278,N_7274);
or U7457 (N_7457,N_7384,N_7294);
xor U7458 (N_7458,N_7386,N_7305);
nand U7459 (N_7459,N_7393,N_7291);
nor U7460 (N_7460,N_7339,N_7302);
nand U7461 (N_7461,N_7259,N_7242);
xnor U7462 (N_7462,N_7347,N_7233);
nand U7463 (N_7463,N_7344,N_7356);
nor U7464 (N_7464,N_7224,N_7366);
or U7465 (N_7465,N_7239,N_7262);
xor U7466 (N_7466,N_7263,N_7350);
xor U7467 (N_7467,N_7315,N_7323);
nor U7468 (N_7468,N_7338,N_7293);
and U7469 (N_7469,N_7317,N_7371);
or U7470 (N_7470,N_7335,N_7203);
or U7471 (N_7471,N_7375,N_7361);
xnor U7472 (N_7472,N_7290,N_7222);
and U7473 (N_7473,N_7201,N_7299);
or U7474 (N_7474,N_7376,N_7362);
xnor U7475 (N_7475,N_7248,N_7298);
and U7476 (N_7476,N_7328,N_7336);
nor U7477 (N_7477,N_7379,N_7389);
and U7478 (N_7478,N_7367,N_7205);
and U7479 (N_7479,N_7253,N_7206);
xor U7480 (N_7480,N_7254,N_7213);
and U7481 (N_7481,N_7349,N_7218);
xnor U7482 (N_7482,N_7240,N_7301);
or U7483 (N_7483,N_7333,N_7275);
or U7484 (N_7484,N_7281,N_7210);
nand U7485 (N_7485,N_7238,N_7232);
nand U7486 (N_7486,N_7322,N_7296);
nor U7487 (N_7487,N_7249,N_7271);
and U7488 (N_7488,N_7326,N_7392);
nor U7489 (N_7489,N_7355,N_7276);
xnor U7490 (N_7490,N_7247,N_7374);
xor U7491 (N_7491,N_7211,N_7319);
and U7492 (N_7492,N_7396,N_7219);
xor U7493 (N_7493,N_7377,N_7229);
nor U7494 (N_7494,N_7313,N_7270);
xnor U7495 (N_7495,N_7303,N_7372);
nand U7496 (N_7496,N_7346,N_7266);
nor U7497 (N_7497,N_7348,N_7209);
xnor U7498 (N_7498,N_7357,N_7359);
xor U7499 (N_7499,N_7399,N_7231);
xnor U7500 (N_7500,N_7213,N_7342);
and U7501 (N_7501,N_7296,N_7316);
nor U7502 (N_7502,N_7272,N_7302);
and U7503 (N_7503,N_7363,N_7334);
nor U7504 (N_7504,N_7271,N_7201);
or U7505 (N_7505,N_7234,N_7311);
or U7506 (N_7506,N_7213,N_7287);
and U7507 (N_7507,N_7264,N_7218);
nand U7508 (N_7508,N_7360,N_7292);
nor U7509 (N_7509,N_7270,N_7275);
xor U7510 (N_7510,N_7265,N_7231);
nor U7511 (N_7511,N_7368,N_7276);
nand U7512 (N_7512,N_7368,N_7242);
nand U7513 (N_7513,N_7212,N_7211);
or U7514 (N_7514,N_7359,N_7259);
nand U7515 (N_7515,N_7209,N_7276);
xnor U7516 (N_7516,N_7332,N_7216);
nand U7517 (N_7517,N_7309,N_7326);
nor U7518 (N_7518,N_7355,N_7364);
or U7519 (N_7519,N_7324,N_7250);
and U7520 (N_7520,N_7345,N_7297);
and U7521 (N_7521,N_7335,N_7240);
nand U7522 (N_7522,N_7213,N_7241);
xor U7523 (N_7523,N_7220,N_7396);
xor U7524 (N_7524,N_7368,N_7305);
and U7525 (N_7525,N_7336,N_7300);
or U7526 (N_7526,N_7283,N_7379);
xor U7527 (N_7527,N_7232,N_7305);
xor U7528 (N_7528,N_7288,N_7222);
xor U7529 (N_7529,N_7264,N_7242);
xnor U7530 (N_7530,N_7346,N_7395);
and U7531 (N_7531,N_7353,N_7382);
nand U7532 (N_7532,N_7342,N_7376);
or U7533 (N_7533,N_7213,N_7297);
nand U7534 (N_7534,N_7266,N_7261);
and U7535 (N_7535,N_7349,N_7201);
nand U7536 (N_7536,N_7365,N_7289);
nor U7537 (N_7537,N_7247,N_7337);
nor U7538 (N_7538,N_7242,N_7372);
nor U7539 (N_7539,N_7387,N_7217);
or U7540 (N_7540,N_7390,N_7307);
nor U7541 (N_7541,N_7246,N_7256);
xnor U7542 (N_7542,N_7260,N_7270);
xor U7543 (N_7543,N_7385,N_7299);
and U7544 (N_7544,N_7233,N_7362);
nand U7545 (N_7545,N_7274,N_7344);
nand U7546 (N_7546,N_7320,N_7303);
xor U7547 (N_7547,N_7275,N_7226);
and U7548 (N_7548,N_7237,N_7311);
nand U7549 (N_7549,N_7319,N_7349);
xnor U7550 (N_7550,N_7234,N_7335);
and U7551 (N_7551,N_7323,N_7260);
xor U7552 (N_7552,N_7208,N_7277);
xor U7553 (N_7553,N_7228,N_7360);
and U7554 (N_7554,N_7235,N_7275);
xnor U7555 (N_7555,N_7207,N_7239);
or U7556 (N_7556,N_7254,N_7205);
nor U7557 (N_7557,N_7233,N_7392);
or U7558 (N_7558,N_7386,N_7266);
and U7559 (N_7559,N_7296,N_7330);
and U7560 (N_7560,N_7350,N_7278);
nor U7561 (N_7561,N_7325,N_7290);
nand U7562 (N_7562,N_7290,N_7302);
and U7563 (N_7563,N_7298,N_7263);
nor U7564 (N_7564,N_7305,N_7277);
nand U7565 (N_7565,N_7229,N_7288);
nand U7566 (N_7566,N_7352,N_7367);
nor U7567 (N_7567,N_7303,N_7205);
and U7568 (N_7568,N_7243,N_7285);
and U7569 (N_7569,N_7357,N_7361);
nor U7570 (N_7570,N_7360,N_7226);
xnor U7571 (N_7571,N_7351,N_7307);
nor U7572 (N_7572,N_7239,N_7350);
or U7573 (N_7573,N_7266,N_7302);
nor U7574 (N_7574,N_7202,N_7374);
and U7575 (N_7575,N_7283,N_7390);
or U7576 (N_7576,N_7208,N_7393);
nor U7577 (N_7577,N_7258,N_7379);
and U7578 (N_7578,N_7213,N_7262);
xor U7579 (N_7579,N_7300,N_7312);
nor U7580 (N_7580,N_7340,N_7360);
nor U7581 (N_7581,N_7214,N_7303);
and U7582 (N_7582,N_7262,N_7299);
or U7583 (N_7583,N_7272,N_7379);
xor U7584 (N_7584,N_7339,N_7281);
or U7585 (N_7585,N_7339,N_7381);
nand U7586 (N_7586,N_7330,N_7246);
and U7587 (N_7587,N_7260,N_7326);
and U7588 (N_7588,N_7364,N_7383);
xor U7589 (N_7589,N_7281,N_7200);
or U7590 (N_7590,N_7216,N_7369);
nor U7591 (N_7591,N_7205,N_7342);
nand U7592 (N_7592,N_7269,N_7298);
xor U7593 (N_7593,N_7254,N_7220);
and U7594 (N_7594,N_7224,N_7212);
and U7595 (N_7595,N_7397,N_7267);
or U7596 (N_7596,N_7318,N_7269);
nor U7597 (N_7597,N_7319,N_7255);
xnor U7598 (N_7598,N_7272,N_7370);
xnor U7599 (N_7599,N_7297,N_7397);
nand U7600 (N_7600,N_7581,N_7528);
xor U7601 (N_7601,N_7427,N_7550);
and U7602 (N_7602,N_7494,N_7569);
xnor U7603 (N_7603,N_7454,N_7442);
or U7604 (N_7604,N_7503,N_7456);
and U7605 (N_7605,N_7546,N_7457);
xnor U7606 (N_7606,N_7598,N_7478);
and U7607 (N_7607,N_7507,N_7439);
and U7608 (N_7608,N_7531,N_7435);
xor U7609 (N_7609,N_7481,N_7539);
xor U7610 (N_7610,N_7558,N_7445);
nand U7611 (N_7611,N_7520,N_7412);
or U7612 (N_7612,N_7583,N_7575);
or U7613 (N_7613,N_7499,N_7580);
or U7614 (N_7614,N_7438,N_7477);
nor U7615 (N_7615,N_7405,N_7538);
nor U7616 (N_7616,N_7571,N_7408);
nand U7617 (N_7617,N_7429,N_7400);
nand U7618 (N_7618,N_7527,N_7555);
or U7619 (N_7619,N_7553,N_7534);
xnor U7620 (N_7620,N_7588,N_7417);
nand U7621 (N_7621,N_7488,N_7430);
xor U7622 (N_7622,N_7548,N_7515);
xnor U7623 (N_7623,N_7463,N_7498);
nor U7624 (N_7624,N_7492,N_7466);
or U7625 (N_7625,N_7495,N_7579);
or U7626 (N_7626,N_7532,N_7403);
or U7627 (N_7627,N_7423,N_7419);
nand U7628 (N_7628,N_7589,N_7522);
xor U7629 (N_7629,N_7563,N_7599);
or U7630 (N_7630,N_7414,N_7592);
or U7631 (N_7631,N_7535,N_7510);
nor U7632 (N_7632,N_7566,N_7491);
or U7633 (N_7633,N_7551,N_7446);
and U7634 (N_7634,N_7406,N_7501);
nand U7635 (N_7635,N_7505,N_7541);
xor U7636 (N_7636,N_7564,N_7542);
nand U7637 (N_7637,N_7497,N_7586);
and U7638 (N_7638,N_7493,N_7476);
and U7639 (N_7639,N_7432,N_7474);
xor U7640 (N_7640,N_7425,N_7426);
or U7641 (N_7641,N_7460,N_7594);
or U7642 (N_7642,N_7407,N_7565);
xor U7643 (N_7643,N_7422,N_7506);
nand U7644 (N_7644,N_7557,N_7473);
xor U7645 (N_7645,N_7573,N_7487);
and U7646 (N_7646,N_7468,N_7544);
nor U7647 (N_7647,N_7533,N_7574);
xor U7648 (N_7648,N_7461,N_7475);
and U7649 (N_7649,N_7496,N_7500);
xor U7650 (N_7650,N_7483,N_7511);
and U7651 (N_7651,N_7570,N_7467);
nand U7652 (N_7652,N_7402,N_7521);
xnor U7653 (N_7653,N_7562,N_7469);
xor U7654 (N_7654,N_7458,N_7420);
xor U7655 (N_7655,N_7509,N_7428);
xnor U7656 (N_7656,N_7540,N_7587);
xnor U7657 (N_7657,N_7559,N_7448);
and U7658 (N_7658,N_7529,N_7443);
nand U7659 (N_7659,N_7591,N_7459);
nand U7660 (N_7660,N_7415,N_7421);
xor U7661 (N_7661,N_7582,N_7572);
nor U7662 (N_7662,N_7547,N_7449);
xor U7663 (N_7663,N_7537,N_7554);
nand U7664 (N_7664,N_7590,N_7595);
and U7665 (N_7665,N_7502,N_7513);
nand U7666 (N_7666,N_7447,N_7523);
nor U7667 (N_7667,N_7451,N_7525);
nor U7668 (N_7668,N_7441,N_7576);
and U7669 (N_7669,N_7455,N_7413);
or U7670 (N_7670,N_7404,N_7504);
nand U7671 (N_7671,N_7440,N_7470);
nand U7672 (N_7672,N_7536,N_7444);
nand U7673 (N_7673,N_7508,N_7519);
and U7674 (N_7674,N_7472,N_7484);
xor U7675 (N_7675,N_7479,N_7518);
xnor U7676 (N_7676,N_7482,N_7549);
nand U7677 (N_7677,N_7560,N_7433);
xor U7678 (N_7678,N_7489,N_7409);
nor U7679 (N_7679,N_7462,N_7567);
xor U7680 (N_7680,N_7486,N_7452);
nor U7681 (N_7681,N_7418,N_7585);
nor U7682 (N_7682,N_7512,N_7568);
and U7683 (N_7683,N_7524,N_7411);
xor U7684 (N_7684,N_7410,N_7577);
xor U7685 (N_7685,N_7437,N_7453);
nand U7686 (N_7686,N_7416,N_7561);
nand U7687 (N_7687,N_7593,N_7401);
or U7688 (N_7688,N_7552,N_7596);
nor U7689 (N_7689,N_7450,N_7436);
and U7690 (N_7690,N_7480,N_7464);
nor U7691 (N_7691,N_7556,N_7434);
or U7692 (N_7692,N_7545,N_7517);
nor U7693 (N_7693,N_7465,N_7584);
and U7694 (N_7694,N_7597,N_7543);
or U7695 (N_7695,N_7578,N_7526);
or U7696 (N_7696,N_7431,N_7424);
nor U7697 (N_7697,N_7514,N_7485);
nand U7698 (N_7698,N_7516,N_7471);
nand U7699 (N_7699,N_7530,N_7490);
nand U7700 (N_7700,N_7434,N_7479);
nor U7701 (N_7701,N_7483,N_7487);
nor U7702 (N_7702,N_7436,N_7534);
nand U7703 (N_7703,N_7571,N_7522);
and U7704 (N_7704,N_7591,N_7524);
nand U7705 (N_7705,N_7435,N_7488);
nor U7706 (N_7706,N_7528,N_7465);
nor U7707 (N_7707,N_7455,N_7446);
nand U7708 (N_7708,N_7407,N_7471);
and U7709 (N_7709,N_7425,N_7493);
nand U7710 (N_7710,N_7475,N_7520);
xor U7711 (N_7711,N_7444,N_7472);
or U7712 (N_7712,N_7559,N_7580);
nor U7713 (N_7713,N_7572,N_7577);
and U7714 (N_7714,N_7406,N_7478);
xor U7715 (N_7715,N_7480,N_7525);
and U7716 (N_7716,N_7536,N_7484);
and U7717 (N_7717,N_7579,N_7538);
and U7718 (N_7718,N_7494,N_7400);
nand U7719 (N_7719,N_7446,N_7423);
or U7720 (N_7720,N_7535,N_7539);
and U7721 (N_7721,N_7441,N_7578);
xor U7722 (N_7722,N_7582,N_7583);
xnor U7723 (N_7723,N_7540,N_7452);
nand U7724 (N_7724,N_7439,N_7568);
and U7725 (N_7725,N_7430,N_7570);
or U7726 (N_7726,N_7458,N_7536);
or U7727 (N_7727,N_7420,N_7412);
or U7728 (N_7728,N_7568,N_7466);
xnor U7729 (N_7729,N_7531,N_7579);
xor U7730 (N_7730,N_7422,N_7447);
nor U7731 (N_7731,N_7407,N_7526);
nor U7732 (N_7732,N_7585,N_7518);
xnor U7733 (N_7733,N_7442,N_7577);
and U7734 (N_7734,N_7401,N_7439);
or U7735 (N_7735,N_7428,N_7494);
nor U7736 (N_7736,N_7468,N_7542);
and U7737 (N_7737,N_7535,N_7455);
or U7738 (N_7738,N_7572,N_7535);
and U7739 (N_7739,N_7433,N_7417);
nor U7740 (N_7740,N_7483,N_7507);
or U7741 (N_7741,N_7471,N_7539);
or U7742 (N_7742,N_7458,N_7547);
or U7743 (N_7743,N_7470,N_7449);
xnor U7744 (N_7744,N_7515,N_7542);
xor U7745 (N_7745,N_7424,N_7530);
nand U7746 (N_7746,N_7575,N_7561);
xor U7747 (N_7747,N_7523,N_7588);
nand U7748 (N_7748,N_7506,N_7474);
and U7749 (N_7749,N_7412,N_7449);
or U7750 (N_7750,N_7565,N_7448);
nand U7751 (N_7751,N_7407,N_7505);
or U7752 (N_7752,N_7481,N_7543);
nor U7753 (N_7753,N_7560,N_7450);
or U7754 (N_7754,N_7578,N_7561);
nor U7755 (N_7755,N_7543,N_7440);
xnor U7756 (N_7756,N_7456,N_7519);
and U7757 (N_7757,N_7454,N_7587);
xnor U7758 (N_7758,N_7544,N_7568);
or U7759 (N_7759,N_7554,N_7435);
or U7760 (N_7760,N_7495,N_7490);
or U7761 (N_7761,N_7497,N_7498);
xnor U7762 (N_7762,N_7519,N_7488);
and U7763 (N_7763,N_7437,N_7520);
and U7764 (N_7764,N_7487,N_7544);
nor U7765 (N_7765,N_7434,N_7596);
and U7766 (N_7766,N_7571,N_7559);
xnor U7767 (N_7767,N_7478,N_7465);
and U7768 (N_7768,N_7509,N_7480);
or U7769 (N_7769,N_7421,N_7413);
and U7770 (N_7770,N_7547,N_7441);
nand U7771 (N_7771,N_7403,N_7474);
or U7772 (N_7772,N_7464,N_7563);
or U7773 (N_7773,N_7578,N_7493);
and U7774 (N_7774,N_7428,N_7411);
nand U7775 (N_7775,N_7524,N_7572);
nor U7776 (N_7776,N_7523,N_7476);
nor U7777 (N_7777,N_7541,N_7448);
nand U7778 (N_7778,N_7403,N_7498);
or U7779 (N_7779,N_7434,N_7511);
or U7780 (N_7780,N_7411,N_7562);
and U7781 (N_7781,N_7415,N_7471);
nand U7782 (N_7782,N_7447,N_7465);
xnor U7783 (N_7783,N_7571,N_7482);
and U7784 (N_7784,N_7529,N_7418);
xnor U7785 (N_7785,N_7414,N_7586);
and U7786 (N_7786,N_7439,N_7599);
nand U7787 (N_7787,N_7446,N_7450);
and U7788 (N_7788,N_7570,N_7478);
nand U7789 (N_7789,N_7508,N_7515);
nand U7790 (N_7790,N_7582,N_7597);
nand U7791 (N_7791,N_7534,N_7562);
and U7792 (N_7792,N_7596,N_7550);
xnor U7793 (N_7793,N_7572,N_7485);
nor U7794 (N_7794,N_7499,N_7430);
nand U7795 (N_7795,N_7431,N_7433);
or U7796 (N_7796,N_7403,N_7542);
nor U7797 (N_7797,N_7495,N_7413);
and U7798 (N_7798,N_7412,N_7544);
nand U7799 (N_7799,N_7526,N_7564);
or U7800 (N_7800,N_7657,N_7615);
nand U7801 (N_7801,N_7646,N_7711);
xnor U7802 (N_7802,N_7664,N_7747);
and U7803 (N_7803,N_7700,N_7710);
xnor U7804 (N_7804,N_7725,N_7652);
or U7805 (N_7805,N_7751,N_7608);
and U7806 (N_7806,N_7697,N_7783);
xor U7807 (N_7807,N_7784,N_7601);
xor U7808 (N_7808,N_7607,N_7739);
or U7809 (N_7809,N_7651,N_7758);
and U7810 (N_7810,N_7684,N_7754);
nand U7811 (N_7811,N_7663,N_7670);
nand U7812 (N_7812,N_7643,N_7775);
and U7813 (N_7813,N_7732,N_7715);
and U7814 (N_7814,N_7704,N_7685);
or U7815 (N_7815,N_7722,N_7666);
and U7816 (N_7816,N_7745,N_7617);
nor U7817 (N_7817,N_7658,N_7750);
or U7818 (N_7818,N_7777,N_7717);
nand U7819 (N_7819,N_7605,N_7609);
nor U7820 (N_7820,N_7671,N_7782);
or U7821 (N_7821,N_7629,N_7702);
or U7822 (N_7822,N_7641,N_7687);
and U7823 (N_7823,N_7659,N_7748);
and U7824 (N_7824,N_7699,N_7637);
and U7825 (N_7825,N_7741,N_7654);
or U7826 (N_7826,N_7786,N_7794);
nand U7827 (N_7827,N_7744,N_7735);
xor U7828 (N_7828,N_7721,N_7613);
or U7829 (N_7829,N_7708,N_7679);
and U7830 (N_7830,N_7639,N_7632);
nor U7831 (N_7831,N_7624,N_7619);
xor U7832 (N_7832,N_7650,N_7680);
nand U7833 (N_7833,N_7630,N_7698);
and U7834 (N_7834,N_7716,N_7764);
and U7835 (N_7835,N_7682,N_7628);
nand U7836 (N_7836,N_7738,N_7603);
and U7837 (N_7837,N_7713,N_7776);
xor U7838 (N_7838,N_7636,N_7719);
nor U7839 (N_7839,N_7771,N_7742);
xor U7840 (N_7840,N_7656,N_7648);
or U7841 (N_7841,N_7626,N_7755);
xor U7842 (N_7842,N_7737,N_7606);
or U7843 (N_7843,N_7779,N_7649);
xnor U7844 (N_7844,N_7778,N_7795);
or U7845 (N_7845,N_7672,N_7634);
and U7846 (N_7846,N_7665,N_7602);
and U7847 (N_7847,N_7757,N_7701);
and U7848 (N_7848,N_7785,N_7712);
xnor U7849 (N_7849,N_7780,N_7734);
nand U7850 (N_7850,N_7774,N_7787);
nor U7851 (N_7851,N_7733,N_7642);
and U7852 (N_7852,N_7767,N_7604);
and U7853 (N_7853,N_7789,N_7610);
and U7854 (N_7854,N_7611,N_7718);
xnor U7855 (N_7855,N_7727,N_7696);
nor U7856 (N_7856,N_7638,N_7724);
nor U7857 (N_7857,N_7761,N_7660);
and U7858 (N_7858,N_7668,N_7720);
nand U7859 (N_7859,N_7695,N_7614);
xor U7860 (N_7860,N_7683,N_7661);
or U7861 (N_7861,N_7769,N_7623);
or U7862 (N_7862,N_7692,N_7644);
or U7863 (N_7863,N_7690,N_7675);
nor U7864 (N_7864,N_7753,N_7798);
or U7865 (N_7865,N_7729,N_7706);
or U7866 (N_7866,N_7770,N_7686);
and U7867 (N_7867,N_7731,N_7625);
and U7868 (N_7868,N_7793,N_7612);
xnor U7869 (N_7869,N_7756,N_7796);
and U7870 (N_7870,N_7762,N_7691);
and U7871 (N_7871,N_7760,N_7620);
and U7872 (N_7872,N_7703,N_7730);
nor U7873 (N_7873,N_7631,N_7678);
nor U7874 (N_7874,N_7743,N_7788);
and U7875 (N_7875,N_7749,N_7709);
and U7876 (N_7876,N_7765,N_7726);
xnor U7877 (N_7877,N_7746,N_7674);
xor U7878 (N_7878,N_7673,N_7707);
or U7879 (N_7879,N_7677,N_7689);
nor U7880 (N_7880,N_7616,N_7752);
nand U7881 (N_7881,N_7600,N_7635);
and U7882 (N_7882,N_7766,N_7768);
xnor U7883 (N_7883,N_7633,N_7662);
and U7884 (N_7884,N_7681,N_7736);
nor U7885 (N_7885,N_7676,N_7790);
or U7886 (N_7886,N_7728,N_7799);
xnor U7887 (N_7887,N_7655,N_7645);
or U7888 (N_7888,N_7694,N_7781);
xor U7889 (N_7889,N_7669,N_7627);
xnor U7890 (N_7890,N_7773,N_7705);
nor U7891 (N_7891,N_7723,N_7618);
xnor U7892 (N_7892,N_7667,N_7791);
or U7893 (N_7893,N_7622,N_7792);
or U7894 (N_7894,N_7647,N_7772);
nor U7895 (N_7895,N_7740,N_7797);
xor U7896 (N_7896,N_7759,N_7688);
or U7897 (N_7897,N_7763,N_7621);
nor U7898 (N_7898,N_7693,N_7653);
nand U7899 (N_7899,N_7714,N_7640);
xor U7900 (N_7900,N_7601,N_7733);
or U7901 (N_7901,N_7673,N_7747);
or U7902 (N_7902,N_7790,N_7799);
or U7903 (N_7903,N_7758,N_7675);
and U7904 (N_7904,N_7618,N_7717);
xor U7905 (N_7905,N_7766,N_7727);
and U7906 (N_7906,N_7726,N_7616);
nor U7907 (N_7907,N_7636,N_7716);
nand U7908 (N_7908,N_7767,N_7700);
nand U7909 (N_7909,N_7707,N_7676);
or U7910 (N_7910,N_7748,N_7721);
nor U7911 (N_7911,N_7620,N_7610);
nor U7912 (N_7912,N_7780,N_7721);
nor U7913 (N_7913,N_7662,N_7787);
and U7914 (N_7914,N_7688,N_7662);
and U7915 (N_7915,N_7774,N_7697);
nand U7916 (N_7916,N_7638,N_7643);
xor U7917 (N_7917,N_7648,N_7617);
or U7918 (N_7918,N_7749,N_7694);
and U7919 (N_7919,N_7765,N_7625);
or U7920 (N_7920,N_7656,N_7794);
or U7921 (N_7921,N_7659,N_7640);
nand U7922 (N_7922,N_7691,N_7675);
or U7923 (N_7923,N_7665,N_7623);
or U7924 (N_7924,N_7696,N_7612);
or U7925 (N_7925,N_7657,N_7707);
or U7926 (N_7926,N_7763,N_7729);
nor U7927 (N_7927,N_7624,N_7600);
nor U7928 (N_7928,N_7675,N_7604);
nand U7929 (N_7929,N_7778,N_7763);
nand U7930 (N_7930,N_7640,N_7779);
and U7931 (N_7931,N_7658,N_7702);
and U7932 (N_7932,N_7743,N_7757);
and U7933 (N_7933,N_7660,N_7626);
and U7934 (N_7934,N_7782,N_7654);
or U7935 (N_7935,N_7799,N_7708);
or U7936 (N_7936,N_7650,N_7707);
nand U7937 (N_7937,N_7767,N_7772);
or U7938 (N_7938,N_7723,N_7765);
nand U7939 (N_7939,N_7600,N_7738);
or U7940 (N_7940,N_7608,N_7636);
nand U7941 (N_7941,N_7714,N_7628);
and U7942 (N_7942,N_7627,N_7683);
or U7943 (N_7943,N_7720,N_7601);
or U7944 (N_7944,N_7612,N_7779);
or U7945 (N_7945,N_7647,N_7625);
and U7946 (N_7946,N_7704,N_7663);
nand U7947 (N_7947,N_7603,N_7705);
nor U7948 (N_7948,N_7644,N_7705);
xor U7949 (N_7949,N_7611,N_7787);
or U7950 (N_7950,N_7653,N_7776);
and U7951 (N_7951,N_7718,N_7766);
xor U7952 (N_7952,N_7634,N_7756);
nand U7953 (N_7953,N_7700,N_7722);
or U7954 (N_7954,N_7724,N_7765);
nand U7955 (N_7955,N_7704,N_7717);
and U7956 (N_7956,N_7711,N_7647);
and U7957 (N_7957,N_7681,N_7639);
and U7958 (N_7958,N_7701,N_7737);
nand U7959 (N_7959,N_7671,N_7747);
nor U7960 (N_7960,N_7669,N_7637);
and U7961 (N_7961,N_7784,N_7661);
and U7962 (N_7962,N_7689,N_7670);
xnor U7963 (N_7963,N_7718,N_7699);
xor U7964 (N_7964,N_7613,N_7622);
and U7965 (N_7965,N_7607,N_7789);
and U7966 (N_7966,N_7692,N_7775);
nor U7967 (N_7967,N_7679,N_7652);
xnor U7968 (N_7968,N_7763,N_7625);
nor U7969 (N_7969,N_7723,N_7698);
and U7970 (N_7970,N_7725,N_7697);
xor U7971 (N_7971,N_7615,N_7662);
or U7972 (N_7972,N_7672,N_7787);
nand U7973 (N_7973,N_7772,N_7602);
nand U7974 (N_7974,N_7759,N_7735);
nand U7975 (N_7975,N_7768,N_7642);
xnor U7976 (N_7976,N_7707,N_7668);
xor U7977 (N_7977,N_7684,N_7698);
or U7978 (N_7978,N_7725,N_7672);
nand U7979 (N_7979,N_7632,N_7681);
nor U7980 (N_7980,N_7622,N_7658);
or U7981 (N_7981,N_7785,N_7717);
or U7982 (N_7982,N_7632,N_7666);
and U7983 (N_7983,N_7775,N_7701);
xnor U7984 (N_7984,N_7779,N_7615);
or U7985 (N_7985,N_7643,N_7791);
or U7986 (N_7986,N_7610,N_7768);
nor U7987 (N_7987,N_7707,N_7632);
nand U7988 (N_7988,N_7606,N_7784);
and U7989 (N_7989,N_7735,N_7714);
nand U7990 (N_7990,N_7604,N_7792);
or U7991 (N_7991,N_7701,N_7642);
nor U7992 (N_7992,N_7719,N_7670);
or U7993 (N_7993,N_7603,N_7663);
or U7994 (N_7994,N_7718,N_7694);
nand U7995 (N_7995,N_7785,N_7633);
or U7996 (N_7996,N_7788,N_7730);
and U7997 (N_7997,N_7642,N_7775);
and U7998 (N_7998,N_7614,N_7751);
or U7999 (N_7999,N_7620,N_7644);
or U8000 (N_8000,N_7923,N_7948);
xor U8001 (N_8001,N_7879,N_7941);
or U8002 (N_8002,N_7970,N_7969);
nor U8003 (N_8003,N_7915,N_7862);
nand U8004 (N_8004,N_7947,N_7940);
or U8005 (N_8005,N_7968,N_7839);
nand U8006 (N_8006,N_7921,N_7860);
xor U8007 (N_8007,N_7863,N_7861);
or U8008 (N_8008,N_7955,N_7815);
nand U8009 (N_8009,N_7820,N_7802);
nand U8010 (N_8010,N_7847,N_7909);
or U8011 (N_8011,N_7977,N_7823);
nand U8012 (N_8012,N_7856,N_7878);
or U8013 (N_8013,N_7900,N_7831);
nand U8014 (N_8014,N_7846,N_7890);
xor U8015 (N_8015,N_7876,N_7934);
xor U8016 (N_8016,N_7945,N_7953);
xor U8017 (N_8017,N_7907,N_7972);
nand U8018 (N_8018,N_7916,N_7819);
or U8019 (N_8019,N_7874,N_7931);
xnor U8020 (N_8020,N_7882,N_7918);
and U8021 (N_8021,N_7987,N_7816);
or U8022 (N_8022,N_7956,N_7985);
nor U8023 (N_8023,N_7999,N_7913);
and U8024 (N_8024,N_7949,N_7853);
and U8025 (N_8025,N_7952,N_7902);
nor U8026 (N_8026,N_7967,N_7929);
and U8027 (N_8027,N_7980,N_7858);
and U8028 (N_8028,N_7927,N_7801);
and U8029 (N_8029,N_7822,N_7933);
and U8030 (N_8030,N_7880,N_7895);
nand U8031 (N_8031,N_7988,N_7870);
or U8032 (N_8032,N_7854,N_7958);
nand U8033 (N_8033,N_7896,N_7982);
nand U8034 (N_8034,N_7964,N_7897);
or U8035 (N_8035,N_7946,N_7849);
or U8036 (N_8036,N_7959,N_7840);
or U8037 (N_8037,N_7836,N_7832);
or U8038 (N_8038,N_7981,N_7807);
xnor U8039 (N_8039,N_7919,N_7818);
and U8040 (N_8040,N_7997,N_7811);
xnor U8041 (N_8041,N_7965,N_7842);
nor U8042 (N_8042,N_7830,N_7996);
nor U8043 (N_8043,N_7838,N_7937);
or U8044 (N_8044,N_7912,N_7914);
and U8045 (N_8045,N_7932,N_7852);
nand U8046 (N_8046,N_7920,N_7859);
nand U8047 (N_8047,N_7814,N_7908);
and U8048 (N_8048,N_7930,N_7865);
or U8049 (N_8049,N_7800,N_7993);
xnor U8050 (N_8050,N_7877,N_7922);
nand U8051 (N_8051,N_7978,N_7813);
xnor U8052 (N_8052,N_7910,N_7867);
nor U8053 (N_8053,N_7808,N_7810);
nand U8054 (N_8054,N_7837,N_7973);
or U8055 (N_8055,N_7935,N_7826);
nor U8056 (N_8056,N_7827,N_7954);
nor U8057 (N_8057,N_7835,N_7841);
xor U8058 (N_8058,N_7950,N_7936);
nand U8059 (N_8059,N_7845,N_7989);
nor U8060 (N_8060,N_7975,N_7855);
nand U8061 (N_8061,N_7963,N_7986);
and U8062 (N_8062,N_7917,N_7809);
and U8063 (N_8063,N_7869,N_7848);
nand U8064 (N_8064,N_7928,N_7990);
nor U8065 (N_8065,N_7911,N_7873);
or U8066 (N_8066,N_7889,N_7817);
and U8067 (N_8067,N_7926,N_7992);
nand U8068 (N_8068,N_7979,N_7939);
and U8069 (N_8069,N_7904,N_7961);
nor U8070 (N_8070,N_7906,N_7957);
nand U8071 (N_8071,N_7850,N_7991);
nor U8072 (N_8072,N_7866,N_7943);
and U8073 (N_8073,N_7905,N_7899);
nor U8074 (N_8074,N_7884,N_7871);
nor U8075 (N_8075,N_7843,N_7888);
xor U8076 (N_8076,N_7892,N_7974);
nor U8077 (N_8077,N_7960,N_7925);
xnor U8078 (N_8078,N_7851,N_7883);
and U8079 (N_8079,N_7829,N_7872);
or U8080 (N_8080,N_7834,N_7891);
nand U8081 (N_8081,N_7966,N_7994);
or U8082 (N_8082,N_7875,N_7805);
xor U8083 (N_8083,N_7864,N_7868);
and U8084 (N_8084,N_7971,N_7844);
and U8085 (N_8085,N_7857,N_7803);
or U8086 (N_8086,N_7942,N_7806);
or U8087 (N_8087,N_7962,N_7995);
nor U8088 (N_8088,N_7825,N_7887);
nand U8089 (N_8089,N_7903,N_7828);
nand U8090 (N_8090,N_7821,N_7944);
xor U8091 (N_8091,N_7998,N_7924);
xor U8092 (N_8092,N_7984,N_7894);
nor U8093 (N_8093,N_7938,N_7886);
xnor U8094 (N_8094,N_7983,N_7804);
and U8095 (N_8095,N_7893,N_7885);
nand U8096 (N_8096,N_7824,N_7898);
nor U8097 (N_8097,N_7881,N_7812);
or U8098 (N_8098,N_7951,N_7833);
xnor U8099 (N_8099,N_7976,N_7901);
nand U8100 (N_8100,N_7807,N_7816);
nor U8101 (N_8101,N_7815,N_7979);
and U8102 (N_8102,N_7892,N_7841);
nor U8103 (N_8103,N_7997,N_7914);
and U8104 (N_8104,N_7952,N_7914);
and U8105 (N_8105,N_7844,N_7871);
xnor U8106 (N_8106,N_7823,N_7856);
and U8107 (N_8107,N_7925,N_7973);
nand U8108 (N_8108,N_7980,N_7891);
nand U8109 (N_8109,N_7942,N_7849);
nand U8110 (N_8110,N_7962,N_7986);
and U8111 (N_8111,N_7885,N_7986);
or U8112 (N_8112,N_7885,N_7808);
nor U8113 (N_8113,N_7956,N_7804);
xor U8114 (N_8114,N_7854,N_7897);
or U8115 (N_8115,N_7915,N_7876);
and U8116 (N_8116,N_7932,N_7934);
and U8117 (N_8117,N_7874,N_7832);
and U8118 (N_8118,N_7933,N_7962);
or U8119 (N_8119,N_7845,N_7875);
xnor U8120 (N_8120,N_7932,N_7809);
xnor U8121 (N_8121,N_7831,N_7972);
xor U8122 (N_8122,N_7875,N_7851);
nand U8123 (N_8123,N_7902,N_7954);
or U8124 (N_8124,N_7997,N_7841);
nand U8125 (N_8125,N_7932,N_7907);
nor U8126 (N_8126,N_7875,N_7823);
xor U8127 (N_8127,N_7820,N_7821);
and U8128 (N_8128,N_7864,N_7832);
and U8129 (N_8129,N_7881,N_7983);
and U8130 (N_8130,N_7878,N_7957);
or U8131 (N_8131,N_7876,N_7954);
xnor U8132 (N_8132,N_7983,N_7872);
nor U8133 (N_8133,N_7812,N_7967);
xnor U8134 (N_8134,N_7889,N_7882);
xor U8135 (N_8135,N_7960,N_7849);
nand U8136 (N_8136,N_7944,N_7972);
nand U8137 (N_8137,N_7930,N_7844);
or U8138 (N_8138,N_7873,N_7902);
xnor U8139 (N_8139,N_7825,N_7937);
nand U8140 (N_8140,N_7831,N_7887);
nand U8141 (N_8141,N_7902,N_7922);
or U8142 (N_8142,N_7954,N_7855);
xnor U8143 (N_8143,N_7914,N_7892);
nor U8144 (N_8144,N_7800,N_7814);
nor U8145 (N_8145,N_7821,N_7849);
nor U8146 (N_8146,N_7875,N_7859);
nand U8147 (N_8147,N_7958,N_7987);
and U8148 (N_8148,N_7992,N_7884);
nor U8149 (N_8149,N_7865,N_7868);
and U8150 (N_8150,N_7921,N_7873);
or U8151 (N_8151,N_7877,N_7897);
xnor U8152 (N_8152,N_7834,N_7870);
xnor U8153 (N_8153,N_7814,N_7989);
nor U8154 (N_8154,N_7874,N_7900);
and U8155 (N_8155,N_7980,N_7811);
nor U8156 (N_8156,N_7983,N_7977);
or U8157 (N_8157,N_7894,N_7844);
nor U8158 (N_8158,N_7874,N_7870);
and U8159 (N_8159,N_7992,N_7991);
and U8160 (N_8160,N_7981,N_7915);
nand U8161 (N_8161,N_7874,N_7871);
nand U8162 (N_8162,N_7986,N_7925);
nand U8163 (N_8163,N_7887,N_7808);
nor U8164 (N_8164,N_7958,N_7870);
or U8165 (N_8165,N_7870,N_7890);
nor U8166 (N_8166,N_7966,N_7856);
xor U8167 (N_8167,N_7824,N_7976);
xnor U8168 (N_8168,N_7829,N_7892);
nor U8169 (N_8169,N_7964,N_7821);
nor U8170 (N_8170,N_7845,N_7821);
nor U8171 (N_8171,N_7876,N_7944);
and U8172 (N_8172,N_7848,N_7980);
or U8173 (N_8173,N_7958,N_7976);
xor U8174 (N_8174,N_7909,N_7835);
or U8175 (N_8175,N_7882,N_7837);
and U8176 (N_8176,N_7871,N_7835);
nor U8177 (N_8177,N_7966,N_7926);
or U8178 (N_8178,N_7834,N_7907);
nand U8179 (N_8179,N_7915,N_7894);
nand U8180 (N_8180,N_7983,N_7924);
xnor U8181 (N_8181,N_7885,N_7902);
xnor U8182 (N_8182,N_7836,N_7885);
or U8183 (N_8183,N_7965,N_7884);
and U8184 (N_8184,N_7987,N_7972);
nand U8185 (N_8185,N_7959,N_7989);
and U8186 (N_8186,N_7855,N_7922);
and U8187 (N_8187,N_7925,N_7913);
and U8188 (N_8188,N_7946,N_7901);
xnor U8189 (N_8189,N_7803,N_7959);
or U8190 (N_8190,N_7998,N_7855);
and U8191 (N_8191,N_7991,N_7928);
xor U8192 (N_8192,N_7964,N_7995);
or U8193 (N_8193,N_7913,N_7839);
or U8194 (N_8194,N_7984,N_7806);
or U8195 (N_8195,N_7895,N_7818);
nand U8196 (N_8196,N_7982,N_7985);
and U8197 (N_8197,N_7909,N_7915);
and U8198 (N_8198,N_7901,N_7952);
nor U8199 (N_8199,N_7823,N_7910);
xor U8200 (N_8200,N_8091,N_8097);
xor U8201 (N_8201,N_8020,N_8189);
xnor U8202 (N_8202,N_8030,N_8100);
or U8203 (N_8203,N_8108,N_8149);
xnor U8204 (N_8204,N_8168,N_8199);
xor U8205 (N_8205,N_8043,N_8092);
or U8206 (N_8206,N_8154,N_8079);
nand U8207 (N_8207,N_8073,N_8031);
or U8208 (N_8208,N_8146,N_8006);
xnor U8209 (N_8209,N_8182,N_8038);
or U8210 (N_8210,N_8082,N_8160);
nor U8211 (N_8211,N_8106,N_8009);
xnor U8212 (N_8212,N_8128,N_8075);
nand U8213 (N_8213,N_8137,N_8187);
or U8214 (N_8214,N_8175,N_8174);
and U8215 (N_8215,N_8044,N_8081);
or U8216 (N_8216,N_8061,N_8041);
nor U8217 (N_8217,N_8156,N_8078);
xnor U8218 (N_8218,N_8164,N_8080);
nand U8219 (N_8219,N_8118,N_8172);
nand U8220 (N_8220,N_8028,N_8093);
or U8221 (N_8221,N_8089,N_8016);
nand U8222 (N_8222,N_8026,N_8011);
or U8223 (N_8223,N_8165,N_8067);
or U8224 (N_8224,N_8005,N_8166);
and U8225 (N_8225,N_8071,N_8003);
nor U8226 (N_8226,N_8138,N_8196);
and U8227 (N_8227,N_8099,N_8004);
nand U8228 (N_8228,N_8103,N_8125);
or U8229 (N_8229,N_8183,N_8008);
and U8230 (N_8230,N_8195,N_8062);
nor U8231 (N_8231,N_8054,N_8070);
nand U8232 (N_8232,N_8069,N_8135);
or U8233 (N_8233,N_8184,N_8169);
nand U8234 (N_8234,N_8139,N_8102);
nor U8235 (N_8235,N_8105,N_8007);
xnor U8236 (N_8236,N_8123,N_8143);
nand U8237 (N_8237,N_8052,N_8046);
nand U8238 (N_8238,N_8142,N_8136);
or U8239 (N_8239,N_8170,N_8173);
nand U8240 (N_8240,N_8059,N_8116);
or U8241 (N_8241,N_8163,N_8076);
nor U8242 (N_8242,N_8167,N_8001);
and U8243 (N_8243,N_8119,N_8110);
xnor U8244 (N_8244,N_8148,N_8086);
xnor U8245 (N_8245,N_8090,N_8177);
nor U8246 (N_8246,N_8095,N_8132);
nor U8247 (N_8247,N_8013,N_8098);
xnor U8248 (N_8248,N_8023,N_8121);
nand U8249 (N_8249,N_8141,N_8057);
nor U8250 (N_8250,N_8042,N_8113);
or U8251 (N_8251,N_8051,N_8131);
or U8252 (N_8252,N_8018,N_8037);
or U8253 (N_8253,N_8014,N_8127);
nand U8254 (N_8254,N_8197,N_8047);
xnor U8255 (N_8255,N_8053,N_8109);
nor U8256 (N_8256,N_8162,N_8120);
or U8257 (N_8257,N_8027,N_8152);
nor U8258 (N_8258,N_8024,N_8050);
nand U8259 (N_8259,N_8194,N_8134);
and U8260 (N_8260,N_8019,N_8151);
and U8261 (N_8261,N_8094,N_8083);
nand U8262 (N_8262,N_8022,N_8039);
nor U8263 (N_8263,N_8049,N_8017);
nand U8264 (N_8264,N_8066,N_8178);
or U8265 (N_8265,N_8180,N_8115);
and U8266 (N_8266,N_8048,N_8153);
nor U8267 (N_8267,N_8012,N_8021);
xor U8268 (N_8268,N_8114,N_8159);
and U8269 (N_8269,N_8029,N_8000);
or U8270 (N_8270,N_8158,N_8157);
nand U8271 (N_8271,N_8101,N_8055);
and U8272 (N_8272,N_8015,N_8058);
xnor U8273 (N_8273,N_8192,N_8181);
nand U8274 (N_8274,N_8033,N_8133);
nand U8275 (N_8275,N_8063,N_8040);
nor U8276 (N_8276,N_8056,N_8129);
or U8277 (N_8277,N_8155,N_8122);
nor U8278 (N_8278,N_8150,N_8104);
and U8279 (N_8279,N_8176,N_8074);
and U8280 (N_8280,N_8117,N_8186);
and U8281 (N_8281,N_8064,N_8112);
nor U8282 (N_8282,N_8198,N_8032);
xnor U8283 (N_8283,N_8060,N_8077);
or U8284 (N_8284,N_8161,N_8193);
xor U8285 (N_8285,N_8096,N_8010);
nand U8286 (N_8286,N_8111,N_8084);
xor U8287 (N_8287,N_8124,N_8179);
and U8288 (N_8288,N_8145,N_8036);
xnor U8289 (N_8289,N_8185,N_8171);
and U8290 (N_8290,N_8087,N_8188);
nand U8291 (N_8291,N_8140,N_8002);
nor U8292 (N_8292,N_8126,N_8130);
and U8293 (N_8293,N_8035,N_8085);
xor U8294 (N_8294,N_8107,N_8191);
nand U8295 (N_8295,N_8147,N_8068);
and U8296 (N_8296,N_8088,N_8025);
nand U8297 (N_8297,N_8190,N_8065);
nor U8298 (N_8298,N_8072,N_8034);
and U8299 (N_8299,N_8144,N_8045);
xnor U8300 (N_8300,N_8071,N_8022);
and U8301 (N_8301,N_8041,N_8094);
xnor U8302 (N_8302,N_8017,N_8133);
nand U8303 (N_8303,N_8115,N_8082);
or U8304 (N_8304,N_8034,N_8170);
xor U8305 (N_8305,N_8138,N_8012);
nand U8306 (N_8306,N_8148,N_8175);
nor U8307 (N_8307,N_8105,N_8178);
nand U8308 (N_8308,N_8161,N_8164);
or U8309 (N_8309,N_8158,N_8043);
or U8310 (N_8310,N_8084,N_8010);
or U8311 (N_8311,N_8107,N_8142);
and U8312 (N_8312,N_8019,N_8108);
or U8313 (N_8313,N_8045,N_8012);
xor U8314 (N_8314,N_8091,N_8108);
or U8315 (N_8315,N_8110,N_8184);
xor U8316 (N_8316,N_8136,N_8103);
nand U8317 (N_8317,N_8103,N_8162);
nor U8318 (N_8318,N_8197,N_8185);
nand U8319 (N_8319,N_8193,N_8067);
and U8320 (N_8320,N_8008,N_8060);
nor U8321 (N_8321,N_8162,N_8000);
nand U8322 (N_8322,N_8198,N_8109);
xnor U8323 (N_8323,N_8045,N_8171);
nand U8324 (N_8324,N_8068,N_8102);
or U8325 (N_8325,N_8045,N_8080);
nor U8326 (N_8326,N_8128,N_8168);
xnor U8327 (N_8327,N_8186,N_8016);
or U8328 (N_8328,N_8075,N_8188);
and U8329 (N_8329,N_8076,N_8056);
nand U8330 (N_8330,N_8154,N_8148);
or U8331 (N_8331,N_8108,N_8021);
or U8332 (N_8332,N_8184,N_8142);
or U8333 (N_8333,N_8044,N_8118);
nor U8334 (N_8334,N_8008,N_8080);
nor U8335 (N_8335,N_8015,N_8108);
xnor U8336 (N_8336,N_8119,N_8023);
and U8337 (N_8337,N_8004,N_8094);
nor U8338 (N_8338,N_8100,N_8009);
or U8339 (N_8339,N_8115,N_8001);
nand U8340 (N_8340,N_8195,N_8138);
nor U8341 (N_8341,N_8119,N_8111);
nor U8342 (N_8342,N_8152,N_8171);
nor U8343 (N_8343,N_8170,N_8008);
nor U8344 (N_8344,N_8002,N_8169);
or U8345 (N_8345,N_8179,N_8035);
and U8346 (N_8346,N_8092,N_8046);
or U8347 (N_8347,N_8185,N_8195);
or U8348 (N_8348,N_8124,N_8189);
and U8349 (N_8349,N_8057,N_8126);
nor U8350 (N_8350,N_8103,N_8016);
xnor U8351 (N_8351,N_8168,N_8186);
xor U8352 (N_8352,N_8088,N_8050);
nand U8353 (N_8353,N_8179,N_8036);
and U8354 (N_8354,N_8096,N_8142);
or U8355 (N_8355,N_8000,N_8195);
and U8356 (N_8356,N_8080,N_8114);
or U8357 (N_8357,N_8155,N_8145);
xnor U8358 (N_8358,N_8155,N_8042);
nand U8359 (N_8359,N_8183,N_8018);
nand U8360 (N_8360,N_8158,N_8194);
or U8361 (N_8361,N_8171,N_8019);
nand U8362 (N_8362,N_8137,N_8061);
and U8363 (N_8363,N_8041,N_8071);
and U8364 (N_8364,N_8109,N_8189);
or U8365 (N_8365,N_8167,N_8093);
nor U8366 (N_8366,N_8184,N_8099);
nor U8367 (N_8367,N_8015,N_8173);
xor U8368 (N_8368,N_8029,N_8070);
xor U8369 (N_8369,N_8126,N_8133);
xor U8370 (N_8370,N_8129,N_8143);
or U8371 (N_8371,N_8158,N_8103);
and U8372 (N_8372,N_8167,N_8000);
and U8373 (N_8373,N_8036,N_8008);
nor U8374 (N_8374,N_8074,N_8153);
or U8375 (N_8375,N_8144,N_8016);
xnor U8376 (N_8376,N_8073,N_8166);
nor U8377 (N_8377,N_8074,N_8037);
xor U8378 (N_8378,N_8006,N_8057);
nand U8379 (N_8379,N_8146,N_8157);
xor U8380 (N_8380,N_8119,N_8002);
and U8381 (N_8381,N_8105,N_8191);
xnor U8382 (N_8382,N_8195,N_8144);
xor U8383 (N_8383,N_8177,N_8169);
nor U8384 (N_8384,N_8033,N_8120);
nand U8385 (N_8385,N_8055,N_8186);
and U8386 (N_8386,N_8188,N_8070);
xnor U8387 (N_8387,N_8000,N_8061);
or U8388 (N_8388,N_8144,N_8043);
xor U8389 (N_8389,N_8078,N_8024);
nor U8390 (N_8390,N_8071,N_8025);
nand U8391 (N_8391,N_8150,N_8051);
or U8392 (N_8392,N_8094,N_8067);
and U8393 (N_8393,N_8187,N_8160);
xnor U8394 (N_8394,N_8197,N_8183);
nor U8395 (N_8395,N_8054,N_8030);
or U8396 (N_8396,N_8195,N_8052);
and U8397 (N_8397,N_8127,N_8180);
nor U8398 (N_8398,N_8096,N_8150);
nand U8399 (N_8399,N_8042,N_8059);
and U8400 (N_8400,N_8283,N_8324);
nor U8401 (N_8401,N_8348,N_8209);
nand U8402 (N_8402,N_8204,N_8264);
or U8403 (N_8403,N_8303,N_8278);
nor U8404 (N_8404,N_8260,N_8369);
xnor U8405 (N_8405,N_8228,N_8289);
nor U8406 (N_8406,N_8393,N_8365);
nor U8407 (N_8407,N_8230,N_8325);
nor U8408 (N_8408,N_8331,N_8231);
or U8409 (N_8409,N_8248,N_8249);
nor U8410 (N_8410,N_8363,N_8342);
and U8411 (N_8411,N_8329,N_8326);
or U8412 (N_8412,N_8272,N_8284);
and U8413 (N_8413,N_8336,N_8310);
and U8414 (N_8414,N_8337,N_8247);
or U8415 (N_8415,N_8382,N_8270);
nor U8416 (N_8416,N_8371,N_8244);
or U8417 (N_8417,N_8350,N_8259);
xnor U8418 (N_8418,N_8216,N_8268);
or U8419 (N_8419,N_8296,N_8275);
nand U8420 (N_8420,N_8306,N_8226);
xor U8421 (N_8421,N_8234,N_8392);
xnor U8422 (N_8422,N_8314,N_8295);
or U8423 (N_8423,N_8355,N_8367);
or U8424 (N_8424,N_8321,N_8307);
nor U8425 (N_8425,N_8288,N_8286);
or U8426 (N_8426,N_8316,N_8273);
xnor U8427 (N_8427,N_8354,N_8225);
and U8428 (N_8428,N_8334,N_8368);
nand U8429 (N_8429,N_8219,N_8323);
and U8430 (N_8430,N_8387,N_8269);
nand U8431 (N_8431,N_8294,N_8338);
xnor U8432 (N_8432,N_8292,N_8300);
or U8433 (N_8433,N_8255,N_8237);
xor U8434 (N_8434,N_8360,N_8281);
nor U8435 (N_8435,N_8266,N_8271);
nand U8436 (N_8436,N_8333,N_8358);
xnor U8437 (N_8437,N_8344,N_8224);
nand U8438 (N_8438,N_8319,N_8227);
nand U8439 (N_8439,N_8267,N_8347);
and U8440 (N_8440,N_8313,N_8362);
nand U8441 (N_8441,N_8318,N_8254);
or U8442 (N_8442,N_8312,N_8299);
nor U8443 (N_8443,N_8357,N_8343);
xnor U8444 (N_8444,N_8257,N_8341);
and U8445 (N_8445,N_8220,N_8239);
nor U8446 (N_8446,N_8398,N_8250);
nand U8447 (N_8447,N_8315,N_8389);
xor U8448 (N_8448,N_8383,N_8339);
and U8449 (N_8449,N_8243,N_8395);
or U8450 (N_8450,N_8322,N_8332);
nor U8451 (N_8451,N_8208,N_8301);
nor U8452 (N_8452,N_8205,N_8399);
xor U8453 (N_8453,N_8297,N_8223);
nor U8454 (N_8454,N_8349,N_8370);
nor U8455 (N_8455,N_8202,N_8235);
nand U8456 (N_8456,N_8374,N_8236);
or U8457 (N_8457,N_8253,N_8251);
nor U8458 (N_8458,N_8364,N_8311);
nor U8459 (N_8459,N_8330,N_8340);
xnor U8460 (N_8460,N_8372,N_8380);
nor U8461 (N_8461,N_8376,N_8391);
nor U8462 (N_8462,N_8386,N_8308);
nor U8463 (N_8463,N_8375,N_8366);
xor U8464 (N_8464,N_8305,N_8252);
nand U8465 (N_8465,N_8302,N_8335);
nor U8466 (N_8466,N_8261,N_8352);
xnor U8467 (N_8467,N_8203,N_8214);
nand U8468 (N_8468,N_8373,N_8291);
nand U8469 (N_8469,N_8298,N_8274);
or U8470 (N_8470,N_8359,N_8206);
or U8471 (N_8471,N_8293,N_8245);
or U8472 (N_8472,N_8282,N_8221);
and U8473 (N_8473,N_8233,N_8232);
nor U8474 (N_8474,N_8240,N_8384);
and U8475 (N_8475,N_8345,N_8263);
nor U8476 (N_8476,N_8356,N_8279);
nand U8477 (N_8477,N_8378,N_8396);
xor U8478 (N_8478,N_8262,N_8328);
nand U8479 (N_8479,N_8377,N_8394);
nand U8480 (N_8480,N_8242,N_8212);
or U8481 (N_8481,N_8229,N_8290);
xnor U8482 (N_8482,N_8276,N_8277);
or U8483 (N_8483,N_8210,N_8346);
and U8484 (N_8484,N_8379,N_8351);
xnor U8485 (N_8485,N_8213,N_8361);
nor U8486 (N_8486,N_8246,N_8238);
xor U8487 (N_8487,N_8390,N_8222);
nand U8488 (N_8488,N_8217,N_8353);
and U8489 (N_8489,N_8280,N_8317);
and U8490 (N_8490,N_8265,N_8397);
xor U8491 (N_8491,N_8309,N_8200);
and U8492 (N_8492,N_8304,N_8258);
nor U8493 (N_8493,N_8327,N_8287);
and U8494 (N_8494,N_8241,N_8256);
or U8495 (N_8495,N_8218,N_8388);
nor U8496 (N_8496,N_8385,N_8207);
and U8497 (N_8497,N_8381,N_8215);
nor U8498 (N_8498,N_8320,N_8201);
and U8499 (N_8499,N_8211,N_8285);
or U8500 (N_8500,N_8312,N_8261);
nand U8501 (N_8501,N_8305,N_8227);
and U8502 (N_8502,N_8361,N_8360);
xor U8503 (N_8503,N_8365,N_8217);
or U8504 (N_8504,N_8378,N_8270);
nor U8505 (N_8505,N_8351,N_8255);
nor U8506 (N_8506,N_8383,N_8350);
or U8507 (N_8507,N_8336,N_8284);
and U8508 (N_8508,N_8343,N_8294);
or U8509 (N_8509,N_8346,N_8364);
nand U8510 (N_8510,N_8220,N_8238);
or U8511 (N_8511,N_8294,N_8293);
nand U8512 (N_8512,N_8315,N_8353);
nor U8513 (N_8513,N_8355,N_8398);
xor U8514 (N_8514,N_8355,N_8378);
and U8515 (N_8515,N_8206,N_8209);
or U8516 (N_8516,N_8324,N_8379);
nor U8517 (N_8517,N_8249,N_8263);
and U8518 (N_8518,N_8202,N_8390);
or U8519 (N_8519,N_8290,N_8287);
xnor U8520 (N_8520,N_8301,N_8225);
or U8521 (N_8521,N_8263,N_8353);
xor U8522 (N_8522,N_8288,N_8251);
nor U8523 (N_8523,N_8320,N_8363);
and U8524 (N_8524,N_8205,N_8359);
nor U8525 (N_8525,N_8297,N_8394);
or U8526 (N_8526,N_8291,N_8390);
nor U8527 (N_8527,N_8351,N_8292);
nand U8528 (N_8528,N_8323,N_8220);
xnor U8529 (N_8529,N_8338,N_8314);
nor U8530 (N_8530,N_8250,N_8263);
nor U8531 (N_8531,N_8208,N_8285);
xnor U8532 (N_8532,N_8302,N_8290);
nor U8533 (N_8533,N_8236,N_8212);
or U8534 (N_8534,N_8264,N_8218);
xor U8535 (N_8535,N_8267,N_8346);
and U8536 (N_8536,N_8262,N_8258);
or U8537 (N_8537,N_8370,N_8392);
nor U8538 (N_8538,N_8343,N_8272);
nand U8539 (N_8539,N_8368,N_8350);
nand U8540 (N_8540,N_8263,N_8339);
xnor U8541 (N_8541,N_8319,N_8299);
nand U8542 (N_8542,N_8219,N_8378);
nor U8543 (N_8543,N_8206,N_8275);
or U8544 (N_8544,N_8244,N_8382);
nor U8545 (N_8545,N_8373,N_8267);
nor U8546 (N_8546,N_8283,N_8219);
nor U8547 (N_8547,N_8220,N_8353);
nor U8548 (N_8548,N_8307,N_8379);
nor U8549 (N_8549,N_8250,N_8260);
or U8550 (N_8550,N_8227,N_8274);
or U8551 (N_8551,N_8326,N_8331);
xnor U8552 (N_8552,N_8397,N_8206);
or U8553 (N_8553,N_8379,N_8212);
xor U8554 (N_8554,N_8373,N_8215);
or U8555 (N_8555,N_8334,N_8338);
and U8556 (N_8556,N_8388,N_8204);
and U8557 (N_8557,N_8228,N_8281);
or U8558 (N_8558,N_8307,N_8345);
and U8559 (N_8559,N_8364,N_8201);
nand U8560 (N_8560,N_8358,N_8305);
nor U8561 (N_8561,N_8247,N_8317);
or U8562 (N_8562,N_8366,N_8221);
xnor U8563 (N_8563,N_8276,N_8256);
and U8564 (N_8564,N_8246,N_8296);
or U8565 (N_8565,N_8356,N_8238);
xnor U8566 (N_8566,N_8293,N_8393);
and U8567 (N_8567,N_8306,N_8327);
xor U8568 (N_8568,N_8387,N_8362);
xor U8569 (N_8569,N_8306,N_8307);
or U8570 (N_8570,N_8355,N_8292);
nand U8571 (N_8571,N_8369,N_8254);
nor U8572 (N_8572,N_8297,N_8373);
xnor U8573 (N_8573,N_8365,N_8264);
nor U8574 (N_8574,N_8201,N_8372);
nor U8575 (N_8575,N_8276,N_8366);
and U8576 (N_8576,N_8223,N_8211);
or U8577 (N_8577,N_8223,N_8391);
or U8578 (N_8578,N_8279,N_8340);
xor U8579 (N_8579,N_8348,N_8390);
and U8580 (N_8580,N_8330,N_8335);
and U8581 (N_8581,N_8321,N_8210);
and U8582 (N_8582,N_8338,N_8216);
or U8583 (N_8583,N_8372,N_8202);
or U8584 (N_8584,N_8247,N_8258);
nand U8585 (N_8585,N_8233,N_8220);
xnor U8586 (N_8586,N_8369,N_8281);
or U8587 (N_8587,N_8212,N_8347);
and U8588 (N_8588,N_8254,N_8335);
or U8589 (N_8589,N_8263,N_8229);
or U8590 (N_8590,N_8232,N_8290);
xor U8591 (N_8591,N_8393,N_8203);
and U8592 (N_8592,N_8305,N_8370);
nand U8593 (N_8593,N_8244,N_8322);
and U8594 (N_8594,N_8355,N_8239);
and U8595 (N_8595,N_8276,N_8310);
and U8596 (N_8596,N_8273,N_8377);
xor U8597 (N_8597,N_8323,N_8239);
nor U8598 (N_8598,N_8326,N_8261);
or U8599 (N_8599,N_8391,N_8295);
or U8600 (N_8600,N_8470,N_8561);
nand U8601 (N_8601,N_8413,N_8580);
nor U8602 (N_8602,N_8548,N_8474);
nor U8603 (N_8603,N_8593,N_8585);
nand U8604 (N_8604,N_8501,N_8571);
nor U8605 (N_8605,N_8459,N_8473);
or U8606 (N_8606,N_8505,N_8402);
xor U8607 (N_8607,N_8407,N_8523);
and U8608 (N_8608,N_8436,N_8556);
xor U8609 (N_8609,N_8451,N_8450);
nand U8610 (N_8610,N_8558,N_8551);
or U8611 (N_8611,N_8524,N_8546);
xnor U8612 (N_8612,N_8599,N_8590);
and U8613 (N_8613,N_8491,N_8447);
and U8614 (N_8614,N_8477,N_8460);
nor U8615 (N_8615,N_8539,N_8515);
or U8616 (N_8616,N_8445,N_8589);
xnor U8617 (N_8617,N_8552,N_8489);
or U8618 (N_8618,N_8442,N_8403);
nor U8619 (N_8619,N_8577,N_8471);
xnor U8620 (N_8620,N_8569,N_8430);
xnor U8621 (N_8621,N_8400,N_8525);
nand U8622 (N_8622,N_8418,N_8527);
and U8623 (N_8623,N_8410,N_8508);
or U8624 (N_8624,N_8519,N_8444);
and U8625 (N_8625,N_8521,N_8578);
or U8626 (N_8626,N_8531,N_8591);
xor U8627 (N_8627,N_8476,N_8554);
and U8628 (N_8628,N_8453,N_8574);
nor U8629 (N_8629,N_8428,N_8411);
or U8630 (N_8630,N_8421,N_8446);
and U8631 (N_8631,N_8542,N_8466);
nand U8632 (N_8632,N_8439,N_8573);
xnor U8633 (N_8633,N_8497,N_8429);
and U8634 (N_8634,N_8467,N_8452);
and U8635 (N_8635,N_8465,N_8435);
xor U8636 (N_8636,N_8425,N_8547);
or U8637 (N_8637,N_8541,N_8555);
and U8638 (N_8638,N_8427,N_8405);
nor U8639 (N_8639,N_8462,N_8495);
xnor U8640 (N_8640,N_8420,N_8543);
and U8641 (N_8641,N_8401,N_8406);
and U8642 (N_8642,N_8480,N_8522);
xor U8643 (N_8643,N_8537,N_8582);
xnor U8644 (N_8644,N_8478,N_8506);
nor U8645 (N_8645,N_8534,N_8550);
and U8646 (N_8646,N_8414,N_8559);
or U8647 (N_8647,N_8468,N_8529);
nand U8648 (N_8648,N_8493,N_8502);
and U8649 (N_8649,N_8499,N_8448);
nor U8650 (N_8650,N_8565,N_8482);
xnor U8651 (N_8651,N_8503,N_8562);
nand U8652 (N_8652,N_8526,N_8423);
and U8653 (N_8653,N_8498,N_8588);
nand U8654 (N_8654,N_8458,N_8504);
or U8655 (N_8655,N_8449,N_8431);
or U8656 (N_8656,N_8422,N_8463);
xnor U8657 (N_8657,N_8479,N_8583);
nor U8658 (N_8658,N_8592,N_8419);
nand U8659 (N_8659,N_8579,N_8520);
and U8660 (N_8660,N_8461,N_8514);
or U8661 (N_8661,N_8440,N_8426);
xor U8662 (N_8662,N_8409,N_8469);
or U8663 (N_8663,N_8416,N_8483);
and U8664 (N_8664,N_8511,N_8454);
nor U8665 (N_8665,N_8566,N_8472);
xor U8666 (N_8666,N_8568,N_8596);
and U8667 (N_8667,N_8581,N_8538);
nand U8668 (N_8668,N_8432,N_8560);
and U8669 (N_8669,N_8507,N_8433);
xor U8670 (N_8670,N_8443,N_8570);
and U8671 (N_8671,N_8487,N_8530);
nand U8672 (N_8672,N_8494,N_8490);
or U8673 (N_8673,N_8481,N_8563);
nand U8674 (N_8674,N_8564,N_8510);
nand U8675 (N_8675,N_8528,N_8485);
nor U8676 (N_8676,N_8572,N_8533);
xor U8677 (N_8677,N_8500,N_8540);
nand U8678 (N_8678,N_8575,N_8532);
nand U8679 (N_8679,N_8584,N_8404);
nand U8680 (N_8680,N_8488,N_8492);
nand U8681 (N_8681,N_8536,N_8516);
or U8682 (N_8682,N_8509,N_8412);
nor U8683 (N_8683,N_8496,N_8484);
and U8684 (N_8684,N_8512,N_8424);
nand U8685 (N_8685,N_8535,N_8417);
or U8686 (N_8686,N_8456,N_8594);
or U8687 (N_8687,N_8557,N_8595);
or U8688 (N_8688,N_8518,N_8437);
xor U8689 (N_8689,N_8553,N_8455);
xor U8690 (N_8690,N_8597,N_8517);
nor U8691 (N_8691,N_8587,N_8576);
nor U8692 (N_8692,N_8457,N_8544);
or U8693 (N_8693,N_8586,N_8438);
and U8694 (N_8694,N_8567,N_8486);
nand U8695 (N_8695,N_8441,N_8513);
or U8696 (N_8696,N_8598,N_8545);
nand U8697 (N_8697,N_8549,N_8475);
and U8698 (N_8698,N_8464,N_8415);
nand U8699 (N_8699,N_8408,N_8434);
and U8700 (N_8700,N_8593,N_8599);
nor U8701 (N_8701,N_8491,N_8514);
or U8702 (N_8702,N_8561,N_8578);
nand U8703 (N_8703,N_8406,N_8502);
nor U8704 (N_8704,N_8497,N_8486);
or U8705 (N_8705,N_8460,N_8591);
or U8706 (N_8706,N_8587,N_8489);
nand U8707 (N_8707,N_8562,N_8446);
nand U8708 (N_8708,N_8585,N_8402);
or U8709 (N_8709,N_8455,N_8558);
or U8710 (N_8710,N_8593,N_8490);
or U8711 (N_8711,N_8471,N_8459);
and U8712 (N_8712,N_8592,N_8561);
nor U8713 (N_8713,N_8481,N_8449);
and U8714 (N_8714,N_8472,N_8512);
or U8715 (N_8715,N_8491,N_8515);
nor U8716 (N_8716,N_8550,N_8451);
xor U8717 (N_8717,N_8503,N_8595);
and U8718 (N_8718,N_8547,N_8583);
or U8719 (N_8719,N_8456,N_8583);
or U8720 (N_8720,N_8563,N_8453);
nand U8721 (N_8721,N_8481,N_8450);
xor U8722 (N_8722,N_8506,N_8438);
nand U8723 (N_8723,N_8557,N_8435);
and U8724 (N_8724,N_8435,N_8509);
nand U8725 (N_8725,N_8414,N_8542);
and U8726 (N_8726,N_8476,N_8435);
or U8727 (N_8727,N_8519,N_8450);
nand U8728 (N_8728,N_8419,N_8543);
nand U8729 (N_8729,N_8417,N_8554);
or U8730 (N_8730,N_8421,N_8490);
nand U8731 (N_8731,N_8555,N_8431);
nor U8732 (N_8732,N_8539,N_8478);
nor U8733 (N_8733,N_8428,N_8592);
xor U8734 (N_8734,N_8401,N_8550);
nor U8735 (N_8735,N_8546,N_8402);
or U8736 (N_8736,N_8514,N_8481);
and U8737 (N_8737,N_8443,N_8486);
or U8738 (N_8738,N_8513,N_8564);
nor U8739 (N_8739,N_8468,N_8598);
or U8740 (N_8740,N_8527,N_8426);
nand U8741 (N_8741,N_8460,N_8488);
or U8742 (N_8742,N_8488,N_8509);
or U8743 (N_8743,N_8556,N_8592);
and U8744 (N_8744,N_8496,N_8508);
nor U8745 (N_8745,N_8599,N_8437);
xor U8746 (N_8746,N_8547,N_8538);
xor U8747 (N_8747,N_8499,N_8554);
nor U8748 (N_8748,N_8503,N_8566);
xor U8749 (N_8749,N_8478,N_8411);
xnor U8750 (N_8750,N_8437,N_8443);
nor U8751 (N_8751,N_8498,N_8473);
and U8752 (N_8752,N_8576,N_8519);
and U8753 (N_8753,N_8493,N_8461);
nor U8754 (N_8754,N_8404,N_8572);
nand U8755 (N_8755,N_8445,N_8558);
nand U8756 (N_8756,N_8562,N_8453);
nor U8757 (N_8757,N_8413,N_8508);
nand U8758 (N_8758,N_8461,N_8400);
xnor U8759 (N_8759,N_8416,N_8428);
nand U8760 (N_8760,N_8541,N_8488);
and U8761 (N_8761,N_8453,N_8591);
nor U8762 (N_8762,N_8417,N_8413);
nand U8763 (N_8763,N_8560,N_8584);
xnor U8764 (N_8764,N_8580,N_8520);
xor U8765 (N_8765,N_8548,N_8487);
or U8766 (N_8766,N_8521,N_8484);
nand U8767 (N_8767,N_8493,N_8576);
xor U8768 (N_8768,N_8439,N_8522);
and U8769 (N_8769,N_8413,N_8541);
and U8770 (N_8770,N_8504,N_8420);
nor U8771 (N_8771,N_8447,N_8477);
nand U8772 (N_8772,N_8495,N_8572);
nand U8773 (N_8773,N_8404,N_8551);
nand U8774 (N_8774,N_8436,N_8524);
nand U8775 (N_8775,N_8452,N_8495);
or U8776 (N_8776,N_8549,N_8472);
and U8777 (N_8777,N_8559,N_8527);
nand U8778 (N_8778,N_8495,N_8571);
or U8779 (N_8779,N_8576,N_8584);
xor U8780 (N_8780,N_8469,N_8560);
and U8781 (N_8781,N_8490,N_8570);
and U8782 (N_8782,N_8587,N_8509);
nor U8783 (N_8783,N_8474,N_8545);
xnor U8784 (N_8784,N_8400,N_8402);
or U8785 (N_8785,N_8475,N_8476);
xnor U8786 (N_8786,N_8550,N_8442);
nand U8787 (N_8787,N_8495,N_8414);
xnor U8788 (N_8788,N_8596,N_8488);
xnor U8789 (N_8789,N_8506,N_8459);
or U8790 (N_8790,N_8513,N_8424);
and U8791 (N_8791,N_8535,N_8520);
or U8792 (N_8792,N_8514,N_8493);
or U8793 (N_8793,N_8413,N_8592);
and U8794 (N_8794,N_8524,N_8548);
or U8795 (N_8795,N_8409,N_8466);
or U8796 (N_8796,N_8542,N_8526);
nand U8797 (N_8797,N_8530,N_8460);
and U8798 (N_8798,N_8507,N_8547);
and U8799 (N_8799,N_8521,N_8512);
or U8800 (N_8800,N_8601,N_8725);
and U8801 (N_8801,N_8747,N_8688);
nor U8802 (N_8802,N_8605,N_8743);
xnor U8803 (N_8803,N_8760,N_8726);
nor U8804 (N_8804,N_8685,N_8625);
nor U8805 (N_8805,N_8604,N_8739);
nor U8806 (N_8806,N_8679,N_8674);
nor U8807 (N_8807,N_8617,N_8650);
or U8808 (N_8808,N_8771,N_8736);
nor U8809 (N_8809,N_8700,N_8733);
and U8810 (N_8810,N_8602,N_8680);
nor U8811 (N_8811,N_8764,N_8699);
nor U8812 (N_8812,N_8657,N_8632);
nand U8813 (N_8813,N_8669,N_8702);
and U8814 (N_8814,N_8682,N_8732);
and U8815 (N_8815,N_8729,N_8609);
and U8816 (N_8816,N_8754,N_8647);
nor U8817 (N_8817,N_8709,N_8681);
and U8818 (N_8818,N_8783,N_8759);
or U8819 (N_8819,N_8621,N_8654);
nor U8820 (N_8820,N_8646,N_8798);
or U8821 (N_8821,N_8797,N_8660);
or U8822 (N_8822,N_8761,N_8766);
xnor U8823 (N_8823,N_8636,N_8786);
and U8824 (N_8824,N_8706,N_8640);
and U8825 (N_8825,N_8762,N_8751);
and U8826 (N_8826,N_8789,N_8607);
nor U8827 (N_8827,N_8757,N_8667);
and U8828 (N_8828,N_8637,N_8626);
nor U8829 (N_8829,N_8794,N_8755);
nor U8830 (N_8830,N_8696,N_8675);
or U8831 (N_8831,N_8666,N_8690);
nand U8832 (N_8832,N_8683,N_8780);
or U8833 (N_8833,N_8738,N_8792);
or U8834 (N_8834,N_8641,N_8689);
nor U8835 (N_8835,N_8718,N_8684);
nor U8836 (N_8836,N_8623,N_8624);
and U8837 (N_8837,N_8779,N_8676);
nor U8838 (N_8838,N_8663,N_8677);
xnor U8839 (N_8839,N_8756,N_8645);
and U8840 (N_8840,N_8701,N_8713);
nor U8841 (N_8841,N_8704,N_8723);
nor U8842 (N_8842,N_8662,N_8740);
nand U8843 (N_8843,N_8672,N_8731);
nand U8844 (N_8844,N_8639,N_8613);
nor U8845 (N_8845,N_8727,N_8734);
and U8846 (N_8846,N_8653,N_8774);
or U8847 (N_8847,N_8777,N_8742);
xor U8848 (N_8848,N_8776,N_8611);
nand U8849 (N_8849,N_8711,N_8785);
and U8850 (N_8850,N_8622,N_8749);
nand U8851 (N_8851,N_8610,N_8630);
nand U8852 (N_8852,N_8796,N_8670);
and U8853 (N_8853,N_8627,N_8678);
nand U8854 (N_8854,N_8620,N_8715);
nor U8855 (N_8855,N_8703,N_8750);
or U8856 (N_8856,N_8722,N_8656);
xor U8857 (N_8857,N_8698,N_8716);
nor U8858 (N_8858,N_8687,N_8746);
nand U8859 (N_8859,N_8788,N_8724);
and U8860 (N_8860,N_8719,N_8695);
or U8861 (N_8861,N_8708,N_8752);
or U8862 (N_8862,N_8795,N_8651);
or U8863 (N_8863,N_8652,N_8763);
or U8864 (N_8864,N_8720,N_8772);
nor U8865 (N_8865,N_8694,N_8730);
and U8866 (N_8866,N_8707,N_8745);
nor U8867 (N_8867,N_8608,N_8778);
and U8868 (N_8868,N_8633,N_8673);
and U8869 (N_8869,N_8668,N_8628);
and U8870 (N_8870,N_8648,N_8642);
nand U8871 (N_8871,N_8692,N_8721);
and U8872 (N_8872,N_8758,N_8741);
nor U8873 (N_8873,N_8655,N_8659);
or U8874 (N_8874,N_8649,N_8635);
or U8875 (N_8875,N_8665,N_8769);
and U8876 (N_8876,N_8705,N_8781);
xor U8877 (N_8877,N_8691,N_8799);
xnor U8878 (N_8878,N_8784,N_8710);
xor U8879 (N_8879,N_8631,N_8671);
and U8880 (N_8880,N_8634,N_8737);
or U8881 (N_8881,N_8728,N_8638);
nor U8882 (N_8882,N_8748,N_8790);
or U8883 (N_8883,N_8717,N_8664);
xor U8884 (N_8884,N_8782,N_8643);
and U8885 (N_8885,N_8658,N_8787);
nand U8886 (N_8886,N_8661,N_8603);
nand U8887 (N_8887,N_8712,N_8791);
nor U8888 (N_8888,N_8618,N_8770);
nand U8889 (N_8889,N_8768,N_8619);
or U8890 (N_8890,N_8765,N_8629);
nor U8891 (N_8891,N_8753,N_8735);
nor U8892 (N_8892,N_8600,N_8612);
xnor U8893 (N_8893,N_8714,N_8686);
xnor U8894 (N_8894,N_8697,N_8744);
or U8895 (N_8895,N_8793,N_8615);
or U8896 (N_8896,N_8693,N_8775);
and U8897 (N_8897,N_8644,N_8606);
and U8898 (N_8898,N_8614,N_8773);
nor U8899 (N_8899,N_8767,N_8616);
nand U8900 (N_8900,N_8692,N_8656);
nor U8901 (N_8901,N_8783,N_8646);
and U8902 (N_8902,N_8714,N_8671);
nand U8903 (N_8903,N_8620,N_8790);
or U8904 (N_8904,N_8604,N_8772);
nand U8905 (N_8905,N_8618,N_8708);
xnor U8906 (N_8906,N_8619,N_8766);
or U8907 (N_8907,N_8670,N_8625);
or U8908 (N_8908,N_8698,N_8611);
nor U8909 (N_8909,N_8677,N_8761);
nor U8910 (N_8910,N_8609,N_8762);
xor U8911 (N_8911,N_8763,N_8762);
nand U8912 (N_8912,N_8693,N_8638);
nor U8913 (N_8913,N_8638,N_8794);
nand U8914 (N_8914,N_8780,N_8755);
xor U8915 (N_8915,N_8767,N_8608);
nor U8916 (N_8916,N_8738,N_8631);
xnor U8917 (N_8917,N_8731,N_8698);
nand U8918 (N_8918,N_8683,N_8773);
nor U8919 (N_8919,N_8613,N_8607);
xnor U8920 (N_8920,N_8799,N_8701);
nor U8921 (N_8921,N_8674,N_8629);
and U8922 (N_8922,N_8745,N_8722);
xnor U8923 (N_8923,N_8786,N_8760);
xnor U8924 (N_8924,N_8602,N_8648);
nor U8925 (N_8925,N_8781,N_8729);
and U8926 (N_8926,N_8602,N_8699);
and U8927 (N_8927,N_8757,N_8608);
and U8928 (N_8928,N_8706,N_8695);
nor U8929 (N_8929,N_8774,N_8798);
and U8930 (N_8930,N_8741,N_8784);
nand U8931 (N_8931,N_8601,N_8655);
xor U8932 (N_8932,N_8618,N_8774);
or U8933 (N_8933,N_8667,N_8660);
xor U8934 (N_8934,N_8633,N_8656);
nand U8935 (N_8935,N_8756,N_8731);
nor U8936 (N_8936,N_8702,N_8760);
nor U8937 (N_8937,N_8718,N_8792);
nand U8938 (N_8938,N_8770,N_8732);
nand U8939 (N_8939,N_8727,N_8625);
xor U8940 (N_8940,N_8727,N_8611);
or U8941 (N_8941,N_8689,N_8797);
and U8942 (N_8942,N_8746,N_8605);
xor U8943 (N_8943,N_8678,N_8743);
and U8944 (N_8944,N_8711,N_8634);
xnor U8945 (N_8945,N_8798,N_8737);
nand U8946 (N_8946,N_8799,N_8696);
nor U8947 (N_8947,N_8719,N_8794);
or U8948 (N_8948,N_8716,N_8693);
nand U8949 (N_8949,N_8786,N_8691);
nor U8950 (N_8950,N_8795,N_8624);
or U8951 (N_8951,N_8629,N_8789);
xnor U8952 (N_8952,N_8747,N_8717);
or U8953 (N_8953,N_8788,N_8624);
nand U8954 (N_8954,N_8700,N_8780);
nand U8955 (N_8955,N_8762,N_8625);
and U8956 (N_8956,N_8749,N_8696);
nand U8957 (N_8957,N_8633,N_8751);
nor U8958 (N_8958,N_8618,N_8649);
xnor U8959 (N_8959,N_8613,N_8796);
nand U8960 (N_8960,N_8686,N_8780);
nor U8961 (N_8961,N_8607,N_8658);
nand U8962 (N_8962,N_8783,N_8788);
or U8963 (N_8963,N_8647,N_8785);
and U8964 (N_8964,N_8685,N_8656);
nor U8965 (N_8965,N_8716,N_8690);
or U8966 (N_8966,N_8649,N_8683);
or U8967 (N_8967,N_8696,N_8691);
xnor U8968 (N_8968,N_8760,N_8725);
nor U8969 (N_8969,N_8769,N_8637);
or U8970 (N_8970,N_8758,N_8622);
and U8971 (N_8971,N_8712,N_8719);
nand U8972 (N_8972,N_8756,N_8608);
or U8973 (N_8973,N_8647,N_8634);
xor U8974 (N_8974,N_8623,N_8753);
and U8975 (N_8975,N_8680,N_8721);
xor U8976 (N_8976,N_8659,N_8733);
nor U8977 (N_8977,N_8740,N_8739);
and U8978 (N_8978,N_8798,N_8640);
or U8979 (N_8979,N_8687,N_8604);
xnor U8980 (N_8980,N_8740,N_8710);
xnor U8981 (N_8981,N_8792,N_8610);
nand U8982 (N_8982,N_8686,N_8600);
xor U8983 (N_8983,N_8691,N_8774);
nor U8984 (N_8984,N_8755,N_8785);
or U8985 (N_8985,N_8755,N_8741);
nor U8986 (N_8986,N_8705,N_8730);
xor U8987 (N_8987,N_8786,N_8772);
nand U8988 (N_8988,N_8741,N_8795);
xnor U8989 (N_8989,N_8732,N_8606);
xnor U8990 (N_8990,N_8630,N_8703);
and U8991 (N_8991,N_8705,N_8696);
nand U8992 (N_8992,N_8690,N_8738);
nor U8993 (N_8993,N_8712,N_8623);
or U8994 (N_8994,N_8723,N_8765);
nor U8995 (N_8995,N_8628,N_8709);
nor U8996 (N_8996,N_8614,N_8690);
and U8997 (N_8997,N_8733,N_8677);
nand U8998 (N_8998,N_8694,N_8606);
and U8999 (N_8999,N_8793,N_8696);
nand U9000 (N_9000,N_8817,N_8915);
nand U9001 (N_9001,N_8898,N_8886);
nor U9002 (N_9002,N_8989,N_8919);
nor U9003 (N_9003,N_8809,N_8905);
nor U9004 (N_9004,N_8845,N_8856);
xnor U9005 (N_9005,N_8991,N_8884);
nand U9006 (N_9006,N_8834,N_8914);
and U9007 (N_9007,N_8978,N_8924);
nor U9008 (N_9008,N_8944,N_8862);
nand U9009 (N_9009,N_8950,N_8811);
nor U9010 (N_9010,N_8822,N_8827);
nand U9011 (N_9011,N_8910,N_8984);
nor U9012 (N_9012,N_8957,N_8952);
and U9013 (N_9013,N_8807,N_8879);
nand U9014 (N_9014,N_8873,N_8876);
nand U9015 (N_9015,N_8987,N_8964);
or U9016 (N_9016,N_8808,N_8930);
nand U9017 (N_9017,N_8891,N_8877);
nand U9018 (N_9018,N_8996,N_8913);
xnor U9019 (N_9019,N_8872,N_8859);
nand U9020 (N_9020,N_8979,N_8870);
or U9021 (N_9021,N_8896,N_8965);
and U9022 (N_9022,N_8970,N_8813);
nor U9023 (N_9023,N_8858,N_8982);
nand U9024 (N_9024,N_8893,N_8823);
nand U9025 (N_9025,N_8954,N_8941);
or U9026 (N_9026,N_8869,N_8820);
nand U9027 (N_9027,N_8985,N_8836);
nand U9028 (N_9028,N_8945,N_8997);
nand U9029 (N_9029,N_8933,N_8909);
and U9030 (N_9030,N_8904,N_8814);
xor U9031 (N_9031,N_8961,N_8816);
or U9032 (N_9032,N_8897,N_8971);
and U9033 (N_9033,N_8882,N_8846);
xnor U9034 (N_9034,N_8889,N_8926);
and U9035 (N_9035,N_8973,N_8912);
or U9036 (N_9036,N_8821,N_8843);
xor U9037 (N_9037,N_8967,N_8900);
or U9038 (N_9038,N_8990,N_8874);
nand U9039 (N_9039,N_8974,N_8931);
and U9040 (N_9040,N_8866,N_8951);
xor U9041 (N_9041,N_8850,N_8806);
or U9042 (N_9042,N_8819,N_8927);
or U9043 (N_9043,N_8980,N_8864);
nand U9044 (N_9044,N_8878,N_8800);
nand U9045 (N_9045,N_8981,N_8894);
and U9046 (N_9046,N_8976,N_8920);
and U9047 (N_9047,N_8956,N_8966);
xor U9048 (N_9048,N_8847,N_8865);
nand U9049 (N_9049,N_8977,N_8962);
nand U9050 (N_9050,N_8815,N_8922);
or U9051 (N_9051,N_8903,N_8867);
nor U9052 (N_9052,N_8881,N_8963);
or U9053 (N_9053,N_8887,N_8828);
xnor U9054 (N_9054,N_8959,N_8929);
xor U9055 (N_9055,N_8852,N_8936);
nor U9056 (N_9056,N_8804,N_8921);
nor U9057 (N_9057,N_8812,N_8824);
nor U9058 (N_9058,N_8983,N_8892);
xnor U9059 (N_9059,N_8937,N_8998);
or U9060 (N_9060,N_8829,N_8994);
nand U9061 (N_9061,N_8838,N_8841);
nand U9062 (N_9062,N_8940,N_8844);
and U9063 (N_9063,N_8953,N_8835);
xor U9064 (N_9064,N_8906,N_8972);
nor U9065 (N_9065,N_8995,N_8888);
and U9066 (N_9066,N_8830,N_8946);
xor U9067 (N_9067,N_8875,N_8938);
nand U9068 (N_9068,N_8999,N_8833);
xnor U9069 (N_9069,N_8960,N_8810);
nand U9070 (N_9070,N_8848,N_8993);
or U9071 (N_9071,N_8975,N_8902);
nor U9072 (N_9072,N_8942,N_8818);
nand U9073 (N_9073,N_8939,N_8840);
or U9074 (N_9074,N_8934,N_8803);
xnor U9075 (N_9075,N_8935,N_8907);
or U9076 (N_9076,N_8880,N_8857);
xnor U9077 (N_9077,N_8868,N_8986);
xor U9078 (N_9078,N_8854,N_8992);
xnor U9079 (N_9079,N_8916,N_8949);
and U9080 (N_9080,N_8918,N_8825);
nand U9081 (N_9081,N_8925,N_8958);
or U9082 (N_9082,N_8901,N_8890);
nand U9083 (N_9083,N_8928,N_8923);
nand U9084 (N_9084,N_8805,N_8801);
nand U9085 (N_9085,N_8899,N_8863);
xnor U9086 (N_9086,N_8871,N_8883);
or U9087 (N_9087,N_8853,N_8948);
nor U9088 (N_9088,N_8826,N_8885);
and U9089 (N_9089,N_8908,N_8932);
nand U9090 (N_9090,N_8832,N_8839);
nand U9091 (N_9091,N_8855,N_8988);
nor U9092 (N_9092,N_8917,N_8861);
xor U9093 (N_9093,N_8968,N_8969);
and U9094 (N_9094,N_8911,N_8860);
nor U9095 (N_9095,N_8831,N_8802);
or U9096 (N_9096,N_8895,N_8837);
xnor U9097 (N_9097,N_8943,N_8851);
nand U9098 (N_9098,N_8842,N_8849);
and U9099 (N_9099,N_8955,N_8947);
nor U9100 (N_9100,N_8939,N_8944);
or U9101 (N_9101,N_8933,N_8993);
xor U9102 (N_9102,N_8917,N_8977);
nand U9103 (N_9103,N_8946,N_8867);
nor U9104 (N_9104,N_8982,N_8979);
nand U9105 (N_9105,N_8851,N_8984);
or U9106 (N_9106,N_8968,N_8809);
or U9107 (N_9107,N_8838,N_8878);
xor U9108 (N_9108,N_8972,N_8869);
and U9109 (N_9109,N_8949,N_8967);
nand U9110 (N_9110,N_8965,N_8935);
xnor U9111 (N_9111,N_8950,N_8994);
xnor U9112 (N_9112,N_8960,N_8821);
or U9113 (N_9113,N_8879,N_8800);
nand U9114 (N_9114,N_8861,N_8865);
nand U9115 (N_9115,N_8947,N_8886);
and U9116 (N_9116,N_8950,N_8921);
and U9117 (N_9117,N_8901,N_8822);
or U9118 (N_9118,N_8898,N_8977);
nor U9119 (N_9119,N_8977,N_8875);
or U9120 (N_9120,N_8956,N_8816);
nor U9121 (N_9121,N_8890,N_8992);
nor U9122 (N_9122,N_8839,N_8908);
or U9123 (N_9123,N_8835,N_8957);
nand U9124 (N_9124,N_8947,N_8875);
xor U9125 (N_9125,N_8938,N_8867);
and U9126 (N_9126,N_8870,N_8845);
nand U9127 (N_9127,N_8997,N_8867);
or U9128 (N_9128,N_8868,N_8893);
nor U9129 (N_9129,N_8842,N_8950);
and U9130 (N_9130,N_8810,N_8824);
nand U9131 (N_9131,N_8937,N_8984);
xnor U9132 (N_9132,N_8915,N_8884);
nor U9133 (N_9133,N_8844,N_8808);
and U9134 (N_9134,N_8985,N_8898);
nand U9135 (N_9135,N_8941,N_8959);
or U9136 (N_9136,N_8891,N_8845);
and U9137 (N_9137,N_8829,N_8973);
or U9138 (N_9138,N_8844,N_8999);
xnor U9139 (N_9139,N_8996,N_8822);
and U9140 (N_9140,N_8950,N_8963);
and U9141 (N_9141,N_8967,N_8938);
and U9142 (N_9142,N_8884,N_8853);
nor U9143 (N_9143,N_8884,N_8995);
or U9144 (N_9144,N_8870,N_8802);
and U9145 (N_9145,N_8906,N_8953);
or U9146 (N_9146,N_8935,N_8855);
xor U9147 (N_9147,N_8968,N_8904);
and U9148 (N_9148,N_8839,N_8991);
and U9149 (N_9149,N_8928,N_8803);
xor U9150 (N_9150,N_8949,N_8806);
or U9151 (N_9151,N_8988,N_8968);
and U9152 (N_9152,N_8928,N_8830);
nand U9153 (N_9153,N_8874,N_8937);
nor U9154 (N_9154,N_8814,N_8890);
nor U9155 (N_9155,N_8834,N_8945);
and U9156 (N_9156,N_8812,N_8866);
xor U9157 (N_9157,N_8930,N_8847);
and U9158 (N_9158,N_8881,N_8998);
or U9159 (N_9159,N_8884,N_8997);
nor U9160 (N_9160,N_8989,N_8982);
nand U9161 (N_9161,N_8957,N_8991);
nor U9162 (N_9162,N_8970,N_8874);
or U9163 (N_9163,N_8827,N_8907);
or U9164 (N_9164,N_8911,N_8861);
or U9165 (N_9165,N_8937,N_8836);
xnor U9166 (N_9166,N_8938,N_8817);
or U9167 (N_9167,N_8955,N_8860);
and U9168 (N_9168,N_8981,N_8874);
and U9169 (N_9169,N_8928,N_8835);
xor U9170 (N_9170,N_8969,N_8888);
nand U9171 (N_9171,N_8940,N_8941);
and U9172 (N_9172,N_8924,N_8842);
xnor U9173 (N_9173,N_8885,N_8855);
nand U9174 (N_9174,N_8904,N_8859);
xnor U9175 (N_9175,N_8942,N_8859);
and U9176 (N_9176,N_8931,N_8927);
nor U9177 (N_9177,N_8986,N_8963);
nand U9178 (N_9178,N_8881,N_8970);
or U9179 (N_9179,N_8880,N_8897);
and U9180 (N_9180,N_8832,N_8945);
xnor U9181 (N_9181,N_8907,N_8865);
nor U9182 (N_9182,N_8841,N_8970);
nand U9183 (N_9183,N_8904,N_8906);
or U9184 (N_9184,N_8899,N_8834);
and U9185 (N_9185,N_8954,N_8832);
xor U9186 (N_9186,N_8956,N_8830);
nand U9187 (N_9187,N_8835,N_8884);
nor U9188 (N_9188,N_8852,N_8871);
or U9189 (N_9189,N_8810,N_8981);
xnor U9190 (N_9190,N_8871,N_8824);
or U9191 (N_9191,N_8807,N_8803);
and U9192 (N_9192,N_8860,N_8945);
xor U9193 (N_9193,N_8952,N_8882);
or U9194 (N_9194,N_8975,N_8961);
xnor U9195 (N_9195,N_8913,N_8869);
xnor U9196 (N_9196,N_8991,N_8962);
or U9197 (N_9197,N_8884,N_8822);
nand U9198 (N_9198,N_8838,N_8800);
nand U9199 (N_9199,N_8969,N_8938);
and U9200 (N_9200,N_9059,N_9101);
nor U9201 (N_9201,N_9079,N_9102);
and U9202 (N_9202,N_9106,N_9069);
or U9203 (N_9203,N_9000,N_9029);
and U9204 (N_9204,N_9030,N_9119);
or U9205 (N_9205,N_9189,N_9111);
and U9206 (N_9206,N_9093,N_9193);
xnor U9207 (N_9207,N_9147,N_9042);
or U9208 (N_9208,N_9050,N_9094);
nor U9209 (N_9209,N_9071,N_9139);
nand U9210 (N_9210,N_9121,N_9188);
or U9211 (N_9211,N_9027,N_9085);
xor U9212 (N_9212,N_9141,N_9108);
or U9213 (N_9213,N_9061,N_9161);
nor U9214 (N_9214,N_9054,N_9198);
xnor U9215 (N_9215,N_9127,N_9033);
xnor U9216 (N_9216,N_9090,N_9049);
xor U9217 (N_9217,N_9180,N_9082);
or U9218 (N_9218,N_9048,N_9126);
nand U9219 (N_9219,N_9105,N_9145);
xor U9220 (N_9220,N_9008,N_9191);
and U9221 (N_9221,N_9052,N_9011);
xor U9222 (N_9222,N_9186,N_9114);
nand U9223 (N_9223,N_9012,N_9159);
xor U9224 (N_9224,N_9063,N_9003);
xor U9225 (N_9225,N_9142,N_9021);
nand U9226 (N_9226,N_9146,N_9080);
xor U9227 (N_9227,N_9129,N_9109);
nand U9228 (N_9228,N_9122,N_9135);
nor U9229 (N_9229,N_9192,N_9024);
nor U9230 (N_9230,N_9091,N_9190);
nand U9231 (N_9231,N_9058,N_9013);
xor U9232 (N_9232,N_9179,N_9037);
xnor U9233 (N_9233,N_9099,N_9113);
xnor U9234 (N_9234,N_9199,N_9047);
and U9235 (N_9235,N_9025,N_9005);
nand U9236 (N_9236,N_9039,N_9112);
nor U9237 (N_9237,N_9034,N_9162);
xnor U9238 (N_9238,N_9177,N_9163);
nor U9239 (N_9239,N_9043,N_9015);
and U9240 (N_9240,N_9194,N_9132);
nand U9241 (N_9241,N_9157,N_9137);
or U9242 (N_9242,N_9140,N_9183);
and U9243 (N_9243,N_9086,N_9004);
and U9244 (N_9244,N_9035,N_9017);
or U9245 (N_9245,N_9060,N_9066);
nand U9246 (N_9246,N_9154,N_9168);
xnor U9247 (N_9247,N_9056,N_9019);
and U9248 (N_9248,N_9081,N_9195);
xor U9249 (N_9249,N_9184,N_9107);
nand U9250 (N_9250,N_9156,N_9124);
nand U9251 (N_9251,N_9149,N_9032);
xnor U9252 (N_9252,N_9152,N_9065);
nor U9253 (N_9253,N_9053,N_9116);
and U9254 (N_9254,N_9169,N_9036);
and U9255 (N_9255,N_9087,N_9153);
and U9256 (N_9256,N_9164,N_9150);
nand U9257 (N_9257,N_9187,N_9170);
nor U9258 (N_9258,N_9028,N_9044);
and U9259 (N_9259,N_9051,N_9062);
xnor U9260 (N_9260,N_9185,N_9040);
and U9261 (N_9261,N_9002,N_9174);
and U9262 (N_9262,N_9128,N_9023);
nand U9263 (N_9263,N_9075,N_9133);
nor U9264 (N_9264,N_9171,N_9144);
or U9265 (N_9265,N_9026,N_9104);
and U9266 (N_9266,N_9092,N_9070);
xor U9267 (N_9267,N_9073,N_9115);
nand U9268 (N_9268,N_9134,N_9098);
xnor U9269 (N_9269,N_9175,N_9097);
nand U9270 (N_9270,N_9136,N_9176);
or U9271 (N_9271,N_9057,N_9077);
nor U9272 (N_9272,N_9178,N_9046);
nand U9273 (N_9273,N_9100,N_9130);
nor U9274 (N_9274,N_9165,N_9088);
nor U9275 (N_9275,N_9181,N_9010);
or U9276 (N_9276,N_9038,N_9173);
nor U9277 (N_9277,N_9064,N_9155);
or U9278 (N_9278,N_9151,N_9160);
nand U9279 (N_9279,N_9196,N_9117);
or U9280 (N_9280,N_9096,N_9110);
nand U9281 (N_9281,N_9083,N_9016);
xnor U9282 (N_9282,N_9045,N_9055);
nor U9283 (N_9283,N_9018,N_9125);
and U9284 (N_9284,N_9148,N_9158);
or U9285 (N_9285,N_9131,N_9103);
xnor U9286 (N_9286,N_9072,N_9084);
xor U9287 (N_9287,N_9167,N_9089);
or U9288 (N_9288,N_9172,N_9067);
nor U9289 (N_9289,N_9074,N_9118);
and U9290 (N_9290,N_9006,N_9014);
xor U9291 (N_9291,N_9078,N_9041);
and U9292 (N_9292,N_9001,N_9197);
xor U9293 (N_9293,N_9143,N_9123);
and U9294 (N_9294,N_9095,N_9076);
nand U9295 (N_9295,N_9138,N_9120);
nand U9296 (N_9296,N_9007,N_9068);
or U9297 (N_9297,N_9182,N_9031);
or U9298 (N_9298,N_9022,N_9009);
xor U9299 (N_9299,N_9020,N_9166);
xnor U9300 (N_9300,N_9151,N_9038);
xnor U9301 (N_9301,N_9158,N_9193);
and U9302 (N_9302,N_9188,N_9018);
and U9303 (N_9303,N_9013,N_9129);
and U9304 (N_9304,N_9161,N_9013);
nor U9305 (N_9305,N_9192,N_9157);
nor U9306 (N_9306,N_9158,N_9050);
and U9307 (N_9307,N_9062,N_9094);
nand U9308 (N_9308,N_9130,N_9121);
nor U9309 (N_9309,N_9053,N_9000);
nand U9310 (N_9310,N_9050,N_9134);
and U9311 (N_9311,N_9017,N_9039);
or U9312 (N_9312,N_9010,N_9171);
nand U9313 (N_9313,N_9076,N_9160);
nor U9314 (N_9314,N_9192,N_9112);
and U9315 (N_9315,N_9113,N_9042);
nand U9316 (N_9316,N_9158,N_9042);
xnor U9317 (N_9317,N_9142,N_9017);
nor U9318 (N_9318,N_9061,N_9005);
and U9319 (N_9319,N_9029,N_9055);
and U9320 (N_9320,N_9194,N_9111);
nor U9321 (N_9321,N_9160,N_9036);
nor U9322 (N_9322,N_9085,N_9120);
nand U9323 (N_9323,N_9187,N_9135);
nor U9324 (N_9324,N_9079,N_9183);
nand U9325 (N_9325,N_9048,N_9079);
or U9326 (N_9326,N_9185,N_9138);
nor U9327 (N_9327,N_9032,N_9189);
nor U9328 (N_9328,N_9184,N_9112);
xnor U9329 (N_9329,N_9195,N_9136);
nand U9330 (N_9330,N_9013,N_9179);
nand U9331 (N_9331,N_9153,N_9195);
xor U9332 (N_9332,N_9061,N_9108);
or U9333 (N_9333,N_9026,N_9173);
nor U9334 (N_9334,N_9166,N_9022);
and U9335 (N_9335,N_9182,N_9032);
and U9336 (N_9336,N_9019,N_9034);
and U9337 (N_9337,N_9141,N_9085);
or U9338 (N_9338,N_9069,N_9186);
or U9339 (N_9339,N_9107,N_9174);
xnor U9340 (N_9340,N_9073,N_9128);
nor U9341 (N_9341,N_9125,N_9073);
and U9342 (N_9342,N_9140,N_9148);
nand U9343 (N_9343,N_9189,N_9020);
nor U9344 (N_9344,N_9134,N_9118);
xor U9345 (N_9345,N_9117,N_9069);
or U9346 (N_9346,N_9035,N_9086);
nand U9347 (N_9347,N_9066,N_9054);
nor U9348 (N_9348,N_9172,N_9100);
and U9349 (N_9349,N_9062,N_9008);
nand U9350 (N_9350,N_9068,N_9128);
nand U9351 (N_9351,N_9195,N_9196);
or U9352 (N_9352,N_9133,N_9107);
xor U9353 (N_9353,N_9168,N_9043);
xor U9354 (N_9354,N_9013,N_9173);
nor U9355 (N_9355,N_9193,N_9126);
or U9356 (N_9356,N_9183,N_9077);
xor U9357 (N_9357,N_9133,N_9039);
and U9358 (N_9358,N_9022,N_9122);
or U9359 (N_9359,N_9162,N_9054);
and U9360 (N_9360,N_9072,N_9019);
xor U9361 (N_9361,N_9163,N_9100);
or U9362 (N_9362,N_9130,N_9052);
or U9363 (N_9363,N_9048,N_9103);
or U9364 (N_9364,N_9041,N_9075);
nand U9365 (N_9365,N_9150,N_9126);
nor U9366 (N_9366,N_9123,N_9020);
nor U9367 (N_9367,N_9148,N_9007);
nor U9368 (N_9368,N_9187,N_9003);
xnor U9369 (N_9369,N_9164,N_9026);
and U9370 (N_9370,N_9075,N_9003);
xor U9371 (N_9371,N_9033,N_9077);
or U9372 (N_9372,N_9106,N_9158);
xor U9373 (N_9373,N_9106,N_9012);
and U9374 (N_9374,N_9132,N_9004);
nand U9375 (N_9375,N_9072,N_9175);
xor U9376 (N_9376,N_9149,N_9195);
or U9377 (N_9377,N_9119,N_9054);
nand U9378 (N_9378,N_9050,N_9172);
xnor U9379 (N_9379,N_9074,N_9038);
and U9380 (N_9380,N_9124,N_9157);
nand U9381 (N_9381,N_9000,N_9079);
nor U9382 (N_9382,N_9153,N_9180);
xnor U9383 (N_9383,N_9061,N_9062);
nor U9384 (N_9384,N_9144,N_9165);
xor U9385 (N_9385,N_9049,N_9170);
or U9386 (N_9386,N_9135,N_9192);
nor U9387 (N_9387,N_9005,N_9014);
or U9388 (N_9388,N_9111,N_9124);
xnor U9389 (N_9389,N_9065,N_9176);
and U9390 (N_9390,N_9059,N_9030);
nor U9391 (N_9391,N_9022,N_9154);
nor U9392 (N_9392,N_9023,N_9064);
nor U9393 (N_9393,N_9187,N_9152);
nand U9394 (N_9394,N_9065,N_9020);
or U9395 (N_9395,N_9147,N_9132);
xnor U9396 (N_9396,N_9178,N_9153);
xnor U9397 (N_9397,N_9198,N_9069);
xor U9398 (N_9398,N_9134,N_9047);
nand U9399 (N_9399,N_9069,N_9103);
xnor U9400 (N_9400,N_9289,N_9384);
nor U9401 (N_9401,N_9242,N_9363);
or U9402 (N_9402,N_9315,N_9306);
or U9403 (N_9403,N_9391,N_9371);
or U9404 (N_9404,N_9308,N_9292);
xor U9405 (N_9405,N_9235,N_9320);
xnor U9406 (N_9406,N_9309,N_9253);
nand U9407 (N_9407,N_9390,N_9265);
nor U9408 (N_9408,N_9204,N_9297);
nor U9409 (N_9409,N_9331,N_9239);
or U9410 (N_9410,N_9268,N_9375);
nor U9411 (N_9411,N_9367,N_9252);
and U9412 (N_9412,N_9365,N_9323);
or U9413 (N_9413,N_9376,N_9351);
and U9414 (N_9414,N_9291,N_9314);
or U9415 (N_9415,N_9219,N_9311);
xnor U9416 (N_9416,N_9322,N_9318);
or U9417 (N_9417,N_9262,N_9260);
or U9418 (N_9418,N_9237,N_9233);
and U9419 (N_9419,N_9283,N_9230);
nor U9420 (N_9420,N_9250,N_9218);
xor U9421 (N_9421,N_9298,N_9310);
or U9422 (N_9422,N_9330,N_9301);
xor U9423 (N_9423,N_9223,N_9340);
or U9424 (N_9424,N_9381,N_9312);
nand U9425 (N_9425,N_9225,N_9334);
xor U9426 (N_9426,N_9339,N_9361);
nor U9427 (N_9427,N_9395,N_9202);
xnor U9428 (N_9428,N_9290,N_9399);
or U9429 (N_9429,N_9373,N_9279);
and U9430 (N_9430,N_9336,N_9208);
or U9431 (N_9431,N_9261,N_9378);
xnor U9432 (N_9432,N_9387,N_9241);
nor U9433 (N_9433,N_9353,N_9350);
nor U9434 (N_9434,N_9358,N_9248);
nand U9435 (N_9435,N_9328,N_9343);
xnor U9436 (N_9436,N_9313,N_9201);
and U9437 (N_9437,N_9346,N_9272);
nand U9438 (N_9438,N_9282,N_9394);
xor U9439 (N_9439,N_9374,N_9277);
nor U9440 (N_9440,N_9303,N_9359);
and U9441 (N_9441,N_9305,N_9333);
or U9442 (N_9442,N_9229,N_9338);
nor U9443 (N_9443,N_9231,N_9299);
xor U9444 (N_9444,N_9383,N_9256);
nand U9445 (N_9445,N_9293,N_9295);
xor U9446 (N_9446,N_9222,N_9213);
nand U9447 (N_9447,N_9388,N_9352);
xor U9448 (N_9448,N_9246,N_9389);
or U9449 (N_9449,N_9232,N_9212);
and U9450 (N_9450,N_9326,N_9258);
nor U9451 (N_9451,N_9294,N_9217);
xor U9452 (N_9452,N_9362,N_9270);
nor U9453 (N_9453,N_9273,N_9251);
and U9454 (N_9454,N_9206,N_9370);
or U9455 (N_9455,N_9327,N_9284);
nor U9456 (N_9456,N_9224,N_9348);
xor U9457 (N_9457,N_9354,N_9203);
and U9458 (N_9458,N_9349,N_9238);
or U9459 (N_9459,N_9274,N_9227);
nor U9460 (N_9460,N_9304,N_9243);
and U9461 (N_9461,N_9382,N_9216);
xnor U9462 (N_9462,N_9316,N_9357);
or U9463 (N_9463,N_9211,N_9356);
nand U9464 (N_9464,N_9377,N_9386);
or U9465 (N_9465,N_9259,N_9278);
and U9466 (N_9466,N_9337,N_9200);
nand U9467 (N_9467,N_9286,N_9267);
or U9468 (N_9468,N_9335,N_9266);
nand U9469 (N_9469,N_9214,N_9285);
xor U9470 (N_9470,N_9302,N_9379);
and U9471 (N_9471,N_9210,N_9236);
nor U9472 (N_9472,N_9226,N_9254);
nor U9473 (N_9473,N_9275,N_9247);
and U9474 (N_9474,N_9344,N_9398);
and U9475 (N_9475,N_9347,N_9325);
nand U9476 (N_9476,N_9307,N_9355);
xnor U9477 (N_9477,N_9341,N_9221);
nand U9478 (N_9478,N_9296,N_9245);
nor U9479 (N_9479,N_9324,N_9255);
nor U9480 (N_9480,N_9385,N_9228);
xor U9481 (N_9481,N_9269,N_9345);
nand U9482 (N_9482,N_9209,N_9205);
nand U9483 (N_9483,N_9396,N_9207);
or U9484 (N_9484,N_9368,N_9319);
nand U9485 (N_9485,N_9234,N_9372);
nor U9486 (N_9486,N_9280,N_9281);
nor U9487 (N_9487,N_9244,N_9257);
or U9488 (N_9488,N_9215,N_9300);
xnor U9489 (N_9489,N_9271,N_9276);
and U9490 (N_9490,N_9240,N_9264);
or U9491 (N_9491,N_9263,N_9287);
nor U9492 (N_9492,N_9380,N_9288);
nor U9493 (N_9493,N_9332,N_9321);
nand U9494 (N_9494,N_9364,N_9220);
nand U9495 (N_9495,N_9360,N_9249);
and U9496 (N_9496,N_9366,N_9397);
and U9497 (N_9497,N_9369,N_9329);
xnor U9498 (N_9498,N_9392,N_9393);
nand U9499 (N_9499,N_9317,N_9342);
nand U9500 (N_9500,N_9298,N_9234);
and U9501 (N_9501,N_9249,N_9250);
nor U9502 (N_9502,N_9316,N_9312);
or U9503 (N_9503,N_9328,N_9356);
and U9504 (N_9504,N_9241,N_9374);
xnor U9505 (N_9505,N_9210,N_9340);
or U9506 (N_9506,N_9249,N_9217);
xnor U9507 (N_9507,N_9200,N_9321);
or U9508 (N_9508,N_9287,N_9341);
and U9509 (N_9509,N_9354,N_9358);
or U9510 (N_9510,N_9217,N_9263);
nand U9511 (N_9511,N_9383,N_9252);
and U9512 (N_9512,N_9374,N_9295);
xor U9513 (N_9513,N_9245,N_9331);
nor U9514 (N_9514,N_9260,N_9349);
xnor U9515 (N_9515,N_9309,N_9345);
xnor U9516 (N_9516,N_9354,N_9392);
and U9517 (N_9517,N_9383,N_9290);
and U9518 (N_9518,N_9267,N_9364);
nand U9519 (N_9519,N_9372,N_9340);
and U9520 (N_9520,N_9213,N_9258);
nor U9521 (N_9521,N_9247,N_9249);
and U9522 (N_9522,N_9258,N_9352);
nor U9523 (N_9523,N_9372,N_9303);
or U9524 (N_9524,N_9289,N_9284);
and U9525 (N_9525,N_9282,N_9378);
and U9526 (N_9526,N_9354,N_9286);
and U9527 (N_9527,N_9258,N_9374);
or U9528 (N_9528,N_9324,N_9398);
xnor U9529 (N_9529,N_9277,N_9351);
nor U9530 (N_9530,N_9293,N_9226);
or U9531 (N_9531,N_9392,N_9223);
xor U9532 (N_9532,N_9345,N_9301);
nand U9533 (N_9533,N_9308,N_9296);
or U9534 (N_9534,N_9238,N_9308);
xnor U9535 (N_9535,N_9284,N_9203);
nand U9536 (N_9536,N_9339,N_9303);
nor U9537 (N_9537,N_9331,N_9233);
or U9538 (N_9538,N_9386,N_9276);
or U9539 (N_9539,N_9218,N_9362);
nand U9540 (N_9540,N_9286,N_9279);
or U9541 (N_9541,N_9361,N_9300);
and U9542 (N_9542,N_9264,N_9278);
xor U9543 (N_9543,N_9371,N_9374);
and U9544 (N_9544,N_9306,N_9282);
nand U9545 (N_9545,N_9248,N_9359);
nand U9546 (N_9546,N_9318,N_9233);
and U9547 (N_9547,N_9205,N_9366);
xnor U9548 (N_9548,N_9212,N_9382);
xnor U9549 (N_9549,N_9337,N_9221);
xnor U9550 (N_9550,N_9388,N_9293);
nor U9551 (N_9551,N_9254,N_9216);
or U9552 (N_9552,N_9341,N_9298);
xnor U9553 (N_9553,N_9221,N_9279);
xnor U9554 (N_9554,N_9399,N_9346);
nand U9555 (N_9555,N_9308,N_9298);
nand U9556 (N_9556,N_9200,N_9300);
or U9557 (N_9557,N_9376,N_9361);
nand U9558 (N_9558,N_9394,N_9285);
xor U9559 (N_9559,N_9321,N_9396);
or U9560 (N_9560,N_9212,N_9372);
and U9561 (N_9561,N_9259,N_9250);
xnor U9562 (N_9562,N_9352,N_9380);
xor U9563 (N_9563,N_9304,N_9289);
xor U9564 (N_9564,N_9273,N_9302);
xor U9565 (N_9565,N_9358,N_9357);
nand U9566 (N_9566,N_9347,N_9312);
or U9567 (N_9567,N_9370,N_9332);
nor U9568 (N_9568,N_9212,N_9252);
nand U9569 (N_9569,N_9244,N_9245);
and U9570 (N_9570,N_9356,N_9266);
or U9571 (N_9571,N_9323,N_9216);
or U9572 (N_9572,N_9330,N_9231);
nand U9573 (N_9573,N_9235,N_9346);
nor U9574 (N_9574,N_9206,N_9201);
and U9575 (N_9575,N_9332,N_9232);
nand U9576 (N_9576,N_9277,N_9389);
nand U9577 (N_9577,N_9200,N_9389);
and U9578 (N_9578,N_9243,N_9273);
and U9579 (N_9579,N_9300,N_9228);
nand U9580 (N_9580,N_9284,N_9282);
and U9581 (N_9581,N_9211,N_9202);
nor U9582 (N_9582,N_9365,N_9285);
nor U9583 (N_9583,N_9259,N_9237);
xor U9584 (N_9584,N_9205,N_9275);
and U9585 (N_9585,N_9205,N_9298);
nand U9586 (N_9586,N_9239,N_9247);
nand U9587 (N_9587,N_9259,N_9332);
nor U9588 (N_9588,N_9247,N_9228);
and U9589 (N_9589,N_9304,N_9366);
xor U9590 (N_9590,N_9351,N_9231);
or U9591 (N_9591,N_9345,N_9234);
nor U9592 (N_9592,N_9263,N_9362);
and U9593 (N_9593,N_9316,N_9326);
nor U9594 (N_9594,N_9268,N_9286);
or U9595 (N_9595,N_9320,N_9221);
nor U9596 (N_9596,N_9225,N_9389);
xnor U9597 (N_9597,N_9294,N_9363);
or U9598 (N_9598,N_9312,N_9281);
nor U9599 (N_9599,N_9333,N_9249);
nor U9600 (N_9600,N_9583,N_9506);
xor U9601 (N_9601,N_9539,N_9490);
xnor U9602 (N_9602,N_9405,N_9439);
or U9603 (N_9603,N_9530,N_9551);
and U9604 (N_9604,N_9521,N_9538);
nand U9605 (N_9605,N_9574,N_9416);
or U9606 (N_9606,N_9565,N_9514);
and U9607 (N_9607,N_9430,N_9508);
nand U9608 (N_9608,N_9510,N_9562);
or U9609 (N_9609,N_9426,N_9444);
or U9610 (N_9610,N_9504,N_9517);
xor U9611 (N_9611,N_9576,N_9423);
or U9612 (N_9612,N_9455,N_9590);
or U9613 (N_9613,N_9499,N_9437);
xnor U9614 (N_9614,N_9594,N_9404);
and U9615 (N_9615,N_9467,N_9407);
or U9616 (N_9616,N_9408,N_9497);
and U9617 (N_9617,N_9520,N_9401);
or U9618 (N_9618,N_9535,N_9546);
nand U9619 (N_9619,N_9454,N_9446);
and U9620 (N_9620,N_9534,N_9585);
xnor U9621 (N_9621,N_9559,N_9478);
nor U9622 (N_9622,N_9457,N_9588);
or U9623 (N_9623,N_9553,N_9519);
xnor U9624 (N_9624,N_9440,N_9509);
nor U9625 (N_9625,N_9463,N_9477);
nand U9626 (N_9626,N_9568,N_9593);
nor U9627 (N_9627,N_9525,N_9481);
nor U9628 (N_9628,N_9484,N_9411);
xnor U9629 (N_9629,N_9458,N_9507);
and U9630 (N_9630,N_9487,N_9533);
or U9631 (N_9631,N_9464,N_9545);
nor U9632 (N_9632,N_9438,N_9433);
xnor U9633 (N_9633,N_9480,N_9575);
nor U9634 (N_9634,N_9406,N_9472);
and U9635 (N_9635,N_9500,N_9486);
and U9636 (N_9636,N_9549,N_9435);
and U9637 (N_9637,N_9536,N_9459);
nand U9638 (N_9638,N_9541,N_9427);
nor U9639 (N_9639,N_9428,N_9456);
or U9640 (N_9640,N_9471,N_9563);
or U9641 (N_9641,N_9577,N_9502);
and U9642 (N_9642,N_9445,N_9578);
nor U9643 (N_9643,N_9400,N_9528);
or U9644 (N_9644,N_9451,N_9489);
xnor U9645 (N_9645,N_9473,N_9526);
xor U9646 (N_9646,N_9548,N_9552);
and U9647 (N_9647,N_9547,N_9479);
or U9648 (N_9648,N_9431,N_9449);
or U9649 (N_9649,N_9544,N_9542);
nor U9650 (N_9650,N_9598,N_9410);
nand U9651 (N_9651,N_9529,N_9409);
nand U9652 (N_9652,N_9524,N_9492);
or U9653 (N_9653,N_9572,N_9554);
or U9654 (N_9654,N_9579,N_9589);
or U9655 (N_9655,N_9503,N_9403);
nor U9656 (N_9656,N_9596,N_9418);
nor U9657 (N_9657,N_9569,N_9470);
and U9658 (N_9658,N_9452,N_9475);
xor U9659 (N_9659,N_9532,N_9441);
nand U9660 (N_9660,N_9581,N_9450);
and U9661 (N_9661,N_9550,N_9573);
or U9662 (N_9662,N_9560,N_9496);
or U9663 (N_9663,N_9498,N_9420);
or U9664 (N_9664,N_9580,N_9527);
and U9665 (N_9665,N_9586,N_9402);
or U9666 (N_9666,N_9488,N_9522);
nand U9667 (N_9667,N_9422,N_9424);
nand U9668 (N_9668,N_9436,N_9462);
nand U9669 (N_9669,N_9469,N_9564);
and U9670 (N_9670,N_9434,N_9555);
and U9671 (N_9671,N_9592,N_9465);
nand U9672 (N_9672,N_9442,N_9556);
nor U9673 (N_9673,N_9505,N_9494);
xor U9674 (N_9674,N_9466,N_9425);
and U9675 (N_9675,N_9482,N_9414);
or U9676 (N_9676,N_9476,N_9558);
or U9677 (N_9677,N_9483,N_9537);
nand U9678 (N_9678,N_9493,N_9468);
xnor U9679 (N_9679,N_9432,N_9557);
or U9680 (N_9680,N_9495,N_9421);
nand U9681 (N_9681,N_9515,N_9523);
and U9682 (N_9682,N_9460,N_9429);
xnor U9683 (N_9683,N_9448,N_9567);
nand U9684 (N_9684,N_9531,N_9511);
xor U9685 (N_9685,N_9582,N_9571);
or U9686 (N_9686,N_9443,N_9461);
nor U9687 (N_9687,N_9587,N_9412);
nor U9688 (N_9688,N_9474,N_9540);
nand U9689 (N_9689,N_9599,N_9561);
nor U9690 (N_9690,N_9543,N_9413);
or U9691 (N_9691,N_9518,N_9512);
nor U9692 (N_9692,N_9491,N_9595);
nor U9693 (N_9693,N_9501,N_9566);
nand U9694 (N_9694,N_9447,N_9417);
xnor U9695 (N_9695,N_9453,N_9584);
nand U9696 (N_9696,N_9570,N_9597);
and U9697 (N_9697,N_9419,N_9516);
and U9698 (N_9698,N_9591,N_9415);
xor U9699 (N_9699,N_9513,N_9485);
nor U9700 (N_9700,N_9439,N_9597);
and U9701 (N_9701,N_9534,N_9565);
or U9702 (N_9702,N_9520,N_9534);
nor U9703 (N_9703,N_9416,N_9438);
xnor U9704 (N_9704,N_9504,N_9554);
xnor U9705 (N_9705,N_9509,N_9482);
xnor U9706 (N_9706,N_9551,N_9404);
nor U9707 (N_9707,N_9428,N_9418);
nand U9708 (N_9708,N_9580,N_9536);
xnor U9709 (N_9709,N_9463,N_9584);
nand U9710 (N_9710,N_9459,N_9522);
xnor U9711 (N_9711,N_9452,N_9473);
xor U9712 (N_9712,N_9429,N_9573);
nor U9713 (N_9713,N_9591,N_9460);
xnor U9714 (N_9714,N_9465,N_9519);
and U9715 (N_9715,N_9504,N_9555);
and U9716 (N_9716,N_9480,N_9511);
nor U9717 (N_9717,N_9403,N_9434);
xor U9718 (N_9718,N_9506,N_9550);
nor U9719 (N_9719,N_9436,N_9458);
or U9720 (N_9720,N_9548,N_9484);
xnor U9721 (N_9721,N_9461,N_9402);
and U9722 (N_9722,N_9404,N_9523);
nor U9723 (N_9723,N_9425,N_9539);
nand U9724 (N_9724,N_9554,N_9556);
and U9725 (N_9725,N_9557,N_9456);
nand U9726 (N_9726,N_9503,N_9453);
nor U9727 (N_9727,N_9489,N_9562);
nand U9728 (N_9728,N_9492,N_9581);
and U9729 (N_9729,N_9436,N_9404);
or U9730 (N_9730,N_9573,N_9509);
nand U9731 (N_9731,N_9489,N_9572);
and U9732 (N_9732,N_9598,N_9458);
or U9733 (N_9733,N_9451,N_9414);
nand U9734 (N_9734,N_9576,N_9562);
nand U9735 (N_9735,N_9411,N_9473);
nor U9736 (N_9736,N_9521,N_9429);
xor U9737 (N_9737,N_9421,N_9493);
or U9738 (N_9738,N_9427,N_9474);
xor U9739 (N_9739,N_9521,N_9585);
or U9740 (N_9740,N_9497,N_9518);
nand U9741 (N_9741,N_9424,N_9414);
nand U9742 (N_9742,N_9432,N_9425);
nor U9743 (N_9743,N_9406,N_9453);
nor U9744 (N_9744,N_9542,N_9583);
or U9745 (N_9745,N_9518,N_9553);
and U9746 (N_9746,N_9537,N_9523);
nand U9747 (N_9747,N_9445,N_9542);
nor U9748 (N_9748,N_9465,N_9554);
and U9749 (N_9749,N_9486,N_9419);
and U9750 (N_9750,N_9547,N_9447);
xnor U9751 (N_9751,N_9410,N_9535);
nor U9752 (N_9752,N_9412,N_9407);
or U9753 (N_9753,N_9576,N_9531);
nand U9754 (N_9754,N_9548,N_9587);
xnor U9755 (N_9755,N_9584,N_9461);
xnor U9756 (N_9756,N_9509,N_9401);
and U9757 (N_9757,N_9552,N_9592);
xor U9758 (N_9758,N_9553,N_9534);
xnor U9759 (N_9759,N_9571,N_9526);
or U9760 (N_9760,N_9539,N_9475);
nor U9761 (N_9761,N_9481,N_9428);
or U9762 (N_9762,N_9400,N_9491);
nor U9763 (N_9763,N_9421,N_9521);
and U9764 (N_9764,N_9430,N_9457);
nor U9765 (N_9765,N_9462,N_9582);
and U9766 (N_9766,N_9457,N_9489);
and U9767 (N_9767,N_9526,N_9452);
nor U9768 (N_9768,N_9588,N_9572);
nor U9769 (N_9769,N_9556,N_9512);
and U9770 (N_9770,N_9592,N_9530);
xnor U9771 (N_9771,N_9479,N_9518);
or U9772 (N_9772,N_9473,N_9443);
nand U9773 (N_9773,N_9565,N_9463);
or U9774 (N_9774,N_9454,N_9577);
or U9775 (N_9775,N_9549,N_9502);
or U9776 (N_9776,N_9585,N_9574);
nand U9777 (N_9777,N_9414,N_9531);
nand U9778 (N_9778,N_9502,N_9535);
nand U9779 (N_9779,N_9569,N_9547);
and U9780 (N_9780,N_9462,N_9449);
or U9781 (N_9781,N_9432,N_9552);
and U9782 (N_9782,N_9530,N_9506);
nand U9783 (N_9783,N_9457,N_9466);
nor U9784 (N_9784,N_9416,N_9500);
nand U9785 (N_9785,N_9566,N_9405);
nand U9786 (N_9786,N_9475,N_9569);
nand U9787 (N_9787,N_9535,N_9446);
xor U9788 (N_9788,N_9497,N_9548);
nor U9789 (N_9789,N_9522,N_9590);
or U9790 (N_9790,N_9469,N_9449);
xor U9791 (N_9791,N_9528,N_9565);
nand U9792 (N_9792,N_9462,N_9492);
xor U9793 (N_9793,N_9585,N_9465);
nor U9794 (N_9794,N_9425,N_9479);
nor U9795 (N_9795,N_9530,N_9526);
or U9796 (N_9796,N_9522,N_9408);
or U9797 (N_9797,N_9554,N_9431);
xnor U9798 (N_9798,N_9517,N_9570);
nand U9799 (N_9799,N_9563,N_9526);
or U9800 (N_9800,N_9616,N_9708);
and U9801 (N_9801,N_9675,N_9662);
nand U9802 (N_9802,N_9628,N_9603);
nor U9803 (N_9803,N_9646,N_9797);
xnor U9804 (N_9804,N_9631,N_9650);
or U9805 (N_9805,N_9767,N_9749);
or U9806 (N_9806,N_9686,N_9752);
nor U9807 (N_9807,N_9746,N_9637);
nor U9808 (N_9808,N_9756,N_9698);
xnor U9809 (N_9809,N_9725,N_9744);
nor U9810 (N_9810,N_9727,N_9694);
xor U9811 (N_9811,N_9717,N_9635);
nand U9812 (N_9812,N_9697,N_9607);
nand U9813 (N_9813,N_9782,N_9762);
nor U9814 (N_9814,N_9633,N_9769);
or U9815 (N_9815,N_9757,N_9645);
or U9816 (N_9816,N_9795,N_9670);
nand U9817 (N_9817,N_9639,N_9719);
nand U9818 (N_9818,N_9617,N_9705);
and U9819 (N_9819,N_9684,N_9702);
nor U9820 (N_9820,N_9612,N_9636);
nor U9821 (N_9821,N_9766,N_9679);
xor U9822 (N_9822,N_9671,N_9732);
nor U9823 (N_9823,N_9680,N_9601);
xor U9824 (N_9824,N_9784,N_9640);
nor U9825 (N_9825,N_9786,N_9739);
or U9826 (N_9826,N_9647,N_9785);
nand U9827 (N_9827,N_9693,N_9642);
and U9828 (N_9828,N_9622,N_9729);
nand U9829 (N_9829,N_9674,N_9665);
nor U9830 (N_9830,N_9711,N_9737);
xnor U9831 (N_9831,N_9666,N_9663);
and U9832 (N_9832,N_9677,N_9676);
and U9833 (N_9833,N_9632,N_9721);
nand U9834 (N_9834,N_9761,N_9602);
xnor U9835 (N_9835,N_9715,N_9611);
xnor U9836 (N_9836,N_9690,N_9687);
xnor U9837 (N_9837,N_9668,N_9672);
nor U9838 (N_9838,N_9630,N_9692);
nand U9839 (N_9839,N_9629,N_9753);
or U9840 (N_9840,N_9652,N_9726);
nand U9841 (N_9841,N_9704,N_9714);
and U9842 (N_9842,N_9619,N_9728);
or U9843 (N_9843,N_9710,N_9758);
xnor U9844 (N_9844,N_9787,N_9649);
and U9845 (N_9845,N_9775,N_9655);
nor U9846 (N_9846,N_9641,N_9618);
nand U9847 (N_9847,N_9667,N_9709);
or U9848 (N_9848,N_9688,N_9735);
nor U9849 (N_9849,N_9754,N_9738);
and U9850 (N_9850,N_9643,N_9627);
nand U9851 (N_9851,N_9760,N_9659);
xor U9852 (N_9852,N_9742,N_9763);
nor U9853 (N_9853,N_9747,N_9773);
nand U9854 (N_9854,N_9712,N_9625);
nor U9855 (N_9855,N_9789,N_9771);
or U9856 (N_9856,N_9736,N_9722);
xnor U9857 (N_9857,N_9613,N_9609);
xor U9858 (N_9858,N_9774,N_9793);
or U9859 (N_9859,N_9730,N_9794);
nor U9860 (N_9860,N_9673,N_9706);
xnor U9861 (N_9861,N_9720,N_9623);
nor U9862 (N_9862,N_9798,N_9707);
nor U9863 (N_9863,N_9654,N_9634);
nor U9864 (N_9864,N_9755,N_9734);
or U9865 (N_9865,N_9678,N_9703);
nor U9866 (N_9866,N_9751,N_9724);
xnor U9867 (N_9867,N_9750,N_9685);
nor U9868 (N_9868,N_9764,N_9791);
nor U9869 (N_9869,N_9606,N_9689);
or U9870 (N_9870,N_9740,N_9661);
or U9871 (N_9871,N_9792,N_9648);
nor U9872 (N_9872,N_9620,N_9695);
and U9873 (N_9873,N_9621,N_9781);
nor U9874 (N_9874,N_9600,N_9615);
nor U9875 (N_9875,N_9745,N_9682);
and U9876 (N_9876,N_9718,N_9731);
nand U9877 (N_9877,N_9776,N_9614);
and U9878 (N_9878,N_9658,N_9765);
nand U9879 (N_9879,N_9669,N_9657);
nand U9880 (N_9880,N_9696,N_9656);
xnor U9881 (N_9881,N_9664,N_9783);
nand U9882 (N_9882,N_9610,N_9796);
xor U9883 (N_9883,N_9605,N_9723);
and U9884 (N_9884,N_9780,N_9713);
or U9885 (N_9885,N_9691,N_9733);
or U9886 (N_9886,N_9604,N_9660);
or U9887 (N_9887,N_9716,N_9653);
nand U9888 (N_9888,N_9699,N_9741);
and U9889 (N_9889,N_9700,N_9701);
and U9890 (N_9890,N_9777,N_9626);
nand U9891 (N_9891,N_9608,N_9790);
or U9892 (N_9892,N_9624,N_9799);
or U9893 (N_9893,N_9768,N_9743);
and U9894 (N_9894,N_9759,N_9788);
nor U9895 (N_9895,N_9778,N_9651);
or U9896 (N_9896,N_9770,N_9644);
nor U9897 (N_9897,N_9638,N_9681);
and U9898 (N_9898,N_9748,N_9772);
nor U9899 (N_9899,N_9779,N_9683);
and U9900 (N_9900,N_9774,N_9719);
or U9901 (N_9901,N_9667,N_9689);
or U9902 (N_9902,N_9644,N_9702);
nand U9903 (N_9903,N_9624,N_9633);
xor U9904 (N_9904,N_9620,N_9716);
nand U9905 (N_9905,N_9653,N_9695);
nand U9906 (N_9906,N_9615,N_9750);
and U9907 (N_9907,N_9623,N_9714);
nor U9908 (N_9908,N_9713,N_9715);
nor U9909 (N_9909,N_9725,N_9675);
nand U9910 (N_9910,N_9658,N_9731);
xor U9911 (N_9911,N_9666,N_9611);
or U9912 (N_9912,N_9741,N_9766);
xnor U9913 (N_9913,N_9788,N_9662);
nand U9914 (N_9914,N_9619,N_9718);
xnor U9915 (N_9915,N_9735,N_9636);
or U9916 (N_9916,N_9734,N_9656);
nor U9917 (N_9917,N_9692,N_9666);
nor U9918 (N_9918,N_9759,N_9745);
and U9919 (N_9919,N_9609,N_9676);
nor U9920 (N_9920,N_9668,N_9634);
and U9921 (N_9921,N_9700,N_9782);
xnor U9922 (N_9922,N_9619,N_9635);
and U9923 (N_9923,N_9732,N_9620);
or U9924 (N_9924,N_9658,N_9778);
or U9925 (N_9925,N_9786,N_9753);
xnor U9926 (N_9926,N_9787,N_9625);
xor U9927 (N_9927,N_9684,N_9663);
or U9928 (N_9928,N_9757,N_9738);
nor U9929 (N_9929,N_9748,N_9771);
and U9930 (N_9930,N_9629,N_9670);
or U9931 (N_9931,N_9652,N_9600);
and U9932 (N_9932,N_9615,N_9611);
or U9933 (N_9933,N_9658,N_9689);
and U9934 (N_9934,N_9772,N_9663);
nand U9935 (N_9935,N_9682,N_9634);
nor U9936 (N_9936,N_9752,N_9719);
nand U9937 (N_9937,N_9606,N_9761);
xor U9938 (N_9938,N_9742,N_9722);
xnor U9939 (N_9939,N_9745,N_9619);
nor U9940 (N_9940,N_9709,N_9674);
xor U9941 (N_9941,N_9645,N_9736);
nand U9942 (N_9942,N_9631,N_9750);
nor U9943 (N_9943,N_9736,N_9750);
or U9944 (N_9944,N_9774,N_9704);
or U9945 (N_9945,N_9799,N_9646);
xor U9946 (N_9946,N_9725,N_9709);
or U9947 (N_9947,N_9783,N_9698);
xnor U9948 (N_9948,N_9712,N_9611);
or U9949 (N_9949,N_9682,N_9614);
and U9950 (N_9950,N_9666,N_9787);
and U9951 (N_9951,N_9711,N_9790);
xnor U9952 (N_9952,N_9744,N_9685);
or U9953 (N_9953,N_9711,N_9748);
and U9954 (N_9954,N_9620,N_9749);
nor U9955 (N_9955,N_9694,N_9783);
or U9956 (N_9956,N_9689,N_9796);
nor U9957 (N_9957,N_9707,N_9626);
and U9958 (N_9958,N_9664,N_9741);
nor U9959 (N_9959,N_9771,N_9667);
or U9960 (N_9960,N_9744,N_9711);
or U9961 (N_9961,N_9625,N_9678);
xor U9962 (N_9962,N_9600,N_9724);
or U9963 (N_9963,N_9662,N_9614);
nand U9964 (N_9964,N_9633,N_9673);
xnor U9965 (N_9965,N_9790,N_9770);
or U9966 (N_9966,N_9709,N_9768);
and U9967 (N_9967,N_9719,N_9621);
or U9968 (N_9968,N_9773,N_9656);
nand U9969 (N_9969,N_9616,N_9753);
xnor U9970 (N_9970,N_9775,N_9657);
xor U9971 (N_9971,N_9639,N_9798);
or U9972 (N_9972,N_9674,N_9627);
and U9973 (N_9973,N_9656,N_9659);
and U9974 (N_9974,N_9682,N_9638);
nor U9975 (N_9975,N_9674,N_9697);
and U9976 (N_9976,N_9623,N_9627);
nand U9977 (N_9977,N_9657,N_9787);
nor U9978 (N_9978,N_9666,N_9646);
nor U9979 (N_9979,N_9703,N_9638);
nand U9980 (N_9980,N_9732,N_9786);
xor U9981 (N_9981,N_9755,N_9737);
xor U9982 (N_9982,N_9630,N_9640);
and U9983 (N_9983,N_9766,N_9789);
nor U9984 (N_9984,N_9733,N_9678);
or U9985 (N_9985,N_9727,N_9783);
nand U9986 (N_9986,N_9634,N_9646);
or U9987 (N_9987,N_9613,N_9634);
xnor U9988 (N_9988,N_9737,N_9622);
xor U9989 (N_9989,N_9686,N_9677);
nor U9990 (N_9990,N_9668,N_9688);
and U9991 (N_9991,N_9648,N_9758);
nor U9992 (N_9992,N_9635,N_9629);
nor U9993 (N_9993,N_9691,N_9615);
nor U9994 (N_9994,N_9632,N_9680);
or U9995 (N_9995,N_9784,N_9751);
nor U9996 (N_9996,N_9799,N_9648);
xor U9997 (N_9997,N_9660,N_9762);
nor U9998 (N_9998,N_9718,N_9698);
and U9999 (N_9999,N_9692,N_9707);
xor U10000 (N_10000,N_9884,N_9956);
and U10001 (N_10001,N_9936,N_9817);
xnor U10002 (N_10002,N_9822,N_9802);
nand U10003 (N_10003,N_9882,N_9910);
and U10004 (N_10004,N_9966,N_9834);
or U10005 (N_10005,N_9988,N_9922);
nand U10006 (N_10006,N_9939,N_9844);
or U10007 (N_10007,N_9809,N_9815);
xor U10008 (N_10008,N_9888,N_9856);
xnor U10009 (N_10009,N_9977,N_9872);
or U10010 (N_10010,N_9804,N_9945);
and U10011 (N_10011,N_9836,N_9800);
xnor U10012 (N_10012,N_9840,N_9897);
or U10013 (N_10013,N_9969,N_9992);
xor U10014 (N_10014,N_9981,N_9807);
and U10015 (N_10015,N_9996,N_9983);
nor U10016 (N_10016,N_9857,N_9994);
or U10017 (N_10017,N_9816,N_9806);
nor U10018 (N_10018,N_9851,N_9980);
nor U10019 (N_10019,N_9876,N_9903);
xnor U10020 (N_10020,N_9932,N_9812);
nor U10021 (N_10021,N_9899,N_9948);
nand U10022 (N_10022,N_9978,N_9926);
and U10023 (N_10023,N_9920,N_9873);
or U10024 (N_10024,N_9864,N_9931);
or U10025 (N_10025,N_9825,N_9801);
and U10026 (N_10026,N_9867,N_9885);
nor U10027 (N_10027,N_9821,N_9918);
nand U10028 (N_10028,N_9805,N_9909);
or U10029 (N_10029,N_9865,N_9826);
nand U10030 (N_10030,N_9984,N_9934);
nand U10031 (N_10031,N_9896,N_9841);
nor U10032 (N_10032,N_9874,N_9892);
nor U10033 (N_10033,N_9820,N_9957);
or U10034 (N_10034,N_9839,N_9852);
and U10035 (N_10035,N_9927,N_9960);
nor U10036 (N_10036,N_9869,N_9877);
nor U10037 (N_10037,N_9814,N_9858);
or U10038 (N_10038,N_9997,N_9900);
or U10039 (N_10039,N_9937,N_9933);
nor U10040 (N_10040,N_9958,N_9972);
or U10041 (N_10041,N_9913,N_9880);
or U10042 (N_10042,N_9989,N_9915);
or U10043 (N_10043,N_9993,N_9944);
and U10044 (N_10044,N_9808,N_9975);
or U10045 (N_10045,N_9819,N_9887);
xor U10046 (N_10046,N_9886,N_9916);
nand U10047 (N_10047,N_9950,N_9965);
or U10048 (N_10048,N_9998,N_9908);
nor U10049 (N_10049,N_9924,N_9828);
and U10050 (N_10050,N_9879,N_9878);
xor U10051 (N_10051,N_9862,N_9875);
nand U10052 (N_10052,N_9853,N_9985);
xnor U10053 (N_10053,N_9827,N_9818);
or U10054 (N_10054,N_9940,N_9835);
nand U10055 (N_10055,N_9871,N_9838);
nand U10056 (N_10056,N_9912,N_9914);
nand U10057 (N_10057,N_9923,N_9847);
xnor U10058 (N_10058,N_9905,N_9894);
and U10059 (N_10059,N_9982,N_9991);
xor U10060 (N_10060,N_9863,N_9898);
nand U10061 (N_10061,N_9995,N_9971);
xor U10062 (N_10062,N_9895,N_9938);
nor U10063 (N_10063,N_9831,N_9999);
xnor U10064 (N_10064,N_9837,N_9963);
and U10065 (N_10065,N_9866,N_9979);
nor U10066 (N_10066,N_9830,N_9850);
and U10067 (N_10067,N_9881,N_9976);
xor U10068 (N_10068,N_9889,N_9870);
nand U10069 (N_10069,N_9942,N_9928);
xor U10070 (N_10070,N_9906,N_9947);
nor U10071 (N_10071,N_9861,N_9832);
nor U10072 (N_10072,N_9955,N_9854);
xnor U10073 (N_10073,N_9890,N_9848);
nand U10074 (N_10074,N_9962,N_9954);
and U10075 (N_10075,N_9811,N_9845);
nand U10076 (N_10076,N_9986,N_9902);
xor U10077 (N_10077,N_9833,N_9846);
and U10078 (N_10078,N_9813,N_9868);
nor U10079 (N_10079,N_9946,N_9959);
xor U10080 (N_10080,N_9964,N_9911);
xnor U10081 (N_10081,N_9901,N_9973);
or U10082 (N_10082,N_9990,N_9970);
nand U10083 (N_10083,N_9904,N_9968);
and U10084 (N_10084,N_9824,N_9951);
nor U10085 (N_10085,N_9967,N_9935);
or U10086 (N_10086,N_9943,N_9803);
and U10087 (N_10087,N_9883,N_9843);
or U10088 (N_10088,N_9842,N_9941);
nor U10089 (N_10089,N_9823,N_9859);
xnor U10090 (N_10090,N_9917,N_9921);
nor U10091 (N_10091,N_9891,N_9855);
xor U10092 (N_10092,N_9860,N_9953);
nand U10093 (N_10093,N_9974,N_9849);
nand U10094 (N_10094,N_9930,N_9949);
and U10095 (N_10095,N_9810,N_9907);
and U10096 (N_10096,N_9893,N_9925);
nand U10097 (N_10097,N_9987,N_9829);
xnor U10098 (N_10098,N_9961,N_9952);
and U10099 (N_10099,N_9919,N_9929);
and U10100 (N_10100,N_9868,N_9870);
nand U10101 (N_10101,N_9873,N_9956);
and U10102 (N_10102,N_9827,N_9955);
nor U10103 (N_10103,N_9848,N_9993);
or U10104 (N_10104,N_9987,N_9900);
and U10105 (N_10105,N_9888,N_9815);
xor U10106 (N_10106,N_9949,N_9919);
nor U10107 (N_10107,N_9909,N_9884);
or U10108 (N_10108,N_9803,N_9835);
or U10109 (N_10109,N_9973,N_9801);
or U10110 (N_10110,N_9831,N_9929);
or U10111 (N_10111,N_9869,N_9984);
xor U10112 (N_10112,N_9856,N_9867);
nand U10113 (N_10113,N_9853,N_9803);
and U10114 (N_10114,N_9968,N_9928);
and U10115 (N_10115,N_9861,N_9949);
and U10116 (N_10116,N_9852,N_9806);
nor U10117 (N_10117,N_9915,N_9801);
nand U10118 (N_10118,N_9800,N_9941);
nand U10119 (N_10119,N_9926,N_9891);
nand U10120 (N_10120,N_9891,N_9917);
or U10121 (N_10121,N_9887,N_9831);
nand U10122 (N_10122,N_9975,N_9898);
or U10123 (N_10123,N_9910,N_9934);
nand U10124 (N_10124,N_9806,N_9937);
and U10125 (N_10125,N_9988,N_9834);
xnor U10126 (N_10126,N_9941,N_9819);
and U10127 (N_10127,N_9898,N_9944);
nand U10128 (N_10128,N_9934,N_9995);
or U10129 (N_10129,N_9894,N_9995);
nor U10130 (N_10130,N_9947,N_9920);
nor U10131 (N_10131,N_9801,N_9928);
and U10132 (N_10132,N_9828,N_9857);
and U10133 (N_10133,N_9858,N_9889);
nor U10134 (N_10134,N_9995,N_9979);
and U10135 (N_10135,N_9931,N_9930);
nand U10136 (N_10136,N_9870,N_9856);
nand U10137 (N_10137,N_9970,N_9846);
nor U10138 (N_10138,N_9814,N_9989);
nor U10139 (N_10139,N_9876,N_9961);
or U10140 (N_10140,N_9835,N_9897);
or U10141 (N_10141,N_9835,N_9933);
nand U10142 (N_10142,N_9815,N_9918);
or U10143 (N_10143,N_9871,N_9945);
nor U10144 (N_10144,N_9973,N_9996);
xor U10145 (N_10145,N_9895,N_9805);
xnor U10146 (N_10146,N_9831,N_9898);
nor U10147 (N_10147,N_9928,N_9966);
xnor U10148 (N_10148,N_9852,N_9904);
xor U10149 (N_10149,N_9912,N_9942);
and U10150 (N_10150,N_9804,N_9991);
xor U10151 (N_10151,N_9841,N_9811);
and U10152 (N_10152,N_9998,N_9835);
nor U10153 (N_10153,N_9990,N_9992);
or U10154 (N_10154,N_9802,N_9886);
nand U10155 (N_10155,N_9914,N_9813);
xnor U10156 (N_10156,N_9820,N_9831);
xnor U10157 (N_10157,N_9834,N_9912);
or U10158 (N_10158,N_9943,N_9883);
and U10159 (N_10159,N_9951,N_9853);
nor U10160 (N_10160,N_9890,N_9926);
and U10161 (N_10161,N_9871,N_9864);
or U10162 (N_10162,N_9931,N_9810);
nand U10163 (N_10163,N_9995,N_9928);
nor U10164 (N_10164,N_9869,N_9912);
or U10165 (N_10165,N_9880,N_9829);
xnor U10166 (N_10166,N_9876,N_9865);
or U10167 (N_10167,N_9983,N_9951);
or U10168 (N_10168,N_9808,N_9885);
and U10169 (N_10169,N_9845,N_9838);
or U10170 (N_10170,N_9987,N_9816);
or U10171 (N_10171,N_9831,N_9859);
and U10172 (N_10172,N_9887,N_9931);
nor U10173 (N_10173,N_9871,N_9860);
nand U10174 (N_10174,N_9903,N_9821);
nor U10175 (N_10175,N_9912,N_9882);
nor U10176 (N_10176,N_9944,N_9901);
nor U10177 (N_10177,N_9897,N_9868);
xnor U10178 (N_10178,N_9913,N_9888);
nor U10179 (N_10179,N_9920,N_9828);
nand U10180 (N_10180,N_9827,N_9829);
xnor U10181 (N_10181,N_9999,N_9914);
nand U10182 (N_10182,N_9949,N_9859);
nor U10183 (N_10183,N_9953,N_9986);
xnor U10184 (N_10184,N_9800,N_9823);
xor U10185 (N_10185,N_9853,N_9807);
or U10186 (N_10186,N_9933,N_9913);
or U10187 (N_10187,N_9896,N_9879);
and U10188 (N_10188,N_9845,N_9824);
or U10189 (N_10189,N_9892,N_9817);
and U10190 (N_10190,N_9987,N_9982);
nor U10191 (N_10191,N_9964,N_9843);
nor U10192 (N_10192,N_9824,N_9809);
or U10193 (N_10193,N_9846,N_9883);
and U10194 (N_10194,N_9966,N_9903);
or U10195 (N_10195,N_9883,N_9997);
and U10196 (N_10196,N_9995,N_9942);
nand U10197 (N_10197,N_9937,N_9889);
or U10198 (N_10198,N_9896,N_9823);
or U10199 (N_10199,N_9820,N_9823);
nand U10200 (N_10200,N_10106,N_10138);
xnor U10201 (N_10201,N_10030,N_10097);
nor U10202 (N_10202,N_10153,N_10051);
nor U10203 (N_10203,N_10099,N_10107);
and U10204 (N_10204,N_10175,N_10019);
and U10205 (N_10205,N_10032,N_10071);
and U10206 (N_10206,N_10193,N_10196);
or U10207 (N_10207,N_10133,N_10011);
xor U10208 (N_10208,N_10180,N_10144);
nand U10209 (N_10209,N_10105,N_10112);
xnor U10210 (N_10210,N_10125,N_10183);
xor U10211 (N_10211,N_10123,N_10058);
nor U10212 (N_10212,N_10146,N_10100);
and U10213 (N_10213,N_10091,N_10087);
nand U10214 (N_10214,N_10132,N_10151);
and U10215 (N_10215,N_10002,N_10092);
nor U10216 (N_10216,N_10197,N_10088);
or U10217 (N_10217,N_10159,N_10041);
and U10218 (N_10218,N_10048,N_10082);
nor U10219 (N_10219,N_10047,N_10073);
xnor U10220 (N_10220,N_10184,N_10093);
and U10221 (N_10221,N_10065,N_10074);
nand U10222 (N_10222,N_10124,N_10182);
nand U10223 (N_10223,N_10186,N_10016);
or U10224 (N_10224,N_10079,N_10101);
and U10225 (N_10225,N_10166,N_10078);
xnor U10226 (N_10226,N_10006,N_10070);
or U10227 (N_10227,N_10143,N_10160);
nor U10228 (N_10228,N_10198,N_10140);
and U10229 (N_10229,N_10167,N_10035);
nor U10230 (N_10230,N_10054,N_10008);
nand U10231 (N_10231,N_10042,N_10031);
nand U10232 (N_10232,N_10033,N_10017);
and U10233 (N_10233,N_10121,N_10076);
nand U10234 (N_10234,N_10057,N_10090);
and U10235 (N_10235,N_10053,N_10150);
and U10236 (N_10236,N_10178,N_10174);
and U10237 (N_10237,N_10045,N_10118);
nor U10238 (N_10238,N_10157,N_10148);
nor U10239 (N_10239,N_10120,N_10134);
or U10240 (N_10240,N_10027,N_10015);
xnor U10241 (N_10241,N_10116,N_10012);
xnor U10242 (N_10242,N_10155,N_10114);
nand U10243 (N_10243,N_10024,N_10023);
nor U10244 (N_10244,N_10001,N_10007);
nand U10245 (N_10245,N_10104,N_10152);
or U10246 (N_10246,N_10108,N_10034);
xor U10247 (N_10247,N_10004,N_10113);
and U10248 (N_10248,N_10028,N_10068);
or U10249 (N_10249,N_10172,N_10064);
nand U10250 (N_10250,N_10095,N_10036);
or U10251 (N_10251,N_10063,N_10158);
xnor U10252 (N_10252,N_10188,N_10136);
nand U10253 (N_10253,N_10111,N_10029);
nand U10254 (N_10254,N_10145,N_10110);
and U10255 (N_10255,N_10096,N_10083);
nor U10256 (N_10256,N_10161,N_10168);
nand U10257 (N_10257,N_10130,N_10185);
or U10258 (N_10258,N_10043,N_10052);
nand U10259 (N_10259,N_10163,N_10069);
nor U10260 (N_10260,N_10187,N_10009);
nand U10261 (N_10261,N_10094,N_10194);
xor U10262 (N_10262,N_10044,N_10179);
or U10263 (N_10263,N_10060,N_10010);
xor U10264 (N_10264,N_10037,N_10171);
nor U10265 (N_10265,N_10086,N_10142);
nor U10266 (N_10266,N_10137,N_10177);
and U10267 (N_10267,N_10089,N_10169);
xnor U10268 (N_10268,N_10170,N_10109);
nor U10269 (N_10269,N_10055,N_10005);
and U10270 (N_10270,N_10039,N_10000);
and U10271 (N_10271,N_10013,N_10128);
xnor U10272 (N_10272,N_10066,N_10129);
and U10273 (N_10273,N_10061,N_10080);
xnor U10274 (N_10274,N_10067,N_10103);
or U10275 (N_10275,N_10156,N_10003);
nand U10276 (N_10276,N_10122,N_10119);
nor U10277 (N_10277,N_10020,N_10059);
nor U10278 (N_10278,N_10077,N_10126);
or U10279 (N_10279,N_10040,N_10115);
xnor U10280 (N_10280,N_10056,N_10139);
nand U10281 (N_10281,N_10050,N_10149);
nor U10282 (N_10282,N_10199,N_10038);
xor U10283 (N_10283,N_10189,N_10195);
xor U10284 (N_10284,N_10127,N_10173);
xnor U10285 (N_10285,N_10102,N_10154);
xor U10286 (N_10286,N_10191,N_10135);
nand U10287 (N_10287,N_10176,N_10085);
nor U10288 (N_10288,N_10046,N_10164);
nor U10289 (N_10289,N_10165,N_10192);
and U10290 (N_10290,N_10084,N_10162);
nand U10291 (N_10291,N_10181,N_10018);
nor U10292 (N_10292,N_10131,N_10075);
nor U10293 (N_10293,N_10026,N_10049);
nand U10294 (N_10294,N_10025,N_10021);
nor U10295 (N_10295,N_10141,N_10062);
or U10296 (N_10296,N_10014,N_10190);
xnor U10297 (N_10297,N_10147,N_10117);
xnor U10298 (N_10298,N_10072,N_10022);
nand U10299 (N_10299,N_10098,N_10081);
nor U10300 (N_10300,N_10055,N_10148);
nor U10301 (N_10301,N_10175,N_10060);
xor U10302 (N_10302,N_10059,N_10022);
nand U10303 (N_10303,N_10052,N_10075);
nand U10304 (N_10304,N_10058,N_10076);
xor U10305 (N_10305,N_10080,N_10190);
xor U10306 (N_10306,N_10031,N_10091);
nor U10307 (N_10307,N_10141,N_10030);
or U10308 (N_10308,N_10143,N_10159);
and U10309 (N_10309,N_10074,N_10022);
xnor U10310 (N_10310,N_10123,N_10012);
xnor U10311 (N_10311,N_10089,N_10115);
nand U10312 (N_10312,N_10174,N_10092);
nor U10313 (N_10313,N_10081,N_10009);
nor U10314 (N_10314,N_10154,N_10168);
xor U10315 (N_10315,N_10004,N_10062);
xnor U10316 (N_10316,N_10068,N_10192);
and U10317 (N_10317,N_10198,N_10155);
or U10318 (N_10318,N_10147,N_10042);
or U10319 (N_10319,N_10120,N_10067);
nand U10320 (N_10320,N_10179,N_10159);
and U10321 (N_10321,N_10002,N_10062);
nand U10322 (N_10322,N_10198,N_10080);
and U10323 (N_10323,N_10188,N_10177);
or U10324 (N_10324,N_10019,N_10054);
and U10325 (N_10325,N_10171,N_10007);
xnor U10326 (N_10326,N_10020,N_10097);
xor U10327 (N_10327,N_10147,N_10078);
and U10328 (N_10328,N_10035,N_10145);
nor U10329 (N_10329,N_10153,N_10162);
nor U10330 (N_10330,N_10169,N_10110);
nand U10331 (N_10331,N_10154,N_10042);
xor U10332 (N_10332,N_10113,N_10077);
nand U10333 (N_10333,N_10189,N_10006);
and U10334 (N_10334,N_10093,N_10032);
nand U10335 (N_10335,N_10031,N_10073);
xor U10336 (N_10336,N_10018,N_10092);
and U10337 (N_10337,N_10083,N_10102);
nor U10338 (N_10338,N_10159,N_10038);
and U10339 (N_10339,N_10189,N_10124);
nand U10340 (N_10340,N_10106,N_10051);
xnor U10341 (N_10341,N_10068,N_10089);
nand U10342 (N_10342,N_10007,N_10184);
and U10343 (N_10343,N_10106,N_10025);
xnor U10344 (N_10344,N_10157,N_10161);
nor U10345 (N_10345,N_10189,N_10178);
nor U10346 (N_10346,N_10007,N_10193);
or U10347 (N_10347,N_10068,N_10178);
and U10348 (N_10348,N_10121,N_10101);
nor U10349 (N_10349,N_10138,N_10186);
or U10350 (N_10350,N_10192,N_10186);
nand U10351 (N_10351,N_10174,N_10113);
xnor U10352 (N_10352,N_10020,N_10130);
nand U10353 (N_10353,N_10026,N_10100);
nand U10354 (N_10354,N_10048,N_10016);
or U10355 (N_10355,N_10107,N_10193);
nand U10356 (N_10356,N_10178,N_10054);
xor U10357 (N_10357,N_10032,N_10067);
nor U10358 (N_10358,N_10016,N_10131);
and U10359 (N_10359,N_10053,N_10151);
and U10360 (N_10360,N_10105,N_10029);
or U10361 (N_10361,N_10082,N_10123);
nor U10362 (N_10362,N_10053,N_10132);
or U10363 (N_10363,N_10107,N_10050);
nor U10364 (N_10364,N_10134,N_10111);
xor U10365 (N_10365,N_10102,N_10129);
xnor U10366 (N_10366,N_10076,N_10054);
nor U10367 (N_10367,N_10005,N_10161);
nand U10368 (N_10368,N_10029,N_10025);
nand U10369 (N_10369,N_10010,N_10083);
xor U10370 (N_10370,N_10175,N_10168);
nand U10371 (N_10371,N_10003,N_10017);
xor U10372 (N_10372,N_10110,N_10134);
nor U10373 (N_10373,N_10128,N_10165);
and U10374 (N_10374,N_10011,N_10058);
xnor U10375 (N_10375,N_10196,N_10153);
nand U10376 (N_10376,N_10091,N_10118);
and U10377 (N_10377,N_10094,N_10130);
xor U10378 (N_10378,N_10185,N_10019);
or U10379 (N_10379,N_10156,N_10172);
nor U10380 (N_10380,N_10177,N_10042);
nor U10381 (N_10381,N_10007,N_10046);
xnor U10382 (N_10382,N_10197,N_10022);
xor U10383 (N_10383,N_10105,N_10030);
nand U10384 (N_10384,N_10130,N_10157);
nand U10385 (N_10385,N_10081,N_10148);
nor U10386 (N_10386,N_10006,N_10159);
xnor U10387 (N_10387,N_10104,N_10051);
nand U10388 (N_10388,N_10132,N_10010);
nand U10389 (N_10389,N_10157,N_10018);
or U10390 (N_10390,N_10121,N_10136);
nor U10391 (N_10391,N_10195,N_10021);
nor U10392 (N_10392,N_10052,N_10166);
xnor U10393 (N_10393,N_10140,N_10094);
xnor U10394 (N_10394,N_10025,N_10093);
and U10395 (N_10395,N_10117,N_10052);
nor U10396 (N_10396,N_10149,N_10094);
nor U10397 (N_10397,N_10001,N_10126);
nand U10398 (N_10398,N_10085,N_10139);
or U10399 (N_10399,N_10119,N_10129);
xnor U10400 (N_10400,N_10254,N_10317);
and U10401 (N_10401,N_10353,N_10358);
nor U10402 (N_10402,N_10334,N_10219);
nand U10403 (N_10403,N_10283,N_10379);
xnor U10404 (N_10404,N_10271,N_10206);
nand U10405 (N_10405,N_10314,N_10276);
or U10406 (N_10406,N_10269,N_10383);
nor U10407 (N_10407,N_10278,N_10273);
and U10408 (N_10408,N_10214,N_10374);
nor U10409 (N_10409,N_10369,N_10343);
or U10410 (N_10410,N_10253,N_10258);
nand U10411 (N_10411,N_10251,N_10325);
xnor U10412 (N_10412,N_10396,N_10244);
or U10413 (N_10413,N_10381,N_10368);
nand U10414 (N_10414,N_10255,N_10393);
nand U10415 (N_10415,N_10313,N_10264);
and U10416 (N_10416,N_10384,N_10280);
or U10417 (N_10417,N_10351,N_10227);
and U10418 (N_10418,N_10247,N_10289);
and U10419 (N_10419,N_10236,N_10388);
and U10420 (N_10420,N_10245,N_10259);
or U10421 (N_10421,N_10286,N_10232);
xnor U10422 (N_10422,N_10208,N_10315);
nor U10423 (N_10423,N_10225,N_10222);
and U10424 (N_10424,N_10332,N_10377);
or U10425 (N_10425,N_10287,N_10346);
nor U10426 (N_10426,N_10339,N_10274);
or U10427 (N_10427,N_10284,N_10341);
or U10428 (N_10428,N_10223,N_10272);
and U10429 (N_10429,N_10306,N_10285);
nor U10430 (N_10430,N_10263,N_10275);
xor U10431 (N_10431,N_10361,N_10266);
nor U10432 (N_10432,N_10270,N_10290);
nor U10433 (N_10433,N_10249,N_10331);
xnor U10434 (N_10434,N_10328,N_10333);
or U10435 (N_10435,N_10395,N_10371);
nand U10436 (N_10436,N_10324,N_10362);
nand U10437 (N_10437,N_10342,N_10252);
nand U10438 (N_10438,N_10399,N_10200);
and U10439 (N_10439,N_10262,N_10323);
and U10440 (N_10440,N_10336,N_10391);
nor U10441 (N_10441,N_10352,N_10218);
or U10442 (N_10442,N_10392,N_10387);
xor U10443 (N_10443,N_10326,N_10318);
or U10444 (N_10444,N_10228,N_10316);
and U10445 (N_10445,N_10338,N_10213);
nand U10446 (N_10446,N_10205,N_10356);
and U10447 (N_10447,N_10217,N_10216);
nand U10448 (N_10448,N_10229,N_10327);
or U10449 (N_10449,N_10364,N_10312);
nor U10450 (N_10450,N_10321,N_10345);
or U10451 (N_10451,N_10367,N_10221);
or U10452 (N_10452,N_10375,N_10237);
or U10453 (N_10453,N_10241,N_10299);
xnor U10454 (N_10454,N_10308,N_10347);
or U10455 (N_10455,N_10360,N_10305);
and U10456 (N_10456,N_10242,N_10261);
nand U10457 (N_10457,N_10335,N_10319);
or U10458 (N_10458,N_10320,N_10382);
and U10459 (N_10459,N_10322,N_10296);
nand U10460 (N_10460,N_10386,N_10380);
nor U10461 (N_10461,N_10240,N_10350);
xor U10462 (N_10462,N_10376,N_10366);
and U10463 (N_10463,N_10355,N_10281);
or U10464 (N_10464,N_10354,N_10265);
nand U10465 (N_10465,N_10268,N_10256);
nor U10466 (N_10466,N_10370,N_10344);
or U10467 (N_10467,N_10202,N_10233);
nor U10468 (N_10468,N_10311,N_10349);
and U10469 (N_10469,N_10300,N_10304);
nand U10470 (N_10470,N_10298,N_10210);
nand U10471 (N_10471,N_10243,N_10373);
nand U10472 (N_10472,N_10389,N_10291);
nand U10473 (N_10473,N_10359,N_10250);
xnor U10474 (N_10474,N_10288,N_10365);
nor U10475 (N_10475,N_10385,N_10230);
xor U10476 (N_10476,N_10310,N_10397);
xor U10477 (N_10477,N_10294,N_10260);
nand U10478 (N_10478,N_10394,N_10248);
and U10479 (N_10479,N_10212,N_10372);
nand U10480 (N_10480,N_10220,N_10282);
nor U10481 (N_10481,N_10215,N_10203);
nand U10482 (N_10482,N_10309,N_10257);
xor U10483 (N_10483,N_10267,N_10302);
or U10484 (N_10484,N_10201,N_10297);
nand U10485 (N_10485,N_10224,N_10292);
xnor U10486 (N_10486,N_10301,N_10293);
or U10487 (N_10487,N_10378,N_10303);
nand U10488 (N_10488,N_10329,N_10279);
nor U10489 (N_10489,N_10277,N_10330);
xnor U10490 (N_10490,N_10239,N_10307);
or U10491 (N_10491,N_10209,N_10238);
xor U10492 (N_10492,N_10207,N_10235);
nand U10493 (N_10493,N_10295,N_10398);
and U10494 (N_10494,N_10211,N_10204);
and U10495 (N_10495,N_10340,N_10337);
nor U10496 (N_10496,N_10231,N_10390);
xor U10497 (N_10497,N_10226,N_10246);
and U10498 (N_10498,N_10363,N_10234);
nor U10499 (N_10499,N_10348,N_10357);
nor U10500 (N_10500,N_10356,N_10325);
nand U10501 (N_10501,N_10368,N_10209);
and U10502 (N_10502,N_10362,N_10348);
or U10503 (N_10503,N_10268,N_10217);
or U10504 (N_10504,N_10207,N_10352);
and U10505 (N_10505,N_10238,N_10273);
nor U10506 (N_10506,N_10396,N_10274);
nor U10507 (N_10507,N_10203,N_10314);
nand U10508 (N_10508,N_10202,N_10240);
or U10509 (N_10509,N_10272,N_10255);
xor U10510 (N_10510,N_10312,N_10346);
nand U10511 (N_10511,N_10275,N_10298);
and U10512 (N_10512,N_10242,N_10296);
and U10513 (N_10513,N_10321,N_10272);
xnor U10514 (N_10514,N_10327,N_10247);
nand U10515 (N_10515,N_10354,N_10391);
and U10516 (N_10516,N_10270,N_10354);
xnor U10517 (N_10517,N_10256,N_10331);
xor U10518 (N_10518,N_10220,N_10264);
nand U10519 (N_10519,N_10399,N_10251);
nor U10520 (N_10520,N_10253,N_10236);
nor U10521 (N_10521,N_10248,N_10371);
and U10522 (N_10522,N_10373,N_10376);
nor U10523 (N_10523,N_10322,N_10207);
or U10524 (N_10524,N_10304,N_10355);
or U10525 (N_10525,N_10270,N_10304);
xnor U10526 (N_10526,N_10279,N_10267);
and U10527 (N_10527,N_10260,N_10358);
nand U10528 (N_10528,N_10341,N_10387);
xnor U10529 (N_10529,N_10374,N_10239);
nand U10530 (N_10530,N_10222,N_10285);
xor U10531 (N_10531,N_10316,N_10298);
nand U10532 (N_10532,N_10309,N_10288);
nor U10533 (N_10533,N_10248,N_10221);
xnor U10534 (N_10534,N_10320,N_10296);
nand U10535 (N_10535,N_10280,N_10292);
nand U10536 (N_10536,N_10315,N_10231);
and U10537 (N_10537,N_10226,N_10372);
or U10538 (N_10538,N_10261,N_10217);
or U10539 (N_10539,N_10201,N_10387);
xor U10540 (N_10540,N_10263,N_10265);
or U10541 (N_10541,N_10228,N_10253);
xnor U10542 (N_10542,N_10225,N_10211);
and U10543 (N_10543,N_10217,N_10275);
and U10544 (N_10544,N_10387,N_10204);
nand U10545 (N_10545,N_10327,N_10368);
nand U10546 (N_10546,N_10250,N_10388);
nor U10547 (N_10547,N_10374,N_10246);
xnor U10548 (N_10548,N_10287,N_10336);
nor U10549 (N_10549,N_10330,N_10309);
nor U10550 (N_10550,N_10336,N_10372);
nand U10551 (N_10551,N_10265,N_10345);
and U10552 (N_10552,N_10286,N_10304);
xor U10553 (N_10553,N_10205,N_10290);
nor U10554 (N_10554,N_10318,N_10391);
xnor U10555 (N_10555,N_10325,N_10205);
nor U10556 (N_10556,N_10333,N_10269);
and U10557 (N_10557,N_10376,N_10226);
xnor U10558 (N_10558,N_10227,N_10361);
and U10559 (N_10559,N_10215,N_10370);
xnor U10560 (N_10560,N_10353,N_10381);
or U10561 (N_10561,N_10360,N_10276);
nor U10562 (N_10562,N_10339,N_10348);
nand U10563 (N_10563,N_10349,N_10339);
and U10564 (N_10564,N_10207,N_10371);
nand U10565 (N_10565,N_10383,N_10263);
nand U10566 (N_10566,N_10240,N_10290);
nor U10567 (N_10567,N_10342,N_10249);
nor U10568 (N_10568,N_10282,N_10266);
nand U10569 (N_10569,N_10250,N_10317);
and U10570 (N_10570,N_10278,N_10286);
xnor U10571 (N_10571,N_10289,N_10389);
nor U10572 (N_10572,N_10364,N_10253);
and U10573 (N_10573,N_10328,N_10336);
nor U10574 (N_10574,N_10295,N_10397);
or U10575 (N_10575,N_10277,N_10318);
nor U10576 (N_10576,N_10342,N_10333);
xnor U10577 (N_10577,N_10200,N_10353);
and U10578 (N_10578,N_10346,N_10358);
and U10579 (N_10579,N_10374,N_10224);
nor U10580 (N_10580,N_10244,N_10231);
xnor U10581 (N_10581,N_10240,N_10221);
xnor U10582 (N_10582,N_10313,N_10217);
or U10583 (N_10583,N_10289,N_10296);
nor U10584 (N_10584,N_10291,N_10276);
and U10585 (N_10585,N_10225,N_10292);
nand U10586 (N_10586,N_10279,N_10367);
nor U10587 (N_10587,N_10256,N_10287);
xnor U10588 (N_10588,N_10285,N_10234);
or U10589 (N_10589,N_10271,N_10245);
nand U10590 (N_10590,N_10392,N_10279);
and U10591 (N_10591,N_10259,N_10252);
or U10592 (N_10592,N_10323,N_10368);
nand U10593 (N_10593,N_10290,N_10215);
nand U10594 (N_10594,N_10279,N_10250);
and U10595 (N_10595,N_10358,N_10271);
nor U10596 (N_10596,N_10308,N_10245);
and U10597 (N_10597,N_10218,N_10221);
nand U10598 (N_10598,N_10268,N_10397);
and U10599 (N_10599,N_10212,N_10231);
xnor U10600 (N_10600,N_10462,N_10542);
nor U10601 (N_10601,N_10553,N_10550);
nor U10602 (N_10602,N_10571,N_10419);
nand U10603 (N_10603,N_10416,N_10405);
or U10604 (N_10604,N_10483,N_10522);
and U10605 (N_10605,N_10516,N_10530);
nor U10606 (N_10606,N_10453,N_10544);
nor U10607 (N_10607,N_10408,N_10525);
nor U10608 (N_10608,N_10572,N_10503);
nand U10609 (N_10609,N_10493,N_10579);
or U10610 (N_10610,N_10593,N_10440);
nand U10611 (N_10611,N_10499,N_10509);
or U10612 (N_10612,N_10528,N_10433);
or U10613 (N_10613,N_10429,N_10497);
nor U10614 (N_10614,N_10545,N_10476);
and U10615 (N_10615,N_10486,N_10535);
nand U10616 (N_10616,N_10576,N_10401);
xor U10617 (N_10617,N_10599,N_10537);
nand U10618 (N_10618,N_10425,N_10541);
nand U10619 (N_10619,N_10507,N_10482);
nand U10620 (N_10620,N_10573,N_10506);
or U10621 (N_10621,N_10466,N_10539);
nand U10622 (N_10622,N_10442,N_10524);
or U10623 (N_10623,N_10508,N_10454);
nand U10624 (N_10624,N_10591,N_10452);
nand U10625 (N_10625,N_10560,N_10410);
and U10626 (N_10626,N_10496,N_10479);
xor U10627 (N_10627,N_10534,N_10489);
xor U10628 (N_10628,N_10494,N_10501);
nor U10629 (N_10629,N_10472,N_10490);
xnor U10630 (N_10630,N_10404,N_10447);
or U10631 (N_10631,N_10465,N_10475);
and U10632 (N_10632,N_10592,N_10484);
or U10633 (N_10633,N_10443,N_10538);
or U10634 (N_10634,N_10449,N_10402);
and U10635 (N_10635,N_10575,N_10540);
nor U10636 (N_10636,N_10510,N_10546);
and U10637 (N_10637,N_10406,N_10557);
or U10638 (N_10638,N_10585,N_10526);
and U10639 (N_10639,N_10423,N_10445);
nor U10640 (N_10640,N_10444,N_10485);
xnor U10641 (N_10641,N_10529,N_10428);
or U10642 (N_10642,N_10418,N_10468);
nor U10643 (N_10643,N_10595,N_10407);
xnor U10644 (N_10644,N_10531,N_10457);
nand U10645 (N_10645,N_10562,N_10597);
and U10646 (N_10646,N_10439,N_10561);
nand U10647 (N_10647,N_10467,N_10463);
nand U10648 (N_10648,N_10556,N_10582);
nand U10649 (N_10649,N_10421,N_10515);
or U10650 (N_10650,N_10450,N_10456);
nor U10651 (N_10651,N_10536,N_10504);
or U10652 (N_10652,N_10413,N_10533);
or U10653 (N_10653,N_10578,N_10474);
and U10654 (N_10654,N_10424,N_10491);
nand U10655 (N_10655,N_10412,N_10566);
nand U10656 (N_10656,N_10437,N_10565);
or U10657 (N_10657,N_10511,N_10470);
or U10658 (N_10658,N_10517,N_10594);
nand U10659 (N_10659,N_10559,N_10568);
or U10660 (N_10660,N_10555,N_10487);
xor U10661 (N_10661,N_10518,N_10481);
xor U10662 (N_10662,N_10581,N_10589);
or U10663 (N_10663,N_10492,N_10434);
nand U10664 (N_10664,N_10549,N_10498);
nand U10665 (N_10665,N_10558,N_10458);
nor U10666 (N_10666,N_10430,N_10426);
and U10667 (N_10667,N_10502,N_10469);
nor U10668 (N_10668,N_10514,N_10415);
xor U10669 (N_10669,N_10422,N_10473);
and U10670 (N_10670,N_10598,N_10435);
xor U10671 (N_10671,N_10587,N_10495);
xor U10672 (N_10672,N_10431,N_10563);
and U10673 (N_10673,N_10551,N_10455);
nor U10674 (N_10674,N_10417,N_10584);
and U10675 (N_10675,N_10480,N_10432);
xor U10676 (N_10676,N_10436,N_10420);
nor U10677 (N_10677,N_10580,N_10570);
nor U10678 (N_10678,N_10567,N_10527);
nand U10679 (N_10679,N_10446,N_10577);
nand U10680 (N_10680,N_10464,N_10548);
xor U10681 (N_10681,N_10403,N_10532);
xor U10682 (N_10682,N_10586,N_10441);
nand U10683 (N_10683,N_10523,N_10513);
and U10684 (N_10684,N_10554,N_10569);
nand U10685 (N_10685,N_10519,N_10414);
and U10686 (N_10686,N_10583,N_10438);
nor U10687 (N_10687,N_10448,N_10459);
nor U10688 (N_10688,N_10505,N_10477);
nor U10689 (N_10689,N_10488,N_10409);
and U10690 (N_10690,N_10512,N_10588);
nand U10691 (N_10691,N_10547,N_10552);
nand U10692 (N_10692,N_10500,N_10411);
and U10693 (N_10693,N_10478,N_10427);
xnor U10694 (N_10694,N_10400,N_10590);
nor U10695 (N_10695,N_10471,N_10521);
xnor U10696 (N_10696,N_10460,N_10520);
or U10697 (N_10697,N_10564,N_10461);
and U10698 (N_10698,N_10543,N_10596);
nor U10699 (N_10699,N_10574,N_10451);
nand U10700 (N_10700,N_10486,N_10595);
or U10701 (N_10701,N_10475,N_10535);
nor U10702 (N_10702,N_10568,N_10490);
and U10703 (N_10703,N_10406,N_10478);
nand U10704 (N_10704,N_10593,N_10532);
nor U10705 (N_10705,N_10439,N_10564);
or U10706 (N_10706,N_10408,N_10449);
nor U10707 (N_10707,N_10576,N_10415);
xnor U10708 (N_10708,N_10402,N_10409);
nand U10709 (N_10709,N_10404,N_10598);
nand U10710 (N_10710,N_10512,N_10576);
xor U10711 (N_10711,N_10495,N_10481);
xor U10712 (N_10712,N_10488,N_10565);
nand U10713 (N_10713,N_10454,N_10589);
nor U10714 (N_10714,N_10497,N_10579);
and U10715 (N_10715,N_10427,N_10588);
nor U10716 (N_10716,N_10453,N_10589);
nor U10717 (N_10717,N_10443,N_10525);
and U10718 (N_10718,N_10485,N_10407);
xnor U10719 (N_10719,N_10445,N_10551);
nand U10720 (N_10720,N_10579,N_10403);
nand U10721 (N_10721,N_10407,N_10572);
xnor U10722 (N_10722,N_10412,N_10435);
nand U10723 (N_10723,N_10499,N_10478);
xnor U10724 (N_10724,N_10557,N_10499);
and U10725 (N_10725,N_10563,N_10438);
xnor U10726 (N_10726,N_10474,N_10555);
or U10727 (N_10727,N_10521,N_10460);
nand U10728 (N_10728,N_10520,N_10436);
or U10729 (N_10729,N_10487,N_10559);
nand U10730 (N_10730,N_10440,N_10570);
nand U10731 (N_10731,N_10580,N_10408);
or U10732 (N_10732,N_10542,N_10518);
nor U10733 (N_10733,N_10422,N_10456);
and U10734 (N_10734,N_10533,N_10565);
xnor U10735 (N_10735,N_10422,N_10538);
nor U10736 (N_10736,N_10549,N_10453);
and U10737 (N_10737,N_10570,N_10523);
and U10738 (N_10738,N_10515,N_10488);
nand U10739 (N_10739,N_10581,N_10400);
or U10740 (N_10740,N_10513,N_10448);
nand U10741 (N_10741,N_10525,N_10564);
nor U10742 (N_10742,N_10457,N_10585);
xnor U10743 (N_10743,N_10445,N_10412);
xnor U10744 (N_10744,N_10527,N_10457);
nand U10745 (N_10745,N_10422,N_10441);
nand U10746 (N_10746,N_10553,N_10453);
nor U10747 (N_10747,N_10405,N_10534);
nand U10748 (N_10748,N_10445,N_10473);
nor U10749 (N_10749,N_10584,N_10596);
and U10750 (N_10750,N_10510,N_10446);
and U10751 (N_10751,N_10471,N_10522);
or U10752 (N_10752,N_10548,N_10578);
or U10753 (N_10753,N_10591,N_10553);
nand U10754 (N_10754,N_10402,N_10515);
xnor U10755 (N_10755,N_10587,N_10588);
and U10756 (N_10756,N_10401,N_10515);
nor U10757 (N_10757,N_10408,N_10412);
and U10758 (N_10758,N_10428,N_10594);
nand U10759 (N_10759,N_10434,N_10448);
nor U10760 (N_10760,N_10498,N_10519);
nor U10761 (N_10761,N_10525,N_10486);
nor U10762 (N_10762,N_10592,N_10479);
or U10763 (N_10763,N_10412,N_10578);
xor U10764 (N_10764,N_10401,N_10455);
xor U10765 (N_10765,N_10474,N_10564);
xnor U10766 (N_10766,N_10503,N_10412);
or U10767 (N_10767,N_10510,N_10545);
and U10768 (N_10768,N_10434,N_10596);
nand U10769 (N_10769,N_10444,N_10501);
nand U10770 (N_10770,N_10532,N_10475);
and U10771 (N_10771,N_10424,N_10506);
xor U10772 (N_10772,N_10423,N_10542);
or U10773 (N_10773,N_10440,N_10594);
and U10774 (N_10774,N_10425,N_10436);
and U10775 (N_10775,N_10530,N_10574);
nor U10776 (N_10776,N_10464,N_10401);
nand U10777 (N_10777,N_10452,N_10556);
or U10778 (N_10778,N_10552,N_10568);
and U10779 (N_10779,N_10429,N_10542);
nand U10780 (N_10780,N_10408,N_10532);
nor U10781 (N_10781,N_10484,N_10595);
xnor U10782 (N_10782,N_10480,N_10452);
nand U10783 (N_10783,N_10535,N_10561);
nand U10784 (N_10784,N_10520,N_10494);
nand U10785 (N_10785,N_10516,N_10599);
nor U10786 (N_10786,N_10474,N_10576);
nor U10787 (N_10787,N_10453,N_10480);
nor U10788 (N_10788,N_10571,N_10459);
and U10789 (N_10789,N_10498,N_10524);
nor U10790 (N_10790,N_10592,N_10527);
xnor U10791 (N_10791,N_10436,N_10493);
or U10792 (N_10792,N_10591,N_10408);
xnor U10793 (N_10793,N_10565,N_10478);
nor U10794 (N_10794,N_10403,N_10450);
nand U10795 (N_10795,N_10552,N_10482);
xor U10796 (N_10796,N_10508,N_10525);
nor U10797 (N_10797,N_10541,N_10585);
nand U10798 (N_10798,N_10590,N_10489);
or U10799 (N_10799,N_10525,N_10524);
xnor U10800 (N_10800,N_10649,N_10624);
nand U10801 (N_10801,N_10600,N_10724);
nor U10802 (N_10802,N_10616,N_10755);
xnor U10803 (N_10803,N_10753,N_10679);
nand U10804 (N_10804,N_10754,N_10794);
nand U10805 (N_10805,N_10634,N_10749);
xor U10806 (N_10806,N_10602,N_10774);
xnor U10807 (N_10807,N_10729,N_10718);
nand U10808 (N_10808,N_10787,N_10623);
xor U10809 (N_10809,N_10711,N_10727);
and U10810 (N_10810,N_10622,N_10780);
nand U10811 (N_10811,N_10702,N_10695);
and U10812 (N_10812,N_10756,N_10767);
nand U10813 (N_10813,N_10715,N_10658);
or U10814 (N_10814,N_10628,N_10725);
nand U10815 (N_10815,N_10763,N_10760);
and U10816 (N_10816,N_10748,N_10721);
xnor U10817 (N_10817,N_10783,N_10762);
nand U10818 (N_10818,N_10666,N_10693);
nand U10819 (N_10819,N_10664,N_10635);
or U10820 (N_10820,N_10647,N_10643);
nand U10821 (N_10821,N_10633,N_10740);
nand U10822 (N_10822,N_10793,N_10722);
nor U10823 (N_10823,N_10686,N_10796);
or U10824 (N_10824,N_10619,N_10687);
nor U10825 (N_10825,N_10683,N_10690);
or U10826 (N_10826,N_10707,N_10610);
nor U10827 (N_10827,N_10714,N_10732);
nand U10828 (N_10828,N_10627,N_10772);
xor U10829 (N_10829,N_10688,N_10663);
and U10830 (N_10830,N_10608,N_10752);
nand U10831 (N_10831,N_10637,N_10680);
and U10832 (N_10832,N_10682,N_10670);
nand U10833 (N_10833,N_10692,N_10632);
or U10834 (N_10834,N_10785,N_10697);
or U10835 (N_10835,N_10605,N_10646);
or U10836 (N_10836,N_10703,N_10795);
nand U10837 (N_10837,N_10782,N_10720);
or U10838 (N_10838,N_10651,N_10764);
nand U10839 (N_10839,N_10644,N_10652);
and U10840 (N_10840,N_10614,N_10773);
nor U10841 (N_10841,N_10639,N_10659);
nor U10842 (N_10842,N_10654,N_10613);
xor U10843 (N_10843,N_10775,N_10789);
xor U10844 (N_10844,N_10641,N_10734);
and U10845 (N_10845,N_10779,N_10751);
xnor U10846 (N_10846,N_10665,N_10750);
and U10847 (N_10847,N_10738,N_10629);
nand U10848 (N_10848,N_10784,N_10747);
xnor U10849 (N_10849,N_10788,N_10672);
nor U10850 (N_10850,N_10798,N_10620);
and U10851 (N_10851,N_10630,N_10735);
xor U10852 (N_10852,N_10769,N_10716);
nand U10853 (N_10853,N_10611,N_10661);
xnor U10854 (N_10854,N_10657,N_10737);
nand U10855 (N_10855,N_10625,N_10696);
nand U10856 (N_10856,N_10704,N_10705);
nand U10857 (N_10857,N_10662,N_10719);
xnor U10858 (N_10858,N_10694,N_10667);
or U10859 (N_10859,N_10621,N_10604);
nand U10860 (N_10860,N_10700,N_10733);
nor U10861 (N_10861,N_10673,N_10757);
xnor U10862 (N_10862,N_10765,N_10742);
and U10863 (N_10863,N_10656,N_10701);
nand U10864 (N_10864,N_10618,N_10636);
nor U10865 (N_10865,N_10678,N_10771);
xor U10866 (N_10866,N_10626,N_10792);
nor U10867 (N_10867,N_10745,N_10744);
and U10868 (N_10868,N_10730,N_10713);
xor U10869 (N_10869,N_10766,N_10759);
and U10870 (N_10870,N_10617,N_10778);
nor U10871 (N_10871,N_10660,N_10712);
nor U10872 (N_10872,N_10655,N_10736);
and U10873 (N_10873,N_10675,N_10741);
nor U10874 (N_10874,N_10676,N_10653);
and U10875 (N_10875,N_10677,N_10640);
nand U10876 (N_10876,N_10706,N_10797);
or U10877 (N_10877,N_10717,N_10786);
and U10878 (N_10878,N_10648,N_10761);
and U10879 (N_10879,N_10746,N_10726);
or U10880 (N_10880,N_10731,N_10743);
and U10881 (N_10881,N_10708,N_10645);
and U10882 (N_10882,N_10698,N_10638);
xnor U10883 (N_10883,N_10709,N_10607);
nand U10884 (N_10884,N_10781,N_10710);
and U10885 (N_10885,N_10681,N_10674);
or U10886 (N_10886,N_10671,N_10684);
and U10887 (N_10887,N_10631,N_10612);
and U10888 (N_10888,N_10650,N_10609);
or U10889 (N_10889,N_10728,N_10777);
and U10890 (N_10890,N_10758,N_10768);
nor U10891 (N_10891,N_10601,N_10791);
or U10892 (N_10892,N_10699,N_10799);
nand U10893 (N_10893,N_10606,N_10776);
nor U10894 (N_10894,N_10668,N_10615);
or U10895 (N_10895,N_10642,N_10739);
and U10896 (N_10896,N_10685,N_10790);
xnor U10897 (N_10897,N_10689,N_10691);
and U10898 (N_10898,N_10603,N_10669);
nand U10899 (N_10899,N_10723,N_10770);
nor U10900 (N_10900,N_10665,N_10676);
or U10901 (N_10901,N_10662,N_10725);
nand U10902 (N_10902,N_10620,N_10726);
nor U10903 (N_10903,N_10767,N_10718);
nor U10904 (N_10904,N_10777,N_10675);
xor U10905 (N_10905,N_10744,N_10656);
nand U10906 (N_10906,N_10688,N_10696);
xnor U10907 (N_10907,N_10703,N_10744);
and U10908 (N_10908,N_10757,N_10739);
nand U10909 (N_10909,N_10746,N_10797);
xor U10910 (N_10910,N_10652,N_10725);
or U10911 (N_10911,N_10788,N_10765);
xor U10912 (N_10912,N_10674,N_10718);
or U10913 (N_10913,N_10750,N_10673);
nor U10914 (N_10914,N_10674,N_10761);
nand U10915 (N_10915,N_10780,N_10702);
nand U10916 (N_10916,N_10622,N_10752);
and U10917 (N_10917,N_10691,N_10788);
nand U10918 (N_10918,N_10629,N_10796);
nor U10919 (N_10919,N_10778,N_10741);
xor U10920 (N_10920,N_10774,N_10603);
nor U10921 (N_10921,N_10603,N_10786);
or U10922 (N_10922,N_10704,N_10760);
nand U10923 (N_10923,N_10664,N_10750);
xor U10924 (N_10924,N_10758,N_10785);
or U10925 (N_10925,N_10600,N_10622);
and U10926 (N_10926,N_10620,N_10696);
nor U10927 (N_10927,N_10678,N_10769);
or U10928 (N_10928,N_10640,N_10758);
nand U10929 (N_10929,N_10613,N_10636);
xnor U10930 (N_10930,N_10726,N_10604);
nand U10931 (N_10931,N_10737,N_10668);
nor U10932 (N_10932,N_10633,N_10710);
or U10933 (N_10933,N_10604,N_10730);
nor U10934 (N_10934,N_10601,N_10646);
or U10935 (N_10935,N_10796,N_10608);
nand U10936 (N_10936,N_10721,N_10657);
xnor U10937 (N_10937,N_10629,N_10751);
xnor U10938 (N_10938,N_10749,N_10632);
nor U10939 (N_10939,N_10643,N_10687);
nand U10940 (N_10940,N_10658,N_10739);
or U10941 (N_10941,N_10791,N_10661);
or U10942 (N_10942,N_10759,N_10605);
xor U10943 (N_10943,N_10724,N_10684);
or U10944 (N_10944,N_10670,N_10789);
or U10945 (N_10945,N_10727,N_10606);
nor U10946 (N_10946,N_10752,N_10743);
xnor U10947 (N_10947,N_10626,N_10741);
and U10948 (N_10948,N_10665,N_10614);
and U10949 (N_10949,N_10606,N_10784);
nand U10950 (N_10950,N_10711,N_10714);
nand U10951 (N_10951,N_10734,N_10626);
nor U10952 (N_10952,N_10656,N_10745);
and U10953 (N_10953,N_10772,N_10796);
and U10954 (N_10954,N_10790,N_10756);
nor U10955 (N_10955,N_10638,N_10681);
xnor U10956 (N_10956,N_10710,N_10711);
nand U10957 (N_10957,N_10771,N_10799);
nand U10958 (N_10958,N_10725,N_10687);
xor U10959 (N_10959,N_10745,N_10616);
and U10960 (N_10960,N_10741,N_10700);
nor U10961 (N_10961,N_10706,N_10643);
xnor U10962 (N_10962,N_10720,N_10718);
or U10963 (N_10963,N_10686,N_10634);
nand U10964 (N_10964,N_10751,N_10748);
xor U10965 (N_10965,N_10760,N_10610);
xnor U10966 (N_10966,N_10678,N_10756);
and U10967 (N_10967,N_10746,N_10753);
nor U10968 (N_10968,N_10696,N_10765);
xnor U10969 (N_10969,N_10726,N_10649);
and U10970 (N_10970,N_10624,N_10740);
xor U10971 (N_10971,N_10621,N_10766);
and U10972 (N_10972,N_10687,N_10709);
xor U10973 (N_10973,N_10647,N_10615);
xnor U10974 (N_10974,N_10783,N_10612);
or U10975 (N_10975,N_10646,N_10614);
and U10976 (N_10976,N_10709,N_10730);
and U10977 (N_10977,N_10697,N_10684);
nand U10978 (N_10978,N_10788,N_10756);
xor U10979 (N_10979,N_10712,N_10762);
xor U10980 (N_10980,N_10717,N_10662);
xnor U10981 (N_10981,N_10796,N_10601);
and U10982 (N_10982,N_10630,N_10758);
and U10983 (N_10983,N_10713,N_10622);
nand U10984 (N_10984,N_10670,N_10777);
or U10985 (N_10985,N_10681,N_10620);
nor U10986 (N_10986,N_10608,N_10711);
nor U10987 (N_10987,N_10733,N_10797);
xor U10988 (N_10988,N_10701,N_10716);
nand U10989 (N_10989,N_10636,N_10602);
xnor U10990 (N_10990,N_10690,N_10642);
xor U10991 (N_10991,N_10667,N_10793);
nand U10992 (N_10992,N_10775,N_10764);
nor U10993 (N_10993,N_10622,N_10744);
nand U10994 (N_10994,N_10773,N_10777);
xnor U10995 (N_10995,N_10674,N_10646);
nor U10996 (N_10996,N_10624,N_10799);
nor U10997 (N_10997,N_10653,N_10787);
nand U10998 (N_10998,N_10616,N_10699);
and U10999 (N_10999,N_10624,N_10690);
and U11000 (N_11000,N_10826,N_10880);
xor U11001 (N_11001,N_10944,N_10966);
or U11002 (N_11002,N_10800,N_10929);
nand U11003 (N_11003,N_10862,N_10946);
or U11004 (N_11004,N_10957,N_10968);
nor U11005 (N_11005,N_10941,N_10899);
nand U11006 (N_11006,N_10834,N_10808);
and U11007 (N_11007,N_10922,N_10937);
nand U11008 (N_11008,N_10902,N_10852);
xnor U11009 (N_11009,N_10934,N_10931);
or U11010 (N_11010,N_10991,N_10848);
nor U11011 (N_11011,N_10953,N_10909);
xnor U11012 (N_11012,N_10894,N_10915);
or U11013 (N_11013,N_10955,N_10866);
and U11014 (N_11014,N_10835,N_10947);
xnor U11015 (N_11015,N_10905,N_10853);
and U11016 (N_11016,N_10847,N_10861);
or U11017 (N_11017,N_10884,N_10986);
xnor U11018 (N_11018,N_10998,N_10978);
nor U11019 (N_11019,N_10839,N_10887);
xnor U11020 (N_11020,N_10833,N_10854);
nand U11021 (N_11021,N_10918,N_10988);
or U11022 (N_11022,N_10948,N_10958);
and U11023 (N_11023,N_10801,N_10867);
nand U11024 (N_11024,N_10802,N_10803);
or U11025 (N_11025,N_10960,N_10858);
xor U11026 (N_11026,N_10821,N_10811);
and U11027 (N_11027,N_10927,N_10885);
and U11028 (N_11028,N_10878,N_10871);
xor U11029 (N_11029,N_10954,N_10964);
nor U11030 (N_11030,N_10806,N_10895);
or U11031 (N_11031,N_10933,N_10889);
nor U11032 (N_11032,N_10831,N_10838);
and U11033 (N_11033,N_10903,N_10805);
and U11034 (N_11034,N_10945,N_10819);
and U11035 (N_11035,N_10837,N_10930);
or U11036 (N_11036,N_10864,N_10897);
nand U11037 (N_11037,N_10928,N_10807);
or U11038 (N_11038,N_10820,N_10891);
xor U11039 (N_11039,N_10976,N_10979);
nor U11040 (N_11040,N_10888,N_10855);
and U11041 (N_11041,N_10896,N_10993);
xor U11042 (N_11042,N_10876,N_10917);
nor U11043 (N_11043,N_10911,N_10812);
nand U11044 (N_11044,N_10875,N_10908);
nand U11045 (N_11045,N_10825,N_10967);
nor U11046 (N_11046,N_10938,N_10824);
and U11047 (N_11047,N_10890,N_10982);
nand U11048 (N_11048,N_10844,N_10935);
and U11049 (N_11049,N_10836,N_10870);
or U11050 (N_11050,N_10886,N_10857);
nor U11051 (N_11051,N_10990,N_10882);
nand U11052 (N_11052,N_10910,N_10921);
and U11053 (N_11053,N_10810,N_10950);
or U11054 (N_11054,N_10974,N_10830);
and U11055 (N_11055,N_10995,N_10850);
or U11056 (N_11056,N_10992,N_10984);
and U11057 (N_11057,N_10865,N_10939);
nand U11058 (N_11058,N_10809,N_10969);
nor U11059 (N_11059,N_10997,N_10814);
nand U11060 (N_11060,N_10999,N_10817);
and U11061 (N_11061,N_10851,N_10841);
nand U11062 (N_11062,N_10913,N_10828);
nand U11063 (N_11063,N_10980,N_10989);
and U11064 (N_11064,N_10822,N_10900);
or U11065 (N_11065,N_10951,N_10912);
or U11066 (N_11066,N_10879,N_10983);
nor U11067 (N_11067,N_10949,N_10985);
xnor U11068 (N_11068,N_10813,N_10972);
or U11069 (N_11069,N_10975,N_10860);
and U11070 (N_11070,N_10914,N_10981);
nor U11071 (N_11071,N_10919,N_10959);
or U11072 (N_11072,N_10881,N_10943);
or U11073 (N_11073,N_10877,N_10859);
nand U11074 (N_11074,N_10827,N_10987);
xor U11075 (N_11075,N_10977,N_10901);
nand U11076 (N_11076,N_10893,N_10904);
or U11077 (N_11077,N_10883,N_10940);
and U11078 (N_11078,N_10869,N_10936);
or U11079 (N_11079,N_10829,N_10868);
xor U11080 (N_11080,N_10823,N_10804);
or U11081 (N_11081,N_10892,N_10962);
xor U11082 (N_11082,N_10994,N_10816);
nand U11083 (N_11083,N_10970,N_10873);
or U11084 (N_11084,N_10872,N_10925);
nand U11085 (N_11085,N_10849,N_10920);
nor U11086 (N_11086,N_10874,N_10996);
and U11087 (N_11087,N_10863,N_10843);
and U11088 (N_11088,N_10842,N_10846);
or U11089 (N_11089,N_10956,N_10961);
xor U11090 (N_11090,N_10845,N_10856);
nor U11091 (N_11091,N_10815,N_10965);
and U11092 (N_11092,N_10840,N_10971);
xnor U11093 (N_11093,N_10907,N_10952);
and U11094 (N_11094,N_10923,N_10963);
or U11095 (N_11095,N_10926,N_10818);
and U11096 (N_11096,N_10898,N_10832);
nand U11097 (N_11097,N_10906,N_10973);
xor U11098 (N_11098,N_10942,N_10932);
nor U11099 (N_11099,N_10924,N_10916);
nor U11100 (N_11100,N_10808,N_10815);
xnor U11101 (N_11101,N_10977,N_10853);
and U11102 (N_11102,N_10924,N_10863);
nand U11103 (N_11103,N_10801,N_10932);
or U11104 (N_11104,N_10842,N_10888);
nand U11105 (N_11105,N_10965,N_10895);
and U11106 (N_11106,N_10844,N_10983);
nor U11107 (N_11107,N_10804,N_10840);
xor U11108 (N_11108,N_10827,N_10998);
or U11109 (N_11109,N_10884,N_10935);
or U11110 (N_11110,N_10854,N_10862);
xor U11111 (N_11111,N_10998,N_10937);
or U11112 (N_11112,N_10845,N_10891);
and U11113 (N_11113,N_10955,N_10946);
and U11114 (N_11114,N_10817,N_10881);
xnor U11115 (N_11115,N_10953,N_10945);
and U11116 (N_11116,N_10963,N_10856);
nand U11117 (N_11117,N_10948,N_10987);
and U11118 (N_11118,N_10997,N_10800);
nand U11119 (N_11119,N_10842,N_10985);
and U11120 (N_11120,N_10891,N_10857);
nand U11121 (N_11121,N_10951,N_10803);
and U11122 (N_11122,N_10939,N_10889);
xor U11123 (N_11123,N_10868,N_10885);
xnor U11124 (N_11124,N_10846,N_10997);
xor U11125 (N_11125,N_10832,N_10987);
and U11126 (N_11126,N_10956,N_10936);
and U11127 (N_11127,N_10878,N_10844);
xnor U11128 (N_11128,N_10808,N_10994);
and U11129 (N_11129,N_10957,N_10978);
xnor U11130 (N_11130,N_10804,N_10927);
and U11131 (N_11131,N_10985,N_10882);
and U11132 (N_11132,N_10962,N_10990);
nor U11133 (N_11133,N_10845,N_10928);
nor U11134 (N_11134,N_10973,N_10959);
nand U11135 (N_11135,N_10853,N_10993);
nor U11136 (N_11136,N_10866,N_10805);
xnor U11137 (N_11137,N_10977,N_10841);
nor U11138 (N_11138,N_10916,N_10901);
or U11139 (N_11139,N_10922,N_10939);
or U11140 (N_11140,N_10848,N_10864);
xor U11141 (N_11141,N_10975,N_10866);
xor U11142 (N_11142,N_10823,N_10826);
nor U11143 (N_11143,N_10999,N_10910);
or U11144 (N_11144,N_10967,N_10940);
and U11145 (N_11145,N_10859,N_10804);
nand U11146 (N_11146,N_10892,N_10898);
or U11147 (N_11147,N_10855,N_10944);
nand U11148 (N_11148,N_10962,N_10952);
xor U11149 (N_11149,N_10928,N_10881);
nand U11150 (N_11150,N_10823,N_10999);
or U11151 (N_11151,N_10968,N_10947);
or U11152 (N_11152,N_10834,N_10804);
xor U11153 (N_11153,N_10854,N_10850);
and U11154 (N_11154,N_10846,N_10879);
nand U11155 (N_11155,N_10942,N_10825);
nor U11156 (N_11156,N_10844,N_10832);
and U11157 (N_11157,N_10896,N_10909);
nor U11158 (N_11158,N_10838,N_10856);
or U11159 (N_11159,N_10856,N_10859);
xnor U11160 (N_11160,N_10802,N_10807);
or U11161 (N_11161,N_10959,N_10816);
nor U11162 (N_11162,N_10848,N_10866);
xor U11163 (N_11163,N_10955,N_10803);
xor U11164 (N_11164,N_10985,N_10926);
and U11165 (N_11165,N_10879,N_10922);
nand U11166 (N_11166,N_10970,N_10907);
nand U11167 (N_11167,N_10808,N_10822);
and U11168 (N_11168,N_10886,N_10842);
nand U11169 (N_11169,N_10812,N_10979);
or U11170 (N_11170,N_10972,N_10829);
nor U11171 (N_11171,N_10941,N_10991);
nor U11172 (N_11172,N_10911,N_10856);
or U11173 (N_11173,N_10960,N_10964);
nor U11174 (N_11174,N_10893,N_10914);
nor U11175 (N_11175,N_10806,N_10971);
xnor U11176 (N_11176,N_10964,N_10847);
xnor U11177 (N_11177,N_10965,N_10996);
and U11178 (N_11178,N_10948,N_10890);
and U11179 (N_11179,N_10972,N_10899);
xor U11180 (N_11180,N_10998,N_10933);
xor U11181 (N_11181,N_10943,N_10973);
xnor U11182 (N_11182,N_10813,N_10808);
and U11183 (N_11183,N_10969,N_10838);
or U11184 (N_11184,N_10935,N_10812);
nor U11185 (N_11185,N_10903,N_10862);
and U11186 (N_11186,N_10820,N_10988);
nor U11187 (N_11187,N_10845,N_10805);
nand U11188 (N_11188,N_10834,N_10986);
nor U11189 (N_11189,N_10826,N_10871);
and U11190 (N_11190,N_10912,N_10940);
xnor U11191 (N_11191,N_10893,N_10864);
or U11192 (N_11192,N_10934,N_10852);
nor U11193 (N_11193,N_10835,N_10904);
and U11194 (N_11194,N_10865,N_10832);
and U11195 (N_11195,N_10939,N_10883);
xor U11196 (N_11196,N_10839,N_10906);
nor U11197 (N_11197,N_10971,N_10829);
nor U11198 (N_11198,N_10874,N_10820);
and U11199 (N_11199,N_10804,N_10952);
nor U11200 (N_11200,N_11001,N_11156);
xnor U11201 (N_11201,N_11187,N_11168);
xor U11202 (N_11202,N_11029,N_11115);
nand U11203 (N_11203,N_11111,N_11157);
nor U11204 (N_11204,N_11191,N_11013);
nand U11205 (N_11205,N_11059,N_11000);
nand U11206 (N_11206,N_11167,N_11148);
and U11207 (N_11207,N_11002,N_11072);
nand U11208 (N_11208,N_11058,N_11186);
or U11209 (N_11209,N_11012,N_11037);
and U11210 (N_11210,N_11033,N_11022);
and U11211 (N_11211,N_11180,N_11026);
nand U11212 (N_11212,N_11052,N_11127);
nand U11213 (N_11213,N_11091,N_11155);
and U11214 (N_11214,N_11147,N_11025);
or U11215 (N_11215,N_11193,N_11032);
nand U11216 (N_11216,N_11090,N_11086);
xor U11217 (N_11217,N_11019,N_11014);
xor U11218 (N_11218,N_11095,N_11093);
xor U11219 (N_11219,N_11131,N_11063);
xor U11220 (N_11220,N_11088,N_11079);
xor U11221 (N_11221,N_11190,N_11015);
nand U11222 (N_11222,N_11182,N_11165);
nor U11223 (N_11223,N_11050,N_11011);
xnor U11224 (N_11224,N_11117,N_11141);
nor U11225 (N_11225,N_11046,N_11134);
xnor U11226 (N_11226,N_11142,N_11023);
nor U11227 (N_11227,N_11192,N_11089);
nand U11228 (N_11228,N_11097,N_11118);
or U11229 (N_11229,N_11101,N_11110);
nand U11230 (N_11230,N_11017,N_11080);
xnor U11231 (N_11231,N_11039,N_11051);
or U11232 (N_11232,N_11060,N_11172);
and U11233 (N_11233,N_11099,N_11040);
nor U11234 (N_11234,N_11116,N_11179);
and U11235 (N_11235,N_11024,N_11020);
nand U11236 (N_11236,N_11126,N_11105);
xor U11237 (N_11237,N_11087,N_11042);
xnor U11238 (N_11238,N_11004,N_11133);
and U11239 (N_11239,N_11043,N_11036);
and U11240 (N_11240,N_11177,N_11076);
and U11241 (N_11241,N_11061,N_11171);
xor U11242 (N_11242,N_11021,N_11034);
nand U11243 (N_11243,N_11189,N_11083);
xor U11244 (N_11244,N_11176,N_11175);
or U11245 (N_11245,N_11008,N_11062);
and U11246 (N_11246,N_11129,N_11082);
xnor U11247 (N_11247,N_11169,N_11140);
nor U11248 (N_11248,N_11085,N_11064);
or U11249 (N_11249,N_11006,N_11109);
nand U11250 (N_11250,N_11010,N_11098);
nor U11251 (N_11251,N_11054,N_11161);
nand U11252 (N_11252,N_11150,N_11130);
nand U11253 (N_11253,N_11031,N_11198);
and U11254 (N_11254,N_11145,N_11070);
xor U11255 (N_11255,N_11038,N_11068);
xnor U11256 (N_11256,N_11158,N_11128);
nor U11257 (N_11257,N_11151,N_11030);
nor U11258 (N_11258,N_11066,N_11112);
or U11259 (N_11259,N_11107,N_11119);
nand U11260 (N_11260,N_11184,N_11199);
nor U11261 (N_11261,N_11160,N_11166);
xnor U11262 (N_11262,N_11120,N_11122);
nand U11263 (N_11263,N_11195,N_11124);
and U11264 (N_11264,N_11188,N_11132);
and U11265 (N_11265,N_11194,N_11144);
nand U11266 (N_11266,N_11103,N_11067);
nand U11267 (N_11267,N_11139,N_11053);
nand U11268 (N_11268,N_11152,N_11009);
xnor U11269 (N_11269,N_11136,N_11041);
and U11270 (N_11270,N_11057,N_11075);
nand U11271 (N_11271,N_11018,N_11146);
nand U11272 (N_11272,N_11092,N_11096);
nor U11273 (N_11273,N_11178,N_11125);
xnor U11274 (N_11274,N_11035,N_11108);
and U11275 (N_11275,N_11028,N_11121);
and U11276 (N_11276,N_11164,N_11143);
xnor U11277 (N_11277,N_11163,N_11135);
nand U11278 (N_11278,N_11077,N_11016);
xor U11279 (N_11279,N_11003,N_11084);
xnor U11280 (N_11280,N_11047,N_11102);
nor U11281 (N_11281,N_11113,N_11069);
nor U11282 (N_11282,N_11170,N_11027);
nor U11283 (N_11283,N_11100,N_11007);
nand U11284 (N_11284,N_11123,N_11149);
xor U11285 (N_11285,N_11173,N_11137);
nand U11286 (N_11286,N_11162,N_11073);
and U11287 (N_11287,N_11159,N_11185);
nor U11288 (N_11288,N_11005,N_11074);
xnor U11289 (N_11289,N_11071,N_11197);
nand U11290 (N_11290,N_11065,N_11081);
nand U11291 (N_11291,N_11174,N_11055);
xnor U11292 (N_11292,N_11104,N_11106);
nand U11293 (N_11293,N_11049,N_11048);
xor U11294 (N_11294,N_11153,N_11094);
and U11295 (N_11295,N_11196,N_11114);
xnor U11296 (N_11296,N_11056,N_11078);
and U11297 (N_11297,N_11154,N_11138);
and U11298 (N_11298,N_11183,N_11044);
nand U11299 (N_11299,N_11045,N_11181);
nor U11300 (N_11300,N_11043,N_11103);
and U11301 (N_11301,N_11142,N_11031);
nand U11302 (N_11302,N_11006,N_11118);
and U11303 (N_11303,N_11029,N_11016);
nor U11304 (N_11304,N_11071,N_11096);
nand U11305 (N_11305,N_11070,N_11113);
nand U11306 (N_11306,N_11009,N_11028);
nand U11307 (N_11307,N_11193,N_11176);
or U11308 (N_11308,N_11177,N_11153);
and U11309 (N_11309,N_11138,N_11168);
nand U11310 (N_11310,N_11115,N_11061);
or U11311 (N_11311,N_11194,N_11029);
and U11312 (N_11312,N_11039,N_11091);
xor U11313 (N_11313,N_11071,N_11072);
or U11314 (N_11314,N_11006,N_11092);
nand U11315 (N_11315,N_11166,N_11059);
nor U11316 (N_11316,N_11013,N_11168);
nor U11317 (N_11317,N_11010,N_11155);
nand U11318 (N_11318,N_11142,N_11145);
and U11319 (N_11319,N_11015,N_11109);
or U11320 (N_11320,N_11019,N_11040);
and U11321 (N_11321,N_11181,N_11153);
nand U11322 (N_11322,N_11130,N_11047);
and U11323 (N_11323,N_11194,N_11117);
and U11324 (N_11324,N_11187,N_11108);
nor U11325 (N_11325,N_11005,N_11048);
and U11326 (N_11326,N_11143,N_11049);
nor U11327 (N_11327,N_11050,N_11093);
and U11328 (N_11328,N_11004,N_11092);
nand U11329 (N_11329,N_11154,N_11064);
nor U11330 (N_11330,N_11079,N_11004);
and U11331 (N_11331,N_11113,N_11141);
or U11332 (N_11332,N_11199,N_11040);
or U11333 (N_11333,N_11061,N_11114);
nor U11334 (N_11334,N_11105,N_11011);
xor U11335 (N_11335,N_11092,N_11083);
or U11336 (N_11336,N_11074,N_11099);
nand U11337 (N_11337,N_11159,N_11101);
nor U11338 (N_11338,N_11079,N_11107);
or U11339 (N_11339,N_11179,N_11088);
xnor U11340 (N_11340,N_11045,N_11191);
nand U11341 (N_11341,N_11108,N_11119);
nor U11342 (N_11342,N_11052,N_11031);
nand U11343 (N_11343,N_11150,N_11114);
and U11344 (N_11344,N_11151,N_11095);
or U11345 (N_11345,N_11188,N_11050);
nor U11346 (N_11346,N_11191,N_11008);
nor U11347 (N_11347,N_11030,N_11059);
or U11348 (N_11348,N_11138,N_11093);
nand U11349 (N_11349,N_11115,N_11043);
nor U11350 (N_11350,N_11003,N_11000);
nand U11351 (N_11351,N_11008,N_11156);
or U11352 (N_11352,N_11045,N_11154);
xnor U11353 (N_11353,N_11130,N_11111);
or U11354 (N_11354,N_11036,N_11121);
nand U11355 (N_11355,N_11122,N_11103);
xor U11356 (N_11356,N_11044,N_11038);
nand U11357 (N_11357,N_11173,N_11136);
or U11358 (N_11358,N_11065,N_11087);
nor U11359 (N_11359,N_11068,N_11023);
or U11360 (N_11360,N_11122,N_11074);
and U11361 (N_11361,N_11194,N_11132);
or U11362 (N_11362,N_11130,N_11021);
and U11363 (N_11363,N_11093,N_11124);
nor U11364 (N_11364,N_11128,N_11090);
nand U11365 (N_11365,N_11096,N_11006);
or U11366 (N_11366,N_11146,N_11092);
or U11367 (N_11367,N_11121,N_11115);
xnor U11368 (N_11368,N_11116,N_11062);
nand U11369 (N_11369,N_11133,N_11012);
or U11370 (N_11370,N_11182,N_11121);
nand U11371 (N_11371,N_11006,N_11113);
or U11372 (N_11372,N_11041,N_11113);
nand U11373 (N_11373,N_11167,N_11020);
and U11374 (N_11374,N_11134,N_11194);
nor U11375 (N_11375,N_11169,N_11009);
nand U11376 (N_11376,N_11170,N_11187);
xor U11377 (N_11377,N_11161,N_11094);
nand U11378 (N_11378,N_11094,N_11099);
or U11379 (N_11379,N_11167,N_11151);
or U11380 (N_11380,N_11168,N_11188);
xor U11381 (N_11381,N_11195,N_11004);
or U11382 (N_11382,N_11006,N_11059);
nand U11383 (N_11383,N_11045,N_11171);
nand U11384 (N_11384,N_11152,N_11080);
nor U11385 (N_11385,N_11058,N_11124);
nand U11386 (N_11386,N_11174,N_11196);
or U11387 (N_11387,N_11030,N_11067);
xnor U11388 (N_11388,N_11097,N_11100);
xor U11389 (N_11389,N_11127,N_11049);
xor U11390 (N_11390,N_11052,N_11185);
nand U11391 (N_11391,N_11171,N_11156);
nor U11392 (N_11392,N_11080,N_11096);
or U11393 (N_11393,N_11191,N_11088);
and U11394 (N_11394,N_11114,N_11131);
and U11395 (N_11395,N_11165,N_11119);
and U11396 (N_11396,N_11173,N_11130);
xnor U11397 (N_11397,N_11001,N_11065);
or U11398 (N_11398,N_11156,N_11190);
and U11399 (N_11399,N_11064,N_11099);
nor U11400 (N_11400,N_11325,N_11252);
or U11401 (N_11401,N_11270,N_11264);
xor U11402 (N_11402,N_11250,N_11365);
nor U11403 (N_11403,N_11315,N_11394);
and U11404 (N_11404,N_11388,N_11342);
xnor U11405 (N_11405,N_11219,N_11338);
nor U11406 (N_11406,N_11208,N_11251);
nor U11407 (N_11407,N_11396,N_11391);
nor U11408 (N_11408,N_11395,N_11268);
and U11409 (N_11409,N_11284,N_11314);
nor U11410 (N_11410,N_11229,N_11383);
xnor U11411 (N_11411,N_11349,N_11234);
nor U11412 (N_11412,N_11231,N_11346);
or U11413 (N_11413,N_11387,N_11202);
nor U11414 (N_11414,N_11347,N_11243);
nand U11415 (N_11415,N_11211,N_11214);
xor U11416 (N_11416,N_11382,N_11205);
xor U11417 (N_11417,N_11262,N_11306);
or U11418 (N_11418,N_11351,N_11369);
nor U11419 (N_11419,N_11294,N_11312);
xor U11420 (N_11420,N_11386,N_11226);
nor U11421 (N_11421,N_11275,N_11267);
and U11422 (N_11422,N_11355,N_11271);
nor U11423 (N_11423,N_11305,N_11381);
nand U11424 (N_11424,N_11299,N_11311);
and U11425 (N_11425,N_11269,N_11255);
and U11426 (N_11426,N_11363,N_11240);
nand U11427 (N_11427,N_11206,N_11204);
nor U11428 (N_11428,N_11374,N_11380);
nand U11429 (N_11429,N_11224,N_11333);
nor U11430 (N_11430,N_11222,N_11225);
nand U11431 (N_11431,N_11335,N_11308);
and U11432 (N_11432,N_11258,N_11296);
and U11433 (N_11433,N_11307,N_11354);
and U11434 (N_11434,N_11377,N_11353);
nand U11435 (N_11435,N_11359,N_11279);
and U11436 (N_11436,N_11336,N_11232);
or U11437 (N_11437,N_11301,N_11272);
nand U11438 (N_11438,N_11261,N_11352);
or U11439 (N_11439,N_11332,N_11276);
xor U11440 (N_11440,N_11337,N_11370);
nor U11441 (N_11441,N_11334,N_11249);
nor U11442 (N_11442,N_11298,N_11357);
nand U11443 (N_11443,N_11227,N_11378);
nand U11444 (N_11444,N_11282,N_11285);
nor U11445 (N_11445,N_11319,N_11239);
nand U11446 (N_11446,N_11253,N_11313);
xor U11447 (N_11447,N_11247,N_11291);
nor U11448 (N_11448,N_11361,N_11260);
xnor U11449 (N_11449,N_11230,N_11274);
nor U11450 (N_11450,N_11310,N_11241);
xnor U11451 (N_11451,N_11340,N_11341);
or U11452 (N_11452,N_11254,N_11398);
and U11453 (N_11453,N_11295,N_11364);
nand U11454 (N_11454,N_11372,N_11280);
xnor U11455 (N_11455,N_11327,N_11287);
or U11456 (N_11456,N_11331,N_11259);
and U11457 (N_11457,N_11366,N_11278);
nor U11458 (N_11458,N_11368,N_11360);
or U11459 (N_11459,N_11302,N_11200);
and U11460 (N_11460,N_11213,N_11290);
nor U11461 (N_11461,N_11236,N_11309);
or U11462 (N_11462,N_11317,N_11246);
nand U11463 (N_11463,N_11242,N_11273);
nor U11464 (N_11464,N_11212,N_11392);
nand U11465 (N_11465,N_11303,N_11304);
or U11466 (N_11466,N_11344,N_11399);
or U11467 (N_11467,N_11283,N_11218);
xor U11468 (N_11468,N_11238,N_11358);
or U11469 (N_11469,N_11318,N_11384);
nor U11470 (N_11470,N_11362,N_11201);
xnor U11471 (N_11471,N_11235,N_11393);
or U11472 (N_11472,N_11356,N_11379);
or U11473 (N_11473,N_11328,N_11286);
xnor U11474 (N_11474,N_11373,N_11376);
and U11475 (N_11475,N_11281,N_11322);
xor U11476 (N_11476,N_11210,N_11220);
and U11477 (N_11477,N_11256,N_11316);
xnor U11478 (N_11478,N_11223,N_11217);
or U11479 (N_11479,N_11324,N_11350);
xnor U11480 (N_11480,N_11266,N_11248);
xor U11481 (N_11481,N_11300,N_11293);
nand U11482 (N_11482,N_11289,N_11339);
and U11483 (N_11483,N_11321,N_11237);
and U11484 (N_11484,N_11367,N_11233);
xnor U11485 (N_11485,N_11209,N_11348);
or U11486 (N_11486,N_11292,N_11390);
xnor U11487 (N_11487,N_11215,N_11297);
nor U11488 (N_11488,N_11323,N_11216);
or U11489 (N_11489,N_11263,N_11320);
nor U11490 (N_11490,N_11371,N_11265);
nand U11491 (N_11491,N_11203,N_11326);
nand U11492 (N_11492,N_11245,N_11288);
nor U11493 (N_11493,N_11330,N_11397);
and U11494 (N_11494,N_11389,N_11345);
nor U11495 (N_11495,N_11375,N_11207);
nor U11496 (N_11496,N_11329,N_11385);
nor U11497 (N_11497,N_11257,N_11277);
xor U11498 (N_11498,N_11221,N_11244);
and U11499 (N_11499,N_11343,N_11228);
and U11500 (N_11500,N_11333,N_11311);
and U11501 (N_11501,N_11301,N_11222);
xnor U11502 (N_11502,N_11252,N_11233);
nor U11503 (N_11503,N_11355,N_11398);
nor U11504 (N_11504,N_11378,N_11310);
nor U11505 (N_11505,N_11217,N_11208);
or U11506 (N_11506,N_11281,N_11394);
xor U11507 (N_11507,N_11363,N_11208);
nor U11508 (N_11508,N_11219,N_11362);
and U11509 (N_11509,N_11325,N_11266);
nor U11510 (N_11510,N_11347,N_11314);
nor U11511 (N_11511,N_11233,N_11227);
or U11512 (N_11512,N_11337,N_11394);
nor U11513 (N_11513,N_11350,N_11300);
nand U11514 (N_11514,N_11325,N_11238);
nand U11515 (N_11515,N_11343,N_11312);
nor U11516 (N_11516,N_11348,N_11246);
xnor U11517 (N_11517,N_11258,N_11321);
nor U11518 (N_11518,N_11232,N_11251);
nor U11519 (N_11519,N_11370,N_11351);
xnor U11520 (N_11520,N_11322,N_11222);
xnor U11521 (N_11521,N_11373,N_11358);
and U11522 (N_11522,N_11313,N_11312);
xnor U11523 (N_11523,N_11380,N_11205);
or U11524 (N_11524,N_11203,N_11202);
xnor U11525 (N_11525,N_11326,N_11295);
nand U11526 (N_11526,N_11321,N_11322);
and U11527 (N_11527,N_11293,N_11330);
and U11528 (N_11528,N_11376,N_11235);
xor U11529 (N_11529,N_11291,N_11361);
and U11530 (N_11530,N_11377,N_11260);
nor U11531 (N_11531,N_11361,N_11326);
and U11532 (N_11532,N_11321,N_11293);
nor U11533 (N_11533,N_11238,N_11315);
and U11534 (N_11534,N_11299,N_11296);
and U11535 (N_11535,N_11396,N_11205);
xor U11536 (N_11536,N_11228,N_11217);
xor U11537 (N_11537,N_11354,N_11390);
xor U11538 (N_11538,N_11333,N_11369);
xor U11539 (N_11539,N_11254,N_11253);
nor U11540 (N_11540,N_11392,N_11250);
nor U11541 (N_11541,N_11309,N_11295);
and U11542 (N_11542,N_11308,N_11325);
or U11543 (N_11543,N_11258,N_11294);
or U11544 (N_11544,N_11262,N_11252);
nand U11545 (N_11545,N_11386,N_11392);
and U11546 (N_11546,N_11357,N_11251);
xnor U11547 (N_11547,N_11336,N_11299);
nor U11548 (N_11548,N_11280,N_11237);
nand U11549 (N_11549,N_11272,N_11351);
xor U11550 (N_11550,N_11319,N_11376);
and U11551 (N_11551,N_11235,N_11367);
nor U11552 (N_11552,N_11225,N_11296);
nand U11553 (N_11553,N_11334,N_11265);
xor U11554 (N_11554,N_11241,N_11219);
or U11555 (N_11555,N_11342,N_11322);
xor U11556 (N_11556,N_11285,N_11367);
or U11557 (N_11557,N_11324,N_11293);
and U11558 (N_11558,N_11280,N_11353);
xor U11559 (N_11559,N_11252,N_11300);
or U11560 (N_11560,N_11238,N_11226);
nor U11561 (N_11561,N_11200,N_11358);
nor U11562 (N_11562,N_11252,N_11200);
nor U11563 (N_11563,N_11273,N_11330);
and U11564 (N_11564,N_11321,N_11308);
or U11565 (N_11565,N_11219,N_11394);
and U11566 (N_11566,N_11365,N_11277);
and U11567 (N_11567,N_11236,N_11390);
nand U11568 (N_11568,N_11286,N_11227);
nand U11569 (N_11569,N_11304,N_11246);
and U11570 (N_11570,N_11370,N_11359);
nor U11571 (N_11571,N_11232,N_11361);
nor U11572 (N_11572,N_11253,N_11334);
or U11573 (N_11573,N_11380,N_11294);
and U11574 (N_11574,N_11275,N_11289);
nor U11575 (N_11575,N_11211,N_11306);
nand U11576 (N_11576,N_11368,N_11369);
or U11577 (N_11577,N_11305,N_11276);
nor U11578 (N_11578,N_11358,N_11225);
and U11579 (N_11579,N_11249,N_11279);
or U11580 (N_11580,N_11266,N_11386);
nand U11581 (N_11581,N_11308,N_11213);
and U11582 (N_11582,N_11201,N_11359);
or U11583 (N_11583,N_11267,N_11264);
nor U11584 (N_11584,N_11316,N_11231);
nand U11585 (N_11585,N_11328,N_11374);
nand U11586 (N_11586,N_11309,N_11227);
nand U11587 (N_11587,N_11278,N_11227);
xnor U11588 (N_11588,N_11368,N_11314);
or U11589 (N_11589,N_11376,N_11225);
and U11590 (N_11590,N_11212,N_11315);
nor U11591 (N_11591,N_11299,N_11335);
and U11592 (N_11592,N_11393,N_11264);
and U11593 (N_11593,N_11295,N_11208);
and U11594 (N_11594,N_11318,N_11289);
and U11595 (N_11595,N_11312,N_11211);
nand U11596 (N_11596,N_11279,N_11271);
or U11597 (N_11597,N_11245,N_11258);
xor U11598 (N_11598,N_11242,N_11295);
and U11599 (N_11599,N_11216,N_11306);
nand U11600 (N_11600,N_11509,N_11598);
nor U11601 (N_11601,N_11450,N_11470);
nand U11602 (N_11602,N_11445,N_11536);
or U11603 (N_11603,N_11503,N_11468);
xnor U11604 (N_11604,N_11540,N_11518);
xor U11605 (N_11605,N_11519,N_11514);
and U11606 (N_11606,N_11500,N_11412);
nand U11607 (N_11607,N_11483,N_11444);
or U11608 (N_11608,N_11501,N_11590);
and U11609 (N_11609,N_11596,N_11471);
nor U11610 (N_11610,N_11581,N_11441);
xnor U11611 (N_11611,N_11517,N_11438);
or U11612 (N_11612,N_11460,N_11406);
xor U11613 (N_11613,N_11543,N_11499);
and U11614 (N_11614,N_11402,N_11548);
or U11615 (N_11615,N_11537,N_11400);
nand U11616 (N_11616,N_11454,N_11510);
and U11617 (N_11617,N_11436,N_11493);
nand U11618 (N_11618,N_11492,N_11439);
nand U11619 (N_11619,N_11549,N_11452);
xnor U11620 (N_11620,N_11588,N_11552);
nor U11621 (N_11621,N_11530,N_11404);
xor U11622 (N_11622,N_11411,N_11472);
xnor U11623 (N_11623,N_11481,N_11521);
or U11624 (N_11624,N_11496,N_11467);
nand U11625 (N_11625,N_11599,N_11557);
or U11626 (N_11626,N_11433,N_11461);
nand U11627 (N_11627,N_11583,N_11463);
nor U11628 (N_11628,N_11574,N_11538);
or U11629 (N_11629,N_11429,N_11531);
and U11630 (N_11630,N_11544,N_11443);
xor U11631 (N_11631,N_11432,N_11416);
nand U11632 (N_11632,N_11527,N_11555);
or U11633 (N_11633,N_11569,N_11423);
and U11634 (N_11634,N_11413,N_11586);
and U11635 (N_11635,N_11448,N_11535);
and U11636 (N_11636,N_11462,N_11449);
and U11637 (N_11637,N_11431,N_11458);
or U11638 (N_11638,N_11560,N_11502);
or U11639 (N_11639,N_11512,N_11559);
nor U11640 (N_11640,N_11484,N_11589);
nand U11641 (N_11641,N_11587,N_11465);
nand U11642 (N_11642,N_11410,N_11524);
nand U11643 (N_11643,N_11504,N_11425);
nand U11644 (N_11644,N_11466,N_11577);
xnor U11645 (N_11645,N_11525,N_11526);
nor U11646 (N_11646,N_11424,N_11422);
or U11647 (N_11647,N_11522,N_11476);
or U11648 (N_11648,N_11533,N_11409);
nand U11649 (N_11649,N_11579,N_11405);
nor U11650 (N_11650,N_11584,N_11447);
or U11651 (N_11651,N_11529,N_11572);
nand U11652 (N_11652,N_11553,N_11515);
nand U11653 (N_11653,N_11506,N_11511);
xnor U11654 (N_11654,N_11539,N_11532);
or U11655 (N_11655,N_11440,N_11457);
xor U11656 (N_11656,N_11428,N_11495);
nor U11657 (N_11657,N_11573,N_11566);
nor U11658 (N_11658,N_11464,N_11480);
and U11659 (N_11659,N_11451,N_11534);
and U11660 (N_11660,N_11592,N_11407);
xnor U11661 (N_11661,N_11561,N_11489);
or U11662 (N_11662,N_11568,N_11547);
nor U11663 (N_11663,N_11528,N_11418);
nand U11664 (N_11664,N_11459,N_11415);
nand U11665 (N_11665,N_11571,N_11508);
xor U11666 (N_11666,N_11497,N_11585);
or U11667 (N_11667,N_11565,N_11490);
xor U11668 (N_11668,N_11437,N_11469);
xor U11669 (N_11669,N_11487,N_11505);
or U11670 (N_11670,N_11550,N_11541);
or U11671 (N_11671,N_11551,N_11419);
and U11672 (N_11672,N_11417,N_11485);
xor U11673 (N_11673,N_11401,N_11414);
and U11674 (N_11674,N_11546,N_11435);
or U11675 (N_11675,N_11478,N_11421);
or U11676 (N_11676,N_11595,N_11523);
nor U11677 (N_11677,N_11580,N_11576);
or U11678 (N_11678,N_11455,N_11430);
and U11679 (N_11679,N_11516,N_11442);
nand U11680 (N_11680,N_11542,N_11426);
nor U11681 (N_11681,N_11403,N_11582);
and U11682 (N_11682,N_11474,N_11507);
nor U11683 (N_11683,N_11498,N_11591);
nor U11684 (N_11684,N_11488,N_11558);
nand U11685 (N_11685,N_11434,N_11570);
or U11686 (N_11686,N_11486,N_11427);
xor U11687 (N_11687,N_11594,N_11562);
or U11688 (N_11688,N_11479,N_11554);
xor U11689 (N_11689,N_11456,N_11491);
or U11690 (N_11690,N_11482,N_11494);
and U11691 (N_11691,N_11597,N_11475);
xor U11692 (N_11692,N_11556,N_11453);
nor U11693 (N_11693,N_11593,N_11477);
nand U11694 (N_11694,N_11563,N_11513);
and U11695 (N_11695,N_11567,N_11578);
nand U11696 (N_11696,N_11420,N_11564);
and U11697 (N_11697,N_11545,N_11473);
nand U11698 (N_11698,N_11408,N_11446);
nor U11699 (N_11699,N_11575,N_11520);
nand U11700 (N_11700,N_11404,N_11403);
and U11701 (N_11701,N_11522,N_11545);
xnor U11702 (N_11702,N_11588,N_11509);
xor U11703 (N_11703,N_11527,N_11420);
nand U11704 (N_11704,N_11492,N_11549);
xnor U11705 (N_11705,N_11525,N_11586);
nor U11706 (N_11706,N_11456,N_11515);
nand U11707 (N_11707,N_11461,N_11488);
xnor U11708 (N_11708,N_11509,N_11407);
nand U11709 (N_11709,N_11404,N_11545);
or U11710 (N_11710,N_11595,N_11551);
and U11711 (N_11711,N_11480,N_11411);
or U11712 (N_11712,N_11525,N_11556);
xnor U11713 (N_11713,N_11502,N_11428);
or U11714 (N_11714,N_11438,N_11590);
and U11715 (N_11715,N_11560,N_11541);
and U11716 (N_11716,N_11443,N_11403);
or U11717 (N_11717,N_11598,N_11584);
and U11718 (N_11718,N_11571,N_11549);
or U11719 (N_11719,N_11501,N_11422);
nor U11720 (N_11720,N_11582,N_11401);
nand U11721 (N_11721,N_11435,N_11564);
nand U11722 (N_11722,N_11560,N_11557);
nand U11723 (N_11723,N_11576,N_11588);
and U11724 (N_11724,N_11570,N_11415);
xnor U11725 (N_11725,N_11446,N_11474);
or U11726 (N_11726,N_11572,N_11472);
nand U11727 (N_11727,N_11413,N_11400);
or U11728 (N_11728,N_11576,N_11489);
nand U11729 (N_11729,N_11517,N_11499);
nor U11730 (N_11730,N_11585,N_11403);
and U11731 (N_11731,N_11535,N_11456);
and U11732 (N_11732,N_11404,N_11572);
xor U11733 (N_11733,N_11571,N_11588);
or U11734 (N_11734,N_11550,N_11428);
xor U11735 (N_11735,N_11538,N_11410);
xor U11736 (N_11736,N_11465,N_11538);
xor U11737 (N_11737,N_11510,N_11550);
and U11738 (N_11738,N_11588,N_11530);
or U11739 (N_11739,N_11539,N_11404);
and U11740 (N_11740,N_11418,N_11590);
or U11741 (N_11741,N_11507,N_11468);
and U11742 (N_11742,N_11539,N_11442);
and U11743 (N_11743,N_11500,N_11486);
and U11744 (N_11744,N_11514,N_11598);
nand U11745 (N_11745,N_11480,N_11594);
and U11746 (N_11746,N_11480,N_11459);
xnor U11747 (N_11747,N_11475,N_11543);
nor U11748 (N_11748,N_11476,N_11410);
nand U11749 (N_11749,N_11578,N_11453);
xor U11750 (N_11750,N_11568,N_11510);
xnor U11751 (N_11751,N_11439,N_11531);
nor U11752 (N_11752,N_11561,N_11524);
xor U11753 (N_11753,N_11447,N_11597);
nor U11754 (N_11754,N_11589,N_11579);
or U11755 (N_11755,N_11539,N_11449);
or U11756 (N_11756,N_11422,N_11575);
xnor U11757 (N_11757,N_11548,N_11497);
or U11758 (N_11758,N_11435,N_11425);
nand U11759 (N_11759,N_11440,N_11561);
nand U11760 (N_11760,N_11519,N_11506);
nand U11761 (N_11761,N_11400,N_11559);
nor U11762 (N_11762,N_11454,N_11521);
xor U11763 (N_11763,N_11531,N_11402);
nand U11764 (N_11764,N_11596,N_11482);
xnor U11765 (N_11765,N_11515,N_11443);
nand U11766 (N_11766,N_11435,N_11414);
or U11767 (N_11767,N_11434,N_11413);
or U11768 (N_11768,N_11473,N_11564);
nand U11769 (N_11769,N_11449,N_11426);
nand U11770 (N_11770,N_11526,N_11517);
nand U11771 (N_11771,N_11591,N_11581);
or U11772 (N_11772,N_11404,N_11514);
and U11773 (N_11773,N_11587,N_11520);
nand U11774 (N_11774,N_11553,N_11543);
nand U11775 (N_11775,N_11497,N_11593);
nor U11776 (N_11776,N_11434,N_11443);
nor U11777 (N_11777,N_11495,N_11414);
xnor U11778 (N_11778,N_11470,N_11415);
nand U11779 (N_11779,N_11433,N_11572);
nor U11780 (N_11780,N_11472,N_11430);
nor U11781 (N_11781,N_11442,N_11572);
nand U11782 (N_11782,N_11413,N_11459);
or U11783 (N_11783,N_11497,N_11571);
xnor U11784 (N_11784,N_11436,N_11495);
or U11785 (N_11785,N_11581,N_11437);
and U11786 (N_11786,N_11518,N_11529);
nor U11787 (N_11787,N_11530,N_11462);
xor U11788 (N_11788,N_11412,N_11563);
nor U11789 (N_11789,N_11502,N_11477);
nand U11790 (N_11790,N_11496,N_11437);
and U11791 (N_11791,N_11584,N_11423);
nand U11792 (N_11792,N_11542,N_11590);
nor U11793 (N_11793,N_11456,N_11510);
xor U11794 (N_11794,N_11440,N_11581);
or U11795 (N_11795,N_11441,N_11443);
nor U11796 (N_11796,N_11439,N_11522);
xnor U11797 (N_11797,N_11461,N_11426);
nor U11798 (N_11798,N_11595,N_11440);
and U11799 (N_11799,N_11575,N_11454);
and U11800 (N_11800,N_11617,N_11712);
and U11801 (N_11801,N_11758,N_11764);
and U11802 (N_11802,N_11766,N_11660);
xor U11803 (N_11803,N_11747,N_11626);
nand U11804 (N_11804,N_11648,N_11615);
or U11805 (N_11805,N_11789,N_11668);
xor U11806 (N_11806,N_11704,N_11724);
nand U11807 (N_11807,N_11769,N_11646);
xnor U11808 (N_11808,N_11672,N_11643);
or U11809 (N_11809,N_11654,N_11651);
or U11810 (N_11810,N_11720,N_11784);
nand U11811 (N_11811,N_11698,N_11703);
nor U11812 (N_11812,N_11708,N_11790);
or U11813 (N_11813,N_11604,N_11701);
and U11814 (N_11814,N_11762,N_11713);
xor U11815 (N_11815,N_11692,N_11787);
xor U11816 (N_11816,N_11602,N_11730);
or U11817 (N_11817,N_11771,N_11669);
xnor U11818 (N_11818,N_11687,N_11773);
nand U11819 (N_11819,N_11661,N_11753);
xor U11820 (N_11820,N_11735,N_11685);
nand U11821 (N_11821,N_11737,N_11746);
or U11822 (N_11822,N_11624,N_11676);
nand U11823 (N_11823,N_11709,N_11638);
nor U11824 (N_11824,N_11745,N_11616);
nor U11825 (N_11825,N_11622,N_11774);
or U11826 (N_11826,N_11722,N_11697);
nor U11827 (N_11827,N_11788,N_11621);
or U11828 (N_11828,N_11628,N_11796);
xor U11829 (N_11829,N_11742,N_11752);
or U11830 (N_11830,N_11641,N_11770);
nand U11831 (N_11831,N_11663,N_11798);
nor U11832 (N_11832,N_11680,N_11711);
and U11833 (N_11833,N_11623,N_11736);
and U11834 (N_11834,N_11652,N_11656);
and U11835 (N_11835,N_11781,N_11734);
nor U11836 (N_11836,N_11755,N_11750);
and U11837 (N_11837,N_11645,N_11792);
nand U11838 (N_11838,N_11657,N_11740);
nor U11839 (N_11839,N_11632,N_11670);
and U11840 (N_11840,N_11760,N_11705);
xnor U11841 (N_11841,N_11639,N_11716);
or U11842 (N_11842,N_11649,N_11797);
nand U11843 (N_11843,N_11761,N_11681);
nor U11844 (N_11844,N_11719,N_11603);
nand U11845 (N_11845,N_11667,N_11674);
nor U11846 (N_11846,N_11637,N_11644);
nor U11847 (N_11847,N_11795,N_11723);
xnor U11848 (N_11848,N_11631,N_11633);
or U11849 (N_11849,N_11664,N_11763);
nor U11850 (N_11850,N_11739,N_11780);
nand U11851 (N_11851,N_11694,N_11725);
or U11852 (N_11852,N_11791,N_11715);
xor U11853 (N_11853,N_11741,N_11690);
nor U11854 (N_11854,N_11749,N_11678);
nand U11855 (N_11855,N_11608,N_11707);
xnor U11856 (N_11856,N_11614,N_11612);
xnor U11857 (N_11857,N_11679,N_11684);
nor U11858 (N_11858,N_11733,N_11702);
and U11859 (N_11859,N_11748,N_11793);
nand U11860 (N_11860,N_11600,N_11611);
nor U11861 (N_11861,N_11688,N_11786);
xnor U11862 (N_11862,N_11779,N_11710);
nand U11863 (N_11863,N_11775,N_11659);
nor U11864 (N_11864,N_11671,N_11609);
or U11865 (N_11865,N_11635,N_11640);
and U11866 (N_11866,N_11744,N_11728);
xnor U11867 (N_11867,N_11768,N_11610);
xnor U11868 (N_11868,N_11642,N_11721);
and U11869 (N_11869,N_11647,N_11682);
xor U11870 (N_11870,N_11717,N_11756);
or U11871 (N_11871,N_11759,N_11605);
and U11872 (N_11872,N_11629,N_11606);
and U11873 (N_11873,N_11662,N_11767);
nor U11874 (N_11874,N_11613,N_11785);
nand U11875 (N_11875,N_11693,N_11625);
xnor U11876 (N_11876,N_11799,N_11655);
nor U11877 (N_11877,N_11630,N_11620);
nor U11878 (N_11878,N_11675,N_11607);
nor U11879 (N_11879,N_11757,N_11772);
xor U11880 (N_11880,N_11691,N_11778);
and U11881 (N_11881,N_11782,N_11650);
xnor U11882 (N_11882,N_11777,N_11738);
or U11883 (N_11883,N_11726,N_11618);
nor U11884 (N_11884,N_11732,N_11689);
and U11885 (N_11885,N_11636,N_11765);
xor U11886 (N_11886,N_11729,N_11666);
or U11887 (N_11887,N_11683,N_11794);
xor U11888 (N_11888,N_11699,N_11627);
or U11889 (N_11889,N_11706,N_11696);
and U11890 (N_11890,N_11695,N_11673);
and U11891 (N_11891,N_11634,N_11718);
and U11892 (N_11892,N_11677,N_11658);
nor U11893 (N_11893,N_11619,N_11754);
nand U11894 (N_11894,N_11783,N_11743);
nand U11895 (N_11895,N_11776,N_11653);
nor U11896 (N_11896,N_11700,N_11714);
and U11897 (N_11897,N_11727,N_11751);
xor U11898 (N_11898,N_11601,N_11686);
xnor U11899 (N_11899,N_11665,N_11731);
nand U11900 (N_11900,N_11790,N_11684);
or U11901 (N_11901,N_11634,N_11735);
nand U11902 (N_11902,N_11699,N_11704);
nand U11903 (N_11903,N_11615,N_11707);
nor U11904 (N_11904,N_11798,N_11605);
and U11905 (N_11905,N_11735,N_11606);
and U11906 (N_11906,N_11631,N_11634);
and U11907 (N_11907,N_11673,N_11781);
xor U11908 (N_11908,N_11691,N_11607);
and U11909 (N_11909,N_11700,N_11767);
nand U11910 (N_11910,N_11678,N_11721);
nand U11911 (N_11911,N_11667,N_11791);
xor U11912 (N_11912,N_11744,N_11662);
nand U11913 (N_11913,N_11734,N_11656);
or U11914 (N_11914,N_11740,N_11604);
or U11915 (N_11915,N_11662,N_11637);
xnor U11916 (N_11916,N_11798,N_11734);
and U11917 (N_11917,N_11765,N_11631);
nor U11918 (N_11918,N_11615,N_11794);
or U11919 (N_11919,N_11718,N_11711);
or U11920 (N_11920,N_11604,N_11623);
and U11921 (N_11921,N_11741,N_11675);
xnor U11922 (N_11922,N_11770,N_11609);
nand U11923 (N_11923,N_11669,N_11796);
nor U11924 (N_11924,N_11791,N_11684);
nor U11925 (N_11925,N_11650,N_11736);
nor U11926 (N_11926,N_11694,N_11649);
nand U11927 (N_11927,N_11665,N_11719);
xnor U11928 (N_11928,N_11732,N_11668);
nand U11929 (N_11929,N_11758,N_11660);
xor U11930 (N_11930,N_11695,N_11736);
nor U11931 (N_11931,N_11632,N_11734);
nor U11932 (N_11932,N_11719,N_11621);
nor U11933 (N_11933,N_11745,N_11744);
or U11934 (N_11934,N_11739,N_11700);
nand U11935 (N_11935,N_11684,N_11676);
nand U11936 (N_11936,N_11723,N_11750);
xor U11937 (N_11937,N_11661,N_11694);
nand U11938 (N_11938,N_11738,N_11663);
or U11939 (N_11939,N_11601,N_11787);
xor U11940 (N_11940,N_11696,N_11680);
nor U11941 (N_11941,N_11757,N_11786);
nor U11942 (N_11942,N_11627,N_11755);
xor U11943 (N_11943,N_11790,N_11700);
nor U11944 (N_11944,N_11624,N_11772);
nor U11945 (N_11945,N_11720,N_11711);
or U11946 (N_11946,N_11608,N_11762);
xnor U11947 (N_11947,N_11644,N_11654);
xnor U11948 (N_11948,N_11632,N_11726);
xnor U11949 (N_11949,N_11758,N_11671);
nand U11950 (N_11950,N_11684,N_11715);
nor U11951 (N_11951,N_11774,N_11626);
or U11952 (N_11952,N_11734,N_11783);
or U11953 (N_11953,N_11691,N_11663);
nand U11954 (N_11954,N_11747,N_11720);
nor U11955 (N_11955,N_11683,N_11731);
or U11956 (N_11956,N_11731,N_11729);
nor U11957 (N_11957,N_11785,N_11610);
nor U11958 (N_11958,N_11710,N_11712);
xnor U11959 (N_11959,N_11721,N_11619);
and U11960 (N_11960,N_11661,N_11673);
xnor U11961 (N_11961,N_11714,N_11791);
xnor U11962 (N_11962,N_11793,N_11783);
xor U11963 (N_11963,N_11700,N_11784);
nand U11964 (N_11964,N_11749,N_11736);
and U11965 (N_11965,N_11621,N_11668);
nand U11966 (N_11966,N_11608,N_11690);
nand U11967 (N_11967,N_11611,N_11788);
xor U11968 (N_11968,N_11610,N_11637);
and U11969 (N_11969,N_11656,N_11688);
and U11970 (N_11970,N_11696,N_11730);
and U11971 (N_11971,N_11796,N_11772);
nor U11972 (N_11972,N_11758,N_11734);
or U11973 (N_11973,N_11746,N_11759);
nor U11974 (N_11974,N_11795,N_11642);
xnor U11975 (N_11975,N_11675,N_11760);
nor U11976 (N_11976,N_11688,N_11637);
nor U11977 (N_11977,N_11681,N_11623);
nand U11978 (N_11978,N_11770,N_11793);
xor U11979 (N_11979,N_11679,N_11708);
and U11980 (N_11980,N_11798,N_11652);
and U11981 (N_11981,N_11793,N_11603);
nand U11982 (N_11982,N_11781,N_11650);
and U11983 (N_11983,N_11794,N_11701);
nand U11984 (N_11984,N_11782,N_11725);
xnor U11985 (N_11985,N_11662,N_11673);
xor U11986 (N_11986,N_11729,N_11607);
and U11987 (N_11987,N_11654,N_11660);
and U11988 (N_11988,N_11676,N_11655);
nor U11989 (N_11989,N_11723,N_11662);
nor U11990 (N_11990,N_11712,N_11752);
and U11991 (N_11991,N_11666,N_11746);
or U11992 (N_11992,N_11740,N_11733);
or U11993 (N_11993,N_11691,N_11633);
nand U11994 (N_11994,N_11765,N_11614);
nor U11995 (N_11995,N_11777,N_11739);
or U11996 (N_11996,N_11679,N_11619);
xor U11997 (N_11997,N_11639,N_11611);
nor U11998 (N_11998,N_11757,N_11627);
xor U11999 (N_11999,N_11727,N_11735);
and U12000 (N_12000,N_11870,N_11934);
nor U12001 (N_12001,N_11962,N_11957);
or U12002 (N_12002,N_11805,N_11857);
nand U12003 (N_12003,N_11856,N_11973);
and U12004 (N_12004,N_11922,N_11827);
nand U12005 (N_12005,N_11916,N_11800);
nand U12006 (N_12006,N_11877,N_11963);
xnor U12007 (N_12007,N_11904,N_11920);
xnor U12008 (N_12008,N_11888,N_11896);
nor U12009 (N_12009,N_11976,N_11863);
and U12010 (N_12010,N_11832,N_11915);
and U12011 (N_12011,N_11807,N_11983);
nand U12012 (N_12012,N_11897,N_11872);
nor U12013 (N_12013,N_11953,N_11844);
or U12014 (N_12014,N_11969,N_11909);
nor U12015 (N_12015,N_11955,N_11997);
nor U12016 (N_12016,N_11862,N_11813);
nor U12017 (N_12017,N_11802,N_11968);
and U12018 (N_12018,N_11944,N_11925);
nor U12019 (N_12019,N_11911,N_11865);
nor U12020 (N_12020,N_11937,N_11906);
nand U12021 (N_12021,N_11956,N_11831);
nand U12022 (N_12022,N_11900,N_11842);
xnor U12023 (N_12023,N_11892,N_11901);
or U12024 (N_12024,N_11986,N_11829);
xnor U12025 (N_12025,N_11891,N_11914);
nor U12026 (N_12026,N_11913,N_11946);
or U12027 (N_12027,N_11918,N_11905);
nor U12028 (N_12028,N_11975,N_11974);
nand U12029 (N_12029,N_11964,N_11853);
nor U12030 (N_12030,N_11887,N_11941);
and U12031 (N_12031,N_11818,N_11803);
and U12032 (N_12032,N_11868,N_11912);
xor U12033 (N_12033,N_11834,N_11855);
xnor U12034 (N_12034,N_11815,N_11902);
nand U12035 (N_12035,N_11826,N_11959);
xor U12036 (N_12036,N_11837,N_11819);
or U12037 (N_12037,N_11812,N_11972);
nor U12038 (N_12038,N_11879,N_11924);
xor U12039 (N_12039,N_11854,N_11951);
and U12040 (N_12040,N_11987,N_11820);
or U12041 (N_12041,N_11821,N_11971);
nand U12042 (N_12042,N_11928,N_11998);
or U12043 (N_12043,N_11871,N_11960);
and U12044 (N_12044,N_11991,N_11895);
xnor U12045 (N_12045,N_11874,N_11993);
or U12046 (N_12046,N_11889,N_11824);
and U12047 (N_12047,N_11977,N_11982);
and U12048 (N_12048,N_11808,N_11940);
or U12049 (N_12049,N_11929,N_11816);
or U12050 (N_12050,N_11876,N_11884);
and U12051 (N_12051,N_11910,N_11943);
and U12052 (N_12052,N_11867,N_11890);
xor U12053 (N_12053,N_11848,N_11878);
nand U12054 (N_12054,N_11994,N_11881);
xnor U12055 (N_12055,N_11858,N_11836);
and U12056 (N_12056,N_11840,N_11822);
and U12057 (N_12057,N_11948,N_11860);
or U12058 (N_12058,N_11980,N_11907);
and U12059 (N_12059,N_11875,N_11979);
or U12060 (N_12060,N_11893,N_11990);
nand U12061 (N_12061,N_11830,N_11961);
and U12062 (N_12062,N_11995,N_11882);
xor U12063 (N_12063,N_11869,N_11898);
and U12064 (N_12064,N_11847,N_11903);
or U12065 (N_12065,N_11978,N_11825);
nor U12066 (N_12066,N_11942,N_11801);
nand U12067 (N_12067,N_11885,N_11845);
nand U12068 (N_12068,N_11967,N_11873);
nand U12069 (N_12069,N_11970,N_11850);
or U12070 (N_12070,N_11930,N_11921);
xnor U12071 (N_12071,N_11849,N_11835);
and U12072 (N_12072,N_11949,N_11981);
or U12073 (N_12073,N_11814,N_11919);
nand U12074 (N_12074,N_11992,N_11952);
or U12075 (N_12075,N_11811,N_11843);
and U12076 (N_12076,N_11932,N_11859);
nor U12077 (N_12077,N_11935,N_11936);
nand U12078 (N_12078,N_11883,N_11939);
nor U12079 (N_12079,N_11861,N_11828);
xnor U12080 (N_12080,N_11846,N_11880);
nor U12081 (N_12081,N_11965,N_11851);
or U12082 (N_12082,N_11894,N_11908);
nand U12083 (N_12083,N_11804,N_11931);
and U12084 (N_12084,N_11886,N_11958);
nand U12085 (N_12085,N_11926,N_11833);
or U12086 (N_12086,N_11999,N_11938);
or U12087 (N_12087,N_11823,N_11864);
nand U12088 (N_12088,N_11806,N_11966);
or U12089 (N_12089,N_11923,N_11899);
nand U12090 (N_12090,N_11988,N_11927);
and U12091 (N_12091,N_11945,N_11950);
or U12092 (N_12092,N_11917,N_11838);
and U12093 (N_12093,N_11841,N_11810);
xnor U12094 (N_12094,N_11985,N_11954);
nor U12095 (N_12095,N_11852,N_11933);
or U12096 (N_12096,N_11989,N_11817);
xor U12097 (N_12097,N_11996,N_11947);
nand U12098 (N_12098,N_11839,N_11866);
or U12099 (N_12099,N_11809,N_11984);
nand U12100 (N_12100,N_11982,N_11867);
or U12101 (N_12101,N_11908,N_11890);
nand U12102 (N_12102,N_11877,N_11845);
nand U12103 (N_12103,N_11919,N_11885);
or U12104 (N_12104,N_11831,N_11820);
nand U12105 (N_12105,N_11805,N_11872);
xor U12106 (N_12106,N_11887,N_11953);
nand U12107 (N_12107,N_11964,N_11922);
or U12108 (N_12108,N_11869,N_11829);
xnor U12109 (N_12109,N_11916,N_11924);
xor U12110 (N_12110,N_11938,N_11985);
nor U12111 (N_12111,N_11923,N_11943);
and U12112 (N_12112,N_11994,N_11844);
nand U12113 (N_12113,N_11888,N_11816);
nand U12114 (N_12114,N_11996,N_11917);
and U12115 (N_12115,N_11889,N_11937);
nor U12116 (N_12116,N_11968,N_11856);
and U12117 (N_12117,N_11840,N_11978);
and U12118 (N_12118,N_11868,N_11923);
or U12119 (N_12119,N_11859,N_11917);
nor U12120 (N_12120,N_11961,N_11882);
and U12121 (N_12121,N_11907,N_11917);
or U12122 (N_12122,N_11968,N_11886);
xnor U12123 (N_12123,N_11866,N_11927);
xor U12124 (N_12124,N_11937,N_11996);
nor U12125 (N_12125,N_11922,N_11876);
nor U12126 (N_12126,N_11962,N_11926);
nand U12127 (N_12127,N_11802,N_11941);
and U12128 (N_12128,N_11842,N_11987);
or U12129 (N_12129,N_11975,N_11992);
or U12130 (N_12130,N_11808,N_11989);
or U12131 (N_12131,N_11975,N_11884);
or U12132 (N_12132,N_11998,N_11831);
nor U12133 (N_12133,N_11881,N_11892);
and U12134 (N_12134,N_11944,N_11959);
nand U12135 (N_12135,N_11912,N_11805);
nor U12136 (N_12136,N_11908,N_11830);
nand U12137 (N_12137,N_11968,N_11927);
nand U12138 (N_12138,N_11830,N_11825);
xnor U12139 (N_12139,N_11865,N_11879);
and U12140 (N_12140,N_11968,N_11881);
and U12141 (N_12141,N_11802,N_11822);
xor U12142 (N_12142,N_11819,N_11931);
or U12143 (N_12143,N_11973,N_11990);
and U12144 (N_12144,N_11987,N_11809);
xnor U12145 (N_12145,N_11944,N_11936);
nand U12146 (N_12146,N_11916,N_11853);
xnor U12147 (N_12147,N_11866,N_11841);
and U12148 (N_12148,N_11880,N_11810);
nor U12149 (N_12149,N_11947,N_11932);
xor U12150 (N_12150,N_11806,N_11896);
xor U12151 (N_12151,N_11874,N_11963);
xnor U12152 (N_12152,N_11937,N_11828);
nand U12153 (N_12153,N_11989,N_11813);
nand U12154 (N_12154,N_11976,N_11901);
nor U12155 (N_12155,N_11973,N_11923);
and U12156 (N_12156,N_11967,N_11804);
nand U12157 (N_12157,N_11956,N_11949);
or U12158 (N_12158,N_11997,N_11833);
nand U12159 (N_12159,N_11988,N_11995);
nand U12160 (N_12160,N_11986,N_11863);
nor U12161 (N_12161,N_11846,N_11967);
xnor U12162 (N_12162,N_11998,N_11921);
nor U12163 (N_12163,N_11804,N_11999);
nand U12164 (N_12164,N_11869,N_11953);
nor U12165 (N_12165,N_11887,N_11976);
nand U12166 (N_12166,N_11809,N_11916);
nor U12167 (N_12167,N_11907,N_11869);
or U12168 (N_12168,N_11930,N_11822);
and U12169 (N_12169,N_11816,N_11932);
and U12170 (N_12170,N_11971,N_11955);
xnor U12171 (N_12171,N_11873,N_11821);
and U12172 (N_12172,N_11883,N_11912);
xor U12173 (N_12173,N_11907,N_11962);
and U12174 (N_12174,N_11826,N_11907);
nand U12175 (N_12175,N_11896,N_11956);
or U12176 (N_12176,N_11984,N_11912);
xnor U12177 (N_12177,N_11866,N_11869);
nand U12178 (N_12178,N_11944,N_11888);
xor U12179 (N_12179,N_11895,N_11807);
or U12180 (N_12180,N_11817,N_11808);
nand U12181 (N_12181,N_11898,N_11989);
or U12182 (N_12182,N_11894,N_11974);
and U12183 (N_12183,N_11888,N_11970);
nor U12184 (N_12184,N_11933,N_11931);
nand U12185 (N_12185,N_11874,N_11871);
nand U12186 (N_12186,N_11978,N_11950);
or U12187 (N_12187,N_11896,N_11811);
nor U12188 (N_12188,N_11845,N_11927);
nor U12189 (N_12189,N_11811,N_11986);
and U12190 (N_12190,N_11958,N_11860);
or U12191 (N_12191,N_11846,N_11847);
and U12192 (N_12192,N_11812,N_11815);
xor U12193 (N_12193,N_11941,N_11844);
xnor U12194 (N_12194,N_11975,N_11837);
or U12195 (N_12195,N_11821,N_11896);
and U12196 (N_12196,N_11923,N_11878);
and U12197 (N_12197,N_11853,N_11961);
nand U12198 (N_12198,N_11821,N_11939);
or U12199 (N_12199,N_11848,N_11919);
and U12200 (N_12200,N_12021,N_12168);
or U12201 (N_12201,N_12138,N_12042);
xor U12202 (N_12202,N_12191,N_12088);
nand U12203 (N_12203,N_12057,N_12169);
nor U12204 (N_12204,N_12166,N_12159);
or U12205 (N_12205,N_12018,N_12133);
and U12206 (N_12206,N_12005,N_12094);
xor U12207 (N_12207,N_12091,N_12025);
xor U12208 (N_12208,N_12126,N_12188);
xor U12209 (N_12209,N_12074,N_12149);
or U12210 (N_12210,N_12006,N_12171);
xor U12211 (N_12211,N_12153,N_12002);
nand U12212 (N_12212,N_12031,N_12199);
and U12213 (N_12213,N_12010,N_12087);
nand U12214 (N_12214,N_12118,N_12061);
nor U12215 (N_12215,N_12064,N_12160);
or U12216 (N_12216,N_12148,N_12045);
nor U12217 (N_12217,N_12181,N_12072);
or U12218 (N_12218,N_12055,N_12154);
and U12219 (N_12219,N_12113,N_12189);
and U12220 (N_12220,N_12195,N_12043);
xnor U12221 (N_12221,N_12106,N_12032);
and U12222 (N_12222,N_12099,N_12077);
and U12223 (N_12223,N_12081,N_12130);
xor U12224 (N_12224,N_12066,N_12150);
nand U12225 (N_12225,N_12157,N_12170);
xnor U12226 (N_12226,N_12089,N_12011);
and U12227 (N_12227,N_12012,N_12140);
or U12228 (N_12228,N_12165,N_12047);
and U12229 (N_12229,N_12053,N_12164);
and U12230 (N_12230,N_12100,N_12052);
nand U12231 (N_12231,N_12039,N_12125);
and U12232 (N_12232,N_12007,N_12013);
nor U12233 (N_12233,N_12177,N_12004);
nand U12234 (N_12234,N_12186,N_12144);
and U12235 (N_12235,N_12070,N_12097);
nand U12236 (N_12236,N_12180,N_12062);
xnor U12237 (N_12237,N_12050,N_12085);
xor U12238 (N_12238,N_12082,N_12173);
xor U12239 (N_12239,N_12156,N_12112);
nor U12240 (N_12240,N_12001,N_12071);
or U12241 (N_12241,N_12029,N_12182);
nor U12242 (N_12242,N_12121,N_12016);
nand U12243 (N_12243,N_12022,N_12158);
xnor U12244 (N_12244,N_12184,N_12187);
nand U12245 (N_12245,N_12193,N_12017);
nand U12246 (N_12246,N_12054,N_12030);
xor U12247 (N_12247,N_12079,N_12178);
nor U12248 (N_12248,N_12101,N_12198);
nor U12249 (N_12249,N_12028,N_12110);
nand U12250 (N_12250,N_12080,N_12117);
and U12251 (N_12251,N_12145,N_12172);
xnor U12252 (N_12252,N_12076,N_12183);
nand U12253 (N_12253,N_12078,N_12034);
and U12254 (N_12254,N_12051,N_12147);
nand U12255 (N_12255,N_12197,N_12063);
and U12256 (N_12256,N_12041,N_12059);
xnor U12257 (N_12257,N_12049,N_12024);
nand U12258 (N_12258,N_12190,N_12015);
or U12259 (N_12259,N_12035,N_12105);
or U12260 (N_12260,N_12111,N_12132);
or U12261 (N_12261,N_12161,N_12037);
and U12262 (N_12262,N_12048,N_12095);
xnor U12263 (N_12263,N_12083,N_12033);
nand U12264 (N_12264,N_12142,N_12129);
nand U12265 (N_12265,N_12124,N_12019);
or U12266 (N_12266,N_12084,N_12155);
nand U12267 (N_12267,N_12162,N_12192);
and U12268 (N_12268,N_12056,N_12058);
or U12269 (N_12269,N_12127,N_12167);
nor U12270 (N_12270,N_12096,N_12067);
and U12271 (N_12271,N_12036,N_12009);
and U12272 (N_12272,N_12136,N_12090);
nor U12273 (N_12273,N_12065,N_12046);
xnor U12274 (N_12274,N_12093,N_12175);
or U12275 (N_12275,N_12073,N_12128);
xnor U12276 (N_12276,N_12040,N_12107);
or U12277 (N_12277,N_12027,N_12185);
xor U12278 (N_12278,N_12141,N_12163);
nand U12279 (N_12279,N_12176,N_12000);
xor U12280 (N_12280,N_12135,N_12060);
xor U12281 (N_12281,N_12120,N_12102);
or U12282 (N_12282,N_12092,N_12026);
nor U12283 (N_12283,N_12038,N_12194);
and U12284 (N_12284,N_12023,N_12008);
and U12285 (N_12285,N_12152,N_12139);
and U12286 (N_12286,N_12108,N_12134);
and U12287 (N_12287,N_12069,N_12151);
xor U12288 (N_12288,N_12122,N_12123);
or U12289 (N_12289,N_12119,N_12179);
nand U12290 (N_12290,N_12131,N_12086);
and U12291 (N_12291,N_12109,N_12115);
and U12292 (N_12292,N_12196,N_12146);
nand U12293 (N_12293,N_12068,N_12137);
xor U12294 (N_12294,N_12104,N_12014);
and U12295 (N_12295,N_12103,N_12044);
xor U12296 (N_12296,N_12003,N_12020);
nor U12297 (N_12297,N_12114,N_12116);
nand U12298 (N_12298,N_12143,N_12075);
or U12299 (N_12299,N_12174,N_12098);
xnor U12300 (N_12300,N_12093,N_12177);
and U12301 (N_12301,N_12081,N_12187);
and U12302 (N_12302,N_12123,N_12176);
xor U12303 (N_12303,N_12198,N_12111);
xnor U12304 (N_12304,N_12176,N_12192);
nand U12305 (N_12305,N_12198,N_12070);
and U12306 (N_12306,N_12135,N_12042);
nand U12307 (N_12307,N_12165,N_12054);
nor U12308 (N_12308,N_12083,N_12091);
nor U12309 (N_12309,N_12086,N_12103);
nand U12310 (N_12310,N_12171,N_12074);
xor U12311 (N_12311,N_12063,N_12185);
xor U12312 (N_12312,N_12135,N_12149);
nand U12313 (N_12313,N_12127,N_12094);
xnor U12314 (N_12314,N_12059,N_12167);
and U12315 (N_12315,N_12113,N_12196);
and U12316 (N_12316,N_12166,N_12165);
nor U12317 (N_12317,N_12183,N_12114);
xnor U12318 (N_12318,N_12036,N_12192);
nand U12319 (N_12319,N_12159,N_12199);
nor U12320 (N_12320,N_12023,N_12128);
and U12321 (N_12321,N_12111,N_12165);
or U12322 (N_12322,N_12137,N_12034);
nand U12323 (N_12323,N_12029,N_12088);
nor U12324 (N_12324,N_12125,N_12136);
nor U12325 (N_12325,N_12041,N_12107);
xor U12326 (N_12326,N_12126,N_12100);
nor U12327 (N_12327,N_12035,N_12028);
and U12328 (N_12328,N_12094,N_12105);
or U12329 (N_12329,N_12111,N_12012);
xnor U12330 (N_12330,N_12091,N_12119);
nor U12331 (N_12331,N_12167,N_12157);
nor U12332 (N_12332,N_12036,N_12135);
nand U12333 (N_12333,N_12064,N_12110);
nor U12334 (N_12334,N_12122,N_12112);
nand U12335 (N_12335,N_12093,N_12077);
or U12336 (N_12336,N_12100,N_12050);
nand U12337 (N_12337,N_12171,N_12049);
xnor U12338 (N_12338,N_12093,N_12072);
xor U12339 (N_12339,N_12197,N_12049);
and U12340 (N_12340,N_12190,N_12136);
or U12341 (N_12341,N_12175,N_12129);
nand U12342 (N_12342,N_12188,N_12180);
xor U12343 (N_12343,N_12086,N_12139);
or U12344 (N_12344,N_12046,N_12179);
nor U12345 (N_12345,N_12047,N_12174);
or U12346 (N_12346,N_12109,N_12155);
nor U12347 (N_12347,N_12003,N_12153);
and U12348 (N_12348,N_12062,N_12147);
or U12349 (N_12349,N_12090,N_12047);
nand U12350 (N_12350,N_12194,N_12002);
or U12351 (N_12351,N_12000,N_12066);
and U12352 (N_12352,N_12000,N_12117);
nor U12353 (N_12353,N_12132,N_12127);
nand U12354 (N_12354,N_12036,N_12038);
nor U12355 (N_12355,N_12134,N_12199);
and U12356 (N_12356,N_12154,N_12164);
nor U12357 (N_12357,N_12004,N_12085);
xor U12358 (N_12358,N_12139,N_12154);
or U12359 (N_12359,N_12000,N_12159);
and U12360 (N_12360,N_12123,N_12106);
nand U12361 (N_12361,N_12172,N_12141);
xnor U12362 (N_12362,N_12045,N_12032);
or U12363 (N_12363,N_12195,N_12005);
xor U12364 (N_12364,N_12111,N_12096);
nand U12365 (N_12365,N_12062,N_12199);
nand U12366 (N_12366,N_12162,N_12176);
nand U12367 (N_12367,N_12163,N_12153);
nor U12368 (N_12368,N_12182,N_12068);
xnor U12369 (N_12369,N_12078,N_12095);
and U12370 (N_12370,N_12183,N_12028);
nor U12371 (N_12371,N_12012,N_12177);
xnor U12372 (N_12372,N_12049,N_12066);
nand U12373 (N_12373,N_12098,N_12036);
nor U12374 (N_12374,N_12000,N_12093);
nand U12375 (N_12375,N_12019,N_12057);
nand U12376 (N_12376,N_12109,N_12172);
nor U12377 (N_12377,N_12133,N_12017);
and U12378 (N_12378,N_12059,N_12017);
nand U12379 (N_12379,N_12184,N_12006);
or U12380 (N_12380,N_12098,N_12195);
nand U12381 (N_12381,N_12057,N_12181);
or U12382 (N_12382,N_12178,N_12089);
xnor U12383 (N_12383,N_12127,N_12130);
nand U12384 (N_12384,N_12191,N_12161);
xnor U12385 (N_12385,N_12123,N_12195);
and U12386 (N_12386,N_12046,N_12051);
and U12387 (N_12387,N_12029,N_12141);
and U12388 (N_12388,N_12075,N_12074);
nor U12389 (N_12389,N_12128,N_12038);
and U12390 (N_12390,N_12052,N_12031);
nor U12391 (N_12391,N_12063,N_12005);
xnor U12392 (N_12392,N_12073,N_12094);
and U12393 (N_12393,N_12157,N_12147);
nand U12394 (N_12394,N_12127,N_12146);
or U12395 (N_12395,N_12100,N_12043);
nand U12396 (N_12396,N_12070,N_12047);
nor U12397 (N_12397,N_12008,N_12036);
nor U12398 (N_12398,N_12066,N_12071);
or U12399 (N_12399,N_12051,N_12044);
or U12400 (N_12400,N_12291,N_12264);
nand U12401 (N_12401,N_12324,N_12357);
or U12402 (N_12402,N_12240,N_12351);
xnor U12403 (N_12403,N_12295,N_12356);
nor U12404 (N_12404,N_12378,N_12304);
nor U12405 (N_12405,N_12346,N_12393);
xnor U12406 (N_12406,N_12321,N_12328);
nand U12407 (N_12407,N_12397,N_12394);
and U12408 (N_12408,N_12213,N_12230);
nor U12409 (N_12409,N_12276,N_12252);
nor U12410 (N_12410,N_12223,N_12358);
xor U12411 (N_12411,N_12238,N_12376);
and U12412 (N_12412,N_12244,N_12363);
nor U12413 (N_12413,N_12206,N_12292);
nand U12414 (N_12414,N_12282,N_12232);
xor U12415 (N_12415,N_12381,N_12314);
nor U12416 (N_12416,N_12391,N_12286);
and U12417 (N_12417,N_12388,N_12399);
and U12418 (N_12418,N_12253,N_12239);
and U12419 (N_12419,N_12260,N_12392);
or U12420 (N_12420,N_12247,N_12256);
nor U12421 (N_12421,N_12214,N_12250);
xor U12422 (N_12422,N_12315,N_12339);
and U12423 (N_12423,N_12348,N_12263);
or U12424 (N_12424,N_12202,N_12389);
nor U12425 (N_12425,N_12365,N_12246);
nor U12426 (N_12426,N_12287,N_12382);
nor U12427 (N_12427,N_12208,N_12320);
nand U12428 (N_12428,N_12267,N_12273);
and U12429 (N_12429,N_12296,N_12262);
nand U12430 (N_12430,N_12285,N_12300);
or U12431 (N_12431,N_12272,N_12369);
nor U12432 (N_12432,N_12241,N_12248);
and U12433 (N_12433,N_12279,N_12200);
and U12434 (N_12434,N_12340,N_12294);
nand U12435 (N_12435,N_12211,N_12362);
nand U12436 (N_12436,N_12234,N_12386);
or U12437 (N_12437,N_12305,N_12209);
xor U12438 (N_12438,N_12364,N_12341);
or U12439 (N_12439,N_12242,N_12281);
xor U12440 (N_12440,N_12205,N_12359);
nand U12441 (N_12441,N_12335,N_12387);
and U12442 (N_12442,N_12265,N_12374);
nand U12443 (N_12443,N_12350,N_12274);
or U12444 (N_12444,N_12227,N_12293);
and U12445 (N_12445,N_12354,N_12220);
nor U12446 (N_12446,N_12283,N_12236);
nand U12447 (N_12447,N_12380,N_12222);
xor U12448 (N_12448,N_12277,N_12210);
and U12449 (N_12449,N_12332,N_12280);
nor U12450 (N_12450,N_12224,N_12255);
nor U12451 (N_12451,N_12370,N_12371);
xnor U12452 (N_12452,N_12216,N_12366);
and U12453 (N_12453,N_12268,N_12311);
or U12454 (N_12454,N_12318,N_12334);
xor U12455 (N_12455,N_12212,N_12245);
and U12456 (N_12456,N_12217,N_12215);
xnor U12457 (N_12457,N_12372,N_12266);
and U12458 (N_12458,N_12322,N_12361);
xnor U12459 (N_12459,N_12390,N_12396);
and U12460 (N_12460,N_12302,N_12343);
nand U12461 (N_12461,N_12251,N_12352);
and U12462 (N_12462,N_12316,N_12275);
and U12463 (N_12463,N_12312,N_12367);
nor U12464 (N_12464,N_12298,N_12329);
or U12465 (N_12465,N_12233,N_12336);
and U12466 (N_12466,N_12383,N_12303);
xnor U12467 (N_12467,N_12338,N_12349);
nor U12468 (N_12468,N_12207,N_12204);
nand U12469 (N_12469,N_12377,N_12288);
or U12470 (N_12470,N_12289,N_12306);
nor U12471 (N_12471,N_12201,N_12375);
nor U12472 (N_12472,N_12385,N_12218);
nor U12473 (N_12473,N_12326,N_12301);
nor U12474 (N_12474,N_12353,N_12225);
nand U12475 (N_12475,N_12290,N_12308);
nand U12476 (N_12476,N_12360,N_12342);
xnor U12477 (N_12477,N_12331,N_12249);
nor U12478 (N_12478,N_12327,N_12309);
nand U12479 (N_12479,N_12313,N_12278);
nor U12480 (N_12480,N_12347,N_12226);
xor U12481 (N_12481,N_12299,N_12284);
and U12482 (N_12482,N_12259,N_12237);
nor U12483 (N_12483,N_12310,N_12254);
or U12484 (N_12484,N_12373,N_12325);
nand U12485 (N_12485,N_12243,N_12337);
nor U12486 (N_12486,N_12395,N_12221);
or U12487 (N_12487,N_12270,N_12319);
nand U12488 (N_12488,N_12333,N_12368);
nor U12489 (N_12489,N_12261,N_12231);
xnor U12490 (N_12490,N_12297,N_12384);
nor U12491 (N_12491,N_12235,N_12323);
nor U12492 (N_12492,N_12258,N_12307);
xor U12493 (N_12493,N_12344,N_12345);
xor U12494 (N_12494,N_12330,N_12269);
nor U12495 (N_12495,N_12219,N_12228);
or U12496 (N_12496,N_12317,N_12229);
and U12497 (N_12497,N_12398,N_12203);
or U12498 (N_12498,N_12271,N_12355);
or U12499 (N_12499,N_12379,N_12257);
nor U12500 (N_12500,N_12389,N_12359);
and U12501 (N_12501,N_12220,N_12260);
nor U12502 (N_12502,N_12353,N_12333);
xnor U12503 (N_12503,N_12298,N_12398);
or U12504 (N_12504,N_12380,N_12336);
nand U12505 (N_12505,N_12376,N_12300);
and U12506 (N_12506,N_12395,N_12359);
and U12507 (N_12507,N_12217,N_12295);
nor U12508 (N_12508,N_12352,N_12344);
xor U12509 (N_12509,N_12201,N_12245);
nand U12510 (N_12510,N_12202,N_12363);
nand U12511 (N_12511,N_12200,N_12359);
nand U12512 (N_12512,N_12263,N_12349);
nor U12513 (N_12513,N_12217,N_12272);
or U12514 (N_12514,N_12246,N_12211);
nor U12515 (N_12515,N_12287,N_12265);
nor U12516 (N_12516,N_12366,N_12311);
or U12517 (N_12517,N_12238,N_12381);
xor U12518 (N_12518,N_12249,N_12384);
and U12519 (N_12519,N_12226,N_12353);
nor U12520 (N_12520,N_12387,N_12231);
nor U12521 (N_12521,N_12231,N_12281);
nand U12522 (N_12522,N_12221,N_12326);
nand U12523 (N_12523,N_12210,N_12313);
nand U12524 (N_12524,N_12362,N_12237);
or U12525 (N_12525,N_12273,N_12326);
nor U12526 (N_12526,N_12307,N_12364);
nand U12527 (N_12527,N_12383,N_12367);
xnor U12528 (N_12528,N_12339,N_12325);
nand U12529 (N_12529,N_12207,N_12224);
xor U12530 (N_12530,N_12255,N_12382);
nor U12531 (N_12531,N_12378,N_12234);
nand U12532 (N_12532,N_12319,N_12350);
nor U12533 (N_12533,N_12387,N_12332);
xnor U12534 (N_12534,N_12265,N_12333);
or U12535 (N_12535,N_12278,N_12392);
xnor U12536 (N_12536,N_12273,N_12226);
xnor U12537 (N_12537,N_12301,N_12213);
and U12538 (N_12538,N_12213,N_12344);
nand U12539 (N_12539,N_12377,N_12321);
and U12540 (N_12540,N_12310,N_12398);
or U12541 (N_12541,N_12297,N_12282);
and U12542 (N_12542,N_12205,N_12349);
nand U12543 (N_12543,N_12268,N_12249);
xor U12544 (N_12544,N_12217,N_12275);
and U12545 (N_12545,N_12249,N_12343);
xnor U12546 (N_12546,N_12376,N_12297);
nand U12547 (N_12547,N_12381,N_12253);
and U12548 (N_12548,N_12278,N_12200);
or U12549 (N_12549,N_12309,N_12377);
or U12550 (N_12550,N_12322,N_12210);
and U12551 (N_12551,N_12341,N_12334);
xor U12552 (N_12552,N_12218,N_12214);
nor U12553 (N_12553,N_12228,N_12236);
or U12554 (N_12554,N_12215,N_12289);
xnor U12555 (N_12555,N_12396,N_12269);
or U12556 (N_12556,N_12296,N_12288);
nand U12557 (N_12557,N_12204,N_12264);
xor U12558 (N_12558,N_12313,N_12317);
or U12559 (N_12559,N_12324,N_12263);
nand U12560 (N_12560,N_12205,N_12249);
or U12561 (N_12561,N_12227,N_12336);
or U12562 (N_12562,N_12260,N_12234);
or U12563 (N_12563,N_12389,N_12203);
and U12564 (N_12564,N_12287,N_12373);
or U12565 (N_12565,N_12296,N_12315);
nor U12566 (N_12566,N_12257,N_12216);
and U12567 (N_12567,N_12220,N_12386);
nor U12568 (N_12568,N_12303,N_12262);
or U12569 (N_12569,N_12388,N_12253);
xnor U12570 (N_12570,N_12349,N_12260);
nand U12571 (N_12571,N_12246,N_12353);
xnor U12572 (N_12572,N_12304,N_12288);
nor U12573 (N_12573,N_12273,N_12207);
nor U12574 (N_12574,N_12342,N_12392);
nand U12575 (N_12575,N_12260,N_12369);
nand U12576 (N_12576,N_12215,N_12283);
nor U12577 (N_12577,N_12241,N_12396);
or U12578 (N_12578,N_12280,N_12395);
xor U12579 (N_12579,N_12200,N_12391);
and U12580 (N_12580,N_12395,N_12385);
xor U12581 (N_12581,N_12295,N_12300);
nand U12582 (N_12582,N_12296,N_12312);
and U12583 (N_12583,N_12309,N_12354);
and U12584 (N_12584,N_12317,N_12238);
and U12585 (N_12585,N_12355,N_12268);
nor U12586 (N_12586,N_12397,N_12352);
and U12587 (N_12587,N_12218,N_12213);
and U12588 (N_12588,N_12390,N_12244);
nand U12589 (N_12589,N_12298,N_12275);
xnor U12590 (N_12590,N_12327,N_12217);
or U12591 (N_12591,N_12300,N_12378);
xnor U12592 (N_12592,N_12273,N_12377);
nor U12593 (N_12593,N_12233,N_12318);
and U12594 (N_12594,N_12208,N_12366);
and U12595 (N_12595,N_12382,N_12236);
or U12596 (N_12596,N_12315,N_12208);
nor U12597 (N_12597,N_12271,N_12296);
nand U12598 (N_12598,N_12336,N_12246);
and U12599 (N_12599,N_12291,N_12342);
and U12600 (N_12600,N_12448,N_12567);
and U12601 (N_12601,N_12507,N_12430);
xor U12602 (N_12602,N_12520,N_12424);
xor U12603 (N_12603,N_12501,N_12511);
and U12604 (N_12604,N_12576,N_12504);
nor U12605 (N_12605,N_12418,N_12405);
nor U12606 (N_12606,N_12498,N_12499);
or U12607 (N_12607,N_12512,N_12515);
and U12608 (N_12608,N_12422,N_12591);
xnor U12609 (N_12609,N_12596,N_12492);
or U12610 (N_12610,N_12408,N_12595);
or U12611 (N_12611,N_12489,N_12525);
xnor U12612 (N_12612,N_12446,N_12407);
or U12613 (N_12613,N_12513,N_12485);
nor U12614 (N_12614,N_12552,N_12428);
or U12615 (N_12615,N_12546,N_12574);
nand U12616 (N_12616,N_12560,N_12548);
and U12617 (N_12617,N_12402,N_12510);
or U12618 (N_12618,N_12528,N_12447);
xnor U12619 (N_12619,N_12592,N_12559);
or U12620 (N_12620,N_12461,N_12438);
xor U12621 (N_12621,N_12468,N_12538);
and U12622 (N_12622,N_12414,N_12458);
nor U12623 (N_12623,N_12524,N_12579);
nor U12624 (N_12624,N_12553,N_12533);
or U12625 (N_12625,N_12565,N_12406);
xor U12626 (N_12626,N_12500,N_12415);
or U12627 (N_12627,N_12523,N_12522);
nand U12628 (N_12628,N_12566,N_12516);
nor U12629 (N_12629,N_12575,N_12420);
or U12630 (N_12630,N_12494,N_12473);
and U12631 (N_12631,N_12588,N_12488);
xor U12632 (N_12632,N_12409,N_12540);
and U12633 (N_12633,N_12587,N_12404);
nand U12634 (N_12634,N_12563,N_12439);
and U12635 (N_12635,N_12466,N_12571);
nand U12636 (N_12636,N_12583,N_12509);
nand U12637 (N_12637,N_12547,N_12435);
xor U12638 (N_12638,N_12539,N_12433);
or U12639 (N_12639,N_12578,N_12429);
and U12640 (N_12640,N_12437,N_12577);
or U12641 (N_12641,N_12454,N_12417);
xor U12642 (N_12642,N_12403,N_12467);
nand U12643 (N_12643,N_12497,N_12541);
nor U12644 (N_12644,N_12419,N_12400);
and U12645 (N_12645,N_12564,N_12464);
nand U12646 (N_12646,N_12502,N_12535);
nand U12647 (N_12647,N_12469,N_12568);
nand U12648 (N_12648,N_12544,N_12561);
or U12649 (N_12649,N_12460,N_12481);
xor U12650 (N_12650,N_12554,N_12475);
or U12651 (N_12651,N_12470,N_12532);
or U12652 (N_12652,N_12590,N_12569);
and U12653 (N_12653,N_12545,N_12580);
xnor U12654 (N_12654,N_12411,N_12531);
or U12655 (N_12655,N_12425,N_12537);
or U12656 (N_12656,N_12480,N_12455);
nand U12657 (N_12657,N_12586,N_12562);
or U12658 (N_12658,N_12457,N_12584);
or U12659 (N_12659,N_12431,N_12505);
or U12660 (N_12660,N_12490,N_12527);
nor U12661 (N_12661,N_12484,N_12413);
xnor U12662 (N_12662,N_12401,N_12599);
or U12663 (N_12663,N_12456,N_12471);
nor U12664 (N_12664,N_12436,N_12443);
xor U12665 (N_12665,N_12594,N_12508);
and U12666 (N_12666,N_12462,N_12518);
and U12667 (N_12667,N_12506,N_12449);
and U12668 (N_12668,N_12451,N_12517);
or U12669 (N_12669,N_12450,N_12534);
xor U12670 (N_12670,N_12549,N_12597);
and U12671 (N_12671,N_12542,N_12558);
nand U12672 (N_12672,N_12453,N_12444);
or U12673 (N_12673,N_12526,N_12556);
nand U12674 (N_12674,N_12474,N_12496);
or U12675 (N_12675,N_12476,N_12482);
or U12676 (N_12676,N_12589,N_12543);
and U12677 (N_12677,N_12573,N_12479);
xor U12678 (N_12678,N_12530,N_12442);
and U12679 (N_12679,N_12519,N_12426);
nor U12680 (N_12680,N_12472,N_12514);
xor U12681 (N_12681,N_12555,N_12581);
nor U12682 (N_12682,N_12410,N_12441);
nor U12683 (N_12683,N_12491,N_12421);
nor U12684 (N_12684,N_12487,N_12550);
nand U12685 (N_12685,N_12593,N_12477);
and U12686 (N_12686,N_12463,N_12423);
or U12687 (N_12687,N_12529,N_12416);
xor U12688 (N_12688,N_12459,N_12445);
nand U12689 (N_12689,N_12452,N_12440);
and U12690 (N_12690,N_12570,N_12483);
xnor U12691 (N_12691,N_12427,N_12493);
nand U12692 (N_12692,N_12598,N_12465);
nand U12693 (N_12693,N_12412,N_12557);
nor U12694 (N_12694,N_12582,N_12434);
and U12695 (N_12695,N_12495,N_12551);
nand U12696 (N_12696,N_12521,N_12503);
xor U12697 (N_12697,N_12536,N_12478);
nor U12698 (N_12698,N_12486,N_12432);
nand U12699 (N_12699,N_12585,N_12572);
nor U12700 (N_12700,N_12411,N_12529);
xnor U12701 (N_12701,N_12586,N_12488);
nand U12702 (N_12702,N_12425,N_12555);
xor U12703 (N_12703,N_12472,N_12452);
nor U12704 (N_12704,N_12514,N_12490);
or U12705 (N_12705,N_12497,N_12417);
or U12706 (N_12706,N_12592,N_12405);
and U12707 (N_12707,N_12429,N_12598);
xor U12708 (N_12708,N_12494,N_12431);
and U12709 (N_12709,N_12495,N_12502);
and U12710 (N_12710,N_12597,N_12483);
nor U12711 (N_12711,N_12403,N_12547);
or U12712 (N_12712,N_12490,N_12477);
xor U12713 (N_12713,N_12553,N_12513);
or U12714 (N_12714,N_12574,N_12592);
nor U12715 (N_12715,N_12535,N_12436);
nand U12716 (N_12716,N_12418,N_12417);
xnor U12717 (N_12717,N_12415,N_12528);
nand U12718 (N_12718,N_12445,N_12574);
and U12719 (N_12719,N_12407,N_12471);
nand U12720 (N_12720,N_12514,N_12499);
nor U12721 (N_12721,N_12580,N_12447);
or U12722 (N_12722,N_12588,N_12523);
and U12723 (N_12723,N_12437,N_12565);
nand U12724 (N_12724,N_12533,N_12556);
nor U12725 (N_12725,N_12555,N_12468);
and U12726 (N_12726,N_12473,N_12466);
and U12727 (N_12727,N_12577,N_12537);
or U12728 (N_12728,N_12581,N_12590);
nor U12729 (N_12729,N_12515,N_12543);
and U12730 (N_12730,N_12526,N_12492);
or U12731 (N_12731,N_12412,N_12547);
nor U12732 (N_12732,N_12483,N_12439);
nand U12733 (N_12733,N_12466,N_12573);
xnor U12734 (N_12734,N_12546,N_12480);
xnor U12735 (N_12735,N_12465,N_12481);
and U12736 (N_12736,N_12486,N_12425);
or U12737 (N_12737,N_12473,N_12517);
xnor U12738 (N_12738,N_12527,N_12488);
xnor U12739 (N_12739,N_12429,N_12425);
xor U12740 (N_12740,N_12528,N_12589);
or U12741 (N_12741,N_12482,N_12501);
or U12742 (N_12742,N_12533,N_12562);
nor U12743 (N_12743,N_12547,N_12551);
nand U12744 (N_12744,N_12560,N_12446);
nor U12745 (N_12745,N_12549,N_12447);
nand U12746 (N_12746,N_12581,N_12431);
and U12747 (N_12747,N_12519,N_12561);
xor U12748 (N_12748,N_12568,N_12508);
nor U12749 (N_12749,N_12414,N_12551);
nand U12750 (N_12750,N_12589,N_12447);
nand U12751 (N_12751,N_12487,N_12498);
or U12752 (N_12752,N_12542,N_12480);
xnor U12753 (N_12753,N_12552,N_12576);
nand U12754 (N_12754,N_12462,N_12549);
or U12755 (N_12755,N_12553,N_12556);
or U12756 (N_12756,N_12581,N_12580);
or U12757 (N_12757,N_12508,N_12585);
nor U12758 (N_12758,N_12507,N_12400);
nand U12759 (N_12759,N_12423,N_12480);
or U12760 (N_12760,N_12432,N_12570);
or U12761 (N_12761,N_12497,N_12585);
nor U12762 (N_12762,N_12467,N_12532);
nand U12763 (N_12763,N_12472,N_12429);
nor U12764 (N_12764,N_12482,N_12484);
xor U12765 (N_12765,N_12541,N_12428);
xor U12766 (N_12766,N_12539,N_12574);
and U12767 (N_12767,N_12586,N_12451);
nor U12768 (N_12768,N_12574,N_12560);
or U12769 (N_12769,N_12514,N_12553);
nor U12770 (N_12770,N_12482,N_12509);
or U12771 (N_12771,N_12555,N_12567);
xnor U12772 (N_12772,N_12402,N_12414);
or U12773 (N_12773,N_12405,N_12461);
or U12774 (N_12774,N_12447,N_12462);
or U12775 (N_12775,N_12525,N_12458);
nand U12776 (N_12776,N_12526,N_12532);
nor U12777 (N_12777,N_12590,N_12485);
and U12778 (N_12778,N_12427,N_12565);
or U12779 (N_12779,N_12418,N_12401);
and U12780 (N_12780,N_12463,N_12591);
or U12781 (N_12781,N_12485,N_12557);
or U12782 (N_12782,N_12536,N_12538);
and U12783 (N_12783,N_12529,N_12426);
nand U12784 (N_12784,N_12422,N_12545);
nand U12785 (N_12785,N_12553,N_12423);
and U12786 (N_12786,N_12521,N_12523);
xor U12787 (N_12787,N_12529,N_12428);
xnor U12788 (N_12788,N_12592,N_12509);
and U12789 (N_12789,N_12513,N_12569);
and U12790 (N_12790,N_12540,N_12478);
xnor U12791 (N_12791,N_12512,N_12536);
or U12792 (N_12792,N_12468,N_12449);
nor U12793 (N_12793,N_12517,N_12430);
nand U12794 (N_12794,N_12417,N_12594);
or U12795 (N_12795,N_12410,N_12484);
nor U12796 (N_12796,N_12448,N_12459);
and U12797 (N_12797,N_12420,N_12427);
nor U12798 (N_12798,N_12485,N_12470);
nor U12799 (N_12799,N_12586,N_12444);
nor U12800 (N_12800,N_12643,N_12628);
or U12801 (N_12801,N_12679,N_12722);
nand U12802 (N_12802,N_12638,N_12712);
nor U12803 (N_12803,N_12682,N_12678);
nor U12804 (N_12804,N_12691,N_12687);
nor U12805 (N_12805,N_12753,N_12680);
xnor U12806 (N_12806,N_12701,N_12721);
nor U12807 (N_12807,N_12613,N_12714);
xor U12808 (N_12808,N_12610,N_12648);
nor U12809 (N_12809,N_12767,N_12644);
xnor U12810 (N_12810,N_12667,N_12622);
and U12811 (N_12811,N_12723,N_12779);
and U12812 (N_12812,N_12602,N_12612);
and U12813 (N_12813,N_12734,N_12744);
nand U12814 (N_12814,N_12663,N_12787);
and U12815 (N_12815,N_12719,N_12651);
and U12816 (N_12816,N_12760,N_12670);
and U12817 (N_12817,N_12609,N_12674);
nand U12818 (N_12818,N_12618,N_12724);
nand U12819 (N_12819,N_12607,N_12639);
or U12820 (N_12820,N_12641,N_12659);
nand U12821 (N_12821,N_12681,N_12795);
or U12822 (N_12822,N_12605,N_12743);
nor U12823 (N_12823,N_12774,N_12632);
nor U12824 (N_12824,N_12750,N_12685);
or U12825 (N_12825,N_12739,N_12683);
nor U12826 (N_12826,N_12725,N_12693);
and U12827 (N_12827,N_12718,N_12621);
xor U12828 (N_12828,N_12730,N_12764);
or U12829 (N_12829,N_12615,N_12798);
nand U12830 (N_12830,N_12688,N_12705);
and U12831 (N_12831,N_12732,N_12709);
nor U12832 (N_12832,N_12792,N_12624);
nor U12833 (N_12833,N_12661,N_12656);
and U12834 (N_12834,N_12634,N_12799);
xnor U12835 (N_12835,N_12755,N_12617);
and U12836 (N_12836,N_12733,N_12713);
nor U12837 (N_12837,N_12700,N_12790);
and U12838 (N_12838,N_12773,N_12735);
xnor U12839 (N_12839,N_12777,N_12704);
nand U12840 (N_12840,N_12776,N_12796);
or U12841 (N_12841,N_12635,N_12740);
or U12842 (N_12842,N_12782,N_12788);
or U12843 (N_12843,N_12707,N_12649);
nand U12844 (N_12844,N_12728,N_12601);
and U12845 (N_12845,N_12671,N_12731);
nor U12846 (N_12846,N_12697,N_12762);
nor U12847 (N_12847,N_12600,N_12666);
nor U12848 (N_12848,N_12784,N_12673);
xor U12849 (N_12849,N_12620,N_12625);
and U12850 (N_12850,N_12747,N_12727);
xor U12851 (N_12851,N_12715,N_12662);
or U12852 (N_12852,N_12654,N_12603);
nor U12853 (N_12853,N_12781,N_12698);
xnor U12854 (N_12854,N_12658,N_12742);
or U12855 (N_12855,N_12637,N_12761);
nand U12856 (N_12856,N_12752,N_12789);
nor U12857 (N_12857,N_12706,N_12716);
and U12858 (N_12858,N_12636,N_12759);
xor U12859 (N_12859,N_12754,N_12769);
nor U12860 (N_12860,N_12645,N_12786);
xnor U12861 (N_12861,N_12652,N_12702);
nand U12862 (N_12862,N_12616,N_12736);
xor U12863 (N_12863,N_12686,N_12703);
and U12864 (N_12864,N_12646,N_12791);
and U12865 (N_12865,N_12692,N_12780);
and U12866 (N_12866,N_12771,N_12737);
and U12867 (N_12867,N_12751,N_12783);
xor U12868 (N_12868,N_12710,N_12749);
xor U12869 (N_12869,N_12717,N_12741);
nor U12870 (N_12870,N_12653,N_12606);
nor U12871 (N_12871,N_12756,N_12640);
nand U12872 (N_12872,N_12672,N_12675);
nor U12873 (N_12873,N_12647,N_12664);
nor U12874 (N_12874,N_12699,N_12614);
and U12875 (N_12875,N_12763,N_12657);
nor U12876 (N_12876,N_12689,N_12668);
nand U12877 (N_12877,N_12695,N_12748);
nand U12878 (N_12878,N_12768,N_12775);
and U12879 (N_12879,N_12729,N_12745);
and U12880 (N_12880,N_12694,N_12785);
nand U12881 (N_12881,N_12669,N_12757);
and U12882 (N_12882,N_12793,N_12650);
nand U12883 (N_12883,N_12772,N_12738);
nand U12884 (N_12884,N_12629,N_12711);
or U12885 (N_12885,N_12626,N_12778);
nand U12886 (N_12886,N_12794,N_12655);
nor U12887 (N_12887,N_12758,N_12676);
nand U12888 (N_12888,N_12623,N_12619);
xor U12889 (N_12889,N_12660,N_12696);
or U12890 (N_12890,N_12631,N_12665);
nor U12891 (N_12891,N_12604,N_12684);
nor U12892 (N_12892,N_12765,N_12608);
xor U12893 (N_12893,N_12746,N_12797);
or U12894 (N_12894,N_12708,N_12677);
xnor U12895 (N_12895,N_12611,N_12633);
and U12896 (N_12896,N_12627,N_12690);
xnor U12897 (N_12897,N_12770,N_12766);
nor U12898 (N_12898,N_12642,N_12726);
xnor U12899 (N_12899,N_12720,N_12630);
or U12900 (N_12900,N_12701,N_12604);
nand U12901 (N_12901,N_12796,N_12623);
nor U12902 (N_12902,N_12655,N_12705);
nand U12903 (N_12903,N_12764,N_12763);
xor U12904 (N_12904,N_12626,N_12681);
and U12905 (N_12905,N_12773,N_12627);
nor U12906 (N_12906,N_12678,N_12715);
or U12907 (N_12907,N_12682,N_12699);
or U12908 (N_12908,N_12669,N_12766);
xnor U12909 (N_12909,N_12739,N_12725);
nor U12910 (N_12910,N_12754,N_12750);
or U12911 (N_12911,N_12684,N_12707);
or U12912 (N_12912,N_12647,N_12779);
xor U12913 (N_12913,N_12795,N_12606);
nor U12914 (N_12914,N_12775,N_12674);
nand U12915 (N_12915,N_12651,N_12607);
nand U12916 (N_12916,N_12677,N_12785);
nand U12917 (N_12917,N_12729,N_12716);
xnor U12918 (N_12918,N_12655,N_12723);
nor U12919 (N_12919,N_12698,N_12644);
xnor U12920 (N_12920,N_12791,N_12788);
and U12921 (N_12921,N_12696,N_12654);
nand U12922 (N_12922,N_12694,N_12768);
nor U12923 (N_12923,N_12637,N_12785);
nor U12924 (N_12924,N_12774,N_12730);
xnor U12925 (N_12925,N_12687,N_12663);
nand U12926 (N_12926,N_12701,N_12638);
and U12927 (N_12927,N_12671,N_12795);
nor U12928 (N_12928,N_12703,N_12654);
and U12929 (N_12929,N_12778,N_12680);
xor U12930 (N_12930,N_12608,N_12757);
nand U12931 (N_12931,N_12787,N_12622);
xor U12932 (N_12932,N_12778,N_12705);
and U12933 (N_12933,N_12789,N_12609);
xnor U12934 (N_12934,N_12772,N_12741);
xor U12935 (N_12935,N_12631,N_12766);
or U12936 (N_12936,N_12714,N_12695);
xnor U12937 (N_12937,N_12725,N_12690);
and U12938 (N_12938,N_12748,N_12700);
or U12939 (N_12939,N_12748,N_12743);
and U12940 (N_12940,N_12662,N_12675);
or U12941 (N_12941,N_12650,N_12773);
and U12942 (N_12942,N_12720,N_12632);
nor U12943 (N_12943,N_12640,N_12750);
nor U12944 (N_12944,N_12738,N_12697);
and U12945 (N_12945,N_12647,N_12763);
xnor U12946 (N_12946,N_12651,N_12693);
xnor U12947 (N_12947,N_12748,N_12616);
xnor U12948 (N_12948,N_12782,N_12641);
or U12949 (N_12949,N_12602,N_12617);
or U12950 (N_12950,N_12631,N_12642);
xnor U12951 (N_12951,N_12797,N_12763);
nor U12952 (N_12952,N_12617,N_12708);
xnor U12953 (N_12953,N_12656,N_12790);
nand U12954 (N_12954,N_12619,N_12634);
nand U12955 (N_12955,N_12690,N_12762);
and U12956 (N_12956,N_12780,N_12636);
xnor U12957 (N_12957,N_12703,N_12696);
nand U12958 (N_12958,N_12693,N_12696);
nor U12959 (N_12959,N_12752,N_12688);
nor U12960 (N_12960,N_12752,N_12630);
nand U12961 (N_12961,N_12693,N_12776);
xor U12962 (N_12962,N_12701,N_12681);
xor U12963 (N_12963,N_12634,N_12723);
or U12964 (N_12964,N_12760,N_12758);
nand U12965 (N_12965,N_12624,N_12719);
or U12966 (N_12966,N_12730,N_12759);
xor U12967 (N_12967,N_12709,N_12761);
and U12968 (N_12968,N_12744,N_12600);
nor U12969 (N_12969,N_12610,N_12694);
nor U12970 (N_12970,N_12602,N_12781);
or U12971 (N_12971,N_12752,N_12613);
and U12972 (N_12972,N_12682,N_12794);
nand U12973 (N_12973,N_12798,N_12630);
nor U12974 (N_12974,N_12654,N_12681);
nor U12975 (N_12975,N_12609,N_12605);
nand U12976 (N_12976,N_12690,N_12704);
and U12977 (N_12977,N_12666,N_12776);
nand U12978 (N_12978,N_12715,N_12701);
and U12979 (N_12979,N_12760,N_12750);
nor U12980 (N_12980,N_12696,N_12671);
and U12981 (N_12981,N_12708,N_12664);
or U12982 (N_12982,N_12643,N_12646);
and U12983 (N_12983,N_12760,N_12700);
nor U12984 (N_12984,N_12706,N_12780);
and U12985 (N_12985,N_12740,N_12778);
nand U12986 (N_12986,N_12722,N_12742);
nor U12987 (N_12987,N_12654,N_12731);
and U12988 (N_12988,N_12695,N_12609);
nor U12989 (N_12989,N_12616,N_12602);
nand U12990 (N_12990,N_12601,N_12611);
nand U12991 (N_12991,N_12662,N_12604);
or U12992 (N_12992,N_12682,N_12744);
xnor U12993 (N_12993,N_12774,N_12610);
xor U12994 (N_12994,N_12705,N_12675);
or U12995 (N_12995,N_12779,N_12655);
and U12996 (N_12996,N_12667,N_12693);
and U12997 (N_12997,N_12716,N_12628);
nand U12998 (N_12998,N_12667,N_12707);
or U12999 (N_12999,N_12605,N_12734);
nor U13000 (N_13000,N_12973,N_12971);
or U13001 (N_13001,N_12994,N_12989);
or U13002 (N_13002,N_12902,N_12962);
nand U13003 (N_13003,N_12852,N_12960);
nand U13004 (N_13004,N_12829,N_12931);
nor U13005 (N_13005,N_12899,N_12945);
nand U13006 (N_13006,N_12996,N_12845);
and U13007 (N_13007,N_12863,N_12943);
nand U13008 (N_13008,N_12813,N_12929);
xor U13009 (N_13009,N_12982,N_12893);
nor U13010 (N_13010,N_12880,N_12846);
nand U13011 (N_13011,N_12867,N_12859);
xor U13012 (N_13012,N_12853,N_12938);
xor U13013 (N_13013,N_12836,N_12951);
xnor U13014 (N_13014,N_12924,N_12828);
or U13015 (N_13015,N_12808,N_12912);
and U13016 (N_13016,N_12810,N_12837);
nor U13017 (N_13017,N_12936,N_12886);
xor U13018 (N_13018,N_12838,N_12882);
or U13019 (N_13019,N_12800,N_12889);
nor U13020 (N_13020,N_12919,N_12975);
nor U13021 (N_13021,N_12986,N_12988);
and U13022 (N_13022,N_12997,N_12884);
xnor U13023 (N_13023,N_12980,N_12878);
nand U13024 (N_13024,N_12881,N_12857);
xnor U13025 (N_13025,N_12825,N_12944);
nand U13026 (N_13026,N_12850,N_12820);
nand U13027 (N_13027,N_12817,N_12869);
nor U13028 (N_13028,N_12923,N_12876);
xnor U13029 (N_13029,N_12842,N_12823);
xor U13030 (N_13030,N_12866,N_12841);
and U13031 (N_13031,N_12955,N_12830);
and U13032 (N_13032,N_12948,N_12967);
xor U13033 (N_13033,N_12819,N_12926);
xor U13034 (N_13034,N_12908,N_12978);
nand U13035 (N_13035,N_12898,N_12993);
or U13036 (N_13036,N_12833,N_12897);
nand U13037 (N_13037,N_12883,N_12934);
and U13038 (N_13038,N_12937,N_12873);
xnor U13039 (N_13039,N_12906,N_12953);
nand U13040 (N_13040,N_12966,N_12821);
nand U13041 (N_13041,N_12981,N_12921);
nand U13042 (N_13042,N_12942,N_12990);
or U13043 (N_13043,N_12887,N_12890);
xor U13044 (N_13044,N_12972,N_12987);
and U13045 (N_13045,N_12849,N_12854);
or U13046 (N_13046,N_12894,N_12965);
nor U13047 (N_13047,N_12920,N_12946);
or U13048 (N_13048,N_12822,N_12875);
xnor U13049 (N_13049,N_12957,N_12803);
nand U13050 (N_13050,N_12847,N_12985);
xor U13051 (N_13051,N_12958,N_12999);
xor U13052 (N_13052,N_12874,N_12895);
or U13053 (N_13053,N_12892,N_12861);
nor U13054 (N_13054,N_12939,N_12848);
or U13055 (N_13055,N_12824,N_12984);
xnor U13056 (N_13056,N_12806,N_12910);
and U13057 (N_13057,N_12826,N_12900);
nand U13058 (N_13058,N_12961,N_12864);
and U13059 (N_13059,N_12839,N_12932);
nand U13060 (N_13060,N_12911,N_12917);
nand U13061 (N_13061,N_12871,N_12843);
nand U13062 (N_13062,N_12969,N_12827);
or U13063 (N_13063,N_12998,N_12995);
or U13064 (N_13064,N_12840,N_12879);
or U13065 (N_13065,N_12844,N_12991);
and U13066 (N_13066,N_12968,N_12925);
and U13067 (N_13067,N_12964,N_12956);
nand U13068 (N_13068,N_12804,N_12976);
nor U13069 (N_13069,N_12927,N_12952);
and U13070 (N_13070,N_12815,N_12940);
xor U13071 (N_13071,N_12855,N_12814);
and U13072 (N_13072,N_12930,N_12891);
nor U13073 (N_13073,N_12909,N_12941);
xnor U13074 (N_13074,N_12963,N_12896);
xnor U13075 (N_13075,N_12865,N_12805);
nor U13076 (N_13076,N_12872,N_12916);
xor U13077 (N_13077,N_12905,N_12915);
xnor U13078 (N_13078,N_12888,N_12914);
xnor U13079 (N_13079,N_12834,N_12856);
xor U13080 (N_13080,N_12862,N_12933);
xnor U13081 (N_13081,N_12979,N_12904);
and U13082 (N_13082,N_12935,N_12901);
and U13083 (N_13083,N_12801,N_12885);
nor U13084 (N_13084,N_12816,N_12907);
and U13085 (N_13085,N_12835,N_12870);
xnor U13086 (N_13086,N_12811,N_12974);
nor U13087 (N_13087,N_12922,N_12860);
and U13088 (N_13088,N_12977,N_12954);
xnor U13089 (N_13089,N_12868,N_12959);
and U13090 (N_13090,N_12913,N_12903);
and U13091 (N_13091,N_12812,N_12851);
and U13092 (N_13092,N_12983,N_12950);
nand U13093 (N_13093,N_12818,N_12947);
xnor U13094 (N_13094,N_12809,N_12970);
nand U13095 (N_13095,N_12832,N_12802);
or U13096 (N_13096,N_12949,N_12831);
and U13097 (N_13097,N_12992,N_12807);
nor U13098 (N_13098,N_12928,N_12877);
nor U13099 (N_13099,N_12858,N_12918);
nor U13100 (N_13100,N_12965,N_12812);
or U13101 (N_13101,N_12927,N_12864);
or U13102 (N_13102,N_12872,N_12964);
xor U13103 (N_13103,N_12976,N_12940);
nor U13104 (N_13104,N_12984,N_12969);
or U13105 (N_13105,N_12947,N_12841);
nor U13106 (N_13106,N_12901,N_12809);
nor U13107 (N_13107,N_12886,N_12992);
and U13108 (N_13108,N_12905,N_12890);
or U13109 (N_13109,N_12858,N_12971);
nand U13110 (N_13110,N_12885,N_12872);
and U13111 (N_13111,N_12942,N_12982);
or U13112 (N_13112,N_12973,N_12905);
or U13113 (N_13113,N_12835,N_12907);
xnor U13114 (N_13114,N_12952,N_12816);
nor U13115 (N_13115,N_12867,N_12822);
nor U13116 (N_13116,N_12948,N_12937);
nand U13117 (N_13117,N_12973,N_12800);
and U13118 (N_13118,N_12933,N_12821);
and U13119 (N_13119,N_12966,N_12853);
nand U13120 (N_13120,N_12996,N_12901);
nor U13121 (N_13121,N_12827,N_12816);
nor U13122 (N_13122,N_12849,N_12879);
xnor U13123 (N_13123,N_12937,N_12817);
nor U13124 (N_13124,N_12974,N_12839);
nor U13125 (N_13125,N_12890,N_12926);
or U13126 (N_13126,N_12899,N_12901);
nand U13127 (N_13127,N_12948,N_12856);
and U13128 (N_13128,N_12866,N_12817);
nor U13129 (N_13129,N_12938,N_12851);
nor U13130 (N_13130,N_12910,N_12853);
nor U13131 (N_13131,N_12859,N_12919);
xnor U13132 (N_13132,N_12835,N_12844);
xor U13133 (N_13133,N_12833,N_12866);
nor U13134 (N_13134,N_12859,N_12945);
nand U13135 (N_13135,N_12912,N_12822);
nor U13136 (N_13136,N_12850,N_12974);
xnor U13137 (N_13137,N_12960,N_12944);
nand U13138 (N_13138,N_12802,N_12941);
xnor U13139 (N_13139,N_12954,N_12807);
nand U13140 (N_13140,N_12940,N_12910);
and U13141 (N_13141,N_12988,N_12831);
or U13142 (N_13142,N_12877,N_12876);
or U13143 (N_13143,N_12813,N_12900);
xor U13144 (N_13144,N_12921,N_12900);
nor U13145 (N_13145,N_12956,N_12884);
xnor U13146 (N_13146,N_12886,N_12970);
nand U13147 (N_13147,N_12907,N_12927);
nand U13148 (N_13148,N_12802,N_12800);
nand U13149 (N_13149,N_12876,N_12861);
nand U13150 (N_13150,N_12844,N_12955);
xnor U13151 (N_13151,N_12810,N_12816);
nand U13152 (N_13152,N_12980,N_12963);
xnor U13153 (N_13153,N_12805,N_12929);
and U13154 (N_13154,N_12862,N_12937);
xnor U13155 (N_13155,N_12903,N_12862);
xor U13156 (N_13156,N_12951,N_12949);
or U13157 (N_13157,N_12940,N_12838);
xor U13158 (N_13158,N_12800,N_12957);
and U13159 (N_13159,N_12872,N_12912);
nand U13160 (N_13160,N_12827,N_12804);
and U13161 (N_13161,N_12925,N_12808);
and U13162 (N_13162,N_12874,N_12893);
nand U13163 (N_13163,N_12846,N_12967);
nand U13164 (N_13164,N_12902,N_12823);
and U13165 (N_13165,N_12958,N_12921);
or U13166 (N_13166,N_12900,N_12992);
xnor U13167 (N_13167,N_12983,N_12900);
nand U13168 (N_13168,N_12868,N_12982);
nor U13169 (N_13169,N_12870,N_12977);
nor U13170 (N_13170,N_12975,N_12936);
xnor U13171 (N_13171,N_12921,N_12980);
nand U13172 (N_13172,N_12998,N_12887);
nor U13173 (N_13173,N_12994,N_12995);
or U13174 (N_13174,N_12889,N_12903);
nor U13175 (N_13175,N_12845,N_12901);
or U13176 (N_13176,N_12854,N_12869);
nand U13177 (N_13177,N_12986,N_12820);
xnor U13178 (N_13178,N_12881,N_12951);
nor U13179 (N_13179,N_12911,N_12936);
and U13180 (N_13180,N_12946,N_12994);
xor U13181 (N_13181,N_12972,N_12924);
or U13182 (N_13182,N_12937,N_12951);
and U13183 (N_13183,N_12838,N_12878);
xnor U13184 (N_13184,N_12810,N_12951);
and U13185 (N_13185,N_12939,N_12962);
xor U13186 (N_13186,N_12904,N_12935);
nor U13187 (N_13187,N_12978,N_12927);
xor U13188 (N_13188,N_12884,N_12974);
or U13189 (N_13189,N_12846,N_12903);
and U13190 (N_13190,N_12871,N_12904);
or U13191 (N_13191,N_12872,N_12835);
xnor U13192 (N_13192,N_12865,N_12947);
or U13193 (N_13193,N_12965,N_12900);
nor U13194 (N_13194,N_12955,N_12841);
or U13195 (N_13195,N_12849,N_12984);
nand U13196 (N_13196,N_12953,N_12814);
and U13197 (N_13197,N_12887,N_12822);
nand U13198 (N_13198,N_12806,N_12850);
nor U13199 (N_13199,N_12886,N_12985);
nand U13200 (N_13200,N_13090,N_13048);
or U13201 (N_13201,N_13105,N_13072);
and U13202 (N_13202,N_13147,N_13036);
and U13203 (N_13203,N_13151,N_13061);
nor U13204 (N_13204,N_13180,N_13089);
nand U13205 (N_13205,N_13120,N_13141);
nor U13206 (N_13206,N_13191,N_13149);
nor U13207 (N_13207,N_13008,N_13116);
nor U13208 (N_13208,N_13161,N_13107);
nor U13209 (N_13209,N_13115,N_13169);
nor U13210 (N_13210,N_13199,N_13137);
nand U13211 (N_13211,N_13065,N_13179);
nor U13212 (N_13212,N_13031,N_13014);
nor U13213 (N_13213,N_13013,N_13084);
or U13214 (N_13214,N_13052,N_13138);
and U13215 (N_13215,N_13101,N_13133);
or U13216 (N_13216,N_13187,N_13119);
nand U13217 (N_13217,N_13175,N_13092);
xnor U13218 (N_13218,N_13177,N_13170);
or U13219 (N_13219,N_13155,N_13011);
or U13220 (N_13220,N_13136,N_13094);
xor U13221 (N_13221,N_13194,N_13005);
and U13222 (N_13222,N_13073,N_13025);
or U13223 (N_13223,N_13123,N_13131);
nor U13224 (N_13224,N_13068,N_13142);
nand U13225 (N_13225,N_13009,N_13188);
nor U13226 (N_13226,N_13148,N_13165);
or U13227 (N_13227,N_13003,N_13000);
or U13228 (N_13228,N_13095,N_13108);
nor U13229 (N_13229,N_13016,N_13004);
xnor U13230 (N_13230,N_13195,N_13171);
nor U13231 (N_13231,N_13069,N_13040);
or U13232 (N_13232,N_13166,N_13096);
xor U13233 (N_13233,N_13196,N_13060);
and U13234 (N_13234,N_13128,N_13046);
nand U13235 (N_13235,N_13109,N_13198);
and U13236 (N_13236,N_13197,N_13099);
nor U13237 (N_13237,N_13082,N_13150);
nor U13238 (N_13238,N_13030,N_13021);
nand U13239 (N_13239,N_13085,N_13033);
nor U13240 (N_13240,N_13132,N_13174);
nand U13241 (N_13241,N_13192,N_13055);
and U13242 (N_13242,N_13158,N_13054);
nor U13243 (N_13243,N_13006,N_13043);
xnor U13244 (N_13244,N_13076,N_13135);
and U13245 (N_13245,N_13044,N_13182);
nor U13246 (N_13246,N_13130,N_13172);
xor U13247 (N_13247,N_13156,N_13049);
and U13248 (N_13248,N_13058,N_13057);
nor U13249 (N_13249,N_13051,N_13117);
nor U13250 (N_13250,N_13080,N_13122);
nor U13251 (N_13251,N_13042,N_13088);
and U13252 (N_13252,N_13034,N_13078);
nand U13253 (N_13253,N_13097,N_13086);
nand U13254 (N_13254,N_13007,N_13178);
or U13255 (N_13255,N_13125,N_13140);
and U13256 (N_13256,N_13162,N_13056);
nand U13257 (N_13257,N_13159,N_13062);
or U13258 (N_13258,N_13127,N_13081);
nand U13259 (N_13259,N_13083,N_13045);
and U13260 (N_13260,N_13121,N_13015);
or U13261 (N_13261,N_13001,N_13067);
nand U13262 (N_13262,N_13038,N_13037);
or U13263 (N_13263,N_13113,N_13039);
or U13264 (N_13264,N_13185,N_13103);
nand U13265 (N_13265,N_13024,N_13020);
and U13266 (N_13266,N_13077,N_13124);
nor U13267 (N_13267,N_13163,N_13026);
and U13268 (N_13268,N_13129,N_13181);
xor U13269 (N_13269,N_13167,N_13193);
and U13270 (N_13270,N_13144,N_13053);
xnor U13271 (N_13271,N_13164,N_13173);
xnor U13272 (N_13272,N_13093,N_13134);
and U13273 (N_13273,N_13059,N_13102);
or U13274 (N_13274,N_13074,N_13010);
nand U13275 (N_13275,N_13063,N_13064);
nor U13276 (N_13276,N_13087,N_13114);
nand U13277 (N_13277,N_13027,N_13098);
nor U13278 (N_13278,N_13111,N_13079);
or U13279 (N_13279,N_13028,N_13153);
or U13280 (N_13280,N_13152,N_13168);
and U13281 (N_13281,N_13126,N_13112);
xor U13282 (N_13282,N_13143,N_13154);
and U13283 (N_13283,N_13183,N_13091);
xor U13284 (N_13284,N_13184,N_13106);
nand U13285 (N_13285,N_13189,N_13023);
or U13286 (N_13286,N_13019,N_13070);
nor U13287 (N_13287,N_13190,N_13066);
and U13288 (N_13288,N_13035,N_13139);
xor U13289 (N_13289,N_13146,N_13032);
nor U13290 (N_13290,N_13186,N_13018);
or U13291 (N_13291,N_13012,N_13100);
or U13292 (N_13292,N_13047,N_13050);
nor U13293 (N_13293,N_13017,N_13176);
or U13294 (N_13294,N_13160,N_13118);
and U13295 (N_13295,N_13110,N_13075);
or U13296 (N_13296,N_13071,N_13022);
and U13297 (N_13297,N_13157,N_13104);
or U13298 (N_13298,N_13041,N_13029);
xnor U13299 (N_13299,N_13002,N_13145);
xor U13300 (N_13300,N_13126,N_13024);
and U13301 (N_13301,N_13177,N_13171);
and U13302 (N_13302,N_13164,N_13002);
nand U13303 (N_13303,N_13170,N_13061);
and U13304 (N_13304,N_13148,N_13102);
nand U13305 (N_13305,N_13013,N_13046);
nor U13306 (N_13306,N_13068,N_13031);
nor U13307 (N_13307,N_13091,N_13105);
nor U13308 (N_13308,N_13139,N_13042);
or U13309 (N_13309,N_13090,N_13116);
nor U13310 (N_13310,N_13187,N_13194);
xor U13311 (N_13311,N_13176,N_13134);
nand U13312 (N_13312,N_13009,N_13181);
nor U13313 (N_13313,N_13122,N_13025);
or U13314 (N_13314,N_13102,N_13006);
nor U13315 (N_13315,N_13034,N_13106);
or U13316 (N_13316,N_13026,N_13043);
or U13317 (N_13317,N_13167,N_13073);
nor U13318 (N_13318,N_13103,N_13095);
xnor U13319 (N_13319,N_13047,N_13144);
nand U13320 (N_13320,N_13036,N_13122);
nand U13321 (N_13321,N_13073,N_13061);
or U13322 (N_13322,N_13065,N_13108);
or U13323 (N_13323,N_13037,N_13029);
nand U13324 (N_13324,N_13051,N_13062);
nor U13325 (N_13325,N_13125,N_13088);
nand U13326 (N_13326,N_13060,N_13088);
or U13327 (N_13327,N_13197,N_13179);
xnor U13328 (N_13328,N_13134,N_13174);
nor U13329 (N_13329,N_13166,N_13165);
or U13330 (N_13330,N_13082,N_13186);
xnor U13331 (N_13331,N_13007,N_13124);
nand U13332 (N_13332,N_13023,N_13016);
and U13333 (N_13333,N_13053,N_13074);
xor U13334 (N_13334,N_13093,N_13148);
and U13335 (N_13335,N_13021,N_13138);
nand U13336 (N_13336,N_13045,N_13128);
and U13337 (N_13337,N_13097,N_13128);
or U13338 (N_13338,N_13118,N_13012);
or U13339 (N_13339,N_13127,N_13131);
or U13340 (N_13340,N_13137,N_13035);
xor U13341 (N_13341,N_13062,N_13052);
nand U13342 (N_13342,N_13038,N_13197);
or U13343 (N_13343,N_13123,N_13078);
xnor U13344 (N_13344,N_13165,N_13080);
and U13345 (N_13345,N_13188,N_13061);
or U13346 (N_13346,N_13133,N_13141);
or U13347 (N_13347,N_13131,N_13038);
and U13348 (N_13348,N_13110,N_13198);
or U13349 (N_13349,N_13052,N_13110);
and U13350 (N_13350,N_13084,N_13055);
and U13351 (N_13351,N_13108,N_13139);
or U13352 (N_13352,N_13122,N_13084);
nand U13353 (N_13353,N_13100,N_13150);
nor U13354 (N_13354,N_13090,N_13077);
and U13355 (N_13355,N_13001,N_13160);
nand U13356 (N_13356,N_13054,N_13170);
nand U13357 (N_13357,N_13054,N_13144);
nand U13358 (N_13358,N_13127,N_13109);
nand U13359 (N_13359,N_13052,N_13121);
xnor U13360 (N_13360,N_13015,N_13051);
and U13361 (N_13361,N_13195,N_13169);
xor U13362 (N_13362,N_13052,N_13177);
or U13363 (N_13363,N_13014,N_13115);
or U13364 (N_13364,N_13107,N_13077);
and U13365 (N_13365,N_13183,N_13080);
or U13366 (N_13366,N_13094,N_13123);
nand U13367 (N_13367,N_13044,N_13095);
or U13368 (N_13368,N_13109,N_13097);
or U13369 (N_13369,N_13098,N_13019);
nor U13370 (N_13370,N_13192,N_13003);
xnor U13371 (N_13371,N_13107,N_13153);
nand U13372 (N_13372,N_13045,N_13009);
xnor U13373 (N_13373,N_13070,N_13135);
xnor U13374 (N_13374,N_13129,N_13199);
nand U13375 (N_13375,N_13102,N_13176);
and U13376 (N_13376,N_13038,N_13105);
or U13377 (N_13377,N_13073,N_13175);
xnor U13378 (N_13378,N_13122,N_13134);
or U13379 (N_13379,N_13184,N_13129);
xor U13380 (N_13380,N_13199,N_13190);
nand U13381 (N_13381,N_13159,N_13030);
or U13382 (N_13382,N_13090,N_13120);
nand U13383 (N_13383,N_13039,N_13159);
and U13384 (N_13384,N_13063,N_13074);
xnor U13385 (N_13385,N_13011,N_13104);
or U13386 (N_13386,N_13058,N_13025);
nor U13387 (N_13387,N_13045,N_13179);
nor U13388 (N_13388,N_13097,N_13113);
xor U13389 (N_13389,N_13094,N_13129);
xor U13390 (N_13390,N_13067,N_13139);
or U13391 (N_13391,N_13183,N_13094);
or U13392 (N_13392,N_13055,N_13195);
nor U13393 (N_13393,N_13037,N_13048);
xor U13394 (N_13394,N_13037,N_13171);
nand U13395 (N_13395,N_13195,N_13087);
xor U13396 (N_13396,N_13047,N_13140);
nor U13397 (N_13397,N_13021,N_13063);
xor U13398 (N_13398,N_13095,N_13005);
nand U13399 (N_13399,N_13004,N_13009);
nor U13400 (N_13400,N_13202,N_13379);
xor U13401 (N_13401,N_13330,N_13316);
xor U13402 (N_13402,N_13246,N_13230);
or U13403 (N_13403,N_13301,N_13238);
xor U13404 (N_13404,N_13315,N_13224);
or U13405 (N_13405,N_13317,N_13253);
xor U13406 (N_13406,N_13241,N_13210);
or U13407 (N_13407,N_13290,N_13376);
or U13408 (N_13408,N_13276,N_13320);
or U13409 (N_13409,N_13300,N_13394);
nand U13410 (N_13410,N_13386,N_13204);
nor U13411 (N_13411,N_13322,N_13321);
nor U13412 (N_13412,N_13207,N_13332);
xnor U13413 (N_13413,N_13351,N_13274);
or U13414 (N_13414,N_13272,N_13213);
nand U13415 (N_13415,N_13356,N_13341);
and U13416 (N_13416,N_13363,N_13340);
nand U13417 (N_13417,N_13364,N_13242);
xnor U13418 (N_13418,N_13333,N_13236);
or U13419 (N_13419,N_13380,N_13319);
or U13420 (N_13420,N_13294,N_13299);
nor U13421 (N_13421,N_13265,N_13293);
and U13422 (N_13422,N_13292,N_13339);
nand U13423 (N_13423,N_13233,N_13302);
and U13424 (N_13424,N_13389,N_13390);
or U13425 (N_13425,N_13261,N_13347);
or U13426 (N_13426,N_13370,N_13227);
nor U13427 (N_13427,N_13212,N_13397);
or U13428 (N_13428,N_13229,N_13280);
and U13429 (N_13429,N_13270,N_13251);
or U13430 (N_13430,N_13239,N_13252);
and U13431 (N_13431,N_13247,N_13279);
nand U13432 (N_13432,N_13346,N_13203);
nand U13433 (N_13433,N_13295,N_13304);
and U13434 (N_13434,N_13361,N_13217);
xnor U13435 (N_13435,N_13255,N_13352);
xnor U13436 (N_13436,N_13374,N_13232);
nand U13437 (N_13437,N_13355,N_13254);
nand U13438 (N_13438,N_13256,N_13214);
and U13439 (N_13439,N_13353,N_13263);
and U13440 (N_13440,N_13296,N_13314);
xor U13441 (N_13441,N_13220,N_13209);
and U13442 (N_13442,N_13358,N_13381);
and U13443 (N_13443,N_13298,N_13206);
or U13444 (N_13444,N_13336,N_13282);
xnor U13445 (N_13445,N_13329,N_13271);
nand U13446 (N_13446,N_13323,N_13366);
or U13447 (N_13447,N_13273,N_13237);
or U13448 (N_13448,N_13369,N_13283);
nor U13449 (N_13449,N_13312,N_13367);
or U13450 (N_13450,N_13342,N_13303);
or U13451 (N_13451,N_13226,N_13219);
nor U13452 (N_13452,N_13215,N_13291);
xnor U13453 (N_13453,N_13331,N_13396);
nor U13454 (N_13454,N_13275,N_13200);
or U13455 (N_13455,N_13338,N_13259);
nor U13456 (N_13456,N_13343,N_13344);
and U13457 (N_13457,N_13308,N_13222);
xnor U13458 (N_13458,N_13260,N_13393);
or U13459 (N_13459,N_13334,N_13399);
nor U13460 (N_13460,N_13234,N_13350);
nor U13461 (N_13461,N_13335,N_13371);
or U13462 (N_13462,N_13245,N_13244);
nor U13463 (N_13463,N_13231,N_13391);
xnor U13464 (N_13464,N_13277,N_13348);
nand U13465 (N_13465,N_13310,N_13377);
nor U13466 (N_13466,N_13359,N_13362);
nand U13467 (N_13467,N_13306,N_13266);
or U13468 (N_13468,N_13327,N_13228);
xor U13469 (N_13469,N_13357,N_13235);
nor U13470 (N_13470,N_13278,N_13385);
and U13471 (N_13471,N_13268,N_13287);
xor U13472 (N_13472,N_13267,N_13387);
nand U13473 (N_13473,N_13269,N_13262);
nand U13474 (N_13474,N_13375,N_13281);
or U13475 (N_13475,N_13284,N_13240);
nor U13476 (N_13476,N_13345,N_13208);
nor U13477 (N_13477,N_13249,N_13326);
nand U13478 (N_13478,N_13305,N_13392);
and U13479 (N_13479,N_13373,N_13257);
nand U13480 (N_13480,N_13288,N_13365);
nor U13481 (N_13481,N_13285,N_13307);
and U13482 (N_13482,N_13328,N_13248);
nand U13483 (N_13483,N_13324,N_13223);
nor U13484 (N_13484,N_13383,N_13395);
nor U13485 (N_13485,N_13218,N_13258);
xnor U13486 (N_13486,N_13354,N_13250);
or U13487 (N_13487,N_13216,N_13205);
xnor U13488 (N_13488,N_13372,N_13388);
nand U13489 (N_13489,N_13360,N_13382);
and U13490 (N_13490,N_13309,N_13289);
nor U13491 (N_13491,N_13243,N_13297);
and U13492 (N_13492,N_13286,N_13211);
or U13493 (N_13493,N_13201,N_13398);
or U13494 (N_13494,N_13311,N_13264);
or U13495 (N_13495,N_13368,N_13349);
or U13496 (N_13496,N_13225,N_13318);
and U13497 (N_13497,N_13313,N_13221);
xor U13498 (N_13498,N_13337,N_13378);
or U13499 (N_13499,N_13325,N_13384);
and U13500 (N_13500,N_13255,N_13240);
nand U13501 (N_13501,N_13311,N_13352);
xnor U13502 (N_13502,N_13297,N_13372);
and U13503 (N_13503,N_13365,N_13234);
xor U13504 (N_13504,N_13392,N_13310);
or U13505 (N_13505,N_13357,N_13391);
nor U13506 (N_13506,N_13341,N_13311);
or U13507 (N_13507,N_13359,N_13314);
nor U13508 (N_13508,N_13302,N_13393);
or U13509 (N_13509,N_13282,N_13225);
xor U13510 (N_13510,N_13312,N_13281);
or U13511 (N_13511,N_13222,N_13274);
nor U13512 (N_13512,N_13207,N_13367);
and U13513 (N_13513,N_13255,N_13211);
nor U13514 (N_13514,N_13353,N_13262);
or U13515 (N_13515,N_13212,N_13317);
nand U13516 (N_13516,N_13341,N_13308);
and U13517 (N_13517,N_13320,N_13258);
nor U13518 (N_13518,N_13378,N_13343);
or U13519 (N_13519,N_13238,N_13231);
nor U13520 (N_13520,N_13279,N_13283);
or U13521 (N_13521,N_13257,N_13308);
or U13522 (N_13522,N_13342,N_13326);
and U13523 (N_13523,N_13360,N_13356);
nand U13524 (N_13524,N_13261,N_13318);
nor U13525 (N_13525,N_13270,N_13240);
and U13526 (N_13526,N_13262,N_13361);
nor U13527 (N_13527,N_13216,N_13249);
nand U13528 (N_13528,N_13263,N_13347);
nor U13529 (N_13529,N_13349,N_13243);
xnor U13530 (N_13530,N_13392,N_13341);
nand U13531 (N_13531,N_13228,N_13364);
nor U13532 (N_13532,N_13369,N_13270);
and U13533 (N_13533,N_13366,N_13337);
nor U13534 (N_13534,N_13206,N_13237);
or U13535 (N_13535,N_13207,N_13250);
nand U13536 (N_13536,N_13366,N_13296);
or U13537 (N_13537,N_13366,N_13305);
nand U13538 (N_13538,N_13278,N_13295);
and U13539 (N_13539,N_13203,N_13328);
nor U13540 (N_13540,N_13350,N_13295);
or U13541 (N_13541,N_13232,N_13334);
nor U13542 (N_13542,N_13382,N_13324);
nor U13543 (N_13543,N_13368,N_13281);
and U13544 (N_13544,N_13263,N_13342);
xor U13545 (N_13545,N_13251,N_13207);
nor U13546 (N_13546,N_13223,N_13289);
or U13547 (N_13547,N_13314,N_13238);
nand U13548 (N_13548,N_13279,N_13230);
and U13549 (N_13549,N_13357,N_13373);
xnor U13550 (N_13550,N_13361,N_13365);
nor U13551 (N_13551,N_13224,N_13233);
xnor U13552 (N_13552,N_13230,N_13330);
nor U13553 (N_13553,N_13278,N_13299);
xnor U13554 (N_13554,N_13385,N_13398);
nand U13555 (N_13555,N_13214,N_13378);
and U13556 (N_13556,N_13351,N_13361);
or U13557 (N_13557,N_13358,N_13317);
and U13558 (N_13558,N_13380,N_13348);
nor U13559 (N_13559,N_13305,N_13313);
and U13560 (N_13560,N_13290,N_13330);
xnor U13561 (N_13561,N_13241,N_13343);
and U13562 (N_13562,N_13261,N_13277);
nand U13563 (N_13563,N_13355,N_13267);
nor U13564 (N_13564,N_13252,N_13315);
nor U13565 (N_13565,N_13300,N_13217);
nor U13566 (N_13566,N_13291,N_13240);
or U13567 (N_13567,N_13337,N_13232);
and U13568 (N_13568,N_13249,N_13337);
and U13569 (N_13569,N_13380,N_13351);
nor U13570 (N_13570,N_13229,N_13245);
xnor U13571 (N_13571,N_13384,N_13204);
nand U13572 (N_13572,N_13364,N_13353);
or U13573 (N_13573,N_13288,N_13324);
nor U13574 (N_13574,N_13343,N_13293);
or U13575 (N_13575,N_13213,N_13211);
nand U13576 (N_13576,N_13388,N_13379);
xor U13577 (N_13577,N_13346,N_13231);
xnor U13578 (N_13578,N_13370,N_13259);
and U13579 (N_13579,N_13293,N_13213);
or U13580 (N_13580,N_13372,N_13327);
or U13581 (N_13581,N_13293,N_13376);
nand U13582 (N_13582,N_13276,N_13328);
or U13583 (N_13583,N_13220,N_13358);
xnor U13584 (N_13584,N_13254,N_13326);
or U13585 (N_13585,N_13309,N_13221);
or U13586 (N_13586,N_13320,N_13375);
and U13587 (N_13587,N_13258,N_13393);
nor U13588 (N_13588,N_13293,N_13379);
xor U13589 (N_13589,N_13331,N_13343);
and U13590 (N_13590,N_13347,N_13363);
nand U13591 (N_13591,N_13365,N_13289);
nor U13592 (N_13592,N_13384,N_13375);
xnor U13593 (N_13593,N_13241,N_13363);
or U13594 (N_13594,N_13308,N_13253);
nor U13595 (N_13595,N_13368,N_13370);
nor U13596 (N_13596,N_13229,N_13320);
xnor U13597 (N_13597,N_13319,N_13337);
xor U13598 (N_13598,N_13272,N_13381);
nand U13599 (N_13599,N_13260,N_13205);
nand U13600 (N_13600,N_13424,N_13490);
and U13601 (N_13601,N_13489,N_13583);
nand U13602 (N_13602,N_13546,N_13476);
nor U13603 (N_13603,N_13582,N_13415);
or U13604 (N_13604,N_13455,N_13511);
or U13605 (N_13605,N_13519,N_13543);
nor U13606 (N_13606,N_13510,N_13497);
nor U13607 (N_13607,N_13515,N_13418);
xor U13608 (N_13608,N_13575,N_13469);
and U13609 (N_13609,N_13570,N_13553);
and U13610 (N_13610,N_13462,N_13531);
nor U13611 (N_13611,N_13473,N_13590);
xnor U13612 (N_13612,N_13508,N_13404);
and U13613 (N_13613,N_13450,N_13485);
or U13614 (N_13614,N_13592,N_13410);
nor U13615 (N_13615,N_13502,N_13571);
or U13616 (N_13616,N_13514,N_13576);
xor U13617 (N_13617,N_13427,N_13506);
or U13618 (N_13618,N_13503,N_13523);
nor U13619 (N_13619,N_13589,N_13573);
nor U13620 (N_13620,N_13527,N_13417);
nor U13621 (N_13621,N_13456,N_13559);
and U13622 (N_13622,N_13438,N_13412);
or U13623 (N_13623,N_13465,N_13414);
nor U13624 (N_13624,N_13593,N_13549);
or U13625 (N_13625,N_13529,N_13596);
xnor U13626 (N_13626,N_13585,N_13588);
nand U13627 (N_13627,N_13597,N_13433);
nor U13628 (N_13628,N_13586,N_13499);
nand U13629 (N_13629,N_13464,N_13406);
and U13630 (N_13630,N_13480,N_13505);
and U13631 (N_13631,N_13548,N_13447);
xnor U13632 (N_13632,N_13555,N_13594);
or U13633 (N_13633,N_13496,N_13537);
and U13634 (N_13634,N_13554,N_13558);
and U13635 (N_13635,N_13491,N_13532);
and U13636 (N_13636,N_13451,N_13401);
and U13637 (N_13637,N_13560,N_13440);
and U13638 (N_13638,N_13521,N_13441);
or U13639 (N_13639,N_13405,N_13507);
xnor U13640 (N_13640,N_13478,N_13439);
xor U13641 (N_13641,N_13577,N_13458);
nor U13642 (N_13642,N_13487,N_13423);
nand U13643 (N_13643,N_13483,N_13477);
nor U13644 (N_13644,N_13518,N_13525);
or U13645 (N_13645,N_13429,N_13443);
xor U13646 (N_13646,N_13470,N_13421);
or U13647 (N_13647,N_13509,N_13461);
nand U13648 (N_13648,N_13472,N_13547);
nor U13649 (N_13649,N_13512,N_13460);
xor U13650 (N_13650,N_13492,N_13598);
and U13651 (N_13651,N_13453,N_13430);
or U13652 (N_13652,N_13516,N_13540);
or U13653 (N_13653,N_13449,N_13479);
xor U13654 (N_13654,N_13530,N_13474);
nand U13655 (N_13655,N_13495,N_13488);
xor U13656 (N_13656,N_13566,N_13467);
and U13657 (N_13657,N_13431,N_13534);
or U13658 (N_13658,N_13556,N_13428);
nand U13659 (N_13659,N_13434,N_13498);
and U13660 (N_13660,N_13599,N_13435);
nor U13661 (N_13661,N_13578,N_13402);
nand U13662 (N_13662,N_13539,N_13426);
nor U13663 (N_13663,N_13457,N_13501);
nand U13664 (N_13664,N_13550,N_13587);
or U13665 (N_13665,N_13463,N_13454);
and U13666 (N_13666,N_13482,N_13408);
or U13667 (N_13667,N_13533,N_13595);
nor U13668 (N_13668,N_13562,N_13494);
nor U13669 (N_13669,N_13538,N_13544);
xnor U13670 (N_13670,N_13568,N_13572);
and U13671 (N_13671,N_13513,N_13471);
nand U13672 (N_13672,N_13484,N_13584);
and U13673 (N_13673,N_13535,N_13557);
nor U13674 (N_13674,N_13448,N_13520);
nor U13675 (N_13675,N_13569,N_13437);
nor U13676 (N_13676,N_13436,N_13403);
or U13677 (N_13677,N_13504,N_13591);
nor U13678 (N_13678,N_13545,N_13445);
or U13679 (N_13679,N_13542,N_13574);
xor U13680 (N_13680,N_13442,N_13552);
or U13681 (N_13681,N_13522,N_13416);
xnor U13682 (N_13682,N_13486,N_13452);
nand U13683 (N_13683,N_13468,N_13409);
and U13684 (N_13684,N_13400,N_13526);
xnor U13685 (N_13685,N_13580,N_13407);
nand U13686 (N_13686,N_13565,N_13551);
nand U13687 (N_13687,N_13444,N_13564);
nor U13688 (N_13688,N_13422,N_13432);
nand U13689 (N_13689,N_13536,N_13493);
nand U13690 (N_13690,N_13517,N_13459);
nor U13691 (N_13691,N_13563,N_13524);
nor U13692 (N_13692,N_13413,N_13481);
nor U13693 (N_13693,N_13579,N_13475);
xnor U13694 (N_13694,N_13581,N_13411);
nand U13695 (N_13695,N_13567,N_13541);
xnor U13696 (N_13696,N_13466,N_13419);
nor U13697 (N_13697,N_13561,N_13420);
xor U13698 (N_13698,N_13500,N_13446);
xnor U13699 (N_13699,N_13425,N_13528);
nor U13700 (N_13700,N_13496,N_13587);
nor U13701 (N_13701,N_13591,N_13425);
nor U13702 (N_13702,N_13553,N_13442);
or U13703 (N_13703,N_13545,N_13441);
or U13704 (N_13704,N_13515,N_13483);
nand U13705 (N_13705,N_13475,N_13539);
or U13706 (N_13706,N_13455,N_13512);
or U13707 (N_13707,N_13580,N_13551);
nand U13708 (N_13708,N_13562,N_13595);
and U13709 (N_13709,N_13445,N_13584);
xnor U13710 (N_13710,N_13542,N_13595);
nor U13711 (N_13711,N_13466,N_13449);
nor U13712 (N_13712,N_13409,N_13596);
or U13713 (N_13713,N_13547,N_13408);
or U13714 (N_13714,N_13541,N_13492);
or U13715 (N_13715,N_13485,N_13520);
xnor U13716 (N_13716,N_13452,N_13463);
nor U13717 (N_13717,N_13559,N_13536);
or U13718 (N_13718,N_13440,N_13512);
or U13719 (N_13719,N_13421,N_13503);
nand U13720 (N_13720,N_13487,N_13448);
and U13721 (N_13721,N_13533,N_13555);
xnor U13722 (N_13722,N_13532,N_13473);
and U13723 (N_13723,N_13530,N_13488);
and U13724 (N_13724,N_13493,N_13450);
nand U13725 (N_13725,N_13558,N_13470);
nand U13726 (N_13726,N_13478,N_13595);
nor U13727 (N_13727,N_13497,N_13519);
or U13728 (N_13728,N_13591,N_13464);
nand U13729 (N_13729,N_13450,N_13580);
xnor U13730 (N_13730,N_13589,N_13519);
nand U13731 (N_13731,N_13424,N_13446);
or U13732 (N_13732,N_13586,N_13597);
nand U13733 (N_13733,N_13558,N_13450);
nand U13734 (N_13734,N_13491,N_13489);
and U13735 (N_13735,N_13521,N_13443);
nor U13736 (N_13736,N_13460,N_13435);
xnor U13737 (N_13737,N_13570,N_13551);
xnor U13738 (N_13738,N_13474,N_13599);
xor U13739 (N_13739,N_13558,N_13552);
xor U13740 (N_13740,N_13546,N_13559);
or U13741 (N_13741,N_13431,N_13531);
and U13742 (N_13742,N_13475,N_13573);
or U13743 (N_13743,N_13568,N_13520);
xor U13744 (N_13744,N_13405,N_13586);
or U13745 (N_13745,N_13587,N_13532);
xnor U13746 (N_13746,N_13509,N_13468);
nor U13747 (N_13747,N_13544,N_13414);
and U13748 (N_13748,N_13432,N_13588);
or U13749 (N_13749,N_13454,N_13571);
nor U13750 (N_13750,N_13472,N_13402);
nor U13751 (N_13751,N_13511,N_13477);
nor U13752 (N_13752,N_13448,N_13485);
nand U13753 (N_13753,N_13460,N_13542);
nor U13754 (N_13754,N_13420,N_13425);
or U13755 (N_13755,N_13490,N_13471);
or U13756 (N_13756,N_13545,N_13400);
or U13757 (N_13757,N_13462,N_13437);
xnor U13758 (N_13758,N_13558,N_13567);
and U13759 (N_13759,N_13477,N_13431);
and U13760 (N_13760,N_13432,N_13527);
nor U13761 (N_13761,N_13517,N_13451);
xnor U13762 (N_13762,N_13434,N_13532);
nor U13763 (N_13763,N_13511,N_13586);
and U13764 (N_13764,N_13498,N_13530);
xor U13765 (N_13765,N_13546,N_13595);
or U13766 (N_13766,N_13485,N_13432);
or U13767 (N_13767,N_13594,N_13441);
and U13768 (N_13768,N_13527,N_13546);
xor U13769 (N_13769,N_13495,N_13565);
or U13770 (N_13770,N_13478,N_13420);
or U13771 (N_13771,N_13470,N_13469);
nor U13772 (N_13772,N_13550,N_13422);
and U13773 (N_13773,N_13565,N_13464);
and U13774 (N_13774,N_13478,N_13563);
nand U13775 (N_13775,N_13526,N_13544);
xor U13776 (N_13776,N_13584,N_13450);
nor U13777 (N_13777,N_13564,N_13541);
or U13778 (N_13778,N_13564,N_13402);
nand U13779 (N_13779,N_13441,N_13546);
nor U13780 (N_13780,N_13427,N_13517);
nor U13781 (N_13781,N_13474,N_13531);
or U13782 (N_13782,N_13532,N_13518);
or U13783 (N_13783,N_13494,N_13420);
nor U13784 (N_13784,N_13476,N_13595);
nand U13785 (N_13785,N_13483,N_13584);
xor U13786 (N_13786,N_13503,N_13562);
or U13787 (N_13787,N_13444,N_13559);
nor U13788 (N_13788,N_13588,N_13581);
or U13789 (N_13789,N_13419,N_13465);
xor U13790 (N_13790,N_13439,N_13476);
or U13791 (N_13791,N_13429,N_13521);
or U13792 (N_13792,N_13440,N_13405);
and U13793 (N_13793,N_13540,N_13598);
and U13794 (N_13794,N_13462,N_13426);
nand U13795 (N_13795,N_13563,N_13465);
or U13796 (N_13796,N_13519,N_13441);
and U13797 (N_13797,N_13438,N_13468);
or U13798 (N_13798,N_13402,N_13572);
and U13799 (N_13799,N_13525,N_13476);
and U13800 (N_13800,N_13692,N_13693);
or U13801 (N_13801,N_13656,N_13707);
nor U13802 (N_13802,N_13783,N_13647);
nor U13803 (N_13803,N_13756,N_13713);
nand U13804 (N_13804,N_13767,N_13651);
and U13805 (N_13805,N_13643,N_13760);
nand U13806 (N_13806,N_13705,N_13711);
and U13807 (N_13807,N_13675,N_13620);
nor U13808 (N_13808,N_13748,N_13610);
xor U13809 (N_13809,N_13726,N_13744);
nand U13810 (N_13810,N_13665,N_13697);
and U13811 (N_13811,N_13634,N_13772);
xor U13812 (N_13812,N_13638,N_13673);
xor U13813 (N_13813,N_13788,N_13633);
nand U13814 (N_13814,N_13771,N_13699);
or U13815 (N_13815,N_13714,N_13703);
xnor U13816 (N_13816,N_13617,N_13600);
or U13817 (N_13817,N_13680,N_13609);
nor U13818 (N_13818,N_13653,N_13779);
and U13819 (N_13819,N_13676,N_13762);
nand U13820 (N_13820,N_13777,N_13613);
and U13821 (N_13821,N_13640,N_13719);
or U13822 (N_13822,N_13745,N_13642);
nor U13823 (N_13823,N_13752,N_13674);
xnor U13824 (N_13824,N_13632,N_13729);
nand U13825 (N_13825,N_13761,N_13795);
nand U13826 (N_13826,N_13612,N_13727);
and U13827 (N_13827,N_13746,N_13679);
and U13828 (N_13828,N_13698,N_13786);
nor U13829 (N_13829,N_13690,N_13768);
nand U13830 (N_13830,N_13796,N_13661);
and U13831 (N_13831,N_13781,N_13657);
xnor U13832 (N_13832,N_13753,N_13734);
nor U13833 (N_13833,N_13616,N_13790);
or U13834 (N_13834,N_13718,N_13784);
nor U13835 (N_13835,N_13700,N_13728);
or U13836 (N_13836,N_13626,N_13798);
and U13837 (N_13837,N_13789,N_13623);
or U13838 (N_13838,N_13664,N_13791);
and U13839 (N_13839,N_13636,N_13793);
or U13840 (N_13840,N_13721,N_13622);
nor U13841 (N_13841,N_13735,N_13797);
or U13842 (N_13842,N_13766,N_13758);
xor U13843 (N_13843,N_13606,N_13694);
and U13844 (N_13844,N_13695,N_13603);
xnor U13845 (N_13845,N_13681,N_13635);
xor U13846 (N_13846,N_13686,N_13644);
and U13847 (N_13847,N_13725,N_13701);
nand U13848 (N_13848,N_13776,N_13778);
or U13849 (N_13849,N_13792,N_13731);
nor U13850 (N_13850,N_13660,N_13627);
and U13851 (N_13851,N_13628,N_13751);
nor U13852 (N_13852,N_13631,N_13706);
and U13853 (N_13853,N_13742,N_13624);
or U13854 (N_13854,N_13654,N_13602);
nor U13855 (N_13855,N_13641,N_13607);
or U13856 (N_13856,N_13671,N_13630);
xnor U13857 (N_13857,N_13658,N_13787);
nor U13858 (N_13858,N_13637,N_13737);
xnor U13859 (N_13859,N_13730,N_13639);
xnor U13860 (N_13860,N_13733,N_13710);
xnor U13861 (N_13861,N_13667,N_13708);
nand U13862 (N_13862,N_13619,N_13782);
xnor U13863 (N_13863,N_13646,N_13655);
and U13864 (N_13864,N_13662,N_13615);
or U13865 (N_13865,N_13605,N_13743);
and U13866 (N_13866,N_13799,N_13738);
xor U13867 (N_13867,N_13720,N_13659);
or U13868 (N_13868,N_13614,N_13732);
nor U13869 (N_13869,N_13669,N_13611);
or U13870 (N_13870,N_13759,N_13763);
nor U13871 (N_13871,N_13670,N_13668);
nor U13872 (N_13872,N_13677,N_13629);
xor U13873 (N_13873,N_13755,N_13750);
or U13874 (N_13874,N_13652,N_13709);
nand U13875 (N_13875,N_13757,N_13650);
xor U13876 (N_13876,N_13747,N_13715);
xor U13877 (N_13877,N_13770,N_13683);
xor U13878 (N_13878,N_13608,N_13666);
and U13879 (N_13879,N_13773,N_13723);
nor U13880 (N_13880,N_13769,N_13740);
or U13881 (N_13881,N_13712,N_13785);
nand U13882 (N_13882,N_13749,N_13604);
nand U13883 (N_13883,N_13684,N_13716);
nand U13884 (N_13884,N_13687,N_13764);
and U13885 (N_13885,N_13724,N_13625);
or U13886 (N_13886,N_13704,N_13618);
nand U13887 (N_13887,N_13774,N_13645);
xnor U13888 (N_13888,N_13775,N_13689);
nand U13889 (N_13889,N_13648,N_13663);
or U13890 (N_13890,N_13688,N_13702);
nand U13891 (N_13891,N_13765,N_13794);
xor U13892 (N_13892,N_13780,N_13672);
or U13893 (N_13893,N_13717,N_13682);
or U13894 (N_13894,N_13722,N_13678);
xor U13895 (N_13895,N_13685,N_13741);
nor U13896 (N_13896,N_13754,N_13601);
xnor U13897 (N_13897,N_13736,N_13621);
xnor U13898 (N_13898,N_13739,N_13696);
xnor U13899 (N_13899,N_13649,N_13691);
nor U13900 (N_13900,N_13721,N_13698);
or U13901 (N_13901,N_13724,N_13722);
nand U13902 (N_13902,N_13717,N_13799);
and U13903 (N_13903,N_13647,N_13679);
and U13904 (N_13904,N_13751,N_13653);
nand U13905 (N_13905,N_13791,N_13779);
or U13906 (N_13906,N_13669,N_13771);
nor U13907 (N_13907,N_13783,N_13641);
or U13908 (N_13908,N_13756,N_13688);
nand U13909 (N_13909,N_13729,N_13792);
or U13910 (N_13910,N_13673,N_13699);
nor U13911 (N_13911,N_13711,N_13734);
nand U13912 (N_13912,N_13629,N_13756);
or U13913 (N_13913,N_13632,N_13745);
or U13914 (N_13914,N_13786,N_13619);
xor U13915 (N_13915,N_13630,N_13600);
xnor U13916 (N_13916,N_13648,N_13620);
or U13917 (N_13917,N_13727,N_13685);
xnor U13918 (N_13918,N_13630,N_13770);
or U13919 (N_13919,N_13678,N_13739);
nor U13920 (N_13920,N_13744,N_13752);
xnor U13921 (N_13921,N_13777,N_13688);
or U13922 (N_13922,N_13731,N_13781);
and U13923 (N_13923,N_13689,N_13645);
nor U13924 (N_13924,N_13740,N_13643);
nor U13925 (N_13925,N_13647,N_13623);
nand U13926 (N_13926,N_13772,N_13780);
nor U13927 (N_13927,N_13633,N_13743);
xor U13928 (N_13928,N_13785,N_13786);
xnor U13929 (N_13929,N_13637,N_13611);
nand U13930 (N_13930,N_13711,N_13647);
or U13931 (N_13931,N_13700,N_13644);
nand U13932 (N_13932,N_13621,N_13735);
nor U13933 (N_13933,N_13682,N_13783);
xor U13934 (N_13934,N_13712,N_13653);
nand U13935 (N_13935,N_13625,N_13631);
nand U13936 (N_13936,N_13693,N_13769);
nand U13937 (N_13937,N_13752,N_13640);
nand U13938 (N_13938,N_13683,N_13699);
and U13939 (N_13939,N_13655,N_13751);
nand U13940 (N_13940,N_13772,N_13732);
nand U13941 (N_13941,N_13748,N_13758);
xor U13942 (N_13942,N_13637,N_13675);
nor U13943 (N_13943,N_13717,N_13600);
xor U13944 (N_13944,N_13755,N_13713);
xnor U13945 (N_13945,N_13699,N_13611);
nor U13946 (N_13946,N_13781,N_13784);
and U13947 (N_13947,N_13732,N_13609);
and U13948 (N_13948,N_13672,N_13607);
and U13949 (N_13949,N_13655,N_13693);
nand U13950 (N_13950,N_13652,N_13627);
nor U13951 (N_13951,N_13654,N_13629);
nand U13952 (N_13952,N_13740,N_13655);
or U13953 (N_13953,N_13746,N_13789);
xnor U13954 (N_13954,N_13653,N_13698);
nor U13955 (N_13955,N_13698,N_13619);
nand U13956 (N_13956,N_13764,N_13604);
and U13957 (N_13957,N_13723,N_13758);
nand U13958 (N_13958,N_13777,N_13639);
xor U13959 (N_13959,N_13601,N_13693);
and U13960 (N_13960,N_13605,N_13777);
and U13961 (N_13961,N_13693,N_13608);
or U13962 (N_13962,N_13771,N_13797);
nand U13963 (N_13963,N_13746,N_13608);
nor U13964 (N_13964,N_13620,N_13629);
nand U13965 (N_13965,N_13609,N_13666);
xnor U13966 (N_13966,N_13649,N_13670);
and U13967 (N_13967,N_13703,N_13751);
or U13968 (N_13968,N_13699,N_13744);
xnor U13969 (N_13969,N_13720,N_13601);
nand U13970 (N_13970,N_13759,N_13799);
nor U13971 (N_13971,N_13654,N_13780);
or U13972 (N_13972,N_13794,N_13689);
nor U13973 (N_13973,N_13658,N_13766);
and U13974 (N_13974,N_13665,N_13602);
nor U13975 (N_13975,N_13716,N_13678);
or U13976 (N_13976,N_13708,N_13636);
and U13977 (N_13977,N_13740,N_13722);
nand U13978 (N_13978,N_13637,N_13621);
or U13979 (N_13979,N_13717,N_13731);
and U13980 (N_13980,N_13724,N_13662);
and U13981 (N_13981,N_13733,N_13736);
and U13982 (N_13982,N_13765,N_13703);
nor U13983 (N_13983,N_13744,N_13746);
nor U13984 (N_13984,N_13625,N_13731);
nand U13985 (N_13985,N_13696,N_13705);
and U13986 (N_13986,N_13716,N_13695);
nand U13987 (N_13987,N_13624,N_13680);
nor U13988 (N_13988,N_13653,N_13781);
or U13989 (N_13989,N_13669,N_13739);
xor U13990 (N_13990,N_13717,N_13759);
nor U13991 (N_13991,N_13719,N_13656);
nand U13992 (N_13992,N_13700,N_13664);
or U13993 (N_13993,N_13773,N_13672);
nand U13994 (N_13994,N_13662,N_13777);
xnor U13995 (N_13995,N_13729,N_13713);
nand U13996 (N_13996,N_13771,N_13713);
or U13997 (N_13997,N_13604,N_13746);
nor U13998 (N_13998,N_13693,N_13600);
or U13999 (N_13999,N_13635,N_13672);
and U14000 (N_14000,N_13972,N_13971);
xor U14001 (N_14001,N_13918,N_13915);
or U14002 (N_14002,N_13820,N_13898);
nor U14003 (N_14003,N_13886,N_13975);
or U14004 (N_14004,N_13834,N_13919);
and U14005 (N_14005,N_13865,N_13933);
xor U14006 (N_14006,N_13987,N_13977);
xnor U14007 (N_14007,N_13961,N_13835);
and U14008 (N_14008,N_13811,N_13872);
or U14009 (N_14009,N_13901,N_13969);
nor U14010 (N_14010,N_13809,N_13962);
and U14011 (N_14011,N_13980,N_13942);
nand U14012 (N_14012,N_13828,N_13803);
or U14013 (N_14013,N_13868,N_13857);
nor U14014 (N_14014,N_13876,N_13997);
nor U14015 (N_14015,N_13801,N_13827);
and U14016 (N_14016,N_13873,N_13922);
nand U14017 (N_14017,N_13985,N_13893);
or U14018 (N_14018,N_13900,N_13874);
or U14019 (N_14019,N_13965,N_13999);
and U14020 (N_14020,N_13846,N_13949);
nand U14021 (N_14021,N_13894,N_13910);
and U14022 (N_14022,N_13936,N_13887);
xnor U14023 (N_14023,N_13884,N_13851);
or U14024 (N_14024,N_13899,N_13862);
nand U14025 (N_14025,N_13804,N_13836);
and U14026 (N_14026,N_13853,N_13882);
xor U14027 (N_14027,N_13946,N_13968);
or U14028 (N_14028,N_13821,N_13990);
nor U14029 (N_14029,N_13907,N_13932);
or U14030 (N_14030,N_13986,N_13831);
xor U14031 (N_14031,N_13940,N_13976);
or U14032 (N_14032,N_13929,N_13814);
xnor U14033 (N_14033,N_13867,N_13974);
xor U14034 (N_14034,N_13914,N_13960);
and U14035 (N_14035,N_13925,N_13870);
nand U14036 (N_14036,N_13879,N_13822);
and U14037 (N_14037,N_13964,N_13802);
nor U14038 (N_14038,N_13864,N_13810);
and U14039 (N_14039,N_13998,N_13916);
xnor U14040 (N_14040,N_13924,N_13993);
nor U14041 (N_14041,N_13805,N_13895);
and U14042 (N_14042,N_13840,N_13889);
or U14043 (N_14043,N_13830,N_13902);
nor U14044 (N_14044,N_13838,N_13994);
nand U14045 (N_14045,N_13806,N_13989);
nand U14046 (N_14046,N_13845,N_13903);
or U14047 (N_14047,N_13913,N_13817);
xor U14048 (N_14048,N_13850,N_13863);
nand U14049 (N_14049,N_13984,N_13982);
nor U14050 (N_14050,N_13988,N_13928);
nor U14051 (N_14051,N_13826,N_13966);
and U14052 (N_14052,N_13935,N_13952);
or U14053 (N_14053,N_13837,N_13906);
xor U14054 (N_14054,N_13888,N_13896);
nor U14055 (N_14055,N_13883,N_13941);
and U14056 (N_14056,N_13812,N_13950);
nand U14057 (N_14057,N_13815,N_13927);
and U14058 (N_14058,N_13930,N_13920);
xnor U14059 (N_14059,N_13816,N_13849);
and U14060 (N_14060,N_13937,N_13943);
nor U14061 (N_14061,N_13897,N_13957);
nor U14062 (N_14062,N_13995,N_13848);
xor U14063 (N_14063,N_13818,N_13819);
or U14064 (N_14064,N_13861,N_13856);
and U14065 (N_14065,N_13892,N_13854);
nand U14066 (N_14066,N_13839,N_13841);
and U14067 (N_14067,N_13931,N_13959);
nand U14068 (N_14068,N_13947,N_13869);
and U14069 (N_14069,N_13909,N_13908);
xor U14070 (N_14070,N_13878,N_13858);
or U14071 (N_14071,N_13800,N_13938);
nor U14072 (N_14072,N_13983,N_13890);
and U14073 (N_14073,N_13880,N_13926);
xor U14074 (N_14074,N_13923,N_13967);
and U14075 (N_14075,N_13905,N_13813);
or U14076 (N_14076,N_13951,N_13945);
xor U14077 (N_14077,N_13981,N_13921);
or U14078 (N_14078,N_13991,N_13829);
xor U14079 (N_14079,N_13825,N_13855);
or U14080 (N_14080,N_13953,N_13956);
nor U14081 (N_14081,N_13917,N_13939);
xnor U14082 (N_14082,N_13911,N_13866);
nand U14083 (N_14083,N_13970,N_13996);
nor U14084 (N_14084,N_13963,N_13992);
or U14085 (N_14085,N_13823,N_13944);
and U14086 (N_14086,N_13973,N_13824);
nor U14087 (N_14087,N_13904,N_13875);
or U14088 (N_14088,N_13871,N_13958);
or U14089 (N_14089,N_13852,N_13859);
nor U14090 (N_14090,N_13860,N_13843);
and U14091 (N_14091,N_13912,N_13832);
nor U14092 (N_14092,N_13807,N_13948);
nand U14093 (N_14093,N_13844,N_13833);
nand U14094 (N_14094,N_13881,N_13877);
nor U14095 (N_14095,N_13954,N_13978);
or U14096 (N_14096,N_13891,N_13955);
nand U14097 (N_14097,N_13885,N_13934);
and U14098 (N_14098,N_13979,N_13808);
xnor U14099 (N_14099,N_13842,N_13847);
and U14100 (N_14100,N_13877,N_13990);
and U14101 (N_14101,N_13850,N_13936);
xor U14102 (N_14102,N_13867,N_13866);
nand U14103 (N_14103,N_13947,N_13964);
and U14104 (N_14104,N_13852,N_13880);
xor U14105 (N_14105,N_13802,N_13856);
nand U14106 (N_14106,N_13820,N_13863);
nand U14107 (N_14107,N_13896,N_13829);
nand U14108 (N_14108,N_13967,N_13872);
xnor U14109 (N_14109,N_13820,N_13958);
nand U14110 (N_14110,N_13870,N_13919);
nand U14111 (N_14111,N_13804,N_13953);
xnor U14112 (N_14112,N_13932,N_13829);
and U14113 (N_14113,N_13931,N_13808);
and U14114 (N_14114,N_13992,N_13967);
nor U14115 (N_14115,N_13899,N_13806);
and U14116 (N_14116,N_13971,N_13831);
and U14117 (N_14117,N_13870,N_13833);
or U14118 (N_14118,N_13814,N_13891);
nand U14119 (N_14119,N_13865,N_13801);
nand U14120 (N_14120,N_13966,N_13951);
xnor U14121 (N_14121,N_13824,N_13918);
xor U14122 (N_14122,N_13830,N_13821);
and U14123 (N_14123,N_13848,N_13833);
nand U14124 (N_14124,N_13818,N_13809);
nand U14125 (N_14125,N_13996,N_13980);
nor U14126 (N_14126,N_13864,N_13908);
nand U14127 (N_14127,N_13898,N_13918);
and U14128 (N_14128,N_13918,N_13905);
nor U14129 (N_14129,N_13898,N_13848);
nand U14130 (N_14130,N_13982,N_13846);
xnor U14131 (N_14131,N_13803,N_13988);
nor U14132 (N_14132,N_13804,N_13999);
and U14133 (N_14133,N_13859,N_13900);
xor U14134 (N_14134,N_13829,N_13828);
xnor U14135 (N_14135,N_13847,N_13862);
or U14136 (N_14136,N_13998,N_13950);
and U14137 (N_14137,N_13938,N_13849);
or U14138 (N_14138,N_13927,N_13869);
nor U14139 (N_14139,N_13979,N_13916);
and U14140 (N_14140,N_13903,N_13991);
and U14141 (N_14141,N_13934,N_13837);
xor U14142 (N_14142,N_13804,N_13996);
and U14143 (N_14143,N_13843,N_13922);
or U14144 (N_14144,N_13962,N_13916);
xnor U14145 (N_14145,N_13930,N_13875);
and U14146 (N_14146,N_13947,N_13854);
nor U14147 (N_14147,N_13904,N_13894);
nand U14148 (N_14148,N_13954,N_13971);
nor U14149 (N_14149,N_13906,N_13905);
nor U14150 (N_14150,N_13983,N_13874);
nor U14151 (N_14151,N_13885,N_13995);
xor U14152 (N_14152,N_13895,N_13926);
nor U14153 (N_14153,N_13831,N_13877);
xnor U14154 (N_14154,N_13964,N_13876);
or U14155 (N_14155,N_13807,N_13997);
nand U14156 (N_14156,N_13905,N_13984);
nor U14157 (N_14157,N_13896,N_13866);
or U14158 (N_14158,N_13879,N_13850);
xnor U14159 (N_14159,N_13890,N_13928);
nand U14160 (N_14160,N_13881,N_13815);
and U14161 (N_14161,N_13891,N_13859);
or U14162 (N_14162,N_13828,N_13866);
or U14163 (N_14163,N_13836,N_13812);
and U14164 (N_14164,N_13968,N_13889);
nand U14165 (N_14165,N_13997,N_13936);
or U14166 (N_14166,N_13857,N_13947);
and U14167 (N_14167,N_13848,N_13831);
xnor U14168 (N_14168,N_13838,N_13945);
nor U14169 (N_14169,N_13971,N_13964);
or U14170 (N_14170,N_13880,N_13922);
nor U14171 (N_14171,N_13997,N_13987);
nand U14172 (N_14172,N_13921,N_13966);
xnor U14173 (N_14173,N_13934,N_13890);
nor U14174 (N_14174,N_13950,N_13993);
xnor U14175 (N_14175,N_13858,N_13840);
xor U14176 (N_14176,N_13800,N_13899);
xnor U14177 (N_14177,N_13815,N_13906);
nor U14178 (N_14178,N_13805,N_13917);
or U14179 (N_14179,N_13880,N_13892);
and U14180 (N_14180,N_13896,N_13865);
xor U14181 (N_14181,N_13824,N_13963);
nand U14182 (N_14182,N_13947,N_13820);
xnor U14183 (N_14183,N_13961,N_13975);
xor U14184 (N_14184,N_13816,N_13930);
or U14185 (N_14185,N_13882,N_13854);
or U14186 (N_14186,N_13855,N_13991);
nor U14187 (N_14187,N_13800,N_13996);
nor U14188 (N_14188,N_13871,N_13913);
and U14189 (N_14189,N_13970,N_13927);
nor U14190 (N_14190,N_13812,N_13957);
nand U14191 (N_14191,N_13929,N_13862);
and U14192 (N_14192,N_13842,N_13943);
nor U14193 (N_14193,N_13876,N_13843);
xor U14194 (N_14194,N_13863,N_13972);
xnor U14195 (N_14195,N_13881,N_13833);
and U14196 (N_14196,N_13896,N_13923);
nor U14197 (N_14197,N_13987,N_13850);
nand U14198 (N_14198,N_13968,N_13969);
and U14199 (N_14199,N_13958,N_13821);
nor U14200 (N_14200,N_14184,N_14171);
nand U14201 (N_14201,N_14060,N_14059);
nor U14202 (N_14202,N_14013,N_14101);
and U14203 (N_14203,N_14092,N_14123);
nand U14204 (N_14204,N_14066,N_14033);
or U14205 (N_14205,N_14121,N_14199);
nor U14206 (N_14206,N_14020,N_14034);
nor U14207 (N_14207,N_14045,N_14192);
xor U14208 (N_14208,N_14135,N_14004);
xnor U14209 (N_14209,N_14076,N_14132);
or U14210 (N_14210,N_14153,N_14021);
nor U14211 (N_14211,N_14129,N_14159);
nor U14212 (N_14212,N_14117,N_14003);
nor U14213 (N_14213,N_14005,N_14111);
nor U14214 (N_14214,N_14134,N_14136);
nor U14215 (N_14215,N_14041,N_14038);
xnor U14216 (N_14216,N_14166,N_14036);
or U14217 (N_14217,N_14031,N_14099);
nor U14218 (N_14218,N_14081,N_14077);
nor U14219 (N_14219,N_14193,N_14185);
nand U14220 (N_14220,N_14182,N_14027);
or U14221 (N_14221,N_14011,N_14023);
nor U14222 (N_14222,N_14176,N_14174);
nor U14223 (N_14223,N_14056,N_14112);
nand U14224 (N_14224,N_14050,N_14030);
nand U14225 (N_14225,N_14120,N_14015);
nand U14226 (N_14226,N_14189,N_14052);
and U14227 (N_14227,N_14032,N_14179);
or U14228 (N_14228,N_14000,N_14178);
and U14229 (N_14229,N_14102,N_14061);
and U14230 (N_14230,N_14150,N_14090);
or U14231 (N_14231,N_14025,N_14043);
nand U14232 (N_14232,N_14188,N_14143);
nor U14233 (N_14233,N_14109,N_14054);
nand U14234 (N_14234,N_14048,N_14149);
xor U14235 (N_14235,N_14139,N_14097);
nand U14236 (N_14236,N_14161,N_14085);
nand U14237 (N_14237,N_14016,N_14100);
xnor U14238 (N_14238,N_14105,N_14187);
xor U14239 (N_14239,N_14009,N_14051);
xor U14240 (N_14240,N_14125,N_14162);
nor U14241 (N_14241,N_14122,N_14116);
or U14242 (N_14242,N_14091,N_14164);
and U14243 (N_14243,N_14177,N_14024);
nand U14244 (N_14244,N_14096,N_14198);
and U14245 (N_14245,N_14010,N_14088);
nand U14246 (N_14246,N_14181,N_14086);
xnor U14247 (N_14247,N_14106,N_14113);
xor U14248 (N_14248,N_14042,N_14062);
and U14249 (N_14249,N_14124,N_14190);
or U14250 (N_14250,N_14186,N_14163);
and U14251 (N_14251,N_14104,N_14014);
nand U14252 (N_14252,N_14007,N_14055);
and U14253 (N_14253,N_14197,N_14058);
xor U14254 (N_14254,N_14047,N_14040);
nand U14255 (N_14255,N_14035,N_14152);
nand U14256 (N_14256,N_14065,N_14167);
or U14257 (N_14257,N_14145,N_14138);
and U14258 (N_14258,N_14080,N_14157);
nand U14259 (N_14259,N_14064,N_14095);
or U14260 (N_14260,N_14070,N_14049);
nand U14261 (N_14261,N_14130,N_14169);
and U14262 (N_14262,N_14039,N_14079);
or U14263 (N_14263,N_14073,N_14175);
and U14264 (N_14264,N_14094,N_14142);
xor U14265 (N_14265,N_14151,N_14156);
xnor U14266 (N_14266,N_14019,N_14063);
xor U14267 (N_14267,N_14180,N_14195);
xor U14268 (N_14268,N_14022,N_14127);
and U14269 (N_14269,N_14026,N_14196);
nor U14270 (N_14270,N_14001,N_14160);
nand U14271 (N_14271,N_14071,N_14147);
xor U14272 (N_14272,N_14119,N_14115);
nor U14273 (N_14273,N_14012,N_14053);
or U14274 (N_14274,N_14170,N_14093);
and U14275 (N_14275,N_14165,N_14069);
nor U14276 (N_14276,N_14046,N_14075);
nor U14277 (N_14277,N_14140,N_14098);
and U14278 (N_14278,N_14148,N_14057);
nor U14279 (N_14279,N_14155,N_14118);
nand U14280 (N_14280,N_14103,N_14078);
or U14281 (N_14281,N_14131,N_14107);
nor U14282 (N_14282,N_14087,N_14083);
and U14283 (N_14283,N_14128,N_14172);
and U14284 (N_14284,N_14002,N_14006);
xnor U14285 (N_14285,N_14037,N_14137);
nor U14286 (N_14286,N_14028,N_14141);
and U14287 (N_14287,N_14158,N_14133);
and U14288 (N_14288,N_14114,N_14017);
nor U14289 (N_14289,N_14110,N_14018);
nand U14290 (N_14290,N_14008,N_14029);
or U14291 (N_14291,N_14068,N_14191);
nor U14292 (N_14292,N_14044,N_14183);
and U14293 (N_14293,N_14168,N_14072);
xnor U14294 (N_14294,N_14089,N_14074);
nor U14295 (N_14295,N_14067,N_14084);
and U14296 (N_14296,N_14173,N_14146);
and U14297 (N_14297,N_14154,N_14144);
nand U14298 (N_14298,N_14194,N_14108);
nor U14299 (N_14299,N_14126,N_14082);
or U14300 (N_14300,N_14129,N_14002);
and U14301 (N_14301,N_14032,N_14149);
nand U14302 (N_14302,N_14196,N_14085);
xnor U14303 (N_14303,N_14141,N_14154);
xor U14304 (N_14304,N_14122,N_14077);
and U14305 (N_14305,N_14054,N_14175);
and U14306 (N_14306,N_14089,N_14187);
nor U14307 (N_14307,N_14018,N_14184);
nor U14308 (N_14308,N_14057,N_14194);
nor U14309 (N_14309,N_14199,N_14150);
and U14310 (N_14310,N_14118,N_14021);
nand U14311 (N_14311,N_14130,N_14045);
nand U14312 (N_14312,N_14104,N_14149);
nand U14313 (N_14313,N_14016,N_14013);
or U14314 (N_14314,N_14039,N_14026);
nand U14315 (N_14315,N_14165,N_14056);
nor U14316 (N_14316,N_14185,N_14161);
xor U14317 (N_14317,N_14196,N_14162);
xnor U14318 (N_14318,N_14108,N_14097);
nor U14319 (N_14319,N_14003,N_14040);
or U14320 (N_14320,N_14003,N_14011);
nor U14321 (N_14321,N_14164,N_14172);
nand U14322 (N_14322,N_14031,N_14015);
xor U14323 (N_14323,N_14120,N_14167);
xor U14324 (N_14324,N_14154,N_14031);
nand U14325 (N_14325,N_14126,N_14052);
nor U14326 (N_14326,N_14150,N_14156);
and U14327 (N_14327,N_14022,N_14035);
and U14328 (N_14328,N_14134,N_14146);
xnor U14329 (N_14329,N_14038,N_14010);
nor U14330 (N_14330,N_14192,N_14119);
nand U14331 (N_14331,N_14092,N_14163);
nor U14332 (N_14332,N_14166,N_14188);
xnor U14333 (N_14333,N_14188,N_14007);
or U14334 (N_14334,N_14081,N_14168);
nand U14335 (N_14335,N_14015,N_14166);
and U14336 (N_14336,N_14123,N_14145);
xnor U14337 (N_14337,N_14118,N_14187);
nand U14338 (N_14338,N_14189,N_14176);
or U14339 (N_14339,N_14180,N_14134);
xnor U14340 (N_14340,N_14148,N_14184);
nor U14341 (N_14341,N_14086,N_14117);
nand U14342 (N_14342,N_14126,N_14012);
or U14343 (N_14343,N_14101,N_14174);
and U14344 (N_14344,N_14003,N_14139);
xor U14345 (N_14345,N_14199,N_14122);
and U14346 (N_14346,N_14078,N_14005);
nand U14347 (N_14347,N_14083,N_14161);
and U14348 (N_14348,N_14184,N_14051);
nor U14349 (N_14349,N_14181,N_14053);
xor U14350 (N_14350,N_14090,N_14097);
and U14351 (N_14351,N_14186,N_14085);
and U14352 (N_14352,N_14124,N_14041);
and U14353 (N_14353,N_14033,N_14016);
nor U14354 (N_14354,N_14141,N_14117);
nor U14355 (N_14355,N_14109,N_14183);
nor U14356 (N_14356,N_14177,N_14060);
and U14357 (N_14357,N_14153,N_14173);
or U14358 (N_14358,N_14186,N_14165);
xor U14359 (N_14359,N_14042,N_14136);
nand U14360 (N_14360,N_14011,N_14068);
xor U14361 (N_14361,N_14196,N_14121);
xnor U14362 (N_14362,N_14009,N_14020);
xor U14363 (N_14363,N_14161,N_14160);
nor U14364 (N_14364,N_14112,N_14162);
and U14365 (N_14365,N_14103,N_14006);
and U14366 (N_14366,N_14172,N_14197);
xnor U14367 (N_14367,N_14112,N_14006);
nand U14368 (N_14368,N_14123,N_14103);
nor U14369 (N_14369,N_14049,N_14014);
and U14370 (N_14370,N_14046,N_14194);
or U14371 (N_14371,N_14188,N_14177);
or U14372 (N_14372,N_14191,N_14109);
nor U14373 (N_14373,N_14074,N_14154);
and U14374 (N_14374,N_14090,N_14140);
xnor U14375 (N_14375,N_14131,N_14100);
and U14376 (N_14376,N_14186,N_14047);
nand U14377 (N_14377,N_14116,N_14004);
xor U14378 (N_14378,N_14081,N_14114);
xnor U14379 (N_14379,N_14081,N_14138);
xnor U14380 (N_14380,N_14136,N_14147);
or U14381 (N_14381,N_14001,N_14123);
and U14382 (N_14382,N_14052,N_14181);
and U14383 (N_14383,N_14118,N_14001);
and U14384 (N_14384,N_14043,N_14023);
xnor U14385 (N_14385,N_14021,N_14007);
xor U14386 (N_14386,N_14038,N_14164);
nor U14387 (N_14387,N_14101,N_14083);
xnor U14388 (N_14388,N_14125,N_14018);
nand U14389 (N_14389,N_14164,N_14001);
or U14390 (N_14390,N_14045,N_14137);
xnor U14391 (N_14391,N_14019,N_14115);
and U14392 (N_14392,N_14137,N_14135);
nor U14393 (N_14393,N_14193,N_14166);
or U14394 (N_14394,N_14021,N_14186);
nand U14395 (N_14395,N_14006,N_14140);
or U14396 (N_14396,N_14034,N_14109);
or U14397 (N_14397,N_14182,N_14003);
nand U14398 (N_14398,N_14092,N_14174);
or U14399 (N_14399,N_14080,N_14067);
nand U14400 (N_14400,N_14344,N_14296);
or U14401 (N_14401,N_14214,N_14376);
or U14402 (N_14402,N_14259,N_14359);
nor U14403 (N_14403,N_14272,N_14279);
nand U14404 (N_14404,N_14233,N_14268);
xor U14405 (N_14405,N_14249,N_14385);
xnor U14406 (N_14406,N_14331,N_14380);
or U14407 (N_14407,N_14384,N_14250);
or U14408 (N_14408,N_14324,N_14243);
xor U14409 (N_14409,N_14394,N_14230);
nand U14410 (N_14410,N_14398,N_14245);
and U14411 (N_14411,N_14289,N_14201);
nor U14412 (N_14412,N_14286,N_14232);
xnor U14413 (N_14413,N_14336,N_14317);
nand U14414 (N_14414,N_14399,N_14310);
nor U14415 (N_14415,N_14262,N_14255);
nor U14416 (N_14416,N_14258,N_14313);
or U14417 (N_14417,N_14276,N_14298);
xor U14418 (N_14418,N_14288,N_14216);
nor U14419 (N_14419,N_14391,N_14383);
xor U14420 (N_14420,N_14274,N_14221);
nand U14421 (N_14421,N_14254,N_14375);
or U14422 (N_14422,N_14370,N_14200);
nand U14423 (N_14423,N_14364,N_14326);
nor U14424 (N_14424,N_14367,N_14278);
xnor U14425 (N_14425,N_14318,N_14323);
and U14426 (N_14426,N_14395,N_14351);
nor U14427 (N_14427,N_14277,N_14382);
and U14428 (N_14428,N_14388,N_14332);
xor U14429 (N_14429,N_14273,N_14379);
nand U14430 (N_14430,N_14307,N_14372);
and U14431 (N_14431,N_14240,N_14284);
and U14432 (N_14432,N_14287,N_14209);
nor U14433 (N_14433,N_14213,N_14347);
xnor U14434 (N_14434,N_14308,N_14354);
xnor U14435 (N_14435,N_14275,N_14361);
nand U14436 (N_14436,N_14334,N_14238);
nor U14437 (N_14437,N_14346,N_14312);
and U14438 (N_14438,N_14363,N_14340);
nor U14439 (N_14439,N_14397,N_14269);
nand U14440 (N_14440,N_14236,N_14231);
or U14441 (N_14441,N_14356,N_14328);
nand U14442 (N_14442,N_14348,N_14244);
nand U14443 (N_14443,N_14319,N_14343);
or U14444 (N_14444,N_14297,N_14208);
and U14445 (N_14445,N_14322,N_14220);
nand U14446 (N_14446,N_14369,N_14271);
and U14447 (N_14447,N_14225,N_14285);
and U14448 (N_14448,N_14325,N_14349);
or U14449 (N_14449,N_14228,N_14373);
and U14450 (N_14450,N_14342,N_14247);
or U14451 (N_14451,N_14335,N_14396);
or U14452 (N_14452,N_14248,N_14282);
nor U14453 (N_14453,N_14360,N_14265);
nor U14454 (N_14454,N_14242,N_14299);
nand U14455 (N_14455,N_14264,N_14329);
and U14456 (N_14456,N_14293,N_14311);
nor U14457 (N_14457,N_14390,N_14235);
nand U14458 (N_14458,N_14305,N_14345);
xnor U14459 (N_14459,N_14314,N_14306);
and U14460 (N_14460,N_14393,N_14229);
xnor U14461 (N_14461,N_14357,N_14392);
or U14462 (N_14462,N_14315,N_14350);
nand U14463 (N_14463,N_14256,N_14212);
and U14464 (N_14464,N_14355,N_14260);
nor U14465 (N_14465,N_14207,N_14251);
or U14466 (N_14466,N_14205,N_14316);
nor U14467 (N_14467,N_14267,N_14283);
nand U14468 (N_14468,N_14327,N_14341);
nor U14469 (N_14469,N_14381,N_14358);
xnor U14470 (N_14470,N_14252,N_14378);
nor U14471 (N_14471,N_14234,N_14215);
and U14472 (N_14472,N_14241,N_14387);
and U14473 (N_14473,N_14222,N_14365);
and U14474 (N_14474,N_14377,N_14263);
xnor U14475 (N_14475,N_14257,N_14294);
nand U14476 (N_14476,N_14295,N_14300);
and U14477 (N_14477,N_14227,N_14320);
or U14478 (N_14478,N_14203,N_14202);
or U14479 (N_14479,N_14371,N_14266);
nor U14480 (N_14480,N_14210,N_14281);
or U14481 (N_14481,N_14211,N_14280);
xnor U14482 (N_14482,N_14338,N_14352);
or U14483 (N_14483,N_14291,N_14309);
nand U14484 (N_14484,N_14292,N_14204);
nor U14485 (N_14485,N_14237,N_14224);
nand U14486 (N_14486,N_14253,N_14246);
xor U14487 (N_14487,N_14206,N_14301);
and U14488 (N_14488,N_14223,N_14226);
and U14489 (N_14489,N_14337,N_14303);
and U14490 (N_14490,N_14333,N_14290);
xor U14491 (N_14491,N_14362,N_14389);
xnor U14492 (N_14492,N_14374,N_14219);
xor U14493 (N_14493,N_14270,N_14353);
xor U14494 (N_14494,N_14386,N_14217);
nand U14495 (N_14495,N_14261,N_14368);
and U14496 (N_14496,N_14239,N_14218);
xor U14497 (N_14497,N_14321,N_14366);
xor U14498 (N_14498,N_14302,N_14304);
xor U14499 (N_14499,N_14339,N_14330);
or U14500 (N_14500,N_14389,N_14370);
and U14501 (N_14501,N_14378,N_14241);
nor U14502 (N_14502,N_14284,N_14328);
nand U14503 (N_14503,N_14314,N_14359);
nand U14504 (N_14504,N_14369,N_14211);
or U14505 (N_14505,N_14326,N_14352);
or U14506 (N_14506,N_14268,N_14297);
nand U14507 (N_14507,N_14312,N_14349);
nor U14508 (N_14508,N_14313,N_14307);
nand U14509 (N_14509,N_14367,N_14250);
nand U14510 (N_14510,N_14230,N_14239);
or U14511 (N_14511,N_14307,N_14314);
xor U14512 (N_14512,N_14375,N_14210);
nand U14513 (N_14513,N_14239,N_14221);
nor U14514 (N_14514,N_14270,N_14249);
xor U14515 (N_14515,N_14256,N_14211);
xnor U14516 (N_14516,N_14222,N_14252);
or U14517 (N_14517,N_14273,N_14335);
xor U14518 (N_14518,N_14217,N_14206);
nor U14519 (N_14519,N_14246,N_14212);
xnor U14520 (N_14520,N_14396,N_14369);
nor U14521 (N_14521,N_14344,N_14290);
nor U14522 (N_14522,N_14215,N_14327);
nor U14523 (N_14523,N_14203,N_14229);
nor U14524 (N_14524,N_14340,N_14370);
nor U14525 (N_14525,N_14252,N_14327);
or U14526 (N_14526,N_14319,N_14287);
and U14527 (N_14527,N_14305,N_14320);
or U14528 (N_14528,N_14254,N_14247);
nor U14529 (N_14529,N_14205,N_14263);
or U14530 (N_14530,N_14209,N_14344);
and U14531 (N_14531,N_14358,N_14212);
nand U14532 (N_14532,N_14300,N_14215);
or U14533 (N_14533,N_14305,N_14297);
or U14534 (N_14534,N_14378,N_14326);
or U14535 (N_14535,N_14347,N_14234);
nand U14536 (N_14536,N_14227,N_14368);
and U14537 (N_14537,N_14290,N_14231);
nor U14538 (N_14538,N_14345,N_14268);
nand U14539 (N_14539,N_14375,N_14310);
and U14540 (N_14540,N_14205,N_14241);
and U14541 (N_14541,N_14274,N_14363);
nor U14542 (N_14542,N_14350,N_14287);
xor U14543 (N_14543,N_14334,N_14214);
or U14544 (N_14544,N_14388,N_14252);
and U14545 (N_14545,N_14351,N_14296);
nor U14546 (N_14546,N_14352,N_14243);
nor U14547 (N_14547,N_14218,N_14357);
and U14548 (N_14548,N_14313,N_14346);
nor U14549 (N_14549,N_14309,N_14221);
nand U14550 (N_14550,N_14338,N_14280);
xor U14551 (N_14551,N_14331,N_14349);
xnor U14552 (N_14552,N_14380,N_14315);
and U14553 (N_14553,N_14283,N_14265);
nor U14554 (N_14554,N_14369,N_14284);
nand U14555 (N_14555,N_14255,N_14324);
nor U14556 (N_14556,N_14343,N_14331);
or U14557 (N_14557,N_14391,N_14370);
xor U14558 (N_14558,N_14203,N_14244);
nand U14559 (N_14559,N_14389,N_14383);
nand U14560 (N_14560,N_14274,N_14326);
and U14561 (N_14561,N_14265,N_14217);
xor U14562 (N_14562,N_14357,N_14361);
or U14563 (N_14563,N_14218,N_14257);
or U14564 (N_14564,N_14380,N_14309);
nand U14565 (N_14565,N_14327,N_14398);
or U14566 (N_14566,N_14344,N_14234);
nand U14567 (N_14567,N_14344,N_14254);
nand U14568 (N_14568,N_14229,N_14271);
or U14569 (N_14569,N_14315,N_14342);
and U14570 (N_14570,N_14371,N_14210);
or U14571 (N_14571,N_14278,N_14326);
nand U14572 (N_14572,N_14274,N_14257);
and U14573 (N_14573,N_14231,N_14233);
nand U14574 (N_14574,N_14226,N_14271);
or U14575 (N_14575,N_14347,N_14349);
xor U14576 (N_14576,N_14285,N_14379);
and U14577 (N_14577,N_14288,N_14375);
nand U14578 (N_14578,N_14374,N_14221);
xnor U14579 (N_14579,N_14387,N_14389);
xnor U14580 (N_14580,N_14264,N_14360);
and U14581 (N_14581,N_14206,N_14295);
xnor U14582 (N_14582,N_14276,N_14224);
nand U14583 (N_14583,N_14251,N_14231);
or U14584 (N_14584,N_14261,N_14388);
and U14585 (N_14585,N_14391,N_14361);
nand U14586 (N_14586,N_14263,N_14375);
or U14587 (N_14587,N_14362,N_14308);
or U14588 (N_14588,N_14324,N_14310);
nor U14589 (N_14589,N_14294,N_14335);
or U14590 (N_14590,N_14325,N_14306);
nor U14591 (N_14591,N_14224,N_14354);
xnor U14592 (N_14592,N_14239,N_14327);
xor U14593 (N_14593,N_14225,N_14240);
and U14594 (N_14594,N_14386,N_14342);
or U14595 (N_14595,N_14214,N_14210);
nor U14596 (N_14596,N_14356,N_14226);
xor U14597 (N_14597,N_14297,N_14316);
or U14598 (N_14598,N_14298,N_14282);
nand U14599 (N_14599,N_14257,N_14362);
xnor U14600 (N_14600,N_14521,N_14439);
nor U14601 (N_14601,N_14487,N_14569);
nor U14602 (N_14602,N_14444,N_14412);
nand U14603 (N_14603,N_14571,N_14411);
nor U14604 (N_14604,N_14574,N_14558);
nand U14605 (N_14605,N_14583,N_14489);
or U14606 (N_14606,N_14564,N_14581);
xor U14607 (N_14607,N_14425,N_14511);
nor U14608 (N_14608,N_14575,N_14495);
xor U14609 (N_14609,N_14585,N_14541);
and U14610 (N_14610,N_14526,N_14502);
and U14611 (N_14611,N_14517,N_14453);
nor U14612 (N_14612,N_14401,N_14553);
xor U14613 (N_14613,N_14480,N_14445);
nor U14614 (N_14614,N_14539,N_14507);
xnor U14615 (N_14615,N_14586,N_14594);
xnor U14616 (N_14616,N_14469,N_14408);
and U14617 (N_14617,N_14400,N_14527);
nor U14618 (N_14618,N_14573,N_14435);
xnor U14619 (N_14619,N_14410,N_14538);
xor U14620 (N_14620,N_14593,N_14457);
or U14621 (N_14621,N_14543,N_14458);
and U14622 (N_14622,N_14447,N_14556);
xnor U14623 (N_14623,N_14560,N_14483);
xor U14624 (N_14624,N_14474,N_14528);
and U14625 (N_14625,N_14509,N_14542);
nand U14626 (N_14626,N_14493,N_14406);
or U14627 (N_14627,N_14578,N_14433);
nor U14628 (N_14628,N_14422,N_14515);
nand U14629 (N_14629,N_14547,N_14580);
nand U14630 (N_14630,N_14468,N_14525);
or U14631 (N_14631,N_14419,N_14530);
nor U14632 (N_14632,N_14471,N_14418);
nor U14633 (N_14633,N_14473,N_14448);
nor U14634 (N_14634,N_14520,N_14464);
nand U14635 (N_14635,N_14529,N_14597);
nand U14636 (N_14636,N_14470,N_14467);
nor U14637 (N_14637,N_14415,N_14478);
xor U14638 (N_14638,N_14563,N_14416);
or U14639 (N_14639,N_14430,N_14442);
nor U14640 (N_14640,N_14544,N_14548);
xor U14641 (N_14641,N_14508,N_14536);
xnor U14642 (N_14642,N_14417,N_14516);
and U14643 (N_14643,N_14554,N_14591);
nand U14644 (N_14644,N_14537,N_14421);
and U14645 (N_14645,N_14588,N_14463);
and U14646 (N_14646,N_14562,N_14452);
and U14647 (N_14647,N_14565,N_14404);
or U14648 (N_14648,N_14598,N_14449);
or U14649 (N_14649,N_14432,N_14555);
nor U14650 (N_14650,N_14518,N_14500);
xnor U14651 (N_14651,N_14407,N_14590);
nor U14652 (N_14652,N_14557,N_14485);
or U14653 (N_14653,N_14545,N_14413);
or U14654 (N_14654,N_14551,N_14595);
or U14655 (N_14655,N_14481,N_14535);
nand U14656 (N_14656,N_14599,N_14426);
nand U14657 (N_14657,N_14497,N_14503);
or U14658 (N_14658,N_14434,N_14486);
or U14659 (N_14659,N_14579,N_14499);
nand U14660 (N_14660,N_14459,N_14559);
nor U14661 (N_14661,N_14567,N_14494);
nand U14662 (N_14662,N_14437,N_14519);
nand U14663 (N_14663,N_14477,N_14550);
xor U14664 (N_14664,N_14587,N_14524);
and U14665 (N_14665,N_14506,N_14491);
nand U14666 (N_14666,N_14462,N_14523);
nor U14667 (N_14667,N_14414,N_14450);
nand U14668 (N_14668,N_14552,N_14451);
nand U14669 (N_14669,N_14561,N_14492);
and U14670 (N_14670,N_14455,N_14436);
xnor U14671 (N_14671,N_14576,N_14505);
nand U14672 (N_14672,N_14566,N_14577);
or U14673 (N_14673,N_14438,N_14596);
nand U14674 (N_14674,N_14472,N_14443);
nor U14675 (N_14675,N_14533,N_14582);
xnor U14676 (N_14676,N_14479,N_14488);
and U14677 (N_14677,N_14475,N_14496);
nand U14678 (N_14678,N_14589,N_14484);
nor U14679 (N_14679,N_14402,N_14428);
or U14680 (N_14680,N_14568,N_14440);
nand U14681 (N_14681,N_14534,N_14531);
or U14682 (N_14682,N_14427,N_14461);
nand U14683 (N_14683,N_14429,N_14456);
nor U14684 (N_14684,N_14504,N_14510);
nor U14685 (N_14685,N_14482,N_14423);
nor U14686 (N_14686,N_14409,N_14465);
or U14687 (N_14687,N_14513,N_14490);
and U14688 (N_14688,N_14498,N_14546);
or U14689 (N_14689,N_14441,N_14431);
nor U14690 (N_14690,N_14522,N_14420);
nor U14691 (N_14691,N_14592,N_14512);
or U14692 (N_14692,N_14514,N_14570);
and U14693 (N_14693,N_14446,N_14424);
or U14694 (N_14694,N_14501,N_14454);
nor U14695 (N_14695,N_14405,N_14549);
and U14696 (N_14696,N_14476,N_14540);
or U14697 (N_14697,N_14572,N_14403);
nor U14698 (N_14698,N_14466,N_14460);
nor U14699 (N_14699,N_14532,N_14584);
or U14700 (N_14700,N_14434,N_14400);
or U14701 (N_14701,N_14499,N_14456);
nand U14702 (N_14702,N_14429,N_14469);
xor U14703 (N_14703,N_14576,N_14560);
xor U14704 (N_14704,N_14409,N_14507);
xor U14705 (N_14705,N_14507,N_14435);
nor U14706 (N_14706,N_14422,N_14566);
nand U14707 (N_14707,N_14427,N_14426);
and U14708 (N_14708,N_14584,N_14424);
xnor U14709 (N_14709,N_14486,N_14463);
nand U14710 (N_14710,N_14417,N_14423);
and U14711 (N_14711,N_14548,N_14481);
nor U14712 (N_14712,N_14496,N_14583);
and U14713 (N_14713,N_14574,N_14485);
and U14714 (N_14714,N_14533,N_14531);
or U14715 (N_14715,N_14400,N_14545);
or U14716 (N_14716,N_14454,N_14442);
or U14717 (N_14717,N_14455,N_14489);
nand U14718 (N_14718,N_14582,N_14513);
or U14719 (N_14719,N_14421,N_14523);
nor U14720 (N_14720,N_14485,N_14519);
and U14721 (N_14721,N_14481,N_14578);
xor U14722 (N_14722,N_14432,N_14481);
xor U14723 (N_14723,N_14509,N_14485);
nand U14724 (N_14724,N_14470,N_14545);
or U14725 (N_14725,N_14508,N_14440);
nand U14726 (N_14726,N_14448,N_14490);
xor U14727 (N_14727,N_14570,N_14591);
nand U14728 (N_14728,N_14547,N_14412);
xor U14729 (N_14729,N_14476,N_14573);
nand U14730 (N_14730,N_14576,N_14447);
and U14731 (N_14731,N_14455,N_14583);
xor U14732 (N_14732,N_14518,N_14465);
and U14733 (N_14733,N_14510,N_14488);
and U14734 (N_14734,N_14588,N_14457);
or U14735 (N_14735,N_14462,N_14451);
or U14736 (N_14736,N_14474,N_14403);
nand U14737 (N_14737,N_14496,N_14464);
and U14738 (N_14738,N_14593,N_14460);
or U14739 (N_14739,N_14578,N_14462);
xor U14740 (N_14740,N_14489,N_14408);
nor U14741 (N_14741,N_14522,N_14543);
nand U14742 (N_14742,N_14514,N_14597);
and U14743 (N_14743,N_14421,N_14549);
and U14744 (N_14744,N_14582,N_14498);
or U14745 (N_14745,N_14579,N_14584);
xor U14746 (N_14746,N_14519,N_14479);
and U14747 (N_14747,N_14444,N_14593);
nor U14748 (N_14748,N_14560,N_14533);
or U14749 (N_14749,N_14469,N_14415);
and U14750 (N_14750,N_14538,N_14429);
nand U14751 (N_14751,N_14537,N_14470);
and U14752 (N_14752,N_14468,N_14417);
and U14753 (N_14753,N_14562,N_14542);
nor U14754 (N_14754,N_14549,N_14568);
and U14755 (N_14755,N_14522,N_14476);
nor U14756 (N_14756,N_14410,N_14575);
nor U14757 (N_14757,N_14503,N_14558);
and U14758 (N_14758,N_14591,N_14579);
or U14759 (N_14759,N_14598,N_14578);
or U14760 (N_14760,N_14596,N_14478);
xor U14761 (N_14761,N_14495,N_14574);
xnor U14762 (N_14762,N_14435,N_14470);
and U14763 (N_14763,N_14417,N_14558);
and U14764 (N_14764,N_14507,N_14504);
and U14765 (N_14765,N_14536,N_14473);
xnor U14766 (N_14766,N_14558,N_14561);
or U14767 (N_14767,N_14591,N_14516);
and U14768 (N_14768,N_14565,N_14478);
xor U14769 (N_14769,N_14470,N_14513);
and U14770 (N_14770,N_14434,N_14472);
and U14771 (N_14771,N_14422,N_14530);
and U14772 (N_14772,N_14599,N_14470);
and U14773 (N_14773,N_14405,N_14550);
xor U14774 (N_14774,N_14464,N_14466);
nor U14775 (N_14775,N_14498,N_14451);
xor U14776 (N_14776,N_14575,N_14572);
nor U14777 (N_14777,N_14490,N_14505);
or U14778 (N_14778,N_14590,N_14463);
nand U14779 (N_14779,N_14474,N_14412);
nor U14780 (N_14780,N_14470,N_14511);
xnor U14781 (N_14781,N_14464,N_14494);
and U14782 (N_14782,N_14404,N_14575);
and U14783 (N_14783,N_14556,N_14435);
xnor U14784 (N_14784,N_14565,N_14559);
nor U14785 (N_14785,N_14584,N_14400);
nor U14786 (N_14786,N_14539,N_14415);
xnor U14787 (N_14787,N_14530,N_14424);
nor U14788 (N_14788,N_14441,N_14412);
and U14789 (N_14789,N_14412,N_14451);
nand U14790 (N_14790,N_14549,N_14451);
or U14791 (N_14791,N_14491,N_14453);
nor U14792 (N_14792,N_14415,N_14419);
and U14793 (N_14793,N_14543,N_14565);
and U14794 (N_14794,N_14566,N_14487);
or U14795 (N_14795,N_14483,N_14519);
xnor U14796 (N_14796,N_14411,N_14532);
and U14797 (N_14797,N_14475,N_14473);
xnor U14798 (N_14798,N_14444,N_14415);
or U14799 (N_14799,N_14583,N_14429);
xnor U14800 (N_14800,N_14705,N_14794);
xor U14801 (N_14801,N_14656,N_14730);
nor U14802 (N_14802,N_14744,N_14662);
nor U14803 (N_14803,N_14682,N_14733);
xnor U14804 (N_14804,N_14661,N_14765);
nor U14805 (N_14805,N_14643,N_14603);
and U14806 (N_14806,N_14612,N_14691);
nand U14807 (N_14807,N_14727,N_14664);
or U14808 (N_14808,N_14622,N_14666);
and U14809 (N_14809,N_14792,N_14609);
or U14810 (N_14810,N_14755,N_14614);
nand U14811 (N_14811,N_14710,N_14639);
or U14812 (N_14812,N_14734,N_14601);
xor U14813 (N_14813,N_14787,N_14665);
nor U14814 (N_14814,N_14752,N_14717);
and U14815 (N_14815,N_14676,N_14715);
or U14816 (N_14816,N_14748,N_14762);
and U14817 (N_14817,N_14753,N_14754);
nor U14818 (N_14818,N_14620,N_14640);
and U14819 (N_14819,N_14736,N_14780);
nor U14820 (N_14820,N_14788,N_14797);
nand U14821 (N_14821,N_14735,N_14627);
nand U14822 (N_14822,N_14740,N_14675);
xnor U14823 (N_14823,N_14677,N_14635);
xor U14824 (N_14824,N_14799,N_14713);
xor U14825 (N_14825,N_14774,N_14625);
nor U14826 (N_14826,N_14701,N_14758);
nor U14827 (N_14827,N_14729,N_14783);
nor U14828 (N_14828,N_14619,N_14667);
nand U14829 (N_14829,N_14658,N_14617);
nor U14830 (N_14830,N_14696,N_14793);
nor U14831 (N_14831,N_14638,N_14618);
nand U14832 (N_14832,N_14721,N_14669);
xor U14833 (N_14833,N_14772,N_14711);
nand U14834 (N_14834,N_14681,N_14771);
xor U14835 (N_14835,N_14764,N_14649);
xor U14836 (N_14836,N_14703,N_14652);
and U14837 (N_14837,N_14659,N_14626);
xor U14838 (N_14838,N_14756,N_14668);
or U14839 (N_14839,N_14773,N_14647);
or U14840 (N_14840,N_14624,N_14692);
nand U14841 (N_14841,N_14644,N_14613);
and U14842 (N_14842,N_14621,N_14611);
and U14843 (N_14843,N_14602,N_14695);
xnor U14844 (N_14844,N_14708,N_14674);
xor U14845 (N_14845,N_14670,N_14776);
nand U14846 (N_14846,N_14702,N_14672);
xnor U14847 (N_14847,N_14751,N_14685);
or U14848 (N_14848,N_14782,N_14610);
nand U14849 (N_14849,N_14634,N_14698);
xnor U14850 (N_14850,N_14616,N_14731);
nor U14851 (N_14851,N_14683,N_14739);
and U14852 (N_14852,N_14798,N_14767);
and U14853 (N_14853,N_14637,N_14732);
nor U14854 (N_14854,N_14690,N_14655);
and U14855 (N_14855,N_14679,N_14678);
and U14856 (N_14856,N_14728,N_14738);
or U14857 (N_14857,N_14795,N_14704);
nand U14858 (N_14858,N_14712,N_14718);
xnor U14859 (N_14859,N_14757,N_14689);
nor U14860 (N_14860,N_14706,N_14746);
xnor U14861 (N_14861,N_14777,N_14651);
and U14862 (N_14862,N_14747,N_14716);
nand U14863 (N_14863,N_14743,N_14600);
and U14864 (N_14864,N_14641,N_14761);
nor U14865 (N_14865,N_14719,N_14605);
nand U14866 (N_14866,N_14629,N_14694);
xor U14867 (N_14867,N_14653,N_14628);
and U14868 (N_14868,N_14749,N_14759);
or U14869 (N_14869,N_14709,N_14723);
and U14870 (N_14870,N_14770,N_14680);
xor U14871 (N_14871,N_14646,N_14631);
and U14872 (N_14872,N_14769,N_14684);
or U14873 (N_14873,N_14791,N_14789);
or U14874 (N_14874,N_14790,N_14650);
or U14875 (N_14875,N_14778,N_14722);
and U14876 (N_14876,N_14768,N_14654);
nand U14877 (N_14877,N_14686,N_14786);
nor U14878 (N_14878,N_14687,N_14714);
nand U14879 (N_14879,N_14781,N_14693);
xnor U14880 (N_14880,N_14726,N_14645);
nor U14881 (N_14881,N_14760,N_14648);
nand U14882 (N_14882,N_14724,N_14707);
and U14883 (N_14883,N_14623,N_14720);
xor U14884 (N_14884,N_14763,N_14725);
xor U14885 (N_14885,N_14660,N_14615);
xor U14886 (N_14886,N_14699,N_14742);
nand U14887 (N_14887,N_14608,N_14606);
xor U14888 (N_14888,N_14632,N_14673);
nand U14889 (N_14889,N_14779,N_14700);
xnor U14890 (N_14890,N_14737,N_14741);
and U14891 (N_14891,N_14604,N_14784);
nand U14892 (N_14892,N_14663,N_14785);
nand U14893 (N_14893,N_14636,N_14657);
xor U14894 (N_14894,N_14671,N_14745);
or U14895 (N_14895,N_14688,N_14697);
or U14896 (N_14896,N_14750,N_14633);
or U14897 (N_14897,N_14607,N_14796);
and U14898 (N_14898,N_14766,N_14630);
xnor U14899 (N_14899,N_14642,N_14775);
nand U14900 (N_14900,N_14612,N_14799);
xor U14901 (N_14901,N_14648,N_14617);
or U14902 (N_14902,N_14624,N_14619);
or U14903 (N_14903,N_14793,N_14672);
nor U14904 (N_14904,N_14798,N_14796);
and U14905 (N_14905,N_14673,N_14777);
or U14906 (N_14906,N_14641,N_14787);
nor U14907 (N_14907,N_14793,N_14759);
nand U14908 (N_14908,N_14672,N_14733);
nand U14909 (N_14909,N_14750,N_14677);
xor U14910 (N_14910,N_14718,N_14797);
xor U14911 (N_14911,N_14616,N_14658);
or U14912 (N_14912,N_14781,N_14717);
nand U14913 (N_14913,N_14765,N_14612);
nand U14914 (N_14914,N_14692,N_14729);
and U14915 (N_14915,N_14668,N_14628);
and U14916 (N_14916,N_14703,N_14661);
nor U14917 (N_14917,N_14706,N_14741);
nor U14918 (N_14918,N_14797,N_14659);
or U14919 (N_14919,N_14610,N_14691);
or U14920 (N_14920,N_14762,N_14670);
and U14921 (N_14921,N_14649,N_14714);
and U14922 (N_14922,N_14755,N_14603);
nor U14923 (N_14923,N_14632,N_14764);
nand U14924 (N_14924,N_14725,N_14743);
and U14925 (N_14925,N_14707,N_14777);
nand U14926 (N_14926,N_14797,N_14668);
nand U14927 (N_14927,N_14668,N_14753);
or U14928 (N_14928,N_14698,N_14782);
xnor U14929 (N_14929,N_14602,N_14656);
or U14930 (N_14930,N_14796,N_14739);
or U14931 (N_14931,N_14761,N_14647);
nor U14932 (N_14932,N_14717,N_14665);
and U14933 (N_14933,N_14760,N_14749);
and U14934 (N_14934,N_14668,N_14687);
and U14935 (N_14935,N_14722,N_14730);
xor U14936 (N_14936,N_14774,N_14607);
and U14937 (N_14937,N_14742,N_14680);
or U14938 (N_14938,N_14660,N_14757);
nand U14939 (N_14939,N_14786,N_14607);
nand U14940 (N_14940,N_14727,N_14725);
and U14941 (N_14941,N_14636,N_14769);
xnor U14942 (N_14942,N_14792,N_14724);
nor U14943 (N_14943,N_14676,N_14767);
or U14944 (N_14944,N_14715,N_14743);
and U14945 (N_14945,N_14622,N_14766);
nand U14946 (N_14946,N_14655,N_14794);
and U14947 (N_14947,N_14716,N_14660);
nand U14948 (N_14948,N_14641,N_14609);
nor U14949 (N_14949,N_14606,N_14742);
or U14950 (N_14950,N_14646,N_14700);
nor U14951 (N_14951,N_14708,N_14764);
and U14952 (N_14952,N_14700,N_14760);
or U14953 (N_14953,N_14711,N_14743);
nor U14954 (N_14954,N_14680,N_14700);
nor U14955 (N_14955,N_14641,N_14639);
and U14956 (N_14956,N_14716,N_14642);
and U14957 (N_14957,N_14612,N_14766);
nand U14958 (N_14958,N_14650,N_14676);
or U14959 (N_14959,N_14735,N_14733);
and U14960 (N_14960,N_14788,N_14641);
xnor U14961 (N_14961,N_14703,N_14735);
nor U14962 (N_14962,N_14623,N_14702);
nand U14963 (N_14963,N_14660,N_14781);
and U14964 (N_14964,N_14783,N_14721);
nand U14965 (N_14965,N_14677,N_14650);
nor U14966 (N_14966,N_14603,N_14638);
nor U14967 (N_14967,N_14637,N_14739);
nand U14968 (N_14968,N_14708,N_14645);
or U14969 (N_14969,N_14608,N_14658);
or U14970 (N_14970,N_14613,N_14697);
nor U14971 (N_14971,N_14712,N_14787);
xnor U14972 (N_14972,N_14792,N_14756);
xor U14973 (N_14973,N_14682,N_14705);
or U14974 (N_14974,N_14651,N_14655);
and U14975 (N_14975,N_14760,N_14641);
or U14976 (N_14976,N_14654,N_14691);
nor U14977 (N_14977,N_14671,N_14787);
nand U14978 (N_14978,N_14631,N_14622);
nor U14979 (N_14979,N_14751,N_14616);
nor U14980 (N_14980,N_14724,N_14624);
xnor U14981 (N_14981,N_14709,N_14693);
or U14982 (N_14982,N_14711,N_14623);
xnor U14983 (N_14983,N_14779,N_14655);
or U14984 (N_14984,N_14617,N_14623);
or U14985 (N_14985,N_14625,N_14736);
nor U14986 (N_14986,N_14709,N_14784);
xor U14987 (N_14987,N_14619,N_14697);
xnor U14988 (N_14988,N_14602,N_14625);
or U14989 (N_14989,N_14734,N_14659);
nand U14990 (N_14990,N_14796,N_14705);
xor U14991 (N_14991,N_14739,N_14756);
nand U14992 (N_14992,N_14651,N_14630);
nor U14993 (N_14993,N_14617,N_14685);
or U14994 (N_14994,N_14728,N_14635);
and U14995 (N_14995,N_14796,N_14658);
nand U14996 (N_14996,N_14726,N_14650);
and U14997 (N_14997,N_14755,N_14799);
nand U14998 (N_14998,N_14722,N_14690);
xor U14999 (N_14999,N_14702,N_14610);
xnor U15000 (N_15000,N_14902,N_14912);
or U15001 (N_15001,N_14987,N_14857);
xnor U15002 (N_15002,N_14974,N_14855);
xor U15003 (N_15003,N_14964,N_14826);
xnor U15004 (N_15004,N_14913,N_14866);
or U15005 (N_15005,N_14877,N_14966);
and U15006 (N_15006,N_14963,N_14888);
xor U15007 (N_15007,N_14864,N_14889);
or U15008 (N_15008,N_14862,N_14839);
nor U15009 (N_15009,N_14805,N_14988);
xnor U15010 (N_15010,N_14978,N_14856);
xnor U15011 (N_15011,N_14882,N_14865);
or U15012 (N_15012,N_14835,N_14926);
and U15013 (N_15013,N_14897,N_14977);
nor U15014 (N_15014,N_14814,N_14983);
and U15015 (N_15015,N_14945,N_14917);
nand U15016 (N_15016,N_14810,N_14871);
nand U15017 (N_15017,N_14885,N_14954);
xor U15018 (N_15018,N_14895,N_14848);
nand U15019 (N_15019,N_14994,N_14904);
nor U15020 (N_15020,N_14903,N_14809);
xor U15021 (N_15021,N_14993,N_14928);
and U15022 (N_15022,N_14841,N_14822);
nor U15023 (N_15023,N_14853,N_14990);
or U15024 (N_15024,N_14803,N_14817);
or U15025 (N_15025,N_14875,N_14995);
nand U15026 (N_15026,N_14833,N_14965);
and U15027 (N_15027,N_14905,N_14976);
xor U15028 (N_15028,N_14956,N_14958);
or U15029 (N_15029,N_14953,N_14911);
xnor U15030 (N_15030,N_14929,N_14867);
nor U15031 (N_15031,N_14802,N_14896);
xor U15032 (N_15032,N_14812,N_14938);
xor U15033 (N_15033,N_14819,N_14872);
xor U15034 (N_15034,N_14942,N_14852);
nor U15035 (N_15035,N_14813,N_14947);
nor U15036 (N_15036,N_14861,N_14827);
nand U15037 (N_15037,N_14893,N_14891);
xnor U15038 (N_15038,N_14816,N_14957);
nor U15039 (N_15039,N_14967,N_14921);
xor U15040 (N_15040,N_14927,N_14836);
nand U15041 (N_15041,N_14894,N_14982);
nand U15042 (N_15042,N_14879,N_14899);
nor U15043 (N_15043,N_14869,N_14820);
xnor U15044 (N_15044,N_14834,N_14874);
xor U15045 (N_15045,N_14858,N_14860);
or U15046 (N_15046,N_14801,N_14919);
or U15047 (N_15047,N_14939,N_14969);
and U15048 (N_15048,N_14870,N_14946);
or U15049 (N_15049,N_14825,N_14811);
and U15050 (N_15050,N_14934,N_14881);
nand U15051 (N_15051,N_14842,N_14892);
nor U15052 (N_15052,N_14849,N_14924);
and U15053 (N_15053,N_14907,N_14806);
or U15054 (N_15054,N_14923,N_14951);
nand U15055 (N_15055,N_14961,N_14901);
or U15056 (N_15056,N_14937,N_14840);
nand U15057 (N_15057,N_14989,N_14886);
or U15058 (N_15058,N_14943,N_14930);
or U15059 (N_15059,N_14890,N_14854);
or U15060 (N_15060,N_14971,N_14979);
xor U15061 (N_15061,N_14916,N_14968);
nand U15062 (N_15062,N_14908,N_14910);
and U15063 (N_15063,N_14915,N_14804);
xnor U15064 (N_15064,N_14851,N_14876);
nor U15065 (N_15065,N_14973,N_14998);
nand U15066 (N_15066,N_14859,N_14838);
or U15067 (N_15067,N_14970,N_14996);
nand U15068 (N_15068,N_14863,N_14932);
nor U15069 (N_15069,N_14800,N_14823);
nor U15070 (N_15070,N_14944,N_14914);
or U15071 (N_15071,N_14940,N_14955);
nor U15072 (N_15072,N_14844,N_14878);
xor U15073 (N_15073,N_14984,N_14980);
or U15074 (N_15074,N_14985,N_14808);
nand U15075 (N_15075,N_14922,N_14935);
and U15076 (N_15076,N_14873,N_14846);
and U15077 (N_15077,N_14824,N_14959);
and U15078 (N_15078,N_14960,N_14936);
nor U15079 (N_15079,N_14900,N_14832);
xnor U15080 (N_15080,N_14952,N_14898);
or U15081 (N_15081,N_14883,N_14941);
nand U15082 (N_15082,N_14845,N_14818);
nand U15083 (N_15083,N_14847,N_14920);
nand U15084 (N_15084,N_14821,N_14837);
xor U15085 (N_15085,N_14828,N_14931);
or U15086 (N_15086,N_14992,N_14815);
or U15087 (N_15087,N_14925,N_14829);
nand U15088 (N_15088,N_14807,N_14831);
nor U15089 (N_15089,N_14949,N_14975);
xnor U15090 (N_15090,N_14950,N_14918);
and U15091 (N_15091,N_14986,N_14948);
xnor U15092 (N_15092,N_14962,N_14997);
nand U15093 (N_15093,N_14843,N_14880);
nor U15094 (N_15094,N_14909,N_14981);
or U15095 (N_15095,N_14830,N_14972);
and U15096 (N_15096,N_14933,N_14906);
xor U15097 (N_15097,N_14991,N_14999);
and U15098 (N_15098,N_14850,N_14868);
xor U15099 (N_15099,N_14887,N_14884);
xor U15100 (N_15100,N_14947,N_14835);
xnor U15101 (N_15101,N_14955,N_14841);
or U15102 (N_15102,N_14944,N_14814);
nand U15103 (N_15103,N_14820,N_14955);
xor U15104 (N_15104,N_14850,N_14820);
nand U15105 (N_15105,N_14957,N_14972);
or U15106 (N_15106,N_14848,N_14815);
xnor U15107 (N_15107,N_14866,N_14940);
nor U15108 (N_15108,N_14997,N_14884);
nor U15109 (N_15109,N_14957,N_14824);
xor U15110 (N_15110,N_14968,N_14870);
nand U15111 (N_15111,N_14845,N_14943);
and U15112 (N_15112,N_14813,N_14808);
nor U15113 (N_15113,N_14983,N_14839);
xor U15114 (N_15114,N_14993,N_14907);
nand U15115 (N_15115,N_14841,N_14979);
xnor U15116 (N_15116,N_14818,N_14867);
nor U15117 (N_15117,N_14884,N_14866);
nand U15118 (N_15118,N_14997,N_14874);
nand U15119 (N_15119,N_14860,N_14992);
nor U15120 (N_15120,N_14826,N_14912);
nor U15121 (N_15121,N_14964,N_14933);
or U15122 (N_15122,N_14931,N_14904);
nor U15123 (N_15123,N_14986,N_14960);
and U15124 (N_15124,N_14871,N_14867);
and U15125 (N_15125,N_14982,N_14969);
nor U15126 (N_15126,N_14813,N_14966);
nand U15127 (N_15127,N_14960,N_14932);
xor U15128 (N_15128,N_14914,N_14946);
and U15129 (N_15129,N_14905,N_14945);
and U15130 (N_15130,N_14854,N_14900);
nor U15131 (N_15131,N_14804,N_14942);
or U15132 (N_15132,N_14989,N_14927);
nand U15133 (N_15133,N_14862,N_14933);
nor U15134 (N_15134,N_14812,N_14993);
nand U15135 (N_15135,N_14814,N_14833);
and U15136 (N_15136,N_14850,N_14873);
and U15137 (N_15137,N_14922,N_14937);
nor U15138 (N_15138,N_14858,N_14837);
and U15139 (N_15139,N_14929,N_14923);
xnor U15140 (N_15140,N_14992,N_14806);
nand U15141 (N_15141,N_14852,N_14958);
or U15142 (N_15142,N_14895,N_14873);
xnor U15143 (N_15143,N_14938,N_14809);
nand U15144 (N_15144,N_14853,N_14813);
nand U15145 (N_15145,N_14843,N_14871);
and U15146 (N_15146,N_14903,N_14827);
nor U15147 (N_15147,N_14916,N_14896);
xnor U15148 (N_15148,N_14994,N_14848);
or U15149 (N_15149,N_14958,N_14871);
or U15150 (N_15150,N_14871,N_14935);
xor U15151 (N_15151,N_14805,N_14947);
xor U15152 (N_15152,N_14942,N_14875);
nand U15153 (N_15153,N_14900,N_14864);
and U15154 (N_15154,N_14885,N_14999);
or U15155 (N_15155,N_14925,N_14940);
xor U15156 (N_15156,N_14842,N_14870);
nand U15157 (N_15157,N_14853,N_14973);
xor U15158 (N_15158,N_14892,N_14976);
nand U15159 (N_15159,N_14817,N_14825);
nor U15160 (N_15160,N_14863,N_14853);
and U15161 (N_15161,N_14972,N_14979);
and U15162 (N_15162,N_14881,N_14828);
and U15163 (N_15163,N_14956,N_14808);
xor U15164 (N_15164,N_14975,N_14832);
and U15165 (N_15165,N_14851,N_14904);
nand U15166 (N_15166,N_14970,N_14966);
nor U15167 (N_15167,N_14987,N_14968);
nand U15168 (N_15168,N_14867,N_14859);
xnor U15169 (N_15169,N_14932,N_14970);
and U15170 (N_15170,N_14909,N_14985);
or U15171 (N_15171,N_14885,N_14946);
nor U15172 (N_15172,N_14854,N_14998);
or U15173 (N_15173,N_14807,N_14993);
nor U15174 (N_15174,N_14874,N_14842);
nor U15175 (N_15175,N_14995,N_14903);
nand U15176 (N_15176,N_14810,N_14936);
xnor U15177 (N_15177,N_14810,N_14873);
and U15178 (N_15178,N_14869,N_14948);
nand U15179 (N_15179,N_14944,N_14975);
xor U15180 (N_15180,N_14890,N_14982);
and U15181 (N_15181,N_14808,N_14914);
nand U15182 (N_15182,N_14977,N_14947);
nand U15183 (N_15183,N_14968,N_14929);
or U15184 (N_15184,N_14807,N_14977);
and U15185 (N_15185,N_14895,N_14953);
or U15186 (N_15186,N_14961,N_14950);
nand U15187 (N_15187,N_14939,N_14964);
xnor U15188 (N_15188,N_14985,N_14972);
nor U15189 (N_15189,N_14996,N_14817);
nand U15190 (N_15190,N_14871,N_14877);
nor U15191 (N_15191,N_14968,N_14873);
nor U15192 (N_15192,N_14873,N_14974);
or U15193 (N_15193,N_14982,N_14990);
nand U15194 (N_15194,N_14960,N_14970);
xnor U15195 (N_15195,N_14864,N_14926);
nor U15196 (N_15196,N_14980,N_14856);
or U15197 (N_15197,N_14925,N_14948);
xor U15198 (N_15198,N_14912,N_14891);
or U15199 (N_15199,N_14916,N_14821);
nand U15200 (N_15200,N_15096,N_15004);
xor U15201 (N_15201,N_15124,N_15119);
or U15202 (N_15202,N_15040,N_15121);
or U15203 (N_15203,N_15047,N_15136);
nor U15204 (N_15204,N_15101,N_15002);
xor U15205 (N_15205,N_15195,N_15060);
nand U15206 (N_15206,N_15090,N_15127);
nand U15207 (N_15207,N_15034,N_15068);
or U15208 (N_15208,N_15011,N_15022);
and U15209 (N_15209,N_15094,N_15151);
nand U15210 (N_15210,N_15044,N_15180);
xor U15211 (N_15211,N_15166,N_15141);
nand U15212 (N_15212,N_15118,N_15051);
or U15213 (N_15213,N_15065,N_15156);
nor U15214 (N_15214,N_15177,N_15008);
and U15215 (N_15215,N_15130,N_15145);
or U15216 (N_15216,N_15098,N_15185);
xnor U15217 (N_15217,N_15014,N_15125);
xnor U15218 (N_15218,N_15134,N_15062);
and U15219 (N_15219,N_15012,N_15153);
nand U15220 (N_15220,N_15021,N_15020);
xor U15221 (N_15221,N_15186,N_15128);
and U15222 (N_15222,N_15138,N_15099);
and U15223 (N_15223,N_15131,N_15042);
nand U15224 (N_15224,N_15078,N_15050);
nor U15225 (N_15225,N_15046,N_15126);
nor U15226 (N_15226,N_15073,N_15074);
nor U15227 (N_15227,N_15175,N_15188);
or U15228 (N_15228,N_15115,N_15059);
xnor U15229 (N_15229,N_15187,N_15033);
and U15230 (N_15230,N_15182,N_15026);
nor U15231 (N_15231,N_15140,N_15103);
xor U15232 (N_15232,N_15189,N_15089);
nand U15233 (N_15233,N_15108,N_15039);
or U15234 (N_15234,N_15066,N_15064);
xnor U15235 (N_15235,N_15072,N_15171);
and U15236 (N_15236,N_15067,N_15041);
and U15237 (N_15237,N_15017,N_15029);
nor U15238 (N_15238,N_15055,N_15163);
and U15239 (N_15239,N_15028,N_15015);
or U15240 (N_15240,N_15043,N_15117);
nor U15241 (N_15241,N_15025,N_15169);
nor U15242 (N_15242,N_15135,N_15174);
xor U15243 (N_15243,N_15173,N_15016);
nand U15244 (N_15244,N_15110,N_15152);
nand U15245 (N_15245,N_15018,N_15070);
and U15246 (N_15246,N_15196,N_15114);
xor U15247 (N_15247,N_15045,N_15161);
and U15248 (N_15248,N_15063,N_15023);
nor U15249 (N_15249,N_15193,N_15097);
nand U15250 (N_15250,N_15198,N_15107);
nand U15251 (N_15251,N_15076,N_15111);
or U15252 (N_15252,N_15058,N_15170);
xnor U15253 (N_15253,N_15092,N_15049);
xnor U15254 (N_15254,N_15071,N_15030);
or U15255 (N_15255,N_15184,N_15053);
nand U15256 (N_15256,N_15087,N_15143);
and U15257 (N_15257,N_15144,N_15150);
nand U15258 (N_15258,N_15149,N_15052);
nand U15259 (N_15259,N_15181,N_15165);
nand U15260 (N_15260,N_15048,N_15056);
or U15261 (N_15261,N_15199,N_15113);
xor U15262 (N_15262,N_15147,N_15035);
nor U15263 (N_15263,N_15183,N_15007);
or U15264 (N_15264,N_15102,N_15075);
and U15265 (N_15265,N_15061,N_15142);
nor U15266 (N_15266,N_15086,N_15027);
nor U15267 (N_15267,N_15088,N_15093);
nand U15268 (N_15268,N_15077,N_15024);
xnor U15269 (N_15269,N_15112,N_15000);
and U15270 (N_15270,N_15013,N_15083);
nor U15271 (N_15271,N_15148,N_15194);
nand U15272 (N_15272,N_15160,N_15105);
nor U15273 (N_15273,N_15095,N_15197);
xnor U15274 (N_15274,N_15085,N_15116);
xnor U15275 (N_15275,N_15154,N_15192);
nand U15276 (N_15276,N_15038,N_15120);
and U15277 (N_15277,N_15162,N_15158);
nand U15278 (N_15278,N_15132,N_15091);
and U15279 (N_15279,N_15005,N_15080);
nand U15280 (N_15280,N_15019,N_15009);
nor U15281 (N_15281,N_15032,N_15139);
or U15282 (N_15282,N_15100,N_15167);
and U15283 (N_15283,N_15146,N_15178);
nand U15284 (N_15284,N_15084,N_15010);
nand U15285 (N_15285,N_15109,N_15155);
nor U15286 (N_15286,N_15079,N_15179);
nor U15287 (N_15287,N_15057,N_15106);
nor U15288 (N_15288,N_15129,N_15172);
nor U15289 (N_15289,N_15168,N_15006);
nand U15290 (N_15290,N_15003,N_15176);
or U15291 (N_15291,N_15036,N_15037);
nand U15292 (N_15292,N_15104,N_15157);
or U15293 (N_15293,N_15001,N_15081);
nand U15294 (N_15294,N_15191,N_15159);
nand U15295 (N_15295,N_15031,N_15069);
nand U15296 (N_15296,N_15054,N_15137);
nor U15297 (N_15297,N_15123,N_15190);
or U15298 (N_15298,N_15164,N_15082);
nand U15299 (N_15299,N_15133,N_15122);
and U15300 (N_15300,N_15115,N_15138);
nor U15301 (N_15301,N_15101,N_15017);
nor U15302 (N_15302,N_15149,N_15144);
and U15303 (N_15303,N_15026,N_15113);
or U15304 (N_15304,N_15132,N_15166);
or U15305 (N_15305,N_15142,N_15055);
and U15306 (N_15306,N_15062,N_15169);
or U15307 (N_15307,N_15058,N_15012);
nand U15308 (N_15308,N_15053,N_15170);
xor U15309 (N_15309,N_15107,N_15169);
nor U15310 (N_15310,N_15143,N_15136);
nand U15311 (N_15311,N_15041,N_15184);
or U15312 (N_15312,N_15140,N_15188);
or U15313 (N_15313,N_15043,N_15103);
and U15314 (N_15314,N_15042,N_15111);
nand U15315 (N_15315,N_15153,N_15187);
nor U15316 (N_15316,N_15199,N_15003);
nand U15317 (N_15317,N_15116,N_15170);
nand U15318 (N_15318,N_15089,N_15115);
or U15319 (N_15319,N_15083,N_15113);
nand U15320 (N_15320,N_15198,N_15022);
nor U15321 (N_15321,N_15142,N_15003);
and U15322 (N_15322,N_15084,N_15055);
xnor U15323 (N_15323,N_15191,N_15178);
or U15324 (N_15324,N_15002,N_15065);
xnor U15325 (N_15325,N_15023,N_15025);
and U15326 (N_15326,N_15090,N_15110);
xor U15327 (N_15327,N_15079,N_15093);
and U15328 (N_15328,N_15140,N_15069);
and U15329 (N_15329,N_15073,N_15096);
nor U15330 (N_15330,N_15132,N_15156);
and U15331 (N_15331,N_15196,N_15040);
and U15332 (N_15332,N_15135,N_15145);
nor U15333 (N_15333,N_15013,N_15169);
and U15334 (N_15334,N_15184,N_15061);
and U15335 (N_15335,N_15079,N_15047);
and U15336 (N_15336,N_15044,N_15081);
and U15337 (N_15337,N_15007,N_15008);
or U15338 (N_15338,N_15138,N_15064);
nor U15339 (N_15339,N_15024,N_15197);
nand U15340 (N_15340,N_15083,N_15181);
and U15341 (N_15341,N_15130,N_15104);
nor U15342 (N_15342,N_15017,N_15067);
xnor U15343 (N_15343,N_15157,N_15012);
nor U15344 (N_15344,N_15081,N_15183);
nand U15345 (N_15345,N_15100,N_15000);
nand U15346 (N_15346,N_15025,N_15167);
nor U15347 (N_15347,N_15121,N_15056);
nand U15348 (N_15348,N_15119,N_15157);
and U15349 (N_15349,N_15075,N_15195);
nand U15350 (N_15350,N_15150,N_15118);
nor U15351 (N_15351,N_15044,N_15139);
xnor U15352 (N_15352,N_15166,N_15041);
xor U15353 (N_15353,N_15175,N_15103);
xor U15354 (N_15354,N_15196,N_15172);
or U15355 (N_15355,N_15152,N_15058);
nand U15356 (N_15356,N_15169,N_15196);
nand U15357 (N_15357,N_15062,N_15011);
nor U15358 (N_15358,N_15194,N_15046);
or U15359 (N_15359,N_15145,N_15092);
xor U15360 (N_15360,N_15158,N_15109);
and U15361 (N_15361,N_15151,N_15164);
and U15362 (N_15362,N_15189,N_15025);
nand U15363 (N_15363,N_15025,N_15066);
nor U15364 (N_15364,N_15045,N_15051);
xor U15365 (N_15365,N_15164,N_15167);
nand U15366 (N_15366,N_15131,N_15078);
and U15367 (N_15367,N_15062,N_15041);
nor U15368 (N_15368,N_15199,N_15097);
nand U15369 (N_15369,N_15095,N_15161);
nand U15370 (N_15370,N_15064,N_15148);
xnor U15371 (N_15371,N_15173,N_15109);
and U15372 (N_15372,N_15029,N_15144);
nor U15373 (N_15373,N_15005,N_15075);
and U15374 (N_15374,N_15195,N_15068);
xnor U15375 (N_15375,N_15196,N_15113);
or U15376 (N_15376,N_15198,N_15182);
nand U15377 (N_15377,N_15143,N_15015);
nor U15378 (N_15378,N_15068,N_15188);
nor U15379 (N_15379,N_15084,N_15082);
nand U15380 (N_15380,N_15050,N_15123);
xnor U15381 (N_15381,N_15150,N_15110);
nor U15382 (N_15382,N_15172,N_15071);
or U15383 (N_15383,N_15025,N_15139);
and U15384 (N_15384,N_15023,N_15122);
and U15385 (N_15385,N_15122,N_15060);
nand U15386 (N_15386,N_15135,N_15052);
xnor U15387 (N_15387,N_15062,N_15018);
and U15388 (N_15388,N_15101,N_15089);
nor U15389 (N_15389,N_15013,N_15060);
nor U15390 (N_15390,N_15164,N_15009);
xnor U15391 (N_15391,N_15118,N_15162);
and U15392 (N_15392,N_15037,N_15147);
nand U15393 (N_15393,N_15099,N_15001);
xnor U15394 (N_15394,N_15192,N_15126);
nand U15395 (N_15395,N_15006,N_15091);
and U15396 (N_15396,N_15052,N_15145);
or U15397 (N_15397,N_15041,N_15049);
or U15398 (N_15398,N_15188,N_15178);
nand U15399 (N_15399,N_15063,N_15188);
or U15400 (N_15400,N_15249,N_15283);
xnor U15401 (N_15401,N_15341,N_15284);
nor U15402 (N_15402,N_15395,N_15396);
nor U15403 (N_15403,N_15262,N_15296);
nor U15404 (N_15404,N_15242,N_15309);
nand U15405 (N_15405,N_15368,N_15329);
xnor U15406 (N_15406,N_15327,N_15220);
or U15407 (N_15407,N_15291,N_15274);
nor U15408 (N_15408,N_15356,N_15357);
xor U15409 (N_15409,N_15346,N_15218);
nand U15410 (N_15410,N_15264,N_15321);
nor U15411 (N_15411,N_15221,N_15393);
xnor U15412 (N_15412,N_15398,N_15281);
or U15413 (N_15413,N_15299,N_15317);
or U15414 (N_15414,N_15383,N_15207);
and U15415 (N_15415,N_15318,N_15371);
nand U15416 (N_15416,N_15211,N_15352);
nor U15417 (N_15417,N_15295,N_15366);
and U15418 (N_15418,N_15394,N_15263);
and U15419 (N_15419,N_15310,N_15345);
nand U15420 (N_15420,N_15201,N_15385);
and U15421 (N_15421,N_15333,N_15348);
nand U15422 (N_15422,N_15238,N_15322);
or U15423 (N_15423,N_15314,N_15256);
nor U15424 (N_15424,N_15257,N_15360);
nor U15425 (N_15425,N_15236,N_15223);
or U15426 (N_15426,N_15231,N_15292);
and U15427 (N_15427,N_15361,N_15278);
xor U15428 (N_15428,N_15212,N_15324);
xnor U15429 (N_15429,N_15229,N_15338);
and U15430 (N_15430,N_15247,N_15234);
or U15431 (N_15431,N_15239,N_15227);
nor U15432 (N_15432,N_15307,N_15344);
nand U15433 (N_15433,N_15378,N_15288);
nand U15434 (N_15434,N_15298,N_15267);
nor U15435 (N_15435,N_15392,N_15331);
or U15436 (N_15436,N_15230,N_15376);
nand U15437 (N_15437,N_15358,N_15266);
and U15438 (N_15438,N_15399,N_15273);
nor U15439 (N_15439,N_15232,N_15293);
or U15440 (N_15440,N_15387,N_15297);
nand U15441 (N_15441,N_15205,N_15347);
or U15442 (N_15442,N_15377,N_15258);
or U15443 (N_15443,N_15375,N_15384);
or U15444 (N_15444,N_15305,N_15332);
nor U15445 (N_15445,N_15233,N_15246);
nand U15446 (N_15446,N_15326,N_15235);
or U15447 (N_15447,N_15320,N_15355);
xnor U15448 (N_15448,N_15277,N_15379);
nor U15449 (N_15449,N_15214,N_15276);
nand U15450 (N_15450,N_15315,N_15272);
or U15451 (N_15451,N_15204,N_15328);
nand U15452 (N_15452,N_15271,N_15269);
nand U15453 (N_15453,N_15351,N_15353);
xor U15454 (N_15454,N_15254,N_15302);
nand U15455 (N_15455,N_15311,N_15280);
nor U15456 (N_15456,N_15365,N_15250);
or U15457 (N_15457,N_15381,N_15373);
or U15458 (N_15458,N_15364,N_15237);
nand U15459 (N_15459,N_15340,N_15286);
or U15460 (N_15460,N_15252,N_15335);
nor U15461 (N_15461,N_15251,N_15363);
nand U15462 (N_15462,N_15209,N_15316);
nand U15463 (N_15463,N_15337,N_15342);
xor U15464 (N_15464,N_15391,N_15388);
xor U15465 (N_15465,N_15215,N_15300);
xnor U15466 (N_15466,N_15369,N_15372);
nor U15467 (N_15467,N_15397,N_15200);
or U15468 (N_15468,N_15306,N_15248);
nor U15469 (N_15469,N_15268,N_15261);
xor U15470 (N_15470,N_15362,N_15343);
and U15471 (N_15471,N_15244,N_15301);
or U15472 (N_15472,N_15290,N_15228);
and U15473 (N_15473,N_15226,N_15224);
xnor U15474 (N_15474,N_15367,N_15203);
nor U15475 (N_15475,N_15217,N_15259);
and U15476 (N_15476,N_15336,N_15225);
or U15477 (N_15477,N_15279,N_15334);
xor U15478 (N_15478,N_15313,N_15202);
xor U15479 (N_15479,N_15308,N_15222);
xnor U15480 (N_15480,N_15282,N_15323);
and U15481 (N_15481,N_15339,N_15354);
and U15482 (N_15482,N_15260,N_15359);
xnor U15483 (N_15483,N_15219,N_15370);
or U15484 (N_15484,N_15304,N_15245);
nor U15485 (N_15485,N_15312,N_15255);
xnor U15486 (N_15486,N_15253,N_15275);
or U15487 (N_15487,N_15350,N_15382);
nand U15488 (N_15488,N_15289,N_15349);
nand U15489 (N_15489,N_15265,N_15389);
nand U15490 (N_15490,N_15325,N_15374);
or U15491 (N_15491,N_15330,N_15285);
and U15492 (N_15492,N_15390,N_15213);
or U15493 (N_15493,N_15319,N_15208);
and U15494 (N_15494,N_15241,N_15380);
xnor U15495 (N_15495,N_15240,N_15243);
or U15496 (N_15496,N_15270,N_15386);
nand U15497 (N_15497,N_15294,N_15206);
xor U15498 (N_15498,N_15216,N_15287);
nor U15499 (N_15499,N_15210,N_15303);
and U15500 (N_15500,N_15251,N_15392);
or U15501 (N_15501,N_15351,N_15258);
and U15502 (N_15502,N_15393,N_15321);
nor U15503 (N_15503,N_15276,N_15374);
and U15504 (N_15504,N_15282,N_15264);
nand U15505 (N_15505,N_15258,N_15386);
nand U15506 (N_15506,N_15345,N_15356);
nor U15507 (N_15507,N_15343,N_15254);
nor U15508 (N_15508,N_15339,N_15394);
and U15509 (N_15509,N_15260,N_15335);
nand U15510 (N_15510,N_15324,N_15220);
xnor U15511 (N_15511,N_15347,N_15365);
and U15512 (N_15512,N_15331,N_15397);
nor U15513 (N_15513,N_15224,N_15251);
and U15514 (N_15514,N_15224,N_15210);
and U15515 (N_15515,N_15207,N_15220);
nor U15516 (N_15516,N_15360,N_15292);
and U15517 (N_15517,N_15300,N_15206);
nor U15518 (N_15518,N_15276,N_15360);
nor U15519 (N_15519,N_15255,N_15347);
nor U15520 (N_15520,N_15328,N_15353);
xor U15521 (N_15521,N_15283,N_15387);
nor U15522 (N_15522,N_15348,N_15328);
and U15523 (N_15523,N_15214,N_15268);
nand U15524 (N_15524,N_15214,N_15267);
and U15525 (N_15525,N_15338,N_15288);
nand U15526 (N_15526,N_15232,N_15306);
and U15527 (N_15527,N_15299,N_15351);
xnor U15528 (N_15528,N_15381,N_15217);
xnor U15529 (N_15529,N_15355,N_15252);
or U15530 (N_15530,N_15355,N_15214);
xnor U15531 (N_15531,N_15387,N_15284);
and U15532 (N_15532,N_15307,N_15304);
or U15533 (N_15533,N_15379,N_15340);
xor U15534 (N_15534,N_15278,N_15398);
nor U15535 (N_15535,N_15306,N_15280);
xnor U15536 (N_15536,N_15294,N_15208);
nand U15537 (N_15537,N_15326,N_15391);
and U15538 (N_15538,N_15203,N_15312);
xnor U15539 (N_15539,N_15249,N_15377);
or U15540 (N_15540,N_15374,N_15360);
xor U15541 (N_15541,N_15323,N_15356);
or U15542 (N_15542,N_15327,N_15227);
nor U15543 (N_15543,N_15250,N_15338);
nand U15544 (N_15544,N_15354,N_15246);
and U15545 (N_15545,N_15290,N_15356);
xnor U15546 (N_15546,N_15238,N_15391);
or U15547 (N_15547,N_15380,N_15266);
nor U15548 (N_15548,N_15347,N_15305);
xor U15549 (N_15549,N_15370,N_15244);
xor U15550 (N_15550,N_15251,N_15384);
xnor U15551 (N_15551,N_15271,N_15204);
xnor U15552 (N_15552,N_15340,N_15378);
nor U15553 (N_15553,N_15353,N_15235);
xnor U15554 (N_15554,N_15393,N_15341);
or U15555 (N_15555,N_15371,N_15335);
and U15556 (N_15556,N_15251,N_15212);
nor U15557 (N_15557,N_15389,N_15281);
nand U15558 (N_15558,N_15219,N_15337);
nor U15559 (N_15559,N_15240,N_15353);
and U15560 (N_15560,N_15284,N_15370);
or U15561 (N_15561,N_15339,N_15330);
and U15562 (N_15562,N_15397,N_15271);
xor U15563 (N_15563,N_15278,N_15362);
and U15564 (N_15564,N_15316,N_15315);
or U15565 (N_15565,N_15317,N_15397);
nand U15566 (N_15566,N_15394,N_15364);
xnor U15567 (N_15567,N_15364,N_15339);
or U15568 (N_15568,N_15208,N_15248);
and U15569 (N_15569,N_15374,N_15317);
or U15570 (N_15570,N_15332,N_15259);
nor U15571 (N_15571,N_15264,N_15240);
nor U15572 (N_15572,N_15222,N_15312);
or U15573 (N_15573,N_15285,N_15202);
nand U15574 (N_15574,N_15361,N_15207);
nor U15575 (N_15575,N_15234,N_15204);
nor U15576 (N_15576,N_15241,N_15245);
nor U15577 (N_15577,N_15301,N_15313);
or U15578 (N_15578,N_15222,N_15366);
and U15579 (N_15579,N_15355,N_15399);
nand U15580 (N_15580,N_15233,N_15284);
xor U15581 (N_15581,N_15327,N_15346);
and U15582 (N_15582,N_15282,N_15204);
and U15583 (N_15583,N_15299,N_15344);
nand U15584 (N_15584,N_15211,N_15285);
or U15585 (N_15585,N_15260,N_15215);
and U15586 (N_15586,N_15215,N_15270);
nand U15587 (N_15587,N_15222,N_15272);
or U15588 (N_15588,N_15393,N_15355);
nand U15589 (N_15589,N_15375,N_15395);
nor U15590 (N_15590,N_15384,N_15270);
nand U15591 (N_15591,N_15262,N_15211);
or U15592 (N_15592,N_15301,N_15304);
and U15593 (N_15593,N_15284,N_15354);
nor U15594 (N_15594,N_15321,N_15244);
nand U15595 (N_15595,N_15257,N_15314);
nor U15596 (N_15596,N_15254,N_15347);
xor U15597 (N_15597,N_15207,N_15310);
nor U15598 (N_15598,N_15265,N_15320);
nand U15599 (N_15599,N_15261,N_15270);
and U15600 (N_15600,N_15502,N_15441);
and U15601 (N_15601,N_15509,N_15526);
and U15602 (N_15602,N_15530,N_15405);
or U15603 (N_15603,N_15587,N_15543);
and U15604 (N_15604,N_15552,N_15581);
and U15605 (N_15605,N_15589,N_15419);
xor U15606 (N_15606,N_15445,N_15482);
and U15607 (N_15607,N_15454,N_15439);
nand U15608 (N_15608,N_15472,N_15418);
nor U15609 (N_15609,N_15555,N_15432);
or U15610 (N_15610,N_15546,N_15446);
or U15611 (N_15611,N_15513,N_15485);
xnor U15612 (N_15612,N_15506,N_15515);
and U15613 (N_15613,N_15544,N_15548);
nand U15614 (N_15614,N_15593,N_15427);
nand U15615 (N_15615,N_15471,N_15475);
and U15616 (N_15616,N_15499,N_15573);
or U15617 (N_15617,N_15578,N_15560);
and U15618 (N_15618,N_15430,N_15551);
nor U15619 (N_15619,N_15508,N_15425);
nand U15620 (N_15620,N_15411,N_15413);
and U15621 (N_15621,N_15568,N_15580);
nor U15622 (N_15622,N_15459,N_15461);
and U15623 (N_15623,N_15534,N_15494);
nand U15624 (N_15624,N_15422,N_15400);
xor U15625 (N_15625,N_15433,N_15582);
nor U15626 (N_15626,N_15599,N_15462);
nand U15627 (N_15627,N_15493,N_15442);
xnor U15628 (N_15628,N_15496,N_15570);
or U15629 (N_15629,N_15504,N_15529);
nand U15630 (N_15630,N_15539,N_15436);
and U15631 (N_15631,N_15596,N_15401);
xnor U15632 (N_15632,N_15557,N_15501);
or U15633 (N_15633,N_15595,N_15484);
and U15634 (N_15634,N_15524,N_15554);
and U15635 (N_15635,N_15594,N_15576);
nor U15636 (N_15636,N_15406,N_15473);
nor U15637 (N_15637,N_15412,N_15518);
or U15638 (N_15638,N_15498,N_15465);
and U15639 (N_15639,N_15572,N_15592);
xor U15640 (N_15640,N_15451,N_15503);
nor U15641 (N_15641,N_15480,N_15569);
nand U15642 (N_15642,N_15564,N_15512);
nand U15643 (N_15643,N_15495,N_15416);
xnor U15644 (N_15644,N_15466,N_15567);
or U15645 (N_15645,N_15542,N_15457);
and U15646 (N_15646,N_15490,N_15553);
nor U15647 (N_15647,N_15467,N_15532);
xor U15648 (N_15648,N_15558,N_15559);
nor U15649 (N_15649,N_15545,N_15478);
nor U15650 (N_15650,N_15528,N_15491);
and U15651 (N_15651,N_15577,N_15426);
or U15652 (N_15652,N_15453,N_15511);
and U15653 (N_15653,N_15510,N_15417);
xor U15654 (N_15654,N_15431,N_15468);
and U15655 (N_15655,N_15523,N_15520);
and U15656 (N_15656,N_15438,N_15541);
and U15657 (N_15657,N_15540,N_15410);
nor U15658 (N_15658,N_15421,N_15415);
nand U15659 (N_15659,N_15483,N_15420);
nand U15660 (N_15660,N_15481,N_15550);
or U15661 (N_15661,N_15447,N_15458);
xnor U15662 (N_15662,N_15574,N_15562);
nor U15663 (N_15663,N_15460,N_15590);
xnor U15664 (N_15664,N_15437,N_15561);
or U15665 (N_15665,N_15448,N_15584);
or U15666 (N_15666,N_15579,N_15571);
xor U15667 (N_15667,N_15474,N_15414);
or U15668 (N_15668,N_15455,N_15538);
nand U15669 (N_15669,N_15535,N_15549);
xnor U15670 (N_15670,N_15440,N_15450);
xor U15671 (N_15671,N_15507,N_15519);
xor U15672 (N_15672,N_15521,N_15497);
nand U15673 (N_15673,N_15452,N_15443);
nand U15674 (N_15674,N_15464,N_15566);
and U15675 (N_15675,N_15522,N_15423);
nor U15676 (N_15676,N_15489,N_15597);
xor U15677 (N_15677,N_15403,N_15429);
and U15678 (N_15678,N_15531,N_15476);
xnor U15679 (N_15679,N_15424,N_15586);
xor U15680 (N_15680,N_15463,N_15525);
nand U15681 (N_15681,N_15547,N_15449);
nand U15682 (N_15682,N_15428,N_15407);
nand U15683 (N_15683,N_15435,N_15598);
nand U15684 (N_15684,N_15556,N_15434);
nor U15685 (N_15685,N_15575,N_15500);
nand U15686 (N_15686,N_15487,N_15563);
nand U15687 (N_15687,N_15565,N_15477);
and U15688 (N_15688,N_15470,N_15479);
nor U15689 (N_15689,N_15527,N_15591);
or U15690 (N_15690,N_15537,N_15536);
and U15691 (N_15691,N_15588,N_15488);
and U15692 (N_15692,N_15444,N_15516);
and U15693 (N_15693,N_15408,N_15469);
nand U15694 (N_15694,N_15409,N_15492);
nand U15695 (N_15695,N_15514,N_15585);
nand U15696 (N_15696,N_15402,N_15533);
nor U15697 (N_15697,N_15583,N_15517);
nand U15698 (N_15698,N_15486,N_15456);
and U15699 (N_15699,N_15404,N_15505);
nor U15700 (N_15700,N_15407,N_15412);
nor U15701 (N_15701,N_15599,N_15597);
nand U15702 (N_15702,N_15473,N_15421);
nand U15703 (N_15703,N_15450,N_15484);
nor U15704 (N_15704,N_15565,N_15512);
nor U15705 (N_15705,N_15457,N_15469);
and U15706 (N_15706,N_15406,N_15430);
nor U15707 (N_15707,N_15432,N_15488);
or U15708 (N_15708,N_15475,N_15479);
nor U15709 (N_15709,N_15460,N_15474);
xnor U15710 (N_15710,N_15499,N_15535);
nand U15711 (N_15711,N_15444,N_15474);
nor U15712 (N_15712,N_15455,N_15522);
or U15713 (N_15713,N_15501,N_15593);
and U15714 (N_15714,N_15593,N_15470);
or U15715 (N_15715,N_15580,N_15481);
xnor U15716 (N_15716,N_15538,N_15563);
and U15717 (N_15717,N_15516,N_15547);
xor U15718 (N_15718,N_15579,N_15534);
xor U15719 (N_15719,N_15522,N_15469);
nand U15720 (N_15720,N_15594,N_15559);
nor U15721 (N_15721,N_15502,N_15545);
xor U15722 (N_15722,N_15595,N_15439);
xnor U15723 (N_15723,N_15575,N_15518);
or U15724 (N_15724,N_15420,N_15468);
or U15725 (N_15725,N_15549,N_15529);
nand U15726 (N_15726,N_15499,N_15473);
xnor U15727 (N_15727,N_15510,N_15532);
nand U15728 (N_15728,N_15458,N_15421);
nor U15729 (N_15729,N_15577,N_15566);
xor U15730 (N_15730,N_15599,N_15520);
nand U15731 (N_15731,N_15469,N_15433);
xnor U15732 (N_15732,N_15572,N_15509);
xor U15733 (N_15733,N_15440,N_15595);
or U15734 (N_15734,N_15413,N_15502);
or U15735 (N_15735,N_15478,N_15526);
xnor U15736 (N_15736,N_15486,N_15595);
nand U15737 (N_15737,N_15485,N_15584);
nor U15738 (N_15738,N_15407,N_15524);
xor U15739 (N_15739,N_15417,N_15441);
xor U15740 (N_15740,N_15409,N_15581);
and U15741 (N_15741,N_15465,N_15556);
and U15742 (N_15742,N_15565,N_15465);
or U15743 (N_15743,N_15414,N_15453);
nor U15744 (N_15744,N_15413,N_15520);
nand U15745 (N_15745,N_15500,N_15573);
nor U15746 (N_15746,N_15405,N_15518);
nor U15747 (N_15747,N_15561,N_15471);
or U15748 (N_15748,N_15539,N_15407);
or U15749 (N_15749,N_15596,N_15459);
or U15750 (N_15750,N_15567,N_15513);
or U15751 (N_15751,N_15541,N_15513);
nor U15752 (N_15752,N_15507,N_15586);
or U15753 (N_15753,N_15599,N_15594);
or U15754 (N_15754,N_15497,N_15593);
or U15755 (N_15755,N_15584,N_15431);
nand U15756 (N_15756,N_15449,N_15537);
and U15757 (N_15757,N_15491,N_15518);
xnor U15758 (N_15758,N_15462,N_15408);
nand U15759 (N_15759,N_15524,N_15501);
nor U15760 (N_15760,N_15441,N_15468);
and U15761 (N_15761,N_15553,N_15465);
xnor U15762 (N_15762,N_15452,N_15563);
nand U15763 (N_15763,N_15440,N_15438);
nand U15764 (N_15764,N_15482,N_15417);
nor U15765 (N_15765,N_15443,N_15460);
or U15766 (N_15766,N_15529,N_15514);
nor U15767 (N_15767,N_15461,N_15577);
xnor U15768 (N_15768,N_15551,N_15528);
xnor U15769 (N_15769,N_15441,N_15497);
and U15770 (N_15770,N_15583,N_15549);
or U15771 (N_15771,N_15491,N_15542);
nor U15772 (N_15772,N_15499,N_15434);
or U15773 (N_15773,N_15400,N_15489);
nand U15774 (N_15774,N_15529,N_15423);
xor U15775 (N_15775,N_15550,N_15484);
nand U15776 (N_15776,N_15546,N_15575);
xnor U15777 (N_15777,N_15469,N_15539);
nor U15778 (N_15778,N_15426,N_15406);
xor U15779 (N_15779,N_15499,N_15590);
or U15780 (N_15780,N_15498,N_15494);
and U15781 (N_15781,N_15486,N_15585);
xnor U15782 (N_15782,N_15510,N_15453);
nor U15783 (N_15783,N_15543,N_15561);
xor U15784 (N_15784,N_15446,N_15459);
nor U15785 (N_15785,N_15473,N_15460);
xor U15786 (N_15786,N_15493,N_15502);
xor U15787 (N_15787,N_15451,N_15464);
nor U15788 (N_15788,N_15581,N_15456);
xor U15789 (N_15789,N_15475,N_15484);
nor U15790 (N_15790,N_15595,N_15523);
nor U15791 (N_15791,N_15498,N_15482);
or U15792 (N_15792,N_15414,N_15554);
nand U15793 (N_15793,N_15535,N_15539);
nor U15794 (N_15794,N_15500,N_15556);
or U15795 (N_15795,N_15461,N_15442);
and U15796 (N_15796,N_15406,N_15515);
nor U15797 (N_15797,N_15435,N_15561);
nor U15798 (N_15798,N_15411,N_15573);
nand U15799 (N_15799,N_15577,N_15516);
nand U15800 (N_15800,N_15677,N_15699);
and U15801 (N_15801,N_15692,N_15682);
nor U15802 (N_15802,N_15757,N_15602);
nor U15803 (N_15803,N_15774,N_15724);
or U15804 (N_15804,N_15672,N_15663);
or U15805 (N_15805,N_15645,N_15646);
and U15806 (N_15806,N_15714,N_15786);
nor U15807 (N_15807,N_15615,N_15641);
and U15808 (N_15808,N_15756,N_15633);
nor U15809 (N_15809,N_15752,N_15632);
nand U15810 (N_15810,N_15618,N_15640);
nand U15811 (N_15811,N_15785,N_15768);
and U15812 (N_15812,N_15755,N_15629);
nor U15813 (N_15813,N_15654,N_15762);
and U15814 (N_15814,N_15731,N_15607);
and U15815 (N_15815,N_15653,N_15691);
or U15816 (N_15816,N_15792,N_15675);
or U15817 (N_15817,N_15773,N_15760);
nand U15818 (N_15818,N_15716,N_15642);
and U15819 (N_15819,N_15687,N_15670);
and U15820 (N_15820,N_15729,N_15624);
and U15821 (N_15821,N_15651,N_15637);
xnor U15822 (N_15822,N_15693,N_15736);
nand U15823 (N_15823,N_15620,N_15779);
xor U15824 (N_15824,N_15643,N_15659);
xnor U15825 (N_15825,N_15656,N_15744);
and U15826 (N_15826,N_15746,N_15770);
or U15827 (N_15827,N_15648,N_15668);
nor U15828 (N_15828,N_15621,N_15715);
xnor U15829 (N_15829,N_15669,N_15718);
or U15830 (N_15830,N_15733,N_15644);
and U15831 (N_15831,N_15685,N_15696);
or U15832 (N_15832,N_15676,N_15743);
xnor U15833 (N_15833,N_15769,N_15761);
nand U15834 (N_15834,N_15612,N_15679);
and U15835 (N_15835,N_15666,N_15738);
nor U15836 (N_15836,N_15741,N_15662);
nand U15837 (N_15837,N_15690,N_15793);
and U15838 (N_15838,N_15778,N_15630);
nor U15839 (N_15839,N_15706,N_15652);
nand U15840 (N_15840,N_15781,N_15712);
xor U15841 (N_15841,N_15775,N_15657);
or U15842 (N_15842,N_15728,N_15771);
xor U15843 (N_15843,N_15742,N_15732);
xnor U15844 (N_15844,N_15754,N_15745);
nor U15845 (N_15845,N_15725,N_15739);
and U15846 (N_15846,N_15636,N_15625);
and U15847 (N_15847,N_15703,N_15787);
xor U15848 (N_15848,N_15681,N_15611);
xnor U15849 (N_15849,N_15776,N_15616);
xnor U15850 (N_15850,N_15711,N_15795);
and U15851 (N_15851,N_15638,N_15766);
xor U15852 (N_15852,N_15680,N_15608);
or U15853 (N_15853,N_15710,N_15717);
nor U15854 (N_15854,N_15601,N_15713);
and U15855 (N_15855,N_15763,N_15609);
or U15856 (N_15856,N_15667,N_15772);
and U15857 (N_15857,N_15619,N_15758);
and U15858 (N_15858,N_15721,N_15723);
xor U15859 (N_15859,N_15683,N_15617);
nand U15860 (N_15860,N_15777,N_15689);
and U15861 (N_15861,N_15797,N_15765);
and U15862 (N_15862,N_15694,N_15665);
nor U15863 (N_15863,N_15791,N_15798);
nand U15864 (N_15864,N_15658,N_15720);
nor U15865 (N_15865,N_15708,N_15719);
nor U15866 (N_15866,N_15734,N_15631);
nor U15867 (N_15867,N_15671,N_15614);
or U15868 (N_15868,N_15790,N_15759);
nand U15869 (N_15869,N_15622,N_15784);
or U15870 (N_15870,N_15606,N_15749);
nand U15871 (N_15871,N_15722,N_15688);
nand U15872 (N_15872,N_15647,N_15750);
nor U15873 (N_15873,N_15788,N_15605);
nor U15874 (N_15874,N_15735,N_15664);
nor U15875 (N_15875,N_15639,N_15780);
or U15876 (N_15876,N_15610,N_15730);
and U15877 (N_15877,N_15709,N_15678);
nor U15878 (N_15878,N_15697,N_15655);
or U15879 (N_15879,N_15623,N_15661);
and U15880 (N_15880,N_15747,N_15674);
or U15881 (N_15881,N_15628,N_15799);
and U15882 (N_15882,N_15695,N_15740);
xnor U15883 (N_15883,N_15783,N_15673);
and U15884 (N_15884,N_15634,N_15737);
xor U15885 (N_15885,N_15726,N_15702);
nand U15886 (N_15886,N_15660,N_15764);
nor U15887 (N_15887,N_15686,N_15794);
nand U15888 (N_15888,N_15707,N_15796);
nor U15889 (N_15889,N_15705,N_15635);
and U15890 (N_15890,N_15704,N_15700);
and U15891 (N_15891,N_15626,N_15753);
xor U15892 (N_15892,N_15748,N_15650);
and U15893 (N_15893,N_15698,N_15603);
xnor U15894 (N_15894,N_15604,N_15782);
and U15895 (N_15895,N_15600,N_15627);
or U15896 (N_15896,N_15789,N_15701);
xnor U15897 (N_15897,N_15751,N_15613);
or U15898 (N_15898,N_15684,N_15649);
xor U15899 (N_15899,N_15727,N_15767);
xor U15900 (N_15900,N_15671,N_15691);
and U15901 (N_15901,N_15765,N_15680);
or U15902 (N_15902,N_15778,N_15615);
nand U15903 (N_15903,N_15707,N_15765);
and U15904 (N_15904,N_15697,N_15783);
nor U15905 (N_15905,N_15606,N_15798);
or U15906 (N_15906,N_15759,N_15797);
and U15907 (N_15907,N_15774,N_15746);
and U15908 (N_15908,N_15731,N_15682);
nor U15909 (N_15909,N_15653,N_15749);
nand U15910 (N_15910,N_15631,N_15618);
and U15911 (N_15911,N_15799,N_15794);
xor U15912 (N_15912,N_15775,N_15642);
or U15913 (N_15913,N_15699,N_15779);
or U15914 (N_15914,N_15629,N_15738);
nor U15915 (N_15915,N_15752,N_15613);
and U15916 (N_15916,N_15611,N_15634);
xor U15917 (N_15917,N_15661,N_15635);
or U15918 (N_15918,N_15795,N_15745);
and U15919 (N_15919,N_15776,N_15684);
nand U15920 (N_15920,N_15720,N_15668);
and U15921 (N_15921,N_15690,N_15698);
and U15922 (N_15922,N_15725,N_15769);
nor U15923 (N_15923,N_15672,N_15766);
and U15924 (N_15924,N_15685,N_15675);
xor U15925 (N_15925,N_15626,N_15655);
nand U15926 (N_15926,N_15787,N_15689);
and U15927 (N_15927,N_15690,N_15689);
nand U15928 (N_15928,N_15727,N_15779);
or U15929 (N_15929,N_15617,N_15704);
xor U15930 (N_15930,N_15749,N_15604);
xnor U15931 (N_15931,N_15600,N_15661);
xnor U15932 (N_15932,N_15734,N_15781);
xor U15933 (N_15933,N_15726,N_15650);
nor U15934 (N_15934,N_15765,N_15644);
and U15935 (N_15935,N_15680,N_15700);
nor U15936 (N_15936,N_15640,N_15796);
nand U15937 (N_15937,N_15767,N_15687);
xnor U15938 (N_15938,N_15731,N_15662);
and U15939 (N_15939,N_15659,N_15740);
nand U15940 (N_15940,N_15691,N_15769);
xnor U15941 (N_15941,N_15613,N_15764);
nand U15942 (N_15942,N_15687,N_15791);
nand U15943 (N_15943,N_15685,N_15726);
and U15944 (N_15944,N_15614,N_15638);
xor U15945 (N_15945,N_15613,N_15682);
and U15946 (N_15946,N_15662,N_15733);
nand U15947 (N_15947,N_15775,N_15764);
and U15948 (N_15948,N_15784,N_15791);
and U15949 (N_15949,N_15617,N_15769);
and U15950 (N_15950,N_15699,N_15749);
or U15951 (N_15951,N_15744,N_15668);
and U15952 (N_15952,N_15699,N_15607);
and U15953 (N_15953,N_15617,N_15783);
xnor U15954 (N_15954,N_15652,N_15704);
and U15955 (N_15955,N_15685,N_15653);
nor U15956 (N_15956,N_15638,N_15761);
or U15957 (N_15957,N_15613,N_15648);
and U15958 (N_15958,N_15640,N_15701);
or U15959 (N_15959,N_15668,N_15673);
and U15960 (N_15960,N_15786,N_15638);
and U15961 (N_15961,N_15703,N_15737);
nor U15962 (N_15962,N_15794,N_15783);
and U15963 (N_15963,N_15732,N_15785);
xor U15964 (N_15964,N_15745,N_15611);
nand U15965 (N_15965,N_15654,N_15658);
nand U15966 (N_15966,N_15774,N_15743);
xnor U15967 (N_15967,N_15654,N_15623);
and U15968 (N_15968,N_15673,N_15726);
nor U15969 (N_15969,N_15633,N_15695);
xnor U15970 (N_15970,N_15625,N_15761);
xnor U15971 (N_15971,N_15600,N_15789);
xnor U15972 (N_15972,N_15668,N_15660);
nor U15973 (N_15973,N_15633,N_15690);
nor U15974 (N_15974,N_15724,N_15753);
or U15975 (N_15975,N_15795,N_15788);
and U15976 (N_15976,N_15762,N_15739);
xnor U15977 (N_15977,N_15726,N_15789);
and U15978 (N_15978,N_15736,N_15755);
xor U15979 (N_15979,N_15630,N_15632);
and U15980 (N_15980,N_15630,N_15722);
xor U15981 (N_15981,N_15794,N_15630);
xnor U15982 (N_15982,N_15685,N_15757);
and U15983 (N_15983,N_15640,N_15655);
nand U15984 (N_15984,N_15756,N_15668);
and U15985 (N_15985,N_15799,N_15781);
xor U15986 (N_15986,N_15766,N_15721);
nor U15987 (N_15987,N_15784,N_15730);
xor U15988 (N_15988,N_15712,N_15676);
or U15989 (N_15989,N_15775,N_15612);
nor U15990 (N_15990,N_15646,N_15773);
and U15991 (N_15991,N_15659,N_15749);
nor U15992 (N_15992,N_15670,N_15726);
and U15993 (N_15993,N_15711,N_15671);
nor U15994 (N_15994,N_15674,N_15639);
nand U15995 (N_15995,N_15644,N_15778);
or U15996 (N_15996,N_15670,N_15739);
and U15997 (N_15997,N_15655,N_15791);
and U15998 (N_15998,N_15647,N_15783);
xnor U15999 (N_15999,N_15600,N_15691);
nor U16000 (N_16000,N_15955,N_15812);
nor U16001 (N_16001,N_15819,N_15885);
or U16002 (N_16002,N_15987,N_15805);
or U16003 (N_16003,N_15869,N_15863);
nand U16004 (N_16004,N_15892,N_15998);
or U16005 (N_16005,N_15963,N_15836);
nor U16006 (N_16006,N_15801,N_15803);
and U16007 (N_16007,N_15938,N_15996);
nand U16008 (N_16008,N_15886,N_15920);
and U16009 (N_16009,N_15860,N_15903);
nand U16010 (N_16010,N_15983,N_15932);
and U16011 (N_16011,N_15808,N_15951);
xnor U16012 (N_16012,N_15807,N_15917);
or U16013 (N_16013,N_15981,N_15929);
nor U16014 (N_16014,N_15939,N_15913);
xnor U16015 (N_16015,N_15935,N_15834);
nor U16016 (N_16016,N_15873,N_15979);
nand U16017 (N_16017,N_15990,N_15956);
and U16018 (N_16018,N_15916,N_15844);
nor U16019 (N_16019,N_15957,N_15822);
or U16020 (N_16020,N_15893,N_15891);
nor U16021 (N_16021,N_15927,N_15904);
and U16022 (N_16022,N_15937,N_15806);
xnor U16023 (N_16023,N_15861,N_15969);
nand U16024 (N_16024,N_15989,N_15868);
nand U16025 (N_16025,N_15826,N_15974);
or U16026 (N_16026,N_15879,N_15889);
xor U16027 (N_16027,N_15881,N_15850);
or U16028 (N_16028,N_15887,N_15942);
nor U16029 (N_16029,N_15899,N_15906);
nor U16030 (N_16030,N_15967,N_15975);
and U16031 (N_16031,N_15950,N_15962);
nand U16032 (N_16032,N_15818,N_15872);
xnor U16033 (N_16033,N_15866,N_15945);
nand U16034 (N_16034,N_15800,N_15825);
and U16035 (N_16035,N_15852,N_15809);
xnor U16036 (N_16036,N_15926,N_15854);
nand U16037 (N_16037,N_15995,N_15882);
and U16038 (N_16038,N_15851,N_15925);
nor U16039 (N_16039,N_15859,N_15977);
nor U16040 (N_16040,N_15833,N_15862);
nand U16041 (N_16041,N_15943,N_15933);
xnor U16042 (N_16042,N_15849,N_15839);
nor U16043 (N_16043,N_15960,N_15911);
or U16044 (N_16044,N_15948,N_15972);
nand U16045 (N_16045,N_15940,N_15853);
or U16046 (N_16046,N_15930,N_15986);
or U16047 (N_16047,N_15902,N_15824);
nor U16048 (N_16048,N_15910,N_15894);
or U16049 (N_16049,N_15867,N_15923);
xnor U16050 (N_16050,N_15876,N_15842);
nand U16051 (N_16051,N_15877,N_15829);
xor U16052 (N_16052,N_15810,N_15835);
xor U16053 (N_16053,N_15890,N_15814);
and U16054 (N_16054,N_15924,N_15895);
or U16055 (N_16055,N_15831,N_15830);
nand U16056 (N_16056,N_15959,N_15804);
or U16057 (N_16057,N_15919,N_15848);
xor U16058 (N_16058,N_15918,N_15936);
and U16059 (N_16059,N_15970,N_15813);
nor U16060 (N_16060,N_15954,N_15909);
or U16061 (N_16061,N_15811,N_15828);
nor U16062 (N_16062,N_15988,N_15843);
xor U16063 (N_16063,N_15880,N_15817);
nor U16064 (N_16064,N_15900,N_15858);
nor U16065 (N_16065,N_15820,N_15934);
nand U16066 (N_16066,N_15897,N_15827);
nand U16067 (N_16067,N_15883,N_15912);
or U16068 (N_16068,N_15837,N_15978);
nand U16069 (N_16069,N_15997,N_15915);
or U16070 (N_16070,N_15944,N_15985);
nor U16071 (N_16071,N_15961,N_15855);
xor U16072 (N_16072,N_15999,N_15949);
nor U16073 (N_16073,N_15878,N_15964);
nand U16074 (N_16074,N_15888,N_15841);
or U16075 (N_16075,N_15993,N_15874);
xor U16076 (N_16076,N_15908,N_15870);
and U16077 (N_16077,N_15821,N_15832);
xnor U16078 (N_16078,N_15865,N_15958);
and U16079 (N_16079,N_15864,N_15802);
or U16080 (N_16080,N_15931,N_15966);
nor U16081 (N_16081,N_15971,N_15907);
or U16082 (N_16082,N_15884,N_15921);
nand U16083 (N_16083,N_15914,N_15928);
nor U16084 (N_16084,N_15968,N_15838);
xor U16085 (N_16085,N_15905,N_15846);
and U16086 (N_16086,N_15847,N_15982);
xnor U16087 (N_16087,N_15840,N_15815);
or U16088 (N_16088,N_15965,N_15901);
nor U16089 (N_16089,N_15952,N_15984);
and U16090 (N_16090,N_15946,N_15898);
and U16091 (N_16091,N_15823,N_15875);
or U16092 (N_16092,N_15896,N_15992);
and U16093 (N_16093,N_15816,N_15856);
nor U16094 (N_16094,N_15976,N_15953);
xnor U16095 (N_16095,N_15980,N_15947);
and U16096 (N_16096,N_15871,N_15994);
nor U16097 (N_16097,N_15857,N_15845);
and U16098 (N_16098,N_15941,N_15991);
nor U16099 (N_16099,N_15973,N_15922);
nor U16100 (N_16100,N_15883,N_15952);
xnor U16101 (N_16101,N_15854,N_15892);
and U16102 (N_16102,N_15812,N_15941);
nand U16103 (N_16103,N_15918,N_15815);
nand U16104 (N_16104,N_15915,N_15993);
or U16105 (N_16105,N_15870,N_15948);
nand U16106 (N_16106,N_15897,N_15917);
and U16107 (N_16107,N_15896,N_15888);
xnor U16108 (N_16108,N_15884,N_15979);
nand U16109 (N_16109,N_15895,N_15898);
nand U16110 (N_16110,N_15823,N_15807);
nand U16111 (N_16111,N_15980,N_15906);
and U16112 (N_16112,N_15804,N_15948);
and U16113 (N_16113,N_15890,N_15878);
xor U16114 (N_16114,N_15938,N_15998);
nand U16115 (N_16115,N_15815,N_15809);
nand U16116 (N_16116,N_15941,N_15879);
xor U16117 (N_16117,N_15972,N_15879);
xor U16118 (N_16118,N_15877,N_15818);
nor U16119 (N_16119,N_15881,N_15846);
nor U16120 (N_16120,N_15960,N_15852);
nor U16121 (N_16121,N_15937,N_15961);
or U16122 (N_16122,N_15957,N_15916);
xnor U16123 (N_16123,N_15996,N_15924);
nor U16124 (N_16124,N_15969,N_15931);
or U16125 (N_16125,N_15973,N_15832);
nor U16126 (N_16126,N_15870,N_15940);
or U16127 (N_16127,N_15833,N_15853);
nand U16128 (N_16128,N_15810,N_15901);
nor U16129 (N_16129,N_15942,N_15865);
nor U16130 (N_16130,N_15935,N_15801);
nand U16131 (N_16131,N_15989,N_15987);
xor U16132 (N_16132,N_15919,N_15872);
and U16133 (N_16133,N_15898,N_15849);
nor U16134 (N_16134,N_15874,N_15965);
xor U16135 (N_16135,N_15960,N_15991);
or U16136 (N_16136,N_15842,N_15863);
and U16137 (N_16137,N_15963,N_15995);
nor U16138 (N_16138,N_15869,N_15992);
nor U16139 (N_16139,N_15830,N_15842);
nor U16140 (N_16140,N_15905,N_15912);
and U16141 (N_16141,N_15821,N_15940);
and U16142 (N_16142,N_15812,N_15854);
or U16143 (N_16143,N_15802,N_15993);
or U16144 (N_16144,N_15919,N_15839);
nand U16145 (N_16145,N_15837,N_15897);
and U16146 (N_16146,N_15948,N_15899);
nor U16147 (N_16147,N_15902,N_15965);
xor U16148 (N_16148,N_15899,N_15807);
nand U16149 (N_16149,N_15961,N_15847);
nand U16150 (N_16150,N_15843,N_15908);
nor U16151 (N_16151,N_15814,N_15915);
and U16152 (N_16152,N_15981,N_15815);
nand U16153 (N_16153,N_15830,N_15861);
and U16154 (N_16154,N_15877,N_15852);
and U16155 (N_16155,N_15854,N_15802);
xor U16156 (N_16156,N_15963,N_15916);
and U16157 (N_16157,N_15835,N_15927);
nor U16158 (N_16158,N_15993,N_15883);
and U16159 (N_16159,N_15957,N_15993);
xor U16160 (N_16160,N_15816,N_15951);
nor U16161 (N_16161,N_15950,N_15863);
nand U16162 (N_16162,N_15964,N_15988);
nand U16163 (N_16163,N_15853,N_15807);
and U16164 (N_16164,N_15899,N_15868);
or U16165 (N_16165,N_15882,N_15915);
and U16166 (N_16166,N_15959,N_15967);
nand U16167 (N_16167,N_15957,N_15912);
nand U16168 (N_16168,N_15944,N_15824);
and U16169 (N_16169,N_15949,N_15821);
or U16170 (N_16170,N_15911,N_15887);
or U16171 (N_16171,N_15985,N_15915);
nand U16172 (N_16172,N_15944,N_15827);
or U16173 (N_16173,N_15984,N_15801);
and U16174 (N_16174,N_15833,N_15953);
nand U16175 (N_16175,N_15973,N_15944);
and U16176 (N_16176,N_15968,N_15880);
xnor U16177 (N_16177,N_15825,N_15951);
and U16178 (N_16178,N_15921,N_15960);
or U16179 (N_16179,N_15882,N_15942);
or U16180 (N_16180,N_15883,N_15860);
nor U16181 (N_16181,N_15891,N_15969);
xnor U16182 (N_16182,N_15940,N_15915);
and U16183 (N_16183,N_15978,N_15928);
or U16184 (N_16184,N_15838,N_15923);
nor U16185 (N_16185,N_15884,N_15853);
xnor U16186 (N_16186,N_15941,N_15922);
or U16187 (N_16187,N_15809,N_15876);
nor U16188 (N_16188,N_15831,N_15992);
nand U16189 (N_16189,N_15913,N_15954);
or U16190 (N_16190,N_15945,N_15889);
xor U16191 (N_16191,N_15948,N_15940);
nand U16192 (N_16192,N_15937,N_15905);
or U16193 (N_16193,N_15810,N_15923);
nor U16194 (N_16194,N_15992,N_15939);
and U16195 (N_16195,N_15946,N_15976);
nand U16196 (N_16196,N_15933,N_15912);
xnor U16197 (N_16197,N_15879,N_15839);
nor U16198 (N_16198,N_15815,N_15850);
or U16199 (N_16199,N_15939,N_15824);
or U16200 (N_16200,N_16181,N_16158);
nor U16201 (N_16201,N_16094,N_16063);
nand U16202 (N_16202,N_16044,N_16168);
xor U16203 (N_16203,N_16129,N_16190);
or U16204 (N_16204,N_16024,N_16100);
nand U16205 (N_16205,N_16057,N_16138);
xnor U16206 (N_16206,N_16139,N_16104);
and U16207 (N_16207,N_16083,N_16193);
nor U16208 (N_16208,N_16022,N_16092);
nand U16209 (N_16209,N_16072,N_16074);
nor U16210 (N_16210,N_16126,N_16175);
and U16211 (N_16211,N_16146,N_16141);
and U16212 (N_16212,N_16053,N_16187);
nor U16213 (N_16213,N_16021,N_16095);
or U16214 (N_16214,N_16000,N_16043);
xnor U16215 (N_16215,N_16183,N_16151);
and U16216 (N_16216,N_16125,N_16089);
nand U16217 (N_16217,N_16199,N_16006);
nand U16218 (N_16218,N_16096,N_16157);
nor U16219 (N_16219,N_16069,N_16163);
nor U16220 (N_16220,N_16037,N_16013);
or U16221 (N_16221,N_16029,N_16123);
xor U16222 (N_16222,N_16048,N_16162);
nor U16223 (N_16223,N_16042,N_16115);
nand U16224 (N_16224,N_16004,N_16142);
and U16225 (N_16225,N_16191,N_16064);
and U16226 (N_16226,N_16012,N_16188);
nand U16227 (N_16227,N_16078,N_16179);
nor U16228 (N_16228,N_16153,N_16035);
xnor U16229 (N_16229,N_16150,N_16001);
and U16230 (N_16230,N_16110,N_16061);
nand U16231 (N_16231,N_16046,N_16066);
or U16232 (N_16232,N_16040,N_16113);
nor U16233 (N_16233,N_16030,N_16065);
xor U16234 (N_16234,N_16137,N_16019);
nor U16235 (N_16235,N_16025,N_16082);
or U16236 (N_16236,N_16184,N_16015);
nor U16237 (N_16237,N_16198,N_16173);
nor U16238 (N_16238,N_16014,N_16131);
nor U16239 (N_16239,N_16020,N_16080);
xnor U16240 (N_16240,N_16180,N_16026);
nand U16241 (N_16241,N_16055,N_16165);
and U16242 (N_16242,N_16195,N_16118);
nand U16243 (N_16243,N_16120,N_16116);
and U16244 (N_16244,N_16102,N_16119);
or U16245 (N_16245,N_16156,N_16008);
or U16246 (N_16246,N_16140,N_16122);
xnor U16247 (N_16247,N_16005,N_16192);
or U16248 (N_16248,N_16134,N_16045);
nor U16249 (N_16249,N_16109,N_16166);
nor U16250 (N_16250,N_16068,N_16145);
xor U16251 (N_16251,N_16169,N_16081);
nor U16252 (N_16252,N_16031,N_16133);
and U16253 (N_16253,N_16027,N_16016);
and U16254 (N_16254,N_16196,N_16091);
and U16255 (N_16255,N_16052,N_16185);
nor U16256 (N_16256,N_16105,N_16086);
nor U16257 (N_16257,N_16160,N_16007);
xnor U16258 (N_16258,N_16017,N_16033);
xor U16259 (N_16259,N_16171,N_16148);
xor U16260 (N_16260,N_16107,N_16018);
nor U16261 (N_16261,N_16039,N_16009);
xnor U16262 (N_16262,N_16127,N_16041);
nand U16263 (N_16263,N_16117,N_16088);
nor U16264 (N_16264,N_16167,N_16121);
or U16265 (N_16265,N_16149,N_16111);
xor U16266 (N_16266,N_16085,N_16093);
nor U16267 (N_16267,N_16036,N_16067);
nand U16268 (N_16268,N_16144,N_16186);
xor U16269 (N_16269,N_16050,N_16103);
nand U16270 (N_16270,N_16058,N_16177);
xor U16271 (N_16271,N_16071,N_16054);
nor U16272 (N_16272,N_16147,N_16084);
xnor U16273 (N_16273,N_16114,N_16038);
xor U16274 (N_16274,N_16194,N_16176);
or U16275 (N_16275,N_16056,N_16003);
or U16276 (N_16276,N_16161,N_16130);
xnor U16277 (N_16277,N_16077,N_16049);
xnor U16278 (N_16278,N_16170,N_16002);
nand U16279 (N_16279,N_16070,N_16023);
and U16280 (N_16280,N_16051,N_16136);
and U16281 (N_16281,N_16098,N_16028);
nor U16282 (N_16282,N_16062,N_16075);
xor U16283 (N_16283,N_16132,N_16087);
nor U16284 (N_16284,N_16101,N_16097);
and U16285 (N_16285,N_16032,N_16159);
nor U16286 (N_16286,N_16073,N_16164);
or U16287 (N_16287,N_16172,N_16197);
or U16288 (N_16288,N_16090,N_16112);
or U16289 (N_16289,N_16010,N_16152);
or U16290 (N_16290,N_16182,N_16011);
nor U16291 (N_16291,N_16178,N_16124);
nand U16292 (N_16292,N_16059,N_16034);
nor U16293 (N_16293,N_16106,N_16189);
and U16294 (N_16294,N_16143,N_16060);
nand U16295 (N_16295,N_16076,N_16128);
xnor U16296 (N_16296,N_16099,N_16154);
xnor U16297 (N_16297,N_16047,N_16174);
nor U16298 (N_16298,N_16155,N_16079);
nand U16299 (N_16299,N_16108,N_16135);
or U16300 (N_16300,N_16194,N_16124);
nand U16301 (N_16301,N_16147,N_16163);
nor U16302 (N_16302,N_16180,N_16008);
and U16303 (N_16303,N_16064,N_16168);
or U16304 (N_16304,N_16003,N_16041);
and U16305 (N_16305,N_16053,N_16170);
nand U16306 (N_16306,N_16058,N_16049);
nor U16307 (N_16307,N_16073,N_16060);
or U16308 (N_16308,N_16186,N_16037);
nor U16309 (N_16309,N_16181,N_16015);
or U16310 (N_16310,N_16118,N_16093);
nor U16311 (N_16311,N_16002,N_16143);
nand U16312 (N_16312,N_16085,N_16110);
nand U16313 (N_16313,N_16030,N_16028);
xor U16314 (N_16314,N_16077,N_16062);
xnor U16315 (N_16315,N_16192,N_16057);
nor U16316 (N_16316,N_16145,N_16118);
xnor U16317 (N_16317,N_16069,N_16148);
nor U16318 (N_16318,N_16028,N_16087);
xor U16319 (N_16319,N_16082,N_16101);
and U16320 (N_16320,N_16175,N_16112);
nand U16321 (N_16321,N_16070,N_16030);
or U16322 (N_16322,N_16034,N_16080);
or U16323 (N_16323,N_16129,N_16187);
nand U16324 (N_16324,N_16033,N_16127);
nand U16325 (N_16325,N_16009,N_16133);
xnor U16326 (N_16326,N_16186,N_16027);
and U16327 (N_16327,N_16178,N_16087);
nand U16328 (N_16328,N_16033,N_16118);
nand U16329 (N_16329,N_16031,N_16124);
nor U16330 (N_16330,N_16089,N_16058);
nand U16331 (N_16331,N_16002,N_16140);
nand U16332 (N_16332,N_16163,N_16090);
nand U16333 (N_16333,N_16195,N_16187);
nand U16334 (N_16334,N_16184,N_16077);
nor U16335 (N_16335,N_16064,N_16081);
or U16336 (N_16336,N_16087,N_16124);
nor U16337 (N_16337,N_16021,N_16156);
nand U16338 (N_16338,N_16172,N_16185);
nand U16339 (N_16339,N_16084,N_16028);
xnor U16340 (N_16340,N_16167,N_16144);
or U16341 (N_16341,N_16156,N_16155);
nor U16342 (N_16342,N_16144,N_16115);
nor U16343 (N_16343,N_16069,N_16077);
nand U16344 (N_16344,N_16075,N_16145);
nand U16345 (N_16345,N_16062,N_16044);
nand U16346 (N_16346,N_16170,N_16134);
nor U16347 (N_16347,N_16085,N_16032);
xnor U16348 (N_16348,N_16146,N_16086);
and U16349 (N_16349,N_16169,N_16159);
nand U16350 (N_16350,N_16125,N_16060);
nor U16351 (N_16351,N_16199,N_16165);
xor U16352 (N_16352,N_16091,N_16143);
or U16353 (N_16353,N_16051,N_16045);
and U16354 (N_16354,N_16082,N_16068);
or U16355 (N_16355,N_16146,N_16032);
and U16356 (N_16356,N_16118,N_16045);
nand U16357 (N_16357,N_16096,N_16003);
and U16358 (N_16358,N_16014,N_16106);
xor U16359 (N_16359,N_16033,N_16030);
nor U16360 (N_16360,N_16068,N_16092);
nand U16361 (N_16361,N_16152,N_16117);
nor U16362 (N_16362,N_16061,N_16024);
xor U16363 (N_16363,N_16054,N_16178);
and U16364 (N_16364,N_16178,N_16120);
or U16365 (N_16365,N_16030,N_16020);
nand U16366 (N_16366,N_16007,N_16046);
nand U16367 (N_16367,N_16194,N_16067);
nor U16368 (N_16368,N_16180,N_16187);
nor U16369 (N_16369,N_16048,N_16009);
or U16370 (N_16370,N_16084,N_16004);
nor U16371 (N_16371,N_16027,N_16028);
and U16372 (N_16372,N_16032,N_16116);
and U16373 (N_16373,N_16126,N_16017);
nand U16374 (N_16374,N_16079,N_16131);
and U16375 (N_16375,N_16053,N_16169);
nor U16376 (N_16376,N_16002,N_16191);
xnor U16377 (N_16377,N_16156,N_16097);
xor U16378 (N_16378,N_16148,N_16124);
nand U16379 (N_16379,N_16026,N_16150);
nor U16380 (N_16380,N_16015,N_16079);
or U16381 (N_16381,N_16054,N_16168);
xnor U16382 (N_16382,N_16095,N_16006);
xor U16383 (N_16383,N_16005,N_16019);
or U16384 (N_16384,N_16133,N_16019);
nand U16385 (N_16385,N_16196,N_16179);
or U16386 (N_16386,N_16116,N_16131);
or U16387 (N_16387,N_16068,N_16085);
nor U16388 (N_16388,N_16141,N_16082);
nand U16389 (N_16389,N_16160,N_16159);
and U16390 (N_16390,N_16088,N_16062);
nand U16391 (N_16391,N_16112,N_16195);
xor U16392 (N_16392,N_16071,N_16113);
and U16393 (N_16393,N_16112,N_16167);
nor U16394 (N_16394,N_16166,N_16197);
and U16395 (N_16395,N_16106,N_16131);
nor U16396 (N_16396,N_16037,N_16182);
and U16397 (N_16397,N_16070,N_16003);
xnor U16398 (N_16398,N_16124,N_16110);
and U16399 (N_16399,N_16003,N_16066);
or U16400 (N_16400,N_16229,N_16373);
xnor U16401 (N_16401,N_16224,N_16288);
xor U16402 (N_16402,N_16234,N_16202);
nand U16403 (N_16403,N_16336,N_16231);
xor U16404 (N_16404,N_16335,N_16332);
xnor U16405 (N_16405,N_16361,N_16278);
xor U16406 (N_16406,N_16296,N_16338);
xor U16407 (N_16407,N_16393,N_16362);
and U16408 (N_16408,N_16232,N_16254);
and U16409 (N_16409,N_16344,N_16307);
xor U16410 (N_16410,N_16273,N_16321);
xnor U16411 (N_16411,N_16241,N_16306);
xor U16412 (N_16412,N_16331,N_16384);
nor U16413 (N_16413,N_16374,N_16385);
or U16414 (N_16414,N_16279,N_16289);
and U16415 (N_16415,N_16255,N_16236);
or U16416 (N_16416,N_16295,N_16359);
nand U16417 (N_16417,N_16282,N_16365);
nor U16418 (N_16418,N_16214,N_16286);
xnor U16419 (N_16419,N_16284,N_16397);
and U16420 (N_16420,N_16376,N_16257);
and U16421 (N_16421,N_16323,N_16248);
or U16422 (N_16422,N_16363,N_16237);
nand U16423 (N_16423,N_16339,N_16266);
or U16424 (N_16424,N_16262,N_16390);
or U16425 (N_16425,N_16326,N_16228);
xor U16426 (N_16426,N_16258,N_16270);
or U16427 (N_16427,N_16205,N_16380);
xnor U16428 (N_16428,N_16219,N_16353);
nand U16429 (N_16429,N_16259,N_16378);
nand U16430 (N_16430,N_16216,N_16244);
nand U16431 (N_16431,N_16293,N_16342);
xor U16432 (N_16432,N_16204,N_16301);
nor U16433 (N_16433,N_16240,N_16225);
nor U16434 (N_16434,N_16267,N_16294);
and U16435 (N_16435,N_16337,N_16386);
xor U16436 (N_16436,N_16250,N_16325);
or U16437 (N_16437,N_16371,N_16360);
and U16438 (N_16438,N_16265,N_16238);
nand U16439 (N_16439,N_16227,N_16366);
nand U16440 (N_16440,N_16372,N_16334);
and U16441 (N_16441,N_16312,N_16313);
nand U16442 (N_16442,N_16395,N_16211);
and U16443 (N_16443,N_16311,N_16281);
and U16444 (N_16444,N_16318,N_16212);
nor U16445 (N_16445,N_16230,N_16268);
xnor U16446 (N_16446,N_16308,N_16328);
nor U16447 (N_16447,N_16347,N_16377);
and U16448 (N_16448,N_16220,N_16388);
or U16449 (N_16449,N_16356,N_16271);
nand U16450 (N_16450,N_16309,N_16261);
nand U16451 (N_16451,N_16382,N_16222);
xnor U16452 (N_16452,N_16310,N_16317);
or U16453 (N_16453,N_16218,N_16389);
nand U16454 (N_16454,N_16235,N_16249);
and U16455 (N_16455,N_16333,N_16351);
xor U16456 (N_16456,N_16276,N_16233);
or U16457 (N_16457,N_16203,N_16246);
nand U16458 (N_16458,N_16221,N_16349);
nand U16459 (N_16459,N_16343,N_16302);
and U16460 (N_16460,N_16275,N_16398);
xor U16461 (N_16461,N_16345,N_16243);
nand U16462 (N_16462,N_16263,N_16217);
or U16463 (N_16463,N_16350,N_16277);
and U16464 (N_16464,N_16322,N_16264);
nor U16465 (N_16465,N_16251,N_16314);
and U16466 (N_16466,N_16392,N_16330);
xor U16467 (N_16467,N_16346,N_16290);
xnor U16468 (N_16468,N_16316,N_16292);
or U16469 (N_16469,N_16200,N_16387);
and U16470 (N_16470,N_16291,N_16226);
nor U16471 (N_16471,N_16209,N_16391);
or U16472 (N_16472,N_16299,N_16367);
and U16473 (N_16473,N_16355,N_16358);
or U16474 (N_16474,N_16260,N_16215);
nor U16475 (N_16475,N_16320,N_16285);
nor U16476 (N_16476,N_16201,N_16207);
and U16477 (N_16477,N_16223,N_16357);
nand U16478 (N_16478,N_16381,N_16369);
nor U16479 (N_16479,N_16383,N_16297);
nand U16480 (N_16480,N_16269,N_16304);
nor U16481 (N_16481,N_16256,N_16364);
and U16482 (N_16482,N_16375,N_16368);
nand U16483 (N_16483,N_16239,N_16245);
xor U16484 (N_16484,N_16210,N_16280);
and U16485 (N_16485,N_16247,N_16315);
or U16486 (N_16486,N_16370,N_16341);
nor U16487 (N_16487,N_16399,N_16305);
nor U16488 (N_16488,N_16329,N_16242);
nor U16489 (N_16489,N_16206,N_16274);
nor U16490 (N_16490,N_16319,N_16340);
xnor U16491 (N_16491,N_16272,N_16396);
xor U16492 (N_16492,N_16379,N_16253);
or U16493 (N_16493,N_16348,N_16287);
nand U16494 (N_16494,N_16394,N_16283);
xnor U16495 (N_16495,N_16354,N_16327);
or U16496 (N_16496,N_16300,N_16298);
or U16497 (N_16497,N_16213,N_16324);
or U16498 (N_16498,N_16208,N_16352);
nand U16499 (N_16499,N_16303,N_16252);
or U16500 (N_16500,N_16311,N_16339);
and U16501 (N_16501,N_16275,N_16379);
nand U16502 (N_16502,N_16236,N_16355);
or U16503 (N_16503,N_16316,N_16363);
and U16504 (N_16504,N_16368,N_16352);
nand U16505 (N_16505,N_16263,N_16282);
and U16506 (N_16506,N_16367,N_16329);
nor U16507 (N_16507,N_16214,N_16320);
xnor U16508 (N_16508,N_16203,N_16345);
and U16509 (N_16509,N_16249,N_16222);
and U16510 (N_16510,N_16358,N_16396);
xor U16511 (N_16511,N_16330,N_16218);
nor U16512 (N_16512,N_16372,N_16273);
nand U16513 (N_16513,N_16276,N_16398);
or U16514 (N_16514,N_16392,N_16212);
nand U16515 (N_16515,N_16307,N_16288);
nand U16516 (N_16516,N_16367,N_16371);
and U16517 (N_16517,N_16337,N_16322);
nor U16518 (N_16518,N_16362,N_16274);
nand U16519 (N_16519,N_16253,N_16385);
nand U16520 (N_16520,N_16312,N_16334);
and U16521 (N_16521,N_16244,N_16220);
or U16522 (N_16522,N_16397,N_16379);
nand U16523 (N_16523,N_16302,N_16363);
and U16524 (N_16524,N_16357,N_16251);
and U16525 (N_16525,N_16240,N_16373);
and U16526 (N_16526,N_16346,N_16331);
xnor U16527 (N_16527,N_16232,N_16236);
xnor U16528 (N_16528,N_16369,N_16244);
nand U16529 (N_16529,N_16312,N_16241);
xor U16530 (N_16530,N_16348,N_16275);
or U16531 (N_16531,N_16342,N_16230);
nand U16532 (N_16532,N_16248,N_16392);
xnor U16533 (N_16533,N_16277,N_16369);
nor U16534 (N_16534,N_16289,N_16316);
nor U16535 (N_16535,N_16387,N_16270);
or U16536 (N_16536,N_16255,N_16285);
and U16537 (N_16537,N_16261,N_16232);
or U16538 (N_16538,N_16236,N_16361);
or U16539 (N_16539,N_16245,N_16278);
or U16540 (N_16540,N_16325,N_16291);
or U16541 (N_16541,N_16379,N_16204);
nor U16542 (N_16542,N_16280,N_16237);
xnor U16543 (N_16543,N_16264,N_16390);
xor U16544 (N_16544,N_16307,N_16341);
nor U16545 (N_16545,N_16319,N_16209);
and U16546 (N_16546,N_16309,N_16272);
xnor U16547 (N_16547,N_16265,N_16219);
nor U16548 (N_16548,N_16242,N_16354);
or U16549 (N_16549,N_16347,N_16307);
and U16550 (N_16550,N_16202,N_16359);
and U16551 (N_16551,N_16297,N_16357);
nor U16552 (N_16552,N_16237,N_16283);
xor U16553 (N_16553,N_16314,N_16298);
nand U16554 (N_16554,N_16294,N_16354);
nand U16555 (N_16555,N_16382,N_16366);
and U16556 (N_16556,N_16269,N_16275);
and U16557 (N_16557,N_16259,N_16351);
nand U16558 (N_16558,N_16355,N_16221);
and U16559 (N_16559,N_16330,N_16219);
nand U16560 (N_16560,N_16351,N_16227);
nand U16561 (N_16561,N_16330,N_16265);
or U16562 (N_16562,N_16279,N_16329);
or U16563 (N_16563,N_16346,N_16358);
and U16564 (N_16564,N_16256,N_16399);
or U16565 (N_16565,N_16262,N_16278);
and U16566 (N_16566,N_16211,N_16296);
or U16567 (N_16567,N_16280,N_16294);
nor U16568 (N_16568,N_16373,N_16371);
and U16569 (N_16569,N_16380,N_16223);
nand U16570 (N_16570,N_16286,N_16338);
xnor U16571 (N_16571,N_16237,N_16276);
nor U16572 (N_16572,N_16208,N_16222);
nor U16573 (N_16573,N_16233,N_16249);
or U16574 (N_16574,N_16216,N_16211);
nor U16575 (N_16575,N_16292,N_16240);
and U16576 (N_16576,N_16286,N_16273);
and U16577 (N_16577,N_16256,N_16392);
nand U16578 (N_16578,N_16305,N_16352);
xnor U16579 (N_16579,N_16303,N_16294);
nand U16580 (N_16580,N_16239,N_16252);
nor U16581 (N_16581,N_16338,N_16280);
nor U16582 (N_16582,N_16343,N_16293);
xor U16583 (N_16583,N_16338,N_16202);
xnor U16584 (N_16584,N_16226,N_16325);
xnor U16585 (N_16585,N_16270,N_16255);
nand U16586 (N_16586,N_16243,N_16355);
nand U16587 (N_16587,N_16299,N_16322);
or U16588 (N_16588,N_16236,N_16371);
or U16589 (N_16589,N_16271,N_16349);
nand U16590 (N_16590,N_16396,N_16376);
nor U16591 (N_16591,N_16262,N_16349);
or U16592 (N_16592,N_16359,N_16266);
and U16593 (N_16593,N_16305,N_16244);
and U16594 (N_16594,N_16367,N_16259);
nor U16595 (N_16595,N_16221,N_16242);
xnor U16596 (N_16596,N_16348,N_16298);
and U16597 (N_16597,N_16354,N_16366);
nor U16598 (N_16598,N_16200,N_16283);
xnor U16599 (N_16599,N_16243,N_16315);
nand U16600 (N_16600,N_16579,N_16485);
or U16601 (N_16601,N_16537,N_16512);
xor U16602 (N_16602,N_16549,N_16594);
nor U16603 (N_16603,N_16598,N_16546);
or U16604 (N_16604,N_16582,N_16500);
and U16605 (N_16605,N_16442,N_16520);
xnor U16606 (N_16606,N_16517,N_16591);
nand U16607 (N_16607,N_16443,N_16490);
or U16608 (N_16608,N_16424,N_16590);
or U16609 (N_16609,N_16489,N_16541);
nor U16610 (N_16610,N_16463,N_16554);
and U16611 (N_16611,N_16418,N_16432);
or U16612 (N_16612,N_16521,N_16505);
nand U16613 (N_16613,N_16561,N_16440);
and U16614 (N_16614,N_16564,N_16559);
nand U16615 (N_16615,N_16461,N_16514);
xnor U16616 (N_16616,N_16419,N_16548);
nor U16617 (N_16617,N_16568,N_16577);
xnor U16618 (N_16618,N_16479,N_16545);
xnor U16619 (N_16619,N_16415,N_16474);
or U16620 (N_16620,N_16563,N_16501);
and U16621 (N_16621,N_16544,N_16431);
or U16622 (N_16622,N_16447,N_16406);
and U16623 (N_16623,N_16426,N_16555);
xnor U16624 (N_16624,N_16475,N_16552);
nor U16625 (N_16625,N_16569,N_16483);
nor U16626 (N_16626,N_16515,N_16436);
and U16627 (N_16627,N_16450,N_16471);
nand U16628 (N_16628,N_16428,N_16538);
nand U16629 (N_16629,N_16456,N_16524);
or U16630 (N_16630,N_16468,N_16416);
xor U16631 (N_16631,N_16444,N_16486);
or U16632 (N_16632,N_16478,N_16513);
xor U16633 (N_16633,N_16566,N_16494);
or U16634 (N_16634,N_16454,N_16526);
nand U16635 (N_16635,N_16581,N_16470);
nand U16636 (N_16636,N_16529,N_16482);
nand U16637 (N_16637,N_16575,N_16451);
nor U16638 (N_16638,N_16534,N_16437);
or U16639 (N_16639,N_16528,N_16457);
nor U16640 (N_16640,N_16495,N_16472);
xor U16641 (N_16641,N_16413,N_16452);
or U16642 (N_16642,N_16469,N_16464);
nand U16643 (N_16643,N_16502,N_16589);
nand U16644 (N_16644,N_16498,N_16459);
xnor U16645 (N_16645,N_16571,N_16466);
and U16646 (N_16646,N_16523,N_16562);
or U16647 (N_16647,N_16412,N_16504);
nand U16648 (N_16648,N_16595,N_16565);
nand U16649 (N_16649,N_16570,N_16580);
or U16650 (N_16650,N_16587,N_16527);
nor U16651 (N_16651,N_16441,N_16496);
xnor U16652 (N_16652,N_16400,N_16558);
xor U16653 (N_16653,N_16531,N_16508);
or U16654 (N_16654,N_16560,N_16574);
xnor U16655 (N_16655,N_16407,N_16530);
nand U16656 (N_16656,N_16522,N_16542);
and U16657 (N_16657,N_16585,N_16578);
nand U16658 (N_16658,N_16532,N_16476);
or U16659 (N_16659,N_16435,N_16410);
and U16660 (N_16660,N_16429,N_16543);
nor U16661 (N_16661,N_16525,N_16448);
nor U16662 (N_16662,N_16593,N_16421);
nor U16663 (N_16663,N_16411,N_16427);
nand U16664 (N_16664,N_16516,N_16491);
xnor U16665 (N_16665,N_16572,N_16481);
or U16666 (N_16666,N_16588,N_16402);
and U16667 (N_16667,N_16473,N_16539);
nor U16668 (N_16668,N_16492,N_16550);
xnor U16669 (N_16669,N_16536,N_16477);
nor U16670 (N_16670,N_16507,N_16405);
or U16671 (N_16671,N_16540,N_16453);
nand U16672 (N_16672,N_16488,N_16433);
nand U16673 (N_16673,N_16556,N_16449);
and U16674 (N_16674,N_16467,N_16434);
nor U16675 (N_16675,N_16576,N_16506);
and U16676 (N_16676,N_16592,N_16518);
nand U16677 (N_16677,N_16445,N_16438);
nor U16678 (N_16678,N_16484,N_16509);
nand U16679 (N_16679,N_16551,N_16493);
and U16680 (N_16680,N_16423,N_16409);
or U16681 (N_16681,N_16573,N_16465);
and U16682 (N_16682,N_16557,N_16586);
nor U16683 (N_16683,N_16547,N_16583);
nor U16684 (N_16684,N_16510,N_16439);
nand U16685 (N_16685,N_16401,N_16480);
xnor U16686 (N_16686,N_16422,N_16460);
or U16687 (N_16687,N_16420,N_16596);
and U16688 (N_16688,N_16584,N_16403);
or U16689 (N_16689,N_16519,N_16417);
nor U16690 (N_16690,N_16535,N_16511);
and U16691 (N_16691,N_16487,N_16458);
xor U16692 (N_16692,N_16567,N_16446);
nor U16693 (N_16693,N_16599,N_16503);
and U16694 (N_16694,N_16553,N_16414);
nand U16695 (N_16695,N_16404,N_16497);
and U16696 (N_16696,N_16425,N_16455);
nand U16697 (N_16697,N_16533,N_16597);
or U16698 (N_16698,N_16499,N_16430);
and U16699 (N_16699,N_16462,N_16408);
xor U16700 (N_16700,N_16427,N_16507);
nor U16701 (N_16701,N_16506,N_16493);
or U16702 (N_16702,N_16591,N_16450);
xnor U16703 (N_16703,N_16535,N_16562);
nand U16704 (N_16704,N_16506,N_16598);
and U16705 (N_16705,N_16558,N_16505);
nand U16706 (N_16706,N_16453,N_16522);
xnor U16707 (N_16707,N_16466,N_16473);
and U16708 (N_16708,N_16513,N_16535);
nand U16709 (N_16709,N_16435,N_16553);
and U16710 (N_16710,N_16479,N_16563);
nor U16711 (N_16711,N_16460,N_16579);
nand U16712 (N_16712,N_16497,N_16488);
nor U16713 (N_16713,N_16445,N_16464);
nor U16714 (N_16714,N_16581,N_16456);
nor U16715 (N_16715,N_16516,N_16414);
or U16716 (N_16716,N_16559,N_16429);
nor U16717 (N_16717,N_16530,N_16430);
or U16718 (N_16718,N_16541,N_16407);
and U16719 (N_16719,N_16581,N_16519);
nand U16720 (N_16720,N_16468,N_16573);
or U16721 (N_16721,N_16514,N_16409);
nand U16722 (N_16722,N_16504,N_16400);
or U16723 (N_16723,N_16528,N_16548);
and U16724 (N_16724,N_16539,N_16544);
nor U16725 (N_16725,N_16428,N_16425);
and U16726 (N_16726,N_16460,N_16488);
or U16727 (N_16727,N_16571,N_16583);
xnor U16728 (N_16728,N_16412,N_16539);
xor U16729 (N_16729,N_16448,N_16406);
and U16730 (N_16730,N_16513,N_16465);
xor U16731 (N_16731,N_16581,N_16550);
and U16732 (N_16732,N_16462,N_16558);
and U16733 (N_16733,N_16415,N_16485);
and U16734 (N_16734,N_16500,N_16498);
nand U16735 (N_16735,N_16435,N_16404);
nand U16736 (N_16736,N_16545,N_16562);
and U16737 (N_16737,N_16538,N_16576);
and U16738 (N_16738,N_16532,N_16530);
or U16739 (N_16739,N_16404,N_16549);
and U16740 (N_16740,N_16542,N_16569);
nand U16741 (N_16741,N_16459,N_16545);
nor U16742 (N_16742,N_16574,N_16405);
nor U16743 (N_16743,N_16425,N_16450);
and U16744 (N_16744,N_16485,N_16585);
nand U16745 (N_16745,N_16447,N_16563);
or U16746 (N_16746,N_16411,N_16559);
or U16747 (N_16747,N_16597,N_16549);
nor U16748 (N_16748,N_16450,N_16510);
nor U16749 (N_16749,N_16440,N_16503);
or U16750 (N_16750,N_16400,N_16511);
and U16751 (N_16751,N_16533,N_16578);
xor U16752 (N_16752,N_16593,N_16507);
or U16753 (N_16753,N_16500,N_16559);
nor U16754 (N_16754,N_16534,N_16495);
nand U16755 (N_16755,N_16497,N_16423);
xor U16756 (N_16756,N_16554,N_16410);
or U16757 (N_16757,N_16523,N_16530);
or U16758 (N_16758,N_16579,N_16529);
nor U16759 (N_16759,N_16555,N_16497);
nor U16760 (N_16760,N_16564,N_16454);
and U16761 (N_16761,N_16555,N_16504);
nand U16762 (N_16762,N_16476,N_16465);
xor U16763 (N_16763,N_16447,N_16518);
or U16764 (N_16764,N_16542,N_16461);
or U16765 (N_16765,N_16478,N_16487);
xnor U16766 (N_16766,N_16518,N_16539);
or U16767 (N_16767,N_16493,N_16487);
nand U16768 (N_16768,N_16451,N_16578);
or U16769 (N_16769,N_16532,N_16539);
xor U16770 (N_16770,N_16584,N_16492);
nand U16771 (N_16771,N_16491,N_16470);
nand U16772 (N_16772,N_16447,N_16454);
nand U16773 (N_16773,N_16582,N_16535);
or U16774 (N_16774,N_16575,N_16473);
nor U16775 (N_16775,N_16562,N_16479);
or U16776 (N_16776,N_16597,N_16512);
nand U16777 (N_16777,N_16416,N_16441);
or U16778 (N_16778,N_16504,N_16437);
nor U16779 (N_16779,N_16448,N_16462);
and U16780 (N_16780,N_16490,N_16416);
nor U16781 (N_16781,N_16519,N_16412);
nor U16782 (N_16782,N_16524,N_16446);
and U16783 (N_16783,N_16549,N_16520);
nand U16784 (N_16784,N_16497,N_16462);
xnor U16785 (N_16785,N_16430,N_16482);
xnor U16786 (N_16786,N_16576,N_16404);
xnor U16787 (N_16787,N_16514,N_16501);
nor U16788 (N_16788,N_16548,N_16590);
nor U16789 (N_16789,N_16411,N_16533);
xor U16790 (N_16790,N_16496,N_16538);
nand U16791 (N_16791,N_16435,N_16465);
nor U16792 (N_16792,N_16434,N_16547);
nor U16793 (N_16793,N_16535,N_16578);
nor U16794 (N_16794,N_16448,N_16441);
nand U16795 (N_16795,N_16543,N_16418);
and U16796 (N_16796,N_16550,N_16544);
nand U16797 (N_16797,N_16551,N_16476);
nand U16798 (N_16798,N_16546,N_16490);
nand U16799 (N_16799,N_16511,N_16450);
nor U16800 (N_16800,N_16622,N_16737);
xnor U16801 (N_16801,N_16728,N_16654);
and U16802 (N_16802,N_16681,N_16623);
xor U16803 (N_16803,N_16783,N_16667);
nand U16804 (N_16804,N_16761,N_16793);
or U16805 (N_16805,N_16735,N_16762);
or U16806 (N_16806,N_16790,N_16754);
xor U16807 (N_16807,N_16684,N_16619);
and U16808 (N_16808,N_16701,N_16756);
nor U16809 (N_16809,N_16605,N_16604);
xnor U16810 (N_16810,N_16657,N_16697);
nor U16811 (N_16811,N_16710,N_16789);
and U16812 (N_16812,N_16677,N_16673);
and U16813 (N_16813,N_16750,N_16645);
or U16814 (N_16814,N_16672,N_16624);
and U16815 (N_16815,N_16600,N_16771);
and U16816 (N_16816,N_16692,N_16743);
and U16817 (N_16817,N_16734,N_16788);
nand U16818 (N_16818,N_16755,N_16746);
or U16819 (N_16819,N_16611,N_16659);
xnor U16820 (N_16820,N_16638,N_16658);
and U16821 (N_16821,N_16794,N_16747);
nand U16822 (N_16822,N_16784,N_16769);
and U16823 (N_16823,N_16644,N_16640);
nand U16824 (N_16824,N_16768,N_16760);
or U16825 (N_16825,N_16633,N_16689);
xor U16826 (N_16826,N_16778,N_16765);
nand U16827 (N_16827,N_16617,N_16676);
and U16828 (N_16828,N_16613,N_16661);
nor U16829 (N_16829,N_16655,N_16625);
and U16830 (N_16830,N_16621,N_16695);
nand U16831 (N_16831,N_16719,N_16650);
and U16832 (N_16832,N_16731,N_16705);
xor U16833 (N_16833,N_16685,N_16628);
nand U16834 (N_16834,N_16740,N_16712);
xor U16835 (N_16835,N_16607,N_16739);
nor U16836 (N_16836,N_16724,N_16610);
nand U16837 (N_16837,N_16716,N_16602);
nand U16838 (N_16838,N_16730,N_16608);
and U16839 (N_16839,N_16635,N_16752);
xnor U16840 (N_16840,N_16636,N_16707);
or U16841 (N_16841,N_16631,N_16714);
nand U16842 (N_16842,N_16649,N_16779);
xor U16843 (N_16843,N_16687,N_16698);
and U16844 (N_16844,N_16703,N_16745);
nand U16845 (N_16845,N_16696,N_16767);
and U16846 (N_16846,N_16632,N_16748);
nand U16847 (N_16847,N_16691,N_16799);
and U16848 (N_16848,N_16706,N_16773);
xor U16849 (N_16849,N_16709,N_16715);
or U16850 (N_16850,N_16609,N_16708);
nor U16851 (N_16851,N_16741,N_16776);
xor U16852 (N_16852,N_16642,N_16637);
nor U16853 (N_16853,N_16626,N_16786);
and U16854 (N_16854,N_16757,N_16656);
nor U16855 (N_16855,N_16720,N_16704);
nand U16856 (N_16856,N_16686,N_16666);
or U16857 (N_16857,N_16723,N_16785);
or U16858 (N_16858,N_16782,N_16653);
and U16859 (N_16859,N_16699,N_16780);
or U16860 (N_16860,N_16718,N_16751);
nand U16861 (N_16861,N_16674,N_16787);
nor U16862 (N_16862,N_16744,N_16679);
or U16863 (N_16863,N_16663,N_16618);
or U16864 (N_16864,N_16601,N_16722);
and U16865 (N_16865,N_16764,N_16766);
nand U16866 (N_16866,N_16668,N_16665);
xor U16867 (N_16867,N_16797,N_16648);
or U16868 (N_16868,N_16758,N_16682);
nor U16869 (N_16869,N_16753,N_16634);
nand U16870 (N_16870,N_16693,N_16664);
and U16871 (N_16871,N_16614,N_16725);
and U16872 (N_16872,N_16688,N_16694);
xnor U16873 (N_16873,N_16702,N_16606);
and U16874 (N_16874,N_16732,N_16603);
nand U16875 (N_16875,N_16612,N_16690);
and U16876 (N_16876,N_16770,N_16738);
nand U16877 (N_16877,N_16717,N_16774);
nor U16878 (N_16878,N_16627,N_16711);
or U16879 (N_16879,N_16763,N_16796);
or U16880 (N_16880,N_16678,N_16772);
nand U16881 (N_16881,N_16643,N_16639);
xnor U16882 (N_16882,N_16729,N_16646);
xnor U16883 (N_16883,N_16660,N_16675);
xnor U16884 (N_16884,N_16662,N_16721);
and U16885 (N_16885,N_16700,N_16791);
nor U16886 (N_16886,N_16727,N_16620);
or U16887 (N_16887,N_16795,N_16733);
or U16888 (N_16888,N_16652,N_16629);
and U16889 (N_16889,N_16726,N_16775);
or U16890 (N_16890,N_16669,N_16742);
or U16891 (N_16891,N_16683,N_16736);
nor U16892 (N_16892,N_16641,N_16647);
nor U16893 (N_16893,N_16777,N_16792);
nor U16894 (N_16894,N_16713,N_16680);
nor U16895 (N_16895,N_16616,N_16671);
nand U16896 (N_16896,N_16759,N_16615);
and U16897 (N_16897,N_16781,N_16630);
nor U16898 (N_16898,N_16670,N_16798);
nand U16899 (N_16899,N_16749,N_16651);
and U16900 (N_16900,N_16689,N_16745);
and U16901 (N_16901,N_16794,N_16789);
xor U16902 (N_16902,N_16657,N_16767);
and U16903 (N_16903,N_16733,N_16724);
nor U16904 (N_16904,N_16643,N_16777);
and U16905 (N_16905,N_16683,N_16653);
nand U16906 (N_16906,N_16701,N_16616);
nand U16907 (N_16907,N_16724,N_16765);
nand U16908 (N_16908,N_16719,N_16608);
or U16909 (N_16909,N_16630,N_16684);
nor U16910 (N_16910,N_16763,N_16719);
xnor U16911 (N_16911,N_16687,N_16684);
or U16912 (N_16912,N_16746,N_16668);
and U16913 (N_16913,N_16787,N_16782);
nand U16914 (N_16914,N_16782,N_16750);
and U16915 (N_16915,N_16682,N_16771);
or U16916 (N_16916,N_16613,N_16643);
xor U16917 (N_16917,N_16605,N_16724);
nand U16918 (N_16918,N_16763,N_16720);
and U16919 (N_16919,N_16790,N_16761);
nand U16920 (N_16920,N_16703,N_16600);
nor U16921 (N_16921,N_16628,N_16712);
and U16922 (N_16922,N_16676,N_16791);
xnor U16923 (N_16923,N_16675,N_16614);
nor U16924 (N_16924,N_16772,N_16688);
nand U16925 (N_16925,N_16621,N_16750);
nor U16926 (N_16926,N_16768,N_16691);
xnor U16927 (N_16927,N_16672,N_16615);
or U16928 (N_16928,N_16772,N_16656);
or U16929 (N_16929,N_16742,N_16713);
nand U16930 (N_16930,N_16679,N_16777);
nor U16931 (N_16931,N_16678,N_16664);
nor U16932 (N_16932,N_16634,N_16705);
xor U16933 (N_16933,N_16750,N_16629);
nand U16934 (N_16934,N_16609,N_16725);
nand U16935 (N_16935,N_16688,N_16668);
nor U16936 (N_16936,N_16781,N_16664);
or U16937 (N_16937,N_16766,N_16697);
nand U16938 (N_16938,N_16797,N_16788);
nand U16939 (N_16939,N_16622,N_16631);
xor U16940 (N_16940,N_16721,N_16667);
and U16941 (N_16941,N_16758,N_16685);
and U16942 (N_16942,N_16746,N_16735);
or U16943 (N_16943,N_16777,N_16659);
xor U16944 (N_16944,N_16748,N_16701);
xnor U16945 (N_16945,N_16750,N_16667);
nand U16946 (N_16946,N_16679,N_16785);
nand U16947 (N_16947,N_16746,N_16666);
or U16948 (N_16948,N_16698,N_16684);
or U16949 (N_16949,N_16653,N_16793);
nand U16950 (N_16950,N_16769,N_16714);
nand U16951 (N_16951,N_16679,N_16620);
xnor U16952 (N_16952,N_16667,N_16794);
xnor U16953 (N_16953,N_16670,N_16634);
nand U16954 (N_16954,N_16792,N_16767);
and U16955 (N_16955,N_16666,N_16683);
xor U16956 (N_16956,N_16618,N_16658);
or U16957 (N_16957,N_16601,N_16707);
nand U16958 (N_16958,N_16788,N_16619);
nor U16959 (N_16959,N_16603,N_16608);
and U16960 (N_16960,N_16635,N_16745);
nand U16961 (N_16961,N_16735,N_16642);
nand U16962 (N_16962,N_16614,N_16770);
nand U16963 (N_16963,N_16765,N_16685);
nand U16964 (N_16964,N_16749,N_16638);
xnor U16965 (N_16965,N_16675,N_16715);
and U16966 (N_16966,N_16636,N_16684);
and U16967 (N_16967,N_16739,N_16652);
xnor U16968 (N_16968,N_16665,N_16620);
nand U16969 (N_16969,N_16785,N_16704);
nand U16970 (N_16970,N_16654,N_16634);
nor U16971 (N_16971,N_16690,N_16663);
and U16972 (N_16972,N_16634,N_16647);
xor U16973 (N_16973,N_16709,N_16657);
nand U16974 (N_16974,N_16735,N_16646);
xor U16975 (N_16975,N_16605,N_16688);
and U16976 (N_16976,N_16718,N_16756);
or U16977 (N_16977,N_16789,N_16675);
or U16978 (N_16978,N_16667,N_16649);
nand U16979 (N_16979,N_16707,N_16763);
xor U16980 (N_16980,N_16759,N_16604);
nor U16981 (N_16981,N_16624,N_16678);
and U16982 (N_16982,N_16764,N_16637);
nand U16983 (N_16983,N_16685,N_16704);
and U16984 (N_16984,N_16797,N_16763);
nand U16985 (N_16985,N_16678,N_16642);
xnor U16986 (N_16986,N_16633,N_16762);
or U16987 (N_16987,N_16691,N_16613);
and U16988 (N_16988,N_16785,N_16672);
or U16989 (N_16989,N_16757,N_16790);
xor U16990 (N_16990,N_16799,N_16751);
or U16991 (N_16991,N_16715,N_16652);
or U16992 (N_16992,N_16641,N_16727);
nand U16993 (N_16993,N_16623,N_16771);
nand U16994 (N_16994,N_16778,N_16709);
nor U16995 (N_16995,N_16719,N_16735);
xnor U16996 (N_16996,N_16653,N_16744);
nor U16997 (N_16997,N_16677,N_16765);
xnor U16998 (N_16998,N_16713,N_16761);
xor U16999 (N_16999,N_16650,N_16741);
nand U17000 (N_17000,N_16815,N_16943);
xor U17001 (N_17001,N_16827,N_16866);
or U17002 (N_17002,N_16819,N_16854);
xnor U17003 (N_17003,N_16898,N_16939);
xor U17004 (N_17004,N_16818,N_16864);
nor U17005 (N_17005,N_16812,N_16869);
or U17006 (N_17006,N_16978,N_16965);
xnor U17007 (N_17007,N_16880,N_16909);
and U17008 (N_17008,N_16901,N_16942);
nand U17009 (N_17009,N_16834,N_16910);
or U17010 (N_17010,N_16875,N_16906);
nor U17011 (N_17011,N_16907,N_16929);
xnor U17012 (N_17012,N_16997,N_16878);
or U17013 (N_17013,N_16853,N_16999);
or U17014 (N_17014,N_16979,N_16991);
or U17015 (N_17015,N_16844,N_16894);
nor U17016 (N_17016,N_16821,N_16881);
or U17017 (N_17017,N_16852,N_16889);
xor U17018 (N_17018,N_16908,N_16813);
nand U17019 (N_17019,N_16849,N_16996);
nor U17020 (N_17020,N_16990,N_16920);
and U17021 (N_17021,N_16856,N_16937);
nor U17022 (N_17022,N_16893,N_16971);
and U17023 (N_17023,N_16967,N_16884);
nor U17024 (N_17024,N_16896,N_16876);
xor U17025 (N_17025,N_16953,N_16987);
nor U17026 (N_17026,N_16919,N_16947);
xor U17027 (N_17027,N_16850,N_16961);
nor U17028 (N_17028,N_16989,N_16868);
xor U17029 (N_17029,N_16941,N_16882);
xnor U17030 (N_17030,N_16822,N_16954);
xnor U17031 (N_17031,N_16826,N_16841);
or U17032 (N_17032,N_16981,N_16934);
or U17033 (N_17033,N_16933,N_16940);
xnor U17034 (N_17034,N_16955,N_16900);
or U17035 (N_17035,N_16982,N_16842);
nor U17036 (N_17036,N_16924,N_16848);
nand U17037 (N_17037,N_16950,N_16994);
nor U17038 (N_17038,N_16923,N_16951);
nor U17039 (N_17039,N_16973,N_16915);
and U17040 (N_17040,N_16857,N_16952);
or U17041 (N_17041,N_16830,N_16807);
nand U17042 (N_17042,N_16816,N_16902);
nor U17043 (N_17043,N_16823,N_16840);
and U17044 (N_17044,N_16970,N_16914);
nand U17045 (N_17045,N_16870,N_16992);
and U17046 (N_17046,N_16845,N_16956);
and U17047 (N_17047,N_16886,N_16873);
and U17048 (N_17048,N_16890,N_16862);
xnor U17049 (N_17049,N_16865,N_16832);
nor U17050 (N_17050,N_16828,N_16925);
nand U17051 (N_17051,N_16858,N_16949);
or U17052 (N_17052,N_16957,N_16879);
or U17053 (N_17053,N_16995,N_16824);
nor U17054 (N_17054,N_16851,N_16839);
or U17055 (N_17055,N_16846,N_16921);
nor U17056 (N_17056,N_16905,N_16930);
nand U17057 (N_17057,N_16847,N_16903);
xor U17058 (N_17058,N_16962,N_16988);
nand U17059 (N_17059,N_16912,N_16963);
and U17060 (N_17060,N_16887,N_16980);
and U17061 (N_17061,N_16946,N_16825);
or U17062 (N_17062,N_16810,N_16803);
nor U17063 (N_17063,N_16872,N_16945);
nand U17064 (N_17064,N_16977,N_16806);
nor U17065 (N_17065,N_16927,N_16833);
and U17066 (N_17066,N_16938,N_16968);
xor U17067 (N_17067,N_16993,N_16829);
or U17068 (N_17068,N_16809,N_16804);
nand U17069 (N_17069,N_16891,N_16897);
and U17070 (N_17070,N_16817,N_16985);
and U17071 (N_17071,N_16918,N_16831);
xor U17072 (N_17072,N_16936,N_16838);
nand U17073 (N_17073,N_16917,N_16855);
nor U17074 (N_17074,N_16972,N_16913);
and U17075 (N_17075,N_16966,N_16811);
nand U17076 (N_17076,N_16861,N_16960);
nand U17077 (N_17077,N_16835,N_16935);
xor U17078 (N_17078,N_16911,N_16892);
xor U17079 (N_17079,N_16888,N_16874);
and U17080 (N_17080,N_16975,N_16932);
or U17081 (N_17081,N_16883,N_16836);
xnor U17082 (N_17082,N_16984,N_16800);
and U17083 (N_17083,N_16801,N_16859);
and U17084 (N_17084,N_16928,N_16871);
and U17085 (N_17085,N_16958,N_16922);
xnor U17086 (N_17086,N_16948,N_16899);
nand U17087 (N_17087,N_16814,N_16808);
xnor U17088 (N_17088,N_16837,N_16904);
and U17089 (N_17089,N_16877,N_16944);
and U17090 (N_17090,N_16805,N_16959);
nor U17091 (N_17091,N_16986,N_16895);
nand U17092 (N_17092,N_16916,N_16926);
nand U17093 (N_17093,N_16969,N_16863);
or U17094 (N_17094,N_16802,N_16860);
or U17095 (N_17095,N_16964,N_16931);
or U17096 (N_17096,N_16976,N_16820);
nand U17097 (N_17097,N_16867,N_16885);
or U17098 (N_17098,N_16843,N_16974);
nor U17099 (N_17099,N_16983,N_16998);
nand U17100 (N_17100,N_16812,N_16825);
and U17101 (N_17101,N_16993,N_16824);
nor U17102 (N_17102,N_16807,N_16835);
or U17103 (N_17103,N_16827,N_16969);
and U17104 (N_17104,N_16907,N_16976);
or U17105 (N_17105,N_16822,N_16876);
or U17106 (N_17106,N_16993,N_16850);
nand U17107 (N_17107,N_16870,N_16910);
nand U17108 (N_17108,N_16825,N_16871);
nand U17109 (N_17109,N_16857,N_16930);
and U17110 (N_17110,N_16829,N_16926);
or U17111 (N_17111,N_16863,N_16981);
nor U17112 (N_17112,N_16883,N_16823);
xnor U17113 (N_17113,N_16903,N_16827);
or U17114 (N_17114,N_16970,N_16899);
and U17115 (N_17115,N_16804,N_16827);
or U17116 (N_17116,N_16885,N_16815);
nor U17117 (N_17117,N_16935,N_16808);
xnor U17118 (N_17118,N_16989,N_16919);
and U17119 (N_17119,N_16906,N_16833);
nand U17120 (N_17120,N_16964,N_16981);
and U17121 (N_17121,N_16926,N_16886);
xor U17122 (N_17122,N_16936,N_16844);
nand U17123 (N_17123,N_16829,N_16947);
and U17124 (N_17124,N_16866,N_16833);
nand U17125 (N_17125,N_16818,N_16894);
and U17126 (N_17126,N_16888,N_16941);
xnor U17127 (N_17127,N_16995,N_16860);
nor U17128 (N_17128,N_16869,N_16828);
and U17129 (N_17129,N_16891,N_16996);
xnor U17130 (N_17130,N_16933,N_16917);
or U17131 (N_17131,N_16804,N_16817);
or U17132 (N_17132,N_16810,N_16956);
xor U17133 (N_17133,N_16922,N_16997);
nor U17134 (N_17134,N_16995,N_16875);
nand U17135 (N_17135,N_16958,N_16900);
nor U17136 (N_17136,N_16820,N_16957);
nor U17137 (N_17137,N_16825,N_16971);
and U17138 (N_17138,N_16840,N_16937);
nand U17139 (N_17139,N_16811,N_16956);
xnor U17140 (N_17140,N_16869,N_16856);
or U17141 (N_17141,N_16909,N_16821);
xor U17142 (N_17142,N_16804,N_16842);
and U17143 (N_17143,N_16801,N_16954);
or U17144 (N_17144,N_16839,N_16923);
nor U17145 (N_17145,N_16970,N_16925);
nand U17146 (N_17146,N_16984,N_16835);
xnor U17147 (N_17147,N_16942,N_16943);
or U17148 (N_17148,N_16850,N_16905);
nand U17149 (N_17149,N_16998,N_16882);
and U17150 (N_17150,N_16992,N_16934);
nor U17151 (N_17151,N_16810,N_16836);
nor U17152 (N_17152,N_16885,N_16874);
nor U17153 (N_17153,N_16936,N_16896);
or U17154 (N_17154,N_16806,N_16816);
or U17155 (N_17155,N_16986,N_16802);
and U17156 (N_17156,N_16950,N_16888);
or U17157 (N_17157,N_16932,N_16814);
nor U17158 (N_17158,N_16890,N_16845);
or U17159 (N_17159,N_16958,N_16825);
or U17160 (N_17160,N_16942,N_16980);
xnor U17161 (N_17161,N_16804,N_16806);
nor U17162 (N_17162,N_16821,N_16907);
nor U17163 (N_17163,N_16966,N_16967);
nor U17164 (N_17164,N_16916,N_16872);
nor U17165 (N_17165,N_16845,N_16876);
nor U17166 (N_17166,N_16940,N_16861);
and U17167 (N_17167,N_16905,N_16879);
and U17168 (N_17168,N_16825,N_16814);
xor U17169 (N_17169,N_16944,N_16928);
nor U17170 (N_17170,N_16928,N_16804);
and U17171 (N_17171,N_16997,N_16882);
xor U17172 (N_17172,N_16820,N_16879);
nand U17173 (N_17173,N_16816,N_16829);
nor U17174 (N_17174,N_16922,N_16888);
xor U17175 (N_17175,N_16871,N_16946);
xor U17176 (N_17176,N_16996,N_16839);
nand U17177 (N_17177,N_16982,N_16896);
nor U17178 (N_17178,N_16962,N_16995);
nor U17179 (N_17179,N_16824,N_16928);
or U17180 (N_17180,N_16966,N_16839);
xor U17181 (N_17181,N_16932,N_16850);
xor U17182 (N_17182,N_16803,N_16978);
nand U17183 (N_17183,N_16954,N_16841);
nor U17184 (N_17184,N_16812,N_16892);
nor U17185 (N_17185,N_16815,N_16820);
xor U17186 (N_17186,N_16807,N_16916);
or U17187 (N_17187,N_16983,N_16967);
xnor U17188 (N_17188,N_16902,N_16935);
nor U17189 (N_17189,N_16858,N_16837);
and U17190 (N_17190,N_16928,N_16849);
or U17191 (N_17191,N_16857,N_16951);
or U17192 (N_17192,N_16949,N_16889);
xor U17193 (N_17193,N_16802,N_16946);
nand U17194 (N_17194,N_16865,N_16960);
and U17195 (N_17195,N_16917,N_16972);
xnor U17196 (N_17196,N_16958,N_16963);
or U17197 (N_17197,N_16901,N_16960);
xnor U17198 (N_17198,N_16930,N_16925);
or U17199 (N_17199,N_16901,N_16975);
or U17200 (N_17200,N_17077,N_17139);
nand U17201 (N_17201,N_17113,N_17120);
nor U17202 (N_17202,N_17065,N_17148);
xnor U17203 (N_17203,N_17076,N_17052);
nand U17204 (N_17204,N_17190,N_17124);
nand U17205 (N_17205,N_17147,N_17016);
and U17206 (N_17206,N_17030,N_17183);
nand U17207 (N_17207,N_17091,N_17137);
nor U17208 (N_17208,N_17020,N_17083);
or U17209 (N_17209,N_17090,N_17038);
xor U17210 (N_17210,N_17097,N_17143);
nand U17211 (N_17211,N_17035,N_17100);
nor U17212 (N_17212,N_17004,N_17041);
nor U17213 (N_17213,N_17096,N_17153);
nand U17214 (N_17214,N_17199,N_17003);
xnor U17215 (N_17215,N_17019,N_17192);
nor U17216 (N_17216,N_17060,N_17015);
nor U17217 (N_17217,N_17178,N_17138);
or U17218 (N_17218,N_17180,N_17051);
or U17219 (N_17219,N_17197,N_17108);
nor U17220 (N_17220,N_17106,N_17122);
or U17221 (N_17221,N_17159,N_17163);
nand U17222 (N_17222,N_17102,N_17025);
nor U17223 (N_17223,N_17009,N_17133);
or U17224 (N_17224,N_17032,N_17006);
nand U17225 (N_17225,N_17021,N_17007);
and U17226 (N_17226,N_17196,N_17054);
xor U17227 (N_17227,N_17087,N_17135);
nor U17228 (N_17228,N_17177,N_17141);
and U17229 (N_17229,N_17114,N_17053);
or U17230 (N_17230,N_17095,N_17093);
or U17231 (N_17231,N_17011,N_17088);
and U17232 (N_17232,N_17118,N_17013);
xor U17233 (N_17233,N_17134,N_17129);
xor U17234 (N_17234,N_17189,N_17098);
and U17235 (N_17235,N_17017,N_17145);
or U17236 (N_17236,N_17101,N_17027);
xnor U17237 (N_17237,N_17061,N_17058);
nor U17238 (N_17238,N_17043,N_17162);
xnor U17239 (N_17239,N_17028,N_17081);
and U17240 (N_17240,N_17000,N_17018);
xnor U17241 (N_17241,N_17002,N_17170);
or U17242 (N_17242,N_17146,N_17086);
xnor U17243 (N_17243,N_17127,N_17115);
nor U17244 (N_17244,N_17105,N_17079);
nor U17245 (N_17245,N_17109,N_17187);
and U17246 (N_17246,N_17085,N_17029);
and U17247 (N_17247,N_17089,N_17042);
and U17248 (N_17248,N_17155,N_17033);
and U17249 (N_17249,N_17181,N_17092);
and U17250 (N_17250,N_17067,N_17059);
nand U17251 (N_17251,N_17062,N_17166);
or U17252 (N_17252,N_17056,N_17144);
or U17253 (N_17253,N_17174,N_17055);
and U17254 (N_17254,N_17130,N_17064);
nor U17255 (N_17255,N_17024,N_17188);
nor U17256 (N_17256,N_17111,N_17057);
and U17257 (N_17257,N_17023,N_17164);
or U17258 (N_17258,N_17152,N_17151);
nand U17259 (N_17259,N_17165,N_17050);
nand U17260 (N_17260,N_17022,N_17103);
xor U17261 (N_17261,N_17049,N_17154);
or U17262 (N_17262,N_17012,N_17168);
xnor U17263 (N_17263,N_17126,N_17161);
nor U17264 (N_17264,N_17099,N_17167);
nor U17265 (N_17265,N_17066,N_17047);
nor U17266 (N_17266,N_17014,N_17082);
nand U17267 (N_17267,N_17010,N_17158);
and U17268 (N_17268,N_17037,N_17198);
nand U17269 (N_17269,N_17080,N_17128);
nor U17270 (N_17270,N_17036,N_17107);
and U17271 (N_17271,N_17045,N_17169);
nand U17272 (N_17272,N_17173,N_17123);
or U17273 (N_17273,N_17182,N_17156);
and U17274 (N_17274,N_17104,N_17070);
nand U17275 (N_17275,N_17039,N_17034);
nor U17276 (N_17276,N_17131,N_17026);
xor U17277 (N_17277,N_17195,N_17110);
xnor U17278 (N_17278,N_17048,N_17008);
or U17279 (N_17279,N_17119,N_17112);
xnor U17280 (N_17280,N_17184,N_17094);
or U17281 (N_17281,N_17160,N_17136);
or U17282 (N_17282,N_17071,N_17149);
and U17283 (N_17283,N_17125,N_17175);
nor U17284 (N_17284,N_17140,N_17072);
nor U17285 (N_17285,N_17117,N_17185);
and U17286 (N_17286,N_17179,N_17001);
and U17287 (N_17287,N_17142,N_17171);
nand U17288 (N_17288,N_17069,N_17046);
xnor U17289 (N_17289,N_17068,N_17044);
xnor U17290 (N_17290,N_17191,N_17116);
xnor U17291 (N_17291,N_17078,N_17176);
nor U17292 (N_17292,N_17172,N_17150);
and U17293 (N_17293,N_17157,N_17031);
and U17294 (N_17294,N_17084,N_17040);
nand U17295 (N_17295,N_17121,N_17186);
and U17296 (N_17296,N_17073,N_17193);
or U17297 (N_17297,N_17194,N_17132);
and U17298 (N_17298,N_17075,N_17063);
and U17299 (N_17299,N_17005,N_17074);
and U17300 (N_17300,N_17094,N_17096);
xnor U17301 (N_17301,N_17112,N_17003);
and U17302 (N_17302,N_17007,N_17139);
or U17303 (N_17303,N_17003,N_17143);
nor U17304 (N_17304,N_17079,N_17019);
xor U17305 (N_17305,N_17040,N_17193);
or U17306 (N_17306,N_17179,N_17159);
and U17307 (N_17307,N_17095,N_17081);
xor U17308 (N_17308,N_17138,N_17026);
or U17309 (N_17309,N_17148,N_17110);
and U17310 (N_17310,N_17199,N_17030);
xor U17311 (N_17311,N_17123,N_17124);
xor U17312 (N_17312,N_17151,N_17185);
xor U17313 (N_17313,N_17089,N_17119);
or U17314 (N_17314,N_17022,N_17057);
and U17315 (N_17315,N_17111,N_17171);
and U17316 (N_17316,N_17196,N_17188);
nand U17317 (N_17317,N_17110,N_17061);
and U17318 (N_17318,N_17178,N_17164);
xor U17319 (N_17319,N_17142,N_17045);
and U17320 (N_17320,N_17171,N_17113);
and U17321 (N_17321,N_17141,N_17024);
xor U17322 (N_17322,N_17110,N_17199);
or U17323 (N_17323,N_17114,N_17048);
nand U17324 (N_17324,N_17175,N_17039);
and U17325 (N_17325,N_17174,N_17060);
nor U17326 (N_17326,N_17114,N_17141);
nand U17327 (N_17327,N_17118,N_17014);
xnor U17328 (N_17328,N_17112,N_17047);
nand U17329 (N_17329,N_17168,N_17108);
nand U17330 (N_17330,N_17063,N_17163);
xnor U17331 (N_17331,N_17052,N_17047);
and U17332 (N_17332,N_17185,N_17039);
xor U17333 (N_17333,N_17010,N_17009);
xor U17334 (N_17334,N_17009,N_17031);
or U17335 (N_17335,N_17160,N_17021);
and U17336 (N_17336,N_17080,N_17175);
xnor U17337 (N_17337,N_17101,N_17040);
nor U17338 (N_17338,N_17079,N_17048);
and U17339 (N_17339,N_17131,N_17145);
nand U17340 (N_17340,N_17008,N_17079);
xnor U17341 (N_17341,N_17123,N_17083);
nand U17342 (N_17342,N_17124,N_17078);
xor U17343 (N_17343,N_17065,N_17102);
xnor U17344 (N_17344,N_17091,N_17028);
xnor U17345 (N_17345,N_17112,N_17005);
nor U17346 (N_17346,N_17020,N_17156);
or U17347 (N_17347,N_17021,N_17018);
nor U17348 (N_17348,N_17087,N_17073);
nand U17349 (N_17349,N_17067,N_17164);
xnor U17350 (N_17350,N_17142,N_17094);
xor U17351 (N_17351,N_17163,N_17049);
or U17352 (N_17352,N_17160,N_17156);
nand U17353 (N_17353,N_17112,N_17176);
and U17354 (N_17354,N_17159,N_17165);
xor U17355 (N_17355,N_17000,N_17128);
xor U17356 (N_17356,N_17160,N_17001);
and U17357 (N_17357,N_17172,N_17011);
or U17358 (N_17358,N_17083,N_17131);
or U17359 (N_17359,N_17144,N_17005);
or U17360 (N_17360,N_17050,N_17002);
nand U17361 (N_17361,N_17097,N_17052);
xnor U17362 (N_17362,N_17179,N_17064);
xor U17363 (N_17363,N_17041,N_17123);
or U17364 (N_17364,N_17182,N_17183);
or U17365 (N_17365,N_17157,N_17097);
or U17366 (N_17366,N_17134,N_17154);
or U17367 (N_17367,N_17138,N_17118);
nand U17368 (N_17368,N_17159,N_17000);
and U17369 (N_17369,N_17090,N_17108);
and U17370 (N_17370,N_17142,N_17143);
nand U17371 (N_17371,N_17190,N_17070);
xnor U17372 (N_17372,N_17017,N_17182);
xnor U17373 (N_17373,N_17105,N_17061);
nand U17374 (N_17374,N_17128,N_17013);
and U17375 (N_17375,N_17012,N_17147);
and U17376 (N_17376,N_17040,N_17029);
nor U17377 (N_17377,N_17074,N_17199);
or U17378 (N_17378,N_17024,N_17146);
xor U17379 (N_17379,N_17039,N_17124);
xor U17380 (N_17380,N_17025,N_17184);
or U17381 (N_17381,N_17197,N_17094);
nand U17382 (N_17382,N_17027,N_17179);
and U17383 (N_17383,N_17079,N_17078);
and U17384 (N_17384,N_17088,N_17198);
or U17385 (N_17385,N_17004,N_17035);
xor U17386 (N_17386,N_17003,N_17191);
xor U17387 (N_17387,N_17128,N_17001);
xnor U17388 (N_17388,N_17098,N_17131);
or U17389 (N_17389,N_17151,N_17141);
and U17390 (N_17390,N_17191,N_17125);
nand U17391 (N_17391,N_17172,N_17034);
nor U17392 (N_17392,N_17158,N_17018);
and U17393 (N_17393,N_17112,N_17107);
xor U17394 (N_17394,N_17117,N_17090);
and U17395 (N_17395,N_17154,N_17138);
nor U17396 (N_17396,N_17091,N_17108);
or U17397 (N_17397,N_17179,N_17082);
nand U17398 (N_17398,N_17103,N_17189);
and U17399 (N_17399,N_17181,N_17091);
xnor U17400 (N_17400,N_17245,N_17388);
xnor U17401 (N_17401,N_17383,N_17370);
xor U17402 (N_17402,N_17330,N_17369);
or U17403 (N_17403,N_17317,N_17286);
xnor U17404 (N_17404,N_17293,N_17313);
nor U17405 (N_17405,N_17247,N_17217);
and U17406 (N_17406,N_17209,N_17375);
or U17407 (N_17407,N_17312,N_17229);
and U17408 (N_17408,N_17233,N_17365);
nor U17409 (N_17409,N_17216,N_17322);
or U17410 (N_17410,N_17328,N_17213);
or U17411 (N_17411,N_17324,N_17239);
nor U17412 (N_17412,N_17351,N_17226);
nor U17413 (N_17413,N_17267,N_17254);
xor U17414 (N_17414,N_17251,N_17300);
xor U17415 (N_17415,N_17234,N_17394);
xnor U17416 (N_17416,N_17345,N_17223);
nor U17417 (N_17417,N_17302,N_17220);
or U17418 (N_17418,N_17341,N_17386);
nand U17419 (N_17419,N_17339,N_17290);
xnor U17420 (N_17420,N_17344,N_17360);
and U17421 (N_17421,N_17225,N_17238);
and U17422 (N_17422,N_17391,N_17261);
nor U17423 (N_17423,N_17361,N_17244);
xor U17424 (N_17424,N_17304,N_17219);
nand U17425 (N_17425,N_17236,N_17347);
or U17426 (N_17426,N_17333,N_17235);
and U17427 (N_17427,N_17399,N_17252);
xor U17428 (N_17428,N_17398,N_17311);
nor U17429 (N_17429,N_17340,N_17268);
nor U17430 (N_17430,N_17241,N_17214);
or U17431 (N_17431,N_17308,N_17207);
xnor U17432 (N_17432,N_17358,N_17274);
and U17433 (N_17433,N_17378,N_17348);
nand U17434 (N_17434,N_17326,N_17385);
and U17435 (N_17435,N_17202,N_17390);
or U17436 (N_17436,N_17362,N_17246);
or U17437 (N_17437,N_17323,N_17368);
or U17438 (N_17438,N_17204,N_17357);
nor U17439 (N_17439,N_17210,N_17319);
or U17440 (N_17440,N_17306,N_17352);
and U17441 (N_17441,N_17335,N_17263);
nand U17442 (N_17442,N_17373,N_17309);
nand U17443 (N_17443,N_17305,N_17240);
nor U17444 (N_17444,N_17260,N_17374);
and U17445 (N_17445,N_17270,N_17354);
nand U17446 (N_17446,N_17264,N_17332);
or U17447 (N_17447,N_17283,N_17366);
or U17448 (N_17448,N_17221,N_17337);
and U17449 (N_17449,N_17342,N_17397);
nand U17450 (N_17450,N_17389,N_17280);
or U17451 (N_17451,N_17381,N_17201);
and U17452 (N_17452,N_17355,N_17208);
nor U17453 (N_17453,N_17376,N_17271);
xnor U17454 (N_17454,N_17346,N_17382);
nor U17455 (N_17455,N_17253,N_17279);
or U17456 (N_17456,N_17297,N_17359);
nand U17457 (N_17457,N_17259,N_17248);
or U17458 (N_17458,N_17257,N_17318);
and U17459 (N_17459,N_17228,N_17242);
and U17460 (N_17460,N_17292,N_17282);
nor U17461 (N_17461,N_17262,N_17316);
or U17462 (N_17462,N_17315,N_17379);
nor U17463 (N_17463,N_17266,N_17231);
nor U17464 (N_17464,N_17255,N_17205);
or U17465 (N_17465,N_17285,N_17307);
nand U17466 (N_17466,N_17258,N_17377);
or U17467 (N_17467,N_17350,N_17343);
or U17468 (N_17468,N_17384,N_17288);
nand U17469 (N_17469,N_17275,N_17303);
nand U17470 (N_17470,N_17338,N_17356);
or U17471 (N_17471,N_17314,N_17287);
nand U17472 (N_17472,N_17296,N_17294);
and U17473 (N_17473,N_17349,N_17295);
and U17474 (N_17474,N_17232,N_17371);
and U17475 (N_17475,N_17277,N_17273);
nor U17476 (N_17476,N_17310,N_17380);
nor U17477 (N_17477,N_17230,N_17284);
or U17478 (N_17478,N_17301,N_17325);
or U17479 (N_17479,N_17387,N_17281);
and U17480 (N_17480,N_17227,N_17396);
and U17481 (N_17481,N_17215,N_17372);
and U17482 (N_17482,N_17272,N_17320);
or U17483 (N_17483,N_17212,N_17291);
xnor U17484 (N_17484,N_17276,N_17203);
nand U17485 (N_17485,N_17298,N_17327);
nand U17486 (N_17486,N_17364,N_17218);
and U17487 (N_17487,N_17211,N_17336);
nor U17488 (N_17488,N_17269,N_17329);
and U17489 (N_17489,N_17363,N_17243);
nor U17490 (N_17490,N_17299,N_17289);
xnor U17491 (N_17491,N_17265,N_17206);
nand U17492 (N_17492,N_17278,N_17331);
nand U17493 (N_17493,N_17353,N_17321);
nor U17494 (N_17494,N_17224,N_17249);
nor U17495 (N_17495,N_17367,N_17200);
and U17496 (N_17496,N_17250,N_17334);
nor U17497 (N_17497,N_17393,N_17237);
or U17498 (N_17498,N_17256,N_17392);
nor U17499 (N_17499,N_17222,N_17395);
xnor U17500 (N_17500,N_17316,N_17341);
and U17501 (N_17501,N_17303,N_17374);
xnor U17502 (N_17502,N_17257,N_17352);
and U17503 (N_17503,N_17238,N_17293);
and U17504 (N_17504,N_17306,N_17226);
nand U17505 (N_17505,N_17264,N_17358);
nor U17506 (N_17506,N_17365,N_17257);
xnor U17507 (N_17507,N_17321,N_17210);
or U17508 (N_17508,N_17305,N_17270);
or U17509 (N_17509,N_17254,N_17363);
and U17510 (N_17510,N_17310,N_17362);
nor U17511 (N_17511,N_17294,N_17231);
xnor U17512 (N_17512,N_17345,N_17362);
or U17513 (N_17513,N_17313,N_17219);
xnor U17514 (N_17514,N_17344,N_17227);
or U17515 (N_17515,N_17383,N_17310);
or U17516 (N_17516,N_17358,N_17340);
nand U17517 (N_17517,N_17227,N_17337);
and U17518 (N_17518,N_17203,N_17349);
xor U17519 (N_17519,N_17210,N_17352);
and U17520 (N_17520,N_17366,N_17364);
or U17521 (N_17521,N_17244,N_17292);
or U17522 (N_17522,N_17254,N_17397);
or U17523 (N_17523,N_17388,N_17389);
and U17524 (N_17524,N_17373,N_17297);
nor U17525 (N_17525,N_17371,N_17320);
nand U17526 (N_17526,N_17381,N_17370);
xnor U17527 (N_17527,N_17396,N_17212);
xnor U17528 (N_17528,N_17237,N_17261);
nor U17529 (N_17529,N_17263,N_17356);
nor U17530 (N_17530,N_17340,N_17320);
nor U17531 (N_17531,N_17220,N_17273);
xnor U17532 (N_17532,N_17230,N_17368);
nor U17533 (N_17533,N_17282,N_17251);
nor U17534 (N_17534,N_17208,N_17322);
xor U17535 (N_17535,N_17314,N_17238);
xor U17536 (N_17536,N_17315,N_17294);
nor U17537 (N_17537,N_17389,N_17238);
nand U17538 (N_17538,N_17226,N_17219);
or U17539 (N_17539,N_17324,N_17243);
xor U17540 (N_17540,N_17349,N_17238);
xor U17541 (N_17541,N_17307,N_17263);
xor U17542 (N_17542,N_17347,N_17362);
nor U17543 (N_17543,N_17348,N_17248);
xnor U17544 (N_17544,N_17231,N_17398);
and U17545 (N_17545,N_17379,N_17376);
xnor U17546 (N_17546,N_17356,N_17216);
and U17547 (N_17547,N_17380,N_17268);
and U17548 (N_17548,N_17226,N_17393);
and U17549 (N_17549,N_17312,N_17205);
xor U17550 (N_17550,N_17366,N_17387);
nand U17551 (N_17551,N_17275,N_17366);
xor U17552 (N_17552,N_17308,N_17202);
nand U17553 (N_17553,N_17362,N_17206);
nand U17554 (N_17554,N_17214,N_17261);
and U17555 (N_17555,N_17327,N_17372);
nand U17556 (N_17556,N_17341,N_17304);
nor U17557 (N_17557,N_17219,N_17383);
nand U17558 (N_17558,N_17279,N_17259);
nand U17559 (N_17559,N_17235,N_17373);
nand U17560 (N_17560,N_17330,N_17328);
or U17561 (N_17561,N_17336,N_17224);
nor U17562 (N_17562,N_17213,N_17265);
nor U17563 (N_17563,N_17250,N_17377);
nand U17564 (N_17564,N_17355,N_17201);
xnor U17565 (N_17565,N_17315,N_17287);
or U17566 (N_17566,N_17213,N_17272);
nor U17567 (N_17567,N_17336,N_17389);
nand U17568 (N_17568,N_17346,N_17352);
and U17569 (N_17569,N_17313,N_17247);
and U17570 (N_17570,N_17277,N_17209);
nor U17571 (N_17571,N_17269,N_17322);
nor U17572 (N_17572,N_17321,N_17205);
nor U17573 (N_17573,N_17245,N_17349);
and U17574 (N_17574,N_17252,N_17300);
nand U17575 (N_17575,N_17357,N_17348);
xor U17576 (N_17576,N_17244,N_17386);
and U17577 (N_17577,N_17222,N_17361);
or U17578 (N_17578,N_17270,N_17282);
or U17579 (N_17579,N_17302,N_17344);
xor U17580 (N_17580,N_17321,N_17280);
and U17581 (N_17581,N_17320,N_17215);
or U17582 (N_17582,N_17323,N_17308);
nor U17583 (N_17583,N_17314,N_17246);
nand U17584 (N_17584,N_17364,N_17372);
nand U17585 (N_17585,N_17231,N_17299);
nor U17586 (N_17586,N_17218,N_17372);
or U17587 (N_17587,N_17371,N_17289);
and U17588 (N_17588,N_17399,N_17280);
nor U17589 (N_17589,N_17367,N_17243);
nand U17590 (N_17590,N_17309,N_17353);
nand U17591 (N_17591,N_17312,N_17281);
or U17592 (N_17592,N_17225,N_17300);
nor U17593 (N_17593,N_17339,N_17288);
xnor U17594 (N_17594,N_17229,N_17233);
nand U17595 (N_17595,N_17247,N_17232);
and U17596 (N_17596,N_17292,N_17213);
nor U17597 (N_17597,N_17251,N_17342);
and U17598 (N_17598,N_17319,N_17365);
xor U17599 (N_17599,N_17263,N_17313);
nand U17600 (N_17600,N_17495,N_17465);
and U17601 (N_17601,N_17595,N_17447);
and U17602 (N_17602,N_17590,N_17545);
or U17603 (N_17603,N_17530,N_17539);
nand U17604 (N_17604,N_17586,N_17565);
nand U17605 (N_17605,N_17458,N_17453);
nand U17606 (N_17606,N_17488,N_17515);
nand U17607 (N_17607,N_17434,N_17521);
nand U17608 (N_17608,N_17415,N_17419);
nor U17609 (N_17609,N_17437,N_17416);
xnor U17610 (N_17610,N_17510,N_17485);
nand U17611 (N_17611,N_17534,N_17536);
and U17612 (N_17612,N_17461,N_17591);
xor U17613 (N_17613,N_17540,N_17552);
nor U17614 (N_17614,N_17529,N_17578);
nor U17615 (N_17615,N_17404,N_17581);
xor U17616 (N_17616,N_17579,N_17441);
nor U17617 (N_17617,N_17599,N_17463);
xnor U17618 (N_17618,N_17499,N_17555);
xnor U17619 (N_17619,N_17474,N_17455);
nor U17620 (N_17620,N_17554,N_17561);
nand U17621 (N_17621,N_17500,N_17496);
or U17622 (N_17622,N_17475,N_17572);
nor U17623 (N_17623,N_17596,N_17598);
nand U17624 (N_17624,N_17484,N_17420);
xor U17625 (N_17625,N_17533,N_17594);
and U17626 (N_17626,N_17473,N_17487);
and U17627 (N_17627,N_17535,N_17584);
nand U17628 (N_17628,N_17589,N_17507);
nand U17629 (N_17629,N_17588,N_17449);
xnor U17630 (N_17630,N_17549,N_17582);
or U17631 (N_17631,N_17508,N_17493);
and U17632 (N_17632,N_17580,N_17479);
or U17633 (N_17633,N_17575,N_17513);
nand U17634 (N_17634,N_17450,N_17568);
nand U17635 (N_17635,N_17576,N_17556);
or U17636 (N_17636,N_17526,N_17563);
nand U17637 (N_17637,N_17412,N_17444);
nand U17638 (N_17638,N_17558,N_17490);
or U17639 (N_17639,N_17574,N_17464);
xnor U17640 (N_17640,N_17592,N_17577);
nor U17641 (N_17641,N_17468,N_17446);
nor U17642 (N_17642,N_17462,N_17560);
nor U17643 (N_17643,N_17481,N_17477);
nand U17644 (N_17644,N_17423,N_17425);
nand U17645 (N_17645,N_17432,N_17512);
nor U17646 (N_17646,N_17497,N_17435);
or U17647 (N_17647,N_17506,N_17405);
xor U17648 (N_17648,N_17411,N_17494);
and U17649 (N_17649,N_17439,N_17551);
and U17650 (N_17650,N_17553,N_17478);
or U17651 (N_17651,N_17505,N_17426);
nor U17652 (N_17652,N_17502,N_17541);
nand U17653 (N_17653,N_17452,N_17459);
xnor U17654 (N_17654,N_17550,N_17402);
nand U17655 (N_17655,N_17509,N_17517);
xnor U17656 (N_17656,N_17476,N_17587);
or U17657 (N_17657,N_17492,N_17456);
nor U17658 (N_17658,N_17538,N_17408);
nand U17659 (N_17659,N_17523,N_17454);
nor U17660 (N_17660,N_17466,N_17413);
or U17661 (N_17661,N_17571,N_17451);
or U17662 (N_17662,N_17520,N_17470);
xnor U17663 (N_17663,N_17406,N_17480);
and U17664 (N_17664,N_17491,N_17544);
nand U17665 (N_17665,N_17407,N_17570);
or U17666 (N_17666,N_17471,N_17525);
nand U17667 (N_17667,N_17597,N_17422);
nor U17668 (N_17668,N_17410,N_17547);
xor U17669 (N_17669,N_17522,N_17414);
nor U17670 (N_17670,N_17519,N_17448);
or U17671 (N_17671,N_17442,N_17469);
or U17672 (N_17672,N_17460,N_17524);
nor U17673 (N_17673,N_17593,N_17518);
or U17674 (N_17674,N_17436,N_17567);
nand U17675 (N_17675,N_17400,N_17527);
or U17676 (N_17676,N_17557,N_17430);
xnor U17677 (N_17677,N_17531,N_17503);
xnor U17678 (N_17678,N_17559,N_17542);
nor U17679 (N_17679,N_17421,N_17433);
or U17680 (N_17680,N_17564,N_17548);
nand U17681 (N_17681,N_17511,N_17424);
and U17682 (N_17682,N_17514,N_17467);
nand U17683 (N_17683,N_17428,N_17417);
nand U17684 (N_17684,N_17528,N_17532);
nand U17685 (N_17685,N_17585,N_17504);
or U17686 (N_17686,N_17501,N_17401);
nand U17687 (N_17687,N_17409,N_17445);
and U17688 (N_17688,N_17427,N_17431);
nand U17689 (N_17689,N_17573,N_17429);
and U17690 (N_17690,N_17498,N_17486);
nand U17691 (N_17691,N_17566,N_17472);
and U17692 (N_17692,N_17489,N_17516);
nor U17693 (N_17693,N_17537,N_17457);
and U17694 (N_17694,N_17438,N_17546);
and U17695 (N_17695,N_17483,N_17482);
xnor U17696 (N_17696,N_17418,N_17403);
xnor U17697 (N_17697,N_17569,N_17562);
nor U17698 (N_17698,N_17543,N_17583);
xor U17699 (N_17699,N_17443,N_17440);
nand U17700 (N_17700,N_17569,N_17504);
nor U17701 (N_17701,N_17494,N_17540);
and U17702 (N_17702,N_17596,N_17558);
or U17703 (N_17703,N_17472,N_17515);
nand U17704 (N_17704,N_17434,N_17478);
nand U17705 (N_17705,N_17424,N_17566);
nand U17706 (N_17706,N_17410,N_17479);
xor U17707 (N_17707,N_17437,N_17538);
and U17708 (N_17708,N_17510,N_17491);
nand U17709 (N_17709,N_17435,N_17539);
and U17710 (N_17710,N_17444,N_17530);
or U17711 (N_17711,N_17403,N_17573);
xnor U17712 (N_17712,N_17527,N_17575);
and U17713 (N_17713,N_17487,N_17594);
or U17714 (N_17714,N_17552,N_17462);
or U17715 (N_17715,N_17408,N_17476);
nor U17716 (N_17716,N_17429,N_17527);
xnor U17717 (N_17717,N_17457,N_17548);
or U17718 (N_17718,N_17530,N_17403);
or U17719 (N_17719,N_17447,N_17505);
nor U17720 (N_17720,N_17417,N_17559);
nor U17721 (N_17721,N_17547,N_17404);
nor U17722 (N_17722,N_17406,N_17592);
xnor U17723 (N_17723,N_17473,N_17424);
nand U17724 (N_17724,N_17536,N_17520);
and U17725 (N_17725,N_17485,N_17499);
and U17726 (N_17726,N_17456,N_17536);
nor U17727 (N_17727,N_17416,N_17411);
and U17728 (N_17728,N_17565,N_17535);
xnor U17729 (N_17729,N_17546,N_17474);
xnor U17730 (N_17730,N_17445,N_17567);
or U17731 (N_17731,N_17585,N_17402);
nor U17732 (N_17732,N_17562,N_17583);
xnor U17733 (N_17733,N_17412,N_17487);
or U17734 (N_17734,N_17583,N_17485);
nor U17735 (N_17735,N_17501,N_17456);
or U17736 (N_17736,N_17445,N_17465);
or U17737 (N_17737,N_17560,N_17417);
and U17738 (N_17738,N_17468,N_17521);
or U17739 (N_17739,N_17530,N_17482);
nor U17740 (N_17740,N_17464,N_17596);
xor U17741 (N_17741,N_17436,N_17405);
xor U17742 (N_17742,N_17444,N_17454);
nand U17743 (N_17743,N_17555,N_17594);
and U17744 (N_17744,N_17559,N_17493);
xor U17745 (N_17745,N_17502,N_17596);
and U17746 (N_17746,N_17453,N_17412);
and U17747 (N_17747,N_17578,N_17567);
nor U17748 (N_17748,N_17578,N_17518);
and U17749 (N_17749,N_17414,N_17576);
xnor U17750 (N_17750,N_17443,N_17555);
nor U17751 (N_17751,N_17406,N_17449);
xor U17752 (N_17752,N_17490,N_17515);
nor U17753 (N_17753,N_17416,N_17596);
nand U17754 (N_17754,N_17545,N_17491);
or U17755 (N_17755,N_17435,N_17528);
and U17756 (N_17756,N_17523,N_17420);
xnor U17757 (N_17757,N_17421,N_17422);
nand U17758 (N_17758,N_17472,N_17560);
nor U17759 (N_17759,N_17443,N_17433);
and U17760 (N_17760,N_17437,N_17526);
nand U17761 (N_17761,N_17495,N_17481);
nand U17762 (N_17762,N_17461,N_17508);
nand U17763 (N_17763,N_17598,N_17518);
or U17764 (N_17764,N_17443,N_17439);
and U17765 (N_17765,N_17545,N_17544);
xnor U17766 (N_17766,N_17519,N_17585);
nor U17767 (N_17767,N_17538,N_17489);
nand U17768 (N_17768,N_17441,N_17426);
or U17769 (N_17769,N_17430,N_17431);
nand U17770 (N_17770,N_17578,N_17450);
nand U17771 (N_17771,N_17508,N_17478);
or U17772 (N_17772,N_17404,N_17474);
nand U17773 (N_17773,N_17543,N_17593);
and U17774 (N_17774,N_17576,N_17426);
nand U17775 (N_17775,N_17510,N_17408);
xnor U17776 (N_17776,N_17504,N_17499);
nand U17777 (N_17777,N_17540,N_17570);
and U17778 (N_17778,N_17420,N_17423);
nor U17779 (N_17779,N_17538,N_17507);
nor U17780 (N_17780,N_17479,N_17539);
xnor U17781 (N_17781,N_17416,N_17409);
nand U17782 (N_17782,N_17401,N_17594);
and U17783 (N_17783,N_17470,N_17400);
and U17784 (N_17784,N_17502,N_17455);
nand U17785 (N_17785,N_17485,N_17441);
and U17786 (N_17786,N_17540,N_17403);
nor U17787 (N_17787,N_17529,N_17528);
xor U17788 (N_17788,N_17479,N_17532);
xor U17789 (N_17789,N_17433,N_17447);
and U17790 (N_17790,N_17471,N_17551);
nand U17791 (N_17791,N_17583,N_17436);
xor U17792 (N_17792,N_17542,N_17511);
nand U17793 (N_17793,N_17461,N_17436);
nand U17794 (N_17794,N_17519,N_17590);
nor U17795 (N_17795,N_17590,N_17544);
or U17796 (N_17796,N_17494,N_17575);
nand U17797 (N_17797,N_17554,N_17529);
nor U17798 (N_17798,N_17416,N_17417);
xor U17799 (N_17799,N_17409,N_17414);
nand U17800 (N_17800,N_17737,N_17689);
nor U17801 (N_17801,N_17713,N_17746);
nor U17802 (N_17802,N_17678,N_17655);
nor U17803 (N_17803,N_17609,N_17602);
nand U17804 (N_17804,N_17624,N_17721);
nor U17805 (N_17805,N_17762,N_17675);
and U17806 (N_17806,N_17622,N_17660);
and U17807 (N_17807,N_17674,N_17728);
nor U17808 (N_17808,N_17668,N_17638);
xnor U17809 (N_17809,N_17779,N_17766);
or U17810 (N_17810,N_17783,N_17724);
or U17811 (N_17811,N_17774,N_17697);
nor U17812 (N_17812,N_17676,N_17742);
nor U17813 (N_17813,N_17773,N_17791);
and U17814 (N_17814,N_17753,N_17665);
xor U17815 (N_17815,N_17680,N_17782);
nand U17816 (N_17816,N_17714,N_17743);
or U17817 (N_17817,N_17701,N_17726);
xor U17818 (N_17818,N_17629,N_17751);
xnor U17819 (N_17819,N_17606,N_17610);
nor U17820 (N_17820,N_17649,N_17672);
nor U17821 (N_17821,N_17772,N_17667);
xor U17822 (N_17822,N_17662,N_17718);
or U17823 (N_17823,N_17699,N_17770);
or U17824 (N_17824,N_17748,N_17647);
and U17825 (N_17825,N_17691,N_17631);
nand U17826 (N_17826,N_17696,N_17789);
nor U17827 (N_17827,N_17763,N_17636);
xor U17828 (N_17828,N_17669,N_17634);
nand U17829 (N_17829,N_17603,N_17776);
nand U17830 (N_17830,N_17716,N_17758);
or U17831 (N_17831,N_17797,N_17684);
xnor U17832 (N_17832,N_17729,N_17652);
xnor U17833 (N_17833,N_17614,N_17605);
nand U17834 (N_17834,N_17788,N_17679);
xor U17835 (N_17835,N_17759,N_17657);
xor U17836 (N_17836,N_17687,N_17641);
nand U17837 (N_17837,N_17769,N_17646);
nor U17838 (N_17838,N_17709,N_17673);
xnor U17839 (N_17839,N_17607,N_17658);
and U17840 (N_17840,N_17741,N_17794);
nand U17841 (N_17841,N_17664,N_17786);
nor U17842 (N_17842,N_17640,N_17739);
and U17843 (N_17843,N_17711,N_17752);
nand U17844 (N_17844,N_17621,N_17677);
nor U17845 (N_17845,N_17616,N_17637);
and U17846 (N_17846,N_17639,N_17644);
or U17847 (N_17847,N_17686,N_17693);
or U17848 (N_17848,N_17683,N_17604);
or U17849 (N_17849,N_17666,N_17747);
nor U17850 (N_17850,N_17732,N_17702);
nand U17851 (N_17851,N_17745,N_17659);
nor U17852 (N_17852,N_17682,N_17694);
or U17853 (N_17853,N_17707,N_17777);
nand U17854 (N_17854,N_17653,N_17715);
and U17855 (N_17855,N_17651,N_17626);
or U17856 (N_17856,N_17719,N_17681);
xnor U17857 (N_17857,N_17613,N_17723);
nor U17858 (N_17858,N_17784,N_17744);
xnor U17859 (N_17859,N_17738,N_17688);
nor U17860 (N_17860,N_17725,N_17760);
nor U17861 (N_17861,N_17780,N_17731);
nor U17862 (N_17862,N_17625,N_17690);
nor U17863 (N_17863,N_17740,N_17757);
and U17864 (N_17864,N_17617,N_17787);
nor U17865 (N_17865,N_17685,N_17648);
nor U17866 (N_17866,N_17643,N_17645);
xor U17867 (N_17867,N_17730,N_17799);
or U17868 (N_17868,N_17671,N_17695);
nor U17869 (N_17869,N_17735,N_17733);
or U17870 (N_17870,N_17619,N_17754);
and U17871 (N_17871,N_17749,N_17771);
nand U17872 (N_17872,N_17736,N_17795);
or U17873 (N_17873,N_17663,N_17705);
nand U17874 (N_17874,N_17755,N_17708);
or U17875 (N_17875,N_17670,N_17722);
and U17876 (N_17876,N_17790,N_17700);
nor U17877 (N_17877,N_17628,N_17781);
xor U17878 (N_17878,N_17734,N_17775);
nand U17879 (N_17879,N_17623,N_17717);
xor U17880 (N_17880,N_17704,N_17750);
or U17881 (N_17881,N_17632,N_17608);
xnor U17882 (N_17882,N_17698,N_17656);
or U17883 (N_17883,N_17620,N_17720);
nand U17884 (N_17884,N_17765,N_17756);
or U17885 (N_17885,N_17633,N_17710);
nand U17886 (N_17886,N_17654,N_17650);
and U17887 (N_17887,N_17703,N_17692);
nand U17888 (N_17888,N_17761,N_17785);
nor U17889 (N_17889,N_17635,N_17661);
or U17890 (N_17890,N_17792,N_17727);
and U17891 (N_17891,N_17601,N_17612);
and U17892 (N_17892,N_17764,N_17630);
xnor U17893 (N_17893,N_17712,N_17796);
nand U17894 (N_17894,N_17618,N_17706);
or U17895 (N_17895,N_17615,N_17642);
and U17896 (N_17896,N_17611,N_17627);
nor U17897 (N_17897,N_17793,N_17778);
and U17898 (N_17898,N_17798,N_17767);
nand U17899 (N_17899,N_17768,N_17600);
or U17900 (N_17900,N_17684,N_17678);
and U17901 (N_17901,N_17644,N_17731);
or U17902 (N_17902,N_17779,N_17659);
xor U17903 (N_17903,N_17789,N_17671);
nand U17904 (N_17904,N_17724,N_17717);
nor U17905 (N_17905,N_17611,N_17610);
or U17906 (N_17906,N_17670,N_17647);
and U17907 (N_17907,N_17659,N_17630);
nand U17908 (N_17908,N_17609,N_17711);
xnor U17909 (N_17909,N_17657,N_17770);
nor U17910 (N_17910,N_17755,N_17740);
or U17911 (N_17911,N_17799,N_17766);
nor U17912 (N_17912,N_17649,N_17627);
or U17913 (N_17913,N_17780,N_17702);
xor U17914 (N_17914,N_17700,N_17651);
nand U17915 (N_17915,N_17780,N_17718);
or U17916 (N_17916,N_17782,N_17729);
xnor U17917 (N_17917,N_17685,N_17686);
or U17918 (N_17918,N_17789,N_17618);
nor U17919 (N_17919,N_17772,N_17746);
xnor U17920 (N_17920,N_17630,N_17799);
nor U17921 (N_17921,N_17685,N_17703);
and U17922 (N_17922,N_17637,N_17796);
nand U17923 (N_17923,N_17616,N_17651);
nor U17924 (N_17924,N_17616,N_17782);
and U17925 (N_17925,N_17623,N_17642);
xnor U17926 (N_17926,N_17671,N_17726);
nand U17927 (N_17927,N_17793,N_17691);
nand U17928 (N_17928,N_17683,N_17789);
nand U17929 (N_17929,N_17633,N_17777);
nor U17930 (N_17930,N_17743,N_17724);
nor U17931 (N_17931,N_17750,N_17689);
or U17932 (N_17932,N_17653,N_17612);
or U17933 (N_17933,N_17780,N_17755);
and U17934 (N_17934,N_17751,N_17795);
or U17935 (N_17935,N_17619,N_17692);
or U17936 (N_17936,N_17621,N_17639);
xnor U17937 (N_17937,N_17677,N_17653);
nand U17938 (N_17938,N_17678,N_17742);
and U17939 (N_17939,N_17715,N_17746);
nand U17940 (N_17940,N_17735,N_17692);
or U17941 (N_17941,N_17718,N_17735);
or U17942 (N_17942,N_17680,N_17603);
nor U17943 (N_17943,N_17769,N_17689);
nor U17944 (N_17944,N_17676,N_17696);
nor U17945 (N_17945,N_17601,N_17770);
and U17946 (N_17946,N_17715,N_17648);
and U17947 (N_17947,N_17661,N_17792);
or U17948 (N_17948,N_17614,N_17677);
and U17949 (N_17949,N_17680,N_17788);
xnor U17950 (N_17950,N_17736,N_17786);
or U17951 (N_17951,N_17628,N_17744);
nand U17952 (N_17952,N_17606,N_17755);
nor U17953 (N_17953,N_17664,N_17646);
nor U17954 (N_17954,N_17607,N_17752);
or U17955 (N_17955,N_17638,N_17714);
and U17956 (N_17956,N_17606,N_17727);
nand U17957 (N_17957,N_17702,N_17616);
nor U17958 (N_17958,N_17797,N_17643);
or U17959 (N_17959,N_17756,N_17607);
xor U17960 (N_17960,N_17615,N_17772);
nand U17961 (N_17961,N_17785,N_17762);
and U17962 (N_17962,N_17654,N_17772);
nand U17963 (N_17963,N_17606,N_17624);
nand U17964 (N_17964,N_17743,N_17723);
and U17965 (N_17965,N_17702,N_17697);
xor U17966 (N_17966,N_17785,N_17615);
nor U17967 (N_17967,N_17653,N_17627);
nand U17968 (N_17968,N_17624,N_17664);
or U17969 (N_17969,N_17647,N_17792);
or U17970 (N_17970,N_17745,N_17763);
nand U17971 (N_17971,N_17679,N_17704);
xor U17972 (N_17972,N_17676,N_17747);
nand U17973 (N_17973,N_17796,N_17635);
or U17974 (N_17974,N_17767,N_17771);
xor U17975 (N_17975,N_17768,N_17609);
nand U17976 (N_17976,N_17703,N_17604);
nor U17977 (N_17977,N_17684,N_17772);
xnor U17978 (N_17978,N_17753,N_17770);
xor U17979 (N_17979,N_17648,N_17753);
or U17980 (N_17980,N_17730,N_17764);
nor U17981 (N_17981,N_17678,N_17797);
and U17982 (N_17982,N_17610,N_17779);
or U17983 (N_17983,N_17658,N_17676);
and U17984 (N_17984,N_17725,N_17780);
and U17985 (N_17985,N_17771,N_17725);
or U17986 (N_17986,N_17760,N_17609);
nor U17987 (N_17987,N_17613,N_17752);
and U17988 (N_17988,N_17783,N_17664);
nor U17989 (N_17989,N_17670,N_17773);
nand U17990 (N_17990,N_17628,N_17677);
or U17991 (N_17991,N_17718,N_17698);
and U17992 (N_17992,N_17632,N_17633);
and U17993 (N_17993,N_17749,N_17704);
nand U17994 (N_17994,N_17773,N_17701);
xnor U17995 (N_17995,N_17768,N_17780);
nand U17996 (N_17996,N_17619,N_17638);
nor U17997 (N_17997,N_17791,N_17686);
nand U17998 (N_17998,N_17727,N_17711);
nor U17999 (N_17999,N_17705,N_17643);
xnor U18000 (N_18000,N_17832,N_17998);
nand U18001 (N_18001,N_17954,N_17824);
nand U18002 (N_18002,N_17801,N_17976);
nand U18003 (N_18003,N_17928,N_17904);
or U18004 (N_18004,N_17988,N_17962);
and U18005 (N_18005,N_17938,N_17885);
xnor U18006 (N_18006,N_17845,N_17987);
nand U18007 (N_18007,N_17808,N_17830);
or U18008 (N_18008,N_17944,N_17929);
nor U18009 (N_18009,N_17868,N_17945);
xor U18010 (N_18010,N_17896,N_17927);
or U18011 (N_18011,N_17936,N_17970);
or U18012 (N_18012,N_17917,N_17865);
xnor U18013 (N_18013,N_17841,N_17992);
and U18014 (N_18014,N_17932,N_17930);
and U18015 (N_18015,N_17946,N_17913);
and U18016 (N_18016,N_17809,N_17922);
and U18017 (N_18017,N_17819,N_17924);
xnor U18018 (N_18018,N_17852,N_17800);
nor U18019 (N_18019,N_17853,N_17862);
and U18020 (N_18020,N_17827,N_17958);
nand U18021 (N_18021,N_17948,N_17934);
nand U18022 (N_18022,N_17919,N_17842);
nand U18023 (N_18023,N_17906,N_17811);
or U18024 (N_18024,N_17940,N_17815);
nand U18025 (N_18025,N_17964,N_17876);
or U18026 (N_18026,N_17912,N_17818);
xor U18027 (N_18027,N_17820,N_17953);
nand U18028 (N_18028,N_17895,N_17967);
or U18029 (N_18029,N_17875,N_17975);
nor U18030 (N_18030,N_17918,N_17880);
and U18031 (N_18031,N_17979,N_17869);
or U18032 (N_18032,N_17963,N_17826);
nor U18033 (N_18033,N_17923,N_17961);
xnor U18034 (N_18034,N_17996,N_17846);
xor U18035 (N_18035,N_17866,N_17851);
and U18036 (N_18036,N_17803,N_17839);
or U18037 (N_18037,N_17882,N_17854);
and U18038 (N_18038,N_17955,N_17823);
xor U18039 (N_18039,N_17864,N_17920);
nor U18040 (N_18040,N_17831,N_17921);
xnor U18041 (N_18041,N_17931,N_17925);
nand U18042 (N_18042,N_17995,N_17994);
and U18043 (N_18043,N_17933,N_17806);
and U18044 (N_18044,N_17802,N_17914);
or U18045 (N_18045,N_17881,N_17903);
xnor U18046 (N_18046,N_17935,N_17833);
xor U18047 (N_18047,N_17890,N_17843);
or U18048 (N_18048,N_17951,N_17942);
nand U18049 (N_18049,N_17829,N_17887);
or U18050 (N_18050,N_17861,N_17997);
nor U18051 (N_18051,N_17937,N_17817);
xor U18052 (N_18052,N_17835,N_17857);
nand U18053 (N_18053,N_17888,N_17898);
and U18054 (N_18054,N_17891,N_17879);
and U18055 (N_18055,N_17863,N_17804);
xor U18056 (N_18056,N_17949,N_17980);
nor U18057 (N_18057,N_17971,N_17969);
and U18058 (N_18058,N_17900,N_17989);
or U18059 (N_18059,N_17821,N_17825);
and U18060 (N_18060,N_17978,N_17897);
and U18061 (N_18061,N_17907,N_17855);
nor U18062 (N_18062,N_17894,N_17959);
or U18063 (N_18063,N_17834,N_17947);
nand U18064 (N_18064,N_17972,N_17816);
and U18065 (N_18065,N_17836,N_17849);
xnor U18066 (N_18066,N_17844,N_17981);
nand U18067 (N_18067,N_17973,N_17941);
nor U18068 (N_18068,N_17915,N_17822);
nor U18069 (N_18069,N_17828,N_17990);
nor U18070 (N_18070,N_17966,N_17986);
nor U18071 (N_18071,N_17871,N_17874);
and U18072 (N_18072,N_17837,N_17840);
or U18073 (N_18073,N_17977,N_17950);
and U18074 (N_18074,N_17867,N_17884);
or U18075 (N_18075,N_17858,N_17902);
nor U18076 (N_18076,N_17965,N_17993);
nor U18077 (N_18077,N_17901,N_17982);
or U18078 (N_18078,N_17859,N_17985);
xnor U18079 (N_18079,N_17908,N_17910);
nand U18080 (N_18080,N_17916,N_17984);
nor U18081 (N_18081,N_17968,N_17999);
or U18082 (N_18082,N_17856,N_17893);
or U18083 (N_18083,N_17892,N_17956);
nand U18084 (N_18084,N_17807,N_17943);
xnor U18085 (N_18085,N_17926,N_17878);
nand U18086 (N_18086,N_17991,N_17860);
and U18087 (N_18087,N_17848,N_17813);
nor U18088 (N_18088,N_17810,N_17957);
or U18089 (N_18089,N_17974,N_17838);
nor U18090 (N_18090,N_17886,N_17850);
nor U18091 (N_18091,N_17877,N_17909);
nor U18092 (N_18092,N_17983,N_17939);
nand U18093 (N_18093,N_17905,N_17911);
nor U18094 (N_18094,N_17814,N_17883);
xor U18095 (N_18095,N_17873,N_17952);
nand U18096 (N_18096,N_17889,N_17812);
nand U18097 (N_18097,N_17847,N_17805);
nor U18098 (N_18098,N_17872,N_17960);
or U18099 (N_18099,N_17870,N_17899);
or U18100 (N_18100,N_17844,N_17984);
and U18101 (N_18101,N_17865,N_17905);
nor U18102 (N_18102,N_17870,N_17882);
nand U18103 (N_18103,N_17972,N_17856);
or U18104 (N_18104,N_17952,N_17831);
nor U18105 (N_18105,N_17814,N_17889);
or U18106 (N_18106,N_17980,N_17906);
xnor U18107 (N_18107,N_17822,N_17974);
nor U18108 (N_18108,N_17830,N_17965);
or U18109 (N_18109,N_17946,N_17866);
nand U18110 (N_18110,N_17890,N_17923);
and U18111 (N_18111,N_17980,N_17808);
nor U18112 (N_18112,N_17862,N_17932);
nand U18113 (N_18113,N_17861,N_17932);
or U18114 (N_18114,N_17967,N_17884);
nand U18115 (N_18115,N_17949,N_17866);
nor U18116 (N_18116,N_17962,N_17915);
nor U18117 (N_18117,N_17803,N_17866);
nand U18118 (N_18118,N_17858,N_17914);
nand U18119 (N_18119,N_17971,N_17857);
or U18120 (N_18120,N_17933,N_17839);
or U18121 (N_18121,N_17837,N_17856);
and U18122 (N_18122,N_17890,N_17812);
or U18123 (N_18123,N_17995,N_17939);
or U18124 (N_18124,N_17850,N_17953);
nor U18125 (N_18125,N_17878,N_17911);
or U18126 (N_18126,N_17854,N_17881);
nand U18127 (N_18127,N_17845,N_17815);
and U18128 (N_18128,N_17927,N_17867);
nand U18129 (N_18129,N_17966,N_17821);
xor U18130 (N_18130,N_17854,N_17888);
xnor U18131 (N_18131,N_17953,N_17861);
xor U18132 (N_18132,N_17854,N_17945);
and U18133 (N_18133,N_17842,N_17872);
nor U18134 (N_18134,N_17900,N_17816);
nand U18135 (N_18135,N_17949,N_17906);
xor U18136 (N_18136,N_17914,N_17889);
nand U18137 (N_18137,N_17930,N_17975);
and U18138 (N_18138,N_17930,N_17858);
and U18139 (N_18139,N_17891,N_17905);
and U18140 (N_18140,N_17963,N_17994);
and U18141 (N_18141,N_17966,N_17935);
or U18142 (N_18142,N_17832,N_17899);
and U18143 (N_18143,N_17922,N_17911);
nor U18144 (N_18144,N_17912,N_17902);
and U18145 (N_18145,N_17985,N_17904);
nor U18146 (N_18146,N_17844,N_17863);
xor U18147 (N_18147,N_17926,N_17820);
xnor U18148 (N_18148,N_17820,N_17914);
and U18149 (N_18149,N_17964,N_17918);
nand U18150 (N_18150,N_17943,N_17855);
nor U18151 (N_18151,N_17881,N_17891);
or U18152 (N_18152,N_17842,N_17817);
nor U18153 (N_18153,N_17806,N_17909);
xor U18154 (N_18154,N_17928,N_17845);
nor U18155 (N_18155,N_17812,N_17968);
nand U18156 (N_18156,N_17839,N_17909);
nand U18157 (N_18157,N_17857,N_17802);
xor U18158 (N_18158,N_17946,N_17910);
nand U18159 (N_18159,N_17981,N_17951);
nor U18160 (N_18160,N_17891,N_17819);
xor U18161 (N_18161,N_17927,N_17956);
nor U18162 (N_18162,N_17979,N_17893);
or U18163 (N_18163,N_17961,N_17871);
nand U18164 (N_18164,N_17897,N_17937);
and U18165 (N_18165,N_17828,N_17963);
and U18166 (N_18166,N_17815,N_17995);
or U18167 (N_18167,N_17877,N_17982);
nand U18168 (N_18168,N_17891,N_17848);
xor U18169 (N_18169,N_17819,N_17946);
xnor U18170 (N_18170,N_17936,N_17943);
nand U18171 (N_18171,N_17992,N_17922);
nor U18172 (N_18172,N_17837,N_17847);
nand U18173 (N_18173,N_17853,N_17851);
xor U18174 (N_18174,N_17909,N_17903);
nor U18175 (N_18175,N_17898,N_17935);
nand U18176 (N_18176,N_17985,N_17911);
and U18177 (N_18177,N_17906,N_17817);
nor U18178 (N_18178,N_17827,N_17819);
and U18179 (N_18179,N_17906,N_17816);
nand U18180 (N_18180,N_17835,N_17818);
xor U18181 (N_18181,N_17969,N_17928);
nand U18182 (N_18182,N_17813,N_17831);
or U18183 (N_18183,N_17886,N_17884);
xor U18184 (N_18184,N_17862,N_17887);
xor U18185 (N_18185,N_17968,N_17945);
and U18186 (N_18186,N_17999,N_17860);
and U18187 (N_18187,N_17949,N_17991);
or U18188 (N_18188,N_17940,N_17816);
nand U18189 (N_18189,N_17839,N_17990);
xor U18190 (N_18190,N_17836,N_17954);
nand U18191 (N_18191,N_17891,N_17857);
or U18192 (N_18192,N_17934,N_17968);
or U18193 (N_18193,N_17991,N_17849);
and U18194 (N_18194,N_17919,N_17812);
xnor U18195 (N_18195,N_17937,N_17950);
or U18196 (N_18196,N_17976,N_17894);
or U18197 (N_18197,N_17962,N_17833);
nand U18198 (N_18198,N_17981,N_17916);
nand U18199 (N_18199,N_17877,N_17808);
and U18200 (N_18200,N_18036,N_18051);
or U18201 (N_18201,N_18035,N_18162);
and U18202 (N_18202,N_18168,N_18092);
xor U18203 (N_18203,N_18049,N_18136);
and U18204 (N_18204,N_18046,N_18074);
xnor U18205 (N_18205,N_18126,N_18000);
nand U18206 (N_18206,N_18073,N_18013);
or U18207 (N_18207,N_18056,N_18159);
and U18208 (N_18208,N_18101,N_18192);
or U18209 (N_18209,N_18132,N_18009);
nand U18210 (N_18210,N_18189,N_18131);
xnor U18211 (N_18211,N_18169,N_18139);
nor U18212 (N_18212,N_18187,N_18118);
xnor U18213 (N_18213,N_18119,N_18019);
xor U18214 (N_18214,N_18174,N_18086);
or U18215 (N_18215,N_18135,N_18180);
nand U18216 (N_18216,N_18157,N_18137);
nand U18217 (N_18217,N_18113,N_18146);
or U18218 (N_18218,N_18178,N_18059);
xor U18219 (N_18219,N_18020,N_18143);
or U18220 (N_18220,N_18140,N_18007);
nand U18221 (N_18221,N_18130,N_18015);
nor U18222 (N_18222,N_18129,N_18199);
nor U18223 (N_18223,N_18028,N_18018);
xor U18224 (N_18224,N_18097,N_18164);
and U18225 (N_18225,N_18191,N_18150);
and U18226 (N_18226,N_18022,N_18183);
nand U18227 (N_18227,N_18105,N_18186);
xor U18228 (N_18228,N_18050,N_18011);
nor U18229 (N_18229,N_18032,N_18195);
nor U18230 (N_18230,N_18003,N_18002);
nand U18231 (N_18231,N_18190,N_18027);
and U18232 (N_18232,N_18075,N_18024);
nor U18233 (N_18233,N_18038,N_18081);
nor U18234 (N_18234,N_18098,N_18179);
xor U18235 (N_18235,N_18005,N_18054);
or U18236 (N_18236,N_18172,N_18084);
or U18237 (N_18237,N_18034,N_18196);
and U18238 (N_18238,N_18001,N_18182);
and U18239 (N_18239,N_18091,N_18184);
xnor U18240 (N_18240,N_18144,N_18112);
nor U18241 (N_18241,N_18111,N_18043);
or U18242 (N_18242,N_18173,N_18044);
nor U18243 (N_18243,N_18156,N_18153);
xor U18244 (N_18244,N_18099,N_18110);
xor U18245 (N_18245,N_18052,N_18181);
xor U18246 (N_18246,N_18088,N_18171);
xor U18247 (N_18247,N_18014,N_18042);
xor U18248 (N_18248,N_18021,N_18039);
and U18249 (N_18249,N_18102,N_18069);
or U18250 (N_18250,N_18103,N_18108);
or U18251 (N_18251,N_18053,N_18040);
xor U18252 (N_18252,N_18104,N_18147);
or U18253 (N_18253,N_18100,N_18078);
xnor U18254 (N_18254,N_18083,N_18026);
nor U18255 (N_18255,N_18127,N_18116);
xnor U18256 (N_18256,N_18160,N_18010);
xnor U18257 (N_18257,N_18062,N_18148);
nor U18258 (N_18258,N_18041,N_18106);
and U18259 (N_18259,N_18058,N_18194);
or U18260 (N_18260,N_18063,N_18064);
nor U18261 (N_18261,N_18198,N_18082);
and U18262 (N_18262,N_18133,N_18166);
nand U18263 (N_18263,N_18163,N_18185);
or U18264 (N_18264,N_18017,N_18117);
nor U18265 (N_18265,N_18109,N_18176);
nor U18266 (N_18266,N_18037,N_18055);
nor U18267 (N_18267,N_18060,N_18151);
or U18268 (N_18268,N_18134,N_18167);
xnor U18269 (N_18269,N_18068,N_18142);
or U18270 (N_18270,N_18095,N_18085);
and U18271 (N_18271,N_18125,N_18066);
nor U18272 (N_18272,N_18128,N_18120);
nand U18273 (N_18273,N_18067,N_18175);
and U18274 (N_18274,N_18161,N_18107);
and U18275 (N_18275,N_18158,N_18145);
and U18276 (N_18276,N_18065,N_18030);
or U18277 (N_18277,N_18077,N_18094);
and U18278 (N_18278,N_18087,N_18029);
nor U18279 (N_18279,N_18070,N_18123);
or U18280 (N_18280,N_18072,N_18096);
nor U18281 (N_18281,N_18057,N_18177);
nand U18282 (N_18282,N_18141,N_18124);
or U18283 (N_18283,N_18154,N_18138);
nand U18284 (N_18284,N_18080,N_18025);
or U18285 (N_18285,N_18115,N_18155);
xor U18286 (N_18286,N_18048,N_18047);
xnor U18287 (N_18287,N_18122,N_18114);
or U18288 (N_18288,N_18006,N_18023);
xor U18289 (N_18289,N_18170,N_18121);
and U18290 (N_18290,N_18165,N_18004);
xor U18291 (N_18291,N_18197,N_18089);
xnor U18292 (N_18292,N_18093,N_18061);
xor U18293 (N_18293,N_18193,N_18031);
and U18294 (N_18294,N_18071,N_18033);
nor U18295 (N_18295,N_18008,N_18149);
and U18296 (N_18296,N_18090,N_18076);
or U18297 (N_18297,N_18045,N_18079);
or U18298 (N_18298,N_18016,N_18152);
xnor U18299 (N_18299,N_18188,N_18012);
nand U18300 (N_18300,N_18131,N_18196);
nor U18301 (N_18301,N_18104,N_18185);
xor U18302 (N_18302,N_18162,N_18095);
or U18303 (N_18303,N_18079,N_18081);
nor U18304 (N_18304,N_18195,N_18106);
nand U18305 (N_18305,N_18131,N_18002);
or U18306 (N_18306,N_18116,N_18175);
and U18307 (N_18307,N_18012,N_18023);
xor U18308 (N_18308,N_18097,N_18071);
nand U18309 (N_18309,N_18187,N_18025);
or U18310 (N_18310,N_18109,N_18098);
nor U18311 (N_18311,N_18001,N_18175);
nand U18312 (N_18312,N_18191,N_18147);
or U18313 (N_18313,N_18070,N_18028);
xnor U18314 (N_18314,N_18066,N_18178);
and U18315 (N_18315,N_18155,N_18141);
nand U18316 (N_18316,N_18018,N_18194);
or U18317 (N_18317,N_18123,N_18149);
nand U18318 (N_18318,N_18112,N_18099);
and U18319 (N_18319,N_18168,N_18156);
xor U18320 (N_18320,N_18159,N_18007);
or U18321 (N_18321,N_18014,N_18179);
and U18322 (N_18322,N_18003,N_18081);
nor U18323 (N_18323,N_18158,N_18192);
and U18324 (N_18324,N_18034,N_18107);
xnor U18325 (N_18325,N_18101,N_18063);
nor U18326 (N_18326,N_18113,N_18151);
and U18327 (N_18327,N_18026,N_18090);
nor U18328 (N_18328,N_18031,N_18009);
and U18329 (N_18329,N_18020,N_18151);
or U18330 (N_18330,N_18029,N_18111);
and U18331 (N_18331,N_18093,N_18081);
and U18332 (N_18332,N_18163,N_18028);
nand U18333 (N_18333,N_18158,N_18184);
or U18334 (N_18334,N_18164,N_18190);
xnor U18335 (N_18335,N_18005,N_18186);
nand U18336 (N_18336,N_18026,N_18056);
nor U18337 (N_18337,N_18022,N_18076);
xor U18338 (N_18338,N_18150,N_18110);
nand U18339 (N_18339,N_18075,N_18077);
or U18340 (N_18340,N_18006,N_18152);
nand U18341 (N_18341,N_18045,N_18007);
nand U18342 (N_18342,N_18191,N_18137);
nor U18343 (N_18343,N_18150,N_18012);
and U18344 (N_18344,N_18047,N_18194);
or U18345 (N_18345,N_18030,N_18096);
or U18346 (N_18346,N_18093,N_18089);
nor U18347 (N_18347,N_18010,N_18043);
nor U18348 (N_18348,N_18015,N_18108);
or U18349 (N_18349,N_18025,N_18061);
xnor U18350 (N_18350,N_18035,N_18109);
or U18351 (N_18351,N_18105,N_18184);
nand U18352 (N_18352,N_18152,N_18118);
or U18353 (N_18353,N_18098,N_18013);
nor U18354 (N_18354,N_18173,N_18128);
nand U18355 (N_18355,N_18089,N_18174);
nand U18356 (N_18356,N_18106,N_18093);
and U18357 (N_18357,N_18043,N_18000);
and U18358 (N_18358,N_18131,N_18147);
xor U18359 (N_18359,N_18098,N_18114);
or U18360 (N_18360,N_18047,N_18077);
nor U18361 (N_18361,N_18059,N_18011);
nor U18362 (N_18362,N_18164,N_18004);
or U18363 (N_18363,N_18157,N_18077);
nor U18364 (N_18364,N_18057,N_18059);
or U18365 (N_18365,N_18011,N_18103);
nand U18366 (N_18366,N_18049,N_18081);
xor U18367 (N_18367,N_18048,N_18136);
and U18368 (N_18368,N_18140,N_18056);
and U18369 (N_18369,N_18129,N_18034);
or U18370 (N_18370,N_18108,N_18035);
nor U18371 (N_18371,N_18184,N_18046);
xor U18372 (N_18372,N_18191,N_18038);
or U18373 (N_18373,N_18063,N_18076);
xnor U18374 (N_18374,N_18035,N_18139);
and U18375 (N_18375,N_18037,N_18109);
xnor U18376 (N_18376,N_18089,N_18141);
nand U18377 (N_18377,N_18130,N_18055);
or U18378 (N_18378,N_18083,N_18022);
or U18379 (N_18379,N_18115,N_18099);
xor U18380 (N_18380,N_18128,N_18105);
nand U18381 (N_18381,N_18122,N_18123);
and U18382 (N_18382,N_18049,N_18148);
and U18383 (N_18383,N_18133,N_18073);
nand U18384 (N_18384,N_18167,N_18163);
nor U18385 (N_18385,N_18074,N_18087);
or U18386 (N_18386,N_18076,N_18068);
or U18387 (N_18387,N_18114,N_18174);
xnor U18388 (N_18388,N_18006,N_18180);
nor U18389 (N_18389,N_18096,N_18179);
nand U18390 (N_18390,N_18197,N_18195);
and U18391 (N_18391,N_18143,N_18104);
nand U18392 (N_18392,N_18049,N_18111);
xor U18393 (N_18393,N_18190,N_18081);
or U18394 (N_18394,N_18077,N_18108);
or U18395 (N_18395,N_18170,N_18142);
nor U18396 (N_18396,N_18110,N_18141);
xor U18397 (N_18397,N_18175,N_18006);
xor U18398 (N_18398,N_18153,N_18144);
xnor U18399 (N_18399,N_18017,N_18116);
and U18400 (N_18400,N_18300,N_18359);
nor U18401 (N_18401,N_18319,N_18219);
and U18402 (N_18402,N_18345,N_18309);
xnor U18403 (N_18403,N_18387,N_18312);
and U18404 (N_18404,N_18358,N_18342);
xor U18405 (N_18405,N_18231,N_18240);
and U18406 (N_18406,N_18390,N_18241);
and U18407 (N_18407,N_18268,N_18378);
xnor U18408 (N_18408,N_18396,N_18281);
nor U18409 (N_18409,N_18311,N_18326);
xor U18410 (N_18410,N_18234,N_18242);
and U18411 (N_18411,N_18363,N_18392);
nand U18412 (N_18412,N_18343,N_18391);
xor U18413 (N_18413,N_18205,N_18285);
and U18414 (N_18414,N_18291,N_18226);
or U18415 (N_18415,N_18244,N_18385);
nor U18416 (N_18416,N_18274,N_18246);
nand U18417 (N_18417,N_18207,N_18284);
or U18418 (N_18418,N_18341,N_18365);
nand U18419 (N_18419,N_18263,N_18315);
or U18420 (N_18420,N_18289,N_18377);
nand U18421 (N_18421,N_18213,N_18208);
xnor U18422 (N_18422,N_18397,N_18203);
and U18423 (N_18423,N_18376,N_18347);
xnor U18424 (N_18424,N_18354,N_18248);
xnor U18425 (N_18425,N_18250,N_18296);
or U18426 (N_18426,N_18221,N_18249);
xnor U18427 (N_18427,N_18295,N_18277);
nand U18428 (N_18428,N_18338,N_18200);
xor U18429 (N_18429,N_18283,N_18384);
nand U18430 (N_18430,N_18202,N_18353);
nand U18431 (N_18431,N_18352,N_18371);
nand U18432 (N_18432,N_18303,N_18273);
nand U18433 (N_18433,N_18317,N_18212);
nor U18434 (N_18434,N_18238,N_18237);
and U18435 (N_18435,N_18394,N_18298);
and U18436 (N_18436,N_18366,N_18262);
or U18437 (N_18437,N_18252,N_18267);
or U18438 (N_18438,N_18220,N_18333);
or U18439 (N_18439,N_18388,N_18236);
and U18440 (N_18440,N_18339,N_18305);
and U18441 (N_18441,N_18386,N_18239);
nand U18442 (N_18442,N_18201,N_18233);
nand U18443 (N_18443,N_18367,N_18322);
or U18444 (N_18444,N_18292,N_18313);
nand U18445 (N_18445,N_18350,N_18258);
and U18446 (N_18446,N_18224,N_18278);
nand U18447 (N_18447,N_18355,N_18362);
nor U18448 (N_18448,N_18370,N_18294);
nand U18449 (N_18449,N_18379,N_18327);
nor U18450 (N_18450,N_18218,N_18368);
xor U18451 (N_18451,N_18308,N_18318);
nor U18452 (N_18452,N_18253,N_18310);
and U18453 (N_18453,N_18323,N_18225);
and U18454 (N_18454,N_18351,N_18314);
nor U18455 (N_18455,N_18395,N_18369);
or U18456 (N_18456,N_18266,N_18216);
nand U18457 (N_18457,N_18229,N_18331);
or U18458 (N_18458,N_18316,N_18275);
nand U18459 (N_18459,N_18375,N_18324);
xor U18460 (N_18460,N_18286,N_18280);
nor U18461 (N_18461,N_18301,N_18257);
or U18462 (N_18462,N_18206,N_18264);
or U18463 (N_18463,N_18336,N_18265);
and U18464 (N_18464,N_18255,N_18306);
and U18465 (N_18465,N_18214,N_18382);
or U18466 (N_18466,N_18349,N_18389);
nand U18467 (N_18467,N_18210,N_18293);
and U18468 (N_18468,N_18256,N_18361);
nor U18469 (N_18469,N_18399,N_18230);
nor U18470 (N_18470,N_18380,N_18383);
xor U18471 (N_18471,N_18271,N_18259);
nor U18472 (N_18472,N_18254,N_18251);
nand U18473 (N_18473,N_18276,N_18243);
nor U18474 (N_18474,N_18381,N_18282);
nand U18475 (N_18475,N_18344,N_18332);
xnor U18476 (N_18476,N_18227,N_18325);
nand U18477 (N_18477,N_18287,N_18334);
nor U18478 (N_18478,N_18337,N_18288);
xor U18479 (N_18479,N_18348,N_18245);
nor U18480 (N_18480,N_18235,N_18304);
nor U18481 (N_18481,N_18223,N_18260);
and U18482 (N_18482,N_18222,N_18374);
xor U18483 (N_18483,N_18328,N_18372);
and U18484 (N_18484,N_18320,N_18335);
or U18485 (N_18485,N_18340,N_18217);
xor U18486 (N_18486,N_18302,N_18228);
or U18487 (N_18487,N_18321,N_18307);
nor U18488 (N_18488,N_18204,N_18299);
or U18489 (N_18489,N_18398,N_18356);
or U18490 (N_18490,N_18297,N_18329);
nand U18491 (N_18491,N_18360,N_18272);
xor U18492 (N_18492,N_18357,N_18261);
nor U18493 (N_18493,N_18270,N_18269);
and U18494 (N_18494,N_18373,N_18247);
and U18495 (N_18495,N_18211,N_18279);
xor U18496 (N_18496,N_18393,N_18215);
and U18497 (N_18497,N_18232,N_18346);
nand U18498 (N_18498,N_18330,N_18364);
or U18499 (N_18499,N_18209,N_18290);
nand U18500 (N_18500,N_18234,N_18239);
or U18501 (N_18501,N_18212,N_18311);
and U18502 (N_18502,N_18310,N_18247);
nor U18503 (N_18503,N_18394,N_18396);
and U18504 (N_18504,N_18316,N_18347);
nor U18505 (N_18505,N_18292,N_18252);
nor U18506 (N_18506,N_18258,N_18339);
or U18507 (N_18507,N_18221,N_18380);
or U18508 (N_18508,N_18260,N_18297);
and U18509 (N_18509,N_18390,N_18331);
nor U18510 (N_18510,N_18211,N_18217);
or U18511 (N_18511,N_18384,N_18355);
and U18512 (N_18512,N_18338,N_18272);
or U18513 (N_18513,N_18273,N_18343);
nand U18514 (N_18514,N_18309,N_18332);
or U18515 (N_18515,N_18374,N_18292);
nand U18516 (N_18516,N_18285,N_18309);
and U18517 (N_18517,N_18352,N_18205);
nor U18518 (N_18518,N_18224,N_18336);
xor U18519 (N_18519,N_18382,N_18221);
xor U18520 (N_18520,N_18310,N_18258);
or U18521 (N_18521,N_18285,N_18354);
and U18522 (N_18522,N_18328,N_18267);
and U18523 (N_18523,N_18396,N_18219);
nor U18524 (N_18524,N_18332,N_18291);
nor U18525 (N_18525,N_18249,N_18312);
nor U18526 (N_18526,N_18200,N_18212);
or U18527 (N_18527,N_18253,N_18235);
nor U18528 (N_18528,N_18274,N_18223);
nor U18529 (N_18529,N_18266,N_18372);
nor U18530 (N_18530,N_18243,N_18299);
nor U18531 (N_18531,N_18361,N_18321);
or U18532 (N_18532,N_18214,N_18314);
or U18533 (N_18533,N_18323,N_18218);
xnor U18534 (N_18534,N_18315,N_18201);
or U18535 (N_18535,N_18236,N_18229);
nor U18536 (N_18536,N_18252,N_18289);
and U18537 (N_18537,N_18249,N_18315);
or U18538 (N_18538,N_18288,N_18246);
and U18539 (N_18539,N_18301,N_18233);
xnor U18540 (N_18540,N_18320,N_18276);
xor U18541 (N_18541,N_18334,N_18298);
and U18542 (N_18542,N_18216,N_18350);
or U18543 (N_18543,N_18204,N_18205);
and U18544 (N_18544,N_18264,N_18318);
and U18545 (N_18545,N_18249,N_18336);
nand U18546 (N_18546,N_18202,N_18344);
xor U18547 (N_18547,N_18362,N_18327);
and U18548 (N_18548,N_18277,N_18356);
and U18549 (N_18549,N_18229,N_18315);
nor U18550 (N_18550,N_18328,N_18335);
nand U18551 (N_18551,N_18338,N_18389);
xnor U18552 (N_18552,N_18289,N_18385);
xnor U18553 (N_18553,N_18298,N_18205);
xnor U18554 (N_18554,N_18370,N_18206);
and U18555 (N_18555,N_18379,N_18337);
nand U18556 (N_18556,N_18268,N_18345);
or U18557 (N_18557,N_18229,N_18249);
xor U18558 (N_18558,N_18294,N_18323);
xor U18559 (N_18559,N_18360,N_18218);
and U18560 (N_18560,N_18254,N_18252);
nor U18561 (N_18561,N_18226,N_18295);
nand U18562 (N_18562,N_18217,N_18397);
or U18563 (N_18563,N_18245,N_18399);
and U18564 (N_18564,N_18238,N_18213);
and U18565 (N_18565,N_18344,N_18374);
and U18566 (N_18566,N_18212,N_18357);
xnor U18567 (N_18567,N_18262,N_18341);
or U18568 (N_18568,N_18365,N_18344);
nand U18569 (N_18569,N_18319,N_18391);
xor U18570 (N_18570,N_18312,N_18376);
or U18571 (N_18571,N_18387,N_18207);
or U18572 (N_18572,N_18281,N_18333);
and U18573 (N_18573,N_18217,N_18290);
or U18574 (N_18574,N_18210,N_18354);
and U18575 (N_18575,N_18286,N_18299);
or U18576 (N_18576,N_18311,N_18364);
or U18577 (N_18577,N_18385,N_18250);
and U18578 (N_18578,N_18291,N_18261);
nor U18579 (N_18579,N_18321,N_18319);
or U18580 (N_18580,N_18202,N_18366);
nor U18581 (N_18581,N_18249,N_18342);
xor U18582 (N_18582,N_18359,N_18333);
and U18583 (N_18583,N_18266,N_18299);
or U18584 (N_18584,N_18284,N_18220);
or U18585 (N_18585,N_18222,N_18378);
nand U18586 (N_18586,N_18350,N_18362);
xor U18587 (N_18587,N_18362,N_18388);
nand U18588 (N_18588,N_18299,N_18304);
nor U18589 (N_18589,N_18322,N_18384);
nand U18590 (N_18590,N_18262,N_18301);
xnor U18591 (N_18591,N_18394,N_18378);
and U18592 (N_18592,N_18379,N_18382);
and U18593 (N_18593,N_18204,N_18368);
and U18594 (N_18594,N_18303,N_18289);
and U18595 (N_18595,N_18256,N_18318);
and U18596 (N_18596,N_18268,N_18368);
nor U18597 (N_18597,N_18294,N_18208);
xnor U18598 (N_18598,N_18278,N_18256);
nand U18599 (N_18599,N_18231,N_18311);
nand U18600 (N_18600,N_18532,N_18465);
nor U18601 (N_18601,N_18536,N_18455);
and U18602 (N_18602,N_18487,N_18450);
nor U18603 (N_18603,N_18580,N_18560);
nand U18604 (N_18604,N_18498,N_18473);
nor U18605 (N_18605,N_18556,N_18583);
xor U18606 (N_18606,N_18521,N_18578);
or U18607 (N_18607,N_18407,N_18575);
nor U18608 (N_18608,N_18571,N_18488);
and U18609 (N_18609,N_18515,N_18494);
or U18610 (N_18610,N_18479,N_18592);
nor U18611 (N_18611,N_18441,N_18484);
and U18612 (N_18612,N_18555,N_18459);
nand U18613 (N_18613,N_18404,N_18509);
nor U18614 (N_18614,N_18570,N_18584);
nand U18615 (N_18615,N_18490,N_18420);
and U18616 (N_18616,N_18561,N_18546);
xnor U18617 (N_18617,N_18475,N_18444);
nor U18618 (N_18618,N_18427,N_18503);
or U18619 (N_18619,N_18492,N_18564);
and U18620 (N_18620,N_18424,N_18426);
and U18621 (N_18621,N_18537,N_18405);
and U18622 (N_18622,N_18510,N_18458);
and U18623 (N_18623,N_18400,N_18542);
and U18624 (N_18624,N_18548,N_18429);
nand U18625 (N_18625,N_18595,N_18508);
and U18626 (N_18626,N_18485,N_18563);
nand U18627 (N_18627,N_18558,N_18468);
and U18628 (N_18628,N_18413,N_18440);
nand U18629 (N_18629,N_18573,N_18464);
nor U18630 (N_18630,N_18599,N_18401);
nand U18631 (N_18631,N_18545,N_18425);
or U18632 (N_18632,N_18528,N_18474);
or U18633 (N_18633,N_18552,N_18448);
xor U18634 (N_18634,N_18520,N_18486);
or U18635 (N_18635,N_18419,N_18534);
xor U18636 (N_18636,N_18456,N_18471);
or U18637 (N_18637,N_18519,N_18453);
xnor U18638 (N_18638,N_18550,N_18551);
and U18639 (N_18639,N_18457,N_18451);
xnor U18640 (N_18640,N_18476,N_18431);
xnor U18641 (N_18641,N_18432,N_18443);
xor U18642 (N_18642,N_18483,N_18449);
or U18643 (N_18643,N_18496,N_18547);
nor U18644 (N_18644,N_18574,N_18461);
and U18645 (N_18645,N_18495,N_18412);
xnor U18646 (N_18646,N_18576,N_18559);
or U18647 (N_18647,N_18582,N_18502);
nand U18648 (N_18648,N_18409,N_18469);
or U18649 (N_18649,N_18415,N_18524);
or U18650 (N_18650,N_18535,N_18539);
and U18651 (N_18651,N_18470,N_18463);
or U18652 (N_18652,N_18522,N_18439);
xnor U18653 (N_18653,N_18410,N_18506);
xnor U18654 (N_18654,N_18543,N_18562);
nor U18655 (N_18655,N_18554,N_18531);
nand U18656 (N_18656,N_18477,N_18418);
nand U18657 (N_18657,N_18587,N_18594);
nor U18658 (N_18658,N_18435,N_18452);
and U18659 (N_18659,N_18541,N_18565);
nand U18660 (N_18660,N_18406,N_18538);
or U18661 (N_18661,N_18598,N_18466);
nor U18662 (N_18662,N_18423,N_18527);
nor U18663 (N_18663,N_18530,N_18499);
nand U18664 (N_18664,N_18544,N_18549);
nand U18665 (N_18665,N_18446,N_18577);
or U18666 (N_18666,N_18586,N_18460);
nand U18667 (N_18667,N_18447,N_18417);
and U18668 (N_18668,N_18416,N_18568);
and U18669 (N_18669,N_18529,N_18408);
or U18670 (N_18670,N_18403,N_18438);
and U18671 (N_18671,N_18481,N_18590);
and U18672 (N_18672,N_18585,N_18581);
nor U18673 (N_18673,N_18589,N_18422);
and U18674 (N_18674,N_18540,N_18430);
xor U18675 (N_18675,N_18478,N_18591);
xnor U18676 (N_18676,N_18414,N_18507);
and U18677 (N_18677,N_18493,N_18436);
xor U18678 (N_18678,N_18480,N_18593);
nor U18679 (N_18679,N_18514,N_18454);
or U18680 (N_18680,N_18513,N_18505);
and U18681 (N_18681,N_18445,N_18421);
and U18682 (N_18682,N_18482,N_18462);
and U18683 (N_18683,N_18566,N_18579);
nand U18684 (N_18684,N_18489,N_18511);
nand U18685 (N_18685,N_18569,N_18434);
nor U18686 (N_18686,N_18533,N_18572);
nor U18687 (N_18687,N_18472,N_18501);
xor U18688 (N_18688,N_18567,N_18437);
nand U18689 (N_18689,N_18491,N_18504);
nor U18690 (N_18690,N_18411,N_18516);
nand U18691 (N_18691,N_18557,N_18512);
nand U18692 (N_18692,N_18526,N_18553);
nor U18693 (N_18693,N_18402,N_18497);
or U18694 (N_18694,N_18588,N_18596);
xnor U18695 (N_18695,N_18428,N_18523);
or U18696 (N_18696,N_18433,N_18525);
nor U18697 (N_18697,N_18597,N_18518);
nand U18698 (N_18698,N_18442,N_18517);
nor U18699 (N_18699,N_18467,N_18500);
xnor U18700 (N_18700,N_18599,N_18530);
nor U18701 (N_18701,N_18445,N_18497);
xnor U18702 (N_18702,N_18529,N_18541);
and U18703 (N_18703,N_18595,N_18478);
and U18704 (N_18704,N_18495,N_18421);
xnor U18705 (N_18705,N_18478,N_18427);
nor U18706 (N_18706,N_18462,N_18499);
xnor U18707 (N_18707,N_18576,N_18423);
or U18708 (N_18708,N_18433,N_18582);
nand U18709 (N_18709,N_18563,N_18452);
and U18710 (N_18710,N_18497,N_18433);
or U18711 (N_18711,N_18595,N_18424);
or U18712 (N_18712,N_18580,N_18521);
nor U18713 (N_18713,N_18467,N_18436);
xnor U18714 (N_18714,N_18403,N_18569);
and U18715 (N_18715,N_18452,N_18475);
or U18716 (N_18716,N_18510,N_18525);
xnor U18717 (N_18717,N_18573,N_18528);
nor U18718 (N_18718,N_18492,N_18508);
xor U18719 (N_18719,N_18561,N_18573);
and U18720 (N_18720,N_18443,N_18458);
and U18721 (N_18721,N_18567,N_18445);
nand U18722 (N_18722,N_18417,N_18522);
nor U18723 (N_18723,N_18466,N_18405);
nor U18724 (N_18724,N_18543,N_18530);
xor U18725 (N_18725,N_18542,N_18503);
nor U18726 (N_18726,N_18494,N_18525);
or U18727 (N_18727,N_18493,N_18530);
nand U18728 (N_18728,N_18474,N_18580);
or U18729 (N_18729,N_18590,N_18575);
xor U18730 (N_18730,N_18560,N_18563);
xnor U18731 (N_18731,N_18501,N_18424);
xnor U18732 (N_18732,N_18525,N_18537);
and U18733 (N_18733,N_18465,N_18427);
and U18734 (N_18734,N_18549,N_18517);
xor U18735 (N_18735,N_18410,N_18420);
nor U18736 (N_18736,N_18457,N_18534);
nor U18737 (N_18737,N_18485,N_18553);
xnor U18738 (N_18738,N_18495,N_18443);
and U18739 (N_18739,N_18497,N_18581);
or U18740 (N_18740,N_18400,N_18471);
and U18741 (N_18741,N_18465,N_18591);
xor U18742 (N_18742,N_18496,N_18433);
nor U18743 (N_18743,N_18532,N_18440);
nand U18744 (N_18744,N_18494,N_18457);
xnor U18745 (N_18745,N_18431,N_18459);
nor U18746 (N_18746,N_18444,N_18546);
nand U18747 (N_18747,N_18499,N_18505);
or U18748 (N_18748,N_18515,N_18418);
nor U18749 (N_18749,N_18517,N_18449);
nor U18750 (N_18750,N_18438,N_18510);
nand U18751 (N_18751,N_18567,N_18554);
nor U18752 (N_18752,N_18508,N_18537);
nor U18753 (N_18753,N_18439,N_18575);
and U18754 (N_18754,N_18496,N_18573);
nor U18755 (N_18755,N_18508,N_18573);
or U18756 (N_18756,N_18584,N_18479);
xor U18757 (N_18757,N_18431,N_18552);
xnor U18758 (N_18758,N_18450,N_18496);
nor U18759 (N_18759,N_18557,N_18561);
nand U18760 (N_18760,N_18508,N_18591);
and U18761 (N_18761,N_18576,N_18527);
or U18762 (N_18762,N_18450,N_18416);
nand U18763 (N_18763,N_18465,N_18579);
nor U18764 (N_18764,N_18458,N_18439);
nand U18765 (N_18765,N_18572,N_18595);
nor U18766 (N_18766,N_18536,N_18598);
and U18767 (N_18767,N_18583,N_18555);
nor U18768 (N_18768,N_18573,N_18557);
nand U18769 (N_18769,N_18544,N_18418);
and U18770 (N_18770,N_18438,N_18461);
and U18771 (N_18771,N_18457,N_18415);
xor U18772 (N_18772,N_18438,N_18559);
and U18773 (N_18773,N_18405,N_18401);
nor U18774 (N_18774,N_18478,N_18535);
or U18775 (N_18775,N_18411,N_18475);
xor U18776 (N_18776,N_18421,N_18480);
xnor U18777 (N_18777,N_18403,N_18471);
or U18778 (N_18778,N_18530,N_18526);
and U18779 (N_18779,N_18521,N_18447);
nand U18780 (N_18780,N_18479,N_18493);
nand U18781 (N_18781,N_18597,N_18450);
or U18782 (N_18782,N_18482,N_18437);
nand U18783 (N_18783,N_18553,N_18415);
nand U18784 (N_18784,N_18591,N_18436);
or U18785 (N_18785,N_18520,N_18407);
xnor U18786 (N_18786,N_18596,N_18558);
xor U18787 (N_18787,N_18560,N_18548);
and U18788 (N_18788,N_18587,N_18582);
nor U18789 (N_18789,N_18413,N_18554);
nor U18790 (N_18790,N_18569,N_18429);
xor U18791 (N_18791,N_18478,N_18521);
or U18792 (N_18792,N_18458,N_18499);
or U18793 (N_18793,N_18416,N_18535);
nand U18794 (N_18794,N_18417,N_18454);
or U18795 (N_18795,N_18564,N_18447);
nand U18796 (N_18796,N_18448,N_18598);
nor U18797 (N_18797,N_18494,N_18568);
xnor U18798 (N_18798,N_18466,N_18522);
xnor U18799 (N_18799,N_18459,N_18484);
nor U18800 (N_18800,N_18620,N_18706);
nand U18801 (N_18801,N_18756,N_18629);
nor U18802 (N_18802,N_18681,N_18766);
nand U18803 (N_18803,N_18742,N_18670);
or U18804 (N_18804,N_18789,N_18744);
or U18805 (N_18805,N_18733,N_18637);
nor U18806 (N_18806,N_18775,N_18728);
or U18807 (N_18807,N_18652,N_18639);
xor U18808 (N_18808,N_18763,N_18748);
and U18809 (N_18809,N_18799,N_18631);
or U18810 (N_18810,N_18772,N_18619);
or U18811 (N_18811,N_18625,N_18716);
or U18812 (N_18812,N_18678,N_18732);
nor U18813 (N_18813,N_18630,N_18721);
and U18814 (N_18814,N_18665,N_18700);
xor U18815 (N_18815,N_18718,N_18692);
and U18816 (N_18816,N_18623,N_18759);
nand U18817 (N_18817,N_18729,N_18693);
and U18818 (N_18818,N_18632,N_18653);
nor U18819 (N_18819,N_18740,N_18642);
xor U18820 (N_18820,N_18663,N_18634);
nor U18821 (N_18821,N_18750,N_18749);
nor U18822 (N_18822,N_18719,N_18798);
or U18823 (N_18823,N_18672,N_18776);
xnor U18824 (N_18824,N_18784,N_18753);
nor U18825 (N_18825,N_18709,N_18644);
nor U18826 (N_18826,N_18701,N_18682);
or U18827 (N_18827,N_18671,N_18697);
or U18828 (N_18828,N_18752,N_18680);
and U18829 (N_18829,N_18794,N_18786);
or U18830 (N_18830,N_18788,N_18616);
xor U18831 (N_18831,N_18796,N_18604);
xnor U18832 (N_18832,N_18731,N_18726);
and U18833 (N_18833,N_18797,N_18661);
and U18834 (N_18834,N_18610,N_18702);
or U18835 (N_18835,N_18765,N_18628);
xnor U18836 (N_18836,N_18677,N_18707);
or U18837 (N_18837,N_18648,N_18601);
xor U18838 (N_18838,N_18687,N_18626);
xor U18839 (N_18839,N_18602,N_18674);
and U18840 (N_18840,N_18715,N_18764);
nor U18841 (N_18841,N_18689,N_18724);
nor U18842 (N_18842,N_18656,N_18771);
xor U18843 (N_18843,N_18641,N_18699);
and U18844 (N_18844,N_18624,N_18679);
and U18845 (N_18845,N_18683,N_18668);
nor U18846 (N_18846,N_18758,N_18767);
nand U18847 (N_18847,N_18605,N_18774);
nand U18848 (N_18848,N_18795,N_18600);
or U18849 (N_18849,N_18710,N_18770);
xor U18850 (N_18850,N_18761,N_18757);
nor U18851 (N_18851,N_18647,N_18618);
nor U18852 (N_18852,N_18611,N_18614);
nand U18853 (N_18853,N_18633,N_18655);
nand U18854 (N_18854,N_18650,N_18603);
or U18855 (N_18855,N_18747,N_18708);
and U18856 (N_18856,N_18792,N_18727);
xor U18857 (N_18857,N_18608,N_18755);
nor U18858 (N_18858,N_18651,N_18645);
or U18859 (N_18859,N_18660,N_18609);
or U18860 (N_18860,N_18695,N_18754);
or U18861 (N_18861,N_18649,N_18606);
or U18862 (N_18862,N_18621,N_18778);
nor U18863 (N_18863,N_18694,N_18745);
and U18864 (N_18864,N_18617,N_18790);
nor U18865 (N_18865,N_18658,N_18643);
nand U18866 (N_18866,N_18720,N_18723);
or U18867 (N_18867,N_18612,N_18714);
nand U18868 (N_18868,N_18646,N_18704);
nand U18869 (N_18869,N_18607,N_18730);
xnor U18870 (N_18870,N_18640,N_18684);
or U18871 (N_18871,N_18780,N_18782);
nor U18872 (N_18872,N_18713,N_18739);
nand U18873 (N_18873,N_18711,N_18717);
nand U18874 (N_18874,N_18736,N_18703);
nand U18875 (N_18875,N_18690,N_18638);
nor U18876 (N_18876,N_18738,N_18627);
nor U18877 (N_18877,N_18666,N_18698);
xnor U18878 (N_18878,N_18615,N_18667);
nand U18879 (N_18879,N_18777,N_18793);
and U18880 (N_18880,N_18676,N_18760);
and U18881 (N_18881,N_18779,N_18635);
or U18882 (N_18882,N_18769,N_18696);
nand U18883 (N_18883,N_18662,N_18734);
and U18884 (N_18884,N_18791,N_18785);
nand U18885 (N_18885,N_18705,N_18613);
nand U18886 (N_18886,N_18712,N_18691);
xnor U18887 (N_18887,N_18659,N_18741);
and U18888 (N_18888,N_18737,N_18746);
or U18889 (N_18889,N_18673,N_18685);
nor U18890 (N_18890,N_18751,N_18743);
nor U18891 (N_18891,N_18622,N_18787);
nor U18892 (N_18892,N_18686,N_18735);
or U18893 (N_18893,N_18669,N_18688);
nand U18894 (N_18894,N_18675,N_18722);
nor U18895 (N_18895,N_18657,N_18762);
nand U18896 (N_18896,N_18636,N_18773);
xor U18897 (N_18897,N_18664,N_18781);
and U18898 (N_18898,N_18768,N_18783);
nand U18899 (N_18899,N_18725,N_18654);
nand U18900 (N_18900,N_18610,N_18798);
or U18901 (N_18901,N_18678,N_18720);
and U18902 (N_18902,N_18644,N_18733);
and U18903 (N_18903,N_18714,N_18674);
and U18904 (N_18904,N_18681,N_18731);
and U18905 (N_18905,N_18636,N_18759);
nor U18906 (N_18906,N_18663,N_18792);
or U18907 (N_18907,N_18797,N_18722);
xnor U18908 (N_18908,N_18631,N_18725);
nor U18909 (N_18909,N_18613,N_18676);
and U18910 (N_18910,N_18602,N_18722);
nor U18911 (N_18911,N_18698,N_18615);
xor U18912 (N_18912,N_18781,N_18793);
nand U18913 (N_18913,N_18748,N_18770);
or U18914 (N_18914,N_18758,N_18717);
xor U18915 (N_18915,N_18755,N_18679);
xor U18916 (N_18916,N_18756,N_18769);
and U18917 (N_18917,N_18683,N_18747);
nand U18918 (N_18918,N_18761,N_18644);
nor U18919 (N_18919,N_18661,N_18722);
xnor U18920 (N_18920,N_18727,N_18612);
xor U18921 (N_18921,N_18622,N_18618);
or U18922 (N_18922,N_18720,N_18793);
nand U18923 (N_18923,N_18701,N_18669);
and U18924 (N_18924,N_18727,N_18796);
or U18925 (N_18925,N_18635,N_18718);
nand U18926 (N_18926,N_18635,N_18772);
and U18927 (N_18927,N_18688,N_18619);
xnor U18928 (N_18928,N_18706,N_18618);
nor U18929 (N_18929,N_18660,N_18792);
and U18930 (N_18930,N_18659,N_18720);
nand U18931 (N_18931,N_18728,N_18620);
and U18932 (N_18932,N_18625,N_18641);
xnor U18933 (N_18933,N_18678,N_18776);
nand U18934 (N_18934,N_18666,N_18697);
or U18935 (N_18935,N_18678,N_18689);
xor U18936 (N_18936,N_18648,N_18615);
nand U18937 (N_18937,N_18608,N_18603);
nor U18938 (N_18938,N_18603,N_18782);
nor U18939 (N_18939,N_18673,N_18793);
nor U18940 (N_18940,N_18792,N_18606);
nand U18941 (N_18941,N_18719,N_18634);
nor U18942 (N_18942,N_18757,N_18737);
or U18943 (N_18943,N_18636,N_18675);
xnor U18944 (N_18944,N_18761,N_18612);
or U18945 (N_18945,N_18667,N_18748);
or U18946 (N_18946,N_18797,N_18672);
and U18947 (N_18947,N_18799,N_18719);
or U18948 (N_18948,N_18744,N_18609);
nor U18949 (N_18949,N_18777,N_18772);
nor U18950 (N_18950,N_18666,N_18623);
and U18951 (N_18951,N_18774,N_18722);
nand U18952 (N_18952,N_18724,N_18783);
nor U18953 (N_18953,N_18681,N_18775);
nand U18954 (N_18954,N_18642,N_18731);
nor U18955 (N_18955,N_18659,N_18689);
xnor U18956 (N_18956,N_18735,N_18768);
nand U18957 (N_18957,N_18693,N_18761);
or U18958 (N_18958,N_18685,N_18776);
nand U18959 (N_18959,N_18629,N_18767);
nand U18960 (N_18960,N_18603,N_18725);
or U18961 (N_18961,N_18692,N_18688);
nor U18962 (N_18962,N_18710,N_18666);
or U18963 (N_18963,N_18789,N_18684);
and U18964 (N_18964,N_18609,N_18623);
or U18965 (N_18965,N_18790,N_18697);
xor U18966 (N_18966,N_18679,N_18719);
xor U18967 (N_18967,N_18667,N_18774);
nor U18968 (N_18968,N_18615,N_18773);
or U18969 (N_18969,N_18701,N_18717);
and U18970 (N_18970,N_18659,N_18691);
xnor U18971 (N_18971,N_18788,N_18659);
nor U18972 (N_18972,N_18735,N_18676);
xor U18973 (N_18973,N_18779,N_18638);
nor U18974 (N_18974,N_18777,N_18791);
xnor U18975 (N_18975,N_18647,N_18637);
xnor U18976 (N_18976,N_18658,N_18668);
nor U18977 (N_18977,N_18716,N_18715);
xnor U18978 (N_18978,N_18658,N_18788);
and U18979 (N_18979,N_18645,N_18690);
xor U18980 (N_18980,N_18639,N_18666);
nand U18981 (N_18981,N_18723,N_18656);
nand U18982 (N_18982,N_18759,N_18757);
and U18983 (N_18983,N_18738,N_18750);
xnor U18984 (N_18984,N_18673,N_18763);
or U18985 (N_18985,N_18680,N_18725);
xor U18986 (N_18986,N_18703,N_18601);
or U18987 (N_18987,N_18721,N_18626);
and U18988 (N_18988,N_18652,N_18625);
nand U18989 (N_18989,N_18720,N_18608);
or U18990 (N_18990,N_18758,N_18748);
or U18991 (N_18991,N_18673,N_18708);
nand U18992 (N_18992,N_18636,N_18742);
xnor U18993 (N_18993,N_18660,N_18683);
and U18994 (N_18994,N_18654,N_18626);
and U18995 (N_18995,N_18631,N_18661);
nand U18996 (N_18996,N_18780,N_18655);
and U18997 (N_18997,N_18754,N_18788);
or U18998 (N_18998,N_18658,N_18671);
xor U18999 (N_18999,N_18680,N_18632);
and U19000 (N_19000,N_18918,N_18962);
or U19001 (N_19001,N_18826,N_18899);
xnor U19002 (N_19002,N_18831,N_18970);
xnor U19003 (N_19003,N_18820,N_18924);
nand U19004 (N_19004,N_18840,N_18828);
or U19005 (N_19005,N_18864,N_18830);
or U19006 (N_19006,N_18916,N_18837);
or U19007 (N_19007,N_18921,N_18809);
nor U19008 (N_19008,N_18926,N_18838);
or U19009 (N_19009,N_18975,N_18994);
nand U19010 (N_19010,N_18834,N_18875);
and U19011 (N_19011,N_18813,N_18836);
and U19012 (N_19012,N_18900,N_18925);
and U19013 (N_19013,N_18877,N_18889);
or U19014 (N_19014,N_18964,N_18846);
nand U19015 (N_19015,N_18818,N_18980);
or U19016 (N_19016,N_18917,N_18863);
xor U19017 (N_19017,N_18893,N_18909);
nor U19018 (N_19018,N_18829,N_18835);
nand U19019 (N_19019,N_18937,N_18876);
nand U19020 (N_19020,N_18800,N_18951);
nor U19021 (N_19021,N_18895,N_18867);
and U19022 (N_19022,N_18928,N_18896);
and U19023 (N_19023,N_18844,N_18849);
nor U19024 (N_19024,N_18966,N_18959);
nand U19025 (N_19025,N_18821,N_18885);
or U19026 (N_19026,N_18982,N_18969);
or U19027 (N_19027,N_18903,N_18940);
nand U19028 (N_19028,N_18906,N_18850);
xnor U19029 (N_19029,N_18802,N_18901);
or U19030 (N_19030,N_18967,N_18948);
nor U19031 (N_19031,N_18833,N_18804);
and U19032 (N_19032,N_18985,N_18858);
nand U19033 (N_19033,N_18816,N_18920);
xor U19034 (N_19034,N_18987,N_18891);
nand U19035 (N_19035,N_18855,N_18988);
nand U19036 (N_19036,N_18897,N_18806);
nor U19037 (N_19037,N_18949,N_18823);
xor U19038 (N_19038,N_18845,N_18848);
and U19039 (N_19039,N_18968,N_18851);
nand U19040 (N_19040,N_18839,N_18868);
and U19041 (N_19041,N_18908,N_18973);
nand U19042 (N_19042,N_18805,N_18871);
xnor U19043 (N_19043,N_18887,N_18983);
nand U19044 (N_19044,N_18999,N_18825);
or U19045 (N_19045,N_18808,N_18857);
nor U19046 (N_19046,N_18963,N_18955);
nor U19047 (N_19047,N_18919,N_18971);
and U19048 (N_19048,N_18856,N_18934);
nand U19049 (N_19049,N_18807,N_18933);
xor U19050 (N_19050,N_18824,N_18907);
nor U19051 (N_19051,N_18812,N_18881);
nor U19052 (N_19052,N_18990,N_18938);
nand U19053 (N_19053,N_18932,N_18873);
nor U19054 (N_19054,N_18946,N_18931);
xor U19055 (N_19055,N_18860,N_18911);
nor U19056 (N_19056,N_18870,N_18953);
nor U19057 (N_19057,N_18892,N_18817);
nand U19058 (N_19058,N_18993,N_18954);
nand U19059 (N_19059,N_18942,N_18810);
nor U19060 (N_19060,N_18989,N_18922);
nor U19061 (N_19061,N_18945,N_18883);
and U19062 (N_19062,N_18986,N_18972);
and U19063 (N_19063,N_18944,N_18902);
nor U19064 (N_19064,N_18827,N_18803);
nand U19065 (N_19065,N_18936,N_18952);
or U19066 (N_19066,N_18865,N_18923);
or U19067 (N_19067,N_18974,N_18976);
or U19068 (N_19068,N_18941,N_18815);
and U19069 (N_19069,N_18978,N_18874);
and U19070 (N_19070,N_18957,N_18910);
or U19071 (N_19071,N_18819,N_18898);
xor U19072 (N_19072,N_18882,N_18822);
or U19073 (N_19073,N_18984,N_18886);
or U19074 (N_19074,N_18996,N_18960);
xor U19075 (N_19075,N_18811,N_18977);
nand U19076 (N_19076,N_18878,N_18981);
nor U19077 (N_19077,N_18843,N_18888);
nor U19078 (N_19078,N_18814,N_18995);
xor U19079 (N_19079,N_18914,N_18947);
nor U19080 (N_19080,N_18929,N_18862);
and U19081 (N_19081,N_18879,N_18847);
xor U19082 (N_19082,N_18861,N_18853);
xnor U19083 (N_19083,N_18997,N_18866);
and U19084 (N_19084,N_18842,N_18852);
nand U19085 (N_19085,N_18958,N_18992);
and U19086 (N_19086,N_18859,N_18979);
or U19087 (N_19087,N_18872,N_18894);
nor U19088 (N_19088,N_18998,N_18927);
nor U19089 (N_19089,N_18890,N_18965);
xnor U19090 (N_19090,N_18950,N_18880);
or U19091 (N_19091,N_18832,N_18869);
nor U19092 (N_19092,N_18912,N_18961);
or U19093 (N_19093,N_18884,N_18905);
xnor U19094 (N_19094,N_18930,N_18939);
nand U19095 (N_19095,N_18943,N_18841);
nor U19096 (N_19096,N_18991,N_18913);
or U19097 (N_19097,N_18915,N_18904);
or U19098 (N_19098,N_18956,N_18854);
xnor U19099 (N_19099,N_18801,N_18935);
and U19100 (N_19100,N_18958,N_18969);
nand U19101 (N_19101,N_18983,N_18895);
xor U19102 (N_19102,N_18825,N_18986);
nor U19103 (N_19103,N_18855,N_18974);
and U19104 (N_19104,N_18802,N_18958);
or U19105 (N_19105,N_18884,N_18958);
xnor U19106 (N_19106,N_18942,N_18835);
nor U19107 (N_19107,N_18867,N_18818);
nand U19108 (N_19108,N_18989,N_18869);
xnor U19109 (N_19109,N_18993,N_18951);
or U19110 (N_19110,N_18894,N_18828);
nand U19111 (N_19111,N_18920,N_18923);
nor U19112 (N_19112,N_18954,N_18872);
xnor U19113 (N_19113,N_18844,N_18887);
or U19114 (N_19114,N_18954,N_18886);
and U19115 (N_19115,N_18933,N_18945);
and U19116 (N_19116,N_18904,N_18967);
or U19117 (N_19117,N_18812,N_18897);
xnor U19118 (N_19118,N_18963,N_18832);
or U19119 (N_19119,N_18991,N_18868);
nand U19120 (N_19120,N_18893,N_18950);
xnor U19121 (N_19121,N_18849,N_18840);
nand U19122 (N_19122,N_18957,N_18987);
and U19123 (N_19123,N_18825,N_18802);
xor U19124 (N_19124,N_18819,N_18800);
nor U19125 (N_19125,N_18923,N_18949);
nand U19126 (N_19126,N_18883,N_18822);
nor U19127 (N_19127,N_18802,N_18883);
xor U19128 (N_19128,N_18914,N_18879);
nor U19129 (N_19129,N_18861,N_18832);
xor U19130 (N_19130,N_18919,N_18994);
or U19131 (N_19131,N_18822,N_18867);
nor U19132 (N_19132,N_18913,N_18877);
or U19133 (N_19133,N_18842,N_18995);
nor U19134 (N_19134,N_18801,N_18844);
xnor U19135 (N_19135,N_18970,N_18886);
and U19136 (N_19136,N_18808,N_18973);
and U19137 (N_19137,N_18864,N_18978);
xnor U19138 (N_19138,N_18910,N_18812);
nand U19139 (N_19139,N_18943,N_18869);
xnor U19140 (N_19140,N_18883,N_18914);
nor U19141 (N_19141,N_18998,N_18885);
xnor U19142 (N_19142,N_18855,N_18922);
nand U19143 (N_19143,N_18834,N_18830);
nor U19144 (N_19144,N_18863,N_18933);
xnor U19145 (N_19145,N_18963,N_18867);
nand U19146 (N_19146,N_18887,N_18829);
xnor U19147 (N_19147,N_18837,N_18961);
or U19148 (N_19148,N_18926,N_18903);
and U19149 (N_19149,N_18854,N_18874);
xor U19150 (N_19150,N_18812,N_18992);
xor U19151 (N_19151,N_18818,N_18804);
and U19152 (N_19152,N_18883,N_18999);
or U19153 (N_19153,N_18801,N_18818);
xor U19154 (N_19154,N_18840,N_18833);
nor U19155 (N_19155,N_18857,N_18981);
and U19156 (N_19156,N_18803,N_18819);
nand U19157 (N_19157,N_18906,N_18968);
nand U19158 (N_19158,N_18919,N_18839);
xnor U19159 (N_19159,N_18921,N_18980);
or U19160 (N_19160,N_18814,N_18921);
nand U19161 (N_19161,N_18856,N_18939);
and U19162 (N_19162,N_18823,N_18922);
and U19163 (N_19163,N_18956,N_18988);
xnor U19164 (N_19164,N_18845,N_18898);
and U19165 (N_19165,N_18905,N_18882);
xor U19166 (N_19166,N_18830,N_18943);
and U19167 (N_19167,N_18852,N_18860);
or U19168 (N_19168,N_18868,N_18983);
or U19169 (N_19169,N_18879,N_18918);
and U19170 (N_19170,N_18926,N_18825);
xor U19171 (N_19171,N_18838,N_18924);
nor U19172 (N_19172,N_18902,N_18903);
nor U19173 (N_19173,N_18984,N_18924);
nand U19174 (N_19174,N_18828,N_18851);
nand U19175 (N_19175,N_18975,N_18992);
and U19176 (N_19176,N_18977,N_18850);
nand U19177 (N_19177,N_18835,N_18871);
xor U19178 (N_19178,N_18813,N_18943);
or U19179 (N_19179,N_18840,N_18855);
nor U19180 (N_19180,N_18835,N_18830);
or U19181 (N_19181,N_18818,N_18906);
xnor U19182 (N_19182,N_18841,N_18993);
xor U19183 (N_19183,N_18859,N_18923);
and U19184 (N_19184,N_18819,N_18804);
nor U19185 (N_19185,N_18858,N_18902);
xor U19186 (N_19186,N_18917,N_18975);
or U19187 (N_19187,N_18970,N_18875);
xor U19188 (N_19188,N_18849,N_18918);
xor U19189 (N_19189,N_18907,N_18818);
nand U19190 (N_19190,N_18974,N_18895);
xor U19191 (N_19191,N_18984,N_18832);
nor U19192 (N_19192,N_18979,N_18987);
xor U19193 (N_19193,N_18821,N_18815);
or U19194 (N_19194,N_18850,N_18925);
nor U19195 (N_19195,N_18940,N_18966);
or U19196 (N_19196,N_18927,N_18849);
or U19197 (N_19197,N_18868,N_18865);
and U19198 (N_19198,N_18821,N_18860);
xnor U19199 (N_19199,N_18978,N_18912);
and U19200 (N_19200,N_19142,N_19169);
and U19201 (N_19201,N_19011,N_19131);
nor U19202 (N_19202,N_19067,N_19019);
or U19203 (N_19203,N_19178,N_19090);
and U19204 (N_19204,N_19110,N_19192);
and U19205 (N_19205,N_19031,N_19144);
nor U19206 (N_19206,N_19030,N_19016);
nand U19207 (N_19207,N_19156,N_19088);
nand U19208 (N_19208,N_19127,N_19133);
and U19209 (N_19209,N_19009,N_19124);
nor U19210 (N_19210,N_19107,N_19176);
and U19211 (N_19211,N_19140,N_19010);
nor U19212 (N_19212,N_19159,N_19155);
nand U19213 (N_19213,N_19021,N_19000);
nor U19214 (N_19214,N_19027,N_19051);
nor U19215 (N_19215,N_19005,N_19062);
and U19216 (N_19216,N_19029,N_19123);
xor U19217 (N_19217,N_19091,N_19056);
or U19218 (N_19218,N_19138,N_19174);
or U19219 (N_19219,N_19053,N_19173);
and U19220 (N_19220,N_19170,N_19194);
nand U19221 (N_19221,N_19046,N_19137);
or U19222 (N_19222,N_19099,N_19177);
or U19223 (N_19223,N_19070,N_19101);
nor U19224 (N_19224,N_19003,N_19085);
nor U19225 (N_19225,N_19007,N_19164);
and U19226 (N_19226,N_19072,N_19092);
nor U19227 (N_19227,N_19055,N_19041);
and U19228 (N_19228,N_19082,N_19077);
xor U19229 (N_19229,N_19081,N_19083);
xnor U19230 (N_19230,N_19069,N_19023);
or U19231 (N_19231,N_19047,N_19108);
nor U19232 (N_19232,N_19198,N_19154);
and U19233 (N_19233,N_19167,N_19017);
and U19234 (N_19234,N_19105,N_19151);
nor U19235 (N_19235,N_19097,N_19008);
nor U19236 (N_19236,N_19139,N_19116);
and U19237 (N_19237,N_19036,N_19112);
xor U19238 (N_19238,N_19106,N_19148);
xor U19239 (N_19239,N_19004,N_19013);
or U19240 (N_19240,N_19060,N_19136);
or U19241 (N_19241,N_19033,N_19002);
or U19242 (N_19242,N_19145,N_19117);
xnor U19243 (N_19243,N_19180,N_19100);
xnor U19244 (N_19244,N_19073,N_19181);
nor U19245 (N_19245,N_19102,N_19187);
or U19246 (N_19246,N_19061,N_19163);
xnor U19247 (N_19247,N_19063,N_19183);
nand U19248 (N_19248,N_19093,N_19121);
nand U19249 (N_19249,N_19084,N_19040);
xnor U19250 (N_19250,N_19015,N_19038);
xnor U19251 (N_19251,N_19050,N_19188);
nand U19252 (N_19252,N_19166,N_19146);
xnor U19253 (N_19253,N_19126,N_19157);
nor U19254 (N_19254,N_19199,N_19043);
or U19255 (N_19255,N_19095,N_19078);
xnor U19256 (N_19256,N_19074,N_19162);
or U19257 (N_19257,N_19119,N_19025);
xor U19258 (N_19258,N_19052,N_19037);
nor U19259 (N_19259,N_19066,N_19186);
or U19260 (N_19260,N_19065,N_19197);
nor U19261 (N_19261,N_19161,N_19068);
nand U19262 (N_19262,N_19184,N_19193);
and U19263 (N_19263,N_19118,N_19039);
nor U19264 (N_19264,N_19014,N_19087);
and U19265 (N_19265,N_19071,N_19185);
xnor U19266 (N_19266,N_19122,N_19135);
xnor U19267 (N_19267,N_19001,N_19160);
or U19268 (N_19268,N_19153,N_19058);
nor U19269 (N_19269,N_19094,N_19191);
xor U19270 (N_19270,N_19149,N_19165);
xor U19271 (N_19271,N_19132,N_19028);
nand U19272 (N_19272,N_19048,N_19018);
xnor U19273 (N_19273,N_19086,N_19006);
and U19274 (N_19274,N_19098,N_19172);
xor U19275 (N_19275,N_19045,N_19075);
xnor U19276 (N_19276,N_19035,N_19147);
and U19277 (N_19277,N_19196,N_19026);
xnor U19278 (N_19278,N_19080,N_19032);
or U19279 (N_19279,N_19054,N_19109);
or U19280 (N_19280,N_19089,N_19022);
nor U19281 (N_19281,N_19076,N_19143);
xor U19282 (N_19282,N_19152,N_19115);
nor U19283 (N_19283,N_19057,N_19130);
nor U19284 (N_19284,N_19044,N_19096);
or U19285 (N_19285,N_19120,N_19141);
nand U19286 (N_19286,N_19079,N_19103);
nand U19287 (N_19287,N_19175,N_19171);
xnor U19288 (N_19288,N_19129,N_19195);
or U19289 (N_19289,N_19104,N_19012);
nand U19290 (N_19290,N_19158,N_19134);
nor U19291 (N_19291,N_19125,N_19168);
or U19292 (N_19292,N_19059,N_19182);
and U19293 (N_19293,N_19064,N_19150);
xor U19294 (N_19294,N_19189,N_19049);
nand U19295 (N_19295,N_19179,N_19042);
and U19296 (N_19296,N_19020,N_19128);
and U19297 (N_19297,N_19190,N_19114);
nand U19298 (N_19298,N_19113,N_19111);
nor U19299 (N_19299,N_19024,N_19034);
nand U19300 (N_19300,N_19087,N_19111);
nand U19301 (N_19301,N_19102,N_19103);
xor U19302 (N_19302,N_19134,N_19087);
or U19303 (N_19303,N_19051,N_19068);
or U19304 (N_19304,N_19046,N_19106);
and U19305 (N_19305,N_19099,N_19123);
nor U19306 (N_19306,N_19118,N_19136);
nand U19307 (N_19307,N_19016,N_19027);
nor U19308 (N_19308,N_19062,N_19132);
and U19309 (N_19309,N_19099,N_19129);
and U19310 (N_19310,N_19135,N_19184);
xnor U19311 (N_19311,N_19114,N_19128);
nand U19312 (N_19312,N_19133,N_19176);
nand U19313 (N_19313,N_19116,N_19064);
and U19314 (N_19314,N_19096,N_19071);
or U19315 (N_19315,N_19022,N_19162);
xnor U19316 (N_19316,N_19097,N_19179);
nor U19317 (N_19317,N_19013,N_19020);
xor U19318 (N_19318,N_19175,N_19152);
or U19319 (N_19319,N_19067,N_19042);
nor U19320 (N_19320,N_19091,N_19018);
nand U19321 (N_19321,N_19022,N_19115);
or U19322 (N_19322,N_19080,N_19060);
nand U19323 (N_19323,N_19016,N_19048);
xor U19324 (N_19324,N_19001,N_19070);
or U19325 (N_19325,N_19010,N_19184);
or U19326 (N_19326,N_19020,N_19179);
nor U19327 (N_19327,N_19174,N_19184);
nand U19328 (N_19328,N_19193,N_19148);
and U19329 (N_19329,N_19052,N_19131);
and U19330 (N_19330,N_19004,N_19064);
nor U19331 (N_19331,N_19193,N_19043);
nand U19332 (N_19332,N_19151,N_19047);
or U19333 (N_19333,N_19086,N_19185);
xnor U19334 (N_19334,N_19137,N_19041);
and U19335 (N_19335,N_19027,N_19162);
xor U19336 (N_19336,N_19191,N_19058);
xor U19337 (N_19337,N_19192,N_19026);
xnor U19338 (N_19338,N_19146,N_19112);
nand U19339 (N_19339,N_19193,N_19172);
xnor U19340 (N_19340,N_19023,N_19177);
xnor U19341 (N_19341,N_19134,N_19093);
and U19342 (N_19342,N_19174,N_19178);
nor U19343 (N_19343,N_19101,N_19005);
and U19344 (N_19344,N_19162,N_19106);
or U19345 (N_19345,N_19032,N_19170);
nor U19346 (N_19346,N_19150,N_19152);
xnor U19347 (N_19347,N_19028,N_19164);
nand U19348 (N_19348,N_19121,N_19178);
nand U19349 (N_19349,N_19140,N_19143);
nor U19350 (N_19350,N_19124,N_19090);
and U19351 (N_19351,N_19015,N_19094);
nor U19352 (N_19352,N_19106,N_19103);
or U19353 (N_19353,N_19095,N_19032);
xnor U19354 (N_19354,N_19048,N_19160);
or U19355 (N_19355,N_19156,N_19084);
or U19356 (N_19356,N_19051,N_19120);
nand U19357 (N_19357,N_19102,N_19154);
or U19358 (N_19358,N_19048,N_19011);
xor U19359 (N_19359,N_19098,N_19043);
nor U19360 (N_19360,N_19011,N_19197);
and U19361 (N_19361,N_19037,N_19133);
and U19362 (N_19362,N_19198,N_19029);
nor U19363 (N_19363,N_19172,N_19062);
or U19364 (N_19364,N_19082,N_19027);
xor U19365 (N_19365,N_19090,N_19126);
xor U19366 (N_19366,N_19088,N_19075);
or U19367 (N_19367,N_19069,N_19047);
nor U19368 (N_19368,N_19158,N_19110);
xor U19369 (N_19369,N_19034,N_19158);
nand U19370 (N_19370,N_19074,N_19147);
or U19371 (N_19371,N_19140,N_19085);
nor U19372 (N_19372,N_19182,N_19169);
and U19373 (N_19373,N_19053,N_19132);
and U19374 (N_19374,N_19127,N_19001);
and U19375 (N_19375,N_19047,N_19139);
xnor U19376 (N_19376,N_19178,N_19069);
xnor U19377 (N_19377,N_19128,N_19105);
and U19378 (N_19378,N_19167,N_19139);
or U19379 (N_19379,N_19168,N_19035);
and U19380 (N_19380,N_19083,N_19017);
or U19381 (N_19381,N_19088,N_19079);
and U19382 (N_19382,N_19010,N_19104);
xnor U19383 (N_19383,N_19058,N_19183);
xor U19384 (N_19384,N_19050,N_19020);
or U19385 (N_19385,N_19180,N_19116);
nand U19386 (N_19386,N_19194,N_19162);
nor U19387 (N_19387,N_19104,N_19063);
nor U19388 (N_19388,N_19054,N_19131);
and U19389 (N_19389,N_19161,N_19092);
nand U19390 (N_19390,N_19010,N_19156);
xor U19391 (N_19391,N_19151,N_19027);
and U19392 (N_19392,N_19197,N_19099);
nor U19393 (N_19393,N_19134,N_19031);
xnor U19394 (N_19394,N_19157,N_19129);
or U19395 (N_19395,N_19102,N_19172);
xnor U19396 (N_19396,N_19153,N_19156);
nor U19397 (N_19397,N_19176,N_19028);
nor U19398 (N_19398,N_19169,N_19112);
xor U19399 (N_19399,N_19089,N_19038);
xor U19400 (N_19400,N_19204,N_19211);
and U19401 (N_19401,N_19203,N_19240);
and U19402 (N_19402,N_19263,N_19361);
or U19403 (N_19403,N_19383,N_19270);
or U19404 (N_19404,N_19286,N_19382);
and U19405 (N_19405,N_19314,N_19300);
and U19406 (N_19406,N_19368,N_19336);
nand U19407 (N_19407,N_19302,N_19224);
nor U19408 (N_19408,N_19290,N_19365);
nand U19409 (N_19409,N_19212,N_19233);
nand U19410 (N_19410,N_19305,N_19310);
nor U19411 (N_19411,N_19251,N_19202);
and U19412 (N_19412,N_19316,N_19200);
xor U19413 (N_19413,N_19265,N_19234);
and U19414 (N_19414,N_19249,N_19289);
nor U19415 (N_19415,N_19298,N_19238);
or U19416 (N_19416,N_19268,N_19397);
xor U19417 (N_19417,N_19210,N_19285);
and U19418 (N_19418,N_19362,N_19245);
and U19419 (N_19419,N_19244,N_19342);
or U19420 (N_19420,N_19225,N_19374);
xnor U19421 (N_19421,N_19283,N_19367);
and U19422 (N_19422,N_19372,N_19333);
and U19423 (N_19423,N_19259,N_19223);
or U19424 (N_19424,N_19272,N_19311);
or U19425 (N_19425,N_19339,N_19214);
xor U19426 (N_19426,N_19381,N_19299);
xnor U19427 (N_19427,N_19222,N_19359);
xor U19428 (N_19428,N_19366,N_19201);
nand U19429 (N_19429,N_19221,N_19261);
or U19430 (N_19430,N_19293,N_19355);
nand U19431 (N_19431,N_19232,N_19328);
nand U19432 (N_19432,N_19294,N_19350);
or U19433 (N_19433,N_19349,N_19247);
and U19434 (N_19434,N_19320,N_19392);
nor U19435 (N_19435,N_19207,N_19390);
or U19436 (N_19436,N_19326,N_19334);
or U19437 (N_19437,N_19216,N_19356);
xor U19438 (N_19438,N_19346,N_19318);
nor U19439 (N_19439,N_19380,N_19242);
xnor U19440 (N_19440,N_19394,N_19275);
nor U19441 (N_19441,N_19288,N_19387);
and U19442 (N_19442,N_19280,N_19279);
xnor U19443 (N_19443,N_19271,N_19277);
nand U19444 (N_19444,N_19291,N_19398);
nor U19445 (N_19445,N_19317,N_19378);
nand U19446 (N_19446,N_19255,N_19227);
xnor U19447 (N_19447,N_19246,N_19254);
nand U19448 (N_19448,N_19231,N_19396);
nand U19449 (N_19449,N_19315,N_19287);
xnor U19450 (N_19450,N_19331,N_19354);
nor U19451 (N_19451,N_19284,N_19330);
xnor U19452 (N_19452,N_19295,N_19309);
nand U19453 (N_19453,N_19377,N_19278);
nor U19454 (N_19454,N_19257,N_19395);
or U19455 (N_19455,N_19357,N_19217);
and U19456 (N_19456,N_19208,N_19229);
or U19457 (N_19457,N_19352,N_19370);
and U19458 (N_19458,N_19371,N_19343);
and U19459 (N_19459,N_19306,N_19351);
and U19460 (N_19460,N_19205,N_19296);
xnor U19461 (N_19461,N_19226,N_19239);
nand U19462 (N_19462,N_19281,N_19258);
nor U19463 (N_19463,N_19376,N_19267);
and U19464 (N_19464,N_19269,N_19319);
nand U19465 (N_19465,N_19358,N_19250);
nor U19466 (N_19466,N_19332,N_19369);
and U19467 (N_19467,N_19219,N_19388);
nand U19468 (N_19468,N_19338,N_19327);
and U19469 (N_19469,N_19364,N_19312);
nand U19470 (N_19470,N_19385,N_19230);
nor U19471 (N_19471,N_19206,N_19266);
nand U19472 (N_19472,N_19304,N_19235);
and U19473 (N_19473,N_19292,N_19253);
xor U19474 (N_19474,N_19347,N_19297);
or U19475 (N_19475,N_19301,N_19373);
nor U19476 (N_19476,N_19220,N_19276);
nor U19477 (N_19477,N_19345,N_19323);
xnor U19478 (N_19478,N_19264,N_19308);
or U19479 (N_19479,N_19391,N_19393);
and U19480 (N_19480,N_19307,N_19236);
xnor U19481 (N_19481,N_19324,N_19344);
nor U19482 (N_19482,N_19260,N_19335);
xnor U19483 (N_19483,N_19379,N_19340);
nand U19484 (N_19484,N_19274,N_19241);
xor U19485 (N_19485,N_19360,N_19389);
or U19486 (N_19486,N_19273,N_19282);
xnor U19487 (N_19487,N_19303,N_19262);
nor U19488 (N_19488,N_19237,N_19322);
nand U19489 (N_19489,N_19313,N_19348);
and U19490 (N_19490,N_19256,N_19386);
and U19491 (N_19491,N_19215,N_19228);
and U19492 (N_19492,N_19353,N_19213);
nor U19493 (N_19493,N_19321,N_19399);
or U19494 (N_19494,N_19248,N_19252);
and U19495 (N_19495,N_19341,N_19243);
nand U19496 (N_19496,N_19384,N_19325);
or U19497 (N_19497,N_19329,N_19218);
and U19498 (N_19498,N_19209,N_19375);
and U19499 (N_19499,N_19363,N_19337);
and U19500 (N_19500,N_19285,N_19248);
or U19501 (N_19501,N_19341,N_19372);
and U19502 (N_19502,N_19255,N_19283);
xor U19503 (N_19503,N_19254,N_19298);
nand U19504 (N_19504,N_19358,N_19333);
xnor U19505 (N_19505,N_19374,N_19357);
nor U19506 (N_19506,N_19223,N_19390);
nor U19507 (N_19507,N_19211,N_19309);
nand U19508 (N_19508,N_19312,N_19248);
nand U19509 (N_19509,N_19312,N_19352);
or U19510 (N_19510,N_19354,N_19294);
nor U19511 (N_19511,N_19362,N_19318);
and U19512 (N_19512,N_19216,N_19318);
or U19513 (N_19513,N_19211,N_19205);
nand U19514 (N_19514,N_19384,N_19276);
or U19515 (N_19515,N_19342,N_19309);
nand U19516 (N_19516,N_19318,N_19251);
or U19517 (N_19517,N_19338,N_19387);
or U19518 (N_19518,N_19223,N_19237);
nor U19519 (N_19519,N_19353,N_19204);
nand U19520 (N_19520,N_19394,N_19313);
or U19521 (N_19521,N_19328,N_19285);
xnor U19522 (N_19522,N_19386,N_19313);
xnor U19523 (N_19523,N_19394,N_19207);
or U19524 (N_19524,N_19237,N_19219);
xnor U19525 (N_19525,N_19306,N_19255);
xor U19526 (N_19526,N_19392,N_19217);
nand U19527 (N_19527,N_19245,N_19240);
nand U19528 (N_19528,N_19272,N_19391);
nand U19529 (N_19529,N_19343,N_19288);
nand U19530 (N_19530,N_19348,N_19289);
or U19531 (N_19531,N_19281,N_19218);
nor U19532 (N_19532,N_19303,N_19235);
or U19533 (N_19533,N_19253,N_19290);
or U19534 (N_19534,N_19380,N_19259);
nor U19535 (N_19535,N_19319,N_19234);
or U19536 (N_19536,N_19228,N_19257);
nand U19537 (N_19537,N_19294,N_19262);
nand U19538 (N_19538,N_19296,N_19367);
xor U19539 (N_19539,N_19211,N_19346);
nand U19540 (N_19540,N_19299,N_19271);
xor U19541 (N_19541,N_19231,N_19328);
nor U19542 (N_19542,N_19275,N_19240);
and U19543 (N_19543,N_19391,N_19242);
nand U19544 (N_19544,N_19372,N_19273);
xor U19545 (N_19545,N_19211,N_19303);
nor U19546 (N_19546,N_19304,N_19282);
or U19547 (N_19547,N_19315,N_19239);
nor U19548 (N_19548,N_19322,N_19369);
and U19549 (N_19549,N_19254,N_19204);
nand U19550 (N_19550,N_19363,N_19364);
xnor U19551 (N_19551,N_19384,N_19355);
xnor U19552 (N_19552,N_19347,N_19373);
nand U19553 (N_19553,N_19278,N_19214);
or U19554 (N_19554,N_19262,N_19285);
nand U19555 (N_19555,N_19224,N_19223);
nand U19556 (N_19556,N_19319,N_19289);
nor U19557 (N_19557,N_19238,N_19372);
xnor U19558 (N_19558,N_19230,N_19249);
or U19559 (N_19559,N_19303,N_19362);
nand U19560 (N_19560,N_19220,N_19380);
and U19561 (N_19561,N_19328,N_19333);
nand U19562 (N_19562,N_19389,N_19245);
or U19563 (N_19563,N_19283,N_19299);
or U19564 (N_19564,N_19209,N_19232);
nor U19565 (N_19565,N_19377,N_19201);
nand U19566 (N_19566,N_19267,N_19365);
xor U19567 (N_19567,N_19203,N_19370);
nor U19568 (N_19568,N_19227,N_19315);
and U19569 (N_19569,N_19232,N_19224);
or U19570 (N_19570,N_19297,N_19304);
and U19571 (N_19571,N_19204,N_19221);
nand U19572 (N_19572,N_19352,N_19349);
nand U19573 (N_19573,N_19343,N_19299);
nor U19574 (N_19574,N_19214,N_19275);
nand U19575 (N_19575,N_19264,N_19285);
nor U19576 (N_19576,N_19258,N_19221);
or U19577 (N_19577,N_19335,N_19272);
xnor U19578 (N_19578,N_19259,N_19340);
xnor U19579 (N_19579,N_19220,N_19350);
or U19580 (N_19580,N_19263,N_19271);
xor U19581 (N_19581,N_19289,N_19363);
nand U19582 (N_19582,N_19306,N_19363);
xnor U19583 (N_19583,N_19365,N_19368);
xor U19584 (N_19584,N_19395,N_19255);
and U19585 (N_19585,N_19282,N_19229);
nor U19586 (N_19586,N_19302,N_19269);
and U19587 (N_19587,N_19344,N_19261);
or U19588 (N_19588,N_19232,N_19230);
and U19589 (N_19589,N_19378,N_19235);
nor U19590 (N_19590,N_19297,N_19355);
nor U19591 (N_19591,N_19377,N_19256);
or U19592 (N_19592,N_19283,N_19372);
or U19593 (N_19593,N_19292,N_19269);
and U19594 (N_19594,N_19251,N_19209);
xnor U19595 (N_19595,N_19230,N_19321);
and U19596 (N_19596,N_19303,N_19285);
and U19597 (N_19597,N_19261,N_19234);
nand U19598 (N_19598,N_19322,N_19307);
or U19599 (N_19599,N_19300,N_19264);
nor U19600 (N_19600,N_19501,N_19410);
nand U19601 (N_19601,N_19563,N_19581);
and U19602 (N_19602,N_19437,N_19522);
and U19603 (N_19603,N_19424,N_19451);
and U19604 (N_19604,N_19405,N_19431);
xnor U19605 (N_19605,N_19535,N_19530);
xnor U19606 (N_19606,N_19597,N_19561);
nor U19607 (N_19607,N_19492,N_19416);
nand U19608 (N_19608,N_19589,N_19433);
and U19609 (N_19609,N_19529,N_19441);
nand U19610 (N_19610,N_19464,N_19432);
nor U19611 (N_19611,N_19578,N_19542);
nand U19612 (N_19612,N_19452,N_19466);
xor U19613 (N_19613,N_19521,N_19468);
nand U19614 (N_19614,N_19478,N_19460);
and U19615 (N_19615,N_19459,N_19557);
xor U19616 (N_19616,N_19423,N_19536);
or U19617 (N_19617,N_19496,N_19584);
xor U19618 (N_19618,N_19485,N_19534);
nand U19619 (N_19619,N_19400,N_19434);
nor U19620 (N_19620,N_19549,N_19541);
or U19621 (N_19621,N_19412,N_19588);
xnor U19622 (N_19622,N_19594,N_19533);
nand U19623 (N_19623,N_19489,N_19463);
nand U19624 (N_19624,N_19573,N_19403);
and U19625 (N_19625,N_19420,N_19560);
nor U19626 (N_19626,N_19553,N_19414);
nand U19627 (N_19627,N_19550,N_19546);
and U19628 (N_19628,N_19487,N_19500);
nand U19629 (N_19629,N_19547,N_19457);
nor U19630 (N_19630,N_19506,N_19590);
nand U19631 (N_19631,N_19537,N_19462);
nor U19632 (N_19632,N_19504,N_19592);
nand U19633 (N_19633,N_19455,N_19598);
xor U19634 (N_19634,N_19568,N_19525);
and U19635 (N_19635,N_19407,N_19572);
or U19636 (N_19636,N_19596,N_19418);
xor U19637 (N_19637,N_19456,N_19454);
or U19638 (N_19638,N_19479,N_19559);
xor U19639 (N_19639,N_19507,N_19404);
or U19640 (N_19640,N_19531,N_19488);
nand U19641 (N_19641,N_19471,N_19562);
nor U19642 (N_19642,N_19427,N_19422);
nand U19643 (N_19643,N_19470,N_19587);
xnor U19644 (N_19644,N_19439,N_19540);
xnor U19645 (N_19645,N_19556,N_19510);
nor U19646 (N_19646,N_19580,N_19551);
nand U19647 (N_19647,N_19490,N_19574);
or U19648 (N_19648,N_19526,N_19583);
and U19649 (N_19649,N_19402,N_19519);
and U19650 (N_19650,N_19435,N_19532);
or U19651 (N_19651,N_19520,N_19458);
nand U19652 (N_19652,N_19419,N_19509);
and U19653 (N_19653,N_19577,N_19512);
nor U19654 (N_19654,N_19453,N_19545);
xor U19655 (N_19655,N_19593,N_19480);
nor U19656 (N_19656,N_19595,N_19428);
or U19657 (N_19657,N_19515,N_19538);
or U19658 (N_19658,N_19513,N_19543);
xnor U19659 (N_19659,N_19415,N_19497);
or U19660 (N_19660,N_19436,N_19444);
nand U19661 (N_19661,N_19586,N_19544);
nand U19662 (N_19662,N_19565,N_19467);
xnor U19663 (N_19663,N_19469,N_19539);
nor U19664 (N_19664,N_19576,N_19445);
and U19665 (N_19665,N_19503,N_19575);
and U19666 (N_19666,N_19484,N_19417);
nand U19667 (N_19667,N_19477,N_19406);
xnor U19668 (N_19668,N_19566,N_19448);
xor U19669 (N_19669,N_19425,N_19493);
xnor U19670 (N_19670,N_19481,N_19571);
xnor U19671 (N_19671,N_19591,N_19440);
and U19672 (N_19672,N_19518,N_19461);
nor U19673 (N_19673,N_19567,N_19472);
xnor U19674 (N_19674,N_19554,N_19450);
and U19675 (N_19675,N_19528,N_19411);
nor U19676 (N_19676,N_19430,N_19482);
or U19677 (N_19677,N_19514,N_19483);
nand U19678 (N_19678,N_19570,N_19409);
or U19679 (N_19679,N_19508,N_19429);
nor U19680 (N_19680,N_19495,N_19446);
or U19681 (N_19681,N_19498,N_19473);
nor U19682 (N_19682,N_19408,N_19491);
xnor U19683 (N_19683,N_19527,N_19401);
nor U19684 (N_19684,N_19585,N_19569);
nand U19685 (N_19685,N_19599,N_19516);
nor U19686 (N_19686,N_19486,N_19421);
xnor U19687 (N_19687,N_19548,N_19499);
nor U19688 (N_19688,N_19474,N_19494);
or U19689 (N_19689,N_19465,N_19426);
nand U19690 (N_19690,N_19502,N_19449);
and U19691 (N_19691,N_19443,N_19582);
nand U19692 (N_19692,N_19476,N_19523);
nor U19693 (N_19693,N_19413,N_19558);
xor U19694 (N_19694,N_19524,N_19475);
or U19695 (N_19695,N_19442,N_19552);
nor U19696 (N_19696,N_19438,N_19511);
xnor U19697 (N_19697,N_19517,N_19447);
nor U19698 (N_19698,N_19579,N_19564);
and U19699 (N_19699,N_19505,N_19555);
xor U19700 (N_19700,N_19550,N_19593);
or U19701 (N_19701,N_19504,N_19452);
nand U19702 (N_19702,N_19443,N_19505);
or U19703 (N_19703,N_19592,N_19497);
or U19704 (N_19704,N_19563,N_19504);
nor U19705 (N_19705,N_19593,N_19545);
nand U19706 (N_19706,N_19409,N_19487);
nand U19707 (N_19707,N_19432,N_19512);
nand U19708 (N_19708,N_19455,N_19424);
nand U19709 (N_19709,N_19540,N_19436);
nand U19710 (N_19710,N_19561,N_19586);
xnor U19711 (N_19711,N_19555,N_19401);
nand U19712 (N_19712,N_19501,N_19548);
xor U19713 (N_19713,N_19421,N_19579);
nand U19714 (N_19714,N_19588,N_19467);
xnor U19715 (N_19715,N_19507,N_19580);
nand U19716 (N_19716,N_19461,N_19494);
xor U19717 (N_19717,N_19418,N_19536);
and U19718 (N_19718,N_19512,N_19513);
and U19719 (N_19719,N_19541,N_19520);
nor U19720 (N_19720,N_19525,N_19567);
nor U19721 (N_19721,N_19578,N_19591);
xor U19722 (N_19722,N_19482,N_19592);
nand U19723 (N_19723,N_19588,N_19423);
and U19724 (N_19724,N_19546,N_19589);
and U19725 (N_19725,N_19419,N_19530);
and U19726 (N_19726,N_19445,N_19446);
nand U19727 (N_19727,N_19404,N_19437);
xor U19728 (N_19728,N_19464,N_19496);
or U19729 (N_19729,N_19460,N_19471);
nand U19730 (N_19730,N_19437,N_19502);
nor U19731 (N_19731,N_19495,N_19438);
nor U19732 (N_19732,N_19513,N_19487);
nor U19733 (N_19733,N_19513,N_19599);
xnor U19734 (N_19734,N_19531,N_19409);
nor U19735 (N_19735,N_19436,N_19448);
nand U19736 (N_19736,N_19450,N_19465);
nand U19737 (N_19737,N_19586,N_19438);
nand U19738 (N_19738,N_19488,N_19482);
nand U19739 (N_19739,N_19460,N_19465);
and U19740 (N_19740,N_19556,N_19438);
xor U19741 (N_19741,N_19419,N_19475);
or U19742 (N_19742,N_19401,N_19547);
nand U19743 (N_19743,N_19471,N_19439);
and U19744 (N_19744,N_19590,N_19479);
xnor U19745 (N_19745,N_19483,N_19557);
xnor U19746 (N_19746,N_19465,N_19405);
nor U19747 (N_19747,N_19547,N_19407);
nand U19748 (N_19748,N_19451,N_19503);
nand U19749 (N_19749,N_19568,N_19598);
nand U19750 (N_19750,N_19482,N_19469);
or U19751 (N_19751,N_19485,N_19566);
and U19752 (N_19752,N_19537,N_19436);
nand U19753 (N_19753,N_19408,N_19492);
xnor U19754 (N_19754,N_19433,N_19492);
nor U19755 (N_19755,N_19550,N_19507);
nand U19756 (N_19756,N_19517,N_19481);
nand U19757 (N_19757,N_19589,N_19540);
nand U19758 (N_19758,N_19426,N_19406);
and U19759 (N_19759,N_19407,N_19525);
nand U19760 (N_19760,N_19541,N_19448);
and U19761 (N_19761,N_19453,N_19419);
nand U19762 (N_19762,N_19536,N_19538);
and U19763 (N_19763,N_19584,N_19510);
and U19764 (N_19764,N_19472,N_19466);
xnor U19765 (N_19765,N_19474,N_19463);
xnor U19766 (N_19766,N_19569,N_19491);
or U19767 (N_19767,N_19576,N_19522);
nor U19768 (N_19768,N_19523,N_19590);
nand U19769 (N_19769,N_19418,N_19403);
nor U19770 (N_19770,N_19517,N_19585);
xnor U19771 (N_19771,N_19577,N_19448);
or U19772 (N_19772,N_19501,N_19568);
and U19773 (N_19773,N_19414,N_19547);
or U19774 (N_19774,N_19581,N_19565);
nor U19775 (N_19775,N_19403,N_19509);
nand U19776 (N_19776,N_19564,N_19449);
nand U19777 (N_19777,N_19415,N_19512);
or U19778 (N_19778,N_19461,N_19414);
and U19779 (N_19779,N_19459,N_19507);
xnor U19780 (N_19780,N_19482,N_19569);
and U19781 (N_19781,N_19403,N_19463);
nand U19782 (N_19782,N_19469,N_19546);
nand U19783 (N_19783,N_19484,N_19522);
or U19784 (N_19784,N_19504,N_19502);
or U19785 (N_19785,N_19415,N_19407);
xor U19786 (N_19786,N_19567,N_19436);
and U19787 (N_19787,N_19413,N_19421);
or U19788 (N_19788,N_19532,N_19403);
and U19789 (N_19789,N_19597,N_19516);
and U19790 (N_19790,N_19499,N_19567);
and U19791 (N_19791,N_19553,N_19555);
nor U19792 (N_19792,N_19496,N_19478);
or U19793 (N_19793,N_19509,N_19544);
and U19794 (N_19794,N_19445,N_19487);
nor U19795 (N_19795,N_19530,N_19526);
or U19796 (N_19796,N_19528,N_19471);
nand U19797 (N_19797,N_19489,N_19470);
nand U19798 (N_19798,N_19522,N_19552);
nor U19799 (N_19799,N_19410,N_19562);
nor U19800 (N_19800,N_19788,N_19775);
or U19801 (N_19801,N_19774,N_19603);
and U19802 (N_19802,N_19798,N_19673);
nand U19803 (N_19803,N_19662,N_19653);
xor U19804 (N_19804,N_19770,N_19696);
xnor U19805 (N_19805,N_19666,N_19638);
xnor U19806 (N_19806,N_19635,N_19694);
xnor U19807 (N_19807,N_19762,N_19741);
nor U19808 (N_19808,N_19738,N_19615);
or U19809 (N_19809,N_19742,N_19684);
and U19810 (N_19810,N_19688,N_19637);
nand U19811 (N_19811,N_19701,N_19730);
nor U19812 (N_19812,N_19699,N_19636);
nor U19813 (N_19813,N_19685,N_19627);
and U19814 (N_19814,N_19654,N_19720);
and U19815 (N_19815,N_19715,N_19795);
and U19816 (N_19816,N_19749,N_19690);
and U19817 (N_19817,N_19668,N_19671);
and U19818 (N_19818,N_19644,N_19607);
nand U19819 (N_19819,N_19723,N_19725);
xor U19820 (N_19820,N_19791,N_19672);
nor U19821 (N_19821,N_19773,N_19618);
nor U19822 (N_19822,N_19729,N_19796);
nand U19823 (N_19823,N_19634,N_19670);
and U19824 (N_19824,N_19744,N_19799);
or U19825 (N_19825,N_19783,N_19691);
xor U19826 (N_19826,N_19789,N_19784);
nand U19827 (N_19827,N_19661,N_19600);
nor U19828 (N_19828,N_19659,N_19612);
and U19829 (N_19829,N_19757,N_19655);
nor U19830 (N_19830,N_19793,N_19679);
and U19831 (N_19831,N_19755,N_19753);
and U19832 (N_19832,N_19728,N_19610);
nand U19833 (N_19833,N_19777,N_19769);
nand U19834 (N_19834,N_19628,N_19633);
nand U19835 (N_19835,N_19790,N_19669);
and U19836 (N_19836,N_19613,N_19781);
nand U19837 (N_19837,N_19665,N_19608);
or U19838 (N_19838,N_19686,N_19767);
xor U19839 (N_19839,N_19745,N_19719);
nand U19840 (N_19840,N_19619,N_19640);
nand U19841 (N_19841,N_19601,N_19766);
nand U19842 (N_19842,N_19717,N_19706);
nor U19843 (N_19843,N_19626,N_19731);
and U19844 (N_19844,N_19697,N_19629);
or U19845 (N_19845,N_19776,N_19754);
nor U19846 (N_19846,N_19782,N_19643);
nand U19847 (N_19847,N_19726,N_19732);
and U19848 (N_19848,N_19602,N_19703);
or U19849 (N_19849,N_19786,N_19737);
nor U19850 (N_19850,N_19747,N_19649);
nor U19851 (N_19851,N_19680,N_19624);
nor U19852 (N_19852,N_19702,N_19724);
or U19853 (N_19853,N_19639,N_19660);
nor U19854 (N_19854,N_19740,N_19713);
or U19855 (N_19855,N_19716,N_19631);
xnor U19856 (N_19856,N_19718,N_19704);
or U19857 (N_19857,N_19761,N_19616);
or U19858 (N_19858,N_19681,N_19642);
or U19859 (N_19859,N_19736,N_19692);
and U19860 (N_19860,N_19710,N_19748);
xor U19861 (N_19861,N_19751,N_19605);
and U19862 (N_19862,N_19746,N_19657);
or U19863 (N_19863,N_19698,N_19641);
nor U19864 (N_19864,N_19768,N_19604);
or U19865 (N_19865,N_19650,N_19722);
xor U19866 (N_19866,N_19647,N_19648);
nand U19867 (N_19867,N_19772,N_19658);
or U19868 (N_19868,N_19667,N_19617);
and U19869 (N_19869,N_19780,N_19709);
nor U19870 (N_19870,N_19727,N_19609);
and U19871 (N_19871,N_19763,N_19651);
and U19872 (N_19872,N_19797,N_19632);
and U19873 (N_19873,N_19625,N_19721);
xnor U19874 (N_19874,N_19792,N_19700);
nor U19875 (N_19875,N_19611,N_19733);
nor U19876 (N_19876,N_19794,N_19752);
xnor U19877 (N_19877,N_19674,N_19645);
nand U19878 (N_19878,N_19785,N_19620);
xor U19879 (N_19879,N_19764,N_19708);
nand U19880 (N_19880,N_19663,N_19676);
nand U19881 (N_19881,N_19622,N_19623);
nand U19882 (N_19882,N_19652,N_19656);
xnor U19883 (N_19883,N_19787,N_19778);
nand U19884 (N_19884,N_19739,N_19750);
nor U19885 (N_19885,N_19758,N_19707);
and U19886 (N_19886,N_19760,N_19743);
xor U19887 (N_19887,N_19614,N_19664);
nor U19888 (N_19888,N_19606,N_19759);
xnor U19889 (N_19889,N_19621,N_19682);
and U19890 (N_19890,N_19693,N_19756);
or U19891 (N_19891,N_19689,N_19675);
nand U19892 (N_19892,N_19646,N_19630);
nand U19893 (N_19893,N_19712,N_19734);
and U19894 (N_19894,N_19695,N_19677);
nand U19895 (N_19895,N_19683,N_19714);
or U19896 (N_19896,N_19678,N_19687);
xnor U19897 (N_19897,N_19771,N_19779);
or U19898 (N_19898,N_19765,N_19705);
and U19899 (N_19899,N_19711,N_19735);
xor U19900 (N_19900,N_19798,N_19739);
nand U19901 (N_19901,N_19620,N_19789);
nand U19902 (N_19902,N_19712,N_19776);
xor U19903 (N_19903,N_19716,N_19673);
and U19904 (N_19904,N_19612,N_19754);
xnor U19905 (N_19905,N_19668,N_19665);
nor U19906 (N_19906,N_19659,N_19720);
and U19907 (N_19907,N_19788,N_19639);
nor U19908 (N_19908,N_19783,N_19727);
and U19909 (N_19909,N_19754,N_19668);
nand U19910 (N_19910,N_19648,N_19714);
and U19911 (N_19911,N_19797,N_19716);
nor U19912 (N_19912,N_19655,N_19762);
or U19913 (N_19913,N_19711,N_19687);
xnor U19914 (N_19914,N_19604,N_19763);
xnor U19915 (N_19915,N_19645,N_19730);
and U19916 (N_19916,N_19682,N_19648);
nor U19917 (N_19917,N_19674,N_19791);
nand U19918 (N_19918,N_19684,N_19672);
and U19919 (N_19919,N_19702,N_19752);
and U19920 (N_19920,N_19796,N_19765);
xnor U19921 (N_19921,N_19705,N_19619);
or U19922 (N_19922,N_19772,N_19799);
and U19923 (N_19923,N_19727,N_19638);
nand U19924 (N_19924,N_19780,N_19783);
or U19925 (N_19925,N_19603,N_19736);
nor U19926 (N_19926,N_19718,N_19741);
and U19927 (N_19927,N_19700,N_19737);
nor U19928 (N_19928,N_19790,N_19711);
nor U19929 (N_19929,N_19717,N_19699);
nor U19930 (N_19930,N_19655,N_19776);
nand U19931 (N_19931,N_19697,N_19718);
xnor U19932 (N_19932,N_19787,N_19731);
nand U19933 (N_19933,N_19780,N_19620);
nand U19934 (N_19934,N_19632,N_19750);
and U19935 (N_19935,N_19729,N_19777);
xor U19936 (N_19936,N_19750,N_19778);
xor U19937 (N_19937,N_19602,N_19603);
nor U19938 (N_19938,N_19627,N_19790);
and U19939 (N_19939,N_19618,N_19686);
and U19940 (N_19940,N_19776,N_19783);
or U19941 (N_19941,N_19688,N_19719);
xnor U19942 (N_19942,N_19740,N_19698);
xnor U19943 (N_19943,N_19690,N_19778);
nand U19944 (N_19944,N_19646,N_19753);
nand U19945 (N_19945,N_19757,N_19666);
nor U19946 (N_19946,N_19732,N_19681);
and U19947 (N_19947,N_19744,N_19650);
nand U19948 (N_19948,N_19631,N_19664);
or U19949 (N_19949,N_19722,N_19656);
nor U19950 (N_19950,N_19726,N_19793);
xor U19951 (N_19951,N_19695,N_19761);
xor U19952 (N_19952,N_19715,N_19718);
or U19953 (N_19953,N_19748,N_19671);
or U19954 (N_19954,N_19694,N_19604);
and U19955 (N_19955,N_19627,N_19681);
nand U19956 (N_19956,N_19771,N_19688);
xnor U19957 (N_19957,N_19619,N_19790);
and U19958 (N_19958,N_19799,N_19642);
nor U19959 (N_19959,N_19673,N_19672);
xnor U19960 (N_19960,N_19790,N_19743);
and U19961 (N_19961,N_19653,N_19788);
or U19962 (N_19962,N_19792,N_19631);
and U19963 (N_19963,N_19600,N_19677);
nand U19964 (N_19964,N_19685,N_19621);
xor U19965 (N_19965,N_19667,N_19753);
or U19966 (N_19966,N_19663,N_19604);
nand U19967 (N_19967,N_19711,N_19647);
nor U19968 (N_19968,N_19720,N_19679);
nor U19969 (N_19969,N_19660,N_19784);
nor U19970 (N_19970,N_19677,N_19616);
nand U19971 (N_19971,N_19703,N_19704);
nor U19972 (N_19972,N_19635,N_19716);
or U19973 (N_19973,N_19681,N_19760);
and U19974 (N_19974,N_19638,N_19716);
or U19975 (N_19975,N_19639,N_19726);
and U19976 (N_19976,N_19653,N_19601);
or U19977 (N_19977,N_19782,N_19685);
nand U19978 (N_19978,N_19670,N_19766);
nand U19979 (N_19979,N_19745,N_19724);
nand U19980 (N_19980,N_19661,N_19627);
or U19981 (N_19981,N_19707,N_19722);
nor U19982 (N_19982,N_19602,N_19704);
xor U19983 (N_19983,N_19755,N_19640);
xnor U19984 (N_19984,N_19637,N_19754);
and U19985 (N_19985,N_19664,N_19727);
nand U19986 (N_19986,N_19700,N_19663);
nand U19987 (N_19987,N_19779,N_19723);
or U19988 (N_19988,N_19652,N_19617);
or U19989 (N_19989,N_19610,N_19770);
nor U19990 (N_19990,N_19740,N_19633);
nand U19991 (N_19991,N_19622,N_19737);
xnor U19992 (N_19992,N_19618,N_19629);
xnor U19993 (N_19993,N_19746,N_19760);
xnor U19994 (N_19994,N_19721,N_19715);
nor U19995 (N_19995,N_19729,N_19601);
and U19996 (N_19996,N_19723,N_19604);
xor U19997 (N_19997,N_19622,N_19710);
xor U19998 (N_19998,N_19796,N_19735);
nand U19999 (N_19999,N_19625,N_19675);
nand U20000 (N_20000,N_19892,N_19839);
and U20001 (N_20001,N_19830,N_19961);
nor U20002 (N_20002,N_19947,N_19949);
and U20003 (N_20003,N_19976,N_19935);
and U20004 (N_20004,N_19818,N_19845);
or U20005 (N_20005,N_19822,N_19856);
nor U20006 (N_20006,N_19966,N_19952);
and U20007 (N_20007,N_19863,N_19859);
and U20008 (N_20008,N_19975,N_19938);
nor U20009 (N_20009,N_19804,N_19862);
and U20010 (N_20010,N_19898,N_19833);
nand U20011 (N_20011,N_19843,N_19867);
nor U20012 (N_20012,N_19944,N_19971);
nor U20013 (N_20013,N_19986,N_19891);
xnor U20014 (N_20014,N_19846,N_19992);
nor U20015 (N_20015,N_19801,N_19873);
nor U20016 (N_20016,N_19817,N_19924);
or U20017 (N_20017,N_19864,N_19942);
xnor U20018 (N_20018,N_19934,N_19920);
nand U20019 (N_20019,N_19894,N_19950);
or U20020 (N_20020,N_19906,N_19878);
and U20021 (N_20021,N_19980,N_19909);
and U20022 (N_20022,N_19943,N_19903);
xnor U20023 (N_20023,N_19884,N_19930);
or U20024 (N_20024,N_19993,N_19893);
nand U20025 (N_20025,N_19923,N_19956);
xor U20026 (N_20026,N_19872,N_19984);
nor U20027 (N_20027,N_19912,N_19805);
xor U20028 (N_20028,N_19854,N_19974);
nor U20029 (N_20029,N_19853,N_19803);
xnor U20030 (N_20030,N_19978,N_19815);
nand U20031 (N_20031,N_19861,N_19905);
xor U20032 (N_20032,N_19904,N_19835);
and U20033 (N_20033,N_19850,N_19800);
nand U20034 (N_20034,N_19998,N_19851);
xor U20035 (N_20035,N_19836,N_19962);
and U20036 (N_20036,N_19911,N_19847);
nor U20037 (N_20037,N_19996,N_19871);
nand U20038 (N_20038,N_19916,N_19838);
nand U20039 (N_20039,N_19951,N_19963);
xnor U20040 (N_20040,N_19931,N_19816);
or U20041 (N_20041,N_19883,N_19810);
or U20042 (N_20042,N_19831,N_19841);
nor U20043 (N_20043,N_19899,N_19985);
nor U20044 (N_20044,N_19896,N_19987);
xor U20045 (N_20045,N_19989,N_19882);
and U20046 (N_20046,N_19828,N_19954);
or U20047 (N_20047,N_19929,N_19844);
xor U20048 (N_20048,N_19933,N_19879);
nand U20049 (N_20049,N_19819,N_19994);
xnor U20050 (N_20050,N_19874,N_19983);
nand U20051 (N_20051,N_19932,N_19890);
xnor U20052 (N_20052,N_19928,N_19870);
nand U20053 (N_20053,N_19922,N_19955);
or U20054 (N_20054,N_19936,N_19813);
nand U20055 (N_20055,N_19868,N_19809);
or U20056 (N_20056,N_19915,N_19999);
or U20057 (N_20057,N_19900,N_19865);
or U20058 (N_20058,N_19965,N_19913);
nand U20059 (N_20059,N_19907,N_19866);
and U20060 (N_20060,N_19808,N_19967);
nor U20061 (N_20061,N_19902,N_19919);
or U20062 (N_20062,N_19941,N_19960);
or U20063 (N_20063,N_19885,N_19973);
xnor U20064 (N_20064,N_19880,N_19889);
nor U20065 (N_20065,N_19926,N_19888);
nor U20066 (N_20066,N_19858,N_19875);
and U20067 (N_20067,N_19802,N_19959);
xnor U20068 (N_20068,N_19820,N_19869);
or U20069 (N_20069,N_19821,N_19832);
and U20070 (N_20070,N_19927,N_19940);
nor U20071 (N_20071,N_19852,N_19877);
xor U20072 (N_20072,N_19855,N_19857);
xor U20073 (N_20073,N_19970,N_19829);
and U20074 (N_20074,N_19848,N_19895);
and U20075 (N_20075,N_19945,N_19968);
xor U20076 (N_20076,N_19886,N_19823);
xor U20077 (N_20077,N_19824,N_19921);
and U20078 (N_20078,N_19953,N_19990);
or U20079 (N_20079,N_19814,N_19939);
and U20080 (N_20080,N_19881,N_19849);
xnor U20081 (N_20081,N_19807,N_19860);
xnor U20082 (N_20082,N_19876,N_19977);
and U20083 (N_20083,N_19991,N_19969);
or U20084 (N_20084,N_19997,N_19842);
and U20085 (N_20085,N_19897,N_19981);
nor U20086 (N_20086,N_19837,N_19946);
or U20087 (N_20087,N_19812,N_19914);
and U20088 (N_20088,N_19979,N_19988);
and U20089 (N_20089,N_19948,N_19910);
nor U20090 (N_20090,N_19826,N_19925);
nor U20091 (N_20091,N_19908,N_19806);
and U20092 (N_20092,N_19834,N_19995);
nor U20093 (N_20093,N_19887,N_19958);
nor U20094 (N_20094,N_19917,N_19972);
nand U20095 (N_20095,N_19840,N_19957);
nand U20096 (N_20096,N_19825,N_19827);
nor U20097 (N_20097,N_19901,N_19811);
xnor U20098 (N_20098,N_19937,N_19982);
nand U20099 (N_20099,N_19918,N_19964);
nand U20100 (N_20100,N_19987,N_19810);
or U20101 (N_20101,N_19901,N_19987);
or U20102 (N_20102,N_19938,N_19881);
xnor U20103 (N_20103,N_19877,N_19963);
xnor U20104 (N_20104,N_19970,N_19897);
or U20105 (N_20105,N_19843,N_19889);
nor U20106 (N_20106,N_19942,N_19985);
and U20107 (N_20107,N_19989,N_19979);
nor U20108 (N_20108,N_19869,N_19843);
or U20109 (N_20109,N_19800,N_19804);
nand U20110 (N_20110,N_19870,N_19868);
and U20111 (N_20111,N_19935,N_19859);
xor U20112 (N_20112,N_19872,N_19852);
or U20113 (N_20113,N_19848,N_19947);
xor U20114 (N_20114,N_19812,N_19905);
and U20115 (N_20115,N_19841,N_19851);
or U20116 (N_20116,N_19999,N_19921);
or U20117 (N_20117,N_19857,N_19917);
and U20118 (N_20118,N_19825,N_19952);
or U20119 (N_20119,N_19820,N_19988);
nor U20120 (N_20120,N_19932,N_19966);
and U20121 (N_20121,N_19945,N_19936);
nor U20122 (N_20122,N_19832,N_19834);
nor U20123 (N_20123,N_19881,N_19856);
nand U20124 (N_20124,N_19911,N_19843);
and U20125 (N_20125,N_19845,N_19959);
or U20126 (N_20126,N_19978,N_19800);
xnor U20127 (N_20127,N_19916,N_19891);
nor U20128 (N_20128,N_19831,N_19864);
nor U20129 (N_20129,N_19852,N_19836);
and U20130 (N_20130,N_19983,N_19807);
or U20131 (N_20131,N_19912,N_19953);
or U20132 (N_20132,N_19843,N_19950);
nand U20133 (N_20133,N_19932,N_19862);
xor U20134 (N_20134,N_19962,N_19945);
and U20135 (N_20135,N_19940,N_19880);
and U20136 (N_20136,N_19978,N_19887);
and U20137 (N_20137,N_19873,N_19875);
or U20138 (N_20138,N_19937,N_19819);
nand U20139 (N_20139,N_19917,N_19849);
xnor U20140 (N_20140,N_19997,N_19948);
nand U20141 (N_20141,N_19946,N_19867);
and U20142 (N_20142,N_19894,N_19925);
and U20143 (N_20143,N_19988,N_19994);
nand U20144 (N_20144,N_19967,N_19857);
xor U20145 (N_20145,N_19803,N_19964);
nand U20146 (N_20146,N_19896,N_19846);
nor U20147 (N_20147,N_19807,N_19922);
xnor U20148 (N_20148,N_19823,N_19872);
nand U20149 (N_20149,N_19996,N_19874);
or U20150 (N_20150,N_19877,N_19987);
nand U20151 (N_20151,N_19985,N_19806);
nand U20152 (N_20152,N_19986,N_19975);
nor U20153 (N_20153,N_19951,N_19823);
or U20154 (N_20154,N_19840,N_19803);
nor U20155 (N_20155,N_19993,N_19938);
nor U20156 (N_20156,N_19806,N_19829);
nor U20157 (N_20157,N_19845,N_19828);
nand U20158 (N_20158,N_19948,N_19989);
and U20159 (N_20159,N_19929,N_19931);
xor U20160 (N_20160,N_19836,N_19984);
xor U20161 (N_20161,N_19814,N_19871);
and U20162 (N_20162,N_19914,N_19907);
or U20163 (N_20163,N_19946,N_19981);
or U20164 (N_20164,N_19965,N_19848);
or U20165 (N_20165,N_19902,N_19993);
nand U20166 (N_20166,N_19857,N_19885);
and U20167 (N_20167,N_19929,N_19989);
xnor U20168 (N_20168,N_19959,N_19828);
xor U20169 (N_20169,N_19806,N_19821);
xor U20170 (N_20170,N_19934,N_19865);
nor U20171 (N_20171,N_19834,N_19891);
and U20172 (N_20172,N_19975,N_19955);
xnor U20173 (N_20173,N_19912,N_19929);
nor U20174 (N_20174,N_19979,N_19905);
or U20175 (N_20175,N_19913,N_19955);
nor U20176 (N_20176,N_19806,N_19879);
or U20177 (N_20177,N_19907,N_19933);
xor U20178 (N_20178,N_19913,N_19806);
and U20179 (N_20179,N_19978,N_19933);
or U20180 (N_20180,N_19900,N_19847);
nand U20181 (N_20181,N_19926,N_19898);
nor U20182 (N_20182,N_19940,N_19897);
nor U20183 (N_20183,N_19837,N_19866);
and U20184 (N_20184,N_19974,N_19812);
and U20185 (N_20185,N_19807,N_19996);
xor U20186 (N_20186,N_19878,N_19931);
nor U20187 (N_20187,N_19894,N_19842);
and U20188 (N_20188,N_19846,N_19898);
nand U20189 (N_20189,N_19821,N_19825);
or U20190 (N_20190,N_19945,N_19948);
nand U20191 (N_20191,N_19807,N_19991);
nand U20192 (N_20192,N_19971,N_19984);
nand U20193 (N_20193,N_19907,N_19910);
or U20194 (N_20194,N_19915,N_19807);
nand U20195 (N_20195,N_19917,N_19996);
or U20196 (N_20196,N_19977,N_19973);
and U20197 (N_20197,N_19837,N_19830);
or U20198 (N_20198,N_19847,N_19994);
or U20199 (N_20199,N_19900,N_19858);
nand U20200 (N_20200,N_20118,N_20128);
nand U20201 (N_20201,N_20003,N_20131);
nor U20202 (N_20202,N_20053,N_20137);
or U20203 (N_20203,N_20020,N_20083);
nor U20204 (N_20204,N_20098,N_20019);
nor U20205 (N_20205,N_20102,N_20038);
nor U20206 (N_20206,N_20163,N_20146);
xnor U20207 (N_20207,N_20110,N_20107);
nor U20208 (N_20208,N_20196,N_20006);
nand U20209 (N_20209,N_20026,N_20180);
and U20210 (N_20210,N_20000,N_20181);
and U20211 (N_20211,N_20125,N_20060);
and U20212 (N_20212,N_20168,N_20139);
xor U20213 (N_20213,N_20112,N_20188);
nor U20214 (N_20214,N_20116,N_20122);
nand U20215 (N_20215,N_20094,N_20075);
or U20216 (N_20216,N_20045,N_20042);
xor U20217 (N_20217,N_20119,N_20143);
and U20218 (N_20218,N_20194,N_20176);
nor U20219 (N_20219,N_20059,N_20166);
nor U20220 (N_20220,N_20070,N_20023);
nand U20221 (N_20221,N_20198,N_20089);
xnor U20222 (N_20222,N_20113,N_20187);
nand U20223 (N_20223,N_20106,N_20174);
nand U20224 (N_20224,N_20104,N_20049);
nand U20225 (N_20225,N_20002,N_20140);
and U20226 (N_20226,N_20078,N_20080);
and U20227 (N_20227,N_20156,N_20037);
or U20228 (N_20228,N_20044,N_20056);
nor U20229 (N_20229,N_20197,N_20088);
nor U20230 (N_20230,N_20065,N_20158);
nand U20231 (N_20231,N_20073,N_20011);
nor U20232 (N_20232,N_20185,N_20012);
and U20233 (N_20233,N_20061,N_20082);
or U20234 (N_20234,N_20024,N_20177);
or U20235 (N_20235,N_20067,N_20154);
xor U20236 (N_20236,N_20048,N_20085);
nand U20237 (N_20237,N_20172,N_20121);
nor U20238 (N_20238,N_20199,N_20064);
xnor U20239 (N_20239,N_20159,N_20141);
xor U20240 (N_20240,N_20090,N_20165);
nor U20241 (N_20241,N_20079,N_20018);
xor U20242 (N_20242,N_20151,N_20057);
nor U20243 (N_20243,N_20150,N_20108);
nor U20244 (N_20244,N_20013,N_20136);
xnor U20245 (N_20245,N_20124,N_20130);
or U20246 (N_20246,N_20157,N_20160);
xnor U20247 (N_20247,N_20051,N_20015);
nand U20248 (N_20248,N_20091,N_20149);
and U20249 (N_20249,N_20126,N_20055);
or U20250 (N_20250,N_20092,N_20008);
xnor U20251 (N_20251,N_20007,N_20195);
xor U20252 (N_20252,N_20170,N_20175);
or U20253 (N_20253,N_20072,N_20111);
or U20254 (N_20254,N_20035,N_20145);
xor U20255 (N_20255,N_20178,N_20167);
xnor U20256 (N_20256,N_20043,N_20109);
and U20257 (N_20257,N_20164,N_20074);
or U20258 (N_20258,N_20148,N_20129);
or U20259 (N_20259,N_20014,N_20100);
and U20260 (N_20260,N_20142,N_20041);
xor U20261 (N_20261,N_20033,N_20147);
or U20262 (N_20262,N_20115,N_20179);
nor U20263 (N_20263,N_20039,N_20077);
nand U20264 (N_20264,N_20173,N_20096);
nand U20265 (N_20265,N_20120,N_20054);
or U20266 (N_20266,N_20021,N_20190);
nor U20267 (N_20267,N_20183,N_20114);
or U20268 (N_20268,N_20068,N_20093);
or U20269 (N_20269,N_20132,N_20087);
nand U20270 (N_20270,N_20022,N_20135);
and U20271 (N_20271,N_20063,N_20081);
or U20272 (N_20272,N_20030,N_20009);
xnor U20273 (N_20273,N_20017,N_20193);
or U20274 (N_20274,N_20162,N_20016);
nor U20275 (N_20275,N_20169,N_20192);
and U20276 (N_20276,N_20032,N_20027);
nor U20277 (N_20277,N_20047,N_20105);
and U20278 (N_20278,N_20028,N_20103);
nor U20279 (N_20279,N_20144,N_20101);
or U20280 (N_20280,N_20071,N_20086);
and U20281 (N_20281,N_20052,N_20152);
or U20282 (N_20282,N_20123,N_20034);
and U20283 (N_20283,N_20134,N_20133);
nor U20284 (N_20284,N_20171,N_20025);
xor U20285 (N_20285,N_20076,N_20184);
nand U20286 (N_20286,N_20069,N_20004);
xor U20287 (N_20287,N_20040,N_20097);
nand U20288 (N_20288,N_20010,N_20153);
nand U20289 (N_20289,N_20050,N_20005);
nor U20290 (N_20290,N_20036,N_20062);
nor U20291 (N_20291,N_20084,N_20117);
nor U20292 (N_20292,N_20058,N_20189);
and U20293 (N_20293,N_20029,N_20066);
or U20294 (N_20294,N_20099,N_20186);
nand U20295 (N_20295,N_20182,N_20001);
nor U20296 (N_20296,N_20095,N_20127);
nor U20297 (N_20297,N_20031,N_20191);
nand U20298 (N_20298,N_20155,N_20161);
nor U20299 (N_20299,N_20138,N_20046);
and U20300 (N_20300,N_20169,N_20107);
and U20301 (N_20301,N_20117,N_20096);
nand U20302 (N_20302,N_20051,N_20053);
nand U20303 (N_20303,N_20016,N_20020);
nor U20304 (N_20304,N_20024,N_20078);
and U20305 (N_20305,N_20049,N_20069);
nand U20306 (N_20306,N_20116,N_20134);
and U20307 (N_20307,N_20022,N_20045);
nor U20308 (N_20308,N_20011,N_20066);
xnor U20309 (N_20309,N_20107,N_20102);
nor U20310 (N_20310,N_20191,N_20143);
nor U20311 (N_20311,N_20057,N_20011);
nand U20312 (N_20312,N_20132,N_20103);
nor U20313 (N_20313,N_20002,N_20042);
nand U20314 (N_20314,N_20105,N_20010);
nand U20315 (N_20315,N_20140,N_20042);
and U20316 (N_20316,N_20000,N_20071);
and U20317 (N_20317,N_20176,N_20152);
xor U20318 (N_20318,N_20014,N_20047);
or U20319 (N_20319,N_20060,N_20129);
xor U20320 (N_20320,N_20070,N_20154);
nor U20321 (N_20321,N_20059,N_20048);
and U20322 (N_20322,N_20111,N_20003);
and U20323 (N_20323,N_20055,N_20180);
and U20324 (N_20324,N_20081,N_20019);
nand U20325 (N_20325,N_20061,N_20026);
nand U20326 (N_20326,N_20116,N_20151);
nand U20327 (N_20327,N_20020,N_20069);
or U20328 (N_20328,N_20057,N_20090);
and U20329 (N_20329,N_20087,N_20192);
or U20330 (N_20330,N_20003,N_20087);
nor U20331 (N_20331,N_20035,N_20089);
and U20332 (N_20332,N_20111,N_20017);
or U20333 (N_20333,N_20013,N_20082);
and U20334 (N_20334,N_20169,N_20156);
and U20335 (N_20335,N_20078,N_20153);
and U20336 (N_20336,N_20185,N_20192);
nand U20337 (N_20337,N_20191,N_20077);
and U20338 (N_20338,N_20080,N_20152);
or U20339 (N_20339,N_20145,N_20069);
xor U20340 (N_20340,N_20022,N_20012);
and U20341 (N_20341,N_20068,N_20188);
xor U20342 (N_20342,N_20059,N_20030);
nand U20343 (N_20343,N_20154,N_20099);
or U20344 (N_20344,N_20177,N_20098);
xor U20345 (N_20345,N_20112,N_20037);
and U20346 (N_20346,N_20193,N_20072);
xor U20347 (N_20347,N_20192,N_20005);
or U20348 (N_20348,N_20045,N_20132);
and U20349 (N_20349,N_20118,N_20164);
and U20350 (N_20350,N_20001,N_20183);
nand U20351 (N_20351,N_20181,N_20124);
and U20352 (N_20352,N_20157,N_20181);
and U20353 (N_20353,N_20102,N_20021);
nor U20354 (N_20354,N_20011,N_20044);
nand U20355 (N_20355,N_20099,N_20182);
nand U20356 (N_20356,N_20175,N_20141);
and U20357 (N_20357,N_20122,N_20080);
and U20358 (N_20358,N_20037,N_20004);
or U20359 (N_20359,N_20175,N_20064);
xor U20360 (N_20360,N_20142,N_20073);
xor U20361 (N_20361,N_20100,N_20170);
or U20362 (N_20362,N_20149,N_20047);
or U20363 (N_20363,N_20080,N_20051);
xor U20364 (N_20364,N_20016,N_20193);
nand U20365 (N_20365,N_20030,N_20153);
xnor U20366 (N_20366,N_20000,N_20033);
xor U20367 (N_20367,N_20123,N_20084);
xnor U20368 (N_20368,N_20040,N_20039);
nor U20369 (N_20369,N_20032,N_20100);
nor U20370 (N_20370,N_20111,N_20037);
nand U20371 (N_20371,N_20022,N_20072);
xor U20372 (N_20372,N_20115,N_20162);
nand U20373 (N_20373,N_20023,N_20127);
and U20374 (N_20374,N_20024,N_20131);
nor U20375 (N_20375,N_20090,N_20120);
xnor U20376 (N_20376,N_20076,N_20182);
nand U20377 (N_20377,N_20151,N_20187);
nor U20378 (N_20378,N_20018,N_20171);
and U20379 (N_20379,N_20133,N_20114);
nand U20380 (N_20380,N_20013,N_20144);
xor U20381 (N_20381,N_20124,N_20078);
xor U20382 (N_20382,N_20132,N_20110);
or U20383 (N_20383,N_20040,N_20178);
xnor U20384 (N_20384,N_20098,N_20123);
nand U20385 (N_20385,N_20031,N_20088);
xnor U20386 (N_20386,N_20084,N_20040);
nor U20387 (N_20387,N_20111,N_20095);
nor U20388 (N_20388,N_20080,N_20037);
and U20389 (N_20389,N_20085,N_20044);
or U20390 (N_20390,N_20152,N_20039);
or U20391 (N_20391,N_20027,N_20020);
nand U20392 (N_20392,N_20068,N_20178);
nand U20393 (N_20393,N_20064,N_20108);
or U20394 (N_20394,N_20135,N_20131);
nand U20395 (N_20395,N_20074,N_20167);
nor U20396 (N_20396,N_20047,N_20093);
nor U20397 (N_20397,N_20133,N_20173);
nand U20398 (N_20398,N_20103,N_20136);
nor U20399 (N_20399,N_20114,N_20030);
or U20400 (N_20400,N_20265,N_20352);
or U20401 (N_20401,N_20276,N_20391);
or U20402 (N_20402,N_20313,N_20215);
and U20403 (N_20403,N_20319,N_20230);
xnor U20404 (N_20404,N_20245,N_20251);
nor U20405 (N_20405,N_20229,N_20301);
and U20406 (N_20406,N_20308,N_20349);
xor U20407 (N_20407,N_20266,N_20343);
xnor U20408 (N_20408,N_20362,N_20360);
nor U20409 (N_20409,N_20398,N_20314);
and U20410 (N_20410,N_20297,N_20305);
nand U20411 (N_20411,N_20318,N_20292);
and U20412 (N_20412,N_20320,N_20397);
and U20413 (N_20413,N_20341,N_20203);
and U20414 (N_20414,N_20326,N_20329);
nor U20415 (N_20415,N_20270,N_20287);
xnor U20416 (N_20416,N_20296,N_20224);
or U20417 (N_20417,N_20261,N_20359);
nand U20418 (N_20418,N_20237,N_20200);
nand U20419 (N_20419,N_20365,N_20275);
xor U20420 (N_20420,N_20376,N_20274);
xor U20421 (N_20421,N_20221,N_20264);
and U20422 (N_20422,N_20307,N_20333);
xor U20423 (N_20423,N_20209,N_20395);
or U20424 (N_20424,N_20227,N_20234);
nand U20425 (N_20425,N_20290,N_20212);
nand U20426 (N_20426,N_20310,N_20220);
or U20427 (N_20427,N_20211,N_20210);
xor U20428 (N_20428,N_20249,N_20348);
or U20429 (N_20429,N_20241,N_20378);
xnor U20430 (N_20430,N_20259,N_20289);
nor U20431 (N_20431,N_20254,N_20280);
xnor U20432 (N_20432,N_20388,N_20337);
nor U20433 (N_20433,N_20207,N_20364);
nor U20434 (N_20434,N_20312,N_20253);
or U20435 (N_20435,N_20347,N_20371);
and U20436 (N_20436,N_20394,N_20380);
xor U20437 (N_20437,N_20255,N_20226);
nor U20438 (N_20438,N_20332,N_20344);
and U20439 (N_20439,N_20316,N_20279);
xor U20440 (N_20440,N_20260,N_20324);
xor U20441 (N_20441,N_20250,N_20322);
or U20442 (N_20442,N_20257,N_20225);
and U20443 (N_20443,N_20206,N_20384);
nand U20444 (N_20444,N_20235,N_20342);
nand U20445 (N_20445,N_20358,N_20258);
or U20446 (N_20446,N_20311,N_20370);
or U20447 (N_20447,N_20354,N_20334);
xor U20448 (N_20448,N_20315,N_20299);
or U20449 (N_20449,N_20294,N_20243);
xnor U20450 (N_20450,N_20351,N_20216);
and U20451 (N_20451,N_20240,N_20223);
nand U20452 (N_20452,N_20338,N_20238);
and U20453 (N_20453,N_20228,N_20377);
and U20454 (N_20454,N_20302,N_20295);
or U20455 (N_20455,N_20381,N_20357);
nand U20456 (N_20456,N_20291,N_20353);
nand U20457 (N_20457,N_20286,N_20217);
xnor U20458 (N_20458,N_20284,N_20214);
and U20459 (N_20459,N_20309,N_20233);
nor U20460 (N_20460,N_20373,N_20285);
nand U20461 (N_20461,N_20390,N_20263);
nor U20462 (N_20462,N_20386,N_20363);
nor U20463 (N_20463,N_20273,N_20303);
and U20464 (N_20464,N_20355,N_20244);
or U20465 (N_20465,N_20350,N_20372);
or U20466 (N_20466,N_20383,N_20246);
nor U20467 (N_20467,N_20361,N_20374);
nand U20468 (N_20468,N_20389,N_20204);
or U20469 (N_20469,N_20345,N_20262);
nor U20470 (N_20470,N_20321,N_20367);
nor U20471 (N_20471,N_20269,N_20239);
nor U20472 (N_20472,N_20325,N_20277);
xor U20473 (N_20473,N_20340,N_20293);
xor U20474 (N_20474,N_20248,N_20366);
xnor U20475 (N_20475,N_20327,N_20252);
or U20476 (N_20476,N_20282,N_20330);
nor U20477 (N_20477,N_20283,N_20346);
xor U20478 (N_20478,N_20201,N_20205);
and U20479 (N_20479,N_20232,N_20271);
nor U20480 (N_20480,N_20306,N_20396);
or U20481 (N_20481,N_20399,N_20213);
nor U20482 (N_20482,N_20219,N_20336);
nand U20483 (N_20483,N_20242,N_20331);
nand U20484 (N_20484,N_20202,N_20379);
and U20485 (N_20485,N_20231,N_20317);
nor U20486 (N_20486,N_20236,N_20304);
xor U20487 (N_20487,N_20356,N_20268);
or U20488 (N_20488,N_20300,N_20392);
xor U20489 (N_20489,N_20281,N_20375);
xor U20490 (N_20490,N_20385,N_20267);
or U20491 (N_20491,N_20222,N_20278);
nand U20492 (N_20492,N_20368,N_20328);
nand U20493 (N_20493,N_20339,N_20247);
nor U20494 (N_20494,N_20208,N_20335);
nand U20495 (N_20495,N_20288,N_20256);
nor U20496 (N_20496,N_20369,N_20382);
nor U20497 (N_20497,N_20393,N_20218);
xor U20498 (N_20498,N_20298,N_20387);
xnor U20499 (N_20499,N_20323,N_20272);
nor U20500 (N_20500,N_20288,N_20239);
and U20501 (N_20501,N_20366,N_20330);
or U20502 (N_20502,N_20296,N_20313);
nor U20503 (N_20503,N_20254,N_20263);
and U20504 (N_20504,N_20315,N_20357);
nand U20505 (N_20505,N_20346,N_20325);
and U20506 (N_20506,N_20310,N_20325);
and U20507 (N_20507,N_20260,N_20274);
nand U20508 (N_20508,N_20284,N_20346);
xor U20509 (N_20509,N_20316,N_20225);
xor U20510 (N_20510,N_20399,N_20214);
or U20511 (N_20511,N_20348,N_20246);
nor U20512 (N_20512,N_20208,N_20270);
nand U20513 (N_20513,N_20367,N_20225);
nand U20514 (N_20514,N_20222,N_20310);
and U20515 (N_20515,N_20384,N_20279);
nand U20516 (N_20516,N_20367,N_20216);
and U20517 (N_20517,N_20370,N_20218);
xnor U20518 (N_20518,N_20278,N_20308);
nand U20519 (N_20519,N_20388,N_20262);
nand U20520 (N_20520,N_20388,N_20216);
nand U20521 (N_20521,N_20340,N_20254);
xor U20522 (N_20522,N_20252,N_20390);
nor U20523 (N_20523,N_20302,N_20284);
or U20524 (N_20524,N_20268,N_20350);
xnor U20525 (N_20525,N_20358,N_20266);
and U20526 (N_20526,N_20362,N_20287);
nand U20527 (N_20527,N_20245,N_20318);
or U20528 (N_20528,N_20383,N_20275);
nand U20529 (N_20529,N_20363,N_20298);
nor U20530 (N_20530,N_20365,N_20200);
nor U20531 (N_20531,N_20237,N_20222);
nor U20532 (N_20532,N_20391,N_20374);
and U20533 (N_20533,N_20323,N_20203);
nor U20534 (N_20534,N_20367,N_20363);
nor U20535 (N_20535,N_20376,N_20333);
xnor U20536 (N_20536,N_20229,N_20370);
or U20537 (N_20537,N_20257,N_20320);
and U20538 (N_20538,N_20352,N_20387);
nand U20539 (N_20539,N_20360,N_20307);
xnor U20540 (N_20540,N_20382,N_20355);
and U20541 (N_20541,N_20279,N_20267);
nand U20542 (N_20542,N_20351,N_20349);
xor U20543 (N_20543,N_20237,N_20346);
and U20544 (N_20544,N_20350,N_20340);
and U20545 (N_20545,N_20294,N_20201);
nand U20546 (N_20546,N_20255,N_20346);
and U20547 (N_20547,N_20259,N_20358);
and U20548 (N_20548,N_20310,N_20205);
and U20549 (N_20549,N_20352,N_20294);
nand U20550 (N_20550,N_20247,N_20334);
nand U20551 (N_20551,N_20235,N_20201);
or U20552 (N_20552,N_20339,N_20378);
and U20553 (N_20553,N_20341,N_20267);
or U20554 (N_20554,N_20330,N_20341);
xor U20555 (N_20555,N_20365,N_20253);
or U20556 (N_20556,N_20260,N_20214);
or U20557 (N_20557,N_20271,N_20386);
or U20558 (N_20558,N_20235,N_20267);
xnor U20559 (N_20559,N_20336,N_20322);
nand U20560 (N_20560,N_20246,N_20379);
and U20561 (N_20561,N_20261,N_20231);
or U20562 (N_20562,N_20369,N_20226);
nand U20563 (N_20563,N_20242,N_20260);
nand U20564 (N_20564,N_20237,N_20334);
and U20565 (N_20565,N_20296,N_20254);
and U20566 (N_20566,N_20354,N_20286);
or U20567 (N_20567,N_20305,N_20210);
nor U20568 (N_20568,N_20318,N_20271);
and U20569 (N_20569,N_20220,N_20398);
xnor U20570 (N_20570,N_20232,N_20301);
nand U20571 (N_20571,N_20346,N_20305);
and U20572 (N_20572,N_20357,N_20257);
nand U20573 (N_20573,N_20355,N_20292);
and U20574 (N_20574,N_20398,N_20322);
or U20575 (N_20575,N_20276,N_20325);
xor U20576 (N_20576,N_20247,N_20254);
nand U20577 (N_20577,N_20273,N_20350);
nand U20578 (N_20578,N_20216,N_20343);
or U20579 (N_20579,N_20376,N_20307);
xor U20580 (N_20580,N_20389,N_20393);
or U20581 (N_20581,N_20288,N_20374);
and U20582 (N_20582,N_20295,N_20315);
nand U20583 (N_20583,N_20348,N_20245);
and U20584 (N_20584,N_20218,N_20231);
nor U20585 (N_20585,N_20242,N_20279);
or U20586 (N_20586,N_20212,N_20329);
xnor U20587 (N_20587,N_20381,N_20360);
nand U20588 (N_20588,N_20351,N_20222);
xor U20589 (N_20589,N_20345,N_20396);
nor U20590 (N_20590,N_20229,N_20359);
xnor U20591 (N_20591,N_20265,N_20226);
nor U20592 (N_20592,N_20283,N_20238);
and U20593 (N_20593,N_20358,N_20260);
nor U20594 (N_20594,N_20295,N_20311);
or U20595 (N_20595,N_20256,N_20244);
nor U20596 (N_20596,N_20263,N_20257);
or U20597 (N_20597,N_20322,N_20318);
nand U20598 (N_20598,N_20238,N_20202);
or U20599 (N_20599,N_20378,N_20392);
and U20600 (N_20600,N_20402,N_20412);
and U20601 (N_20601,N_20590,N_20456);
nor U20602 (N_20602,N_20559,N_20561);
or U20603 (N_20603,N_20499,N_20430);
and U20604 (N_20604,N_20485,N_20481);
xnor U20605 (N_20605,N_20578,N_20471);
and U20606 (N_20606,N_20409,N_20567);
nor U20607 (N_20607,N_20519,N_20426);
or U20608 (N_20608,N_20553,N_20560);
nor U20609 (N_20609,N_20483,N_20515);
nand U20610 (N_20610,N_20546,N_20507);
nor U20611 (N_20611,N_20562,N_20452);
nand U20612 (N_20612,N_20432,N_20551);
or U20613 (N_20613,N_20543,N_20512);
nand U20614 (N_20614,N_20447,N_20487);
and U20615 (N_20615,N_20479,N_20580);
nor U20616 (N_20616,N_20587,N_20407);
nand U20617 (N_20617,N_20522,N_20542);
or U20618 (N_20618,N_20511,N_20453);
and U20619 (N_20619,N_20589,N_20526);
nand U20620 (N_20620,N_20448,N_20540);
xnor U20621 (N_20621,N_20595,N_20464);
or U20622 (N_20622,N_20476,N_20572);
nor U20623 (N_20623,N_20514,N_20575);
and U20624 (N_20624,N_20484,N_20585);
nand U20625 (N_20625,N_20583,N_20556);
nand U20626 (N_20626,N_20529,N_20573);
nand U20627 (N_20627,N_20442,N_20461);
nand U20628 (N_20628,N_20433,N_20474);
xor U20629 (N_20629,N_20552,N_20450);
nand U20630 (N_20630,N_20591,N_20494);
nand U20631 (N_20631,N_20422,N_20523);
or U20632 (N_20632,N_20531,N_20404);
nor U20633 (N_20633,N_20469,N_20574);
xor U20634 (N_20634,N_20405,N_20425);
xor U20635 (N_20635,N_20538,N_20466);
nand U20636 (N_20636,N_20576,N_20581);
xnor U20637 (N_20637,N_20594,N_20586);
xnor U20638 (N_20638,N_20548,N_20557);
nor U20639 (N_20639,N_20416,N_20446);
nor U20640 (N_20640,N_20545,N_20443);
and U20641 (N_20641,N_20457,N_20439);
or U20642 (N_20642,N_20569,N_20537);
xnor U20643 (N_20643,N_20510,N_20534);
nand U20644 (N_20644,N_20525,N_20527);
or U20645 (N_20645,N_20565,N_20536);
and U20646 (N_20646,N_20488,N_20584);
nor U20647 (N_20647,N_20570,N_20504);
or U20648 (N_20648,N_20478,N_20541);
and U20649 (N_20649,N_20493,N_20440);
nand U20650 (N_20650,N_20413,N_20579);
and U20651 (N_20651,N_20418,N_20555);
nand U20652 (N_20652,N_20568,N_20477);
nand U20653 (N_20653,N_20475,N_20500);
or U20654 (N_20654,N_20410,N_20431);
xor U20655 (N_20655,N_20521,N_20518);
or U20656 (N_20656,N_20473,N_20459);
nand U20657 (N_20657,N_20539,N_20592);
and U20658 (N_20658,N_20470,N_20454);
nor U20659 (N_20659,N_20505,N_20554);
or U20660 (N_20660,N_20427,N_20463);
and U20661 (N_20661,N_20490,N_20520);
xor U20662 (N_20662,N_20455,N_20403);
or U20663 (N_20663,N_20417,N_20482);
nand U20664 (N_20664,N_20506,N_20462);
nand U20665 (N_20665,N_20435,N_20444);
xor U20666 (N_20666,N_20419,N_20516);
xor U20667 (N_20667,N_20564,N_20437);
and U20668 (N_20668,N_20434,N_20460);
and U20669 (N_20669,N_20597,N_20550);
xnor U20670 (N_20670,N_20429,N_20492);
nand U20671 (N_20671,N_20401,N_20428);
xnor U20672 (N_20672,N_20502,N_20438);
nand U20673 (N_20673,N_20524,N_20415);
or U20674 (N_20674,N_20495,N_20468);
and U20675 (N_20675,N_20436,N_20549);
or U20676 (N_20676,N_20558,N_20598);
or U20677 (N_20677,N_20577,N_20593);
or U20678 (N_20678,N_20563,N_20599);
nor U20679 (N_20679,N_20486,N_20491);
and U20680 (N_20680,N_20421,N_20596);
nand U20681 (N_20681,N_20414,N_20503);
or U20682 (N_20682,N_20406,N_20420);
or U20683 (N_20683,N_20496,N_20513);
nand U20684 (N_20684,N_20400,N_20535);
xnor U20685 (N_20685,N_20497,N_20472);
xnor U20686 (N_20686,N_20451,N_20480);
nor U20687 (N_20687,N_20509,N_20489);
or U20688 (N_20688,N_20571,N_20467);
nand U20689 (N_20689,N_20408,N_20449);
xnor U20690 (N_20690,N_20445,N_20533);
nor U20691 (N_20691,N_20411,N_20528);
nand U20692 (N_20692,N_20544,N_20465);
or U20693 (N_20693,N_20508,N_20530);
nor U20694 (N_20694,N_20566,N_20547);
nand U20695 (N_20695,N_20458,N_20498);
nor U20696 (N_20696,N_20582,N_20441);
or U20697 (N_20697,N_20588,N_20501);
nor U20698 (N_20698,N_20424,N_20423);
nor U20699 (N_20699,N_20517,N_20532);
or U20700 (N_20700,N_20577,N_20589);
or U20701 (N_20701,N_20555,N_20594);
nand U20702 (N_20702,N_20430,N_20563);
nand U20703 (N_20703,N_20400,N_20585);
and U20704 (N_20704,N_20454,N_20449);
and U20705 (N_20705,N_20517,N_20580);
nor U20706 (N_20706,N_20504,N_20506);
xnor U20707 (N_20707,N_20494,N_20409);
or U20708 (N_20708,N_20557,N_20441);
xor U20709 (N_20709,N_20440,N_20425);
or U20710 (N_20710,N_20423,N_20430);
nand U20711 (N_20711,N_20525,N_20556);
nor U20712 (N_20712,N_20524,N_20580);
and U20713 (N_20713,N_20546,N_20529);
or U20714 (N_20714,N_20544,N_20473);
xnor U20715 (N_20715,N_20533,N_20591);
and U20716 (N_20716,N_20497,N_20517);
nand U20717 (N_20717,N_20469,N_20558);
or U20718 (N_20718,N_20490,N_20518);
nand U20719 (N_20719,N_20545,N_20439);
and U20720 (N_20720,N_20526,N_20515);
nor U20721 (N_20721,N_20547,N_20499);
nand U20722 (N_20722,N_20487,N_20529);
nand U20723 (N_20723,N_20477,N_20503);
xor U20724 (N_20724,N_20553,N_20471);
or U20725 (N_20725,N_20429,N_20433);
nor U20726 (N_20726,N_20556,N_20515);
nand U20727 (N_20727,N_20423,N_20411);
nor U20728 (N_20728,N_20555,N_20559);
xnor U20729 (N_20729,N_20517,N_20455);
xnor U20730 (N_20730,N_20542,N_20548);
and U20731 (N_20731,N_20528,N_20593);
nand U20732 (N_20732,N_20427,N_20457);
xor U20733 (N_20733,N_20525,N_20559);
nor U20734 (N_20734,N_20432,N_20542);
xor U20735 (N_20735,N_20513,N_20582);
or U20736 (N_20736,N_20504,N_20582);
xnor U20737 (N_20737,N_20402,N_20545);
or U20738 (N_20738,N_20597,N_20426);
or U20739 (N_20739,N_20522,N_20474);
and U20740 (N_20740,N_20429,N_20563);
or U20741 (N_20741,N_20459,N_20477);
xor U20742 (N_20742,N_20558,N_20580);
nand U20743 (N_20743,N_20466,N_20576);
and U20744 (N_20744,N_20448,N_20539);
and U20745 (N_20745,N_20424,N_20496);
or U20746 (N_20746,N_20515,N_20423);
and U20747 (N_20747,N_20427,N_20508);
and U20748 (N_20748,N_20498,N_20591);
nor U20749 (N_20749,N_20426,N_20516);
or U20750 (N_20750,N_20409,N_20474);
nor U20751 (N_20751,N_20483,N_20595);
and U20752 (N_20752,N_20481,N_20528);
and U20753 (N_20753,N_20510,N_20515);
nor U20754 (N_20754,N_20473,N_20576);
nor U20755 (N_20755,N_20529,N_20485);
and U20756 (N_20756,N_20581,N_20531);
or U20757 (N_20757,N_20450,N_20525);
and U20758 (N_20758,N_20580,N_20520);
xor U20759 (N_20759,N_20582,N_20554);
or U20760 (N_20760,N_20475,N_20444);
or U20761 (N_20761,N_20561,N_20599);
xnor U20762 (N_20762,N_20427,N_20413);
nand U20763 (N_20763,N_20449,N_20562);
nand U20764 (N_20764,N_20408,N_20465);
nand U20765 (N_20765,N_20435,N_20560);
and U20766 (N_20766,N_20569,N_20455);
xnor U20767 (N_20767,N_20403,N_20409);
or U20768 (N_20768,N_20511,N_20444);
and U20769 (N_20769,N_20470,N_20441);
nand U20770 (N_20770,N_20576,N_20454);
xor U20771 (N_20771,N_20553,N_20570);
nand U20772 (N_20772,N_20583,N_20551);
or U20773 (N_20773,N_20494,N_20484);
nand U20774 (N_20774,N_20574,N_20485);
xnor U20775 (N_20775,N_20410,N_20497);
and U20776 (N_20776,N_20449,N_20471);
nand U20777 (N_20777,N_20474,N_20475);
or U20778 (N_20778,N_20575,N_20533);
xnor U20779 (N_20779,N_20488,N_20568);
nor U20780 (N_20780,N_20431,N_20443);
or U20781 (N_20781,N_20405,N_20500);
xnor U20782 (N_20782,N_20572,N_20571);
or U20783 (N_20783,N_20577,N_20476);
and U20784 (N_20784,N_20445,N_20482);
or U20785 (N_20785,N_20525,N_20477);
nand U20786 (N_20786,N_20595,N_20504);
and U20787 (N_20787,N_20580,N_20585);
or U20788 (N_20788,N_20539,N_20527);
nor U20789 (N_20789,N_20574,N_20505);
or U20790 (N_20790,N_20409,N_20418);
xor U20791 (N_20791,N_20444,N_20455);
xnor U20792 (N_20792,N_20446,N_20499);
nor U20793 (N_20793,N_20477,N_20425);
and U20794 (N_20794,N_20489,N_20466);
or U20795 (N_20795,N_20512,N_20499);
and U20796 (N_20796,N_20490,N_20571);
nand U20797 (N_20797,N_20446,N_20525);
nand U20798 (N_20798,N_20432,N_20464);
nor U20799 (N_20799,N_20410,N_20559);
xor U20800 (N_20800,N_20757,N_20652);
and U20801 (N_20801,N_20638,N_20730);
xor U20802 (N_20802,N_20601,N_20664);
or U20803 (N_20803,N_20752,N_20789);
nand U20804 (N_20804,N_20653,N_20700);
and U20805 (N_20805,N_20764,N_20655);
xnor U20806 (N_20806,N_20703,N_20722);
nor U20807 (N_20807,N_20650,N_20733);
xnor U20808 (N_20808,N_20683,N_20603);
nor U20809 (N_20809,N_20635,N_20748);
xnor U20810 (N_20810,N_20774,N_20696);
and U20811 (N_20811,N_20720,N_20662);
or U20812 (N_20812,N_20646,N_20672);
xor U20813 (N_20813,N_20624,N_20745);
xnor U20814 (N_20814,N_20609,N_20702);
and U20815 (N_20815,N_20681,N_20780);
or U20816 (N_20816,N_20747,N_20616);
nor U20817 (N_20817,N_20677,N_20643);
nor U20818 (N_20818,N_20671,N_20682);
and U20819 (N_20819,N_20791,N_20642);
nand U20820 (N_20820,N_20699,N_20695);
or U20821 (N_20821,N_20763,N_20792);
nand U20822 (N_20822,N_20641,N_20736);
nand U20823 (N_20823,N_20793,N_20607);
nor U20824 (N_20824,N_20644,N_20735);
nand U20825 (N_20825,N_20782,N_20628);
or U20826 (N_20826,N_20670,N_20790);
nand U20827 (N_20827,N_20694,N_20785);
nand U20828 (N_20828,N_20765,N_20654);
nand U20829 (N_20829,N_20719,N_20734);
nor U20830 (N_20830,N_20714,N_20631);
xor U20831 (N_20831,N_20685,N_20770);
nand U20832 (N_20832,N_20731,N_20687);
or U20833 (N_20833,N_20622,N_20726);
xnor U20834 (N_20834,N_20612,N_20648);
xor U20835 (N_20835,N_20718,N_20675);
nand U20836 (N_20836,N_20729,N_20658);
and U20837 (N_20837,N_20740,N_20629);
nor U20838 (N_20838,N_20777,N_20759);
or U20839 (N_20839,N_20794,N_20766);
and U20840 (N_20840,N_20625,N_20620);
nand U20841 (N_20841,N_20713,N_20799);
and U20842 (N_20842,N_20649,N_20787);
and U20843 (N_20843,N_20665,N_20617);
nand U20844 (N_20844,N_20712,N_20636);
and U20845 (N_20845,N_20661,N_20773);
xnor U20846 (N_20846,N_20753,N_20725);
or U20847 (N_20847,N_20632,N_20627);
nand U20848 (N_20848,N_20637,N_20688);
and U20849 (N_20849,N_20769,N_20710);
xnor U20850 (N_20850,N_20760,N_20709);
and U20851 (N_20851,N_20647,N_20723);
nor U20852 (N_20852,N_20678,N_20724);
and U20853 (N_20853,N_20608,N_20684);
nand U20854 (N_20854,N_20744,N_20679);
and U20855 (N_20855,N_20743,N_20772);
or U20856 (N_20856,N_20614,N_20663);
or U20857 (N_20857,N_20640,N_20610);
xnor U20858 (N_20858,N_20676,N_20645);
nand U20859 (N_20859,N_20657,N_20781);
and U20860 (N_20860,N_20613,N_20680);
nor U20861 (N_20861,N_20707,N_20693);
xor U20862 (N_20862,N_20715,N_20758);
and U20863 (N_20863,N_20775,N_20756);
or U20864 (N_20864,N_20600,N_20605);
nor U20865 (N_20865,N_20690,N_20737);
nand U20866 (N_20866,N_20784,N_20630);
xnor U20867 (N_20867,N_20786,N_20674);
and U20868 (N_20868,N_20762,N_20761);
and U20869 (N_20869,N_20746,N_20692);
nor U20870 (N_20870,N_20711,N_20667);
nor U20871 (N_20871,N_20689,N_20669);
or U20872 (N_20872,N_20660,N_20795);
and U20873 (N_20873,N_20656,N_20673);
and U20874 (N_20874,N_20691,N_20615);
and U20875 (N_20875,N_20732,N_20717);
and U20876 (N_20876,N_20704,N_20716);
xor U20877 (N_20877,N_20626,N_20767);
and U20878 (N_20878,N_20755,N_20705);
nand U20879 (N_20879,N_20788,N_20721);
nor U20880 (N_20880,N_20659,N_20779);
xor U20881 (N_20881,N_20771,N_20741);
and U20882 (N_20882,N_20611,N_20604);
xor U20883 (N_20883,N_20639,N_20750);
nor U20884 (N_20884,N_20697,N_20776);
xor U20885 (N_20885,N_20738,N_20602);
or U20886 (N_20886,N_20778,N_20606);
nor U20887 (N_20887,N_20727,N_20618);
or U20888 (N_20888,N_20621,N_20749);
and U20889 (N_20889,N_20633,N_20798);
nand U20890 (N_20890,N_20651,N_20797);
nor U20891 (N_20891,N_20698,N_20796);
xor U20892 (N_20892,N_20783,N_20754);
xor U20893 (N_20893,N_20739,N_20728);
nor U20894 (N_20894,N_20768,N_20668);
or U20895 (N_20895,N_20706,N_20701);
or U20896 (N_20896,N_20623,N_20666);
and U20897 (N_20897,N_20742,N_20634);
xnor U20898 (N_20898,N_20686,N_20708);
or U20899 (N_20899,N_20751,N_20619);
nand U20900 (N_20900,N_20726,N_20754);
nand U20901 (N_20901,N_20751,N_20660);
xor U20902 (N_20902,N_20649,N_20752);
nand U20903 (N_20903,N_20728,N_20743);
nand U20904 (N_20904,N_20775,N_20609);
nor U20905 (N_20905,N_20780,N_20634);
and U20906 (N_20906,N_20671,N_20767);
xnor U20907 (N_20907,N_20644,N_20617);
xnor U20908 (N_20908,N_20659,N_20677);
nor U20909 (N_20909,N_20739,N_20755);
nor U20910 (N_20910,N_20745,N_20662);
or U20911 (N_20911,N_20685,N_20611);
nor U20912 (N_20912,N_20668,N_20715);
nand U20913 (N_20913,N_20756,N_20726);
xnor U20914 (N_20914,N_20773,N_20630);
or U20915 (N_20915,N_20696,N_20766);
nor U20916 (N_20916,N_20795,N_20606);
xnor U20917 (N_20917,N_20689,N_20685);
and U20918 (N_20918,N_20615,N_20686);
xor U20919 (N_20919,N_20687,N_20672);
or U20920 (N_20920,N_20791,N_20708);
and U20921 (N_20921,N_20652,N_20622);
nor U20922 (N_20922,N_20771,N_20618);
and U20923 (N_20923,N_20696,N_20748);
xor U20924 (N_20924,N_20789,N_20695);
xnor U20925 (N_20925,N_20670,N_20783);
or U20926 (N_20926,N_20682,N_20707);
xor U20927 (N_20927,N_20618,N_20764);
nor U20928 (N_20928,N_20760,N_20630);
xnor U20929 (N_20929,N_20679,N_20778);
or U20930 (N_20930,N_20723,N_20738);
and U20931 (N_20931,N_20602,N_20708);
or U20932 (N_20932,N_20722,N_20672);
or U20933 (N_20933,N_20666,N_20687);
and U20934 (N_20934,N_20682,N_20797);
xor U20935 (N_20935,N_20655,N_20635);
or U20936 (N_20936,N_20644,N_20689);
or U20937 (N_20937,N_20720,N_20769);
or U20938 (N_20938,N_20677,N_20753);
or U20939 (N_20939,N_20745,N_20765);
nand U20940 (N_20940,N_20636,N_20655);
and U20941 (N_20941,N_20624,N_20697);
nor U20942 (N_20942,N_20691,N_20759);
and U20943 (N_20943,N_20616,N_20791);
nand U20944 (N_20944,N_20637,N_20763);
nor U20945 (N_20945,N_20726,N_20677);
nor U20946 (N_20946,N_20653,N_20787);
or U20947 (N_20947,N_20744,N_20740);
nor U20948 (N_20948,N_20622,N_20722);
nand U20949 (N_20949,N_20792,N_20775);
nor U20950 (N_20950,N_20684,N_20687);
xnor U20951 (N_20951,N_20745,N_20783);
nand U20952 (N_20952,N_20768,N_20694);
nor U20953 (N_20953,N_20773,N_20645);
nor U20954 (N_20954,N_20690,N_20652);
xnor U20955 (N_20955,N_20769,N_20682);
or U20956 (N_20956,N_20728,N_20782);
and U20957 (N_20957,N_20760,N_20639);
nand U20958 (N_20958,N_20766,N_20666);
or U20959 (N_20959,N_20758,N_20650);
nor U20960 (N_20960,N_20636,N_20600);
and U20961 (N_20961,N_20707,N_20664);
and U20962 (N_20962,N_20608,N_20619);
and U20963 (N_20963,N_20746,N_20644);
or U20964 (N_20964,N_20786,N_20740);
or U20965 (N_20965,N_20619,N_20726);
nor U20966 (N_20966,N_20702,N_20605);
and U20967 (N_20967,N_20627,N_20698);
xnor U20968 (N_20968,N_20744,N_20715);
nand U20969 (N_20969,N_20647,N_20601);
or U20970 (N_20970,N_20782,N_20618);
nand U20971 (N_20971,N_20795,N_20756);
nand U20972 (N_20972,N_20742,N_20647);
nand U20973 (N_20973,N_20686,N_20782);
nand U20974 (N_20974,N_20737,N_20618);
or U20975 (N_20975,N_20605,N_20640);
and U20976 (N_20976,N_20767,N_20715);
and U20977 (N_20977,N_20756,N_20672);
nor U20978 (N_20978,N_20686,N_20683);
xor U20979 (N_20979,N_20652,N_20730);
and U20980 (N_20980,N_20626,N_20695);
nor U20981 (N_20981,N_20617,N_20623);
nand U20982 (N_20982,N_20789,N_20756);
or U20983 (N_20983,N_20620,N_20734);
nand U20984 (N_20984,N_20733,N_20608);
nand U20985 (N_20985,N_20670,N_20671);
nor U20986 (N_20986,N_20687,N_20770);
xnor U20987 (N_20987,N_20750,N_20636);
and U20988 (N_20988,N_20649,N_20668);
or U20989 (N_20989,N_20749,N_20732);
or U20990 (N_20990,N_20676,N_20677);
or U20991 (N_20991,N_20606,N_20672);
nor U20992 (N_20992,N_20765,N_20757);
nor U20993 (N_20993,N_20781,N_20760);
and U20994 (N_20994,N_20624,N_20758);
nor U20995 (N_20995,N_20792,N_20663);
nor U20996 (N_20996,N_20749,N_20737);
and U20997 (N_20997,N_20777,N_20629);
xor U20998 (N_20998,N_20635,N_20694);
nor U20999 (N_20999,N_20738,N_20776);
or U21000 (N_21000,N_20876,N_20993);
and U21001 (N_21001,N_20855,N_20902);
nor U21002 (N_21002,N_20839,N_20975);
nor U21003 (N_21003,N_20892,N_20987);
xnor U21004 (N_21004,N_20906,N_20886);
nor U21005 (N_21005,N_20872,N_20895);
xnor U21006 (N_21006,N_20831,N_20953);
or U21007 (N_21007,N_20933,N_20832);
nand U21008 (N_21008,N_20907,N_20891);
nand U21009 (N_21009,N_20968,N_20835);
xnor U21010 (N_21010,N_20856,N_20900);
xor U21011 (N_21011,N_20901,N_20913);
and U21012 (N_21012,N_20860,N_20946);
or U21013 (N_21013,N_20914,N_20998);
nor U21014 (N_21014,N_20821,N_20814);
and U21015 (N_21015,N_20930,N_20801);
nor U21016 (N_21016,N_20899,N_20807);
xnor U21017 (N_21017,N_20863,N_20820);
and U21018 (N_21018,N_20878,N_20961);
nand U21019 (N_21019,N_20818,N_20828);
nor U21020 (N_21020,N_20875,N_20824);
and U21021 (N_21021,N_20850,N_20843);
or U21022 (N_21022,N_20927,N_20874);
xnor U21023 (N_21023,N_20978,N_20905);
nor U21024 (N_21024,N_20898,N_20981);
nor U21025 (N_21025,N_20962,N_20883);
nor U21026 (N_21026,N_20897,N_20811);
xnor U21027 (N_21027,N_20971,N_20825);
or U21028 (N_21028,N_20880,N_20826);
nand U21029 (N_21029,N_20849,N_20890);
xnor U21030 (N_21030,N_20848,N_20806);
nor U21031 (N_21031,N_20974,N_20887);
nor U21032 (N_21032,N_20857,N_20808);
or U21033 (N_21033,N_20884,N_20859);
or U21034 (N_21034,N_20959,N_20809);
nor U21035 (N_21035,N_20896,N_20924);
and U21036 (N_21036,N_20908,N_20979);
nor U21037 (N_21037,N_20985,N_20973);
nor U21038 (N_21038,N_20869,N_20997);
xnor U21039 (N_21039,N_20847,N_20947);
and U21040 (N_21040,N_20964,N_20939);
nand U21041 (N_21041,N_20800,N_20938);
or U21042 (N_21042,N_20945,N_20912);
nor U21043 (N_21043,N_20911,N_20941);
nor U21044 (N_21044,N_20852,N_20846);
nor U21045 (N_21045,N_20980,N_20858);
or U21046 (N_21046,N_20977,N_20802);
or U21047 (N_21047,N_20804,N_20810);
xnor U21048 (N_21048,N_20982,N_20958);
xor U21049 (N_21049,N_20925,N_20837);
nand U21050 (N_21050,N_20954,N_20816);
and U21051 (N_21051,N_20950,N_20833);
or U21052 (N_21052,N_20935,N_20984);
nor U21053 (N_21053,N_20989,N_20862);
and U21054 (N_21054,N_20937,N_20995);
nand U21055 (N_21055,N_20873,N_20879);
xor U21056 (N_21056,N_20819,N_20991);
nand U21057 (N_21057,N_20822,N_20932);
or U21058 (N_21058,N_20919,N_20903);
nand U21059 (N_21059,N_20836,N_20817);
or U21060 (N_21060,N_20877,N_20894);
nor U21061 (N_21061,N_20923,N_20861);
and U21062 (N_21062,N_20922,N_20909);
nand U21063 (N_21063,N_20868,N_20830);
and U21064 (N_21064,N_20967,N_20917);
xnor U21065 (N_21065,N_20910,N_20842);
nand U21066 (N_21066,N_20803,N_20960);
or U21067 (N_21067,N_20934,N_20823);
nand U21068 (N_21068,N_20996,N_20812);
and U21069 (N_21069,N_20844,N_20885);
nor U21070 (N_21070,N_20936,N_20965);
or U21071 (N_21071,N_20969,N_20867);
xor U21072 (N_21072,N_20841,N_20840);
or U21073 (N_21073,N_20851,N_20918);
xnor U21074 (N_21074,N_20813,N_20882);
or U21075 (N_21075,N_20915,N_20992);
or U21076 (N_21076,N_20949,N_20904);
and U21077 (N_21077,N_20931,N_20952);
and U21078 (N_21078,N_20999,N_20951);
or U21079 (N_21079,N_20955,N_20845);
or U21080 (N_21080,N_20865,N_20976);
and U21081 (N_21081,N_20994,N_20943);
and U21082 (N_21082,N_20815,N_20834);
nand U21083 (N_21083,N_20966,N_20805);
and U21084 (N_21084,N_20948,N_20838);
nor U21085 (N_21085,N_20881,N_20866);
and U21086 (N_21086,N_20983,N_20972);
nand U21087 (N_21087,N_20893,N_20942);
nand U21088 (N_21088,N_20854,N_20940);
xnor U21089 (N_21089,N_20853,N_20944);
xnor U21090 (N_21090,N_20956,N_20990);
nand U21091 (N_21091,N_20963,N_20864);
nor U21092 (N_21092,N_20870,N_20916);
nor U21093 (N_21093,N_20829,N_20929);
nand U21094 (N_21094,N_20889,N_20827);
and U21095 (N_21095,N_20928,N_20988);
nand U21096 (N_21096,N_20986,N_20921);
xor U21097 (N_21097,N_20920,N_20888);
xor U21098 (N_21098,N_20957,N_20970);
nand U21099 (N_21099,N_20926,N_20871);
and U21100 (N_21100,N_20839,N_20864);
nor U21101 (N_21101,N_20946,N_20842);
xor U21102 (N_21102,N_20881,N_20875);
or U21103 (N_21103,N_20833,N_20997);
and U21104 (N_21104,N_20916,N_20967);
or U21105 (N_21105,N_20906,N_20832);
nand U21106 (N_21106,N_20985,N_20815);
and U21107 (N_21107,N_20932,N_20971);
xnor U21108 (N_21108,N_20884,N_20925);
nand U21109 (N_21109,N_20891,N_20992);
nor U21110 (N_21110,N_20845,N_20819);
nand U21111 (N_21111,N_20960,N_20920);
or U21112 (N_21112,N_20840,N_20966);
nand U21113 (N_21113,N_20887,N_20894);
or U21114 (N_21114,N_20967,N_20834);
nor U21115 (N_21115,N_20989,N_20806);
nor U21116 (N_21116,N_20817,N_20947);
nand U21117 (N_21117,N_20954,N_20913);
nor U21118 (N_21118,N_20926,N_20816);
or U21119 (N_21119,N_20822,N_20994);
or U21120 (N_21120,N_20916,N_20850);
xor U21121 (N_21121,N_20820,N_20979);
nand U21122 (N_21122,N_20857,N_20807);
xor U21123 (N_21123,N_20923,N_20822);
xnor U21124 (N_21124,N_20911,N_20910);
or U21125 (N_21125,N_20922,N_20884);
and U21126 (N_21126,N_20869,N_20992);
nand U21127 (N_21127,N_20925,N_20977);
and U21128 (N_21128,N_20898,N_20955);
nor U21129 (N_21129,N_20828,N_20974);
or U21130 (N_21130,N_20996,N_20860);
nor U21131 (N_21131,N_20858,N_20920);
xor U21132 (N_21132,N_20818,N_20815);
nand U21133 (N_21133,N_20850,N_20886);
nand U21134 (N_21134,N_20847,N_20853);
and U21135 (N_21135,N_20940,N_20981);
or U21136 (N_21136,N_20895,N_20965);
xnor U21137 (N_21137,N_20802,N_20905);
and U21138 (N_21138,N_20965,N_20947);
and U21139 (N_21139,N_20940,N_20994);
nand U21140 (N_21140,N_20910,N_20933);
and U21141 (N_21141,N_20899,N_20910);
and U21142 (N_21142,N_20990,N_20910);
and U21143 (N_21143,N_20891,N_20847);
and U21144 (N_21144,N_20904,N_20981);
nand U21145 (N_21145,N_20887,N_20899);
xor U21146 (N_21146,N_20837,N_20884);
and U21147 (N_21147,N_20903,N_20857);
and U21148 (N_21148,N_20969,N_20972);
or U21149 (N_21149,N_20846,N_20883);
nor U21150 (N_21150,N_20968,N_20856);
nor U21151 (N_21151,N_20940,N_20922);
xor U21152 (N_21152,N_20887,N_20948);
nand U21153 (N_21153,N_20965,N_20998);
nor U21154 (N_21154,N_20939,N_20922);
nand U21155 (N_21155,N_20851,N_20842);
xnor U21156 (N_21156,N_20897,N_20921);
and U21157 (N_21157,N_20897,N_20933);
xnor U21158 (N_21158,N_20972,N_20817);
nand U21159 (N_21159,N_20915,N_20935);
and U21160 (N_21160,N_20973,N_20952);
or U21161 (N_21161,N_20910,N_20996);
xnor U21162 (N_21162,N_20999,N_20940);
and U21163 (N_21163,N_20975,N_20901);
nand U21164 (N_21164,N_20892,N_20852);
or U21165 (N_21165,N_20992,N_20978);
and U21166 (N_21166,N_20932,N_20880);
or U21167 (N_21167,N_20892,N_20906);
nor U21168 (N_21168,N_20966,N_20890);
or U21169 (N_21169,N_20952,N_20835);
nor U21170 (N_21170,N_20901,N_20951);
and U21171 (N_21171,N_20903,N_20813);
xnor U21172 (N_21172,N_20971,N_20997);
xnor U21173 (N_21173,N_20814,N_20860);
xnor U21174 (N_21174,N_20833,N_20866);
or U21175 (N_21175,N_20975,N_20815);
xnor U21176 (N_21176,N_20847,N_20951);
or U21177 (N_21177,N_20891,N_20845);
and U21178 (N_21178,N_20956,N_20844);
or U21179 (N_21179,N_20852,N_20849);
nor U21180 (N_21180,N_20954,N_20960);
xor U21181 (N_21181,N_20903,N_20942);
xnor U21182 (N_21182,N_20803,N_20809);
nor U21183 (N_21183,N_20994,N_20896);
xor U21184 (N_21184,N_20849,N_20864);
xor U21185 (N_21185,N_20834,N_20939);
and U21186 (N_21186,N_20988,N_20939);
nor U21187 (N_21187,N_20932,N_20870);
and U21188 (N_21188,N_20851,N_20876);
nor U21189 (N_21189,N_20852,N_20914);
and U21190 (N_21190,N_20806,N_20835);
nor U21191 (N_21191,N_20883,N_20884);
xnor U21192 (N_21192,N_20953,N_20844);
and U21193 (N_21193,N_20938,N_20831);
nor U21194 (N_21194,N_20846,N_20874);
xor U21195 (N_21195,N_20819,N_20820);
xor U21196 (N_21196,N_20948,N_20919);
nor U21197 (N_21197,N_20839,N_20968);
nor U21198 (N_21198,N_20894,N_20864);
and U21199 (N_21199,N_20920,N_20813);
or U21200 (N_21200,N_21099,N_21052);
or U21201 (N_21201,N_21014,N_21075);
or U21202 (N_21202,N_21163,N_21124);
and U21203 (N_21203,N_21059,N_21118);
and U21204 (N_21204,N_21039,N_21072);
nor U21205 (N_21205,N_21162,N_21135);
or U21206 (N_21206,N_21154,N_21069);
nor U21207 (N_21207,N_21189,N_21047);
nand U21208 (N_21208,N_21169,N_21086);
or U21209 (N_21209,N_21087,N_21131);
and U21210 (N_21210,N_21056,N_21134);
nor U21211 (N_21211,N_21027,N_21168);
and U21212 (N_21212,N_21077,N_21031);
xor U21213 (N_21213,N_21007,N_21033);
xnor U21214 (N_21214,N_21187,N_21028);
or U21215 (N_21215,N_21080,N_21019);
or U21216 (N_21216,N_21085,N_21181);
nor U21217 (N_21217,N_21144,N_21100);
or U21218 (N_21218,N_21152,N_21005);
nor U21219 (N_21219,N_21146,N_21018);
and U21220 (N_21220,N_21138,N_21140);
xor U21221 (N_21221,N_21167,N_21042);
and U21222 (N_21222,N_21032,N_21009);
nor U21223 (N_21223,N_21058,N_21066);
xnor U21224 (N_21224,N_21136,N_21143);
nor U21225 (N_21225,N_21081,N_21120);
nand U21226 (N_21226,N_21196,N_21123);
and U21227 (N_21227,N_21068,N_21074);
nor U21228 (N_21228,N_21105,N_21002);
nand U21229 (N_21229,N_21182,N_21071);
and U21230 (N_21230,N_21037,N_21043);
nor U21231 (N_21231,N_21076,N_21096);
and U21232 (N_21232,N_21035,N_21117);
and U21233 (N_21233,N_21156,N_21186);
xor U21234 (N_21234,N_21192,N_21091);
xnor U21235 (N_21235,N_21149,N_21048);
xnor U21236 (N_21236,N_21045,N_21114);
and U21237 (N_21237,N_21015,N_21046);
and U21238 (N_21238,N_21024,N_21004);
or U21239 (N_21239,N_21142,N_21092);
nand U21240 (N_21240,N_21173,N_21020);
and U21241 (N_21241,N_21023,N_21174);
nand U21242 (N_21242,N_21041,N_21155);
nor U21243 (N_21243,N_21097,N_21010);
xnor U21244 (N_21244,N_21116,N_21171);
xnor U21245 (N_21245,N_21060,N_21049);
xnor U21246 (N_21246,N_21106,N_21057);
nand U21247 (N_21247,N_21038,N_21050);
xor U21248 (N_21248,N_21158,N_21191);
xor U21249 (N_21249,N_21176,N_21090);
or U21250 (N_21250,N_21153,N_21129);
nor U21251 (N_21251,N_21121,N_21083);
and U21252 (N_21252,N_21172,N_21065);
nand U21253 (N_21253,N_21064,N_21044);
nand U21254 (N_21254,N_21011,N_21034);
nand U21255 (N_21255,N_21185,N_21006);
nor U21256 (N_21256,N_21108,N_21070);
or U21257 (N_21257,N_21130,N_21150);
or U21258 (N_21258,N_21178,N_21054);
nor U21259 (N_21259,N_21079,N_21132);
nor U21260 (N_21260,N_21093,N_21001);
nor U21261 (N_21261,N_21062,N_21109);
nand U21262 (N_21262,N_21119,N_21040);
xnor U21263 (N_21263,N_21193,N_21113);
nor U21264 (N_21264,N_21133,N_21166);
or U21265 (N_21265,N_21095,N_21082);
xnor U21266 (N_21266,N_21107,N_21073);
xnor U21267 (N_21267,N_21110,N_21175);
nand U21268 (N_21268,N_21188,N_21084);
xnor U21269 (N_21269,N_21190,N_21003);
and U21270 (N_21270,N_21055,N_21063);
or U21271 (N_21271,N_21016,N_21127);
nor U21272 (N_21272,N_21025,N_21122);
nand U21273 (N_21273,N_21164,N_21165);
nor U21274 (N_21274,N_21115,N_21111);
nand U21275 (N_21275,N_21161,N_21000);
or U21276 (N_21276,N_21104,N_21197);
nor U21277 (N_21277,N_21184,N_21195);
nand U21278 (N_21278,N_21101,N_21053);
nand U21279 (N_21279,N_21198,N_21139);
nand U21280 (N_21280,N_21026,N_21128);
and U21281 (N_21281,N_21126,N_21179);
nand U21282 (N_21282,N_21089,N_21013);
or U21283 (N_21283,N_21008,N_21017);
and U21284 (N_21284,N_21029,N_21112);
or U21285 (N_21285,N_21177,N_21151);
xor U21286 (N_21286,N_21012,N_21180);
xor U21287 (N_21287,N_21067,N_21199);
xnor U21288 (N_21288,N_21170,N_21030);
or U21289 (N_21289,N_21088,N_21157);
nand U21290 (N_21290,N_21078,N_21137);
and U21291 (N_21291,N_21147,N_21141);
or U21292 (N_21292,N_21102,N_21021);
or U21293 (N_21293,N_21183,N_21103);
and U21294 (N_21294,N_21061,N_21194);
and U21295 (N_21295,N_21159,N_21145);
nor U21296 (N_21296,N_21094,N_21160);
nand U21297 (N_21297,N_21125,N_21098);
nand U21298 (N_21298,N_21148,N_21036);
and U21299 (N_21299,N_21051,N_21022);
and U21300 (N_21300,N_21140,N_21044);
nor U21301 (N_21301,N_21125,N_21156);
and U21302 (N_21302,N_21104,N_21051);
or U21303 (N_21303,N_21091,N_21069);
xor U21304 (N_21304,N_21017,N_21148);
and U21305 (N_21305,N_21136,N_21004);
xor U21306 (N_21306,N_21110,N_21021);
xnor U21307 (N_21307,N_21135,N_21157);
and U21308 (N_21308,N_21076,N_21190);
and U21309 (N_21309,N_21157,N_21071);
and U21310 (N_21310,N_21191,N_21018);
xnor U21311 (N_21311,N_21163,N_21031);
xor U21312 (N_21312,N_21176,N_21026);
nand U21313 (N_21313,N_21182,N_21032);
and U21314 (N_21314,N_21010,N_21105);
or U21315 (N_21315,N_21091,N_21150);
xnor U21316 (N_21316,N_21077,N_21028);
or U21317 (N_21317,N_21051,N_21031);
or U21318 (N_21318,N_21059,N_21141);
and U21319 (N_21319,N_21198,N_21019);
nor U21320 (N_21320,N_21123,N_21065);
xor U21321 (N_21321,N_21083,N_21038);
nand U21322 (N_21322,N_21197,N_21160);
nand U21323 (N_21323,N_21100,N_21125);
xnor U21324 (N_21324,N_21019,N_21028);
or U21325 (N_21325,N_21076,N_21066);
nand U21326 (N_21326,N_21103,N_21009);
xnor U21327 (N_21327,N_21166,N_21054);
xnor U21328 (N_21328,N_21146,N_21021);
and U21329 (N_21329,N_21063,N_21138);
nand U21330 (N_21330,N_21104,N_21136);
nand U21331 (N_21331,N_21005,N_21178);
xor U21332 (N_21332,N_21098,N_21105);
or U21333 (N_21333,N_21190,N_21186);
or U21334 (N_21334,N_21022,N_21017);
nand U21335 (N_21335,N_21023,N_21086);
nor U21336 (N_21336,N_21021,N_21170);
nor U21337 (N_21337,N_21194,N_21147);
xnor U21338 (N_21338,N_21119,N_21064);
and U21339 (N_21339,N_21078,N_21080);
and U21340 (N_21340,N_21156,N_21121);
xnor U21341 (N_21341,N_21126,N_21041);
or U21342 (N_21342,N_21151,N_21138);
or U21343 (N_21343,N_21117,N_21046);
and U21344 (N_21344,N_21003,N_21175);
xnor U21345 (N_21345,N_21114,N_21031);
xnor U21346 (N_21346,N_21096,N_21055);
nand U21347 (N_21347,N_21141,N_21031);
nand U21348 (N_21348,N_21021,N_21061);
xor U21349 (N_21349,N_21087,N_21042);
or U21350 (N_21350,N_21117,N_21139);
and U21351 (N_21351,N_21067,N_21020);
nor U21352 (N_21352,N_21185,N_21155);
nand U21353 (N_21353,N_21073,N_21056);
nor U21354 (N_21354,N_21104,N_21124);
xor U21355 (N_21355,N_21199,N_21037);
or U21356 (N_21356,N_21070,N_21178);
nand U21357 (N_21357,N_21025,N_21035);
or U21358 (N_21358,N_21183,N_21014);
xor U21359 (N_21359,N_21145,N_21060);
xnor U21360 (N_21360,N_21035,N_21022);
nand U21361 (N_21361,N_21096,N_21128);
or U21362 (N_21362,N_21006,N_21099);
or U21363 (N_21363,N_21061,N_21101);
nand U21364 (N_21364,N_21007,N_21073);
and U21365 (N_21365,N_21115,N_21199);
and U21366 (N_21366,N_21072,N_21109);
nor U21367 (N_21367,N_21165,N_21012);
xor U21368 (N_21368,N_21165,N_21167);
nor U21369 (N_21369,N_21000,N_21150);
or U21370 (N_21370,N_21046,N_21129);
nand U21371 (N_21371,N_21023,N_21156);
nand U21372 (N_21372,N_21178,N_21199);
nand U21373 (N_21373,N_21060,N_21173);
nor U21374 (N_21374,N_21126,N_21154);
nand U21375 (N_21375,N_21115,N_21059);
nor U21376 (N_21376,N_21067,N_21163);
nand U21377 (N_21377,N_21110,N_21167);
or U21378 (N_21378,N_21148,N_21195);
or U21379 (N_21379,N_21041,N_21198);
xor U21380 (N_21380,N_21113,N_21190);
or U21381 (N_21381,N_21155,N_21140);
and U21382 (N_21382,N_21077,N_21000);
nor U21383 (N_21383,N_21035,N_21145);
nor U21384 (N_21384,N_21182,N_21035);
xnor U21385 (N_21385,N_21143,N_21030);
xor U21386 (N_21386,N_21142,N_21195);
nand U21387 (N_21387,N_21018,N_21195);
nor U21388 (N_21388,N_21100,N_21159);
xnor U21389 (N_21389,N_21198,N_21119);
nor U21390 (N_21390,N_21048,N_21165);
or U21391 (N_21391,N_21001,N_21027);
and U21392 (N_21392,N_21121,N_21069);
xnor U21393 (N_21393,N_21045,N_21083);
nor U21394 (N_21394,N_21025,N_21026);
and U21395 (N_21395,N_21034,N_21012);
and U21396 (N_21396,N_21072,N_21013);
or U21397 (N_21397,N_21083,N_21174);
nor U21398 (N_21398,N_21188,N_21099);
and U21399 (N_21399,N_21087,N_21019);
xor U21400 (N_21400,N_21359,N_21239);
xor U21401 (N_21401,N_21294,N_21223);
and U21402 (N_21402,N_21322,N_21297);
or U21403 (N_21403,N_21323,N_21274);
nor U21404 (N_21404,N_21326,N_21316);
nor U21405 (N_21405,N_21291,N_21286);
xnor U21406 (N_21406,N_21324,N_21319);
or U21407 (N_21407,N_21310,N_21260);
xnor U21408 (N_21408,N_21343,N_21331);
and U21409 (N_21409,N_21342,N_21284);
xnor U21410 (N_21410,N_21364,N_21349);
nor U21411 (N_21411,N_21262,N_21237);
or U21412 (N_21412,N_21398,N_21219);
xnor U21413 (N_21413,N_21264,N_21336);
xnor U21414 (N_21414,N_21250,N_21351);
or U21415 (N_21415,N_21386,N_21235);
nor U21416 (N_21416,N_21287,N_21347);
or U21417 (N_21417,N_21207,N_21329);
xor U21418 (N_21418,N_21290,N_21234);
xor U21419 (N_21419,N_21301,N_21275);
and U21420 (N_21420,N_21208,N_21334);
or U21421 (N_21421,N_21354,N_21361);
nor U21422 (N_21422,N_21243,N_21345);
nand U21423 (N_21423,N_21356,N_21232);
nand U21424 (N_21424,N_21244,N_21296);
or U21425 (N_21425,N_21338,N_21302);
or U21426 (N_21426,N_21344,N_21374);
xor U21427 (N_21427,N_21367,N_21371);
or U21428 (N_21428,N_21382,N_21397);
and U21429 (N_21429,N_21267,N_21357);
xnor U21430 (N_21430,N_21391,N_21218);
xor U21431 (N_21431,N_21303,N_21355);
or U21432 (N_21432,N_21362,N_21225);
nor U21433 (N_21433,N_21229,N_21233);
or U21434 (N_21434,N_21293,N_21384);
nand U21435 (N_21435,N_21333,N_21269);
nor U21436 (N_21436,N_21236,N_21273);
and U21437 (N_21437,N_21206,N_21245);
nor U21438 (N_21438,N_21279,N_21381);
and U21439 (N_21439,N_21365,N_21392);
or U21440 (N_21440,N_21380,N_21375);
or U21441 (N_21441,N_21308,N_21315);
xor U21442 (N_21442,N_21350,N_21210);
and U21443 (N_21443,N_21231,N_21268);
nor U21444 (N_21444,N_21266,N_21212);
nand U21445 (N_21445,N_21369,N_21327);
nor U21446 (N_21446,N_21251,N_21325);
nand U21447 (N_21447,N_21304,N_21204);
and U21448 (N_21448,N_21288,N_21242);
or U21449 (N_21449,N_21320,N_21221);
and U21450 (N_21450,N_21201,N_21276);
nand U21451 (N_21451,N_21281,N_21396);
and U21452 (N_21452,N_21282,N_21230);
or U21453 (N_21453,N_21317,N_21265);
or U21454 (N_21454,N_21305,N_21314);
or U21455 (N_21455,N_21256,N_21217);
and U21456 (N_21456,N_21295,N_21348);
nand U21457 (N_21457,N_21278,N_21248);
nor U21458 (N_21458,N_21383,N_21247);
nor U21459 (N_21459,N_21203,N_21280);
nand U21460 (N_21460,N_21259,N_21258);
xor U21461 (N_21461,N_21395,N_21353);
and U21462 (N_21462,N_21241,N_21216);
or U21463 (N_21463,N_21337,N_21388);
or U21464 (N_21464,N_21246,N_21335);
nor U21465 (N_21465,N_21271,N_21332);
xnor U21466 (N_21466,N_21339,N_21283);
or U21467 (N_21467,N_21263,N_21390);
or U21468 (N_21468,N_21224,N_21311);
nor U21469 (N_21469,N_21299,N_21209);
nor U21470 (N_21470,N_21249,N_21358);
and U21471 (N_21471,N_21321,N_21289);
nor U21472 (N_21472,N_21399,N_21376);
or U21473 (N_21473,N_21378,N_21292);
and U21474 (N_21474,N_21363,N_21330);
and U21475 (N_21475,N_21270,N_21346);
or U21476 (N_21476,N_21389,N_21215);
or U21477 (N_21477,N_21385,N_21200);
nand U21478 (N_21478,N_21360,N_21387);
xnor U21479 (N_21479,N_21309,N_21222);
xor U21480 (N_21480,N_21257,N_21306);
xor U21481 (N_21481,N_21252,N_21202);
nand U21482 (N_21482,N_21366,N_21368);
nand U21483 (N_21483,N_21277,N_21272);
xor U21484 (N_21484,N_21312,N_21228);
or U21485 (N_21485,N_21341,N_21328);
xor U21486 (N_21486,N_21307,N_21313);
xor U21487 (N_21487,N_21240,N_21298);
nor U21488 (N_21488,N_21220,N_21370);
or U21489 (N_21489,N_21211,N_21372);
or U21490 (N_21490,N_21352,N_21238);
xnor U21491 (N_21491,N_21253,N_21254);
and U21492 (N_21492,N_21205,N_21213);
nand U21493 (N_21493,N_21394,N_21214);
nor U21494 (N_21494,N_21261,N_21285);
xnor U21495 (N_21495,N_21377,N_21255);
nor U21496 (N_21496,N_21227,N_21318);
and U21497 (N_21497,N_21373,N_21226);
or U21498 (N_21498,N_21300,N_21393);
or U21499 (N_21499,N_21340,N_21379);
nand U21500 (N_21500,N_21227,N_21216);
or U21501 (N_21501,N_21268,N_21225);
xnor U21502 (N_21502,N_21256,N_21303);
xor U21503 (N_21503,N_21217,N_21381);
xnor U21504 (N_21504,N_21300,N_21342);
and U21505 (N_21505,N_21353,N_21275);
and U21506 (N_21506,N_21263,N_21226);
or U21507 (N_21507,N_21297,N_21367);
nor U21508 (N_21508,N_21257,N_21280);
nand U21509 (N_21509,N_21353,N_21363);
xor U21510 (N_21510,N_21240,N_21363);
nor U21511 (N_21511,N_21356,N_21296);
nor U21512 (N_21512,N_21352,N_21280);
and U21513 (N_21513,N_21200,N_21290);
xor U21514 (N_21514,N_21347,N_21293);
or U21515 (N_21515,N_21320,N_21203);
nand U21516 (N_21516,N_21265,N_21374);
or U21517 (N_21517,N_21226,N_21274);
xor U21518 (N_21518,N_21273,N_21281);
xor U21519 (N_21519,N_21375,N_21222);
nor U21520 (N_21520,N_21379,N_21236);
xnor U21521 (N_21521,N_21342,N_21277);
nand U21522 (N_21522,N_21209,N_21335);
nor U21523 (N_21523,N_21213,N_21232);
or U21524 (N_21524,N_21346,N_21392);
nor U21525 (N_21525,N_21231,N_21347);
nor U21526 (N_21526,N_21335,N_21206);
or U21527 (N_21527,N_21220,N_21219);
or U21528 (N_21528,N_21367,N_21269);
xor U21529 (N_21529,N_21285,N_21322);
nor U21530 (N_21530,N_21331,N_21219);
xnor U21531 (N_21531,N_21275,N_21218);
xor U21532 (N_21532,N_21285,N_21246);
or U21533 (N_21533,N_21339,N_21214);
nor U21534 (N_21534,N_21384,N_21317);
nor U21535 (N_21535,N_21245,N_21368);
nand U21536 (N_21536,N_21302,N_21371);
nor U21537 (N_21537,N_21326,N_21232);
nand U21538 (N_21538,N_21341,N_21373);
or U21539 (N_21539,N_21318,N_21388);
nor U21540 (N_21540,N_21359,N_21232);
nand U21541 (N_21541,N_21288,N_21363);
or U21542 (N_21542,N_21307,N_21225);
nor U21543 (N_21543,N_21266,N_21252);
nor U21544 (N_21544,N_21220,N_21310);
nand U21545 (N_21545,N_21264,N_21315);
and U21546 (N_21546,N_21394,N_21351);
and U21547 (N_21547,N_21386,N_21337);
nand U21548 (N_21548,N_21267,N_21309);
xor U21549 (N_21549,N_21200,N_21388);
xnor U21550 (N_21550,N_21287,N_21294);
or U21551 (N_21551,N_21373,N_21241);
nand U21552 (N_21552,N_21270,N_21325);
nand U21553 (N_21553,N_21395,N_21246);
xor U21554 (N_21554,N_21237,N_21230);
or U21555 (N_21555,N_21272,N_21284);
xor U21556 (N_21556,N_21276,N_21216);
xnor U21557 (N_21557,N_21356,N_21230);
nand U21558 (N_21558,N_21238,N_21216);
nor U21559 (N_21559,N_21264,N_21321);
nand U21560 (N_21560,N_21287,N_21332);
and U21561 (N_21561,N_21243,N_21389);
and U21562 (N_21562,N_21331,N_21380);
xor U21563 (N_21563,N_21254,N_21207);
nand U21564 (N_21564,N_21206,N_21399);
nand U21565 (N_21565,N_21213,N_21323);
xor U21566 (N_21566,N_21264,N_21346);
or U21567 (N_21567,N_21384,N_21378);
and U21568 (N_21568,N_21309,N_21316);
or U21569 (N_21569,N_21238,N_21210);
or U21570 (N_21570,N_21319,N_21318);
nand U21571 (N_21571,N_21271,N_21309);
nor U21572 (N_21572,N_21201,N_21363);
or U21573 (N_21573,N_21229,N_21292);
nor U21574 (N_21574,N_21326,N_21381);
and U21575 (N_21575,N_21262,N_21204);
nor U21576 (N_21576,N_21290,N_21301);
nand U21577 (N_21577,N_21373,N_21336);
nor U21578 (N_21578,N_21323,N_21287);
or U21579 (N_21579,N_21372,N_21206);
and U21580 (N_21580,N_21317,N_21207);
nor U21581 (N_21581,N_21284,N_21202);
or U21582 (N_21582,N_21366,N_21349);
and U21583 (N_21583,N_21370,N_21338);
nor U21584 (N_21584,N_21301,N_21302);
and U21585 (N_21585,N_21299,N_21339);
and U21586 (N_21586,N_21276,N_21321);
nor U21587 (N_21587,N_21363,N_21246);
nand U21588 (N_21588,N_21213,N_21275);
or U21589 (N_21589,N_21380,N_21217);
xnor U21590 (N_21590,N_21300,N_21357);
and U21591 (N_21591,N_21253,N_21323);
nand U21592 (N_21592,N_21353,N_21206);
and U21593 (N_21593,N_21367,N_21254);
or U21594 (N_21594,N_21219,N_21276);
and U21595 (N_21595,N_21332,N_21379);
xnor U21596 (N_21596,N_21262,N_21323);
nor U21597 (N_21597,N_21231,N_21302);
and U21598 (N_21598,N_21249,N_21314);
and U21599 (N_21599,N_21259,N_21356);
nand U21600 (N_21600,N_21501,N_21549);
or U21601 (N_21601,N_21599,N_21528);
or U21602 (N_21602,N_21509,N_21593);
or U21603 (N_21603,N_21546,N_21478);
xor U21604 (N_21604,N_21558,N_21552);
nor U21605 (N_21605,N_21459,N_21580);
and U21606 (N_21606,N_21515,N_21531);
nor U21607 (N_21607,N_21581,N_21408);
or U21608 (N_21608,N_21586,N_21555);
or U21609 (N_21609,N_21468,N_21452);
xor U21610 (N_21610,N_21481,N_21411);
or U21611 (N_21611,N_21539,N_21498);
xor U21612 (N_21612,N_21484,N_21409);
and U21613 (N_21613,N_21526,N_21422);
nand U21614 (N_21614,N_21493,N_21461);
xnor U21615 (N_21615,N_21476,N_21517);
nand U21616 (N_21616,N_21569,N_21577);
and U21617 (N_21617,N_21415,N_21535);
and U21618 (N_21618,N_21458,N_21453);
or U21619 (N_21619,N_21592,N_21563);
nor U21620 (N_21620,N_21583,N_21446);
and U21621 (N_21621,N_21585,N_21502);
or U21622 (N_21622,N_21405,N_21544);
xor U21623 (N_21623,N_21406,N_21441);
and U21624 (N_21624,N_21428,N_21564);
nand U21625 (N_21625,N_21407,N_21504);
or U21626 (N_21626,N_21568,N_21485);
nor U21627 (N_21627,N_21514,N_21561);
xnor U21628 (N_21628,N_21518,N_21488);
nor U21629 (N_21629,N_21489,N_21467);
nand U21630 (N_21630,N_21447,N_21594);
nor U21631 (N_21631,N_21425,N_21503);
xor U21632 (N_21632,N_21450,N_21413);
nor U21633 (N_21633,N_21433,N_21559);
or U21634 (N_21634,N_21519,N_21404);
and U21635 (N_21635,N_21554,N_21445);
and U21636 (N_21636,N_21572,N_21466);
xnor U21637 (N_21637,N_21449,N_21551);
nor U21638 (N_21638,N_21543,N_21571);
nor U21639 (N_21639,N_21412,N_21547);
xor U21640 (N_21640,N_21508,N_21448);
or U21641 (N_21641,N_21462,N_21471);
nor U21642 (N_21642,N_21434,N_21556);
and U21643 (N_21643,N_21573,N_21578);
nor U21644 (N_21644,N_21567,N_21419);
nand U21645 (N_21645,N_21427,N_21553);
and U21646 (N_21646,N_21443,N_21465);
xor U21647 (N_21647,N_21474,N_21534);
or U21648 (N_21648,N_21472,N_21492);
nand U21649 (N_21649,N_21538,N_21523);
nor U21650 (N_21650,N_21532,N_21512);
or U21651 (N_21651,N_21588,N_21541);
nand U21652 (N_21652,N_21497,N_21426);
nand U21653 (N_21653,N_21436,N_21424);
and U21654 (N_21654,N_21432,N_21416);
nor U21655 (N_21655,N_21557,N_21494);
or U21656 (N_21656,N_21516,N_21506);
nor U21657 (N_21657,N_21527,N_21524);
nor U21658 (N_21658,N_21595,N_21429);
xnor U21659 (N_21659,N_21421,N_21482);
nand U21660 (N_21660,N_21536,N_21420);
xor U21661 (N_21661,N_21438,N_21521);
nand U21662 (N_21662,N_21469,N_21589);
nor U21663 (N_21663,N_21598,N_21520);
or U21664 (N_21664,N_21401,N_21584);
xor U21665 (N_21665,N_21486,N_21479);
or U21666 (N_21666,N_21431,N_21402);
or U21667 (N_21667,N_21490,N_21575);
xnor U21668 (N_21668,N_21525,N_21456);
and U21669 (N_21669,N_21591,N_21491);
nor U21670 (N_21670,N_21460,N_21570);
nor U21671 (N_21671,N_21545,N_21439);
nor U21672 (N_21672,N_21542,N_21487);
nand U21673 (N_21673,N_21507,N_21418);
xor U21674 (N_21674,N_21464,N_21455);
nand U21675 (N_21675,N_21513,N_21463);
and U21676 (N_21676,N_21566,N_21470);
and U21677 (N_21677,N_21403,N_21562);
nor U21678 (N_21678,N_21510,N_21499);
xnor U21679 (N_21679,N_21457,N_21410);
nand U21680 (N_21680,N_21565,N_21473);
xnor U21681 (N_21681,N_21579,N_21435);
and U21682 (N_21682,N_21511,N_21576);
nor U21683 (N_21683,N_21480,N_21582);
xor U21684 (N_21684,N_21529,N_21437);
nor U21685 (N_21685,N_21548,N_21590);
xnor U21686 (N_21686,N_21550,N_21597);
and U21687 (N_21687,N_21417,N_21587);
xor U21688 (N_21688,N_21522,N_21483);
nor U21689 (N_21689,N_21505,N_21475);
nand U21690 (N_21690,N_21596,N_21540);
or U21691 (N_21691,N_21530,N_21414);
xnor U21692 (N_21692,N_21451,N_21495);
or U21693 (N_21693,N_21423,N_21574);
or U21694 (N_21694,N_21533,N_21560);
or U21695 (N_21695,N_21496,N_21454);
nor U21696 (N_21696,N_21444,N_21500);
nand U21697 (N_21697,N_21400,N_21477);
and U21698 (N_21698,N_21430,N_21442);
nand U21699 (N_21699,N_21537,N_21440);
nand U21700 (N_21700,N_21453,N_21514);
and U21701 (N_21701,N_21435,N_21555);
or U21702 (N_21702,N_21526,N_21505);
or U21703 (N_21703,N_21428,N_21449);
nand U21704 (N_21704,N_21568,N_21439);
or U21705 (N_21705,N_21418,N_21584);
nor U21706 (N_21706,N_21431,N_21495);
xor U21707 (N_21707,N_21537,N_21445);
or U21708 (N_21708,N_21406,N_21482);
xor U21709 (N_21709,N_21470,N_21466);
and U21710 (N_21710,N_21440,N_21560);
and U21711 (N_21711,N_21596,N_21533);
nor U21712 (N_21712,N_21560,N_21484);
nand U21713 (N_21713,N_21531,N_21417);
nand U21714 (N_21714,N_21401,N_21471);
and U21715 (N_21715,N_21574,N_21587);
or U21716 (N_21716,N_21512,N_21534);
and U21717 (N_21717,N_21571,N_21485);
or U21718 (N_21718,N_21411,N_21531);
nor U21719 (N_21719,N_21478,N_21583);
nand U21720 (N_21720,N_21408,N_21403);
xor U21721 (N_21721,N_21565,N_21583);
nand U21722 (N_21722,N_21560,N_21566);
nor U21723 (N_21723,N_21415,N_21412);
nor U21724 (N_21724,N_21544,N_21441);
xnor U21725 (N_21725,N_21444,N_21562);
nor U21726 (N_21726,N_21519,N_21528);
nand U21727 (N_21727,N_21484,N_21598);
and U21728 (N_21728,N_21516,N_21502);
or U21729 (N_21729,N_21567,N_21512);
nand U21730 (N_21730,N_21478,N_21505);
or U21731 (N_21731,N_21563,N_21536);
or U21732 (N_21732,N_21575,N_21460);
nand U21733 (N_21733,N_21498,N_21492);
nand U21734 (N_21734,N_21452,N_21430);
nor U21735 (N_21735,N_21472,N_21414);
xnor U21736 (N_21736,N_21476,N_21496);
xor U21737 (N_21737,N_21561,N_21474);
and U21738 (N_21738,N_21565,N_21529);
nor U21739 (N_21739,N_21431,N_21518);
nand U21740 (N_21740,N_21515,N_21574);
or U21741 (N_21741,N_21553,N_21446);
xor U21742 (N_21742,N_21479,N_21590);
xnor U21743 (N_21743,N_21577,N_21537);
or U21744 (N_21744,N_21489,N_21455);
xor U21745 (N_21745,N_21584,N_21597);
xnor U21746 (N_21746,N_21430,N_21594);
xnor U21747 (N_21747,N_21480,N_21427);
xor U21748 (N_21748,N_21463,N_21487);
or U21749 (N_21749,N_21403,N_21514);
and U21750 (N_21750,N_21534,N_21553);
nand U21751 (N_21751,N_21469,N_21548);
nand U21752 (N_21752,N_21427,N_21450);
and U21753 (N_21753,N_21554,N_21411);
nor U21754 (N_21754,N_21476,N_21539);
xor U21755 (N_21755,N_21402,N_21526);
nand U21756 (N_21756,N_21483,N_21529);
or U21757 (N_21757,N_21599,N_21503);
or U21758 (N_21758,N_21455,N_21545);
nor U21759 (N_21759,N_21462,N_21461);
or U21760 (N_21760,N_21412,N_21404);
or U21761 (N_21761,N_21585,N_21419);
and U21762 (N_21762,N_21424,N_21563);
xor U21763 (N_21763,N_21513,N_21586);
xor U21764 (N_21764,N_21454,N_21422);
xor U21765 (N_21765,N_21471,N_21444);
xor U21766 (N_21766,N_21511,N_21463);
xnor U21767 (N_21767,N_21448,N_21521);
nor U21768 (N_21768,N_21434,N_21421);
or U21769 (N_21769,N_21457,N_21502);
xnor U21770 (N_21770,N_21453,N_21497);
nor U21771 (N_21771,N_21500,N_21475);
nor U21772 (N_21772,N_21519,N_21590);
and U21773 (N_21773,N_21446,N_21434);
or U21774 (N_21774,N_21436,N_21496);
or U21775 (N_21775,N_21407,N_21441);
nor U21776 (N_21776,N_21586,N_21454);
nand U21777 (N_21777,N_21529,N_21469);
and U21778 (N_21778,N_21471,N_21438);
nand U21779 (N_21779,N_21574,N_21421);
xor U21780 (N_21780,N_21423,N_21538);
nand U21781 (N_21781,N_21532,N_21498);
and U21782 (N_21782,N_21534,N_21459);
and U21783 (N_21783,N_21409,N_21522);
nor U21784 (N_21784,N_21512,N_21578);
nor U21785 (N_21785,N_21523,N_21479);
nand U21786 (N_21786,N_21444,N_21567);
nor U21787 (N_21787,N_21483,N_21519);
or U21788 (N_21788,N_21400,N_21568);
nor U21789 (N_21789,N_21468,N_21436);
nand U21790 (N_21790,N_21583,N_21572);
or U21791 (N_21791,N_21525,N_21513);
nor U21792 (N_21792,N_21572,N_21458);
nand U21793 (N_21793,N_21483,N_21552);
or U21794 (N_21794,N_21481,N_21489);
nand U21795 (N_21795,N_21508,N_21480);
nor U21796 (N_21796,N_21542,N_21536);
nor U21797 (N_21797,N_21556,N_21544);
nand U21798 (N_21798,N_21486,N_21582);
xnor U21799 (N_21799,N_21464,N_21552);
or U21800 (N_21800,N_21647,N_21747);
nor U21801 (N_21801,N_21646,N_21761);
and U21802 (N_21802,N_21645,N_21752);
or U21803 (N_21803,N_21795,N_21797);
and U21804 (N_21804,N_21730,N_21739);
and U21805 (N_21805,N_21634,N_21733);
xor U21806 (N_21806,N_21756,N_21608);
nand U21807 (N_21807,N_21695,N_21769);
xnor U21808 (N_21808,N_21628,N_21703);
or U21809 (N_21809,N_21709,N_21686);
nand U21810 (N_21810,N_21796,N_21746);
nor U21811 (N_21811,N_21794,N_21727);
nand U21812 (N_21812,N_21673,N_21741);
and U21813 (N_21813,N_21728,N_21786);
and U21814 (N_21814,N_21731,N_21701);
and U21815 (N_21815,N_21788,N_21722);
xor U21816 (N_21816,N_21720,N_21658);
or U21817 (N_21817,N_21687,N_21783);
xor U21818 (N_21818,N_21631,N_21714);
or U21819 (N_21819,N_21775,N_21780);
and U21820 (N_21820,N_21784,N_21662);
xor U21821 (N_21821,N_21721,N_21663);
or U21822 (N_21822,N_21632,N_21724);
or U21823 (N_21823,N_21671,N_21688);
or U21824 (N_21824,N_21653,N_21770);
xnor U21825 (N_21825,N_21649,N_21787);
or U21826 (N_21826,N_21716,N_21755);
nand U21827 (N_21827,N_21782,N_21738);
or U21828 (N_21828,N_21754,N_21681);
or U21829 (N_21829,N_21707,N_21633);
nand U21830 (N_21830,N_21615,N_21619);
nor U21831 (N_21831,N_21705,N_21702);
nand U21832 (N_21832,N_21719,N_21602);
nand U21833 (N_21833,N_21723,N_21699);
xor U21834 (N_21834,N_21708,N_21768);
or U21835 (N_21835,N_21610,N_21640);
nand U21836 (N_21836,N_21715,N_21630);
nand U21837 (N_21837,N_21762,N_21771);
xor U21838 (N_21838,N_21680,N_21604);
nor U21839 (N_21839,N_21665,N_21789);
and U21840 (N_21840,N_21698,N_21607);
xnor U21841 (N_21841,N_21678,N_21791);
xnor U21842 (N_21842,N_21601,N_21657);
nand U21843 (N_21843,N_21676,N_21736);
xnor U21844 (N_21844,N_21612,N_21776);
nand U21845 (N_21845,N_21605,N_21641);
and U21846 (N_21846,N_21690,N_21758);
or U21847 (N_21847,N_21790,N_21675);
nand U21848 (N_21848,N_21618,N_21664);
xor U21849 (N_21849,N_21700,N_21660);
nor U21850 (N_21850,N_21611,N_21737);
nor U21851 (N_21851,N_21627,N_21749);
nor U21852 (N_21852,N_21751,N_21651);
and U21853 (N_21853,N_21704,N_21620);
xor U21854 (N_21854,N_21718,N_21774);
xor U21855 (N_21855,N_21717,N_21757);
or U21856 (N_21856,N_21767,N_21742);
and U21857 (N_21857,N_21793,N_21696);
nor U21858 (N_21858,N_21711,N_21625);
nand U21859 (N_21859,N_21669,N_21799);
and U21860 (N_21860,N_21765,N_21666);
and U21861 (N_21861,N_21743,N_21694);
xor U21862 (N_21862,N_21679,N_21760);
or U21863 (N_21863,N_21614,N_21689);
nor U21864 (N_21864,N_21637,N_21603);
or U21865 (N_21865,N_21668,N_21781);
nor U21866 (N_21866,N_21750,N_21763);
or U21867 (N_21867,N_21744,N_21652);
nor U21868 (N_21868,N_21622,N_21643);
and U21869 (N_21869,N_21753,N_21785);
nand U21870 (N_21870,N_21644,N_21616);
nand U21871 (N_21871,N_21609,N_21745);
or U21872 (N_21872,N_21732,N_21621);
nor U21873 (N_21873,N_21642,N_21685);
and U21874 (N_21874,N_21638,N_21617);
or U21875 (N_21875,N_21655,N_21667);
xnor U21876 (N_21876,N_21764,N_21735);
xor U21877 (N_21877,N_21697,N_21624);
and U21878 (N_21878,N_21682,N_21623);
nor U21879 (N_21879,N_21629,N_21777);
xor U21880 (N_21880,N_21674,N_21773);
nand U21881 (N_21881,N_21691,N_21659);
and U21882 (N_21882,N_21613,N_21759);
nand U21883 (N_21883,N_21778,N_21713);
and U21884 (N_21884,N_21729,N_21626);
or U21885 (N_21885,N_21710,N_21670);
or U21886 (N_21886,N_21684,N_21636);
nand U21887 (N_21887,N_21656,N_21672);
nor U21888 (N_21888,N_21654,N_21772);
and U21889 (N_21889,N_21766,N_21748);
or U21890 (N_21890,N_21734,N_21648);
nor U21891 (N_21891,N_21692,N_21650);
or U21892 (N_21892,N_21712,N_21725);
xor U21893 (N_21893,N_21677,N_21606);
and U21894 (N_21894,N_21779,N_21600);
and U21895 (N_21895,N_21661,N_21683);
or U21896 (N_21896,N_21706,N_21798);
nor U21897 (N_21897,N_21635,N_21639);
or U21898 (N_21898,N_21726,N_21740);
or U21899 (N_21899,N_21792,N_21693);
or U21900 (N_21900,N_21611,N_21628);
or U21901 (N_21901,N_21743,N_21622);
xnor U21902 (N_21902,N_21731,N_21672);
and U21903 (N_21903,N_21756,N_21674);
and U21904 (N_21904,N_21649,N_21756);
nor U21905 (N_21905,N_21749,N_21780);
or U21906 (N_21906,N_21604,N_21694);
nor U21907 (N_21907,N_21713,N_21680);
and U21908 (N_21908,N_21619,N_21784);
nor U21909 (N_21909,N_21708,N_21733);
xor U21910 (N_21910,N_21631,N_21720);
xor U21911 (N_21911,N_21682,N_21635);
or U21912 (N_21912,N_21600,N_21634);
nor U21913 (N_21913,N_21708,N_21748);
nand U21914 (N_21914,N_21624,N_21754);
and U21915 (N_21915,N_21732,N_21600);
and U21916 (N_21916,N_21625,N_21756);
nand U21917 (N_21917,N_21673,N_21639);
or U21918 (N_21918,N_21776,N_21796);
nand U21919 (N_21919,N_21752,N_21735);
nor U21920 (N_21920,N_21606,N_21655);
or U21921 (N_21921,N_21690,N_21699);
nor U21922 (N_21922,N_21726,N_21692);
nand U21923 (N_21923,N_21640,N_21791);
and U21924 (N_21924,N_21605,N_21710);
and U21925 (N_21925,N_21767,N_21782);
or U21926 (N_21926,N_21716,N_21702);
or U21927 (N_21927,N_21674,N_21601);
nor U21928 (N_21928,N_21633,N_21731);
and U21929 (N_21929,N_21748,N_21676);
and U21930 (N_21930,N_21715,N_21635);
xor U21931 (N_21931,N_21775,N_21650);
xnor U21932 (N_21932,N_21752,N_21664);
nand U21933 (N_21933,N_21624,N_21610);
or U21934 (N_21934,N_21708,N_21605);
nor U21935 (N_21935,N_21666,N_21688);
xor U21936 (N_21936,N_21767,N_21796);
nor U21937 (N_21937,N_21769,N_21629);
and U21938 (N_21938,N_21673,N_21695);
nand U21939 (N_21939,N_21764,N_21609);
or U21940 (N_21940,N_21751,N_21646);
or U21941 (N_21941,N_21795,N_21752);
or U21942 (N_21942,N_21757,N_21744);
nor U21943 (N_21943,N_21728,N_21677);
nand U21944 (N_21944,N_21724,N_21662);
nand U21945 (N_21945,N_21609,N_21630);
and U21946 (N_21946,N_21719,N_21683);
nand U21947 (N_21947,N_21673,N_21603);
xnor U21948 (N_21948,N_21725,N_21726);
and U21949 (N_21949,N_21682,N_21738);
xnor U21950 (N_21950,N_21703,N_21675);
and U21951 (N_21951,N_21697,N_21759);
or U21952 (N_21952,N_21699,N_21641);
nand U21953 (N_21953,N_21684,N_21767);
nand U21954 (N_21954,N_21794,N_21635);
nand U21955 (N_21955,N_21627,N_21799);
and U21956 (N_21956,N_21792,N_21779);
nor U21957 (N_21957,N_21658,N_21662);
xor U21958 (N_21958,N_21672,N_21755);
nor U21959 (N_21959,N_21632,N_21722);
nand U21960 (N_21960,N_21729,N_21790);
nor U21961 (N_21961,N_21703,N_21612);
nand U21962 (N_21962,N_21695,N_21706);
or U21963 (N_21963,N_21729,N_21619);
or U21964 (N_21964,N_21799,N_21780);
nor U21965 (N_21965,N_21676,N_21630);
xor U21966 (N_21966,N_21752,N_21689);
or U21967 (N_21967,N_21689,N_21793);
nand U21968 (N_21968,N_21666,N_21776);
nand U21969 (N_21969,N_21719,N_21619);
nand U21970 (N_21970,N_21649,N_21702);
nand U21971 (N_21971,N_21711,N_21758);
nor U21972 (N_21972,N_21793,N_21618);
nand U21973 (N_21973,N_21652,N_21784);
nand U21974 (N_21974,N_21796,N_21785);
nor U21975 (N_21975,N_21705,N_21614);
and U21976 (N_21976,N_21713,N_21748);
xnor U21977 (N_21977,N_21727,N_21737);
xnor U21978 (N_21978,N_21698,N_21707);
xor U21979 (N_21979,N_21726,N_21733);
nand U21980 (N_21980,N_21782,N_21652);
nor U21981 (N_21981,N_21672,N_21602);
xnor U21982 (N_21982,N_21779,N_21643);
nand U21983 (N_21983,N_21625,N_21712);
nand U21984 (N_21984,N_21676,N_21750);
or U21985 (N_21985,N_21634,N_21788);
nand U21986 (N_21986,N_21778,N_21772);
or U21987 (N_21987,N_21728,N_21602);
nand U21988 (N_21988,N_21690,N_21730);
or U21989 (N_21989,N_21602,N_21663);
or U21990 (N_21990,N_21745,N_21771);
xnor U21991 (N_21991,N_21637,N_21723);
or U21992 (N_21992,N_21684,N_21707);
or U21993 (N_21993,N_21715,N_21749);
nor U21994 (N_21994,N_21752,N_21694);
and U21995 (N_21995,N_21793,N_21628);
and U21996 (N_21996,N_21619,N_21735);
and U21997 (N_21997,N_21796,N_21798);
nand U21998 (N_21998,N_21736,N_21609);
nor U21999 (N_21999,N_21679,N_21766);
nand U22000 (N_22000,N_21847,N_21881);
xnor U22001 (N_22001,N_21914,N_21833);
nor U22002 (N_22002,N_21893,N_21868);
xnor U22003 (N_22003,N_21863,N_21848);
or U22004 (N_22004,N_21979,N_21811);
nor U22005 (N_22005,N_21807,N_21846);
nand U22006 (N_22006,N_21996,N_21928);
and U22007 (N_22007,N_21830,N_21882);
or U22008 (N_22008,N_21982,N_21972);
nand U22009 (N_22009,N_21934,N_21887);
xor U22010 (N_22010,N_21852,N_21944);
nor U22011 (N_22011,N_21925,N_21859);
nand U22012 (N_22012,N_21907,N_21800);
xor U22013 (N_22013,N_21947,N_21990);
and U22014 (N_22014,N_21946,N_21898);
nand U22015 (N_22015,N_21809,N_21929);
nand U22016 (N_22016,N_21957,N_21879);
nor U22017 (N_22017,N_21858,N_21921);
and U22018 (N_22018,N_21981,N_21999);
nor U22019 (N_22019,N_21955,N_21909);
or U22020 (N_22020,N_21867,N_21853);
nor U22021 (N_22021,N_21937,N_21936);
and U22022 (N_22022,N_21978,N_21949);
xor U22023 (N_22023,N_21823,N_21903);
and U22024 (N_22024,N_21857,N_21959);
xor U22025 (N_22025,N_21930,N_21884);
nand U22026 (N_22026,N_21886,N_21839);
xor U22027 (N_22027,N_21860,N_21980);
nand U22028 (N_22028,N_21910,N_21954);
or U22029 (N_22029,N_21973,N_21942);
or U22030 (N_22030,N_21916,N_21922);
nand U22031 (N_22031,N_21950,N_21904);
xnor U22032 (N_22032,N_21984,N_21943);
nor U22033 (N_22033,N_21965,N_21827);
xor U22034 (N_22034,N_21961,N_21968);
xnor U22035 (N_22035,N_21939,N_21831);
nor U22036 (N_22036,N_21828,N_21824);
or U22037 (N_22037,N_21902,N_21854);
or U22038 (N_22038,N_21986,N_21834);
or U22039 (N_22039,N_21927,N_21808);
or U22040 (N_22040,N_21829,N_21964);
nor U22041 (N_22041,N_21871,N_21892);
nor U22042 (N_22042,N_21977,N_21804);
nand U22043 (N_22043,N_21997,N_21931);
nand U22044 (N_22044,N_21958,N_21851);
or U22045 (N_22045,N_21865,N_21819);
nand U22046 (N_22046,N_21872,N_21969);
nor U22047 (N_22047,N_21926,N_21919);
or U22048 (N_22048,N_21880,N_21912);
xnor U22049 (N_22049,N_21814,N_21935);
and U22050 (N_22050,N_21825,N_21995);
xnor U22051 (N_22051,N_21953,N_21988);
or U22052 (N_22052,N_21805,N_21917);
or U22053 (N_22053,N_21835,N_21971);
xnor U22054 (N_22054,N_21822,N_21813);
and U22055 (N_22055,N_21841,N_21960);
or U22056 (N_22056,N_21956,N_21861);
and U22057 (N_22057,N_21876,N_21842);
xnor U22058 (N_22058,N_21963,N_21985);
nor U22059 (N_22059,N_21966,N_21856);
or U22060 (N_22060,N_21818,N_21976);
xor U22061 (N_22061,N_21802,N_21821);
or U22062 (N_22062,N_21883,N_21975);
xor U22063 (N_22063,N_21803,N_21970);
nand U22064 (N_22064,N_21952,N_21889);
nor U22065 (N_22065,N_21915,N_21998);
or U22066 (N_22066,N_21820,N_21945);
and U22067 (N_22067,N_21941,N_21895);
or U22068 (N_22068,N_21890,N_21913);
nor U22069 (N_22069,N_21962,N_21844);
xor U22070 (N_22070,N_21816,N_21836);
nand U22071 (N_22071,N_21874,N_21845);
nor U22072 (N_22072,N_21908,N_21924);
and U22073 (N_22073,N_21983,N_21850);
nand U22074 (N_22074,N_21905,N_21897);
nor U22075 (N_22075,N_21992,N_21901);
nor U22076 (N_22076,N_21869,N_21838);
or U22077 (N_22077,N_21801,N_21948);
and U22078 (N_22078,N_21900,N_21810);
xor U22079 (N_22079,N_21843,N_21967);
nand U22080 (N_22080,N_21837,N_21993);
or U22081 (N_22081,N_21826,N_21987);
xnor U22082 (N_22082,N_21873,N_21877);
and U22083 (N_22083,N_21875,N_21920);
nand U22084 (N_22084,N_21864,N_21866);
xnor U22085 (N_22085,N_21911,N_21906);
and U22086 (N_22086,N_21974,N_21991);
and U22087 (N_22087,N_21994,N_21923);
and U22088 (N_22088,N_21891,N_21855);
nand U22089 (N_22089,N_21878,N_21870);
nand U22090 (N_22090,N_21817,N_21989);
and U22091 (N_22091,N_21849,N_21815);
or U22092 (N_22092,N_21951,N_21888);
nor U22093 (N_22093,N_21812,N_21806);
and U22094 (N_22094,N_21885,N_21862);
or U22095 (N_22095,N_21896,N_21918);
xnor U22096 (N_22096,N_21933,N_21832);
xnor U22097 (N_22097,N_21940,N_21840);
xor U22098 (N_22098,N_21899,N_21932);
xor U22099 (N_22099,N_21894,N_21938);
nor U22100 (N_22100,N_21902,N_21960);
and U22101 (N_22101,N_21928,N_21802);
and U22102 (N_22102,N_21860,N_21861);
xnor U22103 (N_22103,N_21828,N_21983);
xor U22104 (N_22104,N_21957,N_21815);
or U22105 (N_22105,N_21996,N_21926);
and U22106 (N_22106,N_21813,N_21850);
nand U22107 (N_22107,N_21810,N_21847);
nand U22108 (N_22108,N_21954,N_21850);
and U22109 (N_22109,N_21899,N_21911);
nor U22110 (N_22110,N_21823,N_21891);
nor U22111 (N_22111,N_21926,N_21900);
xnor U22112 (N_22112,N_21895,N_21956);
or U22113 (N_22113,N_21965,N_21841);
and U22114 (N_22114,N_21925,N_21834);
nand U22115 (N_22115,N_21881,N_21834);
xor U22116 (N_22116,N_21802,N_21920);
xnor U22117 (N_22117,N_21819,N_21950);
or U22118 (N_22118,N_21819,N_21915);
nor U22119 (N_22119,N_21829,N_21958);
nand U22120 (N_22120,N_21828,N_21873);
or U22121 (N_22121,N_21878,N_21897);
xnor U22122 (N_22122,N_21831,N_21982);
nand U22123 (N_22123,N_21815,N_21934);
nand U22124 (N_22124,N_21952,N_21876);
nor U22125 (N_22125,N_21841,N_21823);
xor U22126 (N_22126,N_21942,N_21843);
nor U22127 (N_22127,N_21814,N_21893);
or U22128 (N_22128,N_21870,N_21892);
nand U22129 (N_22129,N_21907,N_21815);
xor U22130 (N_22130,N_21969,N_21831);
and U22131 (N_22131,N_21862,N_21824);
nand U22132 (N_22132,N_21910,N_21884);
nand U22133 (N_22133,N_21984,N_21940);
nand U22134 (N_22134,N_21906,N_21876);
and U22135 (N_22135,N_21820,N_21955);
or U22136 (N_22136,N_21912,N_21860);
nor U22137 (N_22137,N_21947,N_21924);
and U22138 (N_22138,N_21834,N_21960);
xnor U22139 (N_22139,N_21888,N_21883);
xor U22140 (N_22140,N_21924,N_21951);
and U22141 (N_22141,N_21842,N_21903);
or U22142 (N_22142,N_21957,N_21929);
nor U22143 (N_22143,N_21992,N_21844);
and U22144 (N_22144,N_21830,N_21980);
nand U22145 (N_22145,N_21981,N_21820);
nor U22146 (N_22146,N_21924,N_21882);
and U22147 (N_22147,N_21945,N_21827);
or U22148 (N_22148,N_21975,N_21933);
nor U22149 (N_22149,N_21865,N_21873);
or U22150 (N_22150,N_21902,N_21930);
nand U22151 (N_22151,N_21869,N_21922);
and U22152 (N_22152,N_21992,N_21885);
and U22153 (N_22153,N_21979,N_21885);
xor U22154 (N_22154,N_21870,N_21985);
nand U22155 (N_22155,N_21903,N_21817);
nand U22156 (N_22156,N_21883,N_21915);
or U22157 (N_22157,N_21851,N_21965);
nand U22158 (N_22158,N_21815,N_21806);
nand U22159 (N_22159,N_21811,N_21886);
xor U22160 (N_22160,N_21918,N_21817);
or U22161 (N_22161,N_21904,N_21898);
nor U22162 (N_22162,N_21955,N_21842);
xnor U22163 (N_22163,N_21941,N_21945);
nand U22164 (N_22164,N_21872,N_21828);
xor U22165 (N_22165,N_21987,N_21903);
or U22166 (N_22166,N_21902,N_21954);
xnor U22167 (N_22167,N_21944,N_21878);
xor U22168 (N_22168,N_21939,N_21943);
xor U22169 (N_22169,N_21967,N_21934);
xnor U22170 (N_22170,N_21843,N_21917);
or U22171 (N_22171,N_21888,N_21842);
nor U22172 (N_22172,N_21850,N_21827);
or U22173 (N_22173,N_21905,N_21873);
or U22174 (N_22174,N_21841,N_21969);
xnor U22175 (N_22175,N_21913,N_21955);
xor U22176 (N_22176,N_21951,N_21862);
nand U22177 (N_22177,N_21865,N_21985);
nor U22178 (N_22178,N_21827,N_21860);
xnor U22179 (N_22179,N_21956,N_21965);
or U22180 (N_22180,N_21889,N_21947);
or U22181 (N_22181,N_21877,N_21939);
nand U22182 (N_22182,N_21945,N_21865);
xor U22183 (N_22183,N_21946,N_21892);
nor U22184 (N_22184,N_21866,N_21848);
and U22185 (N_22185,N_21806,N_21878);
or U22186 (N_22186,N_21806,N_21804);
nand U22187 (N_22187,N_21848,N_21895);
and U22188 (N_22188,N_21978,N_21800);
and U22189 (N_22189,N_21930,N_21963);
or U22190 (N_22190,N_21942,N_21844);
or U22191 (N_22191,N_21957,N_21994);
and U22192 (N_22192,N_21996,N_21895);
nand U22193 (N_22193,N_21805,N_21816);
and U22194 (N_22194,N_21926,N_21885);
or U22195 (N_22195,N_21960,N_21952);
and U22196 (N_22196,N_21915,N_21807);
xor U22197 (N_22197,N_21915,N_21972);
nand U22198 (N_22198,N_21842,N_21994);
xnor U22199 (N_22199,N_21878,N_21968);
xnor U22200 (N_22200,N_22165,N_22138);
nor U22201 (N_22201,N_22155,N_22146);
xor U22202 (N_22202,N_22015,N_22090);
and U22203 (N_22203,N_22132,N_22083);
nor U22204 (N_22204,N_22164,N_22075);
or U22205 (N_22205,N_22187,N_22175);
nor U22206 (N_22206,N_22074,N_22169);
or U22207 (N_22207,N_22183,N_22121);
nor U22208 (N_22208,N_22048,N_22031);
nor U22209 (N_22209,N_22013,N_22006);
and U22210 (N_22210,N_22193,N_22087);
or U22211 (N_22211,N_22098,N_22058);
and U22212 (N_22212,N_22039,N_22148);
nor U22213 (N_22213,N_22078,N_22152);
nor U22214 (N_22214,N_22136,N_22184);
and U22215 (N_22215,N_22178,N_22143);
xnor U22216 (N_22216,N_22077,N_22159);
nand U22217 (N_22217,N_22023,N_22072);
and U22218 (N_22218,N_22174,N_22195);
nor U22219 (N_22219,N_22021,N_22004);
and U22220 (N_22220,N_22158,N_22151);
xor U22221 (N_22221,N_22162,N_22047);
or U22222 (N_22222,N_22060,N_22067);
and U22223 (N_22223,N_22166,N_22191);
nor U22224 (N_22224,N_22197,N_22129);
nand U22225 (N_22225,N_22007,N_22186);
nor U22226 (N_22226,N_22046,N_22001);
xor U22227 (N_22227,N_22092,N_22068);
and U22228 (N_22228,N_22055,N_22161);
nand U22229 (N_22229,N_22038,N_22099);
nor U22230 (N_22230,N_22107,N_22194);
xnor U22231 (N_22231,N_22070,N_22199);
or U22232 (N_22232,N_22168,N_22125);
xor U22233 (N_22233,N_22163,N_22156);
nand U22234 (N_22234,N_22120,N_22127);
nand U22235 (N_22235,N_22190,N_22056);
nor U22236 (N_22236,N_22073,N_22118);
xor U22237 (N_22237,N_22035,N_22106);
nand U22238 (N_22238,N_22097,N_22003);
or U22239 (N_22239,N_22008,N_22140);
nor U22240 (N_22240,N_22139,N_22160);
and U22241 (N_22241,N_22086,N_22185);
xnor U22242 (N_22242,N_22126,N_22034);
or U22243 (N_22243,N_22010,N_22064);
xor U22244 (N_22244,N_22094,N_22116);
nand U22245 (N_22245,N_22167,N_22011);
or U22246 (N_22246,N_22032,N_22182);
and U22247 (N_22247,N_22045,N_22128);
or U22248 (N_22248,N_22084,N_22153);
nand U22249 (N_22249,N_22000,N_22133);
and U22250 (N_22250,N_22192,N_22157);
nor U22251 (N_22251,N_22171,N_22022);
nor U22252 (N_22252,N_22054,N_22154);
xnor U22253 (N_22253,N_22012,N_22131);
and U22254 (N_22254,N_22044,N_22170);
or U22255 (N_22255,N_22014,N_22113);
or U22256 (N_22256,N_22123,N_22181);
or U22257 (N_22257,N_22081,N_22069);
nor U22258 (N_22258,N_22111,N_22108);
or U22259 (N_22259,N_22062,N_22063);
and U22260 (N_22260,N_22082,N_22196);
xor U22261 (N_22261,N_22122,N_22052);
and U22262 (N_22262,N_22176,N_22076);
and U22263 (N_22263,N_22095,N_22189);
nand U22264 (N_22264,N_22017,N_22173);
or U22265 (N_22265,N_22061,N_22080);
and U22266 (N_22266,N_22104,N_22109);
or U22267 (N_22267,N_22110,N_22049);
or U22268 (N_22268,N_22117,N_22089);
nor U22269 (N_22269,N_22124,N_22030);
and U22270 (N_22270,N_22042,N_22043);
and U22271 (N_22271,N_22188,N_22144);
nand U22272 (N_22272,N_22147,N_22112);
nor U22273 (N_22273,N_22066,N_22149);
nor U22274 (N_22274,N_22020,N_22051);
or U22275 (N_22275,N_22145,N_22150);
nor U22276 (N_22276,N_22103,N_22025);
and U22277 (N_22277,N_22028,N_22096);
or U22278 (N_22278,N_22130,N_22088);
nand U22279 (N_22279,N_22180,N_22085);
or U22280 (N_22280,N_22179,N_22101);
xor U22281 (N_22281,N_22050,N_22102);
and U22282 (N_22282,N_22105,N_22134);
and U22283 (N_22283,N_22177,N_22009);
or U22284 (N_22284,N_22093,N_22141);
xor U22285 (N_22285,N_22065,N_22019);
nor U22286 (N_22286,N_22115,N_22040);
nor U22287 (N_22287,N_22024,N_22059);
or U22288 (N_22288,N_22027,N_22142);
or U22289 (N_22289,N_22137,N_22033);
nand U22290 (N_22290,N_22198,N_22114);
and U22291 (N_22291,N_22005,N_22071);
and U22292 (N_22292,N_22057,N_22036);
or U22293 (N_22293,N_22002,N_22041);
xor U22294 (N_22294,N_22079,N_22172);
and U22295 (N_22295,N_22029,N_22091);
xnor U22296 (N_22296,N_22018,N_22119);
nor U22297 (N_22297,N_22016,N_22135);
nand U22298 (N_22298,N_22026,N_22037);
and U22299 (N_22299,N_22053,N_22100);
and U22300 (N_22300,N_22079,N_22176);
or U22301 (N_22301,N_22057,N_22103);
nand U22302 (N_22302,N_22030,N_22040);
xor U22303 (N_22303,N_22058,N_22150);
or U22304 (N_22304,N_22011,N_22111);
xnor U22305 (N_22305,N_22071,N_22089);
or U22306 (N_22306,N_22086,N_22118);
nor U22307 (N_22307,N_22084,N_22068);
and U22308 (N_22308,N_22051,N_22162);
and U22309 (N_22309,N_22061,N_22113);
and U22310 (N_22310,N_22055,N_22051);
nand U22311 (N_22311,N_22163,N_22060);
nand U22312 (N_22312,N_22021,N_22115);
and U22313 (N_22313,N_22084,N_22025);
and U22314 (N_22314,N_22117,N_22056);
xor U22315 (N_22315,N_22068,N_22061);
xor U22316 (N_22316,N_22121,N_22084);
nand U22317 (N_22317,N_22071,N_22153);
xor U22318 (N_22318,N_22059,N_22180);
nor U22319 (N_22319,N_22164,N_22156);
and U22320 (N_22320,N_22031,N_22156);
or U22321 (N_22321,N_22077,N_22052);
and U22322 (N_22322,N_22173,N_22074);
nand U22323 (N_22323,N_22191,N_22028);
and U22324 (N_22324,N_22182,N_22110);
nand U22325 (N_22325,N_22095,N_22012);
nor U22326 (N_22326,N_22145,N_22164);
nand U22327 (N_22327,N_22194,N_22183);
and U22328 (N_22328,N_22027,N_22177);
or U22329 (N_22329,N_22123,N_22083);
xor U22330 (N_22330,N_22111,N_22105);
xor U22331 (N_22331,N_22196,N_22012);
xor U22332 (N_22332,N_22107,N_22104);
nand U22333 (N_22333,N_22066,N_22159);
nor U22334 (N_22334,N_22196,N_22002);
xor U22335 (N_22335,N_22151,N_22155);
xnor U22336 (N_22336,N_22174,N_22151);
xnor U22337 (N_22337,N_22176,N_22050);
xor U22338 (N_22338,N_22011,N_22191);
nor U22339 (N_22339,N_22195,N_22015);
nor U22340 (N_22340,N_22114,N_22075);
nor U22341 (N_22341,N_22188,N_22137);
xor U22342 (N_22342,N_22011,N_22120);
nor U22343 (N_22343,N_22093,N_22054);
nor U22344 (N_22344,N_22006,N_22176);
and U22345 (N_22345,N_22197,N_22101);
and U22346 (N_22346,N_22113,N_22196);
nor U22347 (N_22347,N_22020,N_22021);
or U22348 (N_22348,N_22077,N_22061);
or U22349 (N_22349,N_22087,N_22137);
xor U22350 (N_22350,N_22005,N_22174);
nand U22351 (N_22351,N_22012,N_22073);
xnor U22352 (N_22352,N_22185,N_22015);
and U22353 (N_22353,N_22135,N_22021);
xnor U22354 (N_22354,N_22182,N_22122);
xor U22355 (N_22355,N_22054,N_22077);
nor U22356 (N_22356,N_22008,N_22090);
or U22357 (N_22357,N_22080,N_22172);
and U22358 (N_22358,N_22096,N_22002);
nor U22359 (N_22359,N_22090,N_22161);
or U22360 (N_22360,N_22031,N_22012);
and U22361 (N_22361,N_22128,N_22198);
and U22362 (N_22362,N_22097,N_22161);
nor U22363 (N_22363,N_22189,N_22187);
nand U22364 (N_22364,N_22161,N_22171);
and U22365 (N_22365,N_22055,N_22062);
or U22366 (N_22366,N_22065,N_22057);
and U22367 (N_22367,N_22168,N_22066);
xor U22368 (N_22368,N_22084,N_22058);
nand U22369 (N_22369,N_22027,N_22161);
xnor U22370 (N_22370,N_22050,N_22124);
xor U22371 (N_22371,N_22092,N_22102);
nor U22372 (N_22372,N_22035,N_22198);
and U22373 (N_22373,N_22082,N_22135);
and U22374 (N_22374,N_22040,N_22116);
nor U22375 (N_22375,N_22129,N_22176);
and U22376 (N_22376,N_22111,N_22072);
nand U22377 (N_22377,N_22111,N_22121);
and U22378 (N_22378,N_22154,N_22179);
nand U22379 (N_22379,N_22114,N_22140);
or U22380 (N_22380,N_22167,N_22153);
and U22381 (N_22381,N_22115,N_22172);
nand U22382 (N_22382,N_22087,N_22066);
xnor U22383 (N_22383,N_22040,N_22166);
nand U22384 (N_22384,N_22116,N_22056);
and U22385 (N_22385,N_22177,N_22173);
nand U22386 (N_22386,N_22012,N_22177);
or U22387 (N_22387,N_22151,N_22048);
or U22388 (N_22388,N_22073,N_22127);
nand U22389 (N_22389,N_22033,N_22153);
nand U22390 (N_22390,N_22116,N_22156);
nand U22391 (N_22391,N_22022,N_22156);
and U22392 (N_22392,N_22098,N_22136);
xnor U22393 (N_22393,N_22136,N_22137);
nor U22394 (N_22394,N_22165,N_22082);
and U22395 (N_22395,N_22003,N_22049);
and U22396 (N_22396,N_22040,N_22180);
and U22397 (N_22397,N_22101,N_22057);
or U22398 (N_22398,N_22138,N_22105);
nor U22399 (N_22399,N_22144,N_22146);
xnor U22400 (N_22400,N_22250,N_22217);
and U22401 (N_22401,N_22335,N_22321);
nor U22402 (N_22402,N_22366,N_22351);
nand U22403 (N_22403,N_22326,N_22299);
xor U22404 (N_22404,N_22337,N_22387);
or U22405 (N_22405,N_22369,N_22291);
xor U22406 (N_22406,N_22228,N_22333);
nor U22407 (N_22407,N_22345,N_22232);
nor U22408 (N_22408,N_22203,N_22370);
nor U22409 (N_22409,N_22302,N_22378);
and U22410 (N_22410,N_22239,N_22263);
and U22411 (N_22411,N_22295,N_22312);
nor U22412 (N_22412,N_22289,N_22319);
nor U22413 (N_22413,N_22244,N_22390);
or U22414 (N_22414,N_22286,N_22292);
nand U22415 (N_22415,N_22393,N_22355);
nand U22416 (N_22416,N_22243,N_22394);
nand U22417 (N_22417,N_22363,N_22329);
nand U22418 (N_22418,N_22210,N_22266);
nand U22419 (N_22419,N_22222,N_22285);
nand U22420 (N_22420,N_22377,N_22349);
nor U22421 (N_22421,N_22373,N_22270);
xor U22422 (N_22422,N_22208,N_22313);
nor U22423 (N_22423,N_22259,N_22296);
nand U22424 (N_22424,N_22356,N_22354);
and U22425 (N_22425,N_22332,N_22261);
or U22426 (N_22426,N_22267,N_22275);
and U22427 (N_22427,N_22247,N_22290);
nor U22428 (N_22428,N_22281,N_22288);
or U22429 (N_22429,N_22361,N_22308);
nor U22430 (N_22430,N_22223,N_22236);
and U22431 (N_22431,N_22200,N_22323);
nand U22432 (N_22432,N_22316,N_22242);
nand U22433 (N_22433,N_22371,N_22209);
xor U22434 (N_22434,N_22279,N_22314);
nor U22435 (N_22435,N_22317,N_22277);
xor U22436 (N_22436,N_22330,N_22318);
and U22437 (N_22437,N_22205,N_22320);
nor U22438 (N_22438,N_22287,N_22297);
nor U22439 (N_22439,N_22305,N_22220);
nand U22440 (N_22440,N_22358,N_22395);
nor U22441 (N_22441,N_22241,N_22328);
or U22442 (N_22442,N_22338,N_22280);
or U22443 (N_22443,N_22231,N_22327);
or U22444 (N_22444,N_22265,N_22331);
and U22445 (N_22445,N_22233,N_22353);
xnor U22446 (N_22446,N_22360,N_22283);
xor U22447 (N_22447,N_22230,N_22201);
nand U22448 (N_22448,N_22396,N_22229);
xor U22449 (N_22449,N_22399,N_22324);
and U22450 (N_22450,N_22379,N_22234);
and U22451 (N_22451,N_22310,N_22264);
nand U22452 (N_22452,N_22334,N_22352);
xor U22453 (N_22453,N_22315,N_22274);
and U22454 (N_22454,N_22359,N_22284);
xnor U22455 (N_22455,N_22254,N_22375);
nand U22456 (N_22456,N_22212,N_22364);
xor U22457 (N_22457,N_22347,N_22282);
xnor U22458 (N_22458,N_22322,N_22300);
xnor U22459 (N_22459,N_22252,N_22336);
xor U22460 (N_22460,N_22248,N_22372);
nor U22461 (N_22461,N_22268,N_22202);
nor U22462 (N_22462,N_22238,N_22346);
nor U22463 (N_22463,N_22348,N_22255);
or U22464 (N_22464,N_22376,N_22213);
nor U22465 (N_22465,N_22388,N_22381);
nand U22466 (N_22466,N_22342,N_22340);
and U22467 (N_22467,N_22391,N_22272);
or U22468 (N_22468,N_22204,N_22207);
nor U22469 (N_22469,N_22276,N_22219);
nand U22470 (N_22470,N_22251,N_22341);
or U22471 (N_22471,N_22386,N_22211);
and U22472 (N_22472,N_22218,N_22380);
or U22473 (N_22473,N_22397,N_22258);
nor U22474 (N_22474,N_22214,N_22307);
and U22475 (N_22475,N_22385,N_22398);
and U22476 (N_22476,N_22294,N_22293);
and U22477 (N_22477,N_22384,N_22367);
nor U22478 (N_22478,N_22368,N_22389);
and U22479 (N_22479,N_22271,N_22225);
nand U22480 (N_22480,N_22235,N_22227);
nor U22481 (N_22481,N_22256,N_22237);
or U22482 (N_22482,N_22216,N_22221);
xor U22483 (N_22483,N_22339,N_22374);
xnor U22484 (N_22484,N_22245,N_22226);
nor U22485 (N_22485,N_22269,N_22249);
and U22486 (N_22486,N_22382,N_22253);
nand U22487 (N_22487,N_22257,N_22240);
nand U22488 (N_22488,N_22273,N_22215);
xor U22489 (N_22489,N_22304,N_22383);
or U22490 (N_22490,N_22311,N_22325);
nor U22491 (N_22491,N_22344,N_22306);
nor U22492 (N_22492,N_22362,N_22303);
or U22493 (N_22493,N_22224,N_22260);
nand U22494 (N_22494,N_22343,N_22262);
xor U22495 (N_22495,N_22301,N_22246);
and U22496 (N_22496,N_22309,N_22357);
nand U22497 (N_22497,N_22350,N_22278);
nor U22498 (N_22498,N_22392,N_22365);
nor U22499 (N_22499,N_22206,N_22298);
and U22500 (N_22500,N_22213,N_22373);
nor U22501 (N_22501,N_22330,N_22341);
nor U22502 (N_22502,N_22385,N_22233);
nor U22503 (N_22503,N_22361,N_22380);
nand U22504 (N_22504,N_22291,N_22359);
or U22505 (N_22505,N_22394,N_22336);
xnor U22506 (N_22506,N_22239,N_22236);
xnor U22507 (N_22507,N_22315,N_22311);
nand U22508 (N_22508,N_22344,N_22334);
and U22509 (N_22509,N_22211,N_22379);
or U22510 (N_22510,N_22295,N_22224);
and U22511 (N_22511,N_22260,N_22315);
xor U22512 (N_22512,N_22214,N_22312);
or U22513 (N_22513,N_22282,N_22247);
and U22514 (N_22514,N_22318,N_22361);
nor U22515 (N_22515,N_22301,N_22304);
nor U22516 (N_22516,N_22213,N_22352);
and U22517 (N_22517,N_22236,N_22300);
or U22518 (N_22518,N_22206,N_22337);
xor U22519 (N_22519,N_22356,N_22319);
nor U22520 (N_22520,N_22316,N_22344);
nor U22521 (N_22521,N_22280,N_22322);
or U22522 (N_22522,N_22219,N_22314);
and U22523 (N_22523,N_22281,N_22383);
nor U22524 (N_22524,N_22306,N_22202);
and U22525 (N_22525,N_22308,N_22250);
xnor U22526 (N_22526,N_22320,N_22389);
or U22527 (N_22527,N_22395,N_22262);
and U22528 (N_22528,N_22312,N_22377);
or U22529 (N_22529,N_22252,N_22357);
nor U22530 (N_22530,N_22228,N_22331);
and U22531 (N_22531,N_22291,N_22238);
xor U22532 (N_22532,N_22360,N_22397);
xnor U22533 (N_22533,N_22324,N_22276);
nor U22534 (N_22534,N_22232,N_22375);
nor U22535 (N_22535,N_22215,N_22299);
xor U22536 (N_22536,N_22342,N_22337);
or U22537 (N_22537,N_22372,N_22241);
xnor U22538 (N_22538,N_22217,N_22334);
or U22539 (N_22539,N_22268,N_22369);
or U22540 (N_22540,N_22263,N_22381);
nand U22541 (N_22541,N_22210,N_22294);
and U22542 (N_22542,N_22296,N_22237);
nand U22543 (N_22543,N_22342,N_22308);
or U22544 (N_22544,N_22399,N_22248);
xnor U22545 (N_22545,N_22297,N_22249);
nor U22546 (N_22546,N_22306,N_22339);
and U22547 (N_22547,N_22217,N_22252);
xor U22548 (N_22548,N_22329,N_22241);
xor U22549 (N_22549,N_22267,N_22310);
nand U22550 (N_22550,N_22259,N_22363);
xor U22551 (N_22551,N_22304,N_22303);
nor U22552 (N_22552,N_22375,N_22255);
xnor U22553 (N_22553,N_22328,N_22317);
and U22554 (N_22554,N_22223,N_22246);
and U22555 (N_22555,N_22376,N_22391);
and U22556 (N_22556,N_22227,N_22390);
or U22557 (N_22557,N_22353,N_22363);
and U22558 (N_22558,N_22324,N_22233);
nand U22559 (N_22559,N_22240,N_22336);
nor U22560 (N_22560,N_22382,N_22290);
and U22561 (N_22561,N_22200,N_22201);
xnor U22562 (N_22562,N_22285,N_22331);
and U22563 (N_22563,N_22366,N_22314);
nand U22564 (N_22564,N_22239,N_22379);
nor U22565 (N_22565,N_22210,N_22327);
and U22566 (N_22566,N_22363,N_22304);
or U22567 (N_22567,N_22294,N_22211);
xor U22568 (N_22568,N_22240,N_22273);
xor U22569 (N_22569,N_22390,N_22349);
and U22570 (N_22570,N_22359,N_22242);
and U22571 (N_22571,N_22330,N_22219);
and U22572 (N_22572,N_22238,N_22280);
nor U22573 (N_22573,N_22287,N_22255);
or U22574 (N_22574,N_22265,N_22269);
and U22575 (N_22575,N_22346,N_22374);
or U22576 (N_22576,N_22324,N_22204);
nand U22577 (N_22577,N_22358,N_22222);
nor U22578 (N_22578,N_22246,N_22298);
nor U22579 (N_22579,N_22272,N_22289);
xor U22580 (N_22580,N_22327,N_22249);
nor U22581 (N_22581,N_22328,N_22298);
and U22582 (N_22582,N_22253,N_22377);
or U22583 (N_22583,N_22258,N_22317);
nand U22584 (N_22584,N_22264,N_22341);
nand U22585 (N_22585,N_22354,N_22392);
xnor U22586 (N_22586,N_22292,N_22348);
and U22587 (N_22587,N_22213,N_22311);
and U22588 (N_22588,N_22255,N_22225);
xnor U22589 (N_22589,N_22381,N_22261);
nand U22590 (N_22590,N_22295,N_22327);
or U22591 (N_22591,N_22343,N_22384);
nor U22592 (N_22592,N_22341,N_22222);
or U22593 (N_22593,N_22261,N_22372);
or U22594 (N_22594,N_22377,N_22317);
xor U22595 (N_22595,N_22339,N_22261);
nand U22596 (N_22596,N_22258,N_22340);
and U22597 (N_22597,N_22357,N_22274);
nand U22598 (N_22598,N_22373,N_22399);
or U22599 (N_22599,N_22322,N_22370);
nor U22600 (N_22600,N_22475,N_22587);
or U22601 (N_22601,N_22535,N_22466);
and U22602 (N_22602,N_22448,N_22510);
and U22603 (N_22603,N_22492,N_22480);
nor U22604 (N_22604,N_22572,N_22486);
and U22605 (N_22605,N_22549,N_22477);
and U22606 (N_22606,N_22490,N_22457);
and U22607 (N_22607,N_22515,N_22482);
nand U22608 (N_22608,N_22481,N_22425);
xor U22609 (N_22609,N_22459,N_22487);
xor U22610 (N_22610,N_22576,N_22547);
or U22611 (N_22611,N_22520,N_22589);
nor U22612 (N_22612,N_22539,N_22526);
nand U22613 (N_22613,N_22570,N_22546);
nand U22614 (N_22614,N_22584,N_22578);
nor U22615 (N_22615,N_22430,N_22553);
or U22616 (N_22616,N_22527,N_22493);
xnor U22617 (N_22617,N_22577,N_22417);
and U22618 (N_22618,N_22479,N_22519);
xnor U22619 (N_22619,N_22403,N_22593);
nor U22620 (N_22620,N_22504,N_22424);
and U22621 (N_22621,N_22531,N_22597);
nand U22622 (N_22622,N_22582,N_22462);
nand U22623 (N_22623,N_22488,N_22502);
nor U22624 (N_22624,N_22543,N_22423);
nor U22625 (N_22625,N_22561,N_22567);
nor U22626 (N_22626,N_22558,N_22580);
xor U22627 (N_22627,N_22507,N_22565);
nor U22628 (N_22628,N_22552,N_22569);
nor U22629 (N_22629,N_22590,N_22418);
xnor U22630 (N_22630,N_22452,N_22544);
or U22631 (N_22631,N_22536,N_22518);
nor U22632 (N_22632,N_22516,N_22574);
nand U22633 (N_22633,N_22464,N_22528);
nand U22634 (N_22634,N_22420,N_22505);
xnor U22635 (N_22635,N_22460,N_22551);
xnor U22636 (N_22636,N_22440,N_22461);
xnor U22637 (N_22637,N_22598,N_22472);
or U22638 (N_22638,N_22406,N_22412);
and U22639 (N_22639,N_22564,N_22595);
nand U22640 (N_22640,N_22554,N_22451);
xor U22641 (N_22641,N_22579,N_22489);
xor U22642 (N_22642,N_22433,N_22450);
xnor U22643 (N_22643,N_22407,N_22533);
or U22644 (N_22644,N_22458,N_22436);
or U22645 (N_22645,N_22498,N_22434);
or U22646 (N_22646,N_22538,N_22508);
and U22647 (N_22647,N_22563,N_22524);
and U22648 (N_22648,N_22503,N_22427);
and U22649 (N_22649,N_22401,N_22410);
nor U22650 (N_22650,N_22556,N_22494);
nor U22651 (N_22651,N_22497,N_22550);
nor U22652 (N_22652,N_22559,N_22513);
nand U22653 (N_22653,N_22573,N_22537);
nand U22654 (N_22654,N_22548,N_22426);
and U22655 (N_22655,N_22557,N_22444);
nand U22656 (N_22656,N_22517,N_22512);
and U22657 (N_22657,N_22596,N_22439);
nand U22658 (N_22658,N_22408,N_22435);
xnor U22659 (N_22659,N_22514,N_22575);
or U22660 (N_22660,N_22560,N_22530);
nor U22661 (N_22661,N_22453,N_22529);
or U22662 (N_22662,N_22432,N_22588);
or U22663 (N_22663,N_22441,N_22455);
xor U22664 (N_22664,N_22586,N_22419);
xor U22665 (N_22665,N_22416,N_22499);
nand U22666 (N_22666,N_22483,N_22454);
xor U22667 (N_22667,N_22467,N_22534);
and U22668 (N_22668,N_22447,N_22468);
nand U22669 (N_22669,N_22496,N_22471);
or U22670 (N_22670,N_22591,N_22465);
xor U22671 (N_22671,N_22540,N_22449);
nand U22672 (N_22672,N_22456,N_22525);
or U22673 (N_22673,N_22583,N_22562);
nor U22674 (N_22674,N_22443,N_22405);
and U22675 (N_22675,N_22506,N_22421);
and U22676 (N_22676,N_22463,N_22555);
and U22677 (N_22677,N_22500,N_22568);
or U22678 (N_22678,N_22415,N_22437);
and U22679 (N_22679,N_22592,N_22523);
xnor U22680 (N_22680,N_22571,N_22409);
xor U22681 (N_22681,N_22522,N_22478);
or U22682 (N_22682,N_22542,N_22495);
and U22683 (N_22683,N_22446,N_22402);
and U22684 (N_22684,N_22469,N_22541);
or U22685 (N_22685,N_22581,N_22511);
and U22686 (N_22686,N_22429,N_22599);
nand U22687 (N_22687,N_22470,N_22473);
and U22688 (N_22688,N_22438,N_22445);
xor U22689 (N_22689,N_22491,N_22521);
xor U22690 (N_22690,N_22431,N_22400);
or U22691 (N_22691,N_22476,N_22594);
nor U22692 (N_22692,N_22411,N_22509);
and U22693 (N_22693,N_22413,N_22566);
xor U22694 (N_22694,N_22532,N_22585);
xnor U22695 (N_22695,N_22422,N_22484);
nand U22696 (N_22696,N_22474,N_22404);
nor U22697 (N_22697,N_22414,N_22545);
or U22698 (N_22698,N_22501,N_22442);
or U22699 (N_22699,N_22485,N_22428);
and U22700 (N_22700,N_22494,N_22459);
or U22701 (N_22701,N_22494,N_22425);
nand U22702 (N_22702,N_22517,N_22545);
xor U22703 (N_22703,N_22527,N_22432);
or U22704 (N_22704,N_22570,N_22444);
and U22705 (N_22705,N_22482,N_22427);
nor U22706 (N_22706,N_22552,N_22526);
or U22707 (N_22707,N_22465,N_22403);
xor U22708 (N_22708,N_22490,N_22473);
or U22709 (N_22709,N_22586,N_22507);
nand U22710 (N_22710,N_22490,N_22417);
xor U22711 (N_22711,N_22557,N_22569);
nand U22712 (N_22712,N_22467,N_22457);
nor U22713 (N_22713,N_22465,N_22516);
xor U22714 (N_22714,N_22537,N_22440);
xnor U22715 (N_22715,N_22444,N_22493);
and U22716 (N_22716,N_22430,N_22547);
and U22717 (N_22717,N_22552,N_22486);
xor U22718 (N_22718,N_22420,N_22421);
and U22719 (N_22719,N_22491,N_22599);
nand U22720 (N_22720,N_22558,N_22569);
nand U22721 (N_22721,N_22415,N_22594);
and U22722 (N_22722,N_22439,N_22475);
xnor U22723 (N_22723,N_22493,N_22430);
xor U22724 (N_22724,N_22518,N_22567);
xor U22725 (N_22725,N_22460,N_22468);
nor U22726 (N_22726,N_22573,N_22549);
or U22727 (N_22727,N_22495,N_22512);
nand U22728 (N_22728,N_22558,N_22551);
and U22729 (N_22729,N_22511,N_22448);
nand U22730 (N_22730,N_22567,N_22448);
nand U22731 (N_22731,N_22570,N_22514);
and U22732 (N_22732,N_22511,N_22431);
nand U22733 (N_22733,N_22404,N_22468);
and U22734 (N_22734,N_22490,N_22500);
xor U22735 (N_22735,N_22551,N_22419);
nand U22736 (N_22736,N_22550,N_22433);
or U22737 (N_22737,N_22563,N_22458);
xor U22738 (N_22738,N_22565,N_22511);
nor U22739 (N_22739,N_22597,N_22581);
nand U22740 (N_22740,N_22463,N_22585);
and U22741 (N_22741,N_22439,N_22567);
nor U22742 (N_22742,N_22423,N_22527);
nand U22743 (N_22743,N_22404,N_22425);
nand U22744 (N_22744,N_22573,N_22429);
nor U22745 (N_22745,N_22513,N_22534);
or U22746 (N_22746,N_22495,N_22455);
or U22747 (N_22747,N_22508,N_22440);
xnor U22748 (N_22748,N_22489,N_22478);
or U22749 (N_22749,N_22525,N_22441);
and U22750 (N_22750,N_22470,N_22560);
nand U22751 (N_22751,N_22591,N_22485);
or U22752 (N_22752,N_22411,N_22409);
nand U22753 (N_22753,N_22523,N_22563);
or U22754 (N_22754,N_22539,N_22404);
nor U22755 (N_22755,N_22436,N_22563);
nor U22756 (N_22756,N_22417,N_22465);
xnor U22757 (N_22757,N_22565,N_22587);
nor U22758 (N_22758,N_22411,N_22590);
xor U22759 (N_22759,N_22525,N_22410);
xnor U22760 (N_22760,N_22561,N_22438);
nor U22761 (N_22761,N_22587,N_22503);
nand U22762 (N_22762,N_22543,N_22500);
nor U22763 (N_22763,N_22471,N_22552);
xor U22764 (N_22764,N_22539,N_22430);
nand U22765 (N_22765,N_22433,N_22583);
or U22766 (N_22766,N_22426,N_22445);
xnor U22767 (N_22767,N_22406,N_22545);
xnor U22768 (N_22768,N_22438,N_22588);
or U22769 (N_22769,N_22552,N_22470);
and U22770 (N_22770,N_22411,N_22498);
nor U22771 (N_22771,N_22510,N_22503);
or U22772 (N_22772,N_22462,N_22496);
nor U22773 (N_22773,N_22481,N_22488);
xor U22774 (N_22774,N_22400,N_22574);
nand U22775 (N_22775,N_22507,N_22464);
nand U22776 (N_22776,N_22499,N_22430);
xnor U22777 (N_22777,N_22521,N_22462);
nor U22778 (N_22778,N_22400,N_22498);
nand U22779 (N_22779,N_22410,N_22481);
or U22780 (N_22780,N_22418,N_22484);
nand U22781 (N_22781,N_22585,N_22435);
or U22782 (N_22782,N_22476,N_22550);
or U22783 (N_22783,N_22434,N_22407);
nand U22784 (N_22784,N_22448,N_22542);
xnor U22785 (N_22785,N_22578,N_22432);
or U22786 (N_22786,N_22553,N_22528);
nor U22787 (N_22787,N_22592,N_22423);
xor U22788 (N_22788,N_22475,N_22433);
xnor U22789 (N_22789,N_22450,N_22425);
and U22790 (N_22790,N_22593,N_22590);
nand U22791 (N_22791,N_22583,N_22559);
and U22792 (N_22792,N_22419,N_22550);
or U22793 (N_22793,N_22520,N_22582);
and U22794 (N_22794,N_22555,N_22534);
nand U22795 (N_22795,N_22466,N_22465);
xor U22796 (N_22796,N_22447,N_22503);
xor U22797 (N_22797,N_22450,N_22544);
nor U22798 (N_22798,N_22544,N_22465);
or U22799 (N_22799,N_22435,N_22509);
and U22800 (N_22800,N_22604,N_22780);
nor U22801 (N_22801,N_22669,N_22625);
or U22802 (N_22802,N_22690,N_22697);
or U22803 (N_22803,N_22768,N_22742);
xor U22804 (N_22804,N_22785,N_22783);
nand U22805 (N_22805,N_22643,N_22608);
nand U22806 (N_22806,N_22670,N_22776);
or U22807 (N_22807,N_22781,N_22752);
or U22808 (N_22808,N_22760,N_22751);
and U22809 (N_22809,N_22714,N_22661);
and U22810 (N_22810,N_22764,N_22758);
nor U22811 (N_22811,N_22660,N_22700);
xnor U22812 (N_22812,N_22685,N_22729);
or U22813 (N_22813,N_22737,N_22652);
nor U22814 (N_22814,N_22671,N_22735);
xor U22815 (N_22815,N_22716,N_22610);
xor U22816 (N_22816,N_22719,N_22732);
and U22817 (N_22817,N_22644,N_22646);
or U22818 (N_22818,N_22702,N_22756);
and U22819 (N_22819,N_22762,N_22637);
nand U22820 (N_22820,N_22635,N_22754);
and U22821 (N_22821,N_22656,N_22723);
and U22822 (N_22822,N_22706,N_22793);
nand U22823 (N_22823,N_22789,N_22773);
and U22824 (N_22824,N_22639,N_22713);
and U22825 (N_22825,N_22779,N_22761);
nand U22826 (N_22826,N_22653,N_22666);
xnor U22827 (N_22827,N_22708,N_22667);
xnor U22828 (N_22828,N_22607,N_22641);
nor U22829 (N_22829,N_22694,N_22745);
nor U22830 (N_22830,N_22633,N_22617);
nor U22831 (N_22831,N_22634,N_22741);
nor U22832 (N_22832,N_22788,N_22611);
nor U22833 (N_22833,N_22744,N_22774);
nand U22834 (N_22834,N_22695,N_22722);
and U22835 (N_22835,N_22665,N_22740);
and U22836 (N_22836,N_22620,N_22645);
nand U22837 (N_22837,N_22693,N_22632);
nand U22838 (N_22838,N_22790,N_22736);
nor U22839 (N_22839,N_22703,N_22746);
and U22840 (N_22840,N_22794,N_22724);
or U22841 (N_22841,N_22630,N_22629);
nor U22842 (N_22842,N_22682,N_22734);
xor U22843 (N_22843,N_22738,N_22672);
and U22844 (N_22844,N_22763,N_22622);
or U22845 (N_22845,N_22782,N_22609);
nor U22846 (N_22846,N_22698,N_22613);
xnor U22847 (N_22847,N_22709,N_22640);
nor U22848 (N_22848,N_22638,N_22749);
xor U22849 (N_22849,N_22750,N_22771);
nor U22850 (N_22850,N_22733,N_22691);
nor U22851 (N_22851,N_22648,N_22727);
nand U22852 (N_22852,N_22692,N_22636);
and U22853 (N_22853,N_22720,N_22678);
or U22854 (N_22854,N_22730,N_22747);
nand U22855 (N_22855,N_22712,N_22605);
and U22856 (N_22856,N_22799,N_22679);
and U22857 (N_22857,N_22705,N_22673);
or U22858 (N_22858,N_22658,N_22718);
nand U22859 (N_22859,N_22792,N_22663);
nand U22860 (N_22860,N_22784,N_22657);
nor U22861 (N_22861,N_22798,N_22715);
nand U22862 (N_22862,N_22753,N_22618);
nand U22863 (N_22863,N_22649,N_22787);
or U22864 (N_22864,N_22623,N_22786);
nand U22865 (N_22865,N_22707,N_22796);
or U22866 (N_22866,N_22726,N_22757);
or U22867 (N_22867,N_22626,N_22676);
xnor U22868 (N_22868,N_22739,N_22759);
and U22869 (N_22869,N_22721,N_22675);
or U22870 (N_22870,N_22683,N_22674);
nor U22871 (N_22871,N_22680,N_22662);
or U22872 (N_22872,N_22704,N_22664);
and U22873 (N_22873,N_22606,N_22769);
xor U22874 (N_22874,N_22795,N_22686);
nor U22875 (N_22875,N_22654,N_22767);
or U22876 (N_22876,N_22602,N_22710);
nand U22877 (N_22877,N_22668,N_22621);
and U22878 (N_22878,N_22684,N_22701);
xor U22879 (N_22879,N_22687,N_22755);
or U22880 (N_22880,N_22743,N_22650);
or U22881 (N_22881,N_22728,N_22797);
and U22882 (N_22882,N_22689,N_22603);
nor U22883 (N_22883,N_22659,N_22647);
nor U22884 (N_22884,N_22642,N_22711);
xnor U22885 (N_22885,N_22677,N_22778);
nor U22886 (N_22886,N_22696,N_22624);
and U22887 (N_22887,N_22600,N_22601);
nor U22888 (N_22888,N_22688,N_22765);
xnor U22889 (N_22889,N_22699,N_22651);
or U22890 (N_22890,N_22627,N_22717);
xor U22891 (N_22891,N_22791,N_22614);
nand U22892 (N_22892,N_22731,N_22628);
nand U22893 (N_22893,N_22615,N_22770);
nand U22894 (N_22894,N_22612,N_22777);
or U22895 (N_22895,N_22619,N_22766);
or U22896 (N_22896,N_22616,N_22748);
and U22897 (N_22897,N_22631,N_22725);
nand U22898 (N_22898,N_22772,N_22655);
nand U22899 (N_22899,N_22681,N_22775);
xor U22900 (N_22900,N_22781,N_22763);
or U22901 (N_22901,N_22605,N_22742);
and U22902 (N_22902,N_22637,N_22776);
xnor U22903 (N_22903,N_22714,N_22755);
or U22904 (N_22904,N_22774,N_22717);
nand U22905 (N_22905,N_22724,N_22795);
or U22906 (N_22906,N_22769,N_22683);
and U22907 (N_22907,N_22776,N_22686);
and U22908 (N_22908,N_22624,N_22758);
nor U22909 (N_22909,N_22784,N_22637);
or U22910 (N_22910,N_22693,N_22778);
or U22911 (N_22911,N_22770,N_22711);
nor U22912 (N_22912,N_22771,N_22773);
xnor U22913 (N_22913,N_22646,N_22677);
or U22914 (N_22914,N_22632,N_22736);
nor U22915 (N_22915,N_22763,N_22700);
nor U22916 (N_22916,N_22657,N_22630);
nor U22917 (N_22917,N_22692,N_22664);
and U22918 (N_22918,N_22638,N_22690);
nand U22919 (N_22919,N_22674,N_22684);
and U22920 (N_22920,N_22733,N_22674);
xor U22921 (N_22921,N_22709,N_22658);
nor U22922 (N_22922,N_22765,N_22606);
xor U22923 (N_22923,N_22676,N_22621);
and U22924 (N_22924,N_22799,N_22703);
or U22925 (N_22925,N_22671,N_22623);
and U22926 (N_22926,N_22741,N_22666);
and U22927 (N_22927,N_22651,N_22747);
or U22928 (N_22928,N_22636,N_22710);
and U22929 (N_22929,N_22784,N_22672);
or U22930 (N_22930,N_22714,N_22659);
and U22931 (N_22931,N_22698,N_22610);
or U22932 (N_22932,N_22651,N_22620);
or U22933 (N_22933,N_22735,N_22607);
or U22934 (N_22934,N_22745,N_22686);
xnor U22935 (N_22935,N_22688,N_22615);
xor U22936 (N_22936,N_22693,N_22674);
or U22937 (N_22937,N_22611,N_22791);
xor U22938 (N_22938,N_22653,N_22691);
nand U22939 (N_22939,N_22609,N_22664);
xnor U22940 (N_22940,N_22748,N_22621);
xnor U22941 (N_22941,N_22647,N_22741);
xnor U22942 (N_22942,N_22662,N_22636);
and U22943 (N_22943,N_22718,N_22653);
nand U22944 (N_22944,N_22715,N_22649);
nand U22945 (N_22945,N_22746,N_22752);
nor U22946 (N_22946,N_22665,N_22750);
or U22947 (N_22947,N_22692,N_22698);
or U22948 (N_22948,N_22670,N_22783);
and U22949 (N_22949,N_22673,N_22719);
or U22950 (N_22950,N_22645,N_22758);
and U22951 (N_22951,N_22681,N_22707);
xor U22952 (N_22952,N_22661,N_22651);
xnor U22953 (N_22953,N_22798,N_22752);
nand U22954 (N_22954,N_22685,N_22633);
and U22955 (N_22955,N_22721,N_22681);
and U22956 (N_22956,N_22681,N_22630);
nand U22957 (N_22957,N_22705,N_22768);
or U22958 (N_22958,N_22741,N_22658);
and U22959 (N_22959,N_22679,N_22610);
nand U22960 (N_22960,N_22646,N_22658);
nor U22961 (N_22961,N_22649,N_22747);
nor U22962 (N_22962,N_22793,N_22652);
nor U22963 (N_22963,N_22717,N_22639);
nor U22964 (N_22964,N_22720,N_22610);
nand U22965 (N_22965,N_22667,N_22716);
nand U22966 (N_22966,N_22713,N_22683);
nand U22967 (N_22967,N_22785,N_22727);
or U22968 (N_22968,N_22643,N_22691);
xor U22969 (N_22969,N_22701,N_22628);
xnor U22970 (N_22970,N_22757,N_22656);
or U22971 (N_22971,N_22635,N_22692);
and U22972 (N_22972,N_22783,N_22715);
or U22973 (N_22973,N_22635,N_22601);
nand U22974 (N_22974,N_22722,N_22693);
xnor U22975 (N_22975,N_22765,N_22748);
nand U22976 (N_22976,N_22739,N_22619);
xor U22977 (N_22977,N_22715,N_22601);
xor U22978 (N_22978,N_22769,N_22608);
nor U22979 (N_22979,N_22666,N_22637);
or U22980 (N_22980,N_22606,N_22601);
and U22981 (N_22981,N_22730,N_22676);
and U22982 (N_22982,N_22795,N_22629);
xor U22983 (N_22983,N_22782,N_22671);
nand U22984 (N_22984,N_22685,N_22643);
xor U22985 (N_22985,N_22710,N_22609);
nor U22986 (N_22986,N_22781,N_22797);
xnor U22987 (N_22987,N_22624,N_22617);
or U22988 (N_22988,N_22636,N_22708);
nor U22989 (N_22989,N_22700,N_22635);
xnor U22990 (N_22990,N_22624,N_22658);
xor U22991 (N_22991,N_22626,N_22679);
and U22992 (N_22992,N_22734,N_22640);
xnor U22993 (N_22993,N_22679,N_22752);
xnor U22994 (N_22994,N_22780,N_22749);
nor U22995 (N_22995,N_22715,N_22664);
xor U22996 (N_22996,N_22791,N_22695);
nor U22997 (N_22997,N_22602,N_22768);
nand U22998 (N_22998,N_22791,N_22657);
nor U22999 (N_22999,N_22737,N_22661);
or U23000 (N_23000,N_22858,N_22986);
nand U23001 (N_23001,N_22808,N_22874);
nor U23002 (N_23002,N_22895,N_22893);
xor U23003 (N_23003,N_22914,N_22849);
nand U23004 (N_23004,N_22825,N_22953);
nor U23005 (N_23005,N_22976,N_22964);
nand U23006 (N_23006,N_22800,N_22834);
nor U23007 (N_23007,N_22872,N_22896);
and U23008 (N_23008,N_22870,N_22868);
or U23009 (N_23009,N_22859,N_22853);
xnor U23010 (N_23010,N_22862,N_22939);
or U23011 (N_23011,N_22987,N_22933);
and U23012 (N_23012,N_22810,N_22889);
nor U23013 (N_23013,N_22966,N_22906);
or U23014 (N_23014,N_22928,N_22931);
nand U23015 (N_23015,N_22856,N_22865);
and U23016 (N_23016,N_22832,N_22887);
or U23017 (N_23017,N_22821,N_22924);
and U23018 (N_23018,N_22911,N_22845);
and U23019 (N_23019,N_22912,N_22861);
and U23020 (N_23020,N_22881,N_22851);
xor U23021 (N_23021,N_22999,N_22902);
and U23022 (N_23022,N_22869,N_22850);
nand U23023 (N_23023,N_22809,N_22905);
nor U23024 (N_23024,N_22844,N_22946);
or U23025 (N_23025,N_22837,N_22982);
nand U23026 (N_23026,N_22989,N_22927);
and U23027 (N_23027,N_22864,N_22826);
nand U23028 (N_23028,N_22916,N_22975);
nand U23029 (N_23029,N_22814,N_22973);
xnor U23030 (N_23030,N_22945,N_22917);
or U23031 (N_23031,N_22968,N_22995);
or U23032 (N_23032,N_22842,N_22932);
nor U23033 (N_23033,N_22813,N_22835);
and U23034 (N_23034,N_22941,N_22812);
xor U23035 (N_23035,N_22992,N_22833);
nand U23036 (N_23036,N_22959,N_22891);
nand U23037 (N_23037,N_22867,N_22961);
or U23038 (N_23038,N_22805,N_22972);
xnor U23039 (N_23039,N_22957,N_22947);
nor U23040 (N_23040,N_22839,N_22923);
nand U23041 (N_23041,N_22940,N_22822);
and U23042 (N_23042,N_22935,N_22882);
xnor U23043 (N_23043,N_22918,N_22980);
xnor U23044 (N_23044,N_22884,N_22909);
nor U23045 (N_23045,N_22938,N_22948);
nand U23046 (N_23046,N_22846,N_22875);
and U23047 (N_23047,N_22969,N_22942);
nand U23048 (N_23048,N_22877,N_22863);
and U23049 (N_23049,N_22801,N_22960);
or U23050 (N_23050,N_22819,N_22991);
nand U23051 (N_23051,N_22904,N_22866);
nor U23052 (N_23052,N_22841,N_22962);
xnor U23053 (N_23053,N_22900,N_22886);
xor U23054 (N_23054,N_22815,N_22998);
nor U23055 (N_23055,N_22898,N_22970);
xor U23056 (N_23056,N_22929,N_22988);
nor U23057 (N_23057,N_22857,N_22847);
nand U23058 (N_23058,N_22930,N_22876);
nor U23059 (N_23059,N_22919,N_22979);
xor U23060 (N_23060,N_22913,N_22817);
or U23061 (N_23061,N_22829,N_22888);
nor U23062 (N_23062,N_22894,N_22879);
xnor U23063 (N_23063,N_22937,N_22806);
xnor U23064 (N_23064,N_22915,N_22885);
or U23065 (N_23065,N_22910,N_22981);
xor U23066 (N_23066,N_22956,N_22983);
xor U23067 (N_23067,N_22950,N_22848);
and U23068 (N_23068,N_22936,N_22880);
or U23069 (N_23069,N_22804,N_22971);
nand U23070 (N_23070,N_22907,N_22860);
or U23071 (N_23071,N_22944,N_22908);
nor U23072 (N_23072,N_22843,N_22985);
and U23073 (N_23073,N_22831,N_22994);
or U23074 (N_23074,N_22926,N_22883);
xnor U23075 (N_23075,N_22925,N_22965);
xor U23076 (N_23076,N_22943,N_22807);
xor U23077 (N_23077,N_22993,N_22963);
and U23078 (N_23078,N_22922,N_22951);
xor U23079 (N_23079,N_22820,N_22958);
nand U23080 (N_23080,N_22949,N_22978);
and U23081 (N_23081,N_22840,N_22830);
nor U23082 (N_23082,N_22873,N_22855);
nand U23083 (N_23083,N_22811,N_22952);
nand U23084 (N_23084,N_22827,N_22899);
xor U23085 (N_23085,N_22871,N_22838);
nand U23086 (N_23086,N_22824,N_22818);
nor U23087 (N_23087,N_22921,N_22816);
nor U23088 (N_23088,N_22878,N_22890);
xor U23089 (N_23089,N_22852,N_22954);
nand U23090 (N_23090,N_22828,N_22897);
nor U23091 (N_23091,N_22934,N_22974);
nor U23092 (N_23092,N_22803,N_22854);
or U23093 (N_23093,N_22823,N_22920);
xor U23094 (N_23094,N_22997,N_22955);
nand U23095 (N_23095,N_22996,N_22836);
nor U23096 (N_23096,N_22977,N_22802);
nor U23097 (N_23097,N_22901,N_22967);
nor U23098 (N_23098,N_22903,N_22892);
nor U23099 (N_23099,N_22990,N_22984);
xor U23100 (N_23100,N_22836,N_22863);
and U23101 (N_23101,N_22938,N_22892);
xor U23102 (N_23102,N_22948,N_22840);
xnor U23103 (N_23103,N_22874,N_22929);
and U23104 (N_23104,N_22869,N_22971);
nor U23105 (N_23105,N_22989,N_22968);
nor U23106 (N_23106,N_22898,N_22815);
nand U23107 (N_23107,N_22914,N_22861);
and U23108 (N_23108,N_22964,N_22829);
or U23109 (N_23109,N_22822,N_22871);
and U23110 (N_23110,N_22883,N_22922);
and U23111 (N_23111,N_22946,N_22989);
or U23112 (N_23112,N_22901,N_22965);
nor U23113 (N_23113,N_22874,N_22845);
nor U23114 (N_23114,N_22944,N_22934);
nor U23115 (N_23115,N_22983,N_22961);
or U23116 (N_23116,N_22942,N_22977);
xor U23117 (N_23117,N_22889,N_22920);
nand U23118 (N_23118,N_22801,N_22953);
xnor U23119 (N_23119,N_22848,N_22948);
nand U23120 (N_23120,N_22981,N_22989);
nor U23121 (N_23121,N_22995,N_22921);
or U23122 (N_23122,N_22818,N_22925);
nor U23123 (N_23123,N_22847,N_22817);
xor U23124 (N_23124,N_22851,N_22828);
nor U23125 (N_23125,N_22907,N_22843);
nor U23126 (N_23126,N_22823,N_22956);
nand U23127 (N_23127,N_22850,N_22919);
nand U23128 (N_23128,N_22844,N_22877);
or U23129 (N_23129,N_22935,N_22817);
xor U23130 (N_23130,N_22973,N_22986);
or U23131 (N_23131,N_22985,N_22959);
nand U23132 (N_23132,N_22886,N_22920);
nor U23133 (N_23133,N_22863,N_22915);
or U23134 (N_23134,N_22939,N_22900);
and U23135 (N_23135,N_22946,N_22901);
and U23136 (N_23136,N_22890,N_22829);
nor U23137 (N_23137,N_22884,N_22828);
or U23138 (N_23138,N_22947,N_22962);
and U23139 (N_23139,N_22903,N_22801);
nor U23140 (N_23140,N_22980,N_22842);
and U23141 (N_23141,N_22826,N_22964);
and U23142 (N_23142,N_22828,N_22816);
nor U23143 (N_23143,N_22870,N_22998);
nor U23144 (N_23144,N_22943,N_22857);
xnor U23145 (N_23145,N_22957,N_22815);
and U23146 (N_23146,N_22816,N_22929);
nor U23147 (N_23147,N_22934,N_22919);
nor U23148 (N_23148,N_22893,N_22988);
or U23149 (N_23149,N_22976,N_22936);
nand U23150 (N_23150,N_22902,N_22976);
or U23151 (N_23151,N_22948,N_22833);
nand U23152 (N_23152,N_22932,N_22983);
xor U23153 (N_23153,N_22883,N_22957);
and U23154 (N_23154,N_22827,N_22885);
nand U23155 (N_23155,N_22996,N_22890);
nor U23156 (N_23156,N_22937,N_22948);
nor U23157 (N_23157,N_22814,N_22857);
nand U23158 (N_23158,N_22959,N_22872);
nor U23159 (N_23159,N_22899,N_22857);
nor U23160 (N_23160,N_22994,N_22853);
xnor U23161 (N_23161,N_22865,N_22894);
nand U23162 (N_23162,N_22880,N_22939);
and U23163 (N_23163,N_22916,N_22824);
and U23164 (N_23164,N_22818,N_22949);
xor U23165 (N_23165,N_22820,N_22882);
nand U23166 (N_23166,N_22848,N_22952);
xnor U23167 (N_23167,N_22959,N_22867);
nor U23168 (N_23168,N_22997,N_22830);
nand U23169 (N_23169,N_22869,N_22861);
xor U23170 (N_23170,N_22840,N_22944);
nand U23171 (N_23171,N_22867,N_22966);
or U23172 (N_23172,N_22804,N_22873);
xor U23173 (N_23173,N_22980,N_22900);
nand U23174 (N_23174,N_22870,N_22905);
nor U23175 (N_23175,N_22876,N_22880);
xnor U23176 (N_23176,N_22831,N_22939);
nor U23177 (N_23177,N_22889,N_22839);
or U23178 (N_23178,N_22995,N_22867);
xor U23179 (N_23179,N_22950,N_22956);
xnor U23180 (N_23180,N_22918,N_22901);
nand U23181 (N_23181,N_22907,N_22948);
or U23182 (N_23182,N_22853,N_22827);
xor U23183 (N_23183,N_22998,N_22869);
xnor U23184 (N_23184,N_22832,N_22857);
nor U23185 (N_23185,N_22882,N_22856);
nor U23186 (N_23186,N_22954,N_22878);
or U23187 (N_23187,N_22987,N_22888);
xor U23188 (N_23188,N_22942,N_22867);
or U23189 (N_23189,N_22829,N_22896);
nor U23190 (N_23190,N_22966,N_22849);
nor U23191 (N_23191,N_22918,N_22952);
or U23192 (N_23192,N_22824,N_22822);
nand U23193 (N_23193,N_22993,N_22985);
and U23194 (N_23194,N_22875,N_22871);
xor U23195 (N_23195,N_22825,N_22898);
xor U23196 (N_23196,N_22851,N_22951);
or U23197 (N_23197,N_22823,N_22932);
nor U23198 (N_23198,N_22801,N_22916);
nor U23199 (N_23199,N_22832,N_22807);
nor U23200 (N_23200,N_23017,N_23173);
or U23201 (N_23201,N_23123,N_23066);
or U23202 (N_23202,N_23127,N_23145);
nor U23203 (N_23203,N_23042,N_23165);
or U23204 (N_23204,N_23046,N_23096);
and U23205 (N_23205,N_23172,N_23192);
or U23206 (N_23206,N_23113,N_23125);
or U23207 (N_23207,N_23100,N_23159);
or U23208 (N_23208,N_23097,N_23047);
xor U23209 (N_23209,N_23104,N_23164);
and U23210 (N_23210,N_23131,N_23161);
xor U23211 (N_23211,N_23124,N_23033);
nor U23212 (N_23212,N_23037,N_23137);
nand U23213 (N_23213,N_23052,N_23183);
nor U23214 (N_23214,N_23019,N_23011);
or U23215 (N_23215,N_23035,N_23048);
or U23216 (N_23216,N_23006,N_23054);
or U23217 (N_23217,N_23153,N_23149);
nand U23218 (N_23218,N_23069,N_23147);
nor U23219 (N_23219,N_23081,N_23143);
xor U23220 (N_23220,N_23176,N_23195);
nor U23221 (N_23221,N_23032,N_23103);
and U23222 (N_23222,N_23191,N_23030);
and U23223 (N_23223,N_23198,N_23078);
or U23224 (N_23224,N_23169,N_23074);
nor U23225 (N_23225,N_23175,N_23181);
and U23226 (N_23226,N_23013,N_23186);
or U23227 (N_23227,N_23082,N_23063);
xor U23228 (N_23228,N_23133,N_23008);
nand U23229 (N_23229,N_23031,N_23023);
nand U23230 (N_23230,N_23050,N_23062);
or U23231 (N_23231,N_23026,N_23193);
nor U23232 (N_23232,N_23136,N_23053);
and U23233 (N_23233,N_23064,N_23044);
nor U23234 (N_23234,N_23132,N_23068);
nand U23235 (N_23235,N_23197,N_23120);
or U23236 (N_23236,N_23150,N_23085);
nand U23237 (N_23237,N_23094,N_23065);
nor U23238 (N_23238,N_23028,N_23141);
or U23239 (N_23239,N_23199,N_23056);
and U23240 (N_23240,N_23049,N_23177);
or U23241 (N_23241,N_23060,N_23027);
nand U23242 (N_23242,N_23101,N_23025);
or U23243 (N_23243,N_23105,N_23134);
nor U23244 (N_23244,N_23187,N_23111);
and U23245 (N_23245,N_23170,N_23073);
and U23246 (N_23246,N_23142,N_23093);
nor U23247 (N_23247,N_23022,N_23115);
xnor U23248 (N_23248,N_23016,N_23036);
or U23249 (N_23249,N_23171,N_23058);
or U23250 (N_23250,N_23070,N_23041);
nand U23251 (N_23251,N_23189,N_23040);
or U23252 (N_23252,N_23167,N_23014);
nand U23253 (N_23253,N_23039,N_23021);
nand U23254 (N_23254,N_23001,N_23190);
or U23255 (N_23255,N_23106,N_23067);
and U23256 (N_23256,N_23088,N_23148);
nand U23257 (N_23257,N_23015,N_23139);
nand U23258 (N_23258,N_23178,N_23071);
nor U23259 (N_23259,N_23012,N_23122);
nor U23260 (N_23260,N_23018,N_23155);
or U23261 (N_23261,N_23163,N_23154);
xnor U23262 (N_23262,N_23000,N_23144);
or U23263 (N_23263,N_23146,N_23121);
xnor U23264 (N_23264,N_23152,N_23072);
xnor U23265 (N_23265,N_23077,N_23117);
nand U23266 (N_23266,N_23091,N_23188);
and U23267 (N_23267,N_23184,N_23158);
xor U23268 (N_23268,N_23157,N_23003);
xnor U23269 (N_23269,N_23130,N_23057);
xor U23270 (N_23270,N_23180,N_23162);
and U23271 (N_23271,N_23151,N_23095);
nand U23272 (N_23272,N_23090,N_23099);
or U23273 (N_23273,N_23055,N_23107);
nand U23274 (N_23274,N_23084,N_23076);
and U23275 (N_23275,N_23119,N_23002);
nor U23276 (N_23276,N_23138,N_23086);
and U23277 (N_23277,N_23109,N_23034);
nand U23278 (N_23278,N_23112,N_23140);
or U23279 (N_23279,N_23129,N_23004);
and U23280 (N_23280,N_23118,N_23182);
or U23281 (N_23281,N_23079,N_23116);
nor U23282 (N_23282,N_23166,N_23061);
or U23283 (N_23283,N_23098,N_23043);
xnor U23284 (N_23284,N_23092,N_23005);
nor U23285 (N_23285,N_23075,N_23007);
or U23286 (N_23286,N_23196,N_23059);
and U23287 (N_23287,N_23009,N_23179);
nor U23288 (N_23288,N_23114,N_23135);
nor U23289 (N_23289,N_23108,N_23083);
xnor U23290 (N_23290,N_23128,N_23160);
and U23291 (N_23291,N_23051,N_23045);
xnor U23292 (N_23292,N_23185,N_23024);
or U23293 (N_23293,N_23029,N_23126);
xnor U23294 (N_23294,N_23010,N_23174);
and U23295 (N_23295,N_23102,N_23020);
xor U23296 (N_23296,N_23089,N_23038);
and U23297 (N_23297,N_23194,N_23156);
xnor U23298 (N_23298,N_23110,N_23168);
xor U23299 (N_23299,N_23087,N_23080);
and U23300 (N_23300,N_23092,N_23142);
nor U23301 (N_23301,N_23168,N_23040);
xor U23302 (N_23302,N_23052,N_23090);
nand U23303 (N_23303,N_23169,N_23037);
or U23304 (N_23304,N_23075,N_23183);
nand U23305 (N_23305,N_23024,N_23058);
nand U23306 (N_23306,N_23143,N_23115);
and U23307 (N_23307,N_23057,N_23046);
nor U23308 (N_23308,N_23029,N_23132);
nor U23309 (N_23309,N_23186,N_23143);
nand U23310 (N_23310,N_23092,N_23184);
and U23311 (N_23311,N_23147,N_23049);
or U23312 (N_23312,N_23168,N_23089);
and U23313 (N_23313,N_23190,N_23110);
xor U23314 (N_23314,N_23002,N_23160);
and U23315 (N_23315,N_23140,N_23031);
or U23316 (N_23316,N_23133,N_23107);
and U23317 (N_23317,N_23159,N_23074);
or U23318 (N_23318,N_23046,N_23159);
nand U23319 (N_23319,N_23096,N_23001);
nor U23320 (N_23320,N_23109,N_23055);
nor U23321 (N_23321,N_23135,N_23100);
or U23322 (N_23322,N_23133,N_23053);
nor U23323 (N_23323,N_23149,N_23042);
xor U23324 (N_23324,N_23138,N_23148);
or U23325 (N_23325,N_23139,N_23128);
and U23326 (N_23326,N_23044,N_23003);
nand U23327 (N_23327,N_23173,N_23135);
nor U23328 (N_23328,N_23191,N_23199);
or U23329 (N_23329,N_23061,N_23052);
and U23330 (N_23330,N_23063,N_23147);
and U23331 (N_23331,N_23073,N_23122);
xor U23332 (N_23332,N_23042,N_23056);
nand U23333 (N_23333,N_23164,N_23059);
nor U23334 (N_23334,N_23082,N_23134);
nand U23335 (N_23335,N_23187,N_23168);
nand U23336 (N_23336,N_23151,N_23057);
xnor U23337 (N_23337,N_23120,N_23150);
xor U23338 (N_23338,N_23022,N_23129);
nor U23339 (N_23339,N_23179,N_23055);
or U23340 (N_23340,N_23074,N_23015);
xnor U23341 (N_23341,N_23010,N_23066);
xnor U23342 (N_23342,N_23188,N_23104);
or U23343 (N_23343,N_23037,N_23063);
nor U23344 (N_23344,N_23185,N_23095);
or U23345 (N_23345,N_23073,N_23026);
nand U23346 (N_23346,N_23066,N_23132);
or U23347 (N_23347,N_23133,N_23195);
and U23348 (N_23348,N_23115,N_23068);
and U23349 (N_23349,N_23029,N_23171);
or U23350 (N_23350,N_23005,N_23122);
and U23351 (N_23351,N_23185,N_23009);
or U23352 (N_23352,N_23009,N_23076);
nand U23353 (N_23353,N_23009,N_23023);
nor U23354 (N_23354,N_23197,N_23122);
nor U23355 (N_23355,N_23175,N_23138);
or U23356 (N_23356,N_23074,N_23008);
xnor U23357 (N_23357,N_23190,N_23063);
nand U23358 (N_23358,N_23198,N_23085);
or U23359 (N_23359,N_23001,N_23062);
nor U23360 (N_23360,N_23090,N_23005);
or U23361 (N_23361,N_23003,N_23028);
or U23362 (N_23362,N_23192,N_23169);
xor U23363 (N_23363,N_23186,N_23060);
or U23364 (N_23364,N_23148,N_23090);
xor U23365 (N_23365,N_23146,N_23016);
nor U23366 (N_23366,N_23035,N_23059);
nand U23367 (N_23367,N_23056,N_23007);
or U23368 (N_23368,N_23102,N_23124);
and U23369 (N_23369,N_23090,N_23017);
xnor U23370 (N_23370,N_23180,N_23132);
and U23371 (N_23371,N_23192,N_23000);
nor U23372 (N_23372,N_23116,N_23181);
xnor U23373 (N_23373,N_23105,N_23170);
nor U23374 (N_23374,N_23140,N_23014);
or U23375 (N_23375,N_23187,N_23135);
xnor U23376 (N_23376,N_23184,N_23009);
and U23377 (N_23377,N_23160,N_23024);
xor U23378 (N_23378,N_23002,N_23042);
xnor U23379 (N_23379,N_23100,N_23054);
nand U23380 (N_23380,N_23055,N_23142);
nand U23381 (N_23381,N_23091,N_23063);
nor U23382 (N_23382,N_23114,N_23192);
and U23383 (N_23383,N_23003,N_23115);
and U23384 (N_23384,N_23061,N_23190);
nor U23385 (N_23385,N_23095,N_23111);
or U23386 (N_23386,N_23085,N_23026);
or U23387 (N_23387,N_23174,N_23000);
xnor U23388 (N_23388,N_23189,N_23022);
and U23389 (N_23389,N_23037,N_23083);
xor U23390 (N_23390,N_23076,N_23008);
or U23391 (N_23391,N_23178,N_23028);
or U23392 (N_23392,N_23024,N_23183);
xor U23393 (N_23393,N_23016,N_23015);
or U23394 (N_23394,N_23078,N_23107);
nand U23395 (N_23395,N_23145,N_23070);
xor U23396 (N_23396,N_23099,N_23020);
or U23397 (N_23397,N_23106,N_23126);
and U23398 (N_23398,N_23020,N_23031);
nand U23399 (N_23399,N_23041,N_23172);
nand U23400 (N_23400,N_23255,N_23260);
xor U23401 (N_23401,N_23205,N_23304);
nor U23402 (N_23402,N_23363,N_23322);
xnor U23403 (N_23403,N_23334,N_23239);
nand U23404 (N_23404,N_23291,N_23332);
or U23405 (N_23405,N_23387,N_23373);
nand U23406 (N_23406,N_23273,N_23326);
xnor U23407 (N_23407,N_23353,N_23370);
nand U23408 (N_23408,N_23395,N_23390);
nand U23409 (N_23409,N_23323,N_23352);
or U23410 (N_23410,N_23218,N_23252);
nand U23411 (N_23411,N_23271,N_23246);
nor U23412 (N_23412,N_23394,N_23368);
or U23413 (N_23413,N_23241,N_23340);
nor U23414 (N_23414,N_23372,N_23287);
and U23415 (N_23415,N_23357,N_23354);
or U23416 (N_23416,N_23311,N_23336);
or U23417 (N_23417,N_23284,N_23208);
nand U23418 (N_23418,N_23277,N_23207);
xnor U23419 (N_23419,N_23325,N_23283);
and U23420 (N_23420,N_23209,N_23316);
xor U23421 (N_23421,N_23342,N_23347);
nor U23422 (N_23422,N_23393,N_23303);
nand U23423 (N_23423,N_23339,N_23244);
or U23424 (N_23424,N_23221,N_23201);
nor U23425 (N_23425,N_23275,N_23234);
nor U23426 (N_23426,N_23281,N_23220);
or U23427 (N_23427,N_23375,N_23343);
nor U23428 (N_23428,N_23288,N_23219);
nor U23429 (N_23429,N_23389,N_23314);
nor U23430 (N_23430,N_23338,N_23286);
nor U23431 (N_23431,N_23321,N_23381);
nand U23432 (N_23432,N_23297,N_23337);
xnor U23433 (N_23433,N_23214,N_23227);
nand U23434 (N_23434,N_23274,N_23280);
or U23435 (N_23435,N_23315,N_23279);
nor U23436 (N_23436,N_23211,N_23391);
and U23437 (N_23437,N_23240,N_23224);
or U23438 (N_23438,N_23235,N_23242);
nor U23439 (N_23439,N_23309,N_23399);
or U23440 (N_23440,N_23225,N_23230);
or U23441 (N_23441,N_23302,N_23380);
nand U23442 (N_23442,N_23212,N_23362);
and U23443 (N_23443,N_23258,N_23293);
and U23444 (N_23444,N_23251,N_23312);
nand U23445 (N_23445,N_23366,N_23276);
xor U23446 (N_23446,N_23213,N_23327);
nand U23447 (N_23447,N_23261,N_23317);
and U23448 (N_23448,N_23203,N_23383);
nor U23449 (N_23449,N_23268,N_23341);
or U23450 (N_23450,N_23256,N_23346);
or U23451 (N_23451,N_23377,N_23295);
and U23452 (N_23452,N_23266,N_23204);
and U23453 (N_23453,N_23289,N_23324);
nand U23454 (N_23454,N_23229,N_23202);
or U23455 (N_23455,N_23231,N_23200);
xor U23456 (N_23456,N_23247,N_23398);
or U23457 (N_23457,N_23300,N_23365);
and U23458 (N_23458,N_23392,N_23335);
or U23459 (N_23459,N_23360,N_23385);
or U23460 (N_23460,N_23344,N_23249);
xnor U23461 (N_23461,N_23374,N_23358);
and U23462 (N_23462,N_23263,N_23243);
and U23463 (N_23463,N_23259,N_23329);
nand U23464 (N_23464,N_23350,N_23298);
nor U23465 (N_23465,N_23384,N_23310);
or U23466 (N_23466,N_23328,N_23348);
nand U23467 (N_23467,N_23364,N_23376);
nand U23468 (N_23468,N_23278,N_23359);
nand U23469 (N_23469,N_23367,N_23396);
or U23470 (N_23470,N_23330,N_23301);
nor U23471 (N_23471,N_23355,N_23382);
nor U23472 (N_23472,N_23285,N_23228);
nand U23473 (N_23473,N_23257,N_23253);
nor U23474 (N_23474,N_23292,N_23369);
or U23475 (N_23475,N_23371,N_23307);
or U23476 (N_23476,N_23299,N_23351);
xnor U23477 (N_23477,N_23210,N_23215);
nand U23478 (N_23478,N_23319,N_23306);
nand U23479 (N_23479,N_23232,N_23217);
nor U23480 (N_23480,N_23378,N_23356);
nand U23481 (N_23481,N_23272,N_23388);
xnor U23482 (N_23482,N_23379,N_23290);
nor U23483 (N_23483,N_23250,N_23361);
nor U23484 (N_23484,N_23238,N_23245);
nor U23485 (N_23485,N_23222,N_23331);
nor U23486 (N_23486,N_23320,N_23318);
nor U23487 (N_23487,N_23254,N_23397);
nand U23488 (N_23488,N_23237,N_23223);
xnor U23489 (N_23489,N_23269,N_23265);
xnor U23490 (N_23490,N_23305,N_23386);
xor U23491 (N_23491,N_23345,N_23313);
or U23492 (N_23492,N_23226,N_23270);
and U23493 (N_23493,N_23282,N_23206);
and U23494 (N_23494,N_23264,N_23296);
or U23495 (N_23495,N_23216,N_23233);
or U23496 (N_23496,N_23349,N_23333);
nor U23497 (N_23497,N_23236,N_23267);
nand U23498 (N_23498,N_23262,N_23248);
nor U23499 (N_23499,N_23308,N_23294);
or U23500 (N_23500,N_23333,N_23288);
nor U23501 (N_23501,N_23326,N_23206);
nand U23502 (N_23502,N_23282,N_23291);
nand U23503 (N_23503,N_23219,N_23351);
nand U23504 (N_23504,N_23250,N_23350);
nand U23505 (N_23505,N_23292,N_23325);
nand U23506 (N_23506,N_23281,N_23209);
nand U23507 (N_23507,N_23321,N_23338);
nand U23508 (N_23508,N_23275,N_23302);
and U23509 (N_23509,N_23383,N_23330);
nor U23510 (N_23510,N_23217,N_23246);
nand U23511 (N_23511,N_23342,N_23267);
and U23512 (N_23512,N_23257,N_23395);
nor U23513 (N_23513,N_23382,N_23291);
xnor U23514 (N_23514,N_23348,N_23308);
and U23515 (N_23515,N_23373,N_23395);
nand U23516 (N_23516,N_23328,N_23325);
and U23517 (N_23517,N_23321,N_23329);
nand U23518 (N_23518,N_23370,N_23316);
or U23519 (N_23519,N_23313,N_23324);
nand U23520 (N_23520,N_23333,N_23357);
xnor U23521 (N_23521,N_23293,N_23278);
and U23522 (N_23522,N_23361,N_23254);
or U23523 (N_23523,N_23240,N_23234);
or U23524 (N_23524,N_23397,N_23292);
nand U23525 (N_23525,N_23249,N_23377);
or U23526 (N_23526,N_23366,N_23359);
or U23527 (N_23527,N_23346,N_23307);
nand U23528 (N_23528,N_23222,N_23374);
or U23529 (N_23529,N_23296,N_23315);
nor U23530 (N_23530,N_23239,N_23236);
and U23531 (N_23531,N_23394,N_23232);
nand U23532 (N_23532,N_23325,N_23396);
xnor U23533 (N_23533,N_23338,N_23256);
nand U23534 (N_23534,N_23240,N_23218);
and U23535 (N_23535,N_23251,N_23276);
or U23536 (N_23536,N_23340,N_23375);
or U23537 (N_23537,N_23282,N_23284);
xnor U23538 (N_23538,N_23382,N_23290);
nand U23539 (N_23539,N_23328,N_23286);
or U23540 (N_23540,N_23385,N_23291);
xnor U23541 (N_23541,N_23362,N_23234);
xnor U23542 (N_23542,N_23373,N_23346);
and U23543 (N_23543,N_23273,N_23368);
nor U23544 (N_23544,N_23212,N_23391);
nand U23545 (N_23545,N_23388,N_23328);
and U23546 (N_23546,N_23218,N_23345);
nand U23547 (N_23547,N_23388,N_23203);
nand U23548 (N_23548,N_23268,N_23340);
or U23549 (N_23549,N_23272,N_23371);
or U23550 (N_23550,N_23243,N_23364);
nor U23551 (N_23551,N_23260,N_23399);
nor U23552 (N_23552,N_23395,N_23293);
nand U23553 (N_23553,N_23359,N_23228);
nand U23554 (N_23554,N_23313,N_23319);
and U23555 (N_23555,N_23342,N_23212);
nor U23556 (N_23556,N_23228,N_23287);
nand U23557 (N_23557,N_23334,N_23333);
nand U23558 (N_23558,N_23329,N_23335);
and U23559 (N_23559,N_23305,N_23237);
or U23560 (N_23560,N_23340,N_23330);
and U23561 (N_23561,N_23298,N_23394);
and U23562 (N_23562,N_23284,N_23356);
nor U23563 (N_23563,N_23320,N_23325);
and U23564 (N_23564,N_23322,N_23276);
xor U23565 (N_23565,N_23239,N_23203);
or U23566 (N_23566,N_23341,N_23233);
and U23567 (N_23567,N_23360,N_23284);
xnor U23568 (N_23568,N_23262,N_23249);
nand U23569 (N_23569,N_23339,N_23391);
and U23570 (N_23570,N_23382,N_23314);
nand U23571 (N_23571,N_23303,N_23237);
nand U23572 (N_23572,N_23386,N_23366);
nor U23573 (N_23573,N_23391,N_23282);
nand U23574 (N_23574,N_23261,N_23388);
nand U23575 (N_23575,N_23349,N_23337);
nor U23576 (N_23576,N_23333,N_23363);
and U23577 (N_23577,N_23334,N_23367);
and U23578 (N_23578,N_23205,N_23363);
xor U23579 (N_23579,N_23387,N_23230);
and U23580 (N_23580,N_23243,N_23331);
and U23581 (N_23581,N_23384,N_23372);
nor U23582 (N_23582,N_23332,N_23321);
nor U23583 (N_23583,N_23226,N_23383);
xor U23584 (N_23584,N_23202,N_23320);
nand U23585 (N_23585,N_23344,N_23393);
and U23586 (N_23586,N_23270,N_23244);
xor U23587 (N_23587,N_23285,N_23304);
nor U23588 (N_23588,N_23244,N_23316);
xor U23589 (N_23589,N_23289,N_23357);
and U23590 (N_23590,N_23381,N_23318);
nand U23591 (N_23591,N_23369,N_23288);
xnor U23592 (N_23592,N_23334,N_23282);
or U23593 (N_23593,N_23313,N_23232);
xnor U23594 (N_23594,N_23274,N_23356);
nor U23595 (N_23595,N_23327,N_23329);
and U23596 (N_23596,N_23225,N_23280);
xnor U23597 (N_23597,N_23226,N_23279);
and U23598 (N_23598,N_23280,N_23298);
nor U23599 (N_23599,N_23349,N_23264);
xnor U23600 (N_23600,N_23562,N_23583);
nor U23601 (N_23601,N_23505,N_23493);
and U23602 (N_23602,N_23538,N_23530);
and U23603 (N_23603,N_23591,N_23484);
xor U23604 (N_23604,N_23474,N_23407);
or U23605 (N_23605,N_23568,N_23563);
xor U23606 (N_23606,N_23525,N_23461);
nor U23607 (N_23607,N_23464,N_23428);
xor U23608 (N_23608,N_23413,N_23572);
nor U23609 (N_23609,N_23449,N_23501);
nand U23610 (N_23610,N_23536,N_23435);
xor U23611 (N_23611,N_23586,N_23470);
and U23612 (N_23612,N_23520,N_23419);
nand U23613 (N_23613,N_23514,N_23575);
nor U23614 (N_23614,N_23596,N_23448);
xnor U23615 (N_23615,N_23518,N_23479);
and U23616 (N_23616,N_23517,N_23439);
nand U23617 (N_23617,N_23532,N_23422);
nand U23618 (N_23618,N_23414,N_23534);
xor U23619 (N_23619,N_23485,N_23421);
or U23620 (N_23620,N_23537,N_23475);
xnor U23621 (N_23621,N_23565,N_23542);
and U23622 (N_23622,N_23497,N_23547);
nor U23623 (N_23623,N_23406,N_23504);
nand U23624 (N_23624,N_23473,N_23507);
and U23625 (N_23625,N_23543,N_23441);
nor U23626 (N_23626,N_23594,N_23416);
xor U23627 (N_23627,N_23495,N_23432);
nand U23628 (N_23628,N_23533,N_23494);
nand U23629 (N_23629,N_23540,N_23579);
and U23630 (N_23630,N_23593,N_23554);
or U23631 (N_23631,N_23411,N_23451);
and U23632 (N_23632,N_23443,N_23557);
nand U23633 (N_23633,N_23506,N_23477);
or U23634 (N_23634,N_23558,N_23576);
nand U23635 (N_23635,N_23402,N_23412);
nor U23636 (N_23636,N_23427,N_23527);
nand U23637 (N_23637,N_23508,N_23588);
nand U23638 (N_23638,N_23481,N_23552);
nand U23639 (N_23639,N_23555,N_23577);
and U23640 (N_23640,N_23528,N_23444);
and U23641 (N_23641,N_23465,N_23417);
nor U23642 (N_23642,N_23489,N_23569);
nand U23643 (N_23643,N_23560,N_23453);
and U23644 (N_23644,N_23578,N_23456);
or U23645 (N_23645,N_23436,N_23403);
or U23646 (N_23646,N_23483,N_23503);
and U23647 (N_23647,N_23492,N_23437);
xor U23648 (N_23648,N_23467,N_23434);
nand U23649 (N_23649,N_23488,N_23556);
nand U23650 (N_23650,N_23440,N_23400);
nand U23651 (N_23651,N_23500,N_23454);
or U23652 (N_23652,N_23452,N_23580);
nor U23653 (N_23653,N_23460,N_23418);
nor U23654 (N_23654,N_23431,N_23447);
and U23655 (N_23655,N_23438,N_23426);
or U23656 (N_23656,N_23566,N_23468);
or U23657 (N_23657,N_23521,N_23599);
xor U23658 (N_23658,N_23512,N_23564);
nand U23659 (N_23659,N_23545,N_23425);
or U23660 (N_23660,N_23482,N_23574);
or U23661 (N_23661,N_23509,N_23567);
or U23662 (N_23662,N_23478,N_23490);
xor U23663 (N_23663,N_23502,N_23549);
xor U23664 (N_23664,N_23433,N_23598);
xor U23665 (N_23665,N_23582,N_23526);
xor U23666 (N_23666,N_23496,N_23573);
or U23667 (N_23667,N_23523,N_23513);
and U23668 (N_23668,N_23531,N_23510);
and U23669 (N_23669,N_23559,N_23553);
xnor U23670 (N_23670,N_23511,N_23486);
xnor U23671 (N_23671,N_23458,N_23541);
nand U23672 (N_23672,N_23592,N_23404);
or U23673 (N_23673,N_23546,N_23498);
or U23674 (N_23674,N_23408,N_23463);
nand U23675 (N_23675,N_23539,N_23522);
nor U23676 (N_23676,N_23561,N_23471);
and U23677 (N_23677,N_23466,N_23524);
and U23678 (N_23678,N_23405,N_23487);
or U23679 (N_23679,N_23445,N_23491);
or U23680 (N_23680,N_23462,N_23584);
xnor U23681 (N_23681,N_23430,N_23401);
nor U23682 (N_23682,N_23499,N_23420);
and U23683 (N_23683,N_23581,N_23595);
and U23684 (N_23684,N_23535,N_23570);
nor U23685 (N_23685,N_23455,N_23410);
or U23686 (N_23686,N_23415,N_23450);
nand U23687 (N_23687,N_23585,N_23476);
nand U23688 (N_23688,N_23429,N_23544);
nor U23689 (N_23689,N_23457,N_23550);
nor U23690 (N_23690,N_23442,N_23469);
nor U23691 (N_23691,N_23587,N_23529);
nand U23692 (N_23692,N_23597,N_23423);
nor U23693 (N_23693,N_23459,N_23590);
nor U23694 (N_23694,N_23472,N_23409);
or U23695 (N_23695,N_23571,N_23516);
or U23696 (N_23696,N_23519,N_23446);
and U23697 (N_23697,N_23589,N_23480);
xnor U23698 (N_23698,N_23515,N_23548);
and U23699 (N_23699,N_23551,N_23424);
and U23700 (N_23700,N_23454,N_23570);
xnor U23701 (N_23701,N_23563,N_23466);
nor U23702 (N_23702,N_23489,N_23437);
nand U23703 (N_23703,N_23554,N_23548);
xnor U23704 (N_23704,N_23516,N_23463);
nand U23705 (N_23705,N_23519,N_23586);
or U23706 (N_23706,N_23432,N_23409);
or U23707 (N_23707,N_23475,N_23429);
or U23708 (N_23708,N_23567,N_23498);
or U23709 (N_23709,N_23408,N_23492);
nand U23710 (N_23710,N_23461,N_23594);
nand U23711 (N_23711,N_23571,N_23450);
nand U23712 (N_23712,N_23424,N_23433);
nand U23713 (N_23713,N_23427,N_23449);
or U23714 (N_23714,N_23581,N_23529);
or U23715 (N_23715,N_23517,N_23591);
nand U23716 (N_23716,N_23589,N_23484);
nor U23717 (N_23717,N_23587,N_23424);
and U23718 (N_23718,N_23424,N_23549);
and U23719 (N_23719,N_23439,N_23485);
nand U23720 (N_23720,N_23427,N_23514);
xor U23721 (N_23721,N_23533,N_23498);
xnor U23722 (N_23722,N_23466,N_23448);
xnor U23723 (N_23723,N_23488,N_23505);
nand U23724 (N_23724,N_23479,N_23472);
nand U23725 (N_23725,N_23464,N_23504);
or U23726 (N_23726,N_23565,N_23587);
and U23727 (N_23727,N_23545,N_23584);
nand U23728 (N_23728,N_23543,N_23571);
or U23729 (N_23729,N_23456,N_23508);
or U23730 (N_23730,N_23503,N_23485);
and U23731 (N_23731,N_23452,N_23527);
or U23732 (N_23732,N_23551,N_23576);
or U23733 (N_23733,N_23587,N_23434);
or U23734 (N_23734,N_23435,N_23527);
xnor U23735 (N_23735,N_23450,N_23454);
xnor U23736 (N_23736,N_23409,N_23562);
and U23737 (N_23737,N_23499,N_23492);
or U23738 (N_23738,N_23403,N_23531);
or U23739 (N_23739,N_23401,N_23519);
or U23740 (N_23740,N_23589,N_23440);
or U23741 (N_23741,N_23538,N_23463);
nor U23742 (N_23742,N_23461,N_23426);
and U23743 (N_23743,N_23401,N_23557);
nand U23744 (N_23744,N_23447,N_23555);
and U23745 (N_23745,N_23553,N_23420);
or U23746 (N_23746,N_23566,N_23544);
nor U23747 (N_23747,N_23538,N_23413);
nor U23748 (N_23748,N_23525,N_23528);
nand U23749 (N_23749,N_23438,N_23498);
xnor U23750 (N_23750,N_23548,N_23542);
and U23751 (N_23751,N_23460,N_23597);
or U23752 (N_23752,N_23436,N_23569);
nor U23753 (N_23753,N_23417,N_23416);
or U23754 (N_23754,N_23400,N_23419);
nand U23755 (N_23755,N_23460,N_23406);
and U23756 (N_23756,N_23585,N_23425);
nor U23757 (N_23757,N_23539,N_23450);
or U23758 (N_23758,N_23515,N_23583);
nor U23759 (N_23759,N_23595,N_23570);
nand U23760 (N_23760,N_23540,N_23531);
xor U23761 (N_23761,N_23484,N_23486);
nand U23762 (N_23762,N_23425,N_23416);
xnor U23763 (N_23763,N_23530,N_23475);
nor U23764 (N_23764,N_23575,N_23465);
nor U23765 (N_23765,N_23457,N_23416);
and U23766 (N_23766,N_23583,N_23589);
nor U23767 (N_23767,N_23417,N_23433);
xnor U23768 (N_23768,N_23598,N_23418);
nand U23769 (N_23769,N_23512,N_23473);
or U23770 (N_23770,N_23468,N_23470);
xor U23771 (N_23771,N_23497,N_23437);
and U23772 (N_23772,N_23493,N_23407);
or U23773 (N_23773,N_23430,N_23405);
or U23774 (N_23774,N_23501,N_23529);
xnor U23775 (N_23775,N_23514,N_23583);
and U23776 (N_23776,N_23404,N_23424);
xor U23777 (N_23777,N_23460,N_23415);
nor U23778 (N_23778,N_23506,N_23498);
xnor U23779 (N_23779,N_23554,N_23447);
nand U23780 (N_23780,N_23465,N_23522);
and U23781 (N_23781,N_23558,N_23453);
nor U23782 (N_23782,N_23527,N_23422);
and U23783 (N_23783,N_23465,N_23422);
nand U23784 (N_23784,N_23511,N_23438);
nand U23785 (N_23785,N_23409,N_23521);
xor U23786 (N_23786,N_23521,N_23503);
and U23787 (N_23787,N_23400,N_23495);
or U23788 (N_23788,N_23529,N_23497);
or U23789 (N_23789,N_23537,N_23409);
nor U23790 (N_23790,N_23458,N_23582);
xor U23791 (N_23791,N_23407,N_23417);
nor U23792 (N_23792,N_23529,N_23559);
and U23793 (N_23793,N_23472,N_23482);
nand U23794 (N_23794,N_23548,N_23475);
or U23795 (N_23795,N_23598,N_23549);
or U23796 (N_23796,N_23441,N_23558);
or U23797 (N_23797,N_23500,N_23479);
nand U23798 (N_23798,N_23526,N_23473);
and U23799 (N_23799,N_23417,N_23571);
xnor U23800 (N_23800,N_23676,N_23696);
xnor U23801 (N_23801,N_23635,N_23714);
nor U23802 (N_23802,N_23624,N_23703);
nor U23803 (N_23803,N_23617,N_23723);
nand U23804 (N_23804,N_23763,N_23608);
nor U23805 (N_23805,N_23650,N_23636);
and U23806 (N_23806,N_23735,N_23750);
nor U23807 (N_23807,N_23733,N_23737);
nand U23808 (N_23808,N_23616,N_23756);
xnor U23809 (N_23809,N_23773,N_23700);
nand U23810 (N_23810,N_23762,N_23705);
nor U23811 (N_23811,N_23739,N_23660);
or U23812 (N_23812,N_23602,N_23771);
and U23813 (N_23813,N_23693,N_23727);
and U23814 (N_23814,N_23688,N_23686);
nor U23815 (N_23815,N_23767,N_23615);
or U23816 (N_23816,N_23611,N_23760);
nand U23817 (N_23817,N_23781,N_23697);
nor U23818 (N_23818,N_23792,N_23618);
xor U23819 (N_23819,N_23662,N_23674);
or U23820 (N_23820,N_23725,N_23755);
and U23821 (N_23821,N_23659,N_23622);
nand U23822 (N_23822,N_23743,N_23652);
nand U23823 (N_23823,N_23603,N_23729);
and U23824 (N_23824,N_23761,N_23783);
and U23825 (N_23825,N_23790,N_23741);
nand U23826 (N_23826,N_23644,N_23774);
and U23827 (N_23827,N_23621,N_23604);
xor U23828 (N_23828,N_23655,N_23656);
xnor U23829 (N_23829,N_23791,N_23752);
nor U23830 (N_23830,N_23630,N_23775);
or U23831 (N_23831,N_23613,N_23785);
nand U23832 (N_23832,N_23769,N_23661);
xor U23833 (N_23833,N_23744,N_23722);
and U23834 (N_23834,N_23665,N_23787);
and U23835 (N_23835,N_23753,N_23634);
nor U23836 (N_23836,N_23643,N_23742);
xor U23837 (N_23837,N_23724,N_23628);
or U23838 (N_23838,N_23718,N_23715);
and U23839 (N_23839,N_23667,N_23637);
nand U23840 (N_23840,N_23664,N_23759);
nor U23841 (N_23841,N_23779,N_23757);
and U23842 (N_23842,N_23614,N_23709);
xnor U23843 (N_23843,N_23736,N_23766);
or U23844 (N_23844,N_23632,N_23683);
nor U23845 (N_23845,N_23768,N_23695);
nor U23846 (N_23846,N_23788,N_23669);
nor U23847 (N_23847,N_23654,N_23646);
and U23848 (N_23848,N_23680,N_23716);
and U23849 (N_23849,N_23670,N_23708);
and U23850 (N_23850,N_23641,N_23645);
or U23851 (N_23851,N_23607,N_23796);
nor U23852 (N_23852,N_23789,N_23648);
nand U23853 (N_23853,N_23710,N_23786);
or U23854 (N_23854,N_23782,N_23797);
xnor U23855 (N_23855,N_23619,N_23799);
and U23856 (N_23856,N_23620,N_23679);
or U23857 (N_23857,N_23726,N_23706);
nand U23858 (N_23858,N_23631,N_23704);
nand U23859 (N_23859,N_23793,N_23601);
nor U23860 (N_23860,N_23698,N_23649);
and U23861 (N_23861,N_23677,N_23633);
nand U23862 (N_23862,N_23682,N_23663);
nor U23863 (N_23863,N_23711,N_23798);
nor U23864 (N_23864,N_23731,N_23692);
and U23865 (N_23865,N_23610,N_23627);
and U23866 (N_23866,N_23605,N_23638);
or U23867 (N_23867,N_23778,N_23780);
or U23868 (N_23868,N_23600,N_23751);
or U23869 (N_23869,N_23672,N_23747);
nor U23870 (N_23870,N_23758,N_23699);
xnor U23871 (N_23871,N_23690,N_23740);
and U23872 (N_23872,N_23754,N_23748);
nor U23873 (N_23873,N_23707,N_23713);
and U23874 (N_23874,N_23720,N_23626);
and U23875 (N_23875,N_23738,N_23795);
xor U23876 (N_23876,N_23653,N_23685);
nor U23877 (N_23877,N_23777,N_23749);
xnor U23878 (N_23878,N_23732,N_23730);
and U23879 (N_23879,N_23623,N_23678);
xor U23880 (N_23880,N_23784,N_23681);
or U23881 (N_23881,N_23765,N_23651);
xor U23882 (N_23882,N_23745,N_23728);
nand U23883 (N_23883,N_23764,N_23687);
and U23884 (N_23884,N_23657,N_23721);
nor U23885 (N_23885,N_23658,N_23639);
xor U23886 (N_23886,N_23719,N_23673);
and U23887 (N_23887,N_23671,N_23691);
and U23888 (N_23888,N_23772,N_23609);
xor U23889 (N_23889,N_23684,N_23666);
xnor U23890 (N_23890,N_23625,N_23647);
and U23891 (N_23891,N_23629,N_23712);
xor U23892 (N_23892,N_23702,N_23734);
nand U23893 (N_23893,N_23746,N_23794);
or U23894 (N_23894,N_23642,N_23612);
and U23895 (N_23895,N_23689,N_23701);
nand U23896 (N_23896,N_23770,N_23717);
or U23897 (N_23897,N_23640,N_23776);
or U23898 (N_23898,N_23668,N_23675);
nor U23899 (N_23899,N_23694,N_23606);
xor U23900 (N_23900,N_23790,N_23786);
and U23901 (N_23901,N_23640,N_23732);
and U23902 (N_23902,N_23782,N_23768);
xor U23903 (N_23903,N_23770,N_23711);
nand U23904 (N_23904,N_23749,N_23724);
or U23905 (N_23905,N_23721,N_23716);
nand U23906 (N_23906,N_23748,N_23631);
and U23907 (N_23907,N_23699,N_23652);
or U23908 (N_23908,N_23746,N_23775);
and U23909 (N_23909,N_23764,N_23679);
nor U23910 (N_23910,N_23732,N_23720);
nor U23911 (N_23911,N_23665,N_23743);
or U23912 (N_23912,N_23729,N_23675);
nor U23913 (N_23913,N_23748,N_23613);
or U23914 (N_23914,N_23607,N_23675);
xnor U23915 (N_23915,N_23686,N_23791);
or U23916 (N_23916,N_23634,N_23668);
xor U23917 (N_23917,N_23735,N_23601);
xor U23918 (N_23918,N_23762,N_23752);
nand U23919 (N_23919,N_23778,N_23690);
xnor U23920 (N_23920,N_23725,N_23645);
or U23921 (N_23921,N_23665,N_23765);
nand U23922 (N_23922,N_23614,N_23615);
nand U23923 (N_23923,N_23755,N_23614);
nand U23924 (N_23924,N_23663,N_23612);
nor U23925 (N_23925,N_23733,N_23778);
nor U23926 (N_23926,N_23718,N_23685);
or U23927 (N_23927,N_23686,N_23712);
and U23928 (N_23928,N_23646,N_23747);
nor U23929 (N_23929,N_23679,N_23681);
and U23930 (N_23930,N_23610,N_23663);
or U23931 (N_23931,N_23620,N_23610);
xnor U23932 (N_23932,N_23630,N_23627);
and U23933 (N_23933,N_23777,N_23673);
nand U23934 (N_23934,N_23654,N_23734);
or U23935 (N_23935,N_23715,N_23649);
or U23936 (N_23936,N_23717,N_23790);
xnor U23937 (N_23937,N_23640,N_23629);
nand U23938 (N_23938,N_23783,N_23741);
or U23939 (N_23939,N_23699,N_23795);
nand U23940 (N_23940,N_23689,N_23777);
nor U23941 (N_23941,N_23783,N_23719);
nor U23942 (N_23942,N_23692,N_23686);
or U23943 (N_23943,N_23651,N_23630);
xor U23944 (N_23944,N_23605,N_23604);
nor U23945 (N_23945,N_23692,N_23691);
nand U23946 (N_23946,N_23772,N_23765);
and U23947 (N_23947,N_23797,N_23774);
xor U23948 (N_23948,N_23741,N_23601);
xor U23949 (N_23949,N_23713,N_23732);
or U23950 (N_23950,N_23680,N_23726);
nand U23951 (N_23951,N_23635,N_23753);
nand U23952 (N_23952,N_23616,N_23720);
and U23953 (N_23953,N_23759,N_23687);
or U23954 (N_23954,N_23640,N_23674);
and U23955 (N_23955,N_23669,N_23751);
xnor U23956 (N_23956,N_23681,N_23721);
and U23957 (N_23957,N_23793,N_23626);
xor U23958 (N_23958,N_23768,N_23607);
and U23959 (N_23959,N_23744,N_23644);
nor U23960 (N_23960,N_23755,N_23624);
or U23961 (N_23961,N_23712,N_23623);
or U23962 (N_23962,N_23622,N_23682);
nand U23963 (N_23963,N_23688,N_23709);
xor U23964 (N_23964,N_23735,N_23701);
and U23965 (N_23965,N_23646,N_23681);
and U23966 (N_23966,N_23602,N_23765);
xnor U23967 (N_23967,N_23741,N_23661);
xor U23968 (N_23968,N_23625,N_23740);
nand U23969 (N_23969,N_23784,N_23639);
nor U23970 (N_23970,N_23782,N_23714);
nor U23971 (N_23971,N_23611,N_23794);
xor U23972 (N_23972,N_23660,N_23779);
nor U23973 (N_23973,N_23748,N_23755);
and U23974 (N_23974,N_23719,N_23620);
nor U23975 (N_23975,N_23703,N_23772);
nand U23976 (N_23976,N_23608,N_23667);
nor U23977 (N_23977,N_23731,N_23638);
and U23978 (N_23978,N_23776,N_23748);
nor U23979 (N_23979,N_23730,N_23667);
or U23980 (N_23980,N_23706,N_23708);
nand U23981 (N_23981,N_23692,N_23618);
nor U23982 (N_23982,N_23782,N_23622);
or U23983 (N_23983,N_23630,N_23716);
xnor U23984 (N_23984,N_23772,N_23732);
nor U23985 (N_23985,N_23720,N_23768);
and U23986 (N_23986,N_23718,N_23735);
nand U23987 (N_23987,N_23764,N_23782);
xnor U23988 (N_23988,N_23674,N_23713);
and U23989 (N_23989,N_23751,N_23613);
and U23990 (N_23990,N_23602,N_23673);
nand U23991 (N_23991,N_23610,N_23774);
nor U23992 (N_23992,N_23773,N_23747);
nor U23993 (N_23993,N_23799,N_23782);
xnor U23994 (N_23994,N_23798,N_23707);
nor U23995 (N_23995,N_23746,N_23657);
and U23996 (N_23996,N_23693,N_23628);
nand U23997 (N_23997,N_23674,N_23687);
xnor U23998 (N_23998,N_23707,N_23659);
nand U23999 (N_23999,N_23716,N_23683);
nor U24000 (N_24000,N_23842,N_23922);
or U24001 (N_24001,N_23830,N_23865);
and U24002 (N_24002,N_23827,N_23876);
xnor U24003 (N_24003,N_23879,N_23805);
and U24004 (N_24004,N_23951,N_23974);
xnor U24005 (N_24005,N_23993,N_23980);
xnor U24006 (N_24006,N_23819,N_23913);
and U24007 (N_24007,N_23952,N_23933);
and U24008 (N_24008,N_23983,N_23941);
nor U24009 (N_24009,N_23950,N_23943);
and U24010 (N_24010,N_23874,N_23918);
xor U24011 (N_24011,N_23978,N_23906);
xnor U24012 (N_24012,N_23972,N_23853);
nor U24013 (N_24013,N_23889,N_23878);
or U24014 (N_24014,N_23982,N_23945);
and U24015 (N_24015,N_23901,N_23985);
xnor U24016 (N_24016,N_23953,N_23811);
nor U24017 (N_24017,N_23871,N_23802);
nor U24018 (N_24018,N_23939,N_23908);
and U24019 (N_24019,N_23931,N_23815);
or U24020 (N_24020,N_23897,N_23988);
xor U24021 (N_24021,N_23895,N_23991);
nand U24022 (N_24022,N_23930,N_23834);
nor U24023 (N_24023,N_23904,N_23898);
nor U24024 (N_24024,N_23817,N_23832);
nor U24025 (N_24025,N_23979,N_23888);
xnor U24026 (N_24026,N_23856,N_23997);
nand U24027 (N_24027,N_23996,N_23810);
nor U24028 (N_24028,N_23812,N_23860);
and U24029 (N_24029,N_23965,N_23806);
xnor U24030 (N_24030,N_23934,N_23923);
nor U24031 (N_24031,N_23958,N_23970);
or U24032 (N_24032,N_23893,N_23851);
nand U24033 (N_24033,N_23900,N_23818);
nand U24034 (N_24034,N_23959,N_23870);
nand U24035 (N_24035,N_23938,N_23971);
and U24036 (N_24036,N_23854,N_23875);
nand U24037 (N_24037,N_23986,N_23956);
nor U24038 (N_24038,N_23896,N_23846);
xor U24039 (N_24039,N_23847,N_23859);
nor U24040 (N_24040,N_23902,N_23845);
nor U24041 (N_24041,N_23837,N_23987);
and U24042 (N_24042,N_23891,N_23883);
xnor U24043 (N_24043,N_23981,N_23861);
and U24044 (N_24044,N_23814,N_23995);
nand U24045 (N_24045,N_23866,N_23964);
nand U24046 (N_24046,N_23816,N_23867);
nand U24047 (N_24047,N_23820,N_23844);
nor U24048 (N_24048,N_23916,N_23882);
xnor U24049 (N_24049,N_23935,N_23937);
nor U24050 (N_24050,N_23989,N_23977);
and U24051 (N_24051,N_23961,N_23914);
and U24052 (N_24052,N_23915,N_23831);
xor U24053 (N_24053,N_23966,N_23886);
nor U24054 (N_24054,N_23942,N_23926);
and U24055 (N_24055,N_23957,N_23940);
nor U24056 (N_24056,N_23919,N_23881);
nand U24057 (N_24057,N_23849,N_23969);
or U24058 (N_24058,N_23928,N_23821);
and U24059 (N_24059,N_23903,N_23858);
nor U24060 (N_24060,N_23864,N_23976);
and U24061 (N_24061,N_23839,N_23909);
nor U24062 (N_24062,N_23949,N_23826);
or U24063 (N_24063,N_23925,N_23809);
and U24064 (N_24064,N_23868,N_23803);
nor U24065 (N_24065,N_23999,N_23968);
nor U24066 (N_24066,N_23828,N_23973);
nand U24067 (N_24067,N_23823,N_23850);
or U24068 (N_24068,N_23960,N_23822);
and U24069 (N_24069,N_23843,N_23840);
or U24070 (N_24070,N_23998,N_23899);
xnor U24071 (N_24071,N_23836,N_23824);
or U24072 (N_24072,N_23929,N_23833);
xnor U24073 (N_24073,N_23841,N_23808);
nand U24074 (N_24074,N_23863,N_23825);
and U24075 (N_24075,N_23954,N_23800);
nor U24076 (N_24076,N_23920,N_23807);
nand U24077 (N_24077,N_23990,N_23912);
nand U24078 (N_24078,N_23801,N_23877);
nor U24079 (N_24079,N_23921,N_23887);
or U24080 (N_24080,N_23944,N_23890);
or U24081 (N_24081,N_23936,N_23975);
and U24082 (N_24082,N_23905,N_23862);
nor U24083 (N_24083,N_23955,N_23804);
xnor U24084 (N_24084,N_23835,N_23857);
or U24085 (N_24085,N_23994,N_23869);
and U24086 (N_24086,N_23917,N_23884);
nand U24087 (N_24087,N_23872,N_23829);
nor U24088 (N_24088,N_23992,N_23946);
or U24089 (N_24089,N_23907,N_23984);
nor U24090 (N_24090,N_23892,N_23967);
xnor U24091 (N_24091,N_23911,N_23962);
or U24092 (N_24092,N_23813,N_23838);
xor U24093 (N_24093,N_23910,N_23885);
xor U24094 (N_24094,N_23852,N_23947);
xor U24095 (N_24095,N_23948,N_23873);
nand U24096 (N_24096,N_23927,N_23848);
and U24097 (N_24097,N_23880,N_23855);
nand U24098 (N_24098,N_23963,N_23924);
nand U24099 (N_24099,N_23932,N_23894);
or U24100 (N_24100,N_23897,N_23942);
or U24101 (N_24101,N_23961,N_23973);
nand U24102 (N_24102,N_23946,N_23803);
and U24103 (N_24103,N_23931,N_23975);
xnor U24104 (N_24104,N_23960,N_23873);
or U24105 (N_24105,N_23830,N_23823);
xor U24106 (N_24106,N_23978,N_23803);
nand U24107 (N_24107,N_23841,N_23989);
or U24108 (N_24108,N_23990,N_23891);
or U24109 (N_24109,N_23888,N_23915);
or U24110 (N_24110,N_23997,N_23978);
or U24111 (N_24111,N_23918,N_23860);
or U24112 (N_24112,N_23933,N_23912);
or U24113 (N_24113,N_23857,N_23950);
nor U24114 (N_24114,N_23948,N_23874);
and U24115 (N_24115,N_23882,N_23863);
or U24116 (N_24116,N_23915,N_23895);
xor U24117 (N_24117,N_23971,N_23952);
nor U24118 (N_24118,N_23880,N_23885);
xor U24119 (N_24119,N_23951,N_23837);
nor U24120 (N_24120,N_23987,N_23850);
nand U24121 (N_24121,N_23932,N_23863);
and U24122 (N_24122,N_23877,N_23916);
or U24123 (N_24123,N_23973,N_23890);
nor U24124 (N_24124,N_23970,N_23830);
nor U24125 (N_24125,N_23946,N_23841);
xor U24126 (N_24126,N_23855,N_23908);
nor U24127 (N_24127,N_23946,N_23822);
or U24128 (N_24128,N_23968,N_23996);
and U24129 (N_24129,N_23823,N_23914);
or U24130 (N_24130,N_23864,N_23952);
or U24131 (N_24131,N_23874,N_23914);
nand U24132 (N_24132,N_23838,N_23946);
nor U24133 (N_24133,N_23873,N_23986);
and U24134 (N_24134,N_23862,N_23867);
or U24135 (N_24135,N_23987,N_23890);
nor U24136 (N_24136,N_23995,N_23858);
nor U24137 (N_24137,N_23970,N_23976);
xnor U24138 (N_24138,N_23983,N_23845);
and U24139 (N_24139,N_23898,N_23863);
nor U24140 (N_24140,N_23879,N_23987);
nand U24141 (N_24141,N_23972,N_23881);
nor U24142 (N_24142,N_23909,N_23954);
or U24143 (N_24143,N_23972,N_23963);
and U24144 (N_24144,N_23809,N_23969);
nor U24145 (N_24145,N_23901,N_23957);
or U24146 (N_24146,N_23853,N_23862);
nor U24147 (N_24147,N_23856,N_23806);
nand U24148 (N_24148,N_23841,N_23953);
or U24149 (N_24149,N_23832,N_23863);
and U24150 (N_24150,N_23981,N_23937);
or U24151 (N_24151,N_23977,N_23953);
or U24152 (N_24152,N_23873,N_23864);
nor U24153 (N_24153,N_23867,N_23941);
nand U24154 (N_24154,N_23986,N_23857);
nand U24155 (N_24155,N_23855,N_23941);
nor U24156 (N_24156,N_23817,N_23976);
or U24157 (N_24157,N_23963,N_23964);
xor U24158 (N_24158,N_23869,N_23968);
xnor U24159 (N_24159,N_23934,N_23822);
xnor U24160 (N_24160,N_23873,N_23814);
xor U24161 (N_24161,N_23987,N_23824);
and U24162 (N_24162,N_23902,N_23808);
nand U24163 (N_24163,N_23886,N_23963);
nand U24164 (N_24164,N_23856,N_23904);
or U24165 (N_24165,N_23869,N_23912);
and U24166 (N_24166,N_23863,N_23857);
and U24167 (N_24167,N_23840,N_23878);
and U24168 (N_24168,N_23928,N_23886);
nor U24169 (N_24169,N_23993,N_23970);
xor U24170 (N_24170,N_23884,N_23939);
nor U24171 (N_24171,N_23932,N_23998);
and U24172 (N_24172,N_23806,N_23813);
nand U24173 (N_24173,N_23948,N_23882);
or U24174 (N_24174,N_23862,N_23959);
xnor U24175 (N_24175,N_23859,N_23990);
nand U24176 (N_24176,N_23867,N_23817);
nand U24177 (N_24177,N_23964,N_23971);
nor U24178 (N_24178,N_23849,N_23800);
or U24179 (N_24179,N_23999,N_23827);
xnor U24180 (N_24180,N_23938,N_23855);
or U24181 (N_24181,N_23943,N_23897);
xor U24182 (N_24182,N_23813,N_23902);
or U24183 (N_24183,N_23821,N_23939);
nand U24184 (N_24184,N_23960,N_23852);
nor U24185 (N_24185,N_23914,N_23819);
and U24186 (N_24186,N_23801,N_23883);
or U24187 (N_24187,N_23949,N_23870);
nor U24188 (N_24188,N_23995,N_23877);
or U24189 (N_24189,N_23924,N_23821);
xnor U24190 (N_24190,N_23837,N_23942);
nor U24191 (N_24191,N_23993,N_23923);
or U24192 (N_24192,N_23824,N_23920);
or U24193 (N_24193,N_23872,N_23965);
nand U24194 (N_24194,N_23947,N_23944);
or U24195 (N_24195,N_23923,N_23959);
or U24196 (N_24196,N_23876,N_23995);
and U24197 (N_24197,N_23965,N_23973);
nor U24198 (N_24198,N_23802,N_23820);
nor U24199 (N_24199,N_23840,N_23866);
xor U24200 (N_24200,N_24118,N_24074);
nand U24201 (N_24201,N_24002,N_24007);
nand U24202 (N_24202,N_24167,N_24183);
xnor U24203 (N_24203,N_24000,N_24116);
nor U24204 (N_24204,N_24149,N_24108);
or U24205 (N_24205,N_24162,N_24196);
nand U24206 (N_24206,N_24058,N_24190);
nand U24207 (N_24207,N_24168,N_24180);
xnor U24208 (N_24208,N_24052,N_24071);
and U24209 (N_24209,N_24103,N_24156);
nor U24210 (N_24210,N_24101,N_24137);
xnor U24211 (N_24211,N_24176,N_24115);
nor U24212 (N_24212,N_24131,N_24062);
nor U24213 (N_24213,N_24159,N_24066);
nand U24214 (N_24214,N_24135,N_24197);
nor U24215 (N_24215,N_24076,N_24102);
or U24216 (N_24216,N_24037,N_24179);
and U24217 (N_24217,N_24175,N_24029);
and U24218 (N_24218,N_24125,N_24038);
nand U24219 (N_24219,N_24155,N_24048);
nand U24220 (N_24220,N_24046,N_24113);
and U24221 (N_24221,N_24051,N_24041);
or U24222 (N_24222,N_24077,N_24078);
nand U24223 (N_24223,N_24054,N_24154);
and U24224 (N_24224,N_24033,N_24130);
or U24225 (N_24225,N_24065,N_24042);
or U24226 (N_24226,N_24148,N_24129);
and U24227 (N_24227,N_24133,N_24043);
or U24228 (N_24228,N_24006,N_24163);
or U24229 (N_24229,N_24080,N_24186);
and U24230 (N_24230,N_24015,N_24126);
nor U24231 (N_24231,N_24067,N_24121);
nor U24232 (N_24232,N_24050,N_24164);
nor U24233 (N_24233,N_24172,N_24084);
nand U24234 (N_24234,N_24056,N_24112);
xor U24235 (N_24235,N_24193,N_24194);
xnor U24236 (N_24236,N_24057,N_24093);
or U24237 (N_24237,N_24089,N_24017);
nor U24238 (N_24238,N_24107,N_24012);
and U24239 (N_24239,N_24117,N_24001);
nand U24240 (N_24240,N_24110,N_24082);
xor U24241 (N_24241,N_24146,N_24140);
or U24242 (N_24242,N_24086,N_24034);
nor U24243 (N_24243,N_24192,N_24171);
and U24244 (N_24244,N_24153,N_24095);
nand U24245 (N_24245,N_24100,N_24063);
or U24246 (N_24246,N_24022,N_24147);
xor U24247 (N_24247,N_24036,N_24096);
nand U24248 (N_24248,N_24011,N_24173);
or U24249 (N_24249,N_24128,N_24106);
or U24250 (N_24250,N_24143,N_24024);
nor U24251 (N_24251,N_24184,N_24008);
or U24252 (N_24252,N_24144,N_24139);
and U24253 (N_24253,N_24031,N_24187);
or U24254 (N_24254,N_24141,N_24127);
and U24255 (N_24255,N_24152,N_24088);
nor U24256 (N_24256,N_24181,N_24075);
or U24257 (N_24257,N_24014,N_24157);
nand U24258 (N_24258,N_24018,N_24070);
nand U24259 (N_24259,N_24045,N_24114);
nand U24260 (N_24260,N_24005,N_24069);
nor U24261 (N_24261,N_24142,N_24049);
xor U24262 (N_24262,N_24027,N_24013);
or U24263 (N_24263,N_24111,N_24132);
nand U24264 (N_24264,N_24123,N_24169);
nor U24265 (N_24265,N_24195,N_24039);
or U24266 (N_24266,N_24019,N_24160);
nor U24267 (N_24267,N_24028,N_24090);
nor U24268 (N_24268,N_24053,N_24004);
xor U24269 (N_24269,N_24003,N_24174);
nand U24270 (N_24270,N_24191,N_24023);
and U24271 (N_24271,N_24161,N_24104);
xnor U24272 (N_24272,N_24055,N_24145);
or U24273 (N_24273,N_24060,N_24094);
nand U24274 (N_24274,N_24120,N_24064);
or U24275 (N_24275,N_24061,N_24040);
or U24276 (N_24276,N_24030,N_24189);
nand U24277 (N_24277,N_24124,N_24177);
nor U24278 (N_24278,N_24009,N_24119);
nor U24279 (N_24279,N_24170,N_24035);
and U24280 (N_24280,N_24150,N_24092);
or U24281 (N_24281,N_24109,N_24091);
nor U24282 (N_24282,N_24026,N_24032);
nor U24283 (N_24283,N_24068,N_24136);
nor U24284 (N_24284,N_24165,N_24098);
or U24285 (N_24285,N_24020,N_24105);
xnor U24286 (N_24286,N_24182,N_24021);
or U24287 (N_24287,N_24158,N_24185);
nand U24288 (N_24288,N_24010,N_24166);
xnor U24289 (N_24289,N_24097,N_24199);
and U24290 (N_24290,N_24025,N_24083);
or U24291 (N_24291,N_24122,N_24188);
nand U24292 (N_24292,N_24016,N_24198);
xnor U24293 (N_24293,N_24073,N_24134);
and U24294 (N_24294,N_24079,N_24081);
nand U24295 (N_24295,N_24087,N_24178);
or U24296 (N_24296,N_24151,N_24059);
or U24297 (N_24297,N_24099,N_24044);
nor U24298 (N_24298,N_24138,N_24085);
or U24299 (N_24299,N_24072,N_24047);
or U24300 (N_24300,N_24005,N_24042);
nand U24301 (N_24301,N_24172,N_24076);
and U24302 (N_24302,N_24100,N_24074);
and U24303 (N_24303,N_24191,N_24144);
nor U24304 (N_24304,N_24052,N_24190);
nand U24305 (N_24305,N_24189,N_24085);
nand U24306 (N_24306,N_24097,N_24144);
nand U24307 (N_24307,N_24174,N_24134);
xnor U24308 (N_24308,N_24134,N_24192);
nand U24309 (N_24309,N_24192,N_24035);
nor U24310 (N_24310,N_24197,N_24167);
or U24311 (N_24311,N_24080,N_24139);
xnor U24312 (N_24312,N_24144,N_24031);
nand U24313 (N_24313,N_24042,N_24070);
and U24314 (N_24314,N_24081,N_24069);
and U24315 (N_24315,N_24008,N_24171);
nor U24316 (N_24316,N_24087,N_24007);
or U24317 (N_24317,N_24170,N_24137);
xor U24318 (N_24318,N_24106,N_24049);
xnor U24319 (N_24319,N_24144,N_24054);
nor U24320 (N_24320,N_24072,N_24197);
or U24321 (N_24321,N_24092,N_24199);
nand U24322 (N_24322,N_24115,N_24178);
xor U24323 (N_24323,N_24177,N_24192);
nand U24324 (N_24324,N_24164,N_24102);
and U24325 (N_24325,N_24018,N_24123);
nor U24326 (N_24326,N_24062,N_24182);
nand U24327 (N_24327,N_24077,N_24150);
nand U24328 (N_24328,N_24196,N_24141);
nor U24329 (N_24329,N_24102,N_24130);
or U24330 (N_24330,N_24150,N_24046);
and U24331 (N_24331,N_24102,N_24055);
nand U24332 (N_24332,N_24167,N_24137);
nor U24333 (N_24333,N_24192,N_24142);
nor U24334 (N_24334,N_24162,N_24139);
xor U24335 (N_24335,N_24036,N_24175);
and U24336 (N_24336,N_24024,N_24078);
or U24337 (N_24337,N_24197,N_24119);
nor U24338 (N_24338,N_24095,N_24100);
nand U24339 (N_24339,N_24002,N_24155);
or U24340 (N_24340,N_24149,N_24034);
or U24341 (N_24341,N_24094,N_24110);
xnor U24342 (N_24342,N_24116,N_24044);
nor U24343 (N_24343,N_24027,N_24195);
and U24344 (N_24344,N_24085,N_24071);
or U24345 (N_24345,N_24167,N_24194);
nor U24346 (N_24346,N_24044,N_24125);
xnor U24347 (N_24347,N_24166,N_24144);
and U24348 (N_24348,N_24059,N_24166);
xnor U24349 (N_24349,N_24150,N_24175);
nor U24350 (N_24350,N_24197,N_24099);
or U24351 (N_24351,N_24012,N_24198);
nand U24352 (N_24352,N_24145,N_24188);
xor U24353 (N_24353,N_24197,N_24106);
xor U24354 (N_24354,N_24118,N_24189);
or U24355 (N_24355,N_24194,N_24144);
or U24356 (N_24356,N_24070,N_24121);
xnor U24357 (N_24357,N_24088,N_24132);
xor U24358 (N_24358,N_24054,N_24001);
or U24359 (N_24359,N_24142,N_24124);
nand U24360 (N_24360,N_24055,N_24027);
or U24361 (N_24361,N_24055,N_24127);
nand U24362 (N_24362,N_24123,N_24009);
nor U24363 (N_24363,N_24004,N_24133);
xnor U24364 (N_24364,N_24138,N_24129);
or U24365 (N_24365,N_24056,N_24073);
nand U24366 (N_24366,N_24035,N_24106);
nand U24367 (N_24367,N_24153,N_24029);
or U24368 (N_24368,N_24124,N_24083);
nand U24369 (N_24369,N_24040,N_24142);
nor U24370 (N_24370,N_24012,N_24090);
xnor U24371 (N_24371,N_24023,N_24084);
nand U24372 (N_24372,N_24155,N_24102);
and U24373 (N_24373,N_24044,N_24091);
nand U24374 (N_24374,N_24145,N_24091);
nand U24375 (N_24375,N_24084,N_24146);
nand U24376 (N_24376,N_24121,N_24032);
nand U24377 (N_24377,N_24193,N_24111);
and U24378 (N_24378,N_24031,N_24081);
xnor U24379 (N_24379,N_24077,N_24126);
or U24380 (N_24380,N_24087,N_24096);
or U24381 (N_24381,N_24107,N_24076);
nor U24382 (N_24382,N_24051,N_24111);
or U24383 (N_24383,N_24064,N_24026);
xor U24384 (N_24384,N_24038,N_24093);
and U24385 (N_24385,N_24051,N_24073);
nand U24386 (N_24386,N_24188,N_24052);
xnor U24387 (N_24387,N_24043,N_24107);
or U24388 (N_24388,N_24059,N_24163);
xnor U24389 (N_24389,N_24046,N_24050);
nor U24390 (N_24390,N_24111,N_24120);
nor U24391 (N_24391,N_24149,N_24028);
or U24392 (N_24392,N_24052,N_24045);
nand U24393 (N_24393,N_24091,N_24154);
and U24394 (N_24394,N_24010,N_24137);
or U24395 (N_24395,N_24189,N_24049);
nor U24396 (N_24396,N_24176,N_24013);
nor U24397 (N_24397,N_24017,N_24092);
nand U24398 (N_24398,N_24101,N_24146);
and U24399 (N_24399,N_24011,N_24050);
xor U24400 (N_24400,N_24359,N_24297);
and U24401 (N_24401,N_24356,N_24315);
and U24402 (N_24402,N_24296,N_24234);
nand U24403 (N_24403,N_24345,N_24266);
nor U24404 (N_24404,N_24303,N_24369);
xor U24405 (N_24405,N_24244,N_24260);
or U24406 (N_24406,N_24256,N_24295);
xnor U24407 (N_24407,N_24222,N_24311);
and U24408 (N_24408,N_24226,N_24304);
nand U24409 (N_24409,N_24219,N_24211);
xor U24410 (N_24410,N_24380,N_24354);
and U24411 (N_24411,N_24374,N_24362);
nor U24412 (N_24412,N_24341,N_24202);
or U24413 (N_24413,N_24320,N_24262);
or U24414 (N_24414,N_24257,N_24300);
xnor U24415 (N_24415,N_24399,N_24265);
and U24416 (N_24416,N_24241,N_24224);
xnor U24417 (N_24417,N_24355,N_24287);
nor U24418 (N_24418,N_24316,N_24324);
nor U24419 (N_24419,N_24358,N_24213);
nor U24420 (N_24420,N_24288,N_24302);
nand U24421 (N_24421,N_24272,N_24207);
nor U24422 (N_24422,N_24323,N_24333);
or U24423 (N_24423,N_24391,N_24235);
xor U24424 (N_24424,N_24377,N_24229);
nor U24425 (N_24425,N_24238,N_24363);
nand U24426 (N_24426,N_24239,N_24318);
and U24427 (N_24427,N_24210,N_24314);
xor U24428 (N_24428,N_24353,N_24385);
nor U24429 (N_24429,N_24331,N_24278);
nand U24430 (N_24430,N_24309,N_24276);
xor U24431 (N_24431,N_24291,N_24338);
xor U24432 (N_24432,N_24299,N_24242);
nand U24433 (N_24433,N_24236,N_24357);
or U24434 (N_24434,N_24269,N_24387);
and U24435 (N_24435,N_24274,N_24261);
nand U24436 (N_24436,N_24393,N_24306);
and U24437 (N_24437,N_24217,N_24394);
or U24438 (N_24438,N_24371,N_24386);
or U24439 (N_24439,N_24218,N_24398);
nor U24440 (N_24440,N_24372,N_24361);
nor U24441 (N_24441,N_24247,N_24289);
xnor U24442 (N_24442,N_24381,N_24370);
xnor U24443 (N_24443,N_24208,N_24313);
xor U24444 (N_24444,N_24317,N_24347);
nor U24445 (N_24445,N_24263,N_24255);
and U24446 (N_24446,N_24252,N_24365);
nor U24447 (N_24447,N_24204,N_24283);
xor U24448 (N_24448,N_24254,N_24264);
xnor U24449 (N_24449,N_24350,N_24240);
nand U24450 (N_24450,N_24221,N_24366);
nor U24451 (N_24451,N_24308,N_24284);
xor U24452 (N_24452,N_24248,N_24348);
xnor U24453 (N_24453,N_24206,N_24368);
xor U24454 (N_24454,N_24243,N_24389);
and U24455 (N_24455,N_24294,N_24335);
nand U24456 (N_24456,N_24312,N_24349);
or U24457 (N_24457,N_24310,N_24328);
or U24458 (N_24458,N_24258,N_24277);
nand U24459 (N_24459,N_24376,N_24305);
nand U24460 (N_24460,N_24301,N_24205);
xor U24461 (N_24461,N_24200,N_24290);
xnor U24462 (N_24462,N_24351,N_24343);
or U24463 (N_24463,N_24397,N_24327);
nand U24464 (N_24464,N_24228,N_24352);
nand U24465 (N_24465,N_24373,N_24378);
or U24466 (N_24466,N_24279,N_24249);
nand U24467 (N_24467,N_24268,N_24321);
or U24468 (N_24468,N_24326,N_24384);
nor U24469 (N_24469,N_24332,N_24337);
nand U24470 (N_24470,N_24246,N_24360);
xor U24471 (N_24471,N_24325,N_24270);
or U24472 (N_24472,N_24275,N_24367);
xnor U24473 (N_24473,N_24267,N_24285);
xnor U24474 (N_24474,N_24344,N_24280);
and U24475 (N_24475,N_24271,N_24375);
nor U24476 (N_24476,N_24307,N_24216);
nor U24477 (N_24477,N_24383,N_24212);
nor U24478 (N_24478,N_24225,N_24382);
nand U24479 (N_24479,N_24201,N_24339);
nor U24480 (N_24480,N_24364,N_24319);
and U24481 (N_24481,N_24293,N_24379);
nor U24482 (N_24482,N_24388,N_24340);
and U24483 (N_24483,N_24220,N_24203);
nor U24484 (N_24484,N_24251,N_24227);
or U24485 (N_24485,N_24253,N_24209);
xor U24486 (N_24486,N_24231,N_24342);
nand U24487 (N_24487,N_24215,N_24346);
xor U24488 (N_24488,N_24330,N_24273);
xnor U24489 (N_24489,N_24396,N_24298);
nand U24490 (N_24490,N_24223,N_24282);
xor U24491 (N_24491,N_24392,N_24329);
nand U24492 (N_24492,N_24250,N_24233);
nand U24493 (N_24493,N_24336,N_24292);
and U24494 (N_24494,N_24259,N_24281);
nor U24495 (N_24495,N_24232,N_24237);
nand U24496 (N_24496,N_24322,N_24390);
nand U24497 (N_24497,N_24214,N_24230);
and U24498 (N_24498,N_24334,N_24395);
and U24499 (N_24499,N_24286,N_24245);
or U24500 (N_24500,N_24391,N_24361);
nand U24501 (N_24501,N_24319,N_24374);
or U24502 (N_24502,N_24390,N_24281);
nor U24503 (N_24503,N_24317,N_24375);
nand U24504 (N_24504,N_24219,N_24212);
nor U24505 (N_24505,N_24319,N_24394);
or U24506 (N_24506,N_24262,N_24346);
and U24507 (N_24507,N_24397,N_24227);
and U24508 (N_24508,N_24308,N_24259);
nand U24509 (N_24509,N_24274,N_24305);
xnor U24510 (N_24510,N_24295,N_24369);
xor U24511 (N_24511,N_24204,N_24337);
and U24512 (N_24512,N_24380,N_24375);
or U24513 (N_24513,N_24256,N_24389);
and U24514 (N_24514,N_24329,N_24236);
or U24515 (N_24515,N_24283,N_24261);
or U24516 (N_24516,N_24206,N_24341);
nand U24517 (N_24517,N_24303,N_24347);
nand U24518 (N_24518,N_24231,N_24285);
or U24519 (N_24519,N_24305,N_24344);
xnor U24520 (N_24520,N_24269,N_24367);
and U24521 (N_24521,N_24234,N_24246);
xnor U24522 (N_24522,N_24397,N_24263);
nand U24523 (N_24523,N_24244,N_24356);
and U24524 (N_24524,N_24363,N_24330);
nor U24525 (N_24525,N_24279,N_24393);
xor U24526 (N_24526,N_24264,N_24292);
nor U24527 (N_24527,N_24273,N_24347);
or U24528 (N_24528,N_24270,N_24262);
nor U24529 (N_24529,N_24335,N_24281);
nand U24530 (N_24530,N_24357,N_24286);
xor U24531 (N_24531,N_24202,N_24321);
nor U24532 (N_24532,N_24318,N_24283);
or U24533 (N_24533,N_24279,N_24334);
nor U24534 (N_24534,N_24312,N_24286);
nand U24535 (N_24535,N_24222,N_24383);
nor U24536 (N_24536,N_24311,N_24205);
or U24537 (N_24537,N_24274,N_24285);
and U24538 (N_24538,N_24277,N_24290);
and U24539 (N_24539,N_24229,N_24372);
nor U24540 (N_24540,N_24246,N_24267);
xor U24541 (N_24541,N_24240,N_24267);
and U24542 (N_24542,N_24331,N_24234);
or U24543 (N_24543,N_24287,N_24386);
nand U24544 (N_24544,N_24337,N_24290);
nor U24545 (N_24545,N_24348,N_24271);
xor U24546 (N_24546,N_24288,N_24251);
nand U24547 (N_24547,N_24317,N_24271);
nand U24548 (N_24548,N_24237,N_24349);
or U24549 (N_24549,N_24210,N_24260);
and U24550 (N_24550,N_24345,N_24303);
nor U24551 (N_24551,N_24210,N_24262);
or U24552 (N_24552,N_24269,N_24282);
and U24553 (N_24553,N_24239,N_24202);
nand U24554 (N_24554,N_24362,N_24243);
or U24555 (N_24555,N_24318,N_24315);
nand U24556 (N_24556,N_24278,N_24363);
xnor U24557 (N_24557,N_24310,N_24248);
and U24558 (N_24558,N_24227,N_24264);
or U24559 (N_24559,N_24270,N_24370);
nor U24560 (N_24560,N_24383,N_24328);
and U24561 (N_24561,N_24245,N_24273);
nor U24562 (N_24562,N_24269,N_24398);
or U24563 (N_24563,N_24307,N_24399);
xor U24564 (N_24564,N_24327,N_24218);
xnor U24565 (N_24565,N_24390,N_24313);
nor U24566 (N_24566,N_24345,N_24204);
or U24567 (N_24567,N_24375,N_24388);
xnor U24568 (N_24568,N_24249,N_24287);
nor U24569 (N_24569,N_24344,N_24386);
or U24570 (N_24570,N_24278,N_24262);
and U24571 (N_24571,N_24269,N_24246);
nand U24572 (N_24572,N_24383,N_24308);
or U24573 (N_24573,N_24351,N_24390);
and U24574 (N_24574,N_24335,N_24230);
or U24575 (N_24575,N_24256,N_24304);
xor U24576 (N_24576,N_24229,N_24239);
or U24577 (N_24577,N_24375,N_24222);
nor U24578 (N_24578,N_24309,N_24255);
nand U24579 (N_24579,N_24259,N_24338);
nor U24580 (N_24580,N_24391,N_24334);
or U24581 (N_24581,N_24300,N_24284);
xnor U24582 (N_24582,N_24207,N_24399);
nor U24583 (N_24583,N_24225,N_24327);
and U24584 (N_24584,N_24288,N_24260);
nor U24585 (N_24585,N_24206,N_24298);
and U24586 (N_24586,N_24239,N_24380);
or U24587 (N_24587,N_24302,N_24392);
nand U24588 (N_24588,N_24255,N_24347);
xor U24589 (N_24589,N_24332,N_24372);
xnor U24590 (N_24590,N_24325,N_24324);
xor U24591 (N_24591,N_24300,N_24341);
and U24592 (N_24592,N_24363,N_24226);
and U24593 (N_24593,N_24247,N_24215);
nor U24594 (N_24594,N_24243,N_24385);
or U24595 (N_24595,N_24372,N_24306);
xnor U24596 (N_24596,N_24372,N_24298);
xor U24597 (N_24597,N_24386,N_24307);
and U24598 (N_24598,N_24215,N_24260);
nor U24599 (N_24599,N_24207,N_24365);
xor U24600 (N_24600,N_24528,N_24561);
nor U24601 (N_24601,N_24404,N_24541);
nor U24602 (N_24602,N_24515,N_24483);
and U24603 (N_24603,N_24580,N_24597);
xnor U24604 (N_24604,N_24574,N_24522);
nand U24605 (N_24605,N_24419,N_24569);
nor U24606 (N_24606,N_24552,N_24583);
nand U24607 (N_24607,N_24544,N_24430);
xor U24608 (N_24608,N_24531,N_24439);
nor U24609 (N_24609,N_24520,N_24494);
or U24610 (N_24610,N_24493,N_24530);
xor U24611 (N_24611,N_24436,N_24434);
nor U24612 (N_24612,N_24405,N_24554);
nor U24613 (N_24613,N_24406,N_24411);
nor U24614 (N_24614,N_24511,N_24464);
or U24615 (N_24615,N_24590,N_24414);
nand U24616 (N_24616,N_24579,N_24563);
or U24617 (N_24617,N_24420,N_24441);
xor U24618 (N_24618,N_24472,N_24507);
nor U24619 (N_24619,N_24413,N_24485);
and U24620 (N_24620,N_24562,N_24467);
and U24621 (N_24621,N_24460,N_24432);
nor U24622 (N_24622,N_24553,N_24598);
nor U24623 (N_24623,N_24538,N_24537);
or U24624 (N_24624,N_24549,N_24500);
or U24625 (N_24625,N_24465,N_24476);
nand U24626 (N_24626,N_24570,N_24463);
or U24627 (N_24627,N_24421,N_24540);
and U24628 (N_24628,N_24581,N_24525);
nand U24629 (N_24629,N_24435,N_24556);
nand U24630 (N_24630,N_24445,N_24499);
nand U24631 (N_24631,N_24521,N_24408);
and U24632 (N_24632,N_24489,N_24546);
xor U24633 (N_24633,N_24438,N_24573);
nor U24634 (N_24634,N_24450,N_24446);
and U24635 (N_24635,N_24442,N_24459);
xor U24636 (N_24636,N_24417,N_24449);
xnor U24637 (N_24637,N_24468,N_24495);
xor U24638 (N_24638,N_24490,N_24422);
or U24639 (N_24639,N_24455,N_24508);
xnor U24640 (N_24640,N_24481,N_24410);
and U24641 (N_24641,N_24416,N_24482);
nor U24642 (N_24642,N_24576,N_24409);
nor U24643 (N_24643,N_24548,N_24512);
and U24644 (N_24644,N_24504,N_24443);
xnor U24645 (N_24645,N_24565,N_24575);
xnor U24646 (N_24646,N_24571,N_24519);
nor U24647 (N_24647,N_24532,N_24545);
xnor U24648 (N_24648,N_24491,N_24539);
xor U24649 (N_24649,N_24526,N_24401);
nor U24650 (N_24650,N_24529,N_24415);
nor U24651 (N_24651,N_24567,N_24524);
xnor U24652 (N_24652,N_24572,N_24437);
nand U24653 (N_24653,N_24424,N_24577);
or U24654 (N_24654,N_24555,N_24558);
nand U24655 (N_24655,N_24550,N_24403);
nand U24656 (N_24656,N_24587,N_24440);
nand U24657 (N_24657,N_24462,N_24543);
nand U24658 (N_24658,N_24518,N_24492);
xor U24659 (N_24659,N_24517,N_24502);
xor U24660 (N_24660,N_24447,N_24503);
and U24661 (N_24661,N_24454,N_24407);
nand U24662 (N_24662,N_24523,N_24470);
nand U24663 (N_24663,N_24444,N_24559);
nor U24664 (N_24664,N_24534,N_24497);
nand U24665 (N_24665,N_24535,N_24480);
nand U24666 (N_24666,N_24400,N_24426);
nor U24667 (N_24667,N_24536,N_24599);
or U24668 (N_24668,N_24479,N_24458);
nand U24669 (N_24669,N_24560,N_24477);
and U24670 (N_24670,N_24501,N_24510);
nand U24671 (N_24671,N_24429,N_24514);
and U24672 (N_24672,N_24473,N_24428);
nor U24673 (N_24673,N_24589,N_24568);
nor U24674 (N_24674,N_24505,N_24427);
and U24675 (N_24675,N_24551,N_24542);
or U24676 (N_24676,N_24461,N_24584);
or U24677 (N_24677,N_24478,N_24498);
or U24678 (N_24678,N_24452,N_24431);
or U24679 (N_24679,N_24469,N_24487);
or U24680 (N_24680,N_24566,N_24547);
or U24681 (N_24681,N_24595,N_24488);
or U24682 (N_24682,N_24527,N_24453);
xnor U24683 (N_24683,N_24582,N_24591);
nor U24684 (N_24684,N_24564,N_24457);
or U24685 (N_24685,N_24516,N_24533);
or U24686 (N_24686,N_24506,N_24448);
and U24687 (N_24687,N_24475,N_24433);
xnor U24688 (N_24688,N_24474,N_24557);
nor U24689 (N_24689,N_24466,N_24471);
nand U24690 (N_24690,N_24412,N_24586);
xnor U24691 (N_24691,N_24513,N_24423);
or U24692 (N_24692,N_24456,N_24496);
and U24693 (N_24693,N_24509,N_24585);
or U24694 (N_24694,N_24402,N_24592);
nand U24695 (N_24695,N_24588,N_24596);
nor U24696 (N_24696,N_24578,N_24593);
and U24697 (N_24697,N_24425,N_24594);
xnor U24698 (N_24698,N_24451,N_24486);
and U24699 (N_24699,N_24484,N_24418);
nand U24700 (N_24700,N_24490,N_24441);
xor U24701 (N_24701,N_24588,N_24428);
nand U24702 (N_24702,N_24507,N_24463);
or U24703 (N_24703,N_24415,N_24580);
or U24704 (N_24704,N_24467,N_24485);
or U24705 (N_24705,N_24579,N_24526);
and U24706 (N_24706,N_24422,N_24413);
xnor U24707 (N_24707,N_24469,N_24450);
nand U24708 (N_24708,N_24500,N_24433);
nand U24709 (N_24709,N_24509,N_24548);
and U24710 (N_24710,N_24563,N_24417);
xor U24711 (N_24711,N_24417,N_24429);
nor U24712 (N_24712,N_24564,N_24542);
nand U24713 (N_24713,N_24590,N_24544);
nand U24714 (N_24714,N_24479,N_24560);
or U24715 (N_24715,N_24547,N_24468);
and U24716 (N_24716,N_24532,N_24453);
or U24717 (N_24717,N_24542,N_24521);
nand U24718 (N_24718,N_24446,N_24493);
and U24719 (N_24719,N_24519,N_24560);
xnor U24720 (N_24720,N_24539,N_24519);
nand U24721 (N_24721,N_24537,N_24455);
nand U24722 (N_24722,N_24428,N_24549);
xnor U24723 (N_24723,N_24594,N_24484);
xnor U24724 (N_24724,N_24597,N_24400);
or U24725 (N_24725,N_24503,N_24540);
nand U24726 (N_24726,N_24548,N_24485);
nand U24727 (N_24727,N_24540,N_24480);
or U24728 (N_24728,N_24431,N_24507);
or U24729 (N_24729,N_24424,N_24510);
nand U24730 (N_24730,N_24480,N_24544);
and U24731 (N_24731,N_24513,N_24449);
xor U24732 (N_24732,N_24568,N_24533);
and U24733 (N_24733,N_24455,N_24485);
and U24734 (N_24734,N_24427,N_24456);
nor U24735 (N_24735,N_24586,N_24471);
and U24736 (N_24736,N_24595,N_24433);
nand U24737 (N_24737,N_24425,N_24448);
or U24738 (N_24738,N_24427,N_24481);
or U24739 (N_24739,N_24427,N_24468);
and U24740 (N_24740,N_24447,N_24581);
xor U24741 (N_24741,N_24549,N_24415);
and U24742 (N_24742,N_24477,N_24490);
xor U24743 (N_24743,N_24594,N_24574);
xnor U24744 (N_24744,N_24538,N_24536);
nand U24745 (N_24745,N_24420,N_24481);
or U24746 (N_24746,N_24561,N_24431);
nor U24747 (N_24747,N_24404,N_24435);
or U24748 (N_24748,N_24526,N_24431);
or U24749 (N_24749,N_24424,N_24584);
and U24750 (N_24750,N_24403,N_24593);
and U24751 (N_24751,N_24494,N_24571);
nor U24752 (N_24752,N_24468,N_24472);
nand U24753 (N_24753,N_24538,N_24489);
xor U24754 (N_24754,N_24545,N_24597);
nor U24755 (N_24755,N_24448,N_24416);
xor U24756 (N_24756,N_24547,N_24531);
or U24757 (N_24757,N_24441,N_24474);
xor U24758 (N_24758,N_24449,N_24593);
nor U24759 (N_24759,N_24485,N_24481);
and U24760 (N_24760,N_24533,N_24448);
or U24761 (N_24761,N_24438,N_24547);
nand U24762 (N_24762,N_24512,N_24599);
or U24763 (N_24763,N_24553,N_24514);
xnor U24764 (N_24764,N_24559,N_24440);
nand U24765 (N_24765,N_24475,N_24518);
xor U24766 (N_24766,N_24534,N_24441);
or U24767 (N_24767,N_24508,N_24543);
and U24768 (N_24768,N_24442,N_24503);
nand U24769 (N_24769,N_24551,N_24476);
nor U24770 (N_24770,N_24576,N_24493);
and U24771 (N_24771,N_24499,N_24567);
xnor U24772 (N_24772,N_24543,N_24456);
nor U24773 (N_24773,N_24521,N_24503);
nand U24774 (N_24774,N_24499,N_24428);
and U24775 (N_24775,N_24486,N_24501);
nand U24776 (N_24776,N_24495,N_24556);
xor U24777 (N_24777,N_24401,N_24436);
and U24778 (N_24778,N_24528,N_24459);
or U24779 (N_24779,N_24518,N_24406);
nor U24780 (N_24780,N_24423,N_24530);
and U24781 (N_24781,N_24412,N_24498);
xor U24782 (N_24782,N_24578,N_24492);
or U24783 (N_24783,N_24546,N_24572);
xor U24784 (N_24784,N_24538,N_24445);
nand U24785 (N_24785,N_24406,N_24587);
nor U24786 (N_24786,N_24411,N_24421);
or U24787 (N_24787,N_24583,N_24579);
or U24788 (N_24788,N_24572,N_24533);
or U24789 (N_24789,N_24431,N_24564);
nor U24790 (N_24790,N_24430,N_24540);
nand U24791 (N_24791,N_24417,N_24565);
xnor U24792 (N_24792,N_24419,N_24530);
nand U24793 (N_24793,N_24543,N_24445);
and U24794 (N_24794,N_24536,N_24491);
and U24795 (N_24795,N_24597,N_24500);
and U24796 (N_24796,N_24420,N_24439);
nor U24797 (N_24797,N_24515,N_24405);
and U24798 (N_24798,N_24594,N_24427);
or U24799 (N_24799,N_24450,N_24436);
nor U24800 (N_24800,N_24776,N_24627);
and U24801 (N_24801,N_24783,N_24615);
and U24802 (N_24802,N_24605,N_24764);
nand U24803 (N_24803,N_24721,N_24749);
or U24804 (N_24804,N_24667,N_24723);
nand U24805 (N_24805,N_24790,N_24659);
or U24806 (N_24806,N_24628,N_24739);
and U24807 (N_24807,N_24606,N_24611);
nor U24808 (N_24808,N_24738,N_24710);
nor U24809 (N_24809,N_24734,N_24758);
and U24810 (N_24810,N_24674,N_24663);
xor U24811 (N_24811,N_24745,N_24711);
xor U24812 (N_24812,N_24795,N_24625);
nand U24813 (N_24813,N_24716,N_24696);
nand U24814 (N_24814,N_24765,N_24770);
xnor U24815 (N_24815,N_24698,N_24692);
and U24816 (N_24816,N_24702,N_24632);
nand U24817 (N_24817,N_24693,N_24649);
nor U24818 (N_24818,N_24751,N_24630);
nand U24819 (N_24819,N_24680,N_24747);
and U24820 (N_24820,N_24728,N_24791);
and U24821 (N_24821,N_24784,N_24601);
or U24822 (N_24822,N_24631,N_24638);
or U24823 (N_24823,N_24613,N_24757);
or U24824 (N_24824,N_24695,N_24699);
or U24825 (N_24825,N_24731,N_24707);
xor U24826 (N_24826,N_24662,N_24660);
and U24827 (N_24827,N_24727,N_24740);
xor U24828 (N_24828,N_24742,N_24704);
and U24829 (N_24829,N_24655,N_24717);
nand U24830 (N_24830,N_24665,N_24733);
nor U24831 (N_24831,N_24610,N_24619);
nor U24832 (N_24832,N_24639,N_24779);
and U24833 (N_24833,N_24694,N_24766);
xor U24834 (N_24834,N_24651,N_24755);
xnor U24835 (N_24835,N_24635,N_24782);
or U24836 (N_24836,N_24785,N_24767);
nand U24837 (N_24837,N_24768,N_24673);
and U24838 (N_24838,N_24719,N_24691);
or U24839 (N_24839,N_24760,N_24646);
xor U24840 (N_24840,N_24796,N_24647);
and U24841 (N_24841,N_24629,N_24618);
nor U24842 (N_24842,N_24736,N_24633);
or U24843 (N_24843,N_24676,N_24754);
xor U24844 (N_24844,N_24743,N_24792);
nor U24845 (N_24845,N_24634,N_24713);
and U24846 (N_24846,N_24644,N_24617);
xnor U24847 (N_24847,N_24687,N_24756);
nor U24848 (N_24848,N_24697,N_24737);
nand U24849 (N_24849,N_24690,N_24624);
nand U24850 (N_24850,N_24799,N_24744);
or U24851 (N_24851,N_24678,N_24763);
and U24852 (N_24852,N_24677,N_24771);
or U24853 (N_24853,N_24786,N_24735);
or U24854 (N_24854,N_24789,N_24787);
nor U24855 (N_24855,N_24775,N_24712);
or U24856 (N_24856,N_24661,N_24608);
or U24857 (N_24857,N_24772,N_24640);
nand U24858 (N_24858,N_24718,N_24688);
xnor U24859 (N_24859,N_24705,N_24700);
or U24860 (N_24860,N_24614,N_24759);
nand U24861 (N_24861,N_24626,N_24645);
nor U24862 (N_24862,N_24681,N_24774);
nand U24863 (N_24863,N_24686,N_24753);
or U24864 (N_24864,N_24730,N_24650);
and U24865 (N_24865,N_24750,N_24701);
and U24866 (N_24866,N_24656,N_24722);
or U24867 (N_24867,N_24732,N_24752);
xnor U24868 (N_24868,N_24621,N_24726);
nand U24869 (N_24869,N_24797,N_24607);
and U24870 (N_24870,N_24642,N_24623);
nand U24871 (N_24871,N_24668,N_24706);
nor U24872 (N_24872,N_24684,N_24602);
nand U24873 (N_24873,N_24600,N_24604);
xor U24874 (N_24874,N_24780,N_24670);
nand U24875 (N_24875,N_24612,N_24761);
nand U24876 (N_24876,N_24746,N_24773);
and U24877 (N_24877,N_24616,N_24672);
and U24878 (N_24878,N_24769,N_24653);
nand U24879 (N_24879,N_24643,N_24620);
nor U24880 (N_24880,N_24714,N_24641);
nor U24881 (N_24881,N_24679,N_24664);
and U24882 (N_24882,N_24675,N_24703);
xnor U24883 (N_24883,N_24648,N_24708);
nand U24884 (N_24884,N_24778,N_24682);
nor U24885 (N_24885,N_24685,N_24669);
and U24886 (N_24886,N_24658,N_24793);
nand U24887 (N_24887,N_24654,N_24622);
or U24888 (N_24888,N_24666,N_24748);
or U24889 (N_24889,N_24652,N_24671);
nor U24890 (N_24890,N_24715,N_24657);
or U24891 (N_24891,N_24683,N_24741);
xnor U24892 (N_24892,N_24781,N_24798);
and U24893 (N_24893,N_24636,N_24788);
xor U24894 (N_24894,N_24603,N_24725);
nand U24895 (N_24895,N_24609,N_24794);
or U24896 (N_24896,N_24729,N_24709);
and U24897 (N_24897,N_24720,N_24689);
and U24898 (N_24898,N_24777,N_24724);
xnor U24899 (N_24899,N_24762,N_24637);
nand U24900 (N_24900,N_24713,N_24729);
nor U24901 (N_24901,N_24723,N_24779);
xnor U24902 (N_24902,N_24707,N_24789);
nor U24903 (N_24903,N_24698,N_24783);
nand U24904 (N_24904,N_24611,N_24609);
nor U24905 (N_24905,N_24778,N_24732);
nand U24906 (N_24906,N_24646,N_24698);
nor U24907 (N_24907,N_24765,N_24778);
or U24908 (N_24908,N_24621,N_24661);
and U24909 (N_24909,N_24708,N_24717);
xor U24910 (N_24910,N_24603,N_24790);
and U24911 (N_24911,N_24721,N_24769);
and U24912 (N_24912,N_24665,N_24792);
and U24913 (N_24913,N_24779,N_24690);
nor U24914 (N_24914,N_24697,N_24685);
nand U24915 (N_24915,N_24703,N_24710);
nor U24916 (N_24916,N_24703,N_24719);
nand U24917 (N_24917,N_24712,N_24631);
xnor U24918 (N_24918,N_24792,N_24645);
nand U24919 (N_24919,N_24628,N_24748);
and U24920 (N_24920,N_24716,N_24623);
and U24921 (N_24921,N_24726,N_24742);
or U24922 (N_24922,N_24729,N_24624);
nor U24923 (N_24923,N_24673,N_24708);
nor U24924 (N_24924,N_24619,N_24601);
or U24925 (N_24925,N_24655,N_24715);
nor U24926 (N_24926,N_24798,N_24674);
and U24927 (N_24927,N_24683,N_24625);
and U24928 (N_24928,N_24682,N_24799);
nand U24929 (N_24929,N_24761,N_24633);
and U24930 (N_24930,N_24752,N_24647);
and U24931 (N_24931,N_24676,N_24713);
and U24932 (N_24932,N_24685,N_24767);
or U24933 (N_24933,N_24606,N_24653);
and U24934 (N_24934,N_24751,N_24732);
xor U24935 (N_24935,N_24692,N_24625);
and U24936 (N_24936,N_24719,N_24795);
or U24937 (N_24937,N_24737,N_24735);
and U24938 (N_24938,N_24676,N_24690);
nor U24939 (N_24939,N_24662,N_24605);
and U24940 (N_24940,N_24603,N_24671);
xor U24941 (N_24941,N_24629,N_24648);
or U24942 (N_24942,N_24616,N_24718);
or U24943 (N_24943,N_24619,N_24676);
and U24944 (N_24944,N_24688,N_24636);
nor U24945 (N_24945,N_24705,N_24601);
nand U24946 (N_24946,N_24758,N_24726);
or U24947 (N_24947,N_24656,N_24728);
or U24948 (N_24948,N_24746,N_24796);
nor U24949 (N_24949,N_24624,N_24611);
nand U24950 (N_24950,N_24726,N_24657);
or U24951 (N_24951,N_24629,N_24758);
and U24952 (N_24952,N_24673,N_24731);
nand U24953 (N_24953,N_24695,N_24700);
nor U24954 (N_24954,N_24609,N_24683);
or U24955 (N_24955,N_24788,N_24725);
nand U24956 (N_24956,N_24625,N_24680);
nor U24957 (N_24957,N_24797,N_24682);
nor U24958 (N_24958,N_24637,N_24707);
nand U24959 (N_24959,N_24636,N_24614);
nor U24960 (N_24960,N_24715,N_24761);
and U24961 (N_24961,N_24711,N_24688);
nor U24962 (N_24962,N_24679,N_24669);
and U24963 (N_24963,N_24636,N_24673);
xnor U24964 (N_24964,N_24623,N_24767);
nor U24965 (N_24965,N_24622,N_24720);
nand U24966 (N_24966,N_24773,N_24627);
and U24967 (N_24967,N_24700,N_24600);
nor U24968 (N_24968,N_24730,N_24638);
nor U24969 (N_24969,N_24621,N_24790);
xnor U24970 (N_24970,N_24747,N_24746);
nor U24971 (N_24971,N_24649,N_24664);
nand U24972 (N_24972,N_24765,N_24672);
xor U24973 (N_24973,N_24620,N_24627);
or U24974 (N_24974,N_24642,N_24688);
xor U24975 (N_24975,N_24662,N_24632);
xnor U24976 (N_24976,N_24757,N_24641);
xor U24977 (N_24977,N_24638,N_24788);
nor U24978 (N_24978,N_24751,N_24643);
xor U24979 (N_24979,N_24765,N_24642);
nand U24980 (N_24980,N_24664,N_24745);
nand U24981 (N_24981,N_24682,N_24745);
nor U24982 (N_24982,N_24634,N_24740);
nand U24983 (N_24983,N_24700,N_24665);
nand U24984 (N_24984,N_24729,N_24677);
or U24985 (N_24985,N_24707,N_24791);
or U24986 (N_24986,N_24695,N_24691);
nand U24987 (N_24987,N_24798,N_24616);
xor U24988 (N_24988,N_24697,N_24784);
nor U24989 (N_24989,N_24630,N_24725);
or U24990 (N_24990,N_24770,N_24662);
or U24991 (N_24991,N_24681,N_24673);
xor U24992 (N_24992,N_24727,N_24793);
or U24993 (N_24993,N_24702,N_24799);
or U24994 (N_24994,N_24760,N_24703);
nand U24995 (N_24995,N_24760,N_24601);
and U24996 (N_24996,N_24668,N_24666);
or U24997 (N_24997,N_24770,N_24604);
xor U24998 (N_24998,N_24605,N_24795);
xor U24999 (N_24999,N_24663,N_24750);
or U25000 (N_25000,N_24840,N_24829);
xor U25001 (N_25001,N_24864,N_24944);
xnor U25002 (N_25002,N_24990,N_24828);
or U25003 (N_25003,N_24839,N_24848);
nand U25004 (N_25004,N_24887,N_24877);
xnor U25005 (N_25005,N_24918,N_24902);
xnor U25006 (N_25006,N_24997,N_24846);
and U25007 (N_25007,N_24952,N_24979);
or U25008 (N_25008,N_24815,N_24960);
nand U25009 (N_25009,N_24933,N_24950);
xnor U25010 (N_25010,N_24989,N_24913);
or U25011 (N_25011,N_24921,N_24969);
nand U25012 (N_25012,N_24900,N_24888);
xor U25013 (N_25013,N_24996,N_24879);
xor U25014 (N_25014,N_24936,N_24855);
nor U25015 (N_25015,N_24930,N_24819);
nor U25016 (N_25016,N_24852,N_24940);
and U25017 (N_25017,N_24812,N_24860);
and U25018 (N_25018,N_24912,N_24983);
nand U25019 (N_25019,N_24807,N_24869);
xnor U25020 (N_25020,N_24982,N_24897);
nor U25021 (N_25021,N_24995,N_24975);
or U25022 (N_25022,N_24875,N_24810);
nand U25023 (N_25023,N_24842,N_24825);
nor U25024 (N_25024,N_24927,N_24946);
nor U25025 (N_25025,N_24893,N_24925);
xnor U25026 (N_25026,N_24890,N_24826);
xor U25027 (N_25027,N_24891,N_24976);
nand U25028 (N_25028,N_24813,N_24870);
or U25029 (N_25029,N_24863,N_24803);
nor U25030 (N_25030,N_24926,N_24853);
nand U25031 (N_25031,N_24945,N_24800);
nor U25032 (N_25032,N_24949,N_24993);
and U25033 (N_25033,N_24816,N_24967);
or U25034 (N_25034,N_24830,N_24943);
nor U25035 (N_25035,N_24962,N_24981);
xor U25036 (N_25036,N_24885,N_24898);
nor U25037 (N_25037,N_24977,N_24904);
nor U25038 (N_25038,N_24822,N_24858);
or U25039 (N_25039,N_24931,N_24868);
xnor U25040 (N_25040,N_24831,N_24821);
or U25041 (N_25041,N_24961,N_24915);
xnor U25042 (N_25042,N_24905,N_24827);
or U25043 (N_25043,N_24953,N_24974);
xnor U25044 (N_25044,N_24849,N_24854);
nand U25045 (N_25045,N_24935,N_24968);
and U25046 (N_25046,N_24836,N_24861);
or U25047 (N_25047,N_24917,N_24951);
nor U25048 (N_25048,N_24880,N_24886);
nor U25049 (N_25049,N_24934,N_24954);
xnor U25050 (N_25050,N_24994,N_24987);
xor U25051 (N_25051,N_24942,N_24916);
nor U25052 (N_25052,N_24899,N_24851);
nand U25053 (N_25053,N_24957,N_24823);
or U25054 (N_25054,N_24817,N_24865);
nor U25055 (N_25055,N_24901,N_24924);
xor U25056 (N_25056,N_24895,N_24970);
or U25057 (N_25057,N_24866,N_24963);
nand U25058 (N_25058,N_24920,N_24802);
nand U25059 (N_25059,N_24806,N_24850);
and U25060 (N_25060,N_24964,N_24867);
xnor U25061 (N_25061,N_24862,N_24878);
nand U25062 (N_25062,N_24938,N_24811);
xnor U25063 (N_25063,N_24948,N_24818);
nand U25064 (N_25064,N_24844,N_24988);
and U25065 (N_25065,N_24841,N_24937);
and U25066 (N_25066,N_24965,N_24859);
xor U25067 (N_25067,N_24978,N_24835);
xnor U25068 (N_25068,N_24876,N_24972);
or U25069 (N_25069,N_24958,N_24919);
and U25070 (N_25070,N_24922,N_24955);
xnor U25071 (N_25071,N_24966,N_24909);
xnor U25072 (N_25072,N_24973,N_24971);
xnor U25073 (N_25073,N_24906,N_24998);
xor U25074 (N_25074,N_24892,N_24833);
nand U25075 (N_25075,N_24820,N_24874);
nor U25076 (N_25076,N_24837,N_24838);
nor U25077 (N_25077,N_24911,N_24959);
and U25078 (N_25078,N_24847,N_24986);
or U25079 (N_25079,N_24804,N_24856);
nor U25080 (N_25080,N_24805,N_24801);
nor U25081 (N_25081,N_24984,N_24882);
xor U25082 (N_25082,N_24929,N_24991);
or U25083 (N_25083,N_24883,N_24889);
nor U25084 (N_25084,N_24914,N_24923);
nor U25085 (N_25085,N_24871,N_24908);
or U25086 (N_25086,N_24932,N_24834);
nand U25087 (N_25087,N_24896,N_24881);
xor U25088 (N_25088,N_24857,N_24939);
nand U25089 (N_25089,N_24980,N_24985);
nor U25090 (N_25090,N_24873,N_24809);
or U25091 (N_25091,N_24956,N_24992);
nor U25092 (N_25092,N_24928,N_24824);
xor U25093 (N_25093,N_24903,N_24843);
nand U25094 (N_25094,N_24910,N_24872);
and U25095 (N_25095,N_24884,N_24907);
or U25096 (N_25096,N_24832,N_24947);
and U25097 (N_25097,N_24894,N_24941);
or U25098 (N_25098,N_24845,N_24814);
and U25099 (N_25099,N_24808,N_24999);
and U25100 (N_25100,N_24879,N_24811);
xnor U25101 (N_25101,N_24902,N_24807);
xor U25102 (N_25102,N_24977,N_24972);
and U25103 (N_25103,N_24954,N_24992);
nor U25104 (N_25104,N_24817,N_24989);
nor U25105 (N_25105,N_24864,N_24891);
or U25106 (N_25106,N_24892,N_24909);
nor U25107 (N_25107,N_24967,N_24915);
nor U25108 (N_25108,N_24876,N_24982);
or U25109 (N_25109,N_24813,N_24909);
or U25110 (N_25110,N_24921,N_24935);
xnor U25111 (N_25111,N_24922,N_24821);
nand U25112 (N_25112,N_24912,N_24840);
nor U25113 (N_25113,N_24951,N_24878);
xor U25114 (N_25114,N_24947,N_24886);
nor U25115 (N_25115,N_24985,N_24992);
and U25116 (N_25116,N_24868,N_24811);
nor U25117 (N_25117,N_24921,N_24840);
or U25118 (N_25118,N_24839,N_24819);
xnor U25119 (N_25119,N_24895,N_24990);
xor U25120 (N_25120,N_24967,N_24832);
nor U25121 (N_25121,N_24928,N_24804);
nor U25122 (N_25122,N_24858,N_24853);
nor U25123 (N_25123,N_24838,N_24817);
and U25124 (N_25124,N_24828,N_24988);
and U25125 (N_25125,N_24845,N_24909);
xor U25126 (N_25126,N_24921,N_24952);
xor U25127 (N_25127,N_24821,N_24998);
and U25128 (N_25128,N_24988,N_24924);
xor U25129 (N_25129,N_24920,N_24854);
or U25130 (N_25130,N_24979,N_24862);
nor U25131 (N_25131,N_24926,N_24823);
nand U25132 (N_25132,N_24869,N_24992);
nand U25133 (N_25133,N_24905,N_24997);
and U25134 (N_25134,N_24963,N_24875);
and U25135 (N_25135,N_24846,N_24813);
nor U25136 (N_25136,N_24842,N_24898);
and U25137 (N_25137,N_24865,N_24945);
or U25138 (N_25138,N_24886,N_24894);
nand U25139 (N_25139,N_24911,N_24939);
nand U25140 (N_25140,N_24922,N_24836);
or U25141 (N_25141,N_24875,N_24862);
xnor U25142 (N_25142,N_24968,N_24858);
xor U25143 (N_25143,N_24953,N_24843);
nand U25144 (N_25144,N_24979,N_24847);
nand U25145 (N_25145,N_24955,N_24919);
xor U25146 (N_25146,N_24996,N_24944);
nor U25147 (N_25147,N_24882,N_24958);
and U25148 (N_25148,N_24881,N_24859);
or U25149 (N_25149,N_24959,N_24944);
xor U25150 (N_25150,N_24952,N_24867);
xor U25151 (N_25151,N_24948,N_24846);
xor U25152 (N_25152,N_24964,N_24989);
or U25153 (N_25153,N_24844,N_24994);
and U25154 (N_25154,N_24877,N_24886);
and U25155 (N_25155,N_24841,N_24885);
nor U25156 (N_25156,N_24805,N_24832);
nor U25157 (N_25157,N_24823,N_24933);
nor U25158 (N_25158,N_24994,N_24898);
nand U25159 (N_25159,N_24822,N_24936);
or U25160 (N_25160,N_24858,N_24865);
xnor U25161 (N_25161,N_24884,N_24909);
or U25162 (N_25162,N_24883,N_24859);
xor U25163 (N_25163,N_24871,N_24806);
or U25164 (N_25164,N_24847,N_24890);
and U25165 (N_25165,N_24895,N_24803);
and U25166 (N_25166,N_24872,N_24991);
and U25167 (N_25167,N_24874,N_24943);
and U25168 (N_25168,N_24987,N_24880);
and U25169 (N_25169,N_24855,N_24835);
xnor U25170 (N_25170,N_24929,N_24910);
nand U25171 (N_25171,N_24880,N_24919);
nand U25172 (N_25172,N_24916,N_24962);
xor U25173 (N_25173,N_24908,N_24930);
xor U25174 (N_25174,N_24993,N_24965);
xor U25175 (N_25175,N_24947,N_24875);
nand U25176 (N_25176,N_24892,N_24938);
and U25177 (N_25177,N_24966,N_24860);
nand U25178 (N_25178,N_24943,N_24843);
nand U25179 (N_25179,N_24960,N_24972);
nand U25180 (N_25180,N_24972,N_24859);
and U25181 (N_25181,N_24847,N_24843);
nand U25182 (N_25182,N_24912,N_24929);
or U25183 (N_25183,N_24870,N_24950);
nor U25184 (N_25184,N_24892,N_24830);
nand U25185 (N_25185,N_24941,N_24872);
xnor U25186 (N_25186,N_24867,N_24970);
xor U25187 (N_25187,N_24904,N_24850);
nor U25188 (N_25188,N_24900,N_24905);
nand U25189 (N_25189,N_24959,N_24962);
or U25190 (N_25190,N_24899,N_24872);
or U25191 (N_25191,N_24977,N_24880);
and U25192 (N_25192,N_24911,N_24892);
and U25193 (N_25193,N_24905,N_24959);
xor U25194 (N_25194,N_24983,N_24952);
nor U25195 (N_25195,N_24889,N_24909);
and U25196 (N_25196,N_24955,N_24855);
and U25197 (N_25197,N_24835,N_24963);
xnor U25198 (N_25198,N_24927,N_24884);
and U25199 (N_25199,N_24992,N_24923);
or U25200 (N_25200,N_25013,N_25040);
nand U25201 (N_25201,N_25156,N_25159);
or U25202 (N_25202,N_25165,N_25055);
nand U25203 (N_25203,N_25034,N_25078);
nand U25204 (N_25204,N_25080,N_25098);
and U25205 (N_25205,N_25031,N_25076);
or U25206 (N_25206,N_25152,N_25151);
xor U25207 (N_25207,N_25119,N_25154);
xor U25208 (N_25208,N_25103,N_25097);
or U25209 (N_25209,N_25054,N_25092);
nand U25210 (N_25210,N_25135,N_25089);
xnor U25211 (N_25211,N_25161,N_25198);
and U25212 (N_25212,N_25063,N_25058);
and U25213 (N_25213,N_25132,N_25006);
or U25214 (N_25214,N_25102,N_25193);
nor U25215 (N_25215,N_25045,N_25150);
and U25216 (N_25216,N_25148,N_25053);
nand U25217 (N_25217,N_25002,N_25004);
xor U25218 (N_25218,N_25181,N_25039);
or U25219 (N_25219,N_25069,N_25167);
or U25220 (N_25220,N_25026,N_25180);
xnor U25221 (N_25221,N_25021,N_25084);
xnor U25222 (N_25222,N_25065,N_25127);
xor U25223 (N_25223,N_25008,N_25196);
nor U25224 (N_25224,N_25114,N_25178);
or U25225 (N_25225,N_25182,N_25083);
or U25226 (N_25226,N_25033,N_25011);
xnor U25227 (N_25227,N_25066,N_25142);
or U25228 (N_25228,N_25136,N_25175);
nand U25229 (N_25229,N_25126,N_25168);
nor U25230 (N_25230,N_25101,N_25029);
xnor U25231 (N_25231,N_25115,N_25163);
nor U25232 (N_25232,N_25057,N_25007);
nor U25233 (N_25233,N_25070,N_25185);
nand U25234 (N_25234,N_25138,N_25189);
or U25235 (N_25235,N_25199,N_25091);
xor U25236 (N_25236,N_25164,N_25116);
nor U25237 (N_25237,N_25095,N_25162);
nand U25238 (N_25238,N_25197,N_25099);
xor U25239 (N_25239,N_25052,N_25170);
and U25240 (N_25240,N_25022,N_25106);
or U25241 (N_25241,N_25049,N_25068);
nand U25242 (N_25242,N_25048,N_25158);
nor U25243 (N_25243,N_25130,N_25113);
nor U25244 (N_25244,N_25143,N_25096);
nor U25245 (N_25245,N_25001,N_25051);
or U25246 (N_25246,N_25061,N_25191);
nor U25247 (N_25247,N_25017,N_25038);
nor U25248 (N_25248,N_25169,N_25081);
nand U25249 (N_25249,N_25184,N_25157);
or U25250 (N_25250,N_25186,N_25059);
or U25251 (N_25251,N_25036,N_25192);
or U25252 (N_25252,N_25064,N_25079);
xor U25253 (N_25253,N_25062,N_25173);
nor U25254 (N_25254,N_25023,N_25117);
and U25255 (N_25255,N_25035,N_25146);
and U25256 (N_25256,N_25019,N_25129);
and U25257 (N_25257,N_25074,N_25088);
and U25258 (N_25258,N_25124,N_25003);
and U25259 (N_25259,N_25190,N_25118);
and U25260 (N_25260,N_25100,N_25028);
and U25261 (N_25261,N_25010,N_25147);
xor U25262 (N_25262,N_25122,N_25043);
xnor U25263 (N_25263,N_25134,N_25009);
nor U25264 (N_25264,N_25015,N_25149);
nor U25265 (N_25265,N_25176,N_25172);
nand U25266 (N_25266,N_25187,N_25195);
nand U25267 (N_25267,N_25133,N_25166);
nor U25268 (N_25268,N_25108,N_25090);
xor U25269 (N_25269,N_25016,N_25093);
or U25270 (N_25270,N_25042,N_25144);
xnor U25271 (N_25271,N_25044,N_25123);
and U25272 (N_25272,N_25112,N_25073);
nor U25273 (N_25273,N_25183,N_25107);
nand U25274 (N_25274,N_25131,N_25041);
nor U25275 (N_25275,N_25120,N_25014);
nand U25276 (N_25276,N_25139,N_25109);
and U25277 (N_25277,N_25037,N_25025);
xnor U25278 (N_25278,N_25179,N_25171);
and U25279 (N_25279,N_25160,N_25105);
and U25280 (N_25280,N_25032,N_25086);
and U25281 (N_25281,N_25141,N_25174);
and U25282 (N_25282,N_25027,N_25024);
or U25283 (N_25283,N_25005,N_25020);
and U25284 (N_25284,N_25018,N_25121);
nand U25285 (N_25285,N_25056,N_25137);
nor U25286 (N_25286,N_25075,N_25050);
and U25287 (N_25287,N_25145,N_25094);
nand U25288 (N_25288,N_25111,N_25110);
and U25289 (N_25289,N_25067,N_25046);
nor U25290 (N_25290,N_25012,N_25087);
or U25291 (N_25291,N_25030,N_25153);
and U25292 (N_25292,N_25071,N_25155);
and U25293 (N_25293,N_25104,N_25072);
nand U25294 (N_25294,N_25128,N_25188);
xnor U25295 (N_25295,N_25085,N_25140);
and U25296 (N_25296,N_25077,N_25000);
nand U25297 (N_25297,N_25047,N_25082);
nor U25298 (N_25298,N_25060,N_25177);
nand U25299 (N_25299,N_25194,N_25125);
xnor U25300 (N_25300,N_25174,N_25143);
nor U25301 (N_25301,N_25064,N_25035);
nor U25302 (N_25302,N_25060,N_25134);
xor U25303 (N_25303,N_25012,N_25072);
and U25304 (N_25304,N_25036,N_25046);
nand U25305 (N_25305,N_25163,N_25086);
nand U25306 (N_25306,N_25157,N_25086);
and U25307 (N_25307,N_25133,N_25084);
and U25308 (N_25308,N_25151,N_25141);
xor U25309 (N_25309,N_25139,N_25190);
or U25310 (N_25310,N_25138,N_25079);
nor U25311 (N_25311,N_25046,N_25141);
and U25312 (N_25312,N_25063,N_25126);
xor U25313 (N_25313,N_25036,N_25132);
or U25314 (N_25314,N_25011,N_25159);
or U25315 (N_25315,N_25196,N_25187);
nor U25316 (N_25316,N_25191,N_25086);
xor U25317 (N_25317,N_25122,N_25179);
xor U25318 (N_25318,N_25183,N_25007);
and U25319 (N_25319,N_25078,N_25142);
nand U25320 (N_25320,N_25089,N_25070);
nand U25321 (N_25321,N_25170,N_25087);
xor U25322 (N_25322,N_25120,N_25060);
nand U25323 (N_25323,N_25026,N_25033);
xor U25324 (N_25324,N_25112,N_25061);
nor U25325 (N_25325,N_25093,N_25152);
nor U25326 (N_25326,N_25151,N_25071);
nand U25327 (N_25327,N_25181,N_25056);
xor U25328 (N_25328,N_25151,N_25045);
xor U25329 (N_25329,N_25159,N_25010);
or U25330 (N_25330,N_25000,N_25108);
nand U25331 (N_25331,N_25021,N_25183);
nor U25332 (N_25332,N_25101,N_25120);
xnor U25333 (N_25333,N_25050,N_25100);
or U25334 (N_25334,N_25191,N_25063);
or U25335 (N_25335,N_25078,N_25028);
xor U25336 (N_25336,N_25157,N_25075);
nor U25337 (N_25337,N_25062,N_25088);
nor U25338 (N_25338,N_25124,N_25012);
nor U25339 (N_25339,N_25113,N_25158);
nand U25340 (N_25340,N_25029,N_25112);
or U25341 (N_25341,N_25150,N_25098);
xnor U25342 (N_25342,N_25091,N_25038);
xnor U25343 (N_25343,N_25116,N_25047);
or U25344 (N_25344,N_25197,N_25033);
and U25345 (N_25345,N_25009,N_25141);
xnor U25346 (N_25346,N_25070,N_25171);
or U25347 (N_25347,N_25196,N_25034);
and U25348 (N_25348,N_25184,N_25172);
or U25349 (N_25349,N_25187,N_25030);
nand U25350 (N_25350,N_25144,N_25170);
and U25351 (N_25351,N_25073,N_25102);
or U25352 (N_25352,N_25149,N_25059);
xor U25353 (N_25353,N_25047,N_25146);
and U25354 (N_25354,N_25197,N_25019);
xor U25355 (N_25355,N_25181,N_25186);
nand U25356 (N_25356,N_25013,N_25190);
nand U25357 (N_25357,N_25094,N_25110);
nand U25358 (N_25358,N_25081,N_25106);
or U25359 (N_25359,N_25112,N_25078);
xor U25360 (N_25360,N_25095,N_25064);
or U25361 (N_25361,N_25165,N_25116);
nand U25362 (N_25362,N_25030,N_25039);
or U25363 (N_25363,N_25052,N_25043);
nor U25364 (N_25364,N_25008,N_25078);
nor U25365 (N_25365,N_25068,N_25105);
and U25366 (N_25366,N_25139,N_25047);
nor U25367 (N_25367,N_25198,N_25166);
nor U25368 (N_25368,N_25113,N_25085);
xnor U25369 (N_25369,N_25059,N_25193);
nor U25370 (N_25370,N_25092,N_25112);
nand U25371 (N_25371,N_25116,N_25023);
and U25372 (N_25372,N_25013,N_25054);
and U25373 (N_25373,N_25170,N_25026);
and U25374 (N_25374,N_25055,N_25074);
nand U25375 (N_25375,N_25186,N_25167);
nor U25376 (N_25376,N_25059,N_25100);
and U25377 (N_25377,N_25091,N_25142);
nand U25378 (N_25378,N_25057,N_25098);
or U25379 (N_25379,N_25077,N_25172);
nand U25380 (N_25380,N_25011,N_25048);
nor U25381 (N_25381,N_25188,N_25189);
nand U25382 (N_25382,N_25093,N_25125);
nand U25383 (N_25383,N_25095,N_25076);
and U25384 (N_25384,N_25095,N_25158);
xnor U25385 (N_25385,N_25125,N_25016);
and U25386 (N_25386,N_25168,N_25084);
or U25387 (N_25387,N_25050,N_25003);
nand U25388 (N_25388,N_25143,N_25118);
nor U25389 (N_25389,N_25068,N_25120);
or U25390 (N_25390,N_25021,N_25016);
nor U25391 (N_25391,N_25113,N_25070);
nand U25392 (N_25392,N_25097,N_25030);
and U25393 (N_25393,N_25149,N_25066);
xor U25394 (N_25394,N_25107,N_25086);
or U25395 (N_25395,N_25073,N_25119);
or U25396 (N_25396,N_25181,N_25093);
xor U25397 (N_25397,N_25170,N_25133);
nand U25398 (N_25398,N_25107,N_25075);
nor U25399 (N_25399,N_25117,N_25074);
nor U25400 (N_25400,N_25242,N_25214);
or U25401 (N_25401,N_25294,N_25260);
xnor U25402 (N_25402,N_25272,N_25210);
xor U25403 (N_25403,N_25282,N_25361);
and U25404 (N_25404,N_25309,N_25231);
and U25405 (N_25405,N_25261,N_25224);
nand U25406 (N_25406,N_25228,N_25236);
nor U25407 (N_25407,N_25322,N_25232);
nand U25408 (N_25408,N_25312,N_25235);
or U25409 (N_25409,N_25338,N_25342);
or U25410 (N_25410,N_25364,N_25286);
and U25411 (N_25411,N_25324,N_25373);
or U25412 (N_25412,N_25331,N_25360);
and U25413 (N_25413,N_25233,N_25229);
and U25414 (N_25414,N_25247,N_25302);
and U25415 (N_25415,N_25392,N_25305);
or U25416 (N_25416,N_25366,N_25274);
xnor U25417 (N_25417,N_25262,N_25217);
xor U25418 (N_25418,N_25288,N_25240);
nand U25419 (N_25419,N_25268,N_25368);
nand U25420 (N_25420,N_25343,N_25215);
or U25421 (N_25421,N_25378,N_25308);
nand U25422 (N_25422,N_25399,N_25390);
xor U25423 (N_25423,N_25382,N_25213);
nand U25424 (N_25424,N_25299,N_25375);
or U25425 (N_25425,N_25307,N_25269);
xnor U25426 (N_25426,N_25241,N_25347);
nand U25427 (N_25427,N_25396,N_25328);
nand U25428 (N_25428,N_25298,N_25283);
nand U25429 (N_25429,N_25310,N_25320);
nor U25430 (N_25430,N_25264,N_25349);
or U25431 (N_25431,N_25205,N_25234);
nor U25432 (N_25432,N_25358,N_25394);
xor U25433 (N_25433,N_25265,N_25275);
nor U25434 (N_25434,N_25387,N_25389);
and U25435 (N_25435,N_25249,N_25250);
nand U25436 (N_25436,N_25251,N_25271);
xor U25437 (N_25437,N_25263,N_25201);
xnor U25438 (N_25438,N_25222,N_25397);
xor U25439 (N_25439,N_25369,N_25248);
and U25440 (N_25440,N_25336,N_25371);
or U25441 (N_25441,N_25257,N_25395);
nand U25442 (N_25442,N_25359,N_25239);
nor U25443 (N_25443,N_25221,N_25351);
and U25444 (N_25444,N_25206,N_25208);
xnor U25445 (N_25445,N_25334,N_25219);
or U25446 (N_25446,N_25367,N_25204);
xnor U25447 (N_25447,N_25245,N_25393);
and U25448 (N_25448,N_25381,N_25339);
and U25449 (N_25449,N_25212,N_25332);
nand U25450 (N_25450,N_25279,N_25256);
xor U25451 (N_25451,N_25267,N_25345);
or U25452 (N_25452,N_25374,N_25379);
or U25453 (N_25453,N_25281,N_25385);
nor U25454 (N_25454,N_25344,N_25346);
or U25455 (N_25455,N_25252,N_25291);
and U25456 (N_25456,N_25292,N_25277);
xor U25457 (N_25457,N_25316,N_25227);
and U25458 (N_25458,N_25362,N_25230);
or U25459 (N_25459,N_25335,N_25211);
xor U25460 (N_25460,N_25200,N_25293);
nand U25461 (N_25461,N_25377,N_25243);
nor U25462 (N_25462,N_25350,N_25357);
xnor U25463 (N_25463,N_25318,N_25383);
nor U25464 (N_25464,N_25329,N_25319);
xor U25465 (N_25465,N_25391,N_25254);
nand U25466 (N_25466,N_25244,N_25326);
nor U25467 (N_25467,N_25203,N_25304);
nand U25468 (N_25468,N_25273,N_25380);
nor U25469 (N_25469,N_25363,N_25295);
nor U25470 (N_25470,N_25384,N_25388);
or U25471 (N_25471,N_25209,N_25258);
and U25472 (N_25472,N_25365,N_25287);
nand U25473 (N_25473,N_25253,N_25303);
and U25474 (N_25474,N_25372,N_25340);
nor U25475 (N_25475,N_25354,N_25284);
or U25476 (N_25476,N_25280,N_25255);
or U25477 (N_25477,N_25333,N_25348);
nor U25478 (N_25478,N_25306,N_25289);
xnor U25479 (N_25479,N_25218,N_25237);
or U25480 (N_25480,N_25317,N_25301);
and U25481 (N_25481,N_25321,N_25311);
or U25482 (N_25482,N_25313,N_25296);
or U25483 (N_25483,N_25266,N_25297);
or U25484 (N_25484,N_25276,N_25259);
and U25485 (N_25485,N_25290,N_25207);
nand U25486 (N_25486,N_25356,N_25226);
xnor U25487 (N_25487,N_25325,N_25353);
nor U25488 (N_25488,N_25285,N_25352);
or U25489 (N_25489,N_25323,N_25270);
and U25490 (N_25490,N_25202,N_25278);
and U25491 (N_25491,N_25386,N_25398);
nor U25492 (N_25492,N_25300,N_25238);
nor U25493 (N_25493,N_25216,N_25220);
or U25494 (N_25494,N_25330,N_25223);
or U25495 (N_25495,N_25225,N_25341);
and U25496 (N_25496,N_25314,N_25246);
nor U25497 (N_25497,N_25337,N_25370);
and U25498 (N_25498,N_25327,N_25355);
nand U25499 (N_25499,N_25315,N_25376);
nand U25500 (N_25500,N_25330,N_25265);
and U25501 (N_25501,N_25346,N_25294);
or U25502 (N_25502,N_25228,N_25237);
nand U25503 (N_25503,N_25332,N_25386);
xor U25504 (N_25504,N_25299,N_25352);
nor U25505 (N_25505,N_25299,N_25332);
and U25506 (N_25506,N_25383,N_25204);
nor U25507 (N_25507,N_25394,N_25238);
and U25508 (N_25508,N_25292,N_25301);
nor U25509 (N_25509,N_25374,N_25251);
xor U25510 (N_25510,N_25205,N_25340);
xor U25511 (N_25511,N_25280,N_25297);
nor U25512 (N_25512,N_25391,N_25252);
xor U25513 (N_25513,N_25288,N_25238);
or U25514 (N_25514,N_25233,N_25363);
or U25515 (N_25515,N_25326,N_25375);
xor U25516 (N_25516,N_25320,N_25309);
nand U25517 (N_25517,N_25274,N_25252);
nor U25518 (N_25518,N_25354,N_25272);
nor U25519 (N_25519,N_25229,N_25200);
and U25520 (N_25520,N_25356,N_25296);
or U25521 (N_25521,N_25213,N_25233);
xnor U25522 (N_25522,N_25365,N_25394);
and U25523 (N_25523,N_25244,N_25287);
nand U25524 (N_25524,N_25251,N_25299);
or U25525 (N_25525,N_25295,N_25314);
nand U25526 (N_25526,N_25361,N_25264);
and U25527 (N_25527,N_25321,N_25367);
nor U25528 (N_25528,N_25239,N_25376);
nor U25529 (N_25529,N_25238,N_25379);
nor U25530 (N_25530,N_25315,N_25218);
nor U25531 (N_25531,N_25224,N_25392);
or U25532 (N_25532,N_25263,N_25364);
or U25533 (N_25533,N_25210,N_25221);
xnor U25534 (N_25534,N_25215,N_25373);
nor U25535 (N_25535,N_25285,N_25337);
nand U25536 (N_25536,N_25319,N_25376);
and U25537 (N_25537,N_25306,N_25200);
nor U25538 (N_25538,N_25393,N_25389);
and U25539 (N_25539,N_25371,N_25319);
xor U25540 (N_25540,N_25204,N_25301);
nand U25541 (N_25541,N_25356,N_25228);
xor U25542 (N_25542,N_25260,N_25228);
nor U25543 (N_25543,N_25269,N_25260);
or U25544 (N_25544,N_25228,N_25352);
nand U25545 (N_25545,N_25230,N_25288);
nand U25546 (N_25546,N_25350,N_25245);
and U25547 (N_25547,N_25234,N_25281);
nor U25548 (N_25548,N_25217,N_25378);
nor U25549 (N_25549,N_25398,N_25224);
xor U25550 (N_25550,N_25284,N_25201);
or U25551 (N_25551,N_25368,N_25397);
and U25552 (N_25552,N_25279,N_25207);
nand U25553 (N_25553,N_25287,N_25394);
and U25554 (N_25554,N_25397,N_25320);
or U25555 (N_25555,N_25250,N_25227);
nand U25556 (N_25556,N_25290,N_25325);
nand U25557 (N_25557,N_25352,N_25323);
nand U25558 (N_25558,N_25243,N_25308);
nor U25559 (N_25559,N_25380,N_25322);
xnor U25560 (N_25560,N_25378,N_25381);
xor U25561 (N_25561,N_25264,N_25360);
and U25562 (N_25562,N_25318,N_25265);
or U25563 (N_25563,N_25307,N_25261);
or U25564 (N_25564,N_25205,N_25259);
nor U25565 (N_25565,N_25326,N_25383);
or U25566 (N_25566,N_25260,N_25247);
nand U25567 (N_25567,N_25357,N_25264);
or U25568 (N_25568,N_25240,N_25334);
or U25569 (N_25569,N_25219,N_25294);
nand U25570 (N_25570,N_25261,N_25380);
xnor U25571 (N_25571,N_25259,N_25202);
xnor U25572 (N_25572,N_25368,N_25301);
nand U25573 (N_25573,N_25246,N_25266);
xnor U25574 (N_25574,N_25390,N_25218);
and U25575 (N_25575,N_25252,N_25203);
nor U25576 (N_25576,N_25343,N_25259);
xnor U25577 (N_25577,N_25222,N_25255);
and U25578 (N_25578,N_25238,N_25210);
and U25579 (N_25579,N_25385,N_25391);
nand U25580 (N_25580,N_25266,N_25235);
nand U25581 (N_25581,N_25358,N_25365);
nand U25582 (N_25582,N_25395,N_25292);
or U25583 (N_25583,N_25220,N_25207);
nor U25584 (N_25584,N_25214,N_25277);
or U25585 (N_25585,N_25217,N_25328);
or U25586 (N_25586,N_25363,N_25294);
and U25587 (N_25587,N_25286,N_25381);
xnor U25588 (N_25588,N_25372,N_25211);
nand U25589 (N_25589,N_25335,N_25295);
xnor U25590 (N_25590,N_25300,N_25367);
nor U25591 (N_25591,N_25348,N_25317);
xnor U25592 (N_25592,N_25391,N_25359);
or U25593 (N_25593,N_25296,N_25202);
or U25594 (N_25594,N_25382,N_25342);
and U25595 (N_25595,N_25327,N_25350);
nand U25596 (N_25596,N_25346,N_25322);
and U25597 (N_25597,N_25370,N_25386);
or U25598 (N_25598,N_25379,N_25328);
nor U25599 (N_25599,N_25361,N_25306);
and U25600 (N_25600,N_25595,N_25557);
and U25601 (N_25601,N_25571,N_25436);
xnor U25602 (N_25602,N_25424,N_25497);
or U25603 (N_25603,N_25429,N_25585);
nand U25604 (N_25604,N_25517,N_25404);
nand U25605 (N_25605,N_25443,N_25551);
and U25606 (N_25606,N_25584,N_25423);
nand U25607 (N_25607,N_25559,N_25508);
or U25608 (N_25608,N_25572,N_25469);
nand U25609 (N_25609,N_25412,N_25545);
or U25610 (N_25610,N_25428,N_25570);
or U25611 (N_25611,N_25536,N_25460);
nand U25612 (N_25612,N_25566,N_25544);
nor U25613 (N_25613,N_25542,N_25503);
nand U25614 (N_25614,N_25589,N_25513);
and U25615 (N_25615,N_25474,N_25445);
or U25616 (N_25616,N_25512,N_25568);
xnor U25617 (N_25617,N_25507,N_25457);
and U25618 (N_25618,N_25588,N_25531);
xnor U25619 (N_25619,N_25535,N_25440);
and U25620 (N_25620,N_25498,N_25415);
or U25621 (N_25621,N_25519,N_25597);
or U25622 (N_25622,N_25516,N_25420);
nor U25623 (N_25623,N_25478,N_25502);
nand U25624 (N_25624,N_25522,N_25527);
nor U25625 (N_25625,N_25538,N_25549);
nor U25626 (N_25626,N_25598,N_25521);
and U25627 (N_25627,N_25526,N_25400);
and U25628 (N_25628,N_25465,N_25416);
or U25629 (N_25629,N_25447,N_25590);
nand U25630 (N_25630,N_25403,N_25483);
nand U25631 (N_25631,N_25533,N_25406);
or U25632 (N_25632,N_25467,N_25528);
xor U25633 (N_25633,N_25461,N_25435);
nor U25634 (N_25634,N_25427,N_25471);
nand U25635 (N_25635,N_25567,N_25520);
xor U25636 (N_25636,N_25441,N_25450);
xor U25637 (N_25637,N_25456,N_25564);
xnor U25638 (N_25638,N_25599,N_25425);
nand U25639 (N_25639,N_25446,N_25496);
nand U25640 (N_25640,N_25470,N_25401);
xnor U25641 (N_25641,N_25484,N_25488);
xor U25642 (N_25642,N_25472,N_25459);
nand U25643 (N_25643,N_25586,N_25493);
nor U25644 (N_25644,N_25454,N_25405);
nand U25645 (N_25645,N_25539,N_25569);
or U25646 (N_25646,N_25444,N_25431);
nand U25647 (N_25647,N_25560,N_25554);
xnor U25648 (N_25648,N_25552,N_25462);
and U25649 (N_25649,N_25555,N_25558);
nand U25650 (N_25650,N_25473,N_25573);
xor U25651 (N_25651,N_25505,N_25529);
nand U25652 (N_25652,N_25458,N_25562);
xnor U25653 (N_25653,N_25407,N_25408);
nand U25654 (N_25654,N_25534,N_25583);
xor U25655 (N_25655,N_25437,N_25442);
xor U25656 (N_25656,N_25546,N_25587);
xor U25657 (N_25657,N_25550,N_25448);
or U25658 (N_25658,N_25480,N_25490);
and U25659 (N_25659,N_25577,N_25481);
or U25660 (N_25660,N_25579,N_25482);
nor U25661 (N_25661,N_25422,N_25582);
nand U25662 (N_25662,N_25426,N_25409);
xor U25663 (N_25663,N_25455,N_25561);
nor U25664 (N_25664,N_25530,N_25563);
nor U25665 (N_25665,N_25466,N_25402);
or U25666 (N_25666,N_25540,N_25506);
nor U25667 (N_25667,N_25553,N_25479);
nor U25668 (N_25668,N_25477,N_25578);
xor U25669 (N_25669,N_25548,N_25432);
xor U25670 (N_25670,N_25524,N_25451);
nor U25671 (N_25671,N_25565,N_25414);
and U25672 (N_25672,N_25532,N_25452);
nor U25673 (N_25673,N_25434,N_25591);
xor U25674 (N_25674,N_25575,N_25489);
and U25675 (N_25675,N_25543,N_25523);
nand U25676 (N_25676,N_25511,N_25495);
and U25677 (N_25677,N_25492,N_25463);
nand U25678 (N_25678,N_25518,N_25494);
nor U25679 (N_25679,N_25475,N_25491);
nor U25680 (N_25680,N_25439,N_25419);
nor U25681 (N_25681,N_25514,N_25596);
xor U25682 (N_25682,N_25592,N_25417);
xor U25683 (N_25683,N_25464,N_25547);
nor U25684 (N_25684,N_25430,N_25449);
or U25685 (N_25685,N_25509,N_25500);
and U25686 (N_25686,N_25499,N_25485);
xor U25687 (N_25687,N_25433,N_25525);
and U25688 (N_25688,N_25504,N_25510);
nor U25689 (N_25689,N_25576,N_25438);
nor U25690 (N_25690,N_25580,N_25411);
and U25691 (N_25691,N_25468,N_25541);
nand U25692 (N_25692,N_25476,N_25556);
and U25693 (N_25693,N_25593,N_25487);
or U25694 (N_25694,N_25410,N_25413);
nor U25695 (N_25695,N_25486,N_25574);
nor U25696 (N_25696,N_25515,N_25501);
or U25697 (N_25697,N_25537,N_25418);
xor U25698 (N_25698,N_25581,N_25421);
xnor U25699 (N_25699,N_25594,N_25453);
xor U25700 (N_25700,N_25437,N_25569);
nor U25701 (N_25701,N_25573,N_25533);
nor U25702 (N_25702,N_25579,N_25414);
nand U25703 (N_25703,N_25435,N_25551);
nor U25704 (N_25704,N_25495,N_25440);
xnor U25705 (N_25705,N_25420,N_25458);
nor U25706 (N_25706,N_25538,N_25578);
nor U25707 (N_25707,N_25592,N_25486);
xnor U25708 (N_25708,N_25496,N_25583);
xor U25709 (N_25709,N_25551,N_25593);
xor U25710 (N_25710,N_25508,N_25546);
nand U25711 (N_25711,N_25419,N_25412);
xor U25712 (N_25712,N_25597,N_25477);
xnor U25713 (N_25713,N_25520,N_25459);
nor U25714 (N_25714,N_25428,N_25574);
xnor U25715 (N_25715,N_25516,N_25533);
xor U25716 (N_25716,N_25575,N_25551);
and U25717 (N_25717,N_25444,N_25538);
nand U25718 (N_25718,N_25527,N_25406);
nand U25719 (N_25719,N_25511,N_25480);
xnor U25720 (N_25720,N_25489,N_25501);
xor U25721 (N_25721,N_25496,N_25465);
nand U25722 (N_25722,N_25582,N_25415);
and U25723 (N_25723,N_25480,N_25508);
nor U25724 (N_25724,N_25451,N_25444);
nor U25725 (N_25725,N_25447,N_25555);
xor U25726 (N_25726,N_25523,N_25531);
xor U25727 (N_25727,N_25435,N_25477);
or U25728 (N_25728,N_25461,N_25586);
nor U25729 (N_25729,N_25570,N_25596);
or U25730 (N_25730,N_25543,N_25565);
or U25731 (N_25731,N_25485,N_25529);
and U25732 (N_25732,N_25453,N_25478);
nor U25733 (N_25733,N_25528,N_25417);
nand U25734 (N_25734,N_25433,N_25443);
nand U25735 (N_25735,N_25592,N_25574);
nand U25736 (N_25736,N_25564,N_25486);
or U25737 (N_25737,N_25565,N_25510);
or U25738 (N_25738,N_25518,N_25581);
and U25739 (N_25739,N_25591,N_25594);
xor U25740 (N_25740,N_25509,N_25526);
or U25741 (N_25741,N_25543,N_25411);
or U25742 (N_25742,N_25555,N_25533);
nor U25743 (N_25743,N_25445,N_25449);
nor U25744 (N_25744,N_25589,N_25458);
and U25745 (N_25745,N_25599,N_25426);
xnor U25746 (N_25746,N_25517,N_25424);
nand U25747 (N_25747,N_25518,N_25567);
nand U25748 (N_25748,N_25558,N_25486);
nand U25749 (N_25749,N_25556,N_25437);
or U25750 (N_25750,N_25565,N_25488);
nor U25751 (N_25751,N_25505,N_25402);
nor U25752 (N_25752,N_25475,N_25564);
nand U25753 (N_25753,N_25459,N_25449);
xnor U25754 (N_25754,N_25534,N_25541);
nor U25755 (N_25755,N_25471,N_25400);
xnor U25756 (N_25756,N_25592,N_25507);
xor U25757 (N_25757,N_25520,N_25417);
nor U25758 (N_25758,N_25494,N_25598);
xor U25759 (N_25759,N_25470,N_25489);
xnor U25760 (N_25760,N_25458,N_25587);
nor U25761 (N_25761,N_25535,N_25446);
nor U25762 (N_25762,N_25403,N_25506);
xnor U25763 (N_25763,N_25549,N_25564);
and U25764 (N_25764,N_25561,N_25438);
or U25765 (N_25765,N_25478,N_25404);
or U25766 (N_25766,N_25568,N_25508);
or U25767 (N_25767,N_25501,N_25422);
xnor U25768 (N_25768,N_25502,N_25498);
xnor U25769 (N_25769,N_25521,N_25428);
xnor U25770 (N_25770,N_25446,N_25517);
and U25771 (N_25771,N_25409,N_25422);
xnor U25772 (N_25772,N_25502,N_25525);
nand U25773 (N_25773,N_25486,N_25577);
and U25774 (N_25774,N_25413,N_25444);
nand U25775 (N_25775,N_25482,N_25432);
nand U25776 (N_25776,N_25569,N_25480);
nor U25777 (N_25777,N_25456,N_25492);
xnor U25778 (N_25778,N_25437,N_25568);
nand U25779 (N_25779,N_25478,N_25473);
nand U25780 (N_25780,N_25449,N_25447);
xor U25781 (N_25781,N_25590,N_25476);
nand U25782 (N_25782,N_25570,N_25547);
nand U25783 (N_25783,N_25568,N_25550);
nand U25784 (N_25784,N_25595,N_25509);
and U25785 (N_25785,N_25528,N_25574);
nor U25786 (N_25786,N_25595,N_25441);
xor U25787 (N_25787,N_25416,N_25573);
nand U25788 (N_25788,N_25429,N_25514);
and U25789 (N_25789,N_25402,N_25535);
and U25790 (N_25790,N_25562,N_25593);
or U25791 (N_25791,N_25430,N_25518);
and U25792 (N_25792,N_25531,N_25585);
xnor U25793 (N_25793,N_25433,N_25543);
nor U25794 (N_25794,N_25597,N_25507);
nand U25795 (N_25795,N_25520,N_25468);
and U25796 (N_25796,N_25529,N_25524);
or U25797 (N_25797,N_25485,N_25558);
nand U25798 (N_25798,N_25478,N_25586);
or U25799 (N_25799,N_25551,N_25463);
and U25800 (N_25800,N_25768,N_25710);
nand U25801 (N_25801,N_25799,N_25749);
and U25802 (N_25802,N_25697,N_25665);
nor U25803 (N_25803,N_25751,N_25681);
or U25804 (N_25804,N_25714,N_25638);
and U25805 (N_25805,N_25703,N_25625);
and U25806 (N_25806,N_25700,N_25632);
xor U25807 (N_25807,N_25758,N_25605);
and U25808 (N_25808,N_25619,N_25694);
xnor U25809 (N_25809,N_25601,N_25655);
and U25810 (N_25810,N_25740,N_25786);
or U25811 (N_25811,N_25727,N_25676);
and U25812 (N_25812,N_25760,N_25660);
nor U25813 (N_25813,N_25646,N_25645);
xnor U25814 (N_25814,N_25684,N_25622);
xnor U25815 (N_25815,N_25737,N_25766);
nor U25816 (N_25816,N_25636,N_25722);
or U25817 (N_25817,N_25610,N_25721);
or U25818 (N_25818,N_25775,N_25728);
xor U25819 (N_25819,N_25668,N_25790);
or U25820 (N_25820,N_25618,N_25769);
xor U25821 (N_25821,N_25715,N_25725);
nor U25822 (N_25822,N_25653,N_25617);
and U25823 (N_25823,N_25600,N_25757);
and U25824 (N_25824,N_25663,N_25754);
xnor U25825 (N_25825,N_25666,N_25793);
nand U25826 (N_25826,N_25623,N_25650);
nor U25827 (N_25827,N_25673,N_25798);
nand U25828 (N_25828,N_25780,N_25612);
nand U25829 (N_25829,N_25707,N_25664);
or U25830 (N_25830,N_25692,N_25629);
and U25831 (N_25831,N_25762,N_25603);
and U25832 (N_25832,N_25602,N_25723);
xnor U25833 (N_25833,N_25718,N_25687);
and U25834 (N_25834,N_25705,N_25767);
or U25835 (N_25835,N_25677,N_25631);
nand U25836 (N_25836,N_25759,N_25779);
or U25837 (N_25837,N_25736,N_25708);
xnor U25838 (N_25838,N_25686,N_25713);
xnor U25839 (N_25839,N_25761,N_25620);
or U25840 (N_25840,N_25787,N_25739);
nand U25841 (N_25841,N_25792,N_25797);
or U25842 (N_25842,N_25734,N_25672);
xnor U25843 (N_25843,N_25654,N_25614);
and U25844 (N_25844,N_25735,N_25699);
or U25845 (N_25845,N_25777,N_25764);
or U25846 (N_25846,N_25613,N_25695);
and U25847 (N_25847,N_25679,N_25724);
nor U25848 (N_25848,N_25742,N_25685);
nor U25849 (N_25849,N_25782,N_25791);
xnor U25850 (N_25850,N_25752,N_25635);
xor U25851 (N_25851,N_25675,N_25745);
and U25852 (N_25852,N_25604,N_25701);
nand U25853 (N_25853,N_25671,N_25640);
nor U25854 (N_25854,N_25693,N_25744);
and U25855 (N_25855,N_25659,N_25661);
or U25856 (N_25856,N_25678,N_25658);
xor U25857 (N_25857,N_25788,N_25696);
xor U25858 (N_25858,N_25674,N_25639);
nor U25859 (N_25859,N_25709,N_25616);
and U25860 (N_25860,N_25716,N_25726);
xnor U25861 (N_25861,N_25609,N_25633);
xor U25862 (N_25862,N_25748,N_25785);
or U25863 (N_25863,N_25732,N_25648);
nand U25864 (N_25864,N_25719,N_25637);
nand U25865 (N_25865,N_25711,N_25634);
nand U25866 (N_25866,N_25741,N_25649);
nand U25867 (N_25867,N_25772,N_25746);
nand U25868 (N_25868,N_25643,N_25717);
xnor U25869 (N_25869,N_25730,N_25784);
or U25870 (N_25870,N_25712,N_25608);
nor U25871 (N_25871,N_25743,N_25667);
xnor U25872 (N_25872,N_25776,N_25778);
or U25873 (N_25873,N_25763,N_25773);
nand U25874 (N_25874,N_25702,N_25647);
or U25875 (N_25875,N_25669,N_25795);
nand U25876 (N_25876,N_25680,N_25611);
nand U25877 (N_25877,N_25774,N_25755);
or U25878 (N_25878,N_25789,N_25652);
or U25879 (N_25879,N_25738,N_25770);
nor U25880 (N_25880,N_25670,N_25794);
xnor U25881 (N_25881,N_25781,N_25644);
or U25882 (N_25882,N_25656,N_25607);
xnor U25883 (N_25883,N_25689,N_25720);
nand U25884 (N_25884,N_25606,N_25630);
and U25885 (N_25885,N_25756,N_25706);
and U25886 (N_25886,N_25698,N_25796);
and U25887 (N_25887,N_25731,N_25747);
xor U25888 (N_25888,N_25683,N_25729);
and U25889 (N_25889,N_25657,N_25750);
and U25890 (N_25890,N_25682,N_25615);
nor U25891 (N_25891,N_25662,N_25624);
nand U25892 (N_25892,N_25626,N_25627);
or U25893 (N_25893,N_25690,N_25771);
nand U25894 (N_25894,N_25642,N_25783);
nor U25895 (N_25895,N_25765,N_25688);
nor U25896 (N_25896,N_25704,N_25628);
or U25897 (N_25897,N_25641,N_25691);
nand U25898 (N_25898,N_25733,N_25651);
and U25899 (N_25899,N_25753,N_25621);
xnor U25900 (N_25900,N_25787,N_25743);
and U25901 (N_25901,N_25746,N_25790);
nor U25902 (N_25902,N_25697,N_25667);
nand U25903 (N_25903,N_25607,N_25664);
nand U25904 (N_25904,N_25791,N_25753);
or U25905 (N_25905,N_25616,N_25658);
or U25906 (N_25906,N_25631,N_25705);
xor U25907 (N_25907,N_25622,N_25702);
nor U25908 (N_25908,N_25776,N_25705);
xor U25909 (N_25909,N_25741,N_25755);
and U25910 (N_25910,N_25679,N_25728);
nor U25911 (N_25911,N_25693,N_25674);
and U25912 (N_25912,N_25703,N_25632);
nand U25913 (N_25913,N_25638,N_25751);
nor U25914 (N_25914,N_25691,N_25648);
and U25915 (N_25915,N_25741,N_25681);
nor U25916 (N_25916,N_25617,N_25696);
nor U25917 (N_25917,N_25631,N_25799);
and U25918 (N_25918,N_25763,N_25645);
nor U25919 (N_25919,N_25687,N_25697);
xnor U25920 (N_25920,N_25711,N_25797);
nor U25921 (N_25921,N_25746,N_25642);
nand U25922 (N_25922,N_25738,N_25707);
nand U25923 (N_25923,N_25611,N_25701);
and U25924 (N_25924,N_25609,N_25738);
nand U25925 (N_25925,N_25636,N_25672);
nor U25926 (N_25926,N_25628,N_25693);
and U25927 (N_25927,N_25691,N_25746);
or U25928 (N_25928,N_25661,N_25733);
nor U25929 (N_25929,N_25648,N_25601);
and U25930 (N_25930,N_25730,N_25772);
or U25931 (N_25931,N_25621,N_25703);
nor U25932 (N_25932,N_25653,N_25790);
nand U25933 (N_25933,N_25750,N_25668);
or U25934 (N_25934,N_25746,N_25647);
xor U25935 (N_25935,N_25719,N_25651);
xnor U25936 (N_25936,N_25652,N_25782);
nor U25937 (N_25937,N_25649,N_25662);
and U25938 (N_25938,N_25608,N_25615);
nor U25939 (N_25939,N_25747,N_25633);
or U25940 (N_25940,N_25727,N_25642);
nor U25941 (N_25941,N_25602,N_25641);
nor U25942 (N_25942,N_25733,N_25694);
nand U25943 (N_25943,N_25699,N_25788);
nor U25944 (N_25944,N_25622,N_25628);
nor U25945 (N_25945,N_25687,N_25737);
or U25946 (N_25946,N_25674,N_25737);
nor U25947 (N_25947,N_25774,N_25777);
xnor U25948 (N_25948,N_25716,N_25623);
or U25949 (N_25949,N_25653,N_25766);
xor U25950 (N_25950,N_25639,N_25739);
xor U25951 (N_25951,N_25699,N_25707);
nor U25952 (N_25952,N_25616,N_25717);
and U25953 (N_25953,N_25761,N_25733);
and U25954 (N_25954,N_25625,N_25658);
xor U25955 (N_25955,N_25645,N_25785);
nor U25956 (N_25956,N_25791,N_25789);
nor U25957 (N_25957,N_25780,N_25764);
xor U25958 (N_25958,N_25793,N_25621);
nor U25959 (N_25959,N_25765,N_25644);
nor U25960 (N_25960,N_25767,N_25792);
and U25961 (N_25961,N_25799,N_25604);
nor U25962 (N_25962,N_25725,N_25787);
and U25963 (N_25963,N_25665,N_25763);
nand U25964 (N_25964,N_25656,N_25782);
nor U25965 (N_25965,N_25614,N_25612);
xnor U25966 (N_25966,N_25728,N_25751);
nand U25967 (N_25967,N_25737,N_25758);
or U25968 (N_25968,N_25665,N_25639);
nor U25969 (N_25969,N_25694,N_25767);
nor U25970 (N_25970,N_25724,N_25676);
or U25971 (N_25971,N_25794,N_25682);
or U25972 (N_25972,N_25751,N_25754);
nand U25973 (N_25973,N_25667,N_25770);
xor U25974 (N_25974,N_25766,N_25669);
nand U25975 (N_25975,N_25746,N_25611);
and U25976 (N_25976,N_25702,N_25733);
nand U25977 (N_25977,N_25767,N_25791);
nor U25978 (N_25978,N_25682,N_25710);
xnor U25979 (N_25979,N_25688,N_25695);
nor U25980 (N_25980,N_25635,N_25628);
nor U25981 (N_25981,N_25612,N_25777);
or U25982 (N_25982,N_25757,N_25786);
and U25983 (N_25983,N_25650,N_25654);
nor U25984 (N_25984,N_25781,N_25617);
nand U25985 (N_25985,N_25684,N_25697);
nor U25986 (N_25986,N_25616,N_25719);
nand U25987 (N_25987,N_25747,N_25758);
nor U25988 (N_25988,N_25718,N_25699);
nor U25989 (N_25989,N_25665,N_25644);
and U25990 (N_25990,N_25790,N_25788);
or U25991 (N_25991,N_25722,N_25689);
or U25992 (N_25992,N_25674,N_25785);
nor U25993 (N_25993,N_25673,N_25684);
xor U25994 (N_25994,N_25609,N_25681);
xnor U25995 (N_25995,N_25768,N_25783);
xnor U25996 (N_25996,N_25793,N_25731);
xnor U25997 (N_25997,N_25660,N_25694);
or U25998 (N_25998,N_25620,N_25771);
or U25999 (N_25999,N_25724,N_25633);
xnor U26000 (N_26000,N_25814,N_25955);
xnor U26001 (N_26001,N_25802,N_25941);
nor U26002 (N_26002,N_25811,N_25858);
nand U26003 (N_26003,N_25818,N_25987);
nor U26004 (N_26004,N_25888,N_25918);
and U26005 (N_26005,N_25835,N_25871);
nor U26006 (N_26006,N_25856,N_25898);
and U26007 (N_26007,N_25997,N_25966);
or U26008 (N_26008,N_25827,N_25976);
xor U26009 (N_26009,N_25885,N_25800);
nor U26010 (N_26010,N_25882,N_25971);
xor U26011 (N_26011,N_25833,N_25810);
nand U26012 (N_26012,N_25864,N_25916);
and U26013 (N_26013,N_25840,N_25960);
or U26014 (N_26014,N_25889,N_25896);
nand U26015 (N_26015,N_25958,N_25948);
nor U26016 (N_26016,N_25939,N_25875);
nand U26017 (N_26017,N_25934,N_25952);
or U26018 (N_26018,N_25846,N_25894);
nor U26019 (N_26019,N_25911,N_25857);
nor U26020 (N_26020,N_25999,N_25873);
nor U26021 (N_26021,N_25945,N_25947);
nand U26022 (N_26022,N_25957,N_25866);
nor U26023 (N_26023,N_25985,N_25849);
xnor U26024 (N_26024,N_25989,N_25932);
or U26025 (N_26025,N_25964,N_25988);
nand U26026 (N_26026,N_25965,N_25904);
or U26027 (N_26027,N_25986,N_25953);
and U26028 (N_26028,N_25915,N_25829);
nand U26029 (N_26029,N_25807,N_25900);
nor U26030 (N_26030,N_25920,N_25850);
nor U26031 (N_26031,N_25874,N_25867);
xor U26032 (N_26032,N_25862,N_25812);
xnor U26033 (N_26033,N_25891,N_25910);
and U26034 (N_26034,N_25907,N_25927);
or U26035 (N_26035,N_25984,N_25909);
nor U26036 (N_26036,N_25951,N_25847);
and U26037 (N_26037,N_25942,N_25809);
nor U26038 (N_26038,N_25923,N_25935);
nor U26039 (N_26039,N_25826,N_25962);
nand U26040 (N_26040,N_25969,N_25863);
or U26041 (N_26041,N_25876,N_25834);
nor U26042 (N_26042,N_25831,N_25933);
nand U26043 (N_26043,N_25973,N_25925);
or U26044 (N_26044,N_25819,N_25968);
nor U26045 (N_26045,N_25844,N_25924);
or U26046 (N_26046,N_25804,N_25956);
nand U26047 (N_26047,N_25914,N_25908);
xor U26048 (N_26048,N_25817,N_25901);
nor U26049 (N_26049,N_25949,N_25946);
or U26050 (N_26050,N_25893,N_25944);
or U26051 (N_26051,N_25816,N_25981);
or U26052 (N_26052,N_25899,N_25983);
nand U26053 (N_26053,N_25892,N_25998);
xor U26054 (N_26054,N_25852,N_25929);
nor U26055 (N_26055,N_25991,N_25839);
nor U26056 (N_26056,N_25980,N_25859);
xor U26057 (N_26057,N_25851,N_25886);
or U26058 (N_26058,N_25836,N_25903);
nand U26059 (N_26059,N_25975,N_25961);
and U26060 (N_26060,N_25992,N_25841);
nand U26061 (N_26061,N_25993,N_25887);
xnor U26062 (N_26062,N_25830,N_25895);
nor U26063 (N_26063,N_25865,N_25860);
and U26064 (N_26064,N_25912,N_25936);
and U26065 (N_26065,N_25902,N_25843);
nand U26066 (N_26066,N_25880,N_25878);
or U26067 (N_26067,N_25879,N_25825);
and U26068 (N_26068,N_25931,N_25813);
xnor U26069 (N_26069,N_25938,N_25978);
nand U26070 (N_26070,N_25832,N_25837);
nor U26071 (N_26071,N_25928,N_25820);
or U26072 (N_26072,N_25815,N_25838);
nand U26073 (N_26073,N_25982,N_25967);
or U26074 (N_26074,N_25996,N_25848);
xor U26075 (N_26075,N_25970,N_25854);
or U26076 (N_26076,N_25803,N_25919);
nand U26077 (N_26077,N_25979,N_25855);
or U26078 (N_26078,N_25897,N_25943);
or U26079 (N_26079,N_25995,N_25824);
and U26080 (N_26080,N_25921,N_25842);
xnor U26081 (N_26081,N_25872,N_25884);
nand U26082 (N_26082,N_25974,N_25861);
or U26083 (N_26083,N_25977,N_25883);
nor U26084 (N_26084,N_25926,N_25917);
and U26085 (N_26085,N_25950,N_25930);
and U26086 (N_26086,N_25845,N_25922);
or U26087 (N_26087,N_25853,N_25808);
xnor U26088 (N_26088,N_25890,N_25905);
or U26089 (N_26089,N_25906,N_25954);
or U26090 (N_26090,N_25913,N_25877);
or U26091 (N_26091,N_25869,N_25990);
or U26092 (N_26092,N_25823,N_25963);
xnor U26093 (N_26093,N_25937,N_25806);
nor U26094 (N_26094,N_25805,N_25828);
xor U26095 (N_26095,N_25821,N_25868);
xor U26096 (N_26096,N_25801,N_25994);
nand U26097 (N_26097,N_25959,N_25940);
xnor U26098 (N_26098,N_25870,N_25972);
nor U26099 (N_26099,N_25822,N_25881);
and U26100 (N_26100,N_25818,N_25923);
and U26101 (N_26101,N_25870,N_25837);
nand U26102 (N_26102,N_25957,N_25966);
xor U26103 (N_26103,N_25920,N_25911);
or U26104 (N_26104,N_25968,N_25993);
xor U26105 (N_26105,N_25898,N_25827);
or U26106 (N_26106,N_25907,N_25890);
nand U26107 (N_26107,N_25844,N_25886);
or U26108 (N_26108,N_25924,N_25898);
nand U26109 (N_26109,N_25880,N_25948);
nand U26110 (N_26110,N_25801,N_25823);
xor U26111 (N_26111,N_25902,N_25962);
nand U26112 (N_26112,N_25851,N_25859);
and U26113 (N_26113,N_25973,N_25949);
nor U26114 (N_26114,N_25949,N_25858);
and U26115 (N_26115,N_25912,N_25885);
nor U26116 (N_26116,N_25986,N_25923);
or U26117 (N_26117,N_25956,N_25909);
nor U26118 (N_26118,N_25898,N_25901);
or U26119 (N_26119,N_25802,N_25883);
nor U26120 (N_26120,N_25848,N_25913);
xor U26121 (N_26121,N_25881,N_25925);
and U26122 (N_26122,N_25989,N_25804);
nor U26123 (N_26123,N_25997,N_25922);
nand U26124 (N_26124,N_25960,N_25945);
nand U26125 (N_26125,N_25908,N_25935);
or U26126 (N_26126,N_25828,N_25818);
nand U26127 (N_26127,N_25852,N_25897);
nand U26128 (N_26128,N_25889,N_25965);
nand U26129 (N_26129,N_25977,N_25844);
xor U26130 (N_26130,N_25861,N_25918);
and U26131 (N_26131,N_25950,N_25851);
xor U26132 (N_26132,N_25907,N_25803);
or U26133 (N_26133,N_25899,N_25966);
xnor U26134 (N_26134,N_25843,N_25848);
nor U26135 (N_26135,N_25938,N_25821);
nor U26136 (N_26136,N_25933,N_25824);
xor U26137 (N_26137,N_25800,N_25918);
or U26138 (N_26138,N_25866,N_25817);
and U26139 (N_26139,N_25823,N_25889);
nor U26140 (N_26140,N_25969,N_25893);
or U26141 (N_26141,N_25827,N_25916);
or U26142 (N_26142,N_25866,N_25998);
nor U26143 (N_26143,N_25849,N_25995);
or U26144 (N_26144,N_25824,N_25935);
nor U26145 (N_26145,N_25902,N_25910);
or U26146 (N_26146,N_25800,N_25852);
xor U26147 (N_26147,N_25986,N_25909);
nand U26148 (N_26148,N_25855,N_25922);
nor U26149 (N_26149,N_25935,N_25919);
nor U26150 (N_26150,N_25926,N_25956);
xnor U26151 (N_26151,N_25953,N_25907);
xor U26152 (N_26152,N_25906,N_25937);
nand U26153 (N_26153,N_25991,N_25807);
xor U26154 (N_26154,N_25979,N_25807);
or U26155 (N_26155,N_25968,N_25878);
nor U26156 (N_26156,N_25968,N_25942);
and U26157 (N_26157,N_25960,N_25935);
or U26158 (N_26158,N_25910,N_25819);
and U26159 (N_26159,N_25899,N_25896);
or U26160 (N_26160,N_25949,N_25874);
and U26161 (N_26161,N_25898,N_25909);
xor U26162 (N_26162,N_25938,N_25900);
nor U26163 (N_26163,N_25966,N_25939);
nand U26164 (N_26164,N_25821,N_25964);
nand U26165 (N_26165,N_25911,N_25890);
xnor U26166 (N_26166,N_25808,N_25973);
nor U26167 (N_26167,N_25964,N_25922);
nand U26168 (N_26168,N_25912,N_25920);
nor U26169 (N_26169,N_25827,N_25832);
xnor U26170 (N_26170,N_25852,N_25878);
and U26171 (N_26171,N_25821,N_25865);
or U26172 (N_26172,N_25943,N_25851);
and U26173 (N_26173,N_25817,N_25806);
nor U26174 (N_26174,N_25803,N_25870);
and U26175 (N_26175,N_25996,N_25881);
nor U26176 (N_26176,N_25981,N_25970);
nand U26177 (N_26177,N_25818,N_25813);
nor U26178 (N_26178,N_25861,N_25958);
and U26179 (N_26179,N_25905,N_25896);
nor U26180 (N_26180,N_25817,N_25891);
xnor U26181 (N_26181,N_25853,N_25859);
nor U26182 (N_26182,N_25996,N_25861);
nand U26183 (N_26183,N_25892,N_25908);
nor U26184 (N_26184,N_25882,N_25809);
or U26185 (N_26185,N_25891,N_25955);
and U26186 (N_26186,N_25936,N_25919);
nand U26187 (N_26187,N_25893,N_25885);
and U26188 (N_26188,N_25827,N_25926);
xnor U26189 (N_26189,N_25826,N_25929);
or U26190 (N_26190,N_25840,N_25955);
or U26191 (N_26191,N_25816,N_25847);
xnor U26192 (N_26192,N_25936,N_25907);
nand U26193 (N_26193,N_25987,N_25919);
nand U26194 (N_26194,N_25981,N_25857);
xor U26195 (N_26195,N_25954,N_25963);
nand U26196 (N_26196,N_25848,N_25919);
xnor U26197 (N_26197,N_25930,N_25999);
or U26198 (N_26198,N_25821,N_25958);
xnor U26199 (N_26199,N_25915,N_25939);
xor U26200 (N_26200,N_26037,N_26081);
xnor U26201 (N_26201,N_26099,N_26087);
or U26202 (N_26202,N_26086,N_26182);
nor U26203 (N_26203,N_26180,N_26079);
nor U26204 (N_26204,N_26015,N_26193);
and U26205 (N_26205,N_26160,N_26027);
xnor U26206 (N_26206,N_26060,N_26016);
and U26207 (N_26207,N_26006,N_26185);
nand U26208 (N_26208,N_26018,N_26032);
and U26209 (N_26209,N_26052,N_26048);
or U26210 (N_26210,N_26197,N_26059);
xnor U26211 (N_26211,N_26157,N_26108);
nand U26212 (N_26212,N_26111,N_26046);
or U26213 (N_26213,N_26176,N_26192);
nor U26214 (N_26214,N_26088,N_26025);
and U26215 (N_26215,N_26136,N_26011);
or U26216 (N_26216,N_26061,N_26063);
nand U26217 (N_26217,N_26071,N_26023);
and U26218 (N_26218,N_26098,N_26198);
and U26219 (N_26219,N_26004,N_26047);
nand U26220 (N_26220,N_26090,N_26077);
nor U26221 (N_26221,N_26150,N_26091);
and U26222 (N_26222,N_26095,N_26158);
nor U26223 (N_26223,N_26043,N_26021);
nor U26224 (N_26224,N_26128,N_26041);
and U26225 (N_26225,N_26075,N_26138);
nor U26226 (N_26226,N_26042,N_26119);
and U26227 (N_26227,N_26170,N_26070);
nor U26228 (N_26228,N_26068,N_26029);
nor U26229 (N_26229,N_26163,N_26057);
and U26230 (N_26230,N_26147,N_26105);
nand U26231 (N_26231,N_26020,N_26024);
xor U26232 (N_26232,N_26114,N_26199);
nand U26233 (N_26233,N_26159,N_26137);
nand U26234 (N_26234,N_26194,N_26034);
nor U26235 (N_26235,N_26195,N_26022);
nand U26236 (N_26236,N_26053,N_26118);
nand U26237 (N_26237,N_26165,N_26151);
and U26238 (N_26238,N_26100,N_26003);
nor U26239 (N_26239,N_26177,N_26104);
xor U26240 (N_26240,N_26149,N_26115);
xnor U26241 (N_26241,N_26183,N_26000);
and U26242 (N_26242,N_26035,N_26175);
xnor U26243 (N_26243,N_26085,N_26191);
or U26244 (N_26244,N_26155,N_26141);
nand U26245 (N_26245,N_26164,N_26110);
xor U26246 (N_26246,N_26145,N_26044);
or U26247 (N_26247,N_26066,N_26002);
and U26248 (N_26248,N_26133,N_26084);
nor U26249 (N_26249,N_26161,N_26083);
and U26250 (N_26250,N_26186,N_26102);
or U26251 (N_26251,N_26116,N_26196);
and U26252 (N_26252,N_26174,N_26031);
and U26253 (N_26253,N_26168,N_26033);
or U26254 (N_26254,N_26139,N_26117);
and U26255 (N_26255,N_26039,N_26167);
nand U26256 (N_26256,N_26126,N_26062);
xor U26257 (N_26257,N_26096,N_26067);
xnor U26258 (N_26258,N_26012,N_26154);
nor U26259 (N_26259,N_26120,N_26181);
nand U26260 (N_26260,N_26040,N_26072);
nand U26261 (N_26261,N_26045,N_26010);
or U26262 (N_26262,N_26184,N_26188);
xnor U26263 (N_26263,N_26055,N_26038);
nand U26264 (N_26264,N_26132,N_26152);
and U26265 (N_26265,N_26054,N_26028);
xnor U26266 (N_26266,N_26142,N_26166);
and U26267 (N_26267,N_26172,N_26008);
xnor U26268 (N_26268,N_26121,N_26146);
xnor U26269 (N_26269,N_26007,N_26065);
or U26270 (N_26270,N_26156,N_26162);
xor U26271 (N_26271,N_26179,N_26169);
or U26272 (N_26272,N_26171,N_26106);
or U26273 (N_26273,N_26049,N_26078);
or U26274 (N_26274,N_26076,N_26135);
and U26275 (N_26275,N_26190,N_26127);
nor U26276 (N_26276,N_26080,N_26030);
and U26277 (N_26277,N_26092,N_26093);
and U26278 (N_26278,N_26073,N_26148);
nand U26279 (N_26279,N_26005,N_26129);
nor U26280 (N_26280,N_26189,N_26109);
nor U26281 (N_26281,N_26074,N_26014);
or U26282 (N_26282,N_26122,N_26153);
or U26283 (N_26283,N_26173,N_26140);
xor U26284 (N_26284,N_26019,N_26107);
and U26285 (N_26285,N_26089,N_26058);
nor U26286 (N_26286,N_26009,N_26130);
and U26287 (N_26287,N_26097,N_26094);
xor U26288 (N_26288,N_26056,N_26101);
nand U26289 (N_26289,N_26112,N_26036);
xor U26290 (N_26290,N_26131,N_26017);
nand U26291 (N_26291,N_26187,N_26051);
xor U26292 (N_26292,N_26123,N_26069);
nor U26293 (N_26293,N_26178,N_26113);
nor U26294 (N_26294,N_26013,N_26001);
or U26295 (N_26295,N_26026,N_26082);
nor U26296 (N_26296,N_26144,N_26125);
or U26297 (N_26297,N_26103,N_26064);
nand U26298 (N_26298,N_26124,N_26134);
nand U26299 (N_26299,N_26050,N_26143);
nand U26300 (N_26300,N_26142,N_26009);
nand U26301 (N_26301,N_26100,N_26076);
and U26302 (N_26302,N_26054,N_26116);
nor U26303 (N_26303,N_26154,N_26077);
xor U26304 (N_26304,N_26153,N_26011);
nand U26305 (N_26305,N_26013,N_26194);
and U26306 (N_26306,N_26068,N_26180);
or U26307 (N_26307,N_26072,N_26096);
or U26308 (N_26308,N_26011,N_26195);
and U26309 (N_26309,N_26143,N_26170);
xor U26310 (N_26310,N_26036,N_26021);
and U26311 (N_26311,N_26040,N_26185);
nor U26312 (N_26312,N_26044,N_26027);
nor U26313 (N_26313,N_26037,N_26047);
or U26314 (N_26314,N_26134,N_26082);
nor U26315 (N_26315,N_26020,N_26001);
nand U26316 (N_26316,N_26092,N_26080);
or U26317 (N_26317,N_26147,N_26163);
or U26318 (N_26318,N_26124,N_26054);
and U26319 (N_26319,N_26073,N_26132);
nand U26320 (N_26320,N_26131,N_26144);
or U26321 (N_26321,N_26048,N_26127);
or U26322 (N_26322,N_26113,N_26198);
and U26323 (N_26323,N_26036,N_26038);
or U26324 (N_26324,N_26147,N_26119);
xnor U26325 (N_26325,N_26052,N_26018);
xnor U26326 (N_26326,N_26045,N_26133);
or U26327 (N_26327,N_26102,N_26145);
or U26328 (N_26328,N_26189,N_26191);
nor U26329 (N_26329,N_26081,N_26059);
and U26330 (N_26330,N_26028,N_26173);
or U26331 (N_26331,N_26034,N_26099);
or U26332 (N_26332,N_26110,N_26056);
xnor U26333 (N_26333,N_26119,N_26086);
or U26334 (N_26334,N_26178,N_26183);
or U26335 (N_26335,N_26057,N_26173);
nor U26336 (N_26336,N_26094,N_26124);
xnor U26337 (N_26337,N_26049,N_26081);
nor U26338 (N_26338,N_26138,N_26141);
nand U26339 (N_26339,N_26145,N_26056);
or U26340 (N_26340,N_26197,N_26079);
nor U26341 (N_26341,N_26167,N_26193);
or U26342 (N_26342,N_26121,N_26127);
or U26343 (N_26343,N_26108,N_26152);
nand U26344 (N_26344,N_26113,N_26196);
and U26345 (N_26345,N_26151,N_26183);
or U26346 (N_26346,N_26127,N_26077);
and U26347 (N_26347,N_26160,N_26101);
nor U26348 (N_26348,N_26181,N_26160);
or U26349 (N_26349,N_26190,N_26023);
xor U26350 (N_26350,N_26102,N_26162);
nor U26351 (N_26351,N_26110,N_26054);
nor U26352 (N_26352,N_26026,N_26104);
and U26353 (N_26353,N_26021,N_26121);
nand U26354 (N_26354,N_26112,N_26119);
or U26355 (N_26355,N_26187,N_26029);
xor U26356 (N_26356,N_26091,N_26146);
nand U26357 (N_26357,N_26154,N_26061);
or U26358 (N_26358,N_26196,N_26176);
and U26359 (N_26359,N_26112,N_26101);
or U26360 (N_26360,N_26020,N_26065);
or U26361 (N_26361,N_26162,N_26194);
nor U26362 (N_26362,N_26076,N_26035);
xor U26363 (N_26363,N_26199,N_26033);
and U26364 (N_26364,N_26010,N_26073);
or U26365 (N_26365,N_26182,N_26138);
nand U26366 (N_26366,N_26103,N_26120);
and U26367 (N_26367,N_26052,N_26010);
nor U26368 (N_26368,N_26194,N_26093);
xor U26369 (N_26369,N_26037,N_26124);
xor U26370 (N_26370,N_26107,N_26067);
nor U26371 (N_26371,N_26103,N_26186);
or U26372 (N_26372,N_26188,N_26003);
or U26373 (N_26373,N_26070,N_26064);
or U26374 (N_26374,N_26011,N_26198);
and U26375 (N_26375,N_26196,N_26014);
nor U26376 (N_26376,N_26084,N_26105);
xor U26377 (N_26377,N_26045,N_26141);
nor U26378 (N_26378,N_26044,N_26084);
nor U26379 (N_26379,N_26096,N_26113);
and U26380 (N_26380,N_26072,N_26157);
nand U26381 (N_26381,N_26064,N_26107);
and U26382 (N_26382,N_26113,N_26186);
nand U26383 (N_26383,N_26063,N_26126);
and U26384 (N_26384,N_26065,N_26073);
xor U26385 (N_26385,N_26025,N_26017);
or U26386 (N_26386,N_26026,N_26119);
nand U26387 (N_26387,N_26179,N_26166);
and U26388 (N_26388,N_26113,N_26002);
nor U26389 (N_26389,N_26046,N_26043);
nor U26390 (N_26390,N_26145,N_26046);
and U26391 (N_26391,N_26063,N_26084);
xnor U26392 (N_26392,N_26123,N_26016);
nor U26393 (N_26393,N_26018,N_26102);
nor U26394 (N_26394,N_26018,N_26019);
nand U26395 (N_26395,N_26063,N_26117);
or U26396 (N_26396,N_26049,N_26071);
or U26397 (N_26397,N_26164,N_26058);
or U26398 (N_26398,N_26099,N_26176);
and U26399 (N_26399,N_26083,N_26065);
nor U26400 (N_26400,N_26221,N_26290);
xor U26401 (N_26401,N_26267,N_26257);
nand U26402 (N_26402,N_26323,N_26232);
nand U26403 (N_26403,N_26201,N_26295);
nand U26404 (N_26404,N_26256,N_26294);
xnor U26405 (N_26405,N_26377,N_26331);
or U26406 (N_26406,N_26247,N_26214);
nand U26407 (N_26407,N_26398,N_26246);
and U26408 (N_26408,N_26272,N_26355);
xnor U26409 (N_26409,N_26207,N_26315);
nand U26410 (N_26410,N_26324,N_26284);
and U26411 (N_26411,N_26329,N_26371);
or U26412 (N_26412,N_26236,N_26305);
nand U26413 (N_26413,N_26343,N_26309);
nor U26414 (N_26414,N_26227,N_26291);
nand U26415 (N_26415,N_26338,N_26361);
nor U26416 (N_26416,N_26359,N_26357);
nor U26417 (N_26417,N_26336,N_26314);
xnor U26418 (N_26418,N_26226,N_26333);
nor U26419 (N_26419,N_26362,N_26360);
and U26420 (N_26420,N_26386,N_26238);
nand U26421 (N_26421,N_26202,N_26328);
or U26422 (N_26422,N_26397,N_26234);
nor U26423 (N_26423,N_26363,N_26356);
nor U26424 (N_26424,N_26235,N_26379);
or U26425 (N_26425,N_26337,N_26270);
or U26426 (N_26426,N_26297,N_26348);
nor U26427 (N_26427,N_26277,N_26203);
or U26428 (N_26428,N_26366,N_26384);
xor U26429 (N_26429,N_26399,N_26390);
and U26430 (N_26430,N_26392,N_26320);
nor U26431 (N_26431,N_26223,N_26326);
xor U26432 (N_26432,N_26387,N_26391);
nand U26433 (N_26433,N_26293,N_26354);
nor U26434 (N_26434,N_26322,N_26298);
xnor U26435 (N_26435,N_26358,N_26266);
nand U26436 (N_26436,N_26282,N_26306);
nor U26437 (N_26437,N_26327,N_26375);
xnor U26438 (N_26438,N_26222,N_26278);
nor U26439 (N_26439,N_26318,N_26292);
nor U26440 (N_26440,N_26310,N_26313);
or U26441 (N_26441,N_26239,N_26204);
and U26442 (N_26442,N_26319,N_26243);
nor U26443 (N_26443,N_26273,N_26385);
and U26444 (N_26444,N_26342,N_26286);
nor U26445 (N_26445,N_26351,N_26210);
and U26446 (N_26446,N_26265,N_26353);
or U26447 (N_26447,N_26347,N_26251);
nor U26448 (N_26448,N_26248,N_26261);
or U26449 (N_26449,N_26219,N_26276);
xor U26450 (N_26450,N_26296,N_26394);
nor U26451 (N_26451,N_26301,N_26395);
nor U26452 (N_26452,N_26285,N_26346);
and U26453 (N_26453,N_26264,N_26280);
and U26454 (N_26454,N_26349,N_26378);
or U26455 (N_26455,N_26289,N_26206);
xnor U26456 (N_26456,N_26317,N_26245);
or U26457 (N_26457,N_26274,N_26209);
and U26458 (N_26458,N_26269,N_26205);
or U26459 (N_26459,N_26240,N_26255);
or U26460 (N_26460,N_26350,N_26259);
nand U26461 (N_26461,N_26254,N_26241);
or U26462 (N_26462,N_26340,N_26367);
nand U26463 (N_26463,N_26263,N_26224);
xor U26464 (N_26464,N_26321,N_26258);
nand U26465 (N_26465,N_26396,N_26370);
and U26466 (N_26466,N_26271,N_26368);
or U26467 (N_26467,N_26299,N_26303);
xnor U26468 (N_26468,N_26381,N_26288);
or U26469 (N_26469,N_26339,N_26218);
nand U26470 (N_26470,N_26262,N_26307);
nor U26471 (N_26471,N_26200,N_26228);
nand U26472 (N_26472,N_26325,N_26389);
nor U26473 (N_26473,N_26260,N_26283);
nor U26474 (N_26474,N_26345,N_26330);
and U26475 (N_26475,N_26253,N_26300);
nand U26476 (N_26476,N_26388,N_26217);
nand U26477 (N_26477,N_26279,N_26334);
xor U26478 (N_26478,N_26275,N_26304);
xor U26479 (N_26479,N_26244,N_26211);
or U26480 (N_26480,N_26220,N_26312);
xnor U26481 (N_26481,N_26281,N_26225);
or U26482 (N_26482,N_26216,N_26369);
or U26483 (N_26483,N_26373,N_26382);
or U26484 (N_26484,N_26365,N_26233);
nand U26485 (N_26485,N_26344,N_26268);
nand U26486 (N_26486,N_26237,N_26252);
nor U26487 (N_26487,N_26332,N_26249);
nor U26488 (N_26488,N_26393,N_26308);
or U26489 (N_26489,N_26372,N_26380);
or U26490 (N_26490,N_26213,N_26383);
nor U26491 (N_26491,N_26231,N_26230);
or U26492 (N_26492,N_26212,N_26229);
xnor U26493 (N_26493,N_26374,N_26316);
and U26494 (N_26494,N_26242,N_26364);
xnor U26495 (N_26495,N_26302,N_26287);
or U26496 (N_26496,N_26335,N_26311);
nand U26497 (N_26497,N_26215,N_26341);
nor U26498 (N_26498,N_26250,N_26376);
or U26499 (N_26499,N_26352,N_26208);
or U26500 (N_26500,N_26238,N_26223);
xnor U26501 (N_26501,N_26247,N_26218);
nor U26502 (N_26502,N_26310,N_26392);
nand U26503 (N_26503,N_26390,N_26256);
or U26504 (N_26504,N_26345,N_26213);
nor U26505 (N_26505,N_26278,N_26246);
nor U26506 (N_26506,N_26388,N_26307);
nor U26507 (N_26507,N_26239,N_26223);
xnor U26508 (N_26508,N_26244,N_26254);
or U26509 (N_26509,N_26315,N_26236);
nor U26510 (N_26510,N_26234,N_26252);
nand U26511 (N_26511,N_26265,N_26307);
nor U26512 (N_26512,N_26354,N_26303);
xor U26513 (N_26513,N_26254,N_26345);
or U26514 (N_26514,N_26200,N_26218);
or U26515 (N_26515,N_26308,N_26390);
xnor U26516 (N_26516,N_26368,N_26348);
nand U26517 (N_26517,N_26229,N_26356);
xnor U26518 (N_26518,N_26256,N_26230);
and U26519 (N_26519,N_26221,N_26389);
xnor U26520 (N_26520,N_26377,N_26393);
nand U26521 (N_26521,N_26299,N_26368);
nand U26522 (N_26522,N_26227,N_26355);
nor U26523 (N_26523,N_26201,N_26350);
or U26524 (N_26524,N_26241,N_26390);
nand U26525 (N_26525,N_26280,N_26277);
nand U26526 (N_26526,N_26274,N_26391);
and U26527 (N_26527,N_26245,N_26354);
or U26528 (N_26528,N_26274,N_26251);
and U26529 (N_26529,N_26308,N_26350);
and U26530 (N_26530,N_26299,N_26302);
and U26531 (N_26531,N_26349,N_26220);
or U26532 (N_26532,N_26201,N_26376);
or U26533 (N_26533,N_26293,N_26204);
nor U26534 (N_26534,N_26235,N_26222);
or U26535 (N_26535,N_26266,N_26310);
nor U26536 (N_26536,N_26230,N_26238);
and U26537 (N_26537,N_26256,N_26300);
xor U26538 (N_26538,N_26327,N_26200);
or U26539 (N_26539,N_26335,N_26254);
or U26540 (N_26540,N_26343,N_26390);
and U26541 (N_26541,N_26389,N_26213);
and U26542 (N_26542,N_26216,N_26242);
xnor U26543 (N_26543,N_26377,N_26323);
xnor U26544 (N_26544,N_26398,N_26366);
and U26545 (N_26545,N_26273,N_26223);
xnor U26546 (N_26546,N_26360,N_26206);
nand U26547 (N_26547,N_26324,N_26320);
and U26548 (N_26548,N_26351,N_26355);
nor U26549 (N_26549,N_26205,N_26399);
nor U26550 (N_26550,N_26391,N_26292);
xnor U26551 (N_26551,N_26316,N_26399);
or U26552 (N_26552,N_26250,N_26373);
xnor U26553 (N_26553,N_26308,N_26337);
and U26554 (N_26554,N_26210,N_26353);
or U26555 (N_26555,N_26347,N_26284);
nand U26556 (N_26556,N_26289,N_26305);
nand U26557 (N_26557,N_26277,N_26244);
or U26558 (N_26558,N_26345,N_26231);
nand U26559 (N_26559,N_26321,N_26283);
and U26560 (N_26560,N_26269,N_26399);
and U26561 (N_26561,N_26271,N_26258);
xnor U26562 (N_26562,N_26262,N_26391);
nor U26563 (N_26563,N_26324,N_26281);
xor U26564 (N_26564,N_26395,N_26260);
nor U26565 (N_26565,N_26335,N_26299);
or U26566 (N_26566,N_26272,N_26385);
xor U26567 (N_26567,N_26228,N_26297);
and U26568 (N_26568,N_26382,N_26398);
xor U26569 (N_26569,N_26326,N_26383);
xnor U26570 (N_26570,N_26349,N_26323);
xnor U26571 (N_26571,N_26281,N_26201);
or U26572 (N_26572,N_26344,N_26302);
nand U26573 (N_26573,N_26341,N_26392);
nor U26574 (N_26574,N_26308,N_26311);
and U26575 (N_26575,N_26257,N_26214);
and U26576 (N_26576,N_26386,N_26226);
or U26577 (N_26577,N_26205,N_26345);
nand U26578 (N_26578,N_26357,N_26264);
nand U26579 (N_26579,N_26314,N_26332);
xor U26580 (N_26580,N_26227,N_26280);
and U26581 (N_26581,N_26269,N_26244);
or U26582 (N_26582,N_26275,N_26234);
or U26583 (N_26583,N_26374,N_26375);
and U26584 (N_26584,N_26296,N_26242);
nor U26585 (N_26585,N_26391,N_26247);
xnor U26586 (N_26586,N_26376,N_26317);
or U26587 (N_26587,N_26226,N_26283);
or U26588 (N_26588,N_26294,N_26285);
xor U26589 (N_26589,N_26259,N_26376);
nor U26590 (N_26590,N_26203,N_26263);
and U26591 (N_26591,N_26281,N_26275);
nor U26592 (N_26592,N_26396,N_26302);
and U26593 (N_26593,N_26391,N_26356);
nand U26594 (N_26594,N_26327,N_26293);
and U26595 (N_26595,N_26346,N_26269);
nor U26596 (N_26596,N_26386,N_26369);
xor U26597 (N_26597,N_26208,N_26264);
nor U26598 (N_26598,N_26271,N_26207);
nor U26599 (N_26599,N_26235,N_26345);
or U26600 (N_26600,N_26493,N_26536);
xnor U26601 (N_26601,N_26404,N_26503);
nand U26602 (N_26602,N_26518,N_26446);
or U26603 (N_26603,N_26474,N_26579);
nor U26604 (N_26604,N_26409,N_26531);
xnor U26605 (N_26605,N_26402,N_26436);
nor U26606 (N_26606,N_26408,N_26471);
or U26607 (N_26607,N_26459,N_26547);
nand U26608 (N_26608,N_26560,N_26400);
nor U26609 (N_26609,N_26424,N_26407);
or U26610 (N_26610,N_26438,N_26462);
xnor U26611 (N_26611,N_26458,N_26585);
nand U26612 (N_26612,N_26555,N_26559);
xor U26613 (N_26613,N_26577,N_26440);
nand U26614 (N_26614,N_26535,N_26401);
nand U26615 (N_26615,N_26479,N_26496);
nor U26616 (N_26616,N_26550,N_26466);
xor U26617 (N_26617,N_26476,N_26472);
or U26618 (N_26618,N_26425,N_26580);
or U26619 (N_26619,N_26565,N_26539);
and U26620 (N_26620,N_26428,N_26467);
nand U26621 (N_26621,N_26522,N_26500);
nand U26622 (N_26622,N_26574,N_26514);
and U26623 (N_26623,N_26418,N_26566);
or U26624 (N_26624,N_26567,N_26598);
or U26625 (N_26625,N_26572,N_26526);
or U26626 (N_26626,N_26501,N_26506);
or U26627 (N_26627,N_26413,N_26412);
nor U26628 (N_26628,N_26557,N_26530);
nor U26629 (N_26629,N_26549,N_26406);
xnor U26630 (N_26630,N_26517,N_26461);
and U26631 (N_26631,N_26449,N_26582);
and U26632 (N_26632,N_26590,N_26468);
nand U26633 (N_26633,N_26544,N_26502);
nand U26634 (N_26634,N_26504,N_26521);
and U26635 (N_26635,N_26511,N_26581);
or U26636 (N_26636,N_26548,N_26507);
nand U26637 (N_26637,N_26469,N_26515);
nor U26638 (N_26638,N_26450,N_26498);
xor U26639 (N_26639,N_26437,N_26587);
and U26640 (N_26640,N_26525,N_26519);
nor U26641 (N_26641,N_26588,N_26433);
and U26642 (N_26642,N_26516,N_26512);
and U26643 (N_26643,N_26552,N_26495);
and U26644 (N_26644,N_26529,N_26543);
xor U26645 (N_26645,N_26403,N_26455);
xor U26646 (N_26646,N_26465,N_26571);
or U26647 (N_26647,N_26509,N_26435);
nand U26648 (N_26648,N_26480,N_26451);
xor U26649 (N_26649,N_26597,N_26575);
nor U26650 (N_26650,N_26532,N_26494);
or U26651 (N_26651,N_26593,N_26563);
nand U26652 (N_26652,N_26594,N_26473);
and U26653 (N_26653,N_26528,N_26464);
xor U26654 (N_26654,N_26420,N_26524);
xnor U26655 (N_26655,N_26460,N_26452);
xnor U26656 (N_26656,N_26538,N_26554);
nor U26657 (N_26657,N_26444,N_26540);
and U26658 (N_26658,N_26520,N_26589);
xor U26659 (N_26659,N_26475,N_26583);
xor U26660 (N_26660,N_26569,N_26421);
xnor U26661 (N_26661,N_26426,N_26499);
nand U26662 (N_26662,N_26488,N_26445);
and U26663 (N_26663,N_26595,N_26564);
nand U26664 (N_26664,N_26423,N_26576);
and U26665 (N_26665,N_26483,N_26553);
and U26666 (N_26666,N_26591,N_26596);
or U26667 (N_26667,N_26430,N_26411);
xor U26668 (N_26668,N_26492,N_26546);
xnor U26669 (N_26669,N_26545,N_26523);
nand U26670 (N_26670,N_26478,N_26584);
nor U26671 (N_26671,N_26434,N_26482);
nor U26672 (N_26672,N_26537,N_26586);
nand U26673 (N_26673,N_26463,N_26562);
xnor U26674 (N_26674,N_26447,N_26573);
or U26675 (N_26675,N_26419,N_26416);
nor U26676 (N_26676,N_26487,N_26510);
and U26677 (N_26677,N_26497,N_26551);
nand U26678 (N_26678,N_26448,N_26417);
and U26679 (N_26679,N_26542,N_26527);
and U26680 (N_26680,N_26442,N_26456);
and U26681 (N_26681,N_26568,N_26481);
xnor U26682 (N_26682,N_26592,N_26570);
and U26683 (N_26683,N_26453,N_26484);
nor U26684 (N_26684,N_26489,N_26534);
xnor U26685 (N_26685,N_26439,N_26505);
xor U26686 (N_26686,N_26541,N_26429);
nand U26687 (N_26687,N_26533,N_26561);
xnor U26688 (N_26688,N_26441,N_26431);
and U26689 (N_26689,N_26599,N_26477);
and U26690 (N_26690,N_26415,N_26405);
and U26691 (N_26691,N_26432,N_26410);
or U26692 (N_26692,N_26490,N_26558);
xor U26693 (N_26693,N_26485,N_26486);
nand U26694 (N_26694,N_26443,N_26556);
and U26695 (N_26695,N_26470,N_26422);
nand U26696 (N_26696,N_26414,N_26427);
xnor U26697 (N_26697,N_26513,N_26491);
nor U26698 (N_26698,N_26454,N_26508);
nand U26699 (N_26699,N_26578,N_26457);
xnor U26700 (N_26700,N_26595,N_26541);
or U26701 (N_26701,N_26475,N_26562);
xor U26702 (N_26702,N_26542,N_26485);
or U26703 (N_26703,N_26566,N_26427);
xor U26704 (N_26704,N_26476,N_26467);
nand U26705 (N_26705,N_26456,N_26555);
or U26706 (N_26706,N_26505,N_26574);
xnor U26707 (N_26707,N_26558,N_26573);
or U26708 (N_26708,N_26587,N_26494);
and U26709 (N_26709,N_26586,N_26419);
nand U26710 (N_26710,N_26585,N_26521);
nor U26711 (N_26711,N_26502,N_26475);
nor U26712 (N_26712,N_26506,N_26519);
nand U26713 (N_26713,N_26563,N_26415);
nor U26714 (N_26714,N_26531,N_26405);
nor U26715 (N_26715,N_26446,N_26538);
and U26716 (N_26716,N_26595,N_26480);
and U26717 (N_26717,N_26446,N_26577);
nor U26718 (N_26718,N_26535,N_26550);
xnor U26719 (N_26719,N_26511,N_26416);
and U26720 (N_26720,N_26580,N_26576);
and U26721 (N_26721,N_26406,N_26450);
or U26722 (N_26722,N_26414,N_26514);
and U26723 (N_26723,N_26460,N_26448);
or U26724 (N_26724,N_26443,N_26476);
or U26725 (N_26725,N_26526,N_26457);
nand U26726 (N_26726,N_26454,N_26498);
xnor U26727 (N_26727,N_26422,N_26487);
nor U26728 (N_26728,N_26583,N_26578);
and U26729 (N_26729,N_26528,N_26462);
or U26730 (N_26730,N_26572,N_26594);
nand U26731 (N_26731,N_26474,N_26584);
or U26732 (N_26732,N_26410,N_26493);
nor U26733 (N_26733,N_26541,N_26467);
and U26734 (N_26734,N_26485,N_26523);
or U26735 (N_26735,N_26563,N_26533);
xnor U26736 (N_26736,N_26548,N_26423);
nand U26737 (N_26737,N_26430,N_26537);
nand U26738 (N_26738,N_26521,N_26461);
nor U26739 (N_26739,N_26424,N_26500);
and U26740 (N_26740,N_26514,N_26578);
nor U26741 (N_26741,N_26489,N_26464);
and U26742 (N_26742,N_26538,N_26551);
nand U26743 (N_26743,N_26434,N_26487);
or U26744 (N_26744,N_26561,N_26450);
and U26745 (N_26745,N_26417,N_26416);
nor U26746 (N_26746,N_26525,N_26586);
and U26747 (N_26747,N_26547,N_26470);
xor U26748 (N_26748,N_26506,N_26504);
nor U26749 (N_26749,N_26567,N_26578);
xor U26750 (N_26750,N_26558,N_26485);
xor U26751 (N_26751,N_26577,N_26545);
nor U26752 (N_26752,N_26404,N_26510);
xnor U26753 (N_26753,N_26473,N_26511);
and U26754 (N_26754,N_26584,N_26452);
nor U26755 (N_26755,N_26459,N_26493);
and U26756 (N_26756,N_26576,N_26411);
or U26757 (N_26757,N_26407,N_26430);
nor U26758 (N_26758,N_26593,N_26465);
xnor U26759 (N_26759,N_26566,N_26589);
nand U26760 (N_26760,N_26502,N_26401);
and U26761 (N_26761,N_26541,N_26430);
xnor U26762 (N_26762,N_26471,N_26553);
nor U26763 (N_26763,N_26418,N_26574);
and U26764 (N_26764,N_26560,N_26529);
or U26765 (N_26765,N_26547,N_26583);
xnor U26766 (N_26766,N_26426,N_26457);
xor U26767 (N_26767,N_26459,N_26449);
nand U26768 (N_26768,N_26404,N_26502);
and U26769 (N_26769,N_26549,N_26421);
xor U26770 (N_26770,N_26430,N_26493);
xnor U26771 (N_26771,N_26497,N_26415);
nor U26772 (N_26772,N_26438,N_26536);
nor U26773 (N_26773,N_26488,N_26421);
or U26774 (N_26774,N_26416,N_26478);
nand U26775 (N_26775,N_26454,N_26488);
nand U26776 (N_26776,N_26403,N_26495);
and U26777 (N_26777,N_26451,N_26402);
xor U26778 (N_26778,N_26435,N_26481);
nor U26779 (N_26779,N_26464,N_26497);
or U26780 (N_26780,N_26421,N_26492);
and U26781 (N_26781,N_26582,N_26467);
and U26782 (N_26782,N_26545,N_26569);
nand U26783 (N_26783,N_26594,N_26492);
xnor U26784 (N_26784,N_26485,N_26505);
nand U26785 (N_26785,N_26452,N_26503);
nand U26786 (N_26786,N_26572,N_26489);
nand U26787 (N_26787,N_26501,N_26409);
nor U26788 (N_26788,N_26451,N_26436);
nand U26789 (N_26789,N_26446,N_26434);
and U26790 (N_26790,N_26528,N_26406);
or U26791 (N_26791,N_26537,N_26575);
or U26792 (N_26792,N_26564,N_26550);
and U26793 (N_26793,N_26411,N_26589);
nor U26794 (N_26794,N_26560,N_26454);
xor U26795 (N_26795,N_26465,N_26598);
and U26796 (N_26796,N_26542,N_26505);
xnor U26797 (N_26797,N_26452,N_26587);
nor U26798 (N_26798,N_26427,N_26588);
and U26799 (N_26799,N_26488,N_26491);
nor U26800 (N_26800,N_26651,N_26624);
and U26801 (N_26801,N_26649,N_26614);
nor U26802 (N_26802,N_26701,N_26702);
nand U26803 (N_26803,N_26683,N_26632);
and U26804 (N_26804,N_26663,N_26754);
xnor U26805 (N_26805,N_26640,N_26694);
and U26806 (N_26806,N_26669,N_26719);
or U26807 (N_26807,N_26672,N_26771);
nand U26808 (N_26808,N_26689,N_26773);
or U26809 (N_26809,N_26781,N_26787);
nand U26810 (N_26810,N_26637,N_26610);
or U26811 (N_26811,N_26648,N_26668);
nand U26812 (N_26812,N_26767,N_26627);
and U26813 (N_26813,N_26710,N_26794);
xor U26814 (N_26814,N_26607,N_26774);
xnor U26815 (N_26815,N_26739,N_26655);
nand U26816 (N_26816,N_26602,N_26709);
nor U26817 (N_26817,N_26733,N_26633);
nor U26818 (N_26818,N_26641,N_26662);
nor U26819 (N_26819,N_26639,N_26714);
nor U26820 (N_26820,N_26691,N_26616);
nand U26821 (N_26821,N_26617,N_26612);
nor U26822 (N_26822,N_26705,N_26777);
xor U26823 (N_26823,N_26670,N_26775);
nor U26824 (N_26824,N_26722,N_26644);
nor U26825 (N_26825,N_26763,N_26686);
xnor U26826 (N_26826,N_26665,N_26798);
or U26827 (N_26827,N_26647,N_26625);
or U26828 (N_26828,N_26724,N_26780);
xnor U26829 (N_26829,N_26772,N_26606);
nor U26830 (N_26830,N_26785,N_26711);
or U26831 (N_26831,N_26677,N_26789);
xnor U26832 (N_26832,N_26721,N_26764);
nor U26833 (N_26833,N_26784,N_26603);
or U26834 (N_26834,N_26712,N_26769);
or U26835 (N_26835,N_26635,N_26736);
xnor U26836 (N_26836,N_26759,N_26729);
nand U26837 (N_26837,N_26782,N_26797);
nand U26838 (N_26838,N_26783,N_26690);
nor U26839 (N_26839,N_26786,N_26636);
or U26840 (N_26840,N_26611,N_26750);
and U26841 (N_26841,N_26730,N_26756);
xnor U26842 (N_26842,N_26629,N_26758);
or U26843 (N_26843,N_26718,N_26643);
nand U26844 (N_26844,N_26695,N_26715);
nor U26845 (N_26845,N_26747,N_26744);
nand U26846 (N_26846,N_26792,N_26790);
or U26847 (N_26847,N_26652,N_26713);
xnor U26848 (N_26848,N_26613,N_26755);
xnor U26849 (N_26849,N_26791,N_26731);
and U26850 (N_26850,N_26734,N_26760);
nor U26851 (N_26851,N_26628,N_26742);
and U26852 (N_26852,N_26723,N_26660);
or U26853 (N_26853,N_26799,N_26765);
and U26854 (N_26854,N_26762,N_26673);
and U26855 (N_26855,N_26745,N_26717);
or U26856 (N_26856,N_26678,N_26605);
nor U26857 (N_26857,N_26658,N_26688);
xor U26858 (N_26858,N_26738,N_26676);
nor U26859 (N_26859,N_26681,N_26674);
nor U26860 (N_26860,N_26726,N_26638);
and U26861 (N_26861,N_26685,N_26650);
or U26862 (N_26862,N_26703,N_26666);
nand U26863 (N_26863,N_26630,N_26679);
and U26864 (N_26864,N_26761,N_26740);
xnor U26865 (N_26865,N_26748,N_26601);
nor U26866 (N_26866,N_26646,N_26698);
xnor U26867 (N_26867,N_26659,N_26743);
or U26868 (N_26868,N_26779,N_26661);
nor U26869 (N_26869,N_26687,N_26727);
and U26870 (N_26870,N_26631,N_26621);
and U26871 (N_26871,N_26716,N_26693);
and U26872 (N_26872,N_26675,N_26704);
xor U26873 (N_26873,N_26620,N_26696);
and U26874 (N_26874,N_26657,N_26671);
or U26875 (N_26875,N_26776,N_26707);
nor U26876 (N_26876,N_26664,N_26692);
or U26877 (N_26877,N_26735,N_26757);
nor U26878 (N_26878,N_26622,N_26645);
nor U26879 (N_26879,N_26770,N_26766);
xor U26880 (N_26880,N_26623,N_26795);
nor U26881 (N_26881,N_26752,N_26682);
or U26882 (N_26882,N_26609,N_26725);
and U26883 (N_26883,N_26749,N_26699);
nor U26884 (N_26884,N_26619,N_26728);
nor U26885 (N_26885,N_26654,N_26796);
and U26886 (N_26886,N_26788,N_26751);
nand U26887 (N_26887,N_26768,N_26737);
nand U26888 (N_26888,N_26746,N_26604);
nor U26889 (N_26889,N_26708,N_26753);
and U26890 (N_26890,N_26667,N_26720);
and U26891 (N_26891,N_26741,N_26626);
and U26892 (N_26892,N_26706,N_26793);
nand U26893 (N_26893,N_26778,N_26684);
and U26894 (N_26894,N_26700,N_26680);
xnor U26895 (N_26895,N_26600,N_26697);
and U26896 (N_26896,N_26608,N_26634);
and U26897 (N_26897,N_26653,N_26656);
xnor U26898 (N_26898,N_26615,N_26642);
and U26899 (N_26899,N_26618,N_26732);
and U26900 (N_26900,N_26774,N_26615);
or U26901 (N_26901,N_26669,N_26624);
and U26902 (N_26902,N_26629,N_26749);
or U26903 (N_26903,N_26678,N_26611);
nor U26904 (N_26904,N_26759,N_26779);
and U26905 (N_26905,N_26645,N_26763);
nand U26906 (N_26906,N_26744,N_26685);
xnor U26907 (N_26907,N_26718,N_26706);
and U26908 (N_26908,N_26775,N_26687);
nor U26909 (N_26909,N_26721,N_26669);
or U26910 (N_26910,N_26643,N_26621);
xnor U26911 (N_26911,N_26778,N_26640);
xnor U26912 (N_26912,N_26714,N_26763);
nand U26913 (N_26913,N_26624,N_26723);
nand U26914 (N_26914,N_26691,N_26666);
and U26915 (N_26915,N_26666,N_26793);
nand U26916 (N_26916,N_26666,N_26692);
nand U26917 (N_26917,N_26710,N_26635);
nor U26918 (N_26918,N_26799,N_26629);
xnor U26919 (N_26919,N_26780,N_26773);
xor U26920 (N_26920,N_26746,N_26608);
and U26921 (N_26921,N_26746,N_26744);
xor U26922 (N_26922,N_26718,N_26683);
nor U26923 (N_26923,N_26681,N_26634);
nand U26924 (N_26924,N_26744,N_26668);
xor U26925 (N_26925,N_26695,N_26796);
xor U26926 (N_26926,N_26669,N_26605);
nand U26927 (N_26927,N_26695,N_26601);
and U26928 (N_26928,N_26663,N_26752);
xor U26929 (N_26929,N_26751,N_26617);
nand U26930 (N_26930,N_26666,N_26632);
or U26931 (N_26931,N_26636,N_26655);
and U26932 (N_26932,N_26701,N_26696);
nand U26933 (N_26933,N_26794,N_26648);
nor U26934 (N_26934,N_26654,N_26683);
or U26935 (N_26935,N_26606,N_26631);
xor U26936 (N_26936,N_26667,N_26709);
xor U26937 (N_26937,N_26767,N_26670);
or U26938 (N_26938,N_26612,N_26684);
or U26939 (N_26939,N_26746,N_26779);
nor U26940 (N_26940,N_26743,N_26650);
xor U26941 (N_26941,N_26650,N_26642);
and U26942 (N_26942,N_26727,N_26638);
or U26943 (N_26943,N_26769,N_26633);
nand U26944 (N_26944,N_26639,N_26614);
nor U26945 (N_26945,N_26611,N_26789);
xnor U26946 (N_26946,N_26748,N_26766);
and U26947 (N_26947,N_26784,N_26610);
xnor U26948 (N_26948,N_26699,N_26700);
nand U26949 (N_26949,N_26650,N_26665);
and U26950 (N_26950,N_26725,N_26738);
xnor U26951 (N_26951,N_26656,N_26794);
nor U26952 (N_26952,N_26792,N_26682);
nor U26953 (N_26953,N_26673,N_26654);
and U26954 (N_26954,N_26787,N_26665);
nor U26955 (N_26955,N_26730,N_26608);
xor U26956 (N_26956,N_26769,N_26679);
or U26957 (N_26957,N_26656,N_26720);
xnor U26958 (N_26958,N_26600,N_26658);
nand U26959 (N_26959,N_26638,N_26737);
nor U26960 (N_26960,N_26609,N_26786);
or U26961 (N_26961,N_26785,N_26635);
nor U26962 (N_26962,N_26622,N_26749);
or U26963 (N_26963,N_26693,N_26791);
nor U26964 (N_26964,N_26620,N_26669);
nand U26965 (N_26965,N_26622,N_26638);
nor U26966 (N_26966,N_26797,N_26692);
and U26967 (N_26967,N_26687,N_26669);
xnor U26968 (N_26968,N_26700,N_26753);
or U26969 (N_26969,N_26713,N_26788);
nand U26970 (N_26970,N_26613,N_26747);
nand U26971 (N_26971,N_26636,N_26796);
nand U26972 (N_26972,N_26661,N_26680);
and U26973 (N_26973,N_26720,N_26663);
or U26974 (N_26974,N_26678,N_26739);
and U26975 (N_26975,N_26614,N_26659);
and U26976 (N_26976,N_26795,N_26655);
xnor U26977 (N_26977,N_26677,N_26778);
nor U26978 (N_26978,N_26632,N_26771);
nand U26979 (N_26979,N_26750,N_26796);
xor U26980 (N_26980,N_26766,N_26712);
and U26981 (N_26981,N_26649,N_26650);
xor U26982 (N_26982,N_26640,N_26615);
and U26983 (N_26983,N_26649,N_26745);
nor U26984 (N_26984,N_26702,N_26695);
or U26985 (N_26985,N_26775,N_26777);
or U26986 (N_26986,N_26608,N_26762);
and U26987 (N_26987,N_26731,N_26793);
nor U26988 (N_26988,N_26684,N_26605);
or U26989 (N_26989,N_26681,N_26640);
and U26990 (N_26990,N_26757,N_26773);
or U26991 (N_26991,N_26782,N_26631);
xnor U26992 (N_26992,N_26711,N_26660);
nor U26993 (N_26993,N_26786,N_26606);
nor U26994 (N_26994,N_26721,N_26742);
and U26995 (N_26995,N_26690,N_26776);
nor U26996 (N_26996,N_26636,N_26712);
and U26997 (N_26997,N_26627,N_26635);
and U26998 (N_26998,N_26722,N_26733);
nor U26999 (N_26999,N_26679,N_26699);
nor U27000 (N_27000,N_26991,N_26888);
or U27001 (N_27001,N_26857,N_26975);
xor U27002 (N_27002,N_26887,N_26870);
nor U27003 (N_27003,N_26818,N_26950);
xnor U27004 (N_27004,N_26886,N_26881);
or U27005 (N_27005,N_26873,N_26931);
and U27006 (N_27006,N_26845,N_26929);
or U27007 (N_27007,N_26942,N_26851);
nand U27008 (N_27008,N_26913,N_26976);
xnor U27009 (N_27009,N_26856,N_26841);
xor U27010 (N_27010,N_26892,N_26863);
nor U27011 (N_27011,N_26923,N_26930);
nand U27012 (N_27012,N_26821,N_26938);
nand U27013 (N_27013,N_26829,N_26914);
nor U27014 (N_27014,N_26868,N_26898);
and U27015 (N_27015,N_26884,N_26831);
xor U27016 (N_27016,N_26895,N_26911);
or U27017 (N_27017,N_26838,N_26830);
nor U27018 (N_27018,N_26853,N_26947);
xnor U27019 (N_27019,N_26973,N_26939);
nor U27020 (N_27020,N_26960,N_26935);
xor U27021 (N_27021,N_26859,N_26817);
or U27022 (N_27022,N_26977,N_26835);
xnor U27023 (N_27023,N_26910,N_26943);
nor U27024 (N_27024,N_26912,N_26849);
xnor U27025 (N_27025,N_26815,N_26917);
and U27026 (N_27026,N_26876,N_26906);
and U27027 (N_27027,N_26963,N_26860);
nor U27028 (N_27028,N_26806,N_26986);
nor U27029 (N_27029,N_26985,N_26993);
and U27030 (N_27030,N_26984,N_26901);
and U27031 (N_27031,N_26826,N_26812);
and U27032 (N_27032,N_26918,N_26957);
nor U27033 (N_27033,N_26941,N_26944);
nand U27034 (N_27034,N_26832,N_26896);
or U27035 (N_27035,N_26840,N_26869);
nor U27036 (N_27036,N_26996,N_26897);
nor U27037 (N_27037,N_26894,N_26937);
or U27038 (N_27038,N_26925,N_26965);
xnor U27039 (N_27039,N_26948,N_26858);
nor U27040 (N_27040,N_26839,N_26825);
xor U27041 (N_27041,N_26934,N_26919);
xnor U27042 (N_27042,N_26862,N_26811);
nand U27043 (N_27043,N_26922,N_26899);
nand U27044 (N_27044,N_26964,N_26819);
xnor U27045 (N_27045,N_26834,N_26978);
nor U27046 (N_27046,N_26933,N_26878);
and U27047 (N_27047,N_26828,N_26883);
and U27048 (N_27048,N_26967,N_26992);
nand U27049 (N_27049,N_26864,N_26970);
and U27050 (N_27050,N_26969,N_26836);
or U27051 (N_27051,N_26983,N_26842);
or U27052 (N_27052,N_26871,N_26879);
and U27053 (N_27053,N_26974,N_26877);
xor U27054 (N_27054,N_26875,N_26885);
xor U27055 (N_27055,N_26997,N_26833);
nor U27056 (N_27056,N_26916,N_26808);
xnor U27057 (N_27057,N_26909,N_26874);
nand U27058 (N_27058,N_26903,N_26924);
and U27059 (N_27059,N_26915,N_26861);
nand U27060 (N_27060,N_26890,N_26952);
nand U27061 (N_27061,N_26837,N_26981);
and U27062 (N_27062,N_26972,N_26907);
and U27063 (N_27063,N_26900,N_26848);
and U27064 (N_27064,N_26971,N_26814);
nand U27065 (N_27065,N_26928,N_26953);
nand U27066 (N_27066,N_26823,N_26946);
nand U27067 (N_27067,N_26982,N_26801);
xnor U27068 (N_27068,N_26905,N_26921);
or U27069 (N_27069,N_26940,N_26802);
nand U27070 (N_27070,N_26805,N_26882);
xnor U27071 (N_27071,N_26813,N_26908);
xor U27072 (N_27072,N_26920,N_26803);
nor U27073 (N_27073,N_26980,N_26804);
or U27074 (N_27074,N_26961,N_26847);
nor U27075 (N_27075,N_26956,N_26987);
and U27076 (N_27076,N_26959,N_26807);
and U27077 (N_27077,N_26958,N_26865);
or U27078 (N_27078,N_26990,N_26880);
nor U27079 (N_27079,N_26904,N_26867);
nand U27080 (N_27080,N_26945,N_26800);
nor U27081 (N_27081,N_26810,N_26843);
xor U27082 (N_27082,N_26998,N_26816);
xnor U27083 (N_27083,N_26893,N_26824);
and U27084 (N_27084,N_26932,N_26926);
xnor U27085 (N_27085,N_26822,N_26995);
or U27086 (N_27086,N_26949,N_26820);
nand U27087 (N_27087,N_26988,N_26966);
nand U27088 (N_27088,N_26844,N_26855);
nor U27089 (N_27089,N_26854,N_26809);
nor U27090 (N_27090,N_26955,N_26872);
nor U27091 (N_27091,N_26979,N_26902);
and U27092 (N_27092,N_26866,N_26994);
nand U27093 (N_27093,N_26989,N_26936);
or U27094 (N_27094,N_26852,N_26968);
nor U27095 (N_27095,N_26927,N_26846);
xnor U27096 (N_27096,N_26850,N_26951);
or U27097 (N_27097,N_26827,N_26999);
nand U27098 (N_27098,N_26962,N_26954);
xor U27099 (N_27099,N_26891,N_26889);
nand U27100 (N_27100,N_26812,N_26824);
nor U27101 (N_27101,N_26909,N_26948);
and U27102 (N_27102,N_26810,N_26947);
and U27103 (N_27103,N_26893,N_26960);
nor U27104 (N_27104,N_26903,N_26871);
or U27105 (N_27105,N_26947,N_26975);
or U27106 (N_27106,N_26900,N_26835);
and U27107 (N_27107,N_26905,N_26879);
xnor U27108 (N_27108,N_26828,N_26882);
nand U27109 (N_27109,N_26855,N_26912);
nand U27110 (N_27110,N_26968,N_26844);
xnor U27111 (N_27111,N_26821,N_26888);
nor U27112 (N_27112,N_26990,N_26995);
or U27113 (N_27113,N_26978,N_26938);
nand U27114 (N_27114,N_26918,N_26942);
and U27115 (N_27115,N_26994,N_26913);
xor U27116 (N_27116,N_26984,N_26912);
nand U27117 (N_27117,N_26974,N_26946);
nor U27118 (N_27118,N_26965,N_26848);
nor U27119 (N_27119,N_26936,N_26910);
nand U27120 (N_27120,N_26903,N_26846);
xor U27121 (N_27121,N_26863,N_26951);
xor U27122 (N_27122,N_26932,N_26968);
nor U27123 (N_27123,N_26853,N_26963);
xnor U27124 (N_27124,N_26901,N_26851);
nand U27125 (N_27125,N_26940,N_26938);
nand U27126 (N_27126,N_26882,N_26984);
nand U27127 (N_27127,N_26958,N_26903);
nand U27128 (N_27128,N_26872,N_26983);
nor U27129 (N_27129,N_26913,N_26811);
or U27130 (N_27130,N_26866,N_26949);
nand U27131 (N_27131,N_26845,N_26962);
nor U27132 (N_27132,N_26829,N_26983);
nand U27133 (N_27133,N_26899,N_26938);
and U27134 (N_27134,N_26886,N_26898);
and U27135 (N_27135,N_26807,N_26947);
and U27136 (N_27136,N_26921,N_26962);
nand U27137 (N_27137,N_26959,N_26896);
or U27138 (N_27138,N_26802,N_26930);
nor U27139 (N_27139,N_26922,N_26860);
or U27140 (N_27140,N_26947,N_26954);
nand U27141 (N_27141,N_26844,N_26806);
nand U27142 (N_27142,N_26845,N_26939);
or U27143 (N_27143,N_26993,N_26894);
nor U27144 (N_27144,N_26806,N_26905);
nor U27145 (N_27145,N_26984,N_26823);
and U27146 (N_27146,N_26833,N_26801);
nor U27147 (N_27147,N_26991,N_26963);
xnor U27148 (N_27148,N_26893,N_26919);
or U27149 (N_27149,N_26925,N_26883);
nand U27150 (N_27150,N_26865,N_26864);
and U27151 (N_27151,N_26966,N_26812);
or U27152 (N_27152,N_26834,N_26916);
nor U27153 (N_27153,N_26933,N_26867);
nand U27154 (N_27154,N_26978,N_26846);
nor U27155 (N_27155,N_26894,N_26871);
nand U27156 (N_27156,N_26871,N_26816);
and U27157 (N_27157,N_26995,N_26825);
nand U27158 (N_27158,N_26919,N_26818);
and U27159 (N_27159,N_26946,N_26864);
nand U27160 (N_27160,N_26962,N_26893);
xnor U27161 (N_27161,N_26887,N_26885);
and U27162 (N_27162,N_26953,N_26948);
or U27163 (N_27163,N_26900,N_26926);
and U27164 (N_27164,N_26894,N_26900);
nand U27165 (N_27165,N_26905,N_26814);
and U27166 (N_27166,N_26975,N_26803);
nor U27167 (N_27167,N_26929,N_26861);
or U27168 (N_27168,N_26809,N_26966);
nor U27169 (N_27169,N_26826,N_26913);
and U27170 (N_27170,N_26833,N_26980);
nand U27171 (N_27171,N_26855,N_26895);
nor U27172 (N_27172,N_26932,N_26910);
nor U27173 (N_27173,N_26949,N_26897);
nor U27174 (N_27174,N_26856,N_26937);
nor U27175 (N_27175,N_26896,N_26901);
xor U27176 (N_27176,N_26808,N_26809);
or U27177 (N_27177,N_26963,N_26946);
and U27178 (N_27178,N_26952,N_26928);
or U27179 (N_27179,N_26816,N_26859);
nor U27180 (N_27180,N_26866,N_26943);
xor U27181 (N_27181,N_26987,N_26908);
and U27182 (N_27182,N_26982,N_26986);
and U27183 (N_27183,N_26964,N_26804);
xor U27184 (N_27184,N_26917,N_26982);
and U27185 (N_27185,N_26836,N_26989);
nand U27186 (N_27186,N_26998,N_26901);
nand U27187 (N_27187,N_26834,N_26995);
or U27188 (N_27188,N_26945,N_26920);
nor U27189 (N_27189,N_26801,N_26973);
or U27190 (N_27190,N_26934,N_26994);
or U27191 (N_27191,N_26888,N_26994);
xor U27192 (N_27192,N_26830,N_26828);
nand U27193 (N_27193,N_26838,N_26987);
or U27194 (N_27194,N_26817,N_26946);
nand U27195 (N_27195,N_26873,N_26810);
nand U27196 (N_27196,N_26894,N_26969);
xor U27197 (N_27197,N_26988,N_26918);
or U27198 (N_27198,N_26902,N_26945);
nor U27199 (N_27199,N_26810,N_26837);
nand U27200 (N_27200,N_27194,N_27132);
or U27201 (N_27201,N_27147,N_27026);
or U27202 (N_27202,N_27167,N_27109);
and U27203 (N_27203,N_27172,N_27096);
or U27204 (N_27204,N_27074,N_27037);
or U27205 (N_27205,N_27168,N_27193);
nor U27206 (N_27206,N_27104,N_27134);
and U27207 (N_27207,N_27185,N_27116);
or U27208 (N_27208,N_27153,N_27094);
nand U27209 (N_27209,N_27117,N_27012);
or U27210 (N_27210,N_27097,N_27158);
or U27211 (N_27211,N_27051,N_27061);
nand U27212 (N_27212,N_27098,N_27190);
or U27213 (N_27213,N_27019,N_27161);
nor U27214 (N_27214,N_27048,N_27013);
and U27215 (N_27215,N_27059,N_27038);
nor U27216 (N_27216,N_27092,N_27049);
nor U27217 (N_27217,N_27126,N_27191);
and U27218 (N_27218,N_27197,N_27075);
xnor U27219 (N_27219,N_27040,N_27196);
xnor U27220 (N_27220,N_27103,N_27064);
nor U27221 (N_27221,N_27009,N_27159);
nand U27222 (N_27222,N_27175,N_27043);
and U27223 (N_27223,N_27138,N_27127);
and U27224 (N_27224,N_27189,N_27160);
or U27225 (N_27225,N_27001,N_27078);
and U27226 (N_27226,N_27028,N_27107);
and U27227 (N_27227,N_27198,N_27021);
xnor U27228 (N_27228,N_27195,N_27140);
xor U27229 (N_27229,N_27030,N_27093);
nand U27230 (N_27230,N_27118,N_27120);
nand U27231 (N_27231,N_27004,N_27016);
nor U27232 (N_27232,N_27182,N_27099);
and U27233 (N_27233,N_27010,N_27129);
nor U27234 (N_27234,N_27068,N_27020);
or U27235 (N_27235,N_27035,N_27079);
or U27236 (N_27236,N_27188,N_27174);
or U27237 (N_27237,N_27192,N_27003);
nor U27238 (N_27238,N_27089,N_27027);
xor U27239 (N_27239,N_27178,N_27151);
nor U27240 (N_27240,N_27053,N_27155);
and U27241 (N_27241,N_27014,N_27162);
xor U27242 (N_27242,N_27083,N_27146);
or U27243 (N_27243,N_27110,N_27022);
nor U27244 (N_27244,N_27055,N_27101);
and U27245 (N_27245,N_27137,N_27177);
or U27246 (N_27246,N_27112,N_27154);
and U27247 (N_27247,N_27057,N_27071);
or U27248 (N_27248,N_27102,N_27045);
or U27249 (N_27249,N_27006,N_27100);
or U27250 (N_27250,N_27067,N_27018);
and U27251 (N_27251,N_27062,N_27113);
or U27252 (N_27252,N_27157,N_27011);
nor U27253 (N_27253,N_27046,N_27184);
xor U27254 (N_27254,N_27169,N_27091);
and U27255 (N_27255,N_27166,N_27056);
and U27256 (N_27256,N_27150,N_27077);
xnor U27257 (N_27257,N_27032,N_27039);
nor U27258 (N_27258,N_27058,N_27052);
nand U27259 (N_27259,N_27123,N_27187);
xnor U27260 (N_27260,N_27063,N_27133);
or U27261 (N_27261,N_27119,N_27042);
and U27262 (N_27262,N_27080,N_27076);
and U27263 (N_27263,N_27017,N_27148);
and U27264 (N_27264,N_27007,N_27199);
xnor U27265 (N_27265,N_27125,N_27165);
xor U27266 (N_27266,N_27144,N_27087);
or U27267 (N_27267,N_27029,N_27085);
and U27268 (N_27268,N_27170,N_27008);
xnor U27269 (N_27269,N_27044,N_27005);
xnor U27270 (N_27270,N_27176,N_27124);
and U27271 (N_27271,N_27082,N_27141);
xor U27272 (N_27272,N_27115,N_27108);
xor U27273 (N_27273,N_27086,N_27084);
nor U27274 (N_27274,N_27130,N_27163);
or U27275 (N_27275,N_27180,N_27066);
nor U27276 (N_27276,N_27073,N_27041);
nor U27277 (N_27277,N_27072,N_27156);
xnor U27278 (N_27278,N_27186,N_27023);
nand U27279 (N_27279,N_27033,N_27069);
or U27280 (N_27280,N_27143,N_27131);
nand U27281 (N_27281,N_27114,N_27065);
nor U27282 (N_27282,N_27149,N_27135);
or U27283 (N_27283,N_27152,N_27060);
xor U27284 (N_27284,N_27171,N_27164);
xor U27285 (N_27285,N_27090,N_27036);
and U27286 (N_27286,N_27081,N_27050);
nor U27287 (N_27287,N_27122,N_27139);
and U27288 (N_27288,N_27002,N_27088);
and U27289 (N_27289,N_27034,N_27136);
and U27290 (N_27290,N_27111,N_27095);
and U27291 (N_27291,N_27105,N_27145);
xnor U27292 (N_27292,N_27024,N_27070);
nand U27293 (N_27293,N_27025,N_27015);
nand U27294 (N_27294,N_27181,N_27183);
and U27295 (N_27295,N_27179,N_27121);
or U27296 (N_27296,N_27142,N_27000);
and U27297 (N_27297,N_27054,N_27031);
and U27298 (N_27298,N_27173,N_27047);
nand U27299 (N_27299,N_27128,N_27106);
or U27300 (N_27300,N_27190,N_27083);
nor U27301 (N_27301,N_27156,N_27151);
xnor U27302 (N_27302,N_27147,N_27169);
and U27303 (N_27303,N_27066,N_27183);
nand U27304 (N_27304,N_27133,N_27011);
xnor U27305 (N_27305,N_27108,N_27033);
and U27306 (N_27306,N_27024,N_27148);
or U27307 (N_27307,N_27172,N_27135);
nor U27308 (N_27308,N_27184,N_27047);
nand U27309 (N_27309,N_27020,N_27177);
or U27310 (N_27310,N_27134,N_27024);
nand U27311 (N_27311,N_27175,N_27079);
or U27312 (N_27312,N_27111,N_27197);
xor U27313 (N_27313,N_27185,N_27001);
or U27314 (N_27314,N_27084,N_27164);
nand U27315 (N_27315,N_27157,N_27070);
nor U27316 (N_27316,N_27123,N_27061);
nand U27317 (N_27317,N_27166,N_27150);
or U27318 (N_27318,N_27030,N_27004);
and U27319 (N_27319,N_27118,N_27102);
and U27320 (N_27320,N_27004,N_27044);
or U27321 (N_27321,N_27174,N_27149);
or U27322 (N_27322,N_27137,N_27108);
or U27323 (N_27323,N_27136,N_27166);
or U27324 (N_27324,N_27160,N_27143);
nor U27325 (N_27325,N_27193,N_27183);
or U27326 (N_27326,N_27149,N_27008);
xnor U27327 (N_27327,N_27148,N_27042);
or U27328 (N_27328,N_27075,N_27025);
xnor U27329 (N_27329,N_27024,N_27170);
and U27330 (N_27330,N_27190,N_27032);
nor U27331 (N_27331,N_27135,N_27099);
or U27332 (N_27332,N_27051,N_27108);
and U27333 (N_27333,N_27129,N_27164);
or U27334 (N_27334,N_27118,N_27009);
nand U27335 (N_27335,N_27147,N_27136);
nand U27336 (N_27336,N_27084,N_27149);
and U27337 (N_27337,N_27071,N_27020);
nand U27338 (N_27338,N_27159,N_27158);
and U27339 (N_27339,N_27190,N_27059);
nor U27340 (N_27340,N_27070,N_27182);
xnor U27341 (N_27341,N_27178,N_27165);
and U27342 (N_27342,N_27199,N_27142);
nor U27343 (N_27343,N_27067,N_27121);
nor U27344 (N_27344,N_27031,N_27178);
nand U27345 (N_27345,N_27114,N_27136);
nand U27346 (N_27346,N_27009,N_27005);
or U27347 (N_27347,N_27197,N_27060);
xor U27348 (N_27348,N_27165,N_27025);
and U27349 (N_27349,N_27109,N_27036);
or U27350 (N_27350,N_27171,N_27190);
and U27351 (N_27351,N_27142,N_27036);
or U27352 (N_27352,N_27020,N_27166);
xor U27353 (N_27353,N_27160,N_27186);
and U27354 (N_27354,N_27069,N_27024);
nor U27355 (N_27355,N_27038,N_27091);
nor U27356 (N_27356,N_27114,N_27008);
or U27357 (N_27357,N_27122,N_27178);
nand U27358 (N_27358,N_27115,N_27048);
nand U27359 (N_27359,N_27061,N_27021);
or U27360 (N_27360,N_27063,N_27058);
or U27361 (N_27361,N_27046,N_27070);
and U27362 (N_27362,N_27107,N_27066);
nand U27363 (N_27363,N_27052,N_27181);
xor U27364 (N_27364,N_27105,N_27068);
or U27365 (N_27365,N_27136,N_27048);
or U27366 (N_27366,N_27125,N_27198);
nor U27367 (N_27367,N_27182,N_27041);
nor U27368 (N_27368,N_27088,N_27139);
xnor U27369 (N_27369,N_27060,N_27193);
or U27370 (N_27370,N_27021,N_27032);
nand U27371 (N_27371,N_27162,N_27116);
nand U27372 (N_27372,N_27030,N_27089);
and U27373 (N_27373,N_27181,N_27197);
xnor U27374 (N_27374,N_27006,N_27000);
or U27375 (N_27375,N_27132,N_27113);
or U27376 (N_27376,N_27025,N_27009);
xor U27377 (N_27377,N_27015,N_27189);
and U27378 (N_27378,N_27071,N_27151);
and U27379 (N_27379,N_27066,N_27195);
xor U27380 (N_27380,N_27197,N_27007);
and U27381 (N_27381,N_27085,N_27147);
xnor U27382 (N_27382,N_27100,N_27113);
or U27383 (N_27383,N_27094,N_27174);
nand U27384 (N_27384,N_27177,N_27035);
xor U27385 (N_27385,N_27065,N_27174);
and U27386 (N_27386,N_27038,N_27153);
nand U27387 (N_27387,N_27197,N_27003);
or U27388 (N_27388,N_27082,N_27006);
or U27389 (N_27389,N_27029,N_27138);
and U27390 (N_27390,N_27036,N_27122);
and U27391 (N_27391,N_27175,N_27061);
nor U27392 (N_27392,N_27037,N_27115);
and U27393 (N_27393,N_27011,N_27111);
nand U27394 (N_27394,N_27044,N_27197);
or U27395 (N_27395,N_27162,N_27022);
nand U27396 (N_27396,N_27113,N_27144);
nand U27397 (N_27397,N_27034,N_27169);
and U27398 (N_27398,N_27103,N_27144);
xor U27399 (N_27399,N_27137,N_27169);
nor U27400 (N_27400,N_27316,N_27200);
nor U27401 (N_27401,N_27389,N_27398);
xor U27402 (N_27402,N_27352,N_27257);
and U27403 (N_27403,N_27268,N_27294);
xor U27404 (N_27404,N_27302,N_27350);
nand U27405 (N_27405,N_27299,N_27386);
or U27406 (N_27406,N_27369,N_27228);
nor U27407 (N_27407,N_27303,N_27295);
or U27408 (N_27408,N_27203,N_27229);
nor U27409 (N_27409,N_27277,N_27355);
and U27410 (N_27410,N_27337,N_27298);
nor U27411 (N_27411,N_27358,N_27248);
nor U27412 (N_27412,N_27212,N_27368);
and U27413 (N_27413,N_27318,N_27222);
and U27414 (N_27414,N_27395,N_27282);
or U27415 (N_27415,N_27237,N_27312);
and U27416 (N_27416,N_27380,N_27283);
or U27417 (N_27417,N_27366,N_27309);
or U27418 (N_27418,N_27367,N_27278);
nand U27419 (N_27419,N_27258,N_27216);
nand U27420 (N_27420,N_27327,N_27361);
nand U27421 (N_27421,N_27250,N_27347);
and U27422 (N_27422,N_27285,N_27365);
and U27423 (N_27423,N_27322,N_27315);
or U27424 (N_27424,N_27245,N_27232);
xor U27425 (N_27425,N_27383,N_27332);
xnor U27426 (N_27426,N_27213,N_27307);
and U27427 (N_27427,N_27391,N_27382);
or U27428 (N_27428,N_27210,N_27267);
nor U27429 (N_27429,N_27390,N_27218);
nand U27430 (N_27430,N_27255,N_27331);
xor U27431 (N_27431,N_27351,N_27215);
nand U27432 (N_27432,N_27291,N_27239);
or U27433 (N_27433,N_27304,N_27279);
nor U27434 (N_27434,N_27234,N_27362);
nand U27435 (N_27435,N_27266,N_27354);
and U27436 (N_27436,N_27231,N_27345);
and U27437 (N_27437,N_27290,N_27253);
nor U27438 (N_27438,N_27370,N_27204);
nand U27439 (N_27439,N_27264,N_27296);
or U27440 (N_27440,N_27224,N_27297);
xnor U27441 (N_27441,N_27392,N_27385);
and U27442 (N_27442,N_27305,N_27306);
or U27443 (N_27443,N_27293,N_27396);
or U27444 (N_27444,N_27348,N_27270);
xnor U27445 (N_27445,N_27372,N_27289);
nor U27446 (N_27446,N_27211,N_27205);
nand U27447 (N_27447,N_27319,N_27397);
or U27448 (N_27448,N_27284,N_27281);
or U27449 (N_27449,N_27321,N_27252);
xor U27450 (N_27450,N_27244,N_27286);
xnor U27451 (N_27451,N_27346,N_27251);
or U27452 (N_27452,N_27311,N_27226);
or U27453 (N_27453,N_27262,N_27220);
or U27454 (N_27454,N_27326,N_27399);
and U27455 (N_27455,N_27353,N_27259);
nor U27456 (N_27456,N_27256,N_27300);
or U27457 (N_27457,N_27217,N_27208);
nor U27458 (N_27458,N_27374,N_27276);
nor U27459 (N_27459,N_27323,N_27376);
nor U27460 (N_27460,N_27330,N_27314);
xnor U27461 (N_27461,N_27263,N_27292);
nor U27462 (N_27462,N_27338,N_27393);
and U27463 (N_27463,N_27359,N_27335);
and U27464 (N_27464,N_27371,N_27377);
nor U27465 (N_27465,N_27333,N_27342);
nand U27466 (N_27466,N_27340,N_27328);
and U27467 (N_27467,N_27388,N_27273);
xnor U27468 (N_27468,N_27339,N_27394);
or U27469 (N_27469,N_27356,N_27223);
or U27470 (N_27470,N_27206,N_27381);
nor U27471 (N_27471,N_27364,N_27357);
xnor U27472 (N_27472,N_27363,N_27238);
nand U27473 (N_27473,N_27301,N_27320);
nand U27474 (N_27474,N_27275,N_27241);
or U27475 (N_27475,N_27201,N_27243);
nand U27476 (N_27476,N_27219,N_27310);
xnor U27477 (N_27477,N_27384,N_27246);
nand U27478 (N_27478,N_27214,N_27269);
xor U27479 (N_27479,N_27341,N_27379);
and U27480 (N_27480,N_27207,N_27387);
nor U27481 (N_27481,N_27236,N_27344);
nand U27482 (N_27482,N_27343,N_27254);
and U27483 (N_27483,N_27274,N_27225);
and U27484 (N_27484,N_27324,N_27227);
or U27485 (N_27485,N_27209,N_27329);
xnor U27486 (N_27486,N_27202,N_27373);
nand U27487 (N_27487,N_27233,N_27325);
xnor U27488 (N_27488,N_27260,N_27240);
nand U27489 (N_27489,N_27221,N_27249);
xnor U27490 (N_27490,N_27247,N_27336);
nor U27491 (N_27491,N_27261,N_27360);
and U27492 (N_27492,N_27334,N_27235);
nand U27493 (N_27493,N_27288,N_27280);
and U27494 (N_27494,N_27271,N_27272);
nand U27495 (N_27495,N_27265,N_27287);
nand U27496 (N_27496,N_27378,N_27313);
nor U27497 (N_27497,N_27230,N_27349);
xnor U27498 (N_27498,N_27375,N_27242);
and U27499 (N_27499,N_27317,N_27308);
xnor U27500 (N_27500,N_27329,N_27380);
nor U27501 (N_27501,N_27261,N_27381);
or U27502 (N_27502,N_27322,N_27238);
and U27503 (N_27503,N_27291,N_27270);
nand U27504 (N_27504,N_27347,N_27261);
nor U27505 (N_27505,N_27331,N_27382);
xnor U27506 (N_27506,N_27327,N_27211);
xor U27507 (N_27507,N_27340,N_27256);
xor U27508 (N_27508,N_27289,N_27232);
or U27509 (N_27509,N_27221,N_27379);
or U27510 (N_27510,N_27212,N_27205);
or U27511 (N_27511,N_27397,N_27230);
or U27512 (N_27512,N_27266,N_27207);
or U27513 (N_27513,N_27299,N_27313);
and U27514 (N_27514,N_27304,N_27321);
or U27515 (N_27515,N_27207,N_27222);
nand U27516 (N_27516,N_27265,N_27377);
nor U27517 (N_27517,N_27327,N_27235);
and U27518 (N_27518,N_27200,N_27370);
nor U27519 (N_27519,N_27336,N_27253);
nor U27520 (N_27520,N_27309,N_27362);
nand U27521 (N_27521,N_27377,N_27356);
and U27522 (N_27522,N_27286,N_27285);
and U27523 (N_27523,N_27328,N_27258);
or U27524 (N_27524,N_27335,N_27309);
nand U27525 (N_27525,N_27355,N_27270);
nor U27526 (N_27526,N_27397,N_27291);
xor U27527 (N_27527,N_27285,N_27310);
or U27528 (N_27528,N_27233,N_27399);
or U27529 (N_27529,N_27269,N_27357);
nor U27530 (N_27530,N_27399,N_27368);
xor U27531 (N_27531,N_27367,N_27379);
nor U27532 (N_27532,N_27287,N_27219);
nor U27533 (N_27533,N_27318,N_27367);
xnor U27534 (N_27534,N_27219,N_27224);
or U27535 (N_27535,N_27253,N_27266);
nand U27536 (N_27536,N_27211,N_27284);
and U27537 (N_27537,N_27291,N_27394);
or U27538 (N_27538,N_27222,N_27286);
nand U27539 (N_27539,N_27335,N_27343);
or U27540 (N_27540,N_27363,N_27265);
nand U27541 (N_27541,N_27350,N_27366);
or U27542 (N_27542,N_27232,N_27260);
nand U27543 (N_27543,N_27242,N_27374);
nor U27544 (N_27544,N_27231,N_27266);
xor U27545 (N_27545,N_27347,N_27291);
and U27546 (N_27546,N_27350,N_27328);
nand U27547 (N_27547,N_27362,N_27357);
nor U27548 (N_27548,N_27233,N_27250);
or U27549 (N_27549,N_27216,N_27249);
and U27550 (N_27550,N_27338,N_27241);
or U27551 (N_27551,N_27358,N_27324);
and U27552 (N_27552,N_27344,N_27357);
xnor U27553 (N_27553,N_27376,N_27216);
nand U27554 (N_27554,N_27313,N_27236);
and U27555 (N_27555,N_27267,N_27348);
nor U27556 (N_27556,N_27282,N_27332);
and U27557 (N_27557,N_27263,N_27334);
nor U27558 (N_27558,N_27234,N_27319);
or U27559 (N_27559,N_27372,N_27231);
nand U27560 (N_27560,N_27385,N_27228);
nor U27561 (N_27561,N_27337,N_27304);
xor U27562 (N_27562,N_27324,N_27377);
or U27563 (N_27563,N_27231,N_27224);
and U27564 (N_27564,N_27335,N_27244);
nand U27565 (N_27565,N_27372,N_27237);
and U27566 (N_27566,N_27255,N_27324);
nor U27567 (N_27567,N_27246,N_27263);
nand U27568 (N_27568,N_27304,N_27306);
xor U27569 (N_27569,N_27264,N_27272);
xnor U27570 (N_27570,N_27343,N_27220);
and U27571 (N_27571,N_27335,N_27289);
nor U27572 (N_27572,N_27267,N_27238);
or U27573 (N_27573,N_27334,N_27343);
and U27574 (N_27574,N_27394,N_27317);
and U27575 (N_27575,N_27256,N_27359);
nand U27576 (N_27576,N_27392,N_27354);
or U27577 (N_27577,N_27359,N_27399);
or U27578 (N_27578,N_27307,N_27329);
nor U27579 (N_27579,N_27208,N_27266);
or U27580 (N_27580,N_27226,N_27319);
nand U27581 (N_27581,N_27381,N_27343);
nor U27582 (N_27582,N_27242,N_27323);
and U27583 (N_27583,N_27334,N_27375);
or U27584 (N_27584,N_27210,N_27380);
nand U27585 (N_27585,N_27371,N_27247);
or U27586 (N_27586,N_27302,N_27353);
or U27587 (N_27587,N_27319,N_27356);
nand U27588 (N_27588,N_27388,N_27218);
and U27589 (N_27589,N_27335,N_27241);
nor U27590 (N_27590,N_27308,N_27242);
xor U27591 (N_27591,N_27346,N_27300);
nand U27592 (N_27592,N_27260,N_27264);
or U27593 (N_27593,N_27343,N_27282);
and U27594 (N_27594,N_27259,N_27227);
nand U27595 (N_27595,N_27291,N_27325);
or U27596 (N_27596,N_27337,N_27270);
or U27597 (N_27597,N_27207,N_27216);
nor U27598 (N_27598,N_27360,N_27284);
or U27599 (N_27599,N_27297,N_27229);
xnor U27600 (N_27600,N_27531,N_27542);
nand U27601 (N_27601,N_27509,N_27544);
nor U27602 (N_27602,N_27422,N_27416);
and U27603 (N_27603,N_27441,N_27584);
or U27604 (N_27604,N_27472,N_27559);
nor U27605 (N_27605,N_27405,N_27456);
nor U27606 (N_27606,N_27511,N_27508);
nor U27607 (N_27607,N_27486,N_27476);
xnor U27608 (N_27608,N_27591,N_27497);
and U27609 (N_27609,N_27575,N_27526);
and U27610 (N_27610,N_27406,N_27403);
nor U27611 (N_27611,N_27500,N_27477);
nor U27612 (N_27612,N_27572,N_27564);
and U27613 (N_27613,N_27555,N_27588);
nor U27614 (N_27614,N_27549,N_27440);
or U27615 (N_27615,N_27415,N_27465);
and U27616 (N_27616,N_27593,N_27528);
xor U27617 (N_27617,N_27505,N_27453);
nor U27618 (N_27618,N_27499,N_27556);
nand U27619 (N_27619,N_27443,N_27444);
nor U27620 (N_27620,N_27518,N_27451);
xor U27621 (N_27621,N_27567,N_27523);
or U27622 (N_27622,N_27578,N_27562);
nand U27623 (N_27623,N_27570,N_27479);
nand U27624 (N_27624,N_27543,N_27513);
nand U27625 (N_27625,N_27546,N_27548);
and U27626 (N_27626,N_27494,N_27565);
and U27627 (N_27627,N_27534,N_27424);
nor U27628 (N_27628,N_27428,N_27487);
nor U27629 (N_27629,N_27576,N_27557);
nand U27630 (N_27630,N_27492,N_27402);
nor U27631 (N_27631,N_27400,N_27458);
and U27632 (N_27632,N_27495,N_27470);
and U27633 (N_27633,N_27437,N_27480);
and U27634 (N_27634,N_27408,N_27461);
xnor U27635 (N_27635,N_27420,N_27558);
xnor U27636 (N_27636,N_27459,N_27413);
and U27637 (N_27637,N_27407,N_27507);
and U27638 (N_27638,N_27524,N_27447);
xor U27639 (N_27639,N_27580,N_27585);
and U27640 (N_27640,N_27412,N_27550);
xnor U27641 (N_27641,N_27582,N_27488);
or U27642 (N_27642,N_27596,N_27599);
nand U27643 (N_27643,N_27595,N_27404);
and U27644 (N_27644,N_27411,N_27410);
nand U27645 (N_27645,N_27490,N_27538);
nand U27646 (N_27646,N_27587,N_27435);
nor U27647 (N_27647,N_27506,N_27423);
xnor U27648 (N_27648,N_27473,N_27429);
nand U27649 (N_27649,N_27577,N_27442);
or U27650 (N_27650,N_27571,N_27552);
nand U27651 (N_27651,N_27566,N_27468);
nand U27652 (N_27652,N_27597,N_27502);
nor U27653 (N_27653,N_27484,N_27541);
nor U27654 (N_27654,N_27478,N_27517);
nand U27655 (N_27655,N_27535,N_27482);
nand U27656 (N_27656,N_27449,N_27498);
xnor U27657 (N_27657,N_27433,N_27592);
nand U27658 (N_27658,N_27417,N_27469);
or U27659 (N_27659,N_27519,N_27450);
nor U27660 (N_27660,N_27434,N_27527);
and U27661 (N_27661,N_27551,N_27563);
or U27662 (N_27662,N_27419,N_27452);
nor U27663 (N_27663,N_27568,N_27460);
nand U27664 (N_27664,N_27503,N_27466);
nand U27665 (N_27665,N_27579,N_27454);
nand U27666 (N_27666,N_27409,N_27427);
or U27667 (N_27667,N_27431,N_27540);
and U27668 (N_27668,N_27493,N_27573);
or U27669 (N_27669,N_27485,N_27522);
nand U27670 (N_27670,N_27462,N_27512);
nand U27671 (N_27671,N_27475,N_27421);
xnor U27672 (N_27672,N_27569,N_27426);
xnor U27673 (N_27673,N_27455,N_27590);
xor U27674 (N_27674,N_27463,N_27530);
nand U27675 (N_27675,N_27401,N_27586);
nor U27676 (N_27676,N_27561,N_27448);
nand U27677 (N_27677,N_27432,N_27520);
and U27678 (N_27678,N_27533,N_27529);
and U27679 (N_27679,N_27539,N_27439);
nor U27680 (N_27680,N_27504,N_27414);
nor U27681 (N_27681,N_27583,N_27481);
nor U27682 (N_27682,N_27521,N_27589);
xor U27683 (N_27683,N_27496,N_27425);
nor U27684 (N_27684,N_27514,N_27536);
and U27685 (N_27685,N_27501,N_27554);
xor U27686 (N_27686,N_27510,N_27547);
nor U27687 (N_27687,N_27483,N_27574);
and U27688 (N_27688,N_27594,N_27471);
xnor U27689 (N_27689,N_27581,N_27553);
nor U27690 (N_27690,N_27532,N_27418);
or U27691 (N_27691,N_27525,N_27489);
and U27692 (N_27692,N_27438,N_27446);
xor U27693 (N_27693,N_27467,N_27560);
nand U27694 (N_27694,N_27598,N_27464);
nor U27695 (N_27695,N_27516,N_27430);
xor U27696 (N_27696,N_27445,N_27436);
xnor U27697 (N_27697,N_27515,N_27457);
nand U27698 (N_27698,N_27491,N_27474);
xor U27699 (N_27699,N_27545,N_27537);
or U27700 (N_27700,N_27579,N_27446);
nor U27701 (N_27701,N_27470,N_27426);
xnor U27702 (N_27702,N_27580,N_27456);
and U27703 (N_27703,N_27466,N_27415);
and U27704 (N_27704,N_27589,N_27464);
and U27705 (N_27705,N_27497,N_27515);
or U27706 (N_27706,N_27565,N_27414);
and U27707 (N_27707,N_27492,N_27532);
or U27708 (N_27708,N_27593,N_27589);
and U27709 (N_27709,N_27457,N_27571);
nand U27710 (N_27710,N_27565,N_27442);
nand U27711 (N_27711,N_27433,N_27577);
nor U27712 (N_27712,N_27547,N_27422);
and U27713 (N_27713,N_27592,N_27574);
xor U27714 (N_27714,N_27523,N_27529);
xor U27715 (N_27715,N_27534,N_27554);
nand U27716 (N_27716,N_27520,N_27525);
or U27717 (N_27717,N_27457,N_27532);
and U27718 (N_27718,N_27482,N_27593);
xor U27719 (N_27719,N_27445,N_27591);
or U27720 (N_27720,N_27556,N_27502);
xor U27721 (N_27721,N_27493,N_27413);
or U27722 (N_27722,N_27584,N_27498);
or U27723 (N_27723,N_27519,N_27459);
nand U27724 (N_27724,N_27547,N_27490);
xnor U27725 (N_27725,N_27519,N_27406);
xor U27726 (N_27726,N_27599,N_27591);
and U27727 (N_27727,N_27401,N_27486);
nor U27728 (N_27728,N_27582,N_27590);
xnor U27729 (N_27729,N_27564,N_27450);
and U27730 (N_27730,N_27405,N_27517);
or U27731 (N_27731,N_27471,N_27491);
xor U27732 (N_27732,N_27449,N_27440);
or U27733 (N_27733,N_27548,N_27566);
nor U27734 (N_27734,N_27596,N_27543);
nor U27735 (N_27735,N_27548,N_27539);
or U27736 (N_27736,N_27515,N_27561);
nor U27737 (N_27737,N_27514,N_27427);
xor U27738 (N_27738,N_27520,N_27497);
and U27739 (N_27739,N_27529,N_27581);
nor U27740 (N_27740,N_27420,N_27578);
nor U27741 (N_27741,N_27534,N_27406);
nor U27742 (N_27742,N_27575,N_27540);
xnor U27743 (N_27743,N_27461,N_27449);
nor U27744 (N_27744,N_27530,N_27533);
xnor U27745 (N_27745,N_27513,N_27490);
xor U27746 (N_27746,N_27552,N_27564);
xor U27747 (N_27747,N_27564,N_27587);
nand U27748 (N_27748,N_27518,N_27414);
nand U27749 (N_27749,N_27523,N_27459);
and U27750 (N_27750,N_27597,N_27524);
nor U27751 (N_27751,N_27503,N_27476);
nand U27752 (N_27752,N_27406,N_27423);
xor U27753 (N_27753,N_27492,N_27405);
xnor U27754 (N_27754,N_27503,N_27444);
nand U27755 (N_27755,N_27516,N_27547);
and U27756 (N_27756,N_27474,N_27570);
or U27757 (N_27757,N_27542,N_27492);
and U27758 (N_27758,N_27565,N_27531);
nand U27759 (N_27759,N_27587,N_27559);
xnor U27760 (N_27760,N_27423,N_27427);
or U27761 (N_27761,N_27547,N_27572);
nand U27762 (N_27762,N_27472,N_27554);
and U27763 (N_27763,N_27461,N_27465);
xor U27764 (N_27764,N_27401,N_27547);
xor U27765 (N_27765,N_27461,N_27570);
nor U27766 (N_27766,N_27484,N_27576);
and U27767 (N_27767,N_27520,N_27553);
and U27768 (N_27768,N_27488,N_27591);
or U27769 (N_27769,N_27400,N_27410);
and U27770 (N_27770,N_27518,N_27550);
xnor U27771 (N_27771,N_27589,N_27523);
and U27772 (N_27772,N_27519,N_27505);
or U27773 (N_27773,N_27419,N_27569);
nand U27774 (N_27774,N_27473,N_27486);
and U27775 (N_27775,N_27416,N_27551);
and U27776 (N_27776,N_27514,N_27412);
xor U27777 (N_27777,N_27588,N_27473);
xor U27778 (N_27778,N_27443,N_27483);
xor U27779 (N_27779,N_27502,N_27481);
and U27780 (N_27780,N_27444,N_27467);
and U27781 (N_27781,N_27579,N_27489);
or U27782 (N_27782,N_27434,N_27520);
nand U27783 (N_27783,N_27508,N_27494);
xor U27784 (N_27784,N_27442,N_27535);
xor U27785 (N_27785,N_27429,N_27405);
nor U27786 (N_27786,N_27537,N_27477);
or U27787 (N_27787,N_27514,N_27552);
or U27788 (N_27788,N_27546,N_27531);
nor U27789 (N_27789,N_27414,N_27588);
xor U27790 (N_27790,N_27596,N_27540);
or U27791 (N_27791,N_27551,N_27543);
or U27792 (N_27792,N_27418,N_27455);
xor U27793 (N_27793,N_27491,N_27423);
nand U27794 (N_27794,N_27510,N_27593);
nand U27795 (N_27795,N_27542,N_27590);
or U27796 (N_27796,N_27534,N_27464);
nor U27797 (N_27797,N_27451,N_27519);
nor U27798 (N_27798,N_27463,N_27408);
nand U27799 (N_27799,N_27549,N_27481);
and U27800 (N_27800,N_27735,N_27604);
or U27801 (N_27801,N_27773,N_27642);
xor U27802 (N_27802,N_27667,N_27613);
nand U27803 (N_27803,N_27679,N_27633);
nand U27804 (N_27804,N_27745,N_27699);
or U27805 (N_27805,N_27662,N_27719);
or U27806 (N_27806,N_27713,N_27686);
xor U27807 (N_27807,N_27704,N_27720);
xnor U27808 (N_27808,N_27723,N_27619);
nand U27809 (N_27809,N_27792,N_27691);
or U27810 (N_27810,N_27643,N_27660);
and U27811 (N_27811,N_27779,N_27612);
or U27812 (N_27812,N_27651,N_27672);
or U27813 (N_27813,N_27718,N_27728);
xnor U27814 (N_27814,N_27734,N_27602);
nor U27815 (N_27815,N_27659,N_27764);
xnor U27816 (N_27816,N_27702,N_27614);
xor U27817 (N_27817,N_27684,N_27761);
nand U27818 (N_27818,N_27778,N_27716);
or U27819 (N_27819,N_27750,N_27653);
xor U27820 (N_27820,N_27776,N_27796);
or U27821 (N_27821,N_27687,N_27656);
nor U27822 (N_27822,N_27741,N_27682);
or U27823 (N_27823,N_27756,N_27798);
nor U27824 (N_27824,N_27603,N_27782);
xor U27825 (N_27825,N_27769,N_27799);
nor U27826 (N_27826,N_27695,N_27610);
nand U27827 (N_27827,N_27705,N_27710);
nor U27828 (N_27828,N_27664,N_27729);
xor U27829 (N_27829,N_27742,N_27657);
and U27830 (N_27830,N_27683,N_27738);
xor U27831 (N_27831,N_27681,N_27701);
nand U27832 (N_27832,N_27789,N_27712);
nor U27833 (N_27833,N_27675,N_27618);
or U27834 (N_27834,N_27673,N_27722);
nor U27835 (N_27835,N_27771,N_27639);
nand U27836 (N_27836,N_27770,N_27606);
nand U27837 (N_27837,N_27665,N_27632);
or U27838 (N_27838,N_27647,N_27755);
or U27839 (N_27839,N_27669,N_27670);
nor U27840 (N_27840,N_27746,N_27630);
nor U27841 (N_27841,N_27600,N_27760);
and U27842 (N_27842,N_27706,N_27752);
or U27843 (N_27843,N_27624,N_27644);
and U27844 (N_27844,N_27768,N_27617);
nor U27845 (N_27845,N_27703,N_27724);
and U27846 (N_27846,N_27715,N_27783);
nor U27847 (N_27847,N_27786,N_27766);
nor U27848 (N_27848,N_27652,N_27790);
nand U27849 (N_27849,N_27747,N_27793);
or U27850 (N_27850,N_27698,N_27607);
nand U27851 (N_27851,N_27711,N_27621);
nor U27852 (N_27852,N_27616,N_27772);
nor U27853 (N_27853,N_27692,N_27655);
and U27854 (N_27854,N_27787,N_27737);
or U27855 (N_27855,N_27753,N_27744);
or U27856 (N_27856,N_27714,N_27775);
nor U27857 (N_27857,N_27763,N_27676);
xor U27858 (N_27858,N_27707,N_27688);
nor U27859 (N_27859,N_27725,N_27641);
and U27860 (N_27860,N_27663,N_27748);
nor U27861 (N_27861,N_27661,N_27700);
or U27862 (N_27862,N_27726,N_27650);
xnor U27863 (N_27863,N_27637,N_27762);
and U27864 (N_27864,N_27629,N_27791);
nor U27865 (N_27865,N_27757,N_27777);
and U27866 (N_27866,N_27674,N_27636);
and U27867 (N_27867,N_27708,N_27645);
nand U27868 (N_27868,N_27709,N_27611);
and U27869 (N_27869,N_27623,N_27781);
nand U27870 (N_27870,N_27758,N_27654);
nand U27871 (N_27871,N_27767,N_27615);
or U27872 (N_27872,N_27733,N_27740);
and U27873 (N_27873,N_27626,N_27795);
or U27874 (N_27874,N_27690,N_27666);
nor U27875 (N_27875,N_27658,N_27634);
nand U27876 (N_27876,N_27731,N_27794);
nor U27877 (N_27877,N_27622,N_27627);
xor U27878 (N_27878,N_27721,N_27727);
or U27879 (N_27879,N_27739,N_27668);
and U27880 (N_27880,N_27736,N_27749);
nand U27881 (N_27881,N_27671,N_27717);
xor U27882 (N_27882,N_27696,N_27765);
and U27883 (N_27883,N_27774,N_27677);
or U27884 (N_27884,N_27620,N_27678);
xor U27885 (N_27885,N_27635,N_27638);
nor U27886 (N_27886,N_27693,N_27759);
and U27887 (N_27887,N_27625,N_27743);
nand U27888 (N_27888,N_27730,N_27689);
nand U27889 (N_27889,N_27780,N_27649);
and U27890 (N_27890,N_27694,N_27732);
and U27891 (N_27891,N_27785,N_27605);
and U27892 (N_27892,N_27640,N_27609);
and U27893 (N_27893,N_27628,N_27697);
xor U27894 (N_27894,N_27648,N_27646);
xor U27895 (N_27895,N_27631,N_27754);
xor U27896 (N_27896,N_27751,N_27788);
or U27897 (N_27897,N_27680,N_27608);
nand U27898 (N_27898,N_27601,N_27797);
nor U27899 (N_27899,N_27685,N_27784);
nand U27900 (N_27900,N_27742,N_27698);
xnor U27901 (N_27901,N_27713,N_27620);
nor U27902 (N_27902,N_27727,N_27603);
nor U27903 (N_27903,N_27746,N_27601);
or U27904 (N_27904,N_27602,N_27699);
xor U27905 (N_27905,N_27659,N_27664);
xnor U27906 (N_27906,N_27681,N_27664);
or U27907 (N_27907,N_27763,N_27632);
and U27908 (N_27908,N_27667,N_27755);
nor U27909 (N_27909,N_27610,N_27708);
or U27910 (N_27910,N_27771,N_27791);
nand U27911 (N_27911,N_27669,N_27731);
nor U27912 (N_27912,N_27688,N_27612);
and U27913 (N_27913,N_27701,N_27762);
nand U27914 (N_27914,N_27707,N_27712);
xnor U27915 (N_27915,N_27709,N_27641);
xor U27916 (N_27916,N_27766,N_27623);
and U27917 (N_27917,N_27659,N_27742);
xor U27918 (N_27918,N_27759,N_27622);
or U27919 (N_27919,N_27752,N_27794);
nand U27920 (N_27920,N_27771,N_27681);
nor U27921 (N_27921,N_27697,N_27603);
and U27922 (N_27922,N_27794,N_27705);
or U27923 (N_27923,N_27644,N_27697);
nor U27924 (N_27924,N_27743,N_27674);
and U27925 (N_27925,N_27705,N_27784);
nor U27926 (N_27926,N_27736,N_27647);
xnor U27927 (N_27927,N_27604,N_27644);
nand U27928 (N_27928,N_27702,N_27706);
or U27929 (N_27929,N_27697,N_27777);
nor U27930 (N_27930,N_27622,N_27707);
nor U27931 (N_27931,N_27654,N_27636);
nand U27932 (N_27932,N_27749,N_27635);
nor U27933 (N_27933,N_27681,N_27776);
nor U27934 (N_27934,N_27696,N_27776);
and U27935 (N_27935,N_27795,N_27720);
and U27936 (N_27936,N_27621,N_27749);
or U27937 (N_27937,N_27768,N_27733);
xor U27938 (N_27938,N_27601,N_27661);
nor U27939 (N_27939,N_27743,N_27745);
or U27940 (N_27940,N_27628,N_27740);
nor U27941 (N_27941,N_27680,N_27692);
and U27942 (N_27942,N_27795,N_27610);
and U27943 (N_27943,N_27742,N_27669);
xnor U27944 (N_27944,N_27696,N_27690);
nor U27945 (N_27945,N_27686,N_27726);
or U27946 (N_27946,N_27740,N_27795);
and U27947 (N_27947,N_27651,N_27774);
nand U27948 (N_27948,N_27690,N_27633);
xor U27949 (N_27949,N_27796,N_27618);
nand U27950 (N_27950,N_27681,N_27794);
nand U27951 (N_27951,N_27602,N_27792);
nand U27952 (N_27952,N_27784,N_27736);
nor U27953 (N_27953,N_27750,N_27627);
nor U27954 (N_27954,N_27648,N_27695);
nand U27955 (N_27955,N_27776,N_27741);
or U27956 (N_27956,N_27626,N_27791);
xor U27957 (N_27957,N_27636,N_27657);
xnor U27958 (N_27958,N_27726,N_27709);
nor U27959 (N_27959,N_27641,N_27626);
and U27960 (N_27960,N_27695,N_27758);
nand U27961 (N_27961,N_27694,N_27728);
nor U27962 (N_27962,N_27760,N_27715);
xor U27963 (N_27963,N_27643,N_27762);
or U27964 (N_27964,N_27739,N_27797);
or U27965 (N_27965,N_27706,N_27693);
nand U27966 (N_27966,N_27683,N_27674);
and U27967 (N_27967,N_27768,N_27787);
nand U27968 (N_27968,N_27794,N_27648);
nor U27969 (N_27969,N_27681,N_27761);
and U27970 (N_27970,N_27665,N_27739);
nor U27971 (N_27971,N_27724,N_27799);
nor U27972 (N_27972,N_27643,N_27773);
xnor U27973 (N_27973,N_27764,N_27627);
nand U27974 (N_27974,N_27602,N_27637);
nand U27975 (N_27975,N_27651,N_27683);
nand U27976 (N_27976,N_27694,N_27782);
or U27977 (N_27977,N_27722,N_27689);
nor U27978 (N_27978,N_27663,N_27618);
xnor U27979 (N_27979,N_27614,N_27762);
nand U27980 (N_27980,N_27781,N_27783);
nand U27981 (N_27981,N_27606,N_27603);
xor U27982 (N_27982,N_27780,N_27788);
or U27983 (N_27983,N_27617,N_27798);
xor U27984 (N_27984,N_27734,N_27625);
and U27985 (N_27985,N_27712,N_27646);
and U27986 (N_27986,N_27764,N_27682);
nor U27987 (N_27987,N_27635,N_27710);
and U27988 (N_27988,N_27787,N_27730);
and U27989 (N_27989,N_27704,N_27694);
nand U27990 (N_27990,N_27658,N_27654);
and U27991 (N_27991,N_27640,N_27743);
or U27992 (N_27992,N_27680,N_27623);
nand U27993 (N_27993,N_27600,N_27772);
nand U27994 (N_27994,N_27690,N_27677);
xor U27995 (N_27995,N_27776,N_27740);
nand U27996 (N_27996,N_27714,N_27705);
or U27997 (N_27997,N_27782,N_27712);
and U27998 (N_27998,N_27737,N_27618);
and U27999 (N_27999,N_27745,N_27617);
or U28000 (N_28000,N_27853,N_27812);
or U28001 (N_28001,N_27939,N_27978);
or U28002 (N_28002,N_27870,N_27886);
nor U28003 (N_28003,N_27893,N_27864);
xor U28004 (N_28004,N_27969,N_27865);
and U28005 (N_28005,N_27968,N_27894);
nand U28006 (N_28006,N_27892,N_27847);
and U28007 (N_28007,N_27973,N_27842);
nor U28008 (N_28008,N_27945,N_27900);
nand U28009 (N_28009,N_27962,N_27868);
and U28010 (N_28010,N_27856,N_27983);
and U28011 (N_28011,N_27899,N_27952);
xor U28012 (N_28012,N_27819,N_27876);
nor U28013 (N_28013,N_27902,N_27937);
xnor U28014 (N_28014,N_27875,N_27990);
nand U28015 (N_28015,N_27877,N_27951);
nor U28016 (N_28016,N_27974,N_27841);
or U28017 (N_28017,N_27979,N_27928);
and U28018 (N_28018,N_27848,N_27882);
and U28019 (N_28019,N_27906,N_27963);
nand U28020 (N_28020,N_27895,N_27820);
xnor U28021 (N_28021,N_27992,N_27904);
or U28022 (N_28022,N_27985,N_27913);
xnor U28023 (N_28023,N_27924,N_27843);
and U28024 (N_28024,N_27956,N_27949);
xor U28025 (N_28025,N_27818,N_27933);
xnor U28026 (N_28026,N_27869,N_27891);
xor U28027 (N_28027,N_27827,N_27830);
or U28028 (N_28028,N_27833,N_27946);
nand U28029 (N_28029,N_27936,N_27917);
nor U28030 (N_28030,N_27821,N_27878);
xnor U28031 (N_28031,N_27845,N_27887);
nor U28032 (N_28032,N_27911,N_27925);
and U28033 (N_28033,N_27994,N_27871);
nor U28034 (N_28034,N_27972,N_27987);
or U28035 (N_28035,N_27800,N_27953);
or U28036 (N_28036,N_27822,N_27955);
nor U28037 (N_28037,N_27826,N_27967);
or U28038 (N_28038,N_27890,N_27942);
and U28039 (N_28039,N_27857,N_27885);
nand U28040 (N_28040,N_27998,N_27941);
or U28041 (N_28041,N_27816,N_27808);
xor U28042 (N_28042,N_27971,N_27834);
or U28043 (N_28043,N_27835,N_27923);
xnor U28044 (N_28044,N_27991,N_27806);
or U28045 (N_28045,N_27813,N_27996);
and U28046 (N_28046,N_27907,N_27844);
or U28047 (N_28047,N_27918,N_27919);
xnor U28048 (N_28048,N_27839,N_27881);
xnor U28049 (N_28049,N_27914,N_27932);
or U28050 (N_28050,N_27905,N_27889);
xor U28051 (N_28051,N_27873,N_27921);
or U28052 (N_28052,N_27961,N_27926);
xnor U28053 (N_28053,N_27836,N_27849);
nor U28054 (N_28054,N_27929,N_27840);
or U28055 (N_28055,N_27807,N_27938);
or U28056 (N_28056,N_27901,N_27986);
or U28057 (N_28057,N_27935,N_27815);
nand U28058 (N_28058,N_27993,N_27898);
xor U28059 (N_28059,N_27954,N_27861);
and U28060 (N_28060,N_27838,N_27984);
nor U28061 (N_28061,N_27947,N_27960);
and U28062 (N_28062,N_27872,N_27817);
nand U28063 (N_28063,N_27866,N_27980);
and U28064 (N_28064,N_27988,N_27943);
or U28065 (N_28065,N_27888,N_27896);
nand U28066 (N_28066,N_27837,N_27803);
nand U28067 (N_28067,N_27897,N_27977);
and U28068 (N_28068,N_27832,N_27964);
xnor U28069 (N_28069,N_27852,N_27965);
nand U28070 (N_28070,N_27805,N_27916);
nor U28071 (N_28071,N_27809,N_27874);
nor U28072 (N_28072,N_27940,N_27884);
or U28073 (N_28073,N_27944,N_27831);
nand U28074 (N_28074,N_27824,N_27959);
nand U28075 (N_28075,N_27851,N_27846);
nor U28076 (N_28076,N_27966,N_27999);
nor U28077 (N_28077,N_27931,N_27920);
nor U28078 (N_28078,N_27934,N_27860);
xnor U28079 (N_28079,N_27976,N_27981);
or U28080 (N_28080,N_27829,N_27854);
or U28081 (N_28081,N_27867,N_27850);
or U28082 (N_28082,N_27823,N_27950);
nand U28083 (N_28083,N_27863,N_27948);
or U28084 (N_28084,N_27903,N_27862);
nor U28085 (N_28085,N_27982,N_27927);
or U28086 (N_28086,N_27915,N_27912);
nand U28087 (N_28087,N_27814,N_27957);
and U28088 (N_28088,N_27930,N_27810);
nand U28089 (N_28089,N_27811,N_27958);
xor U28090 (N_28090,N_27855,N_27802);
or U28091 (N_28091,N_27995,N_27970);
xnor U28092 (N_28092,N_27989,N_27828);
nand U28093 (N_28093,N_27909,N_27879);
nor U28094 (N_28094,N_27997,N_27858);
xnor U28095 (N_28095,N_27883,N_27801);
xor U28096 (N_28096,N_27908,N_27922);
and U28097 (N_28097,N_27859,N_27804);
xnor U28098 (N_28098,N_27975,N_27910);
nand U28099 (N_28099,N_27880,N_27825);
nor U28100 (N_28100,N_27941,N_27815);
and U28101 (N_28101,N_27870,N_27842);
or U28102 (N_28102,N_27823,N_27828);
nor U28103 (N_28103,N_27983,N_27864);
and U28104 (N_28104,N_27908,N_27845);
or U28105 (N_28105,N_27913,N_27870);
or U28106 (N_28106,N_27940,N_27831);
nor U28107 (N_28107,N_27957,N_27952);
and U28108 (N_28108,N_27929,N_27822);
nor U28109 (N_28109,N_27965,N_27866);
nor U28110 (N_28110,N_27969,N_27938);
and U28111 (N_28111,N_27806,N_27891);
and U28112 (N_28112,N_27970,N_27806);
and U28113 (N_28113,N_27887,N_27964);
or U28114 (N_28114,N_27909,N_27978);
xnor U28115 (N_28115,N_27910,N_27839);
nor U28116 (N_28116,N_27830,N_27813);
and U28117 (N_28117,N_27849,N_27949);
nor U28118 (N_28118,N_27985,N_27992);
and U28119 (N_28119,N_27848,N_27904);
and U28120 (N_28120,N_27877,N_27815);
xnor U28121 (N_28121,N_27871,N_27824);
nand U28122 (N_28122,N_27851,N_27844);
and U28123 (N_28123,N_27928,N_27938);
nand U28124 (N_28124,N_27957,N_27802);
and U28125 (N_28125,N_27829,N_27913);
nand U28126 (N_28126,N_27992,N_27990);
xnor U28127 (N_28127,N_27947,N_27907);
or U28128 (N_28128,N_27847,N_27849);
nand U28129 (N_28129,N_27980,N_27812);
and U28130 (N_28130,N_27899,N_27984);
and U28131 (N_28131,N_27922,N_27945);
and U28132 (N_28132,N_27983,N_27885);
xnor U28133 (N_28133,N_27883,N_27924);
nor U28134 (N_28134,N_27807,N_27867);
and U28135 (N_28135,N_27900,N_27924);
nor U28136 (N_28136,N_27873,N_27946);
and U28137 (N_28137,N_27821,N_27931);
and U28138 (N_28138,N_27991,N_27860);
xnor U28139 (N_28139,N_27814,N_27822);
nor U28140 (N_28140,N_27937,N_27849);
and U28141 (N_28141,N_27824,N_27955);
nor U28142 (N_28142,N_27937,N_27882);
xor U28143 (N_28143,N_27935,N_27849);
nor U28144 (N_28144,N_27804,N_27855);
or U28145 (N_28145,N_27823,N_27811);
xnor U28146 (N_28146,N_27961,N_27851);
xor U28147 (N_28147,N_27917,N_27896);
nand U28148 (N_28148,N_27912,N_27979);
nand U28149 (N_28149,N_27983,N_27806);
xor U28150 (N_28150,N_27987,N_27857);
or U28151 (N_28151,N_27929,N_27939);
xor U28152 (N_28152,N_27892,N_27984);
or U28153 (N_28153,N_27917,N_27987);
nand U28154 (N_28154,N_27860,N_27863);
nor U28155 (N_28155,N_27888,N_27994);
nand U28156 (N_28156,N_27890,N_27826);
or U28157 (N_28157,N_27995,N_27893);
nand U28158 (N_28158,N_27975,N_27922);
nand U28159 (N_28159,N_27835,N_27891);
or U28160 (N_28160,N_27866,N_27989);
xnor U28161 (N_28161,N_27975,N_27946);
and U28162 (N_28162,N_27904,N_27835);
and U28163 (N_28163,N_27895,N_27957);
or U28164 (N_28164,N_27802,N_27902);
nor U28165 (N_28165,N_27831,N_27966);
and U28166 (N_28166,N_27940,N_27871);
xor U28167 (N_28167,N_27899,N_27939);
or U28168 (N_28168,N_27917,N_27814);
nor U28169 (N_28169,N_27950,N_27943);
xor U28170 (N_28170,N_27930,N_27851);
and U28171 (N_28171,N_27921,N_27964);
nand U28172 (N_28172,N_27840,N_27826);
and U28173 (N_28173,N_27910,N_27982);
nand U28174 (N_28174,N_27849,N_27960);
or U28175 (N_28175,N_27943,N_27847);
xnor U28176 (N_28176,N_27890,N_27944);
nor U28177 (N_28177,N_27950,N_27884);
nor U28178 (N_28178,N_27969,N_27810);
and U28179 (N_28179,N_27850,N_27946);
nand U28180 (N_28180,N_27962,N_27816);
and U28181 (N_28181,N_27897,N_27989);
and U28182 (N_28182,N_27954,N_27841);
nand U28183 (N_28183,N_27967,N_27801);
xor U28184 (N_28184,N_27822,N_27896);
nand U28185 (N_28185,N_27901,N_27991);
and U28186 (N_28186,N_27827,N_27923);
or U28187 (N_28187,N_27864,N_27900);
or U28188 (N_28188,N_27872,N_27969);
and U28189 (N_28189,N_27936,N_27995);
nor U28190 (N_28190,N_27831,N_27904);
nor U28191 (N_28191,N_27971,N_27970);
or U28192 (N_28192,N_27881,N_27965);
or U28193 (N_28193,N_27893,N_27980);
and U28194 (N_28194,N_27990,N_27901);
xor U28195 (N_28195,N_27802,N_27987);
or U28196 (N_28196,N_27832,N_27939);
and U28197 (N_28197,N_27985,N_27951);
xor U28198 (N_28198,N_27889,N_27945);
and U28199 (N_28199,N_27924,N_27960);
nand U28200 (N_28200,N_28107,N_28135);
or U28201 (N_28201,N_28067,N_28109);
or U28202 (N_28202,N_28184,N_28087);
xor U28203 (N_28203,N_28185,N_28144);
nor U28204 (N_28204,N_28122,N_28098);
nand U28205 (N_28205,N_28027,N_28175);
nor U28206 (N_28206,N_28069,N_28156);
nor U28207 (N_28207,N_28128,N_28177);
and U28208 (N_28208,N_28035,N_28052);
and U28209 (N_28209,N_28031,N_28081);
xnor U28210 (N_28210,N_28149,N_28108);
or U28211 (N_28211,N_28025,N_28024);
xor U28212 (N_28212,N_28050,N_28017);
xor U28213 (N_28213,N_28152,N_28068);
nor U28214 (N_28214,N_28145,N_28103);
nor U28215 (N_28215,N_28170,N_28089);
and U28216 (N_28216,N_28001,N_28125);
and U28217 (N_28217,N_28095,N_28080);
and U28218 (N_28218,N_28142,N_28009);
nor U28219 (N_28219,N_28139,N_28063);
or U28220 (N_28220,N_28193,N_28061);
nor U28221 (N_28221,N_28096,N_28165);
nor U28222 (N_28222,N_28046,N_28190);
nor U28223 (N_28223,N_28037,N_28118);
or U28224 (N_28224,N_28121,N_28032);
nor U28225 (N_28225,N_28070,N_28016);
nand U28226 (N_28226,N_28191,N_28143);
nor U28227 (N_28227,N_28011,N_28041);
or U28228 (N_28228,N_28124,N_28051);
and U28229 (N_28229,N_28137,N_28075);
xnor U28230 (N_28230,N_28010,N_28198);
xnor U28231 (N_28231,N_28100,N_28073);
nor U28232 (N_28232,N_28166,N_28043);
and U28233 (N_28233,N_28040,N_28072);
nor U28234 (N_28234,N_28172,N_28120);
nand U28235 (N_28235,N_28059,N_28181);
or U28236 (N_28236,N_28000,N_28048);
xnor U28237 (N_28237,N_28007,N_28130);
or U28238 (N_28238,N_28173,N_28162);
nor U28239 (N_28239,N_28161,N_28008);
nor U28240 (N_28240,N_28044,N_28183);
nand U28241 (N_28241,N_28134,N_28133);
nor U28242 (N_28242,N_28150,N_28058);
or U28243 (N_28243,N_28112,N_28110);
or U28244 (N_28244,N_28084,N_28082);
and U28245 (N_28245,N_28187,N_28194);
nand U28246 (N_28246,N_28160,N_28003);
xor U28247 (N_28247,N_28029,N_28049);
and U28248 (N_28248,N_28105,N_28138);
nand U28249 (N_28249,N_28101,N_28151);
nand U28250 (N_28250,N_28195,N_28197);
nand U28251 (N_28251,N_28126,N_28086);
and U28252 (N_28252,N_28127,N_28053);
xor U28253 (N_28253,N_28180,N_28039);
and U28254 (N_28254,N_28093,N_28113);
xor U28255 (N_28255,N_28056,N_28085);
or U28256 (N_28256,N_28147,N_28074);
nand U28257 (N_28257,N_28163,N_28178);
xor U28258 (N_28258,N_28083,N_28090);
xor U28259 (N_28259,N_28182,N_28167);
or U28260 (N_28260,N_28088,N_28077);
nand U28261 (N_28261,N_28034,N_28057);
and U28262 (N_28262,N_28091,N_28132);
or U28263 (N_28263,N_28131,N_28140);
xor U28264 (N_28264,N_28021,N_28168);
or U28265 (N_28265,N_28060,N_28028);
nand U28266 (N_28266,N_28111,N_28176);
and U28267 (N_28267,N_28171,N_28064);
nor U28268 (N_28268,N_28079,N_28076);
nor U28269 (N_28269,N_28045,N_28155);
xnor U28270 (N_28270,N_28136,N_28106);
nand U28271 (N_28271,N_28119,N_28097);
nor U28272 (N_28272,N_28006,N_28023);
and U28273 (N_28273,N_28146,N_28141);
nor U28274 (N_28274,N_28099,N_28174);
xnor U28275 (N_28275,N_28129,N_28164);
nand U28276 (N_28276,N_28192,N_28158);
nand U28277 (N_28277,N_28196,N_28123);
and U28278 (N_28278,N_28116,N_28199);
or U28279 (N_28279,N_28015,N_28047);
xnor U28280 (N_28280,N_28018,N_28154);
and U28281 (N_28281,N_28114,N_28033);
xor U28282 (N_28282,N_28022,N_28012);
xor U28283 (N_28283,N_28102,N_28071);
nand U28284 (N_28284,N_28159,N_28117);
nand U28285 (N_28285,N_28094,N_28054);
xor U28286 (N_28286,N_28188,N_28019);
nand U28287 (N_28287,N_28169,N_28153);
nand U28288 (N_28288,N_28014,N_28038);
and U28289 (N_28289,N_28179,N_28013);
or U28290 (N_28290,N_28002,N_28004);
nand U28291 (N_28291,N_28078,N_28042);
or U28292 (N_28292,N_28026,N_28066);
or U28293 (N_28293,N_28020,N_28036);
nand U28294 (N_28294,N_28104,N_28189);
nand U28295 (N_28295,N_28005,N_28065);
nand U28296 (N_28296,N_28055,N_28115);
nor U28297 (N_28297,N_28030,N_28092);
xor U28298 (N_28298,N_28148,N_28157);
or U28299 (N_28299,N_28186,N_28062);
xor U28300 (N_28300,N_28129,N_28118);
nand U28301 (N_28301,N_28136,N_28176);
and U28302 (N_28302,N_28097,N_28134);
nor U28303 (N_28303,N_28179,N_28109);
or U28304 (N_28304,N_28184,N_28068);
nor U28305 (N_28305,N_28052,N_28068);
or U28306 (N_28306,N_28116,N_28011);
xor U28307 (N_28307,N_28135,N_28126);
and U28308 (N_28308,N_28060,N_28188);
nand U28309 (N_28309,N_28119,N_28015);
and U28310 (N_28310,N_28030,N_28158);
or U28311 (N_28311,N_28026,N_28115);
nor U28312 (N_28312,N_28016,N_28138);
xnor U28313 (N_28313,N_28009,N_28141);
xor U28314 (N_28314,N_28183,N_28154);
nand U28315 (N_28315,N_28095,N_28199);
xor U28316 (N_28316,N_28073,N_28124);
nand U28317 (N_28317,N_28161,N_28104);
or U28318 (N_28318,N_28128,N_28088);
xor U28319 (N_28319,N_28148,N_28075);
xnor U28320 (N_28320,N_28181,N_28097);
nor U28321 (N_28321,N_28072,N_28039);
nor U28322 (N_28322,N_28177,N_28139);
xor U28323 (N_28323,N_28069,N_28183);
nor U28324 (N_28324,N_28082,N_28121);
xor U28325 (N_28325,N_28193,N_28090);
xor U28326 (N_28326,N_28027,N_28053);
nor U28327 (N_28327,N_28106,N_28060);
and U28328 (N_28328,N_28079,N_28034);
and U28329 (N_28329,N_28046,N_28197);
xor U28330 (N_28330,N_28166,N_28103);
and U28331 (N_28331,N_28018,N_28157);
or U28332 (N_28332,N_28180,N_28129);
xnor U28333 (N_28333,N_28180,N_28089);
xor U28334 (N_28334,N_28188,N_28182);
xnor U28335 (N_28335,N_28005,N_28193);
nor U28336 (N_28336,N_28091,N_28043);
nand U28337 (N_28337,N_28056,N_28136);
nand U28338 (N_28338,N_28194,N_28048);
nand U28339 (N_28339,N_28148,N_28188);
nor U28340 (N_28340,N_28082,N_28114);
xor U28341 (N_28341,N_28179,N_28137);
or U28342 (N_28342,N_28010,N_28079);
nor U28343 (N_28343,N_28008,N_28118);
and U28344 (N_28344,N_28109,N_28103);
nor U28345 (N_28345,N_28141,N_28140);
or U28346 (N_28346,N_28051,N_28116);
xor U28347 (N_28347,N_28017,N_28086);
nor U28348 (N_28348,N_28063,N_28120);
and U28349 (N_28349,N_28035,N_28078);
nand U28350 (N_28350,N_28091,N_28089);
nand U28351 (N_28351,N_28104,N_28125);
or U28352 (N_28352,N_28031,N_28123);
nor U28353 (N_28353,N_28174,N_28117);
or U28354 (N_28354,N_28100,N_28016);
xor U28355 (N_28355,N_28000,N_28128);
and U28356 (N_28356,N_28111,N_28156);
and U28357 (N_28357,N_28134,N_28149);
xor U28358 (N_28358,N_28018,N_28052);
or U28359 (N_28359,N_28186,N_28114);
xor U28360 (N_28360,N_28030,N_28033);
and U28361 (N_28361,N_28017,N_28021);
and U28362 (N_28362,N_28120,N_28149);
nor U28363 (N_28363,N_28149,N_28088);
xnor U28364 (N_28364,N_28087,N_28073);
or U28365 (N_28365,N_28081,N_28100);
nor U28366 (N_28366,N_28187,N_28059);
nor U28367 (N_28367,N_28012,N_28081);
nand U28368 (N_28368,N_28031,N_28143);
or U28369 (N_28369,N_28121,N_28031);
nor U28370 (N_28370,N_28092,N_28058);
and U28371 (N_28371,N_28024,N_28043);
or U28372 (N_28372,N_28121,N_28034);
and U28373 (N_28373,N_28000,N_28028);
or U28374 (N_28374,N_28063,N_28069);
nor U28375 (N_28375,N_28081,N_28137);
xnor U28376 (N_28376,N_28129,N_28173);
nor U28377 (N_28377,N_28043,N_28002);
nand U28378 (N_28378,N_28086,N_28029);
or U28379 (N_28379,N_28045,N_28187);
and U28380 (N_28380,N_28113,N_28005);
nor U28381 (N_28381,N_28188,N_28172);
and U28382 (N_28382,N_28063,N_28056);
nand U28383 (N_28383,N_28029,N_28104);
nor U28384 (N_28384,N_28055,N_28022);
nor U28385 (N_28385,N_28181,N_28141);
xor U28386 (N_28386,N_28040,N_28023);
xor U28387 (N_28387,N_28052,N_28063);
or U28388 (N_28388,N_28094,N_28179);
or U28389 (N_28389,N_28054,N_28014);
xor U28390 (N_28390,N_28147,N_28002);
nand U28391 (N_28391,N_28102,N_28087);
and U28392 (N_28392,N_28137,N_28121);
xnor U28393 (N_28393,N_28052,N_28112);
or U28394 (N_28394,N_28100,N_28004);
and U28395 (N_28395,N_28034,N_28009);
or U28396 (N_28396,N_28026,N_28167);
xor U28397 (N_28397,N_28028,N_28118);
nor U28398 (N_28398,N_28107,N_28022);
nor U28399 (N_28399,N_28053,N_28089);
and U28400 (N_28400,N_28327,N_28361);
xor U28401 (N_28401,N_28366,N_28378);
and U28402 (N_28402,N_28301,N_28250);
and U28403 (N_28403,N_28395,N_28226);
and U28404 (N_28404,N_28217,N_28305);
nor U28405 (N_28405,N_28314,N_28285);
nand U28406 (N_28406,N_28221,N_28238);
nor U28407 (N_28407,N_28251,N_28295);
and U28408 (N_28408,N_28213,N_28368);
nor U28409 (N_28409,N_28304,N_28362);
nand U28410 (N_28410,N_28287,N_28268);
and U28411 (N_28411,N_28339,N_28271);
nor U28412 (N_28412,N_28324,N_28310);
nand U28413 (N_28413,N_28311,N_28234);
xnor U28414 (N_28414,N_28255,N_28222);
xor U28415 (N_28415,N_28261,N_28272);
or U28416 (N_28416,N_28203,N_28206);
xor U28417 (N_28417,N_28386,N_28210);
xor U28418 (N_28418,N_28244,N_28208);
nor U28419 (N_28419,N_28321,N_28320);
nand U28420 (N_28420,N_28354,N_28283);
xnor U28421 (N_28421,N_28214,N_28262);
and U28422 (N_28422,N_28307,N_28349);
and U28423 (N_28423,N_28230,N_28293);
nand U28424 (N_28424,N_28263,N_28325);
xnor U28425 (N_28425,N_28254,N_28298);
or U28426 (N_28426,N_28373,N_28355);
or U28427 (N_28427,N_28390,N_28278);
nor U28428 (N_28428,N_28236,N_28277);
and U28429 (N_28429,N_28223,N_28331);
and U28430 (N_28430,N_28359,N_28350);
and U28431 (N_28431,N_28356,N_28360);
and U28432 (N_28432,N_28227,N_28215);
xor U28433 (N_28433,N_28280,N_28351);
nand U28434 (N_28434,N_28205,N_28228);
or U28435 (N_28435,N_28302,N_28264);
nand U28436 (N_28436,N_28396,N_28201);
nor U28437 (N_28437,N_28398,N_28309);
nor U28438 (N_28438,N_28231,N_28303);
xnor U28439 (N_28439,N_28340,N_28383);
or U28440 (N_28440,N_28384,N_28211);
xor U28441 (N_28441,N_28367,N_28282);
xnor U28442 (N_28442,N_28241,N_28348);
nor U28443 (N_28443,N_28389,N_28218);
nor U28444 (N_28444,N_28393,N_28224);
nor U28445 (N_28445,N_28371,N_28300);
nand U28446 (N_28446,N_28358,N_28294);
xnor U28447 (N_28447,N_28332,N_28200);
nand U28448 (N_28448,N_28375,N_28265);
or U28449 (N_28449,N_28316,N_28353);
nand U28450 (N_28450,N_28388,N_28299);
or U28451 (N_28451,N_28275,N_28239);
or U28452 (N_28452,N_28394,N_28246);
or U28453 (N_28453,N_28343,N_28328);
or U28454 (N_28454,N_28336,N_28219);
or U28455 (N_28455,N_28240,N_28372);
nor U28456 (N_28456,N_28237,N_28274);
nor U28457 (N_28457,N_28399,N_28288);
nor U28458 (N_28458,N_28233,N_28382);
and U28459 (N_28459,N_28308,N_28247);
and U28460 (N_28460,N_28312,N_28212);
nand U28461 (N_28461,N_28345,N_28344);
nor U28462 (N_28462,N_28289,N_28334);
nor U28463 (N_28463,N_28209,N_28252);
or U28464 (N_28464,N_28204,N_28365);
or U28465 (N_28465,N_28267,N_28323);
and U28466 (N_28466,N_28270,N_28379);
nand U28467 (N_28467,N_28232,N_28259);
nor U28468 (N_28468,N_28260,N_28337);
and U28469 (N_28469,N_28296,N_28248);
xor U28470 (N_28470,N_28376,N_28229);
or U28471 (N_28471,N_28385,N_28392);
and U28472 (N_28472,N_28202,N_28306);
and U28473 (N_28473,N_28266,N_28290);
xnor U28474 (N_28474,N_28391,N_28346);
and U28475 (N_28475,N_28207,N_28342);
nand U28476 (N_28476,N_28319,N_28363);
or U28477 (N_28477,N_28397,N_28273);
nor U28478 (N_28478,N_28242,N_28225);
nor U28479 (N_28479,N_28317,N_28322);
nand U28480 (N_28480,N_28369,N_28370);
nor U28481 (N_28481,N_28284,N_28281);
or U28482 (N_28482,N_28381,N_28249);
or U28483 (N_28483,N_28326,N_28253);
xor U28484 (N_28484,N_28313,N_28286);
nor U28485 (N_28485,N_28243,N_28333);
xor U28486 (N_28486,N_28315,N_28220);
or U28487 (N_28487,N_28269,N_28352);
or U28488 (N_28488,N_28380,N_28338);
xnor U28489 (N_28489,N_28330,N_28335);
nor U28490 (N_28490,N_28374,N_28364);
nand U28491 (N_28491,N_28279,N_28257);
and U28492 (N_28492,N_28318,N_28387);
or U28493 (N_28493,N_28256,N_28291);
or U28494 (N_28494,N_28377,N_28329);
and U28495 (N_28495,N_28347,N_28292);
nor U28496 (N_28496,N_28341,N_28276);
nor U28497 (N_28497,N_28357,N_28297);
nand U28498 (N_28498,N_28258,N_28235);
and U28499 (N_28499,N_28216,N_28245);
or U28500 (N_28500,N_28368,N_28380);
xnor U28501 (N_28501,N_28305,N_28331);
or U28502 (N_28502,N_28251,N_28327);
nand U28503 (N_28503,N_28235,N_28257);
nand U28504 (N_28504,N_28269,N_28243);
or U28505 (N_28505,N_28270,N_28223);
or U28506 (N_28506,N_28288,N_28290);
or U28507 (N_28507,N_28321,N_28275);
nand U28508 (N_28508,N_28288,N_28295);
or U28509 (N_28509,N_28399,N_28365);
or U28510 (N_28510,N_28215,N_28336);
and U28511 (N_28511,N_28357,N_28235);
or U28512 (N_28512,N_28269,N_28383);
and U28513 (N_28513,N_28388,N_28306);
xor U28514 (N_28514,N_28328,N_28215);
nor U28515 (N_28515,N_28273,N_28266);
nor U28516 (N_28516,N_28344,N_28376);
and U28517 (N_28517,N_28219,N_28380);
and U28518 (N_28518,N_28380,N_28320);
xnor U28519 (N_28519,N_28216,N_28370);
nand U28520 (N_28520,N_28294,N_28338);
or U28521 (N_28521,N_28280,N_28265);
nor U28522 (N_28522,N_28235,N_28308);
nor U28523 (N_28523,N_28325,N_28396);
nand U28524 (N_28524,N_28347,N_28238);
nand U28525 (N_28525,N_28378,N_28272);
nand U28526 (N_28526,N_28293,N_28363);
xor U28527 (N_28527,N_28268,N_28214);
nor U28528 (N_28528,N_28368,N_28385);
or U28529 (N_28529,N_28318,N_28393);
xnor U28530 (N_28530,N_28272,N_28217);
nand U28531 (N_28531,N_28351,N_28272);
nor U28532 (N_28532,N_28258,N_28295);
nor U28533 (N_28533,N_28294,N_28323);
nand U28534 (N_28534,N_28390,N_28277);
nor U28535 (N_28535,N_28354,N_28323);
nand U28536 (N_28536,N_28212,N_28396);
xnor U28537 (N_28537,N_28370,N_28209);
or U28538 (N_28538,N_28345,N_28330);
nor U28539 (N_28539,N_28366,N_28370);
and U28540 (N_28540,N_28347,N_28297);
xnor U28541 (N_28541,N_28207,N_28352);
and U28542 (N_28542,N_28294,N_28370);
and U28543 (N_28543,N_28398,N_28260);
or U28544 (N_28544,N_28369,N_28264);
nand U28545 (N_28545,N_28349,N_28376);
and U28546 (N_28546,N_28241,N_28293);
nand U28547 (N_28547,N_28242,N_28265);
nor U28548 (N_28548,N_28221,N_28308);
xor U28549 (N_28549,N_28228,N_28390);
nand U28550 (N_28550,N_28378,N_28232);
and U28551 (N_28551,N_28333,N_28369);
nor U28552 (N_28552,N_28202,N_28293);
nand U28553 (N_28553,N_28280,N_28382);
xor U28554 (N_28554,N_28375,N_28315);
and U28555 (N_28555,N_28249,N_28241);
nor U28556 (N_28556,N_28395,N_28213);
and U28557 (N_28557,N_28389,N_28359);
nor U28558 (N_28558,N_28220,N_28333);
nor U28559 (N_28559,N_28318,N_28288);
and U28560 (N_28560,N_28390,N_28350);
or U28561 (N_28561,N_28249,N_28328);
nor U28562 (N_28562,N_28307,N_28324);
xor U28563 (N_28563,N_28316,N_28324);
or U28564 (N_28564,N_28368,N_28322);
nand U28565 (N_28565,N_28317,N_28210);
xor U28566 (N_28566,N_28361,N_28234);
nand U28567 (N_28567,N_28313,N_28341);
nand U28568 (N_28568,N_28311,N_28278);
nand U28569 (N_28569,N_28246,N_28389);
or U28570 (N_28570,N_28391,N_28300);
nand U28571 (N_28571,N_28249,N_28281);
nand U28572 (N_28572,N_28288,N_28226);
and U28573 (N_28573,N_28270,N_28229);
and U28574 (N_28574,N_28222,N_28202);
nand U28575 (N_28575,N_28247,N_28317);
and U28576 (N_28576,N_28391,N_28393);
nand U28577 (N_28577,N_28248,N_28311);
nand U28578 (N_28578,N_28390,N_28355);
and U28579 (N_28579,N_28338,N_28322);
xnor U28580 (N_28580,N_28240,N_28302);
nand U28581 (N_28581,N_28338,N_28397);
xor U28582 (N_28582,N_28315,N_28365);
nand U28583 (N_28583,N_28257,N_28337);
nor U28584 (N_28584,N_28240,N_28276);
xnor U28585 (N_28585,N_28389,N_28214);
and U28586 (N_28586,N_28227,N_28266);
and U28587 (N_28587,N_28248,N_28234);
nor U28588 (N_28588,N_28377,N_28365);
nor U28589 (N_28589,N_28327,N_28277);
xnor U28590 (N_28590,N_28309,N_28366);
or U28591 (N_28591,N_28280,N_28287);
nor U28592 (N_28592,N_28301,N_28330);
nand U28593 (N_28593,N_28356,N_28329);
and U28594 (N_28594,N_28243,N_28257);
and U28595 (N_28595,N_28228,N_28371);
and U28596 (N_28596,N_28203,N_28221);
and U28597 (N_28597,N_28242,N_28237);
or U28598 (N_28598,N_28258,N_28276);
and U28599 (N_28599,N_28240,N_28263);
nor U28600 (N_28600,N_28494,N_28422);
xor U28601 (N_28601,N_28534,N_28499);
and U28602 (N_28602,N_28408,N_28536);
or U28603 (N_28603,N_28511,N_28519);
xor U28604 (N_28604,N_28532,N_28509);
and U28605 (N_28605,N_28415,N_28501);
or U28606 (N_28606,N_28571,N_28587);
and U28607 (N_28607,N_28419,N_28555);
or U28608 (N_28608,N_28473,N_28487);
and U28609 (N_28609,N_28469,N_28481);
and U28610 (N_28610,N_28505,N_28569);
nor U28611 (N_28611,N_28504,N_28517);
nor U28612 (N_28612,N_28521,N_28586);
nand U28613 (N_28613,N_28438,N_28593);
nor U28614 (N_28614,N_28440,N_28576);
and U28615 (N_28615,N_28441,N_28558);
xnor U28616 (N_28616,N_28550,N_28560);
nor U28617 (N_28617,N_28414,N_28489);
nor U28618 (N_28618,N_28453,N_28407);
nand U28619 (N_28619,N_28500,N_28512);
and U28620 (N_28620,N_28426,N_28518);
nand U28621 (N_28621,N_28424,N_28470);
xnor U28622 (N_28622,N_28435,N_28527);
nand U28623 (N_28623,N_28471,N_28412);
or U28624 (N_28624,N_28482,N_28540);
xnor U28625 (N_28625,N_28483,N_28556);
or U28626 (N_28626,N_28572,N_28480);
and U28627 (N_28627,N_28561,N_28516);
nand U28628 (N_28628,N_28584,N_28545);
or U28629 (N_28629,N_28403,N_28522);
nor U28630 (N_28630,N_28462,N_28485);
xor U28631 (N_28631,N_28493,N_28530);
or U28632 (N_28632,N_28590,N_28537);
xor U28633 (N_28633,N_28484,N_28428);
nand U28634 (N_28634,N_28458,N_28570);
xor U28635 (N_28635,N_28463,N_28541);
and U28636 (N_28636,N_28496,N_28478);
nor U28637 (N_28637,N_28575,N_28594);
nand U28638 (N_28638,N_28579,N_28507);
nand U28639 (N_28639,N_28433,N_28448);
or U28640 (N_28640,N_28531,N_28554);
and U28641 (N_28641,N_28502,N_28529);
nand U28642 (N_28642,N_28539,N_28479);
nor U28643 (N_28643,N_28523,N_28420);
or U28644 (N_28644,N_28423,N_28520);
nor U28645 (N_28645,N_28559,N_28400);
nor U28646 (N_28646,N_28526,N_28595);
or U28647 (N_28647,N_28533,N_28552);
nor U28648 (N_28648,N_28513,N_28429);
and U28649 (N_28649,N_28446,N_28465);
nor U28650 (N_28650,N_28491,N_28430);
nand U28651 (N_28651,N_28551,N_28583);
nor U28652 (N_28652,N_28592,N_28460);
nand U28653 (N_28653,N_28436,N_28442);
nor U28654 (N_28654,N_28425,N_28409);
and U28655 (N_28655,N_28542,N_28454);
or U28656 (N_28656,N_28475,N_28417);
nor U28657 (N_28657,N_28450,N_28524);
nor U28658 (N_28658,N_28573,N_28401);
xnor U28659 (N_28659,N_28466,N_28596);
or U28660 (N_28660,N_28538,N_28567);
or U28661 (N_28661,N_28416,N_28447);
xor U28662 (N_28662,N_28457,N_28445);
nand U28663 (N_28663,N_28566,N_28563);
nor U28664 (N_28664,N_28599,N_28546);
nor U28665 (N_28665,N_28411,N_28410);
xor U28666 (N_28666,N_28580,N_28515);
xor U28667 (N_28667,N_28508,N_28451);
and U28668 (N_28668,N_28459,N_28421);
nor U28669 (N_28669,N_28553,N_28486);
or U28670 (N_28670,N_28468,N_28449);
xnor U28671 (N_28671,N_28405,N_28413);
xor U28672 (N_28672,N_28577,N_28439);
nor U28673 (N_28673,N_28581,N_28443);
and U28674 (N_28674,N_28565,N_28589);
xor U28675 (N_28675,N_28427,N_28503);
xnor U28676 (N_28676,N_28452,N_28568);
and U28677 (N_28677,N_28456,N_28598);
nor U28678 (N_28678,N_28514,N_28544);
nand U28679 (N_28679,N_28472,N_28418);
and U28680 (N_28680,N_28464,N_28431);
or U28681 (N_28681,N_28591,N_28476);
nand U28682 (N_28682,N_28547,N_28497);
xnor U28683 (N_28683,N_28455,N_28528);
nor U28684 (N_28684,N_28548,N_28495);
xnor U28685 (N_28685,N_28488,N_28510);
and U28686 (N_28686,N_28525,N_28588);
and U28687 (N_28687,N_28474,N_28506);
nor U28688 (N_28688,N_28597,N_28535);
xnor U28689 (N_28689,N_28406,N_28432);
nor U28690 (N_28690,N_28543,N_28549);
nand U28691 (N_28691,N_28404,N_28562);
nand U28692 (N_28692,N_28467,N_28564);
nand U28693 (N_28693,N_28492,N_28434);
nor U28694 (N_28694,N_28557,N_28490);
or U28695 (N_28695,N_28498,N_28578);
or U28696 (N_28696,N_28461,N_28582);
nor U28697 (N_28697,N_28574,N_28444);
xor U28698 (N_28698,N_28477,N_28402);
xnor U28699 (N_28699,N_28437,N_28585);
xor U28700 (N_28700,N_28599,N_28586);
xor U28701 (N_28701,N_28404,N_28432);
or U28702 (N_28702,N_28539,N_28444);
nand U28703 (N_28703,N_28519,N_28504);
nand U28704 (N_28704,N_28591,N_28483);
or U28705 (N_28705,N_28530,N_28584);
nand U28706 (N_28706,N_28570,N_28580);
and U28707 (N_28707,N_28496,N_28489);
nand U28708 (N_28708,N_28574,N_28484);
nor U28709 (N_28709,N_28589,N_28443);
xor U28710 (N_28710,N_28571,N_28450);
xnor U28711 (N_28711,N_28437,N_28506);
or U28712 (N_28712,N_28577,N_28512);
nand U28713 (N_28713,N_28542,N_28449);
xor U28714 (N_28714,N_28535,N_28467);
nand U28715 (N_28715,N_28589,N_28458);
and U28716 (N_28716,N_28502,N_28517);
nor U28717 (N_28717,N_28546,N_28527);
or U28718 (N_28718,N_28581,N_28402);
nand U28719 (N_28719,N_28440,N_28417);
nor U28720 (N_28720,N_28456,N_28542);
and U28721 (N_28721,N_28485,N_28534);
and U28722 (N_28722,N_28549,N_28474);
nand U28723 (N_28723,N_28536,N_28473);
and U28724 (N_28724,N_28512,N_28523);
xor U28725 (N_28725,N_28446,N_28438);
and U28726 (N_28726,N_28421,N_28433);
xor U28727 (N_28727,N_28580,N_28555);
nor U28728 (N_28728,N_28462,N_28407);
and U28729 (N_28729,N_28527,N_28544);
nor U28730 (N_28730,N_28520,N_28546);
and U28731 (N_28731,N_28463,N_28530);
xor U28732 (N_28732,N_28595,N_28400);
or U28733 (N_28733,N_28413,N_28451);
nand U28734 (N_28734,N_28566,N_28592);
nand U28735 (N_28735,N_28515,N_28549);
or U28736 (N_28736,N_28533,N_28515);
nor U28737 (N_28737,N_28531,N_28523);
xor U28738 (N_28738,N_28441,N_28411);
nand U28739 (N_28739,N_28510,N_28505);
or U28740 (N_28740,N_28459,N_28492);
xor U28741 (N_28741,N_28446,N_28570);
or U28742 (N_28742,N_28511,N_28434);
or U28743 (N_28743,N_28520,N_28412);
or U28744 (N_28744,N_28558,N_28578);
nor U28745 (N_28745,N_28487,N_28403);
or U28746 (N_28746,N_28424,N_28526);
xor U28747 (N_28747,N_28475,N_28551);
xor U28748 (N_28748,N_28484,N_28579);
xor U28749 (N_28749,N_28524,N_28414);
or U28750 (N_28750,N_28462,N_28591);
xor U28751 (N_28751,N_28448,N_28510);
xor U28752 (N_28752,N_28460,N_28403);
nand U28753 (N_28753,N_28460,N_28586);
and U28754 (N_28754,N_28557,N_28565);
nand U28755 (N_28755,N_28548,N_28598);
and U28756 (N_28756,N_28417,N_28429);
nand U28757 (N_28757,N_28480,N_28448);
nand U28758 (N_28758,N_28497,N_28487);
nor U28759 (N_28759,N_28468,N_28541);
nor U28760 (N_28760,N_28531,N_28430);
or U28761 (N_28761,N_28454,N_28420);
nor U28762 (N_28762,N_28502,N_28443);
xnor U28763 (N_28763,N_28472,N_28572);
and U28764 (N_28764,N_28548,N_28462);
nor U28765 (N_28765,N_28430,N_28496);
nand U28766 (N_28766,N_28583,N_28567);
nand U28767 (N_28767,N_28428,N_28456);
xnor U28768 (N_28768,N_28406,N_28460);
xor U28769 (N_28769,N_28554,N_28468);
xnor U28770 (N_28770,N_28474,N_28490);
nor U28771 (N_28771,N_28483,N_28575);
xor U28772 (N_28772,N_28548,N_28529);
nor U28773 (N_28773,N_28572,N_28456);
xor U28774 (N_28774,N_28495,N_28564);
nor U28775 (N_28775,N_28423,N_28575);
or U28776 (N_28776,N_28451,N_28421);
or U28777 (N_28777,N_28577,N_28573);
xor U28778 (N_28778,N_28512,N_28548);
nand U28779 (N_28779,N_28513,N_28416);
or U28780 (N_28780,N_28470,N_28451);
nor U28781 (N_28781,N_28403,N_28582);
xor U28782 (N_28782,N_28499,N_28572);
or U28783 (N_28783,N_28425,N_28520);
nand U28784 (N_28784,N_28553,N_28471);
nand U28785 (N_28785,N_28462,N_28541);
nand U28786 (N_28786,N_28542,N_28525);
nand U28787 (N_28787,N_28413,N_28411);
or U28788 (N_28788,N_28597,N_28432);
nand U28789 (N_28789,N_28557,N_28432);
and U28790 (N_28790,N_28452,N_28483);
xor U28791 (N_28791,N_28439,N_28581);
xnor U28792 (N_28792,N_28548,N_28599);
nand U28793 (N_28793,N_28495,N_28439);
nor U28794 (N_28794,N_28437,N_28582);
and U28795 (N_28795,N_28597,N_28416);
or U28796 (N_28796,N_28565,N_28522);
nor U28797 (N_28797,N_28594,N_28431);
nor U28798 (N_28798,N_28540,N_28435);
xor U28799 (N_28799,N_28538,N_28466);
xnor U28800 (N_28800,N_28639,N_28733);
xnor U28801 (N_28801,N_28748,N_28796);
or U28802 (N_28802,N_28688,N_28722);
or U28803 (N_28803,N_28661,N_28783);
nand U28804 (N_28804,N_28678,N_28792);
nor U28805 (N_28805,N_28721,N_28705);
nor U28806 (N_28806,N_28777,N_28602);
nor U28807 (N_28807,N_28667,N_28647);
nand U28808 (N_28808,N_28773,N_28669);
or U28809 (N_28809,N_28666,N_28630);
nor U28810 (N_28810,N_28640,N_28717);
and U28811 (N_28811,N_28702,N_28761);
and U28812 (N_28812,N_28635,N_28648);
nand U28813 (N_28813,N_28716,N_28742);
nor U28814 (N_28814,N_28618,N_28634);
and U28815 (N_28815,N_28739,N_28627);
nand U28816 (N_28816,N_28660,N_28760);
nand U28817 (N_28817,N_28798,N_28664);
nor U28818 (N_28818,N_28654,N_28747);
nand U28819 (N_28819,N_28726,N_28613);
xnor U28820 (N_28820,N_28746,N_28711);
xor U28821 (N_28821,N_28692,N_28782);
or U28822 (N_28822,N_28632,N_28644);
or U28823 (N_28823,N_28779,N_28780);
nor U28824 (N_28824,N_28764,N_28767);
or U28825 (N_28825,N_28681,N_28745);
nand U28826 (N_28826,N_28741,N_28772);
nor U28827 (N_28827,N_28759,N_28673);
xor U28828 (N_28828,N_28663,N_28700);
xor U28829 (N_28829,N_28677,N_28616);
and U28830 (N_28830,N_28710,N_28658);
nand U28831 (N_28831,N_28794,N_28607);
and U28832 (N_28832,N_28625,N_28642);
or U28833 (N_28833,N_28615,N_28775);
or U28834 (N_28834,N_28671,N_28696);
xor U28835 (N_28835,N_28638,N_28708);
nor U28836 (N_28836,N_28699,N_28765);
nor U28837 (N_28837,N_28672,N_28799);
nand U28838 (N_28838,N_28628,N_28651);
nor U28839 (N_28839,N_28762,N_28734);
or U28840 (N_28840,N_28737,N_28797);
nor U28841 (N_28841,N_28679,N_28729);
nand U28842 (N_28842,N_28771,N_28675);
nand U28843 (N_28843,N_28793,N_28788);
xor U28844 (N_28844,N_28695,N_28606);
or U28845 (N_28845,N_28624,N_28724);
or U28846 (N_28846,N_28609,N_28735);
xnor U28847 (N_28847,N_28684,N_28753);
and U28848 (N_28848,N_28685,N_28603);
nand U28849 (N_28849,N_28789,N_28730);
nor U28850 (N_28850,N_28655,N_28689);
and U28851 (N_28851,N_28752,N_28707);
nand U28852 (N_28852,N_28633,N_28645);
xor U28853 (N_28853,N_28662,N_28680);
xor U28854 (N_28854,N_28687,N_28786);
nor U28855 (N_28855,N_28768,N_28693);
nand U28856 (N_28856,N_28715,N_28690);
nand U28857 (N_28857,N_28795,N_28646);
nor U28858 (N_28858,N_28659,N_28732);
xor U28859 (N_28859,N_28698,N_28723);
and U28860 (N_28860,N_28727,N_28620);
nor U28861 (N_28861,N_28763,N_28653);
or U28862 (N_28862,N_28712,N_28751);
nand U28863 (N_28863,N_28749,N_28714);
xor U28864 (N_28864,N_28750,N_28718);
and U28865 (N_28865,N_28637,N_28604);
nor U28866 (N_28866,N_28622,N_28614);
and U28867 (N_28867,N_28756,N_28778);
nor U28868 (N_28868,N_28691,N_28757);
or U28869 (N_28869,N_28719,N_28611);
or U28870 (N_28870,N_28736,N_28641);
or U28871 (N_28871,N_28787,N_28713);
or U28872 (N_28872,N_28725,N_28623);
xor U28873 (N_28873,N_28758,N_28670);
and U28874 (N_28874,N_28709,N_28649);
nor U28875 (N_28875,N_28643,N_28697);
nand U28876 (N_28876,N_28770,N_28605);
nor U28877 (N_28877,N_28781,N_28683);
nor U28878 (N_28878,N_28704,N_28600);
nor U28879 (N_28879,N_28650,N_28612);
nand U28880 (N_28880,N_28686,N_28743);
nand U28881 (N_28881,N_28728,N_28682);
and U28882 (N_28882,N_28608,N_28766);
nor U28883 (N_28883,N_28652,N_28610);
nor U28884 (N_28884,N_28631,N_28731);
nor U28885 (N_28885,N_28674,N_28626);
and U28886 (N_28886,N_28694,N_28740);
nand U28887 (N_28887,N_28657,N_28720);
or U28888 (N_28888,N_28703,N_28665);
nor U28889 (N_28889,N_28619,N_28701);
nand U28890 (N_28890,N_28769,N_28656);
and U28891 (N_28891,N_28668,N_28636);
and U28892 (N_28892,N_28790,N_28738);
and U28893 (N_28893,N_28785,N_28676);
xor U28894 (N_28894,N_28776,N_28755);
or U28895 (N_28895,N_28754,N_28791);
or U28896 (N_28896,N_28706,N_28617);
nand U28897 (N_28897,N_28629,N_28744);
and U28898 (N_28898,N_28621,N_28601);
nand U28899 (N_28899,N_28774,N_28784);
xor U28900 (N_28900,N_28700,N_28758);
or U28901 (N_28901,N_28606,N_28776);
xnor U28902 (N_28902,N_28646,N_28749);
or U28903 (N_28903,N_28613,N_28760);
or U28904 (N_28904,N_28775,N_28686);
xor U28905 (N_28905,N_28783,N_28738);
or U28906 (N_28906,N_28786,N_28611);
or U28907 (N_28907,N_28771,N_28679);
xnor U28908 (N_28908,N_28778,N_28743);
or U28909 (N_28909,N_28730,N_28718);
and U28910 (N_28910,N_28700,N_28798);
nor U28911 (N_28911,N_28730,N_28736);
or U28912 (N_28912,N_28673,N_28787);
nor U28913 (N_28913,N_28655,N_28634);
xnor U28914 (N_28914,N_28725,N_28629);
or U28915 (N_28915,N_28702,N_28686);
nor U28916 (N_28916,N_28603,N_28699);
or U28917 (N_28917,N_28626,N_28648);
and U28918 (N_28918,N_28712,N_28687);
and U28919 (N_28919,N_28685,N_28690);
or U28920 (N_28920,N_28664,N_28768);
or U28921 (N_28921,N_28765,N_28608);
or U28922 (N_28922,N_28682,N_28647);
or U28923 (N_28923,N_28769,N_28786);
nor U28924 (N_28924,N_28778,N_28738);
and U28925 (N_28925,N_28755,N_28605);
nor U28926 (N_28926,N_28700,N_28797);
or U28927 (N_28927,N_28698,N_28612);
nor U28928 (N_28928,N_28635,N_28783);
and U28929 (N_28929,N_28739,N_28675);
and U28930 (N_28930,N_28757,N_28783);
or U28931 (N_28931,N_28798,N_28753);
or U28932 (N_28932,N_28749,N_28764);
xor U28933 (N_28933,N_28756,N_28678);
or U28934 (N_28934,N_28653,N_28766);
or U28935 (N_28935,N_28718,N_28639);
nand U28936 (N_28936,N_28772,N_28783);
nor U28937 (N_28937,N_28640,N_28684);
and U28938 (N_28938,N_28727,N_28687);
xnor U28939 (N_28939,N_28796,N_28775);
xor U28940 (N_28940,N_28681,N_28628);
nor U28941 (N_28941,N_28776,N_28662);
and U28942 (N_28942,N_28797,N_28655);
or U28943 (N_28943,N_28666,N_28690);
and U28944 (N_28944,N_28691,N_28694);
or U28945 (N_28945,N_28651,N_28779);
nor U28946 (N_28946,N_28784,N_28744);
nand U28947 (N_28947,N_28763,N_28666);
xor U28948 (N_28948,N_28770,N_28757);
and U28949 (N_28949,N_28648,N_28602);
xor U28950 (N_28950,N_28612,N_28735);
or U28951 (N_28951,N_28781,N_28652);
or U28952 (N_28952,N_28603,N_28684);
nand U28953 (N_28953,N_28787,N_28684);
or U28954 (N_28954,N_28765,N_28633);
xnor U28955 (N_28955,N_28625,N_28671);
nor U28956 (N_28956,N_28723,N_28626);
or U28957 (N_28957,N_28771,N_28637);
xnor U28958 (N_28958,N_28639,N_28735);
or U28959 (N_28959,N_28696,N_28771);
xnor U28960 (N_28960,N_28768,N_28699);
nor U28961 (N_28961,N_28781,N_28688);
nor U28962 (N_28962,N_28756,N_28640);
nor U28963 (N_28963,N_28617,N_28631);
or U28964 (N_28964,N_28605,N_28660);
and U28965 (N_28965,N_28674,N_28662);
nand U28966 (N_28966,N_28714,N_28765);
nor U28967 (N_28967,N_28617,N_28760);
or U28968 (N_28968,N_28655,N_28660);
or U28969 (N_28969,N_28624,N_28606);
and U28970 (N_28970,N_28793,N_28658);
xnor U28971 (N_28971,N_28647,N_28733);
and U28972 (N_28972,N_28710,N_28623);
or U28973 (N_28973,N_28684,N_28699);
xor U28974 (N_28974,N_28647,N_28701);
nor U28975 (N_28975,N_28724,N_28606);
or U28976 (N_28976,N_28796,N_28692);
nor U28977 (N_28977,N_28684,N_28657);
and U28978 (N_28978,N_28709,N_28625);
xor U28979 (N_28979,N_28766,N_28691);
xor U28980 (N_28980,N_28693,N_28646);
or U28981 (N_28981,N_28635,N_28662);
nand U28982 (N_28982,N_28770,N_28696);
xor U28983 (N_28983,N_28730,N_28720);
nand U28984 (N_28984,N_28794,N_28604);
xnor U28985 (N_28985,N_28650,N_28611);
or U28986 (N_28986,N_28734,N_28760);
nand U28987 (N_28987,N_28657,N_28744);
nand U28988 (N_28988,N_28657,N_28690);
nor U28989 (N_28989,N_28666,N_28733);
nor U28990 (N_28990,N_28769,N_28717);
and U28991 (N_28991,N_28688,N_28626);
xor U28992 (N_28992,N_28707,N_28672);
and U28993 (N_28993,N_28713,N_28648);
nand U28994 (N_28994,N_28663,N_28743);
or U28995 (N_28995,N_28650,N_28778);
xnor U28996 (N_28996,N_28632,N_28627);
or U28997 (N_28997,N_28731,N_28611);
and U28998 (N_28998,N_28675,N_28622);
xor U28999 (N_28999,N_28727,N_28696);
or U29000 (N_29000,N_28867,N_28977);
nand U29001 (N_29001,N_28907,N_28935);
nor U29002 (N_29002,N_28944,N_28850);
and U29003 (N_29003,N_28818,N_28961);
xnor U29004 (N_29004,N_28942,N_28816);
and U29005 (N_29005,N_28830,N_28819);
and U29006 (N_29006,N_28888,N_28894);
nor U29007 (N_29007,N_28988,N_28910);
nor U29008 (N_29008,N_28955,N_28918);
or U29009 (N_29009,N_28842,N_28854);
nor U29010 (N_29010,N_28897,N_28925);
or U29011 (N_29011,N_28875,N_28948);
nand U29012 (N_29012,N_28951,N_28962);
nor U29013 (N_29013,N_28880,N_28828);
xnor U29014 (N_29014,N_28864,N_28860);
nor U29015 (N_29015,N_28932,N_28914);
xnor U29016 (N_29016,N_28998,N_28803);
xor U29017 (N_29017,N_28990,N_28909);
xor U29018 (N_29018,N_28874,N_28808);
nor U29019 (N_29019,N_28811,N_28931);
nor U29020 (N_29020,N_28855,N_28911);
and U29021 (N_29021,N_28889,N_28916);
nor U29022 (N_29022,N_28841,N_28891);
or U29023 (N_29023,N_28883,N_28934);
and U29024 (N_29024,N_28893,N_28873);
xnor U29025 (N_29025,N_28901,N_28817);
nor U29026 (N_29026,N_28835,N_28947);
nand U29027 (N_29027,N_28913,N_28807);
or U29028 (N_29028,N_28965,N_28964);
xor U29029 (N_29029,N_28967,N_28829);
and U29030 (N_29030,N_28941,N_28877);
nand U29031 (N_29031,N_28969,N_28892);
nand U29032 (N_29032,N_28974,N_28912);
and U29033 (N_29033,N_28992,N_28972);
nor U29034 (N_29034,N_28994,N_28823);
xnor U29035 (N_29035,N_28986,N_28997);
and U29036 (N_29036,N_28959,N_28921);
nor U29037 (N_29037,N_28956,N_28895);
nand U29038 (N_29038,N_28866,N_28989);
nand U29039 (N_29039,N_28939,N_28834);
nand U29040 (N_29040,N_28851,N_28971);
or U29041 (N_29041,N_28946,N_28810);
nor U29042 (N_29042,N_28805,N_28973);
xor U29043 (N_29043,N_28831,N_28954);
nor U29044 (N_29044,N_28976,N_28832);
nor U29045 (N_29045,N_28905,N_28885);
nor U29046 (N_29046,N_28814,N_28843);
nand U29047 (N_29047,N_28825,N_28923);
and U29048 (N_29048,N_28887,N_28837);
nand U29049 (N_29049,N_28982,N_28898);
nand U29050 (N_29050,N_28822,N_28848);
nor U29051 (N_29051,N_28862,N_28900);
nor U29052 (N_29052,N_28804,N_28847);
nand U29053 (N_29053,N_28827,N_28852);
or U29054 (N_29054,N_28917,N_28865);
xnor U29055 (N_29055,N_28940,N_28919);
nor U29056 (N_29056,N_28991,N_28869);
xnor U29057 (N_29057,N_28927,N_28958);
and U29058 (N_29058,N_28800,N_28966);
nand U29059 (N_29059,N_28870,N_28987);
xor U29060 (N_29060,N_28908,N_28936);
and U29061 (N_29061,N_28809,N_28920);
xor U29062 (N_29062,N_28981,N_28815);
xnor U29063 (N_29063,N_28938,N_28943);
nor U29064 (N_29064,N_28863,N_28963);
and U29065 (N_29065,N_28821,N_28980);
nand U29066 (N_29066,N_28957,N_28933);
nor U29067 (N_29067,N_28878,N_28806);
xnor U29068 (N_29068,N_28882,N_28824);
nor U29069 (N_29069,N_28995,N_28950);
xor U29070 (N_29070,N_28970,N_28858);
nor U29071 (N_29071,N_28928,N_28833);
and U29072 (N_29072,N_28838,N_28846);
nor U29073 (N_29073,N_28881,N_28984);
nand U29074 (N_29074,N_28924,N_28999);
xor U29075 (N_29075,N_28953,N_28813);
or U29076 (N_29076,N_28826,N_28945);
nand U29077 (N_29077,N_28879,N_28996);
xor U29078 (N_29078,N_28906,N_28968);
or U29079 (N_29079,N_28949,N_28861);
or U29080 (N_29080,N_28904,N_28836);
xor U29081 (N_29081,N_28840,N_28978);
nor U29082 (N_29082,N_28845,N_28929);
and U29083 (N_29083,N_28876,N_28979);
or U29084 (N_29084,N_28926,N_28985);
xor U29085 (N_29085,N_28856,N_28915);
nor U29086 (N_29086,N_28853,N_28820);
nor U29087 (N_29087,N_28849,N_28952);
and U29088 (N_29088,N_28839,N_28903);
nand U29089 (N_29089,N_28922,N_28857);
and U29090 (N_29090,N_28802,N_28993);
nand U29091 (N_29091,N_28983,N_28812);
and U29092 (N_29092,N_28902,N_28896);
and U29093 (N_29093,N_28844,N_28899);
and U29094 (N_29094,N_28871,N_28868);
or U29095 (N_29095,N_28886,N_28975);
nor U29096 (N_29096,N_28884,N_28960);
and U29097 (N_29097,N_28859,N_28872);
nor U29098 (N_29098,N_28937,N_28930);
xnor U29099 (N_29099,N_28890,N_28801);
nor U29100 (N_29100,N_28809,N_28971);
nor U29101 (N_29101,N_28846,N_28921);
and U29102 (N_29102,N_28972,N_28851);
nor U29103 (N_29103,N_28868,N_28811);
or U29104 (N_29104,N_28845,N_28874);
xnor U29105 (N_29105,N_28905,N_28866);
nor U29106 (N_29106,N_28900,N_28850);
or U29107 (N_29107,N_28851,N_28850);
nor U29108 (N_29108,N_28839,N_28847);
or U29109 (N_29109,N_28942,N_28908);
nor U29110 (N_29110,N_28974,N_28858);
nand U29111 (N_29111,N_28898,N_28834);
or U29112 (N_29112,N_28906,N_28853);
nand U29113 (N_29113,N_28977,N_28931);
xnor U29114 (N_29114,N_28878,N_28999);
or U29115 (N_29115,N_28816,N_28960);
nand U29116 (N_29116,N_28807,N_28819);
xnor U29117 (N_29117,N_28880,N_28931);
xor U29118 (N_29118,N_28913,N_28820);
and U29119 (N_29119,N_28878,N_28861);
or U29120 (N_29120,N_28815,N_28952);
xnor U29121 (N_29121,N_28867,N_28858);
nand U29122 (N_29122,N_28919,N_28845);
nor U29123 (N_29123,N_28987,N_28990);
nand U29124 (N_29124,N_28993,N_28967);
nand U29125 (N_29125,N_28847,N_28939);
xor U29126 (N_29126,N_28954,N_28984);
nand U29127 (N_29127,N_28827,N_28909);
nor U29128 (N_29128,N_28888,N_28877);
or U29129 (N_29129,N_28825,N_28856);
or U29130 (N_29130,N_28959,N_28825);
nand U29131 (N_29131,N_28868,N_28952);
or U29132 (N_29132,N_28975,N_28829);
nand U29133 (N_29133,N_28823,N_28855);
xor U29134 (N_29134,N_28971,N_28995);
or U29135 (N_29135,N_28981,N_28948);
nand U29136 (N_29136,N_28914,N_28998);
xor U29137 (N_29137,N_28841,N_28905);
nand U29138 (N_29138,N_28814,N_28818);
nand U29139 (N_29139,N_28893,N_28946);
or U29140 (N_29140,N_28989,N_28806);
nand U29141 (N_29141,N_28805,N_28856);
xnor U29142 (N_29142,N_28946,N_28947);
xnor U29143 (N_29143,N_28917,N_28862);
nand U29144 (N_29144,N_28803,N_28850);
or U29145 (N_29145,N_28863,N_28937);
or U29146 (N_29146,N_28966,N_28929);
nor U29147 (N_29147,N_28813,N_28943);
or U29148 (N_29148,N_28892,N_28851);
or U29149 (N_29149,N_28938,N_28874);
xnor U29150 (N_29150,N_28911,N_28848);
nor U29151 (N_29151,N_28972,N_28849);
and U29152 (N_29152,N_28942,N_28841);
xor U29153 (N_29153,N_28877,N_28828);
and U29154 (N_29154,N_28866,N_28844);
and U29155 (N_29155,N_28900,N_28914);
nand U29156 (N_29156,N_28956,N_28946);
nand U29157 (N_29157,N_28987,N_28838);
nand U29158 (N_29158,N_28999,N_28982);
and U29159 (N_29159,N_28889,N_28802);
nor U29160 (N_29160,N_28829,N_28885);
and U29161 (N_29161,N_28828,N_28897);
xor U29162 (N_29162,N_28951,N_28881);
or U29163 (N_29163,N_28864,N_28926);
nor U29164 (N_29164,N_28965,N_28949);
nor U29165 (N_29165,N_28870,N_28849);
and U29166 (N_29166,N_28871,N_28900);
xnor U29167 (N_29167,N_28800,N_28801);
nor U29168 (N_29168,N_28822,N_28827);
nor U29169 (N_29169,N_28995,N_28867);
nor U29170 (N_29170,N_28970,N_28953);
and U29171 (N_29171,N_28802,N_28886);
and U29172 (N_29172,N_28985,N_28959);
nand U29173 (N_29173,N_28829,N_28815);
and U29174 (N_29174,N_28998,N_28820);
or U29175 (N_29175,N_28966,N_28965);
nor U29176 (N_29176,N_28851,N_28939);
and U29177 (N_29177,N_28978,N_28970);
xor U29178 (N_29178,N_28898,N_28967);
and U29179 (N_29179,N_28811,N_28841);
and U29180 (N_29180,N_28852,N_28930);
nand U29181 (N_29181,N_28924,N_28913);
and U29182 (N_29182,N_28998,N_28829);
xor U29183 (N_29183,N_28963,N_28962);
and U29184 (N_29184,N_28918,N_28911);
or U29185 (N_29185,N_28818,N_28962);
nor U29186 (N_29186,N_28831,N_28985);
or U29187 (N_29187,N_28864,N_28801);
and U29188 (N_29188,N_28830,N_28906);
nand U29189 (N_29189,N_28858,N_28942);
nor U29190 (N_29190,N_28823,N_28979);
nand U29191 (N_29191,N_28930,N_28847);
xnor U29192 (N_29192,N_28991,N_28875);
xnor U29193 (N_29193,N_28911,N_28938);
xnor U29194 (N_29194,N_28886,N_28835);
or U29195 (N_29195,N_28827,N_28987);
xnor U29196 (N_29196,N_28815,N_28902);
and U29197 (N_29197,N_28917,N_28989);
and U29198 (N_29198,N_28840,N_28939);
or U29199 (N_29199,N_28847,N_28991);
and U29200 (N_29200,N_29061,N_29036);
or U29201 (N_29201,N_29006,N_29051);
and U29202 (N_29202,N_29059,N_29044);
nand U29203 (N_29203,N_29030,N_29152);
xnor U29204 (N_29204,N_29147,N_29180);
nor U29205 (N_29205,N_29186,N_29129);
nor U29206 (N_29206,N_29192,N_29089);
or U29207 (N_29207,N_29118,N_29169);
or U29208 (N_29208,N_29060,N_29076);
or U29209 (N_29209,N_29151,N_29143);
nand U29210 (N_29210,N_29097,N_29033);
nand U29211 (N_29211,N_29073,N_29140);
xor U29212 (N_29212,N_29177,N_29032);
xor U29213 (N_29213,N_29092,N_29122);
or U29214 (N_29214,N_29047,N_29190);
and U29215 (N_29215,N_29173,N_29009);
and U29216 (N_29216,N_29138,N_29017);
and U29217 (N_29217,N_29175,N_29109);
and U29218 (N_29218,N_29154,N_29081);
nor U29219 (N_29219,N_29142,N_29132);
or U29220 (N_29220,N_29099,N_29102);
nor U29221 (N_29221,N_29071,N_29185);
nor U29222 (N_29222,N_29056,N_29095);
xnor U29223 (N_29223,N_29085,N_29016);
nand U29224 (N_29224,N_29157,N_29063);
nor U29225 (N_29225,N_29058,N_29098);
and U29226 (N_29226,N_29068,N_29183);
and U29227 (N_29227,N_29057,N_29199);
or U29228 (N_29228,N_29015,N_29176);
xnor U29229 (N_29229,N_29166,N_29079);
xnor U29230 (N_29230,N_29083,N_29027);
nor U29231 (N_29231,N_29104,N_29050);
nor U29232 (N_29232,N_29112,N_29008);
nand U29233 (N_29233,N_29086,N_29034);
and U29234 (N_29234,N_29084,N_29082);
nor U29235 (N_29235,N_29149,N_29179);
xor U29236 (N_29236,N_29123,N_29158);
xor U29237 (N_29237,N_29002,N_29054);
nand U29238 (N_29238,N_29014,N_29191);
and U29239 (N_29239,N_29029,N_29193);
xnor U29240 (N_29240,N_29119,N_29196);
nor U29241 (N_29241,N_29131,N_29135);
nand U29242 (N_29242,N_29165,N_29114);
and U29243 (N_29243,N_29062,N_29198);
and U29244 (N_29244,N_29181,N_29174);
or U29245 (N_29245,N_29133,N_29172);
nor U29246 (N_29246,N_29100,N_29020);
nor U29247 (N_29247,N_29110,N_29090);
nor U29248 (N_29248,N_29080,N_29003);
or U29249 (N_29249,N_29023,N_29025);
nand U29250 (N_29250,N_29188,N_29011);
and U29251 (N_29251,N_29024,N_29072);
and U29252 (N_29252,N_29184,N_29019);
nor U29253 (N_29253,N_29087,N_29127);
nand U29254 (N_29254,N_29012,N_29148);
and U29255 (N_29255,N_29146,N_29045);
and U29256 (N_29256,N_29004,N_29106);
or U29257 (N_29257,N_29101,N_29162);
nand U29258 (N_29258,N_29096,N_29039);
nor U29259 (N_29259,N_29111,N_29139);
or U29260 (N_29260,N_29066,N_29164);
and U29261 (N_29261,N_29121,N_29168);
xor U29262 (N_29262,N_29141,N_29150);
nor U29263 (N_29263,N_29046,N_29075);
nand U29264 (N_29264,N_29155,N_29010);
nand U29265 (N_29265,N_29128,N_29108);
and U29266 (N_29266,N_29007,N_29125);
nor U29267 (N_29267,N_29064,N_29031);
and U29268 (N_29268,N_29070,N_29153);
nor U29269 (N_29269,N_29013,N_29091);
or U29270 (N_29270,N_29117,N_29053);
and U29271 (N_29271,N_29093,N_29116);
nand U29272 (N_29272,N_29005,N_29120);
and U29273 (N_29273,N_29163,N_29040);
nor U29274 (N_29274,N_29022,N_29038);
or U29275 (N_29275,N_29094,N_29171);
and U29276 (N_29276,N_29144,N_29078);
nand U29277 (N_29277,N_29126,N_29170);
nand U29278 (N_29278,N_29069,N_29115);
and U29279 (N_29279,N_29136,N_29130);
and U29280 (N_29280,N_29065,N_29055);
or U29281 (N_29281,N_29067,N_29074);
nor U29282 (N_29282,N_29042,N_29021);
nand U29283 (N_29283,N_29088,N_29037);
and U29284 (N_29284,N_29137,N_29113);
nand U29285 (N_29285,N_29134,N_29189);
nor U29286 (N_29286,N_29161,N_29160);
nand U29287 (N_29287,N_29028,N_29182);
or U29288 (N_29288,N_29049,N_29001);
xnor U29289 (N_29289,N_29041,N_29103);
xnor U29290 (N_29290,N_29035,N_29052);
nand U29291 (N_29291,N_29178,N_29197);
xor U29292 (N_29292,N_29018,N_29187);
or U29293 (N_29293,N_29156,N_29194);
and U29294 (N_29294,N_29105,N_29195);
xnor U29295 (N_29295,N_29026,N_29167);
nand U29296 (N_29296,N_29043,N_29077);
nor U29297 (N_29297,N_29107,N_29048);
nor U29298 (N_29298,N_29145,N_29000);
nand U29299 (N_29299,N_29124,N_29159);
and U29300 (N_29300,N_29170,N_29104);
nand U29301 (N_29301,N_29025,N_29108);
and U29302 (N_29302,N_29055,N_29113);
nor U29303 (N_29303,N_29124,N_29151);
nor U29304 (N_29304,N_29001,N_29068);
or U29305 (N_29305,N_29179,N_29011);
or U29306 (N_29306,N_29193,N_29017);
or U29307 (N_29307,N_29008,N_29099);
or U29308 (N_29308,N_29033,N_29082);
nor U29309 (N_29309,N_29117,N_29138);
nor U29310 (N_29310,N_29002,N_29151);
nor U29311 (N_29311,N_29020,N_29018);
nor U29312 (N_29312,N_29067,N_29096);
nor U29313 (N_29313,N_29077,N_29135);
and U29314 (N_29314,N_29148,N_29195);
xnor U29315 (N_29315,N_29053,N_29008);
or U29316 (N_29316,N_29128,N_29156);
and U29317 (N_29317,N_29067,N_29118);
and U29318 (N_29318,N_29017,N_29042);
nor U29319 (N_29319,N_29167,N_29113);
and U29320 (N_29320,N_29027,N_29104);
nand U29321 (N_29321,N_29077,N_29191);
or U29322 (N_29322,N_29178,N_29195);
or U29323 (N_29323,N_29018,N_29147);
nor U29324 (N_29324,N_29145,N_29090);
or U29325 (N_29325,N_29032,N_29070);
xor U29326 (N_29326,N_29019,N_29055);
and U29327 (N_29327,N_29143,N_29155);
xor U29328 (N_29328,N_29078,N_29002);
xor U29329 (N_29329,N_29180,N_29027);
or U29330 (N_29330,N_29191,N_29015);
xnor U29331 (N_29331,N_29162,N_29117);
nor U29332 (N_29332,N_29080,N_29096);
nand U29333 (N_29333,N_29057,N_29048);
and U29334 (N_29334,N_29043,N_29082);
xnor U29335 (N_29335,N_29096,N_29078);
nand U29336 (N_29336,N_29057,N_29056);
nor U29337 (N_29337,N_29005,N_29031);
nor U29338 (N_29338,N_29085,N_29078);
nand U29339 (N_29339,N_29002,N_29035);
or U29340 (N_29340,N_29149,N_29093);
xor U29341 (N_29341,N_29109,N_29008);
nor U29342 (N_29342,N_29053,N_29194);
nand U29343 (N_29343,N_29132,N_29156);
nor U29344 (N_29344,N_29139,N_29001);
xor U29345 (N_29345,N_29170,N_29056);
nand U29346 (N_29346,N_29145,N_29110);
or U29347 (N_29347,N_29121,N_29085);
and U29348 (N_29348,N_29056,N_29145);
or U29349 (N_29349,N_29162,N_29102);
nand U29350 (N_29350,N_29199,N_29156);
nor U29351 (N_29351,N_29097,N_29011);
nand U29352 (N_29352,N_29023,N_29172);
xor U29353 (N_29353,N_29177,N_29038);
or U29354 (N_29354,N_29164,N_29101);
xor U29355 (N_29355,N_29157,N_29103);
xnor U29356 (N_29356,N_29184,N_29185);
or U29357 (N_29357,N_29011,N_29118);
and U29358 (N_29358,N_29065,N_29101);
nand U29359 (N_29359,N_29129,N_29012);
and U29360 (N_29360,N_29025,N_29013);
and U29361 (N_29361,N_29131,N_29090);
xnor U29362 (N_29362,N_29160,N_29132);
or U29363 (N_29363,N_29006,N_29014);
or U29364 (N_29364,N_29027,N_29056);
or U29365 (N_29365,N_29094,N_29072);
xnor U29366 (N_29366,N_29024,N_29180);
xnor U29367 (N_29367,N_29153,N_29052);
or U29368 (N_29368,N_29145,N_29060);
nor U29369 (N_29369,N_29195,N_29115);
and U29370 (N_29370,N_29094,N_29017);
nand U29371 (N_29371,N_29042,N_29132);
xor U29372 (N_29372,N_29189,N_29163);
or U29373 (N_29373,N_29068,N_29185);
xnor U29374 (N_29374,N_29181,N_29023);
and U29375 (N_29375,N_29032,N_29036);
or U29376 (N_29376,N_29198,N_29032);
nand U29377 (N_29377,N_29085,N_29068);
nand U29378 (N_29378,N_29039,N_29072);
nand U29379 (N_29379,N_29158,N_29042);
nor U29380 (N_29380,N_29091,N_29074);
xnor U29381 (N_29381,N_29003,N_29063);
nand U29382 (N_29382,N_29186,N_29138);
nor U29383 (N_29383,N_29094,N_29015);
or U29384 (N_29384,N_29108,N_29016);
nand U29385 (N_29385,N_29003,N_29109);
nand U29386 (N_29386,N_29076,N_29128);
or U29387 (N_29387,N_29009,N_29010);
xor U29388 (N_29388,N_29081,N_29006);
or U29389 (N_29389,N_29048,N_29031);
or U29390 (N_29390,N_29002,N_29014);
or U29391 (N_29391,N_29185,N_29195);
xnor U29392 (N_29392,N_29188,N_29095);
nor U29393 (N_29393,N_29140,N_29198);
nand U29394 (N_29394,N_29116,N_29126);
nand U29395 (N_29395,N_29164,N_29043);
nor U29396 (N_29396,N_29084,N_29167);
nor U29397 (N_29397,N_29081,N_29035);
nand U29398 (N_29398,N_29150,N_29139);
xor U29399 (N_29399,N_29023,N_29021);
and U29400 (N_29400,N_29252,N_29353);
nor U29401 (N_29401,N_29330,N_29205);
or U29402 (N_29402,N_29337,N_29278);
and U29403 (N_29403,N_29253,N_29362);
xor U29404 (N_29404,N_29225,N_29285);
nor U29405 (N_29405,N_29383,N_29327);
nand U29406 (N_29406,N_29316,N_29206);
nor U29407 (N_29407,N_29314,N_29377);
nor U29408 (N_29408,N_29392,N_29334);
nand U29409 (N_29409,N_29222,N_29232);
and U29410 (N_29410,N_29311,N_29333);
and U29411 (N_29411,N_29323,N_29250);
or U29412 (N_29412,N_29338,N_29216);
nand U29413 (N_29413,N_29320,N_29295);
nand U29414 (N_29414,N_29254,N_29223);
nand U29415 (N_29415,N_29321,N_29275);
nor U29416 (N_29416,N_29374,N_29261);
nor U29417 (N_29417,N_29266,N_29209);
or U29418 (N_29418,N_29276,N_29345);
or U29419 (N_29419,N_29235,N_29240);
xnor U29420 (N_29420,N_29298,N_29260);
xor U29421 (N_29421,N_29279,N_29390);
xnor U29422 (N_29422,N_29322,N_29291);
or U29423 (N_29423,N_29282,N_29259);
or U29424 (N_29424,N_29356,N_29239);
or U29425 (N_29425,N_29247,N_29245);
nor U29426 (N_29426,N_29251,N_29227);
and U29427 (N_29427,N_29219,N_29286);
nand U29428 (N_29428,N_29280,N_29309);
and U29429 (N_29429,N_29344,N_29257);
and U29430 (N_29430,N_29357,N_29350);
nand U29431 (N_29431,N_29326,N_29397);
and U29432 (N_29432,N_29366,N_29290);
and U29433 (N_29433,N_29301,N_29379);
xnor U29434 (N_29434,N_29224,N_29307);
nor U29435 (N_29435,N_29358,N_29297);
or U29436 (N_29436,N_29264,N_29241);
nor U29437 (N_29437,N_29213,N_29217);
nor U29438 (N_29438,N_29233,N_29306);
nor U29439 (N_29439,N_29394,N_29207);
nor U29440 (N_29440,N_29210,N_29354);
nand U29441 (N_29441,N_29325,N_29229);
nor U29442 (N_29442,N_29317,N_29391);
nand U29443 (N_29443,N_29273,N_29352);
nand U29444 (N_29444,N_29293,N_29267);
nor U29445 (N_29445,N_29367,N_29360);
and U29446 (N_29446,N_29349,N_29339);
or U29447 (N_29447,N_29270,N_29336);
xnor U29448 (N_29448,N_29389,N_29212);
nor U29449 (N_29449,N_29200,N_29384);
xnor U29450 (N_29450,N_29343,N_29271);
nor U29451 (N_29451,N_29340,N_29378);
xnor U29452 (N_29452,N_29248,N_29371);
nand U29453 (N_29453,N_29300,N_29332);
nor U29454 (N_29454,N_29228,N_29395);
nor U29455 (N_29455,N_29364,N_29363);
and U29456 (N_29456,N_29299,N_29369);
and U29457 (N_29457,N_29399,N_29201);
xnor U29458 (N_29458,N_29351,N_29376);
or U29459 (N_29459,N_29346,N_29226);
nor U29460 (N_29460,N_29305,N_29312);
nor U29461 (N_29461,N_29368,N_29258);
nand U29462 (N_29462,N_29387,N_29236);
and U29463 (N_29463,N_29341,N_29218);
and U29464 (N_29464,N_29202,N_29361);
nor U29465 (N_29465,N_29380,N_29294);
xnor U29466 (N_29466,N_29211,N_29230);
xnor U29467 (N_29467,N_29335,N_29214);
or U29468 (N_29468,N_29234,N_29313);
nand U29469 (N_29469,N_29272,N_29302);
and U29470 (N_29470,N_29388,N_29249);
or U29471 (N_29471,N_29342,N_29382);
or U29472 (N_29472,N_29393,N_29355);
or U29473 (N_29473,N_29318,N_29396);
and U29474 (N_29474,N_29215,N_29242);
or U29475 (N_29475,N_29277,N_29329);
xor U29476 (N_29476,N_29347,N_29386);
nand U29477 (N_29477,N_29231,N_29246);
or U29478 (N_29478,N_29372,N_29373);
xor U29479 (N_29479,N_29203,N_29208);
xnor U29480 (N_29480,N_29304,N_29289);
xnor U29481 (N_29481,N_29265,N_29308);
and U29482 (N_29482,N_29237,N_29310);
xor U29483 (N_29483,N_29292,N_29263);
nor U29484 (N_29484,N_29256,N_29370);
xnor U29485 (N_29485,N_29269,N_29262);
xnor U29486 (N_29486,N_29281,N_29315);
or U29487 (N_29487,N_29255,N_29268);
and U29488 (N_29488,N_29284,N_29348);
or U29489 (N_29489,N_29287,N_29221);
or U29490 (N_29490,N_29296,N_29238);
nor U29491 (N_29491,N_29365,N_29303);
xnor U29492 (N_29492,N_29385,N_29220);
nor U29493 (N_29493,N_29328,N_29398);
or U29494 (N_29494,N_29375,N_29204);
xnor U29495 (N_29495,N_29381,N_29274);
nand U29496 (N_29496,N_29331,N_29288);
and U29497 (N_29497,N_29359,N_29244);
nand U29498 (N_29498,N_29243,N_29319);
nor U29499 (N_29499,N_29324,N_29283);
nand U29500 (N_29500,N_29345,N_29396);
or U29501 (N_29501,N_29323,N_29386);
xor U29502 (N_29502,N_29270,N_29321);
nand U29503 (N_29503,N_29335,N_29248);
nand U29504 (N_29504,N_29371,N_29312);
or U29505 (N_29505,N_29269,N_29246);
xnor U29506 (N_29506,N_29213,N_29277);
or U29507 (N_29507,N_29220,N_29311);
or U29508 (N_29508,N_29256,N_29325);
and U29509 (N_29509,N_29290,N_29271);
and U29510 (N_29510,N_29264,N_29360);
xnor U29511 (N_29511,N_29261,N_29219);
xnor U29512 (N_29512,N_29308,N_29284);
xor U29513 (N_29513,N_29270,N_29245);
nor U29514 (N_29514,N_29312,N_29366);
nor U29515 (N_29515,N_29298,N_29374);
and U29516 (N_29516,N_29309,N_29273);
and U29517 (N_29517,N_29281,N_29358);
nor U29518 (N_29518,N_29373,N_29210);
xnor U29519 (N_29519,N_29275,N_29286);
nand U29520 (N_29520,N_29392,N_29323);
xor U29521 (N_29521,N_29320,N_29205);
xor U29522 (N_29522,N_29282,N_29337);
xor U29523 (N_29523,N_29245,N_29351);
nand U29524 (N_29524,N_29214,N_29211);
nand U29525 (N_29525,N_29350,N_29236);
and U29526 (N_29526,N_29308,N_29218);
xnor U29527 (N_29527,N_29235,N_29286);
or U29528 (N_29528,N_29304,N_29373);
nand U29529 (N_29529,N_29313,N_29380);
xor U29530 (N_29530,N_29233,N_29304);
nand U29531 (N_29531,N_29349,N_29297);
xor U29532 (N_29532,N_29347,N_29283);
and U29533 (N_29533,N_29291,N_29207);
or U29534 (N_29534,N_29369,N_29200);
nor U29535 (N_29535,N_29226,N_29260);
or U29536 (N_29536,N_29278,N_29334);
or U29537 (N_29537,N_29337,N_29360);
and U29538 (N_29538,N_29205,N_29364);
and U29539 (N_29539,N_29320,N_29243);
and U29540 (N_29540,N_29221,N_29301);
and U29541 (N_29541,N_29324,N_29350);
or U29542 (N_29542,N_29335,N_29251);
or U29543 (N_29543,N_29294,N_29265);
nor U29544 (N_29544,N_29359,N_29383);
nand U29545 (N_29545,N_29289,N_29261);
nor U29546 (N_29546,N_29314,N_29341);
nand U29547 (N_29547,N_29381,N_29253);
xnor U29548 (N_29548,N_29382,N_29276);
xnor U29549 (N_29549,N_29379,N_29240);
or U29550 (N_29550,N_29250,N_29260);
and U29551 (N_29551,N_29314,N_29258);
or U29552 (N_29552,N_29226,N_29239);
nand U29553 (N_29553,N_29345,N_29337);
and U29554 (N_29554,N_29229,N_29356);
or U29555 (N_29555,N_29289,N_29298);
nor U29556 (N_29556,N_29254,N_29302);
nor U29557 (N_29557,N_29270,N_29381);
and U29558 (N_29558,N_29213,N_29334);
nor U29559 (N_29559,N_29301,N_29279);
and U29560 (N_29560,N_29223,N_29248);
nor U29561 (N_29561,N_29397,N_29369);
nor U29562 (N_29562,N_29302,N_29314);
or U29563 (N_29563,N_29315,N_29220);
xnor U29564 (N_29564,N_29369,N_29251);
and U29565 (N_29565,N_29321,N_29313);
nor U29566 (N_29566,N_29325,N_29219);
nor U29567 (N_29567,N_29317,N_29243);
nor U29568 (N_29568,N_29241,N_29392);
nor U29569 (N_29569,N_29222,N_29233);
xor U29570 (N_29570,N_29232,N_29392);
xor U29571 (N_29571,N_29357,N_29301);
and U29572 (N_29572,N_29280,N_29234);
nor U29573 (N_29573,N_29391,N_29290);
xnor U29574 (N_29574,N_29336,N_29329);
and U29575 (N_29575,N_29370,N_29278);
and U29576 (N_29576,N_29310,N_29291);
or U29577 (N_29577,N_29279,N_29364);
nor U29578 (N_29578,N_29269,N_29318);
or U29579 (N_29579,N_29206,N_29262);
xor U29580 (N_29580,N_29223,N_29287);
or U29581 (N_29581,N_29362,N_29380);
xnor U29582 (N_29582,N_29362,N_29394);
or U29583 (N_29583,N_29284,N_29342);
and U29584 (N_29584,N_29317,N_29365);
nand U29585 (N_29585,N_29357,N_29237);
nand U29586 (N_29586,N_29318,N_29209);
xor U29587 (N_29587,N_29347,N_29238);
or U29588 (N_29588,N_29214,N_29349);
nor U29589 (N_29589,N_29382,N_29286);
xnor U29590 (N_29590,N_29291,N_29239);
or U29591 (N_29591,N_29317,N_29249);
xor U29592 (N_29592,N_29319,N_29382);
xor U29593 (N_29593,N_29388,N_29251);
nand U29594 (N_29594,N_29270,N_29272);
or U29595 (N_29595,N_29395,N_29200);
xor U29596 (N_29596,N_29237,N_29358);
or U29597 (N_29597,N_29254,N_29256);
or U29598 (N_29598,N_29338,N_29221);
nand U29599 (N_29599,N_29225,N_29274);
nor U29600 (N_29600,N_29493,N_29541);
nand U29601 (N_29601,N_29467,N_29561);
nor U29602 (N_29602,N_29421,N_29411);
and U29603 (N_29603,N_29573,N_29563);
xnor U29604 (N_29604,N_29484,N_29524);
nand U29605 (N_29605,N_29526,N_29437);
nand U29606 (N_29606,N_29456,N_29431);
or U29607 (N_29607,N_29504,N_29587);
nand U29608 (N_29608,N_29550,N_29470);
xor U29609 (N_29609,N_29428,N_29507);
or U29610 (N_29610,N_29487,N_29405);
and U29611 (N_29611,N_29513,N_29511);
nor U29612 (N_29612,N_29546,N_29555);
xor U29613 (N_29613,N_29506,N_29400);
nor U29614 (N_29614,N_29407,N_29464);
nor U29615 (N_29615,N_29429,N_29551);
nand U29616 (N_29616,N_29562,N_29420);
and U29617 (N_29617,N_29443,N_29589);
nand U29618 (N_29618,N_29434,N_29578);
nand U29619 (N_29619,N_29517,N_29460);
or U29620 (N_29620,N_29591,N_29527);
nand U29621 (N_29621,N_29538,N_29455);
or U29622 (N_29622,N_29414,N_29557);
or U29623 (N_29623,N_29423,N_29415);
xnor U29624 (N_29624,N_29572,N_29536);
nor U29625 (N_29625,N_29425,N_29486);
nand U29626 (N_29626,N_29597,N_29596);
xor U29627 (N_29627,N_29522,N_29539);
xnor U29628 (N_29628,N_29413,N_29501);
nor U29629 (N_29629,N_29468,N_29595);
and U29630 (N_29630,N_29530,N_29476);
and U29631 (N_29631,N_29590,N_29445);
nand U29632 (N_29632,N_29462,N_29579);
and U29633 (N_29633,N_29548,N_29490);
or U29634 (N_29634,N_29469,N_29503);
nor U29635 (N_29635,N_29454,N_29540);
or U29636 (N_29636,N_29593,N_29565);
xor U29637 (N_29637,N_29547,N_29599);
nor U29638 (N_29638,N_29575,N_29435);
xor U29639 (N_29639,N_29520,N_29500);
nand U29640 (N_29640,N_29465,N_29427);
xor U29641 (N_29641,N_29566,N_29466);
xor U29642 (N_29642,N_29545,N_29461);
or U29643 (N_29643,N_29478,N_29471);
nand U29644 (N_29644,N_29559,N_29438);
nor U29645 (N_29645,N_29439,N_29594);
xor U29646 (N_29646,N_29577,N_29598);
nor U29647 (N_29647,N_29528,N_29518);
and U29648 (N_29648,N_29453,N_29444);
xor U29649 (N_29649,N_29446,N_29586);
nand U29650 (N_29650,N_29416,N_29406);
nand U29651 (N_29651,N_29576,N_29485);
xnor U29652 (N_29652,N_29534,N_29403);
or U29653 (N_29653,N_29404,N_29449);
xor U29654 (N_29654,N_29567,N_29532);
xor U29655 (N_29655,N_29516,N_29531);
nand U29656 (N_29656,N_29496,N_29473);
nor U29657 (N_29657,N_29521,N_29417);
nor U29658 (N_29658,N_29533,N_29560);
nor U29659 (N_29659,N_29424,N_29544);
and U29660 (N_29660,N_29489,N_29447);
nor U29661 (N_29661,N_29554,N_29479);
and U29662 (N_29662,N_29515,N_29580);
nor U29663 (N_29663,N_29452,N_29553);
and U29664 (N_29664,N_29502,N_29457);
nand U29665 (N_29665,N_29537,N_29409);
or U29666 (N_29666,N_29402,N_29477);
nor U29667 (N_29667,N_29523,N_29512);
or U29668 (N_29668,N_29472,N_29481);
nor U29669 (N_29669,N_29430,N_29574);
or U29670 (N_29670,N_29440,N_29463);
nand U29671 (N_29671,N_29535,N_29436);
or U29672 (N_29672,N_29492,N_29558);
or U29673 (N_29673,N_29571,N_29442);
xor U29674 (N_29674,N_29497,N_29418);
and U29675 (N_29675,N_29488,N_29480);
xnor U29676 (N_29676,N_29482,N_29552);
or U29677 (N_29677,N_29581,N_29529);
xor U29678 (N_29678,N_29495,N_29458);
xnor U29679 (N_29679,N_29542,N_29433);
or U29680 (N_29680,N_29491,N_29509);
and U29681 (N_29681,N_29412,N_29450);
xor U29682 (N_29682,N_29568,N_29505);
nor U29683 (N_29683,N_29525,N_29459);
nor U29684 (N_29684,N_29510,N_29583);
nor U29685 (N_29685,N_29410,N_29564);
and U29686 (N_29686,N_29419,N_29549);
or U29687 (N_29687,N_29592,N_29588);
or U29688 (N_29688,N_29475,N_29499);
nor U29689 (N_29689,N_29519,N_29508);
or U29690 (N_29690,N_29582,N_29474);
xor U29691 (N_29691,N_29422,N_29570);
nor U29692 (N_29692,N_29432,N_29584);
nand U29693 (N_29693,N_29448,N_29585);
nor U29694 (N_29694,N_29401,N_29498);
or U29695 (N_29695,N_29408,N_29514);
xnor U29696 (N_29696,N_29441,N_29451);
nor U29697 (N_29697,N_29543,N_29494);
and U29698 (N_29698,N_29426,N_29483);
or U29699 (N_29699,N_29569,N_29556);
xor U29700 (N_29700,N_29515,N_29496);
nand U29701 (N_29701,N_29419,N_29572);
xnor U29702 (N_29702,N_29409,N_29570);
xor U29703 (N_29703,N_29538,N_29471);
or U29704 (N_29704,N_29585,N_29400);
nand U29705 (N_29705,N_29474,N_29596);
nor U29706 (N_29706,N_29405,N_29536);
xnor U29707 (N_29707,N_29439,N_29575);
nor U29708 (N_29708,N_29470,N_29494);
and U29709 (N_29709,N_29449,N_29433);
and U29710 (N_29710,N_29517,N_29591);
or U29711 (N_29711,N_29430,N_29423);
and U29712 (N_29712,N_29519,N_29407);
xor U29713 (N_29713,N_29557,N_29444);
and U29714 (N_29714,N_29581,N_29461);
or U29715 (N_29715,N_29405,N_29522);
nor U29716 (N_29716,N_29519,N_29422);
nand U29717 (N_29717,N_29579,N_29437);
and U29718 (N_29718,N_29545,N_29441);
nand U29719 (N_29719,N_29458,N_29596);
or U29720 (N_29720,N_29434,N_29555);
nand U29721 (N_29721,N_29481,N_29598);
nand U29722 (N_29722,N_29482,N_29460);
or U29723 (N_29723,N_29533,N_29404);
and U29724 (N_29724,N_29431,N_29592);
and U29725 (N_29725,N_29515,N_29468);
and U29726 (N_29726,N_29441,N_29551);
nor U29727 (N_29727,N_29467,N_29547);
or U29728 (N_29728,N_29599,N_29546);
nor U29729 (N_29729,N_29521,N_29434);
xor U29730 (N_29730,N_29461,N_29544);
or U29731 (N_29731,N_29443,N_29469);
nor U29732 (N_29732,N_29552,N_29402);
xor U29733 (N_29733,N_29414,N_29582);
xnor U29734 (N_29734,N_29562,N_29556);
xnor U29735 (N_29735,N_29530,N_29565);
nand U29736 (N_29736,N_29451,N_29592);
or U29737 (N_29737,N_29450,N_29421);
xnor U29738 (N_29738,N_29542,N_29447);
nand U29739 (N_29739,N_29546,N_29590);
and U29740 (N_29740,N_29595,N_29450);
or U29741 (N_29741,N_29568,N_29411);
and U29742 (N_29742,N_29470,N_29405);
nand U29743 (N_29743,N_29405,N_29428);
xnor U29744 (N_29744,N_29426,N_29589);
nand U29745 (N_29745,N_29425,N_29540);
and U29746 (N_29746,N_29455,N_29544);
and U29747 (N_29747,N_29424,N_29558);
nand U29748 (N_29748,N_29584,N_29454);
or U29749 (N_29749,N_29443,N_29458);
xor U29750 (N_29750,N_29462,N_29464);
or U29751 (N_29751,N_29461,N_29543);
xnor U29752 (N_29752,N_29451,N_29415);
and U29753 (N_29753,N_29581,N_29561);
xor U29754 (N_29754,N_29540,N_29470);
xor U29755 (N_29755,N_29518,N_29568);
xnor U29756 (N_29756,N_29401,N_29423);
nand U29757 (N_29757,N_29550,N_29460);
nor U29758 (N_29758,N_29480,N_29402);
nand U29759 (N_29759,N_29489,N_29528);
nor U29760 (N_29760,N_29589,N_29454);
nor U29761 (N_29761,N_29423,N_29406);
nand U29762 (N_29762,N_29561,N_29508);
nor U29763 (N_29763,N_29506,N_29538);
nor U29764 (N_29764,N_29571,N_29501);
nand U29765 (N_29765,N_29503,N_29432);
nand U29766 (N_29766,N_29406,N_29414);
or U29767 (N_29767,N_29492,N_29519);
nor U29768 (N_29768,N_29459,N_29533);
nor U29769 (N_29769,N_29573,N_29591);
nor U29770 (N_29770,N_29568,N_29546);
xnor U29771 (N_29771,N_29413,N_29438);
xor U29772 (N_29772,N_29587,N_29554);
or U29773 (N_29773,N_29495,N_29463);
xor U29774 (N_29774,N_29472,N_29590);
xor U29775 (N_29775,N_29565,N_29505);
nor U29776 (N_29776,N_29585,N_29482);
nand U29777 (N_29777,N_29410,N_29572);
or U29778 (N_29778,N_29433,N_29505);
nor U29779 (N_29779,N_29436,N_29516);
xor U29780 (N_29780,N_29511,N_29493);
nand U29781 (N_29781,N_29576,N_29519);
xnor U29782 (N_29782,N_29566,N_29506);
or U29783 (N_29783,N_29587,N_29579);
xnor U29784 (N_29784,N_29515,N_29561);
xor U29785 (N_29785,N_29444,N_29511);
nor U29786 (N_29786,N_29553,N_29468);
or U29787 (N_29787,N_29569,N_29590);
nor U29788 (N_29788,N_29461,N_29595);
nor U29789 (N_29789,N_29437,N_29402);
and U29790 (N_29790,N_29435,N_29488);
xnor U29791 (N_29791,N_29457,N_29479);
and U29792 (N_29792,N_29538,N_29511);
or U29793 (N_29793,N_29402,N_29414);
and U29794 (N_29794,N_29417,N_29573);
or U29795 (N_29795,N_29496,N_29490);
and U29796 (N_29796,N_29444,N_29591);
and U29797 (N_29797,N_29455,N_29493);
xor U29798 (N_29798,N_29458,N_29422);
or U29799 (N_29799,N_29573,N_29575);
nor U29800 (N_29800,N_29773,N_29790);
xnor U29801 (N_29801,N_29761,N_29613);
nor U29802 (N_29802,N_29661,N_29635);
nor U29803 (N_29803,N_29693,N_29627);
nor U29804 (N_29804,N_29614,N_29733);
nor U29805 (N_29805,N_29641,N_29700);
xnor U29806 (N_29806,N_29665,N_29750);
nor U29807 (N_29807,N_29739,N_29651);
nor U29808 (N_29808,N_29616,N_29763);
nor U29809 (N_29809,N_29619,N_29779);
nand U29810 (N_29810,N_29685,N_29769);
and U29811 (N_29811,N_29659,N_29702);
nor U29812 (N_29812,N_29798,N_29767);
and U29813 (N_29813,N_29723,N_29724);
and U29814 (N_29814,N_29615,N_29780);
nand U29815 (N_29815,N_29755,N_29671);
or U29816 (N_29816,N_29729,N_29783);
nor U29817 (N_29817,N_29720,N_29673);
or U29818 (N_29818,N_29740,N_29623);
xor U29819 (N_29819,N_29684,N_29731);
or U29820 (N_29820,N_29725,N_29762);
or U29821 (N_29821,N_29766,N_29753);
xnor U29822 (N_29822,N_29666,N_29631);
xor U29823 (N_29823,N_29710,N_29734);
and U29824 (N_29824,N_29713,N_29620);
or U29825 (N_29825,N_29654,N_29686);
or U29826 (N_29826,N_29632,N_29677);
nor U29827 (N_29827,N_29745,N_29608);
xnor U29828 (N_29828,N_29645,N_29668);
nor U29829 (N_29829,N_29747,N_29629);
nor U29830 (N_29830,N_29704,N_29732);
nor U29831 (N_29831,N_29730,N_29652);
xor U29832 (N_29832,N_29743,N_29776);
and U29833 (N_29833,N_29751,N_29610);
or U29834 (N_29834,N_29636,N_29703);
nor U29835 (N_29835,N_29669,N_29757);
xor U29836 (N_29836,N_29716,N_29722);
nand U29837 (N_29837,N_29618,N_29603);
and U29838 (N_29838,N_29786,N_29625);
xnor U29839 (N_29839,N_29748,N_29648);
nor U29840 (N_29840,N_29737,N_29787);
and U29841 (N_29841,N_29717,N_29647);
xor U29842 (N_29842,N_29658,N_29741);
and U29843 (N_29843,N_29707,N_29656);
xor U29844 (N_29844,N_29794,N_29628);
xor U29845 (N_29845,N_29642,N_29655);
nor U29846 (N_29846,N_29676,N_29795);
nand U29847 (N_29847,N_29797,N_29672);
or U29848 (N_29848,N_29604,N_29602);
nand U29849 (N_29849,N_29742,N_29612);
or U29850 (N_29850,N_29626,N_29785);
and U29851 (N_29851,N_29774,N_29711);
and U29852 (N_29852,N_29772,N_29784);
and U29853 (N_29853,N_29796,N_29791);
nand U29854 (N_29854,N_29644,N_29775);
nand U29855 (N_29855,N_29727,N_29714);
or U29856 (N_29856,N_29678,N_29650);
xor U29857 (N_29857,N_29670,N_29736);
nand U29858 (N_29858,N_29781,N_29782);
xnor U29859 (N_29859,N_29756,N_29735);
nor U29860 (N_29860,N_29611,N_29622);
and U29861 (N_29861,N_29643,N_29709);
or U29862 (N_29862,N_29770,N_29697);
nor U29863 (N_29863,N_29768,N_29667);
and U29864 (N_29864,N_29663,N_29662);
xnor U29865 (N_29865,N_29738,N_29617);
nand U29866 (N_29866,N_29758,N_29771);
and U29867 (N_29867,N_29712,N_29696);
nor U29868 (N_29868,N_29664,N_29692);
and U29869 (N_29869,N_29701,N_29789);
or U29870 (N_29870,N_29638,N_29799);
or U29871 (N_29871,N_29752,N_29706);
nand U29872 (N_29872,N_29601,N_29721);
nor U29873 (N_29873,N_29681,N_29765);
nand U29874 (N_29874,N_29674,N_29630);
nor U29875 (N_29875,N_29675,N_29744);
xnor U29876 (N_29876,N_29690,N_29778);
and U29877 (N_29877,N_29660,N_29680);
xnor U29878 (N_29878,N_29657,N_29637);
or U29879 (N_29879,N_29705,N_29719);
and U29880 (N_29880,N_29699,N_29726);
xor U29881 (N_29881,N_29746,N_29600);
or U29882 (N_29882,N_29653,N_29760);
nor U29883 (N_29883,N_29777,N_29689);
and U29884 (N_29884,N_29640,N_29695);
nand U29885 (N_29885,N_29621,N_29633);
nor U29886 (N_29886,N_29698,N_29639);
nor U29887 (N_29887,N_29679,N_29792);
nand U29888 (N_29888,N_29788,N_29606);
xnor U29889 (N_29889,N_29759,N_29718);
or U29890 (N_29890,N_29764,N_29624);
xnor U29891 (N_29891,N_29694,N_29688);
or U29892 (N_29892,N_29609,N_29634);
or U29893 (N_29893,N_29682,N_29691);
or U29894 (N_29894,N_29646,N_29605);
or U29895 (N_29895,N_29708,N_29715);
xnor U29896 (N_29896,N_29793,N_29728);
nor U29897 (N_29897,N_29607,N_29649);
and U29898 (N_29898,N_29754,N_29687);
and U29899 (N_29899,N_29749,N_29683);
nand U29900 (N_29900,N_29653,N_29662);
xor U29901 (N_29901,N_29687,N_29706);
and U29902 (N_29902,N_29684,N_29638);
xor U29903 (N_29903,N_29789,N_29695);
nor U29904 (N_29904,N_29624,N_29715);
xnor U29905 (N_29905,N_29605,N_29627);
or U29906 (N_29906,N_29661,N_29736);
nor U29907 (N_29907,N_29750,N_29706);
or U29908 (N_29908,N_29787,N_29664);
nand U29909 (N_29909,N_29654,N_29691);
and U29910 (N_29910,N_29689,N_29731);
nor U29911 (N_29911,N_29723,N_29717);
and U29912 (N_29912,N_29665,N_29631);
or U29913 (N_29913,N_29780,N_29697);
or U29914 (N_29914,N_29630,N_29638);
nand U29915 (N_29915,N_29702,N_29791);
xnor U29916 (N_29916,N_29745,N_29740);
xor U29917 (N_29917,N_29733,N_29651);
or U29918 (N_29918,N_29788,N_29628);
nand U29919 (N_29919,N_29655,N_29737);
nand U29920 (N_29920,N_29634,N_29758);
or U29921 (N_29921,N_29635,N_29781);
and U29922 (N_29922,N_29615,N_29623);
nor U29923 (N_29923,N_29716,N_29694);
nor U29924 (N_29924,N_29610,N_29628);
nor U29925 (N_29925,N_29793,N_29798);
nand U29926 (N_29926,N_29604,N_29777);
nand U29927 (N_29927,N_29787,N_29746);
xnor U29928 (N_29928,N_29718,N_29781);
xor U29929 (N_29929,N_29778,N_29757);
nand U29930 (N_29930,N_29697,N_29783);
or U29931 (N_29931,N_29609,N_29732);
nand U29932 (N_29932,N_29794,N_29602);
or U29933 (N_29933,N_29788,N_29671);
or U29934 (N_29934,N_29717,N_29711);
nand U29935 (N_29935,N_29765,N_29744);
nor U29936 (N_29936,N_29730,N_29644);
and U29937 (N_29937,N_29729,N_29621);
or U29938 (N_29938,N_29777,N_29690);
or U29939 (N_29939,N_29734,N_29744);
or U29940 (N_29940,N_29640,N_29656);
nand U29941 (N_29941,N_29799,N_29631);
and U29942 (N_29942,N_29661,N_29654);
nand U29943 (N_29943,N_29799,N_29669);
and U29944 (N_29944,N_29751,N_29694);
or U29945 (N_29945,N_29610,N_29756);
and U29946 (N_29946,N_29754,N_29603);
and U29947 (N_29947,N_29677,N_29684);
or U29948 (N_29948,N_29745,N_29794);
and U29949 (N_29949,N_29650,N_29720);
nor U29950 (N_29950,N_29736,N_29636);
xor U29951 (N_29951,N_29746,N_29683);
and U29952 (N_29952,N_29730,N_29779);
nor U29953 (N_29953,N_29698,N_29679);
or U29954 (N_29954,N_29603,N_29793);
and U29955 (N_29955,N_29740,N_29795);
xor U29956 (N_29956,N_29708,N_29686);
nor U29957 (N_29957,N_29637,N_29631);
and U29958 (N_29958,N_29797,N_29747);
and U29959 (N_29959,N_29742,N_29619);
nor U29960 (N_29960,N_29620,N_29668);
or U29961 (N_29961,N_29770,N_29772);
or U29962 (N_29962,N_29655,N_29792);
and U29963 (N_29963,N_29711,N_29695);
xor U29964 (N_29964,N_29601,N_29671);
and U29965 (N_29965,N_29692,N_29777);
nand U29966 (N_29966,N_29793,N_29631);
nor U29967 (N_29967,N_29723,N_29698);
or U29968 (N_29968,N_29763,N_29790);
xnor U29969 (N_29969,N_29609,N_29674);
nor U29970 (N_29970,N_29643,N_29644);
or U29971 (N_29971,N_29794,N_29650);
or U29972 (N_29972,N_29768,N_29619);
xor U29973 (N_29973,N_29667,N_29707);
nor U29974 (N_29974,N_29601,N_29747);
xor U29975 (N_29975,N_29637,N_29739);
nor U29976 (N_29976,N_29656,N_29612);
xor U29977 (N_29977,N_29734,N_29633);
xnor U29978 (N_29978,N_29652,N_29666);
nor U29979 (N_29979,N_29632,N_29767);
xor U29980 (N_29980,N_29694,N_29770);
nor U29981 (N_29981,N_29657,N_29792);
or U29982 (N_29982,N_29779,N_29648);
nor U29983 (N_29983,N_29690,N_29702);
xnor U29984 (N_29984,N_29724,N_29630);
xnor U29985 (N_29985,N_29674,N_29693);
nand U29986 (N_29986,N_29632,N_29672);
nand U29987 (N_29987,N_29637,N_29644);
or U29988 (N_29988,N_29604,N_29611);
nand U29989 (N_29989,N_29702,N_29755);
xor U29990 (N_29990,N_29777,N_29770);
nor U29991 (N_29991,N_29702,N_29673);
nand U29992 (N_29992,N_29688,N_29676);
xor U29993 (N_29993,N_29608,N_29798);
xnor U29994 (N_29994,N_29607,N_29773);
and U29995 (N_29995,N_29764,N_29753);
nand U29996 (N_29996,N_29683,N_29653);
and U29997 (N_29997,N_29760,N_29640);
nor U29998 (N_29998,N_29791,N_29742);
nor U29999 (N_29999,N_29672,N_29624);
xor UO_0 (O_0,N_29841,N_29864);
xor UO_1 (O_1,N_29948,N_29925);
and UO_2 (O_2,N_29858,N_29904);
nand UO_3 (O_3,N_29827,N_29896);
xnor UO_4 (O_4,N_29870,N_29873);
or UO_5 (O_5,N_29990,N_29850);
or UO_6 (O_6,N_29851,N_29881);
nand UO_7 (O_7,N_29903,N_29820);
nand UO_8 (O_8,N_29821,N_29844);
nand UO_9 (O_9,N_29940,N_29847);
nand UO_10 (O_10,N_29938,N_29933);
and UO_11 (O_11,N_29970,N_29916);
nand UO_12 (O_12,N_29853,N_29969);
xnor UO_13 (O_13,N_29952,N_29834);
nand UO_14 (O_14,N_29900,N_29884);
or UO_15 (O_15,N_29878,N_29967);
nand UO_16 (O_16,N_29985,N_29917);
and UO_17 (O_17,N_29830,N_29800);
xnor UO_18 (O_18,N_29983,N_29959);
xnor UO_19 (O_19,N_29816,N_29951);
and UO_20 (O_20,N_29891,N_29865);
nor UO_21 (O_21,N_29910,N_29949);
nor UO_22 (O_22,N_29897,N_29918);
nand UO_23 (O_23,N_29802,N_29855);
xor UO_24 (O_24,N_29926,N_29929);
or UO_25 (O_25,N_29968,N_29857);
and UO_26 (O_26,N_29808,N_29943);
and UO_27 (O_27,N_29919,N_29845);
xor UO_28 (O_28,N_29860,N_29931);
nor UO_29 (O_29,N_29836,N_29869);
nand UO_30 (O_30,N_29861,N_29812);
and UO_31 (O_31,N_29890,N_29913);
xnor UO_32 (O_32,N_29942,N_29960);
and UO_33 (O_33,N_29965,N_29859);
or UO_34 (O_34,N_29915,N_29806);
or UO_35 (O_35,N_29912,N_29862);
and UO_36 (O_36,N_29999,N_29978);
and UO_37 (O_37,N_29976,N_29989);
nor UO_38 (O_38,N_29835,N_29966);
nor UO_39 (O_39,N_29991,N_29839);
and UO_40 (O_40,N_29901,N_29977);
nand UO_41 (O_41,N_29946,N_29921);
xor UO_42 (O_42,N_29979,N_29956);
or UO_43 (O_43,N_29838,N_29992);
nor UO_44 (O_44,N_29889,N_29930);
nand UO_45 (O_45,N_29840,N_29846);
or UO_46 (O_46,N_29981,N_29935);
and UO_47 (O_47,N_29958,N_29825);
and UO_48 (O_48,N_29909,N_29819);
nor UO_49 (O_49,N_29974,N_29975);
and UO_50 (O_50,N_29957,N_29810);
nand UO_51 (O_51,N_29815,N_29932);
nor UO_52 (O_52,N_29829,N_29934);
or UO_53 (O_53,N_29987,N_29892);
or UO_54 (O_54,N_29814,N_29995);
xor UO_55 (O_55,N_29875,N_29872);
and UO_56 (O_56,N_29818,N_29805);
and UO_57 (O_57,N_29898,N_29863);
or UO_58 (O_58,N_29843,N_29866);
or UO_59 (O_59,N_29895,N_29984);
and UO_60 (O_60,N_29950,N_29883);
and UO_61 (O_61,N_29848,N_29907);
or UO_62 (O_62,N_29964,N_29988);
nand UO_63 (O_63,N_29887,N_29828);
and UO_64 (O_64,N_29849,N_29826);
xor UO_65 (O_65,N_29945,N_29832);
xnor UO_66 (O_66,N_29920,N_29817);
and UO_67 (O_67,N_29856,N_29854);
nand UO_68 (O_68,N_29871,N_29911);
nand UO_69 (O_69,N_29971,N_29955);
xnor UO_70 (O_70,N_29982,N_29804);
nor UO_71 (O_71,N_29941,N_29868);
xnor UO_72 (O_72,N_29908,N_29824);
and UO_73 (O_73,N_29922,N_29993);
nand UO_74 (O_74,N_29962,N_29899);
and UO_75 (O_75,N_29807,N_29852);
nand UO_76 (O_76,N_29822,N_29837);
xor UO_77 (O_77,N_29998,N_29803);
nor UO_78 (O_78,N_29801,N_29980);
and UO_79 (O_79,N_29927,N_29885);
and UO_80 (O_80,N_29842,N_29973);
nand UO_81 (O_81,N_29906,N_29867);
nand UO_82 (O_82,N_29939,N_29874);
and UO_83 (O_83,N_29831,N_29823);
xor UO_84 (O_84,N_29879,N_29809);
nor UO_85 (O_85,N_29986,N_29997);
nand UO_86 (O_86,N_29963,N_29877);
xor UO_87 (O_87,N_29914,N_29876);
or UO_88 (O_88,N_29936,N_29894);
xor UO_89 (O_89,N_29880,N_29953);
and UO_90 (O_90,N_29923,N_29905);
nand UO_91 (O_91,N_29954,N_29944);
nand UO_92 (O_92,N_29937,N_29947);
nand UO_93 (O_93,N_29924,N_29928);
nor UO_94 (O_94,N_29833,N_29996);
nand UO_95 (O_95,N_29811,N_29886);
nand UO_96 (O_96,N_29972,N_29902);
nand UO_97 (O_97,N_29961,N_29882);
or UO_98 (O_98,N_29813,N_29893);
xor UO_99 (O_99,N_29888,N_29994);
nand UO_100 (O_100,N_29970,N_29995);
xnor UO_101 (O_101,N_29815,N_29903);
xnor UO_102 (O_102,N_29957,N_29808);
or UO_103 (O_103,N_29982,N_29998);
nand UO_104 (O_104,N_29989,N_29802);
nand UO_105 (O_105,N_29824,N_29963);
and UO_106 (O_106,N_29964,N_29965);
and UO_107 (O_107,N_29915,N_29854);
and UO_108 (O_108,N_29946,N_29949);
nand UO_109 (O_109,N_29998,N_29839);
xor UO_110 (O_110,N_29845,N_29896);
or UO_111 (O_111,N_29865,N_29822);
nor UO_112 (O_112,N_29845,N_29931);
xnor UO_113 (O_113,N_29975,N_29973);
or UO_114 (O_114,N_29906,N_29982);
or UO_115 (O_115,N_29821,N_29859);
or UO_116 (O_116,N_29853,N_29872);
or UO_117 (O_117,N_29943,N_29973);
or UO_118 (O_118,N_29811,N_29877);
or UO_119 (O_119,N_29956,N_29971);
and UO_120 (O_120,N_29866,N_29824);
nor UO_121 (O_121,N_29852,N_29890);
and UO_122 (O_122,N_29806,N_29819);
and UO_123 (O_123,N_29826,N_29912);
and UO_124 (O_124,N_29967,N_29832);
nor UO_125 (O_125,N_29930,N_29945);
or UO_126 (O_126,N_29977,N_29909);
and UO_127 (O_127,N_29917,N_29903);
or UO_128 (O_128,N_29993,N_29818);
and UO_129 (O_129,N_29923,N_29847);
and UO_130 (O_130,N_29849,N_29884);
nand UO_131 (O_131,N_29890,N_29843);
or UO_132 (O_132,N_29816,N_29848);
or UO_133 (O_133,N_29988,N_29808);
and UO_134 (O_134,N_29822,N_29953);
nor UO_135 (O_135,N_29885,N_29998);
nand UO_136 (O_136,N_29907,N_29841);
or UO_137 (O_137,N_29937,N_29903);
nand UO_138 (O_138,N_29936,N_29984);
nand UO_139 (O_139,N_29948,N_29817);
xor UO_140 (O_140,N_29874,N_29926);
nand UO_141 (O_141,N_29861,N_29814);
nor UO_142 (O_142,N_29872,N_29847);
xor UO_143 (O_143,N_29886,N_29852);
xnor UO_144 (O_144,N_29931,N_29894);
nand UO_145 (O_145,N_29994,N_29828);
or UO_146 (O_146,N_29800,N_29977);
and UO_147 (O_147,N_29922,N_29947);
nand UO_148 (O_148,N_29846,N_29892);
or UO_149 (O_149,N_29921,N_29962);
or UO_150 (O_150,N_29960,N_29956);
or UO_151 (O_151,N_29996,N_29897);
and UO_152 (O_152,N_29906,N_29909);
or UO_153 (O_153,N_29957,N_29982);
or UO_154 (O_154,N_29936,N_29804);
nand UO_155 (O_155,N_29954,N_29971);
or UO_156 (O_156,N_29898,N_29988);
nand UO_157 (O_157,N_29972,N_29847);
nor UO_158 (O_158,N_29914,N_29957);
nor UO_159 (O_159,N_29859,N_29959);
nor UO_160 (O_160,N_29978,N_29851);
and UO_161 (O_161,N_29891,N_29913);
nand UO_162 (O_162,N_29835,N_29976);
xnor UO_163 (O_163,N_29860,N_29803);
nor UO_164 (O_164,N_29855,N_29981);
nor UO_165 (O_165,N_29962,N_29813);
nand UO_166 (O_166,N_29896,N_29999);
or UO_167 (O_167,N_29923,N_29914);
xor UO_168 (O_168,N_29978,N_29823);
nand UO_169 (O_169,N_29906,N_29908);
and UO_170 (O_170,N_29895,N_29987);
and UO_171 (O_171,N_29811,N_29875);
or UO_172 (O_172,N_29916,N_29881);
nand UO_173 (O_173,N_29857,N_29881);
xor UO_174 (O_174,N_29928,N_29911);
xnor UO_175 (O_175,N_29836,N_29858);
nand UO_176 (O_176,N_29867,N_29809);
nor UO_177 (O_177,N_29806,N_29919);
and UO_178 (O_178,N_29823,N_29889);
nor UO_179 (O_179,N_29881,N_29967);
and UO_180 (O_180,N_29965,N_29998);
nand UO_181 (O_181,N_29802,N_29932);
xnor UO_182 (O_182,N_29866,N_29985);
nand UO_183 (O_183,N_29819,N_29942);
xnor UO_184 (O_184,N_29843,N_29881);
and UO_185 (O_185,N_29888,N_29966);
xnor UO_186 (O_186,N_29816,N_29900);
xor UO_187 (O_187,N_29954,N_29958);
or UO_188 (O_188,N_29808,N_29967);
and UO_189 (O_189,N_29906,N_29904);
nand UO_190 (O_190,N_29963,N_29883);
and UO_191 (O_191,N_29855,N_29865);
nor UO_192 (O_192,N_29833,N_29932);
and UO_193 (O_193,N_29914,N_29956);
xor UO_194 (O_194,N_29900,N_29908);
and UO_195 (O_195,N_29899,N_29854);
and UO_196 (O_196,N_29802,N_29922);
nor UO_197 (O_197,N_29801,N_29857);
xor UO_198 (O_198,N_29977,N_29861);
xnor UO_199 (O_199,N_29811,N_29922);
nand UO_200 (O_200,N_29812,N_29903);
or UO_201 (O_201,N_29853,N_29917);
or UO_202 (O_202,N_29889,N_29976);
nor UO_203 (O_203,N_29897,N_29809);
nand UO_204 (O_204,N_29932,N_29803);
nor UO_205 (O_205,N_29817,N_29952);
nand UO_206 (O_206,N_29876,N_29948);
nor UO_207 (O_207,N_29842,N_29904);
xnor UO_208 (O_208,N_29867,N_29856);
nand UO_209 (O_209,N_29987,N_29967);
and UO_210 (O_210,N_29927,N_29963);
and UO_211 (O_211,N_29989,N_29970);
or UO_212 (O_212,N_29933,N_29843);
or UO_213 (O_213,N_29963,N_29823);
nand UO_214 (O_214,N_29819,N_29871);
nor UO_215 (O_215,N_29914,N_29814);
or UO_216 (O_216,N_29917,N_29866);
nand UO_217 (O_217,N_29954,N_29984);
nor UO_218 (O_218,N_29902,N_29976);
and UO_219 (O_219,N_29944,N_29902);
nand UO_220 (O_220,N_29871,N_29942);
xor UO_221 (O_221,N_29899,N_29980);
nor UO_222 (O_222,N_29826,N_29954);
and UO_223 (O_223,N_29955,N_29902);
and UO_224 (O_224,N_29876,N_29826);
nand UO_225 (O_225,N_29927,N_29903);
nand UO_226 (O_226,N_29832,N_29848);
and UO_227 (O_227,N_29887,N_29800);
or UO_228 (O_228,N_29802,N_29903);
nor UO_229 (O_229,N_29976,N_29942);
nor UO_230 (O_230,N_29998,N_29873);
nand UO_231 (O_231,N_29863,N_29982);
and UO_232 (O_232,N_29800,N_29959);
and UO_233 (O_233,N_29859,N_29911);
nor UO_234 (O_234,N_29911,N_29901);
and UO_235 (O_235,N_29965,N_29867);
nor UO_236 (O_236,N_29837,N_29971);
and UO_237 (O_237,N_29956,N_29819);
nor UO_238 (O_238,N_29980,N_29918);
nand UO_239 (O_239,N_29881,N_29845);
or UO_240 (O_240,N_29985,N_29995);
or UO_241 (O_241,N_29908,N_29800);
xnor UO_242 (O_242,N_29948,N_29835);
or UO_243 (O_243,N_29850,N_29949);
and UO_244 (O_244,N_29856,N_29954);
nand UO_245 (O_245,N_29933,N_29918);
and UO_246 (O_246,N_29829,N_29910);
and UO_247 (O_247,N_29801,N_29874);
xor UO_248 (O_248,N_29996,N_29952);
or UO_249 (O_249,N_29926,N_29889);
nand UO_250 (O_250,N_29930,N_29813);
xnor UO_251 (O_251,N_29871,N_29864);
nand UO_252 (O_252,N_29927,N_29968);
and UO_253 (O_253,N_29932,N_29879);
or UO_254 (O_254,N_29854,N_29805);
nand UO_255 (O_255,N_29872,N_29933);
nor UO_256 (O_256,N_29979,N_29818);
nand UO_257 (O_257,N_29919,N_29947);
nand UO_258 (O_258,N_29898,N_29975);
xor UO_259 (O_259,N_29820,N_29861);
and UO_260 (O_260,N_29898,N_29938);
and UO_261 (O_261,N_29926,N_29853);
nor UO_262 (O_262,N_29894,N_29868);
xor UO_263 (O_263,N_29999,N_29939);
and UO_264 (O_264,N_29906,N_29888);
or UO_265 (O_265,N_29859,N_29994);
nor UO_266 (O_266,N_29829,N_29957);
nand UO_267 (O_267,N_29830,N_29837);
and UO_268 (O_268,N_29808,N_29906);
nor UO_269 (O_269,N_29950,N_29821);
nor UO_270 (O_270,N_29948,N_29836);
and UO_271 (O_271,N_29844,N_29907);
xnor UO_272 (O_272,N_29871,N_29939);
xor UO_273 (O_273,N_29874,N_29965);
xnor UO_274 (O_274,N_29906,N_29800);
or UO_275 (O_275,N_29857,N_29927);
nor UO_276 (O_276,N_29869,N_29973);
or UO_277 (O_277,N_29878,N_29921);
nand UO_278 (O_278,N_29865,N_29898);
nand UO_279 (O_279,N_29966,N_29864);
nor UO_280 (O_280,N_29926,N_29859);
nor UO_281 (O_281,N_29808,N_29953);
and UO_282 (O_282,N_29967,N_29838);
nor UO_283 (O_283,N_29918,N_29828);
xnor UO_284 (O_284,N_29910,N_29973);
xor UO_285 (O_285,N_29924,N_29806);
and UO_286 (O_286,N_29930,N_29996);
and UO_287 (O_287,N_29859,N_29891);
and UO_288 (O_288,N_29835,N_29860);
nor UO_289 (O_289,N_29984,N_29973);
xor UO_290 (O_290,N_29811,N_29841);
nand UO_291 (O_291,N_29939,N_29954);
and UO_292 (O_292,N_29939,N_29847);
and UO_293 (O_293,N_29903,N_29929);
nor UO_294 (O_294,N_29831,N_29857);
or UO_295 (O_295,N_29845,N_29828);
and UO_296 (O_296,N_29939,N_29968);
xnor UO_297 (O_297,N_29804,N_29865);
and UO_298 (O_298,N_29809,N_29991);
xor UO_299 (O_299,N_29923,N_29833);
and UO_300 (O_300,N_29892,N_29841);
nand UO_301 (O_301,N_29872,N_29944);
xnor UO_302 (O_302,N_29827,N_29830);
xor UO_303 (O_303,N_29826,N_29807);
nor UO_304 (O_304,N_29806,N_29953);
or UO_305 (O_305,N_29945,N_29897);
and UO_306 (O_306,N_29973,N_29922);
nand UO_307 (O_307,N_29981,N_29847);
nand UO_308 (O_308,N_29953,N_29858);
or UO_309 (O_309,N_29817,N_29802);
and UO_310 (O_310,N_29830,N_29843);
xnor UO_311 (O_311,N_29965,N_29961);
nor UO_312 (O_312,N_29806,N_29809);
xnor UO_313 (O_313,N_29902,N_29993);
nor UO_314 (O_314,N_29841,N_29895);
and UO_315 (O_315,N_29839,N_29864);
nor UO_316 (O_316,N_29880,N_29957);
nor UO_317 (O_317,N_29954,N_29983);
xor UO_318 (O_318,N_29938,N_29972);
and UO_319 (O_319,N_29952,N_29830);
nand UO_320 (O_320,N_29850,N_29964);
or UO_321 (O_321,N_29984,N_29902);
and UO_322 (O_322,N_29800,N_29816);
or UO_323 (O_323,N_29867,N_29992);
and UO_324 (O_324,N_29968,N_29928);
and UO_325 (O_325,N_29894,N_29976);
nor UO_326 (O_326,N_29902,N_29986);
nand UO_327 (O_327,N_29883,N_29984);
or UO_328 (O_328,N_29995,N_29848);
or UO_329 (O_329,N_29910,N_29805);
nand UO_330 (O_330,N_29805,N_29969);
nand UO_331 (O_331,N_29900,N_29851);
nor UO_332 (O_332,N_29856,N_29841);
xnor UO_333 (O_333,N_29824,N_29999);
and UO_334 (O_334,N_29987,N_29907);
and UO_335 (O_335,N_29951,N_29979);
or UO_336 (O_336,N_29903,N_29804);
or UO_337 (O_337,N_29827,N_29816);
nor UO_338 (O_338,N_29903,N_29928);
xnor UO_339 (O_339,N_29953,N_29968);
xor UO_340 (O_340,N_29960,N_29859);
nand UO_341 (O_341,N_29860,N_29944);
xor UO_342 (O_342,N_29917,N_29812);
nand UO_343 (O_343,N_29900,N_29945);
xor UO_344 (O_344,N_29807,N_29997);
nor UO_345 (O_345,N_29841,N_29887);
or UO_346 (O_346,N_29959,N_29809);
nor UO_347 (O_347,N_29978,N_29965);
or UO_348 (O_348,N_29808,N_29978);
nand UO_349 (O_349,N_29926,N_29877);
nor UO_350 (O_350,N_29835,N_29899);
nor UO_351 (O_351,N_29858,N_29865);
nand UO_352 (O_352,N_29848,N_29900);
xnor UO_353 (O_353,N_29831,N_29824);
or UO_354 (O_354,N_29924,N_29945);
nor UO_355 (O_355,N_29847,N_29886);
nor UO_356 (O_356,N_29857,N_29817);
nor UO_357 (O_357,N_29857,N_29833);
or UO_358 (O_358,N_29817,N_29880);
xnor UO_359 (O_359,N_29902,N_29883);
and UO_360 (O_360,N_29978,N_29853);
and UO_361 (O_361,N_29923,N_29995);
nor UO_362 (O_362,N_29879,N_29805);
nand UO_363 (O_363,N_29866,N_29946);
nand UO_364 (O_364,N_29834,N_29945);
nor UO_365 (O_365,N_29990,N_29804);
and UO_366 (O_366,N_29902,N_29962);
xnor UO_367 (O_367,N_29807,N_29820);
or UO_368 (O_368,N_29945,N_29858);
xnor UO_369 (O_369,N_29830,N_29924);
or UO_370 (O_370,N_29825,N_29867);
and UO_371 (O_371,N_29947,N_29966);
nor UO_372 (O_372,N_29846,N_29811);
nor UO_373 (O_373,N_29869,N_29893);
xor UO_374 (O_374,N_29874,N_29881);
or UO_375 (O_375,N_29808,N_29842);
xor UO_376 (O_376,N_29891,N_29964);
xor UO_377 (O_377,N_29818,N_29971);
nand UO_378 (O_378,N_29924,N_29925);
and UO_379 (O_379,N_29985,N_29958);
nor UO_380 (O_380,N_29868,N_29878);
and UO_381 (O_381,N_29829,N_29871);
nand UO_382 (O_382,N_29880,N_29995);
or UO_383 (O_383,N_29848,N_29841);
and UO_384 (O_384,N_29851,N_29862);
or UO_385 (O_385,N_29844,N_29861);
nor UO_386 (O_386,N_29859,N_29920);
nand UO_387 (O_387,N_29863,N_29932);
or UO_388 (O_388,N_29877,N_29863);
nor UO_389 (O_389,N_29901,N_29934);
xor UO_390 (O_390,N_29824,N_29872);
nor UO_391 (O_391,N_29975,N_29806);
xnor UO_392 (O_392,N_29930,N_29894);
xor UO_393 (O_393,N_29849,N_29823);
xor UO_394 (O_394,N_29980,N_29932);
or UO_395 (O_395,N_29925,N_29893);
nand UO_396 (O_396,N_29832,N_29870);
xnor UO_397 (O_397,N_29998,N_29941);
nor UO_398 (O_398,N_29892,N_29869);
nand UO_399 (O_399,N_29846,N_29895);
nand UO_400 (O_400,N_29893,N_29989);
or UO_401 (O_401,N_29812,N_29870);
or UO_402 (O_402,N_29811,N_29876);
and UO_403 (O_403,N_29848,N_29847);
and UO_404 (O_404,N_29984,N_29937);
nand UO_405 (O_405,N_29958,N_29992);
xnor UO_406 (O_406,N_29966,N_29945);
nor UO_407 (O_407,N_29987,N_29852);
xnor UO_408 (O_408,N_29906,N_29990);
or UO_409 (O_409,N_29917,N_29844);
nor UO_410 (O_410,N_29949,N_29935);
nor UO_411 (O_411,N_29854,N_29932);
nor UO_412 (O_412,N_29872,N_29922);
nor UO_413 (O_413,N_29964,N_29967);
nor UO_414 (O_414,N_29827,N_29867);
xnor UO_415 (O_415,N_29869,N_29857);
nor UO_416 (O_416,N_29972,N_29950);
nand UO_417 (O_417,N_29928,N_29804);
and UO_418 (O_418,N_29808,N_29932);
and UO_419 (O_419,N_29951,N_29909);
nor UO_420 (O_420,N_29823,N_29808);
or UO_421 (O_421,N_29892,N_29977);
or UO_422 (O_422,N_29894,N_29967);
nand UO_423 (O_423,N_29932,N_29979);
and UO_424 (O_424,N_29901,N_29971);
and UO_425 (O_425,N_29825,N_29813);
nor UO_426 (O_426,N_29906,N_29823);
xor UO_427 (O_427,N_29964,N_29821);
xor UO_428 (O_428,N_29902,N_29837);
or UO_429 (O_429,N_29967,N_29889);
nor UO_430 (O_430,N_29925,N_29858);
or UO_431 (O_431,N_29901,N_29805);
nand UO_432 (O_432,N_29994,N_29820);
nor UO_433 (O_433,N_29883,N_29975);
or UO_434 (O_434,N_29911,N_29920);
xor UO_435 (O_435,N_29811,N_29860);
and UO_436 (O_436,N_29903,N_29959);
and UO_437 (O_437,N_29917,N_29938);
nor UO_438 (O_438,N_29994,N_29870);
nand UO_439 (O_439,N_29989,N_29923);
and UO_440 (O_440,N_29952,N_29818);
or UO_441 (O_441,N_29818,N_29847);
nand UO_442 (O_442,N_29830,N_29977);
and UO_443 (O_443,N_29917,N_29849);
nand UO_444 (O_444,N_29967,N_29916);
nand UO_445 (O_445,N_29812,N_29826);
nor UO_446 (O_446,N_29936,N_29819);
and UO_447 (O_447,N_29944,N_29843);
or UO_448 (O_448,N_29823,N_29883);
xor UO_449 (O_449,N_29945,N_29804);
nand UO_450 (O_450,N_29861,N_29915);
and UO_451 (O_451,N_29826,N_29864);
nand UO_452 (O_452,N_29845,N_29818);
nor UO_453 (O_453,N_29984,N_29980);
nor UO_454 (O_454,N_29867,N_29969);
xor UO_455 (O_455,N_29871,N_29818);
nand UO_456 (O_456,N_29896,N_29930);
and UO_457 (O_457,N_29982,N_29846);
nor UO_458 (O_458,N_29914,N_29856);
and UO_459 (O_459,N_29902,N_29999);
nor UO_460 (O_460,N_29972,N_29841);
or UO_461 (O_461,N_29904,N_29871);
nand UO_462 (O_462,N_29902,N_29835);
and UO_463 (O_463,N_29838,N_29862);
or UO_464 (O_464,N_29820,N_29803);
nor UO_465 (O_465,N_29899,N_29827);
xnor UO_466 (O_466,N_29987,N_29931);
nand UO_467 (O_467,N_29828,N_29980);
or UO_468 (O_468,N_29834,N_29857);
xor UO_469 (O_469,N_29881,N_29962);
and UO_470 (O_470,N_29890,N_29849);
or UO_471 (O_471,N_29856,N_29925);
nand UO_472 (O_472,N_29972,N_29998);
and UO_473 (O_473,N_29986,N_29822);
nor UO_474 (O_474,N_29854,N_29801);
or UO_475 (O_475,N_29985,N_29963);
and UO_476 (O_476,N_29914,N_29853);
or UO_477 (O_477,N_29920,N_29842);
and UO_478 (O_478,N_29817,N_29865);
and UO_479 (O_479,N_29986,N_29914);
nor UO_480 (O_480,N_29936,N_29885);
nand UO_481 (O_481,N_29962,N_29977);
xor UO_482 (O_482,N_29838,N_29801);
and UO_483 (O_483,N_29997,N_29966);
nor UO_484 (O_484,N_29944,N_29937);
or UO_485 (O_485,N_29859,N_29834);
xor UO_486 (O_486,N_29911,N_29818);
xnor UO_487 (O_487,N_29923,N_29849);
xor UO_488 (O_488,N_29903,N_29849);
xor UO_489 (O_489,N_29991,N_29973);
xor UO_490 (O_490,N_29882,N_29936);
nor UO_491 (O_491,N_29847,N_29808);
xor UO_492 (O_492,N_29908,N_29947);
nor UO_493 (O_493,N_29830,N_29851);
nor UO_494 (O_494,N_29896,N_29892);
nor UO_495 (O_495,N_29891,N_29836);
nor UO_496 (O_496,N_29955,N_29990);
and UO_497 (O_497,N_29875,N_29834);
xnor UO_498 (O_498,N_29938,N_29874);
and UO_499 (O_499,N_29865,N_29967);
nor UO_500 (O_500,N_29889,N_29995);
nor UO_501 (O_501,N_29946,N_29889);
or UO_502 (O_502,N_29903,N_29890);
or UO_503 (O_503,N_29995,N_29992);
or UO_504 (O_504,N_29857,N_29906);
and UO_505 (O_505,N_29817,N_29834);
or UO_506 (O_506,N_29862,N_29992);
or UO_507 (O_507,N_29922,N_29921);
nor UO_508 (O_508,N_29894,N_29877);
xor UO_509 (O_509,N_29910,N_29958);
and UO_510 (O_510,N_29999,N_29911);
nand UO_511 (O_511,N_29892,N_29847);
nor UO_512 (O_512,N_29969,N_29968);
nor UO_513 (O_513,N_29845,N_29840);
xnor UO_514 (O_514,N_29940,N_29928);
nor UO_515 (O_515,N_29809,N_29862);
nand UO_516 (O_516,N_29951,N_29940);
nand UO_517 (O_517,N_29928,N_29963);
or UO_518 (O_518,N_29952,N_29801);
nor UO_519 (O_519,N_29899,N_29892);
or UO_520 (O_520,N_29918,N_29932);
xor UO_521 (O_521,N_29918,N_29948);
or UO_522 (O_522,N_29850,N_29925);
nor UO_523 (O_523,N_29847,N_29958);
nor UO_524 (O_524,N_29998,N_29994);
or UO_525 (O_525,N_29863,N_29995);
nor UO_526 (O_526,N_29962,N_29954);
nand UO_527 (O_527,N_29931,N_29969);
and UO_528 (O_528,N_29915,N_29980);
and UO_529 (O_529,N_29863,N_29856);
or UO_530 (O_530,N_29861,N_29841);
nor UO_531 (O_531,N_29931,N_29992);
nand UO_532 (O_532,N_29916,N_29810);
or UO_533 (O_533,N_29821,N_29812);
nor UO_534 (O_534,N_29999,N_29817);
xor UO_535 (O_535,N_29937,N_29871);
or UO_536 (O_536,N_29920,N_29830);
or UO_537 (O_537,N_29891,N_29981);
nand UO_538 (O_538,N_29943,N_29889);
or UO_539 (O_539,N_29979,N_29920);
or UO_540 (O_540,N_29999,N_29918);
nor UO_541 (O_541,N_29836,N_29801);
nor UO_542 (O_542,N_29992,N_29959);
nor UO_543 (O_543,N_29892,N_29944);
or UO_544 (O_544,N_29898,N_29847);
or UO_545 (O_545,N_29835,N_29984);
nand UO_546 (O_546,N_29999,N_29897);
nor UO_547 (O_547,N_29995,N_29894);
or UO_548 (O_548,N_29877,N_29976);
nand UO_549 (O_549,N_29998,N_29970);
and UO_550 (O_550,N_29975,N_29801);
and UO_551 (O_551,N_29999,N_29941);
and UO_552 (O_552,N_29961,N_29840);
and UO_553 (O_553,N_29805,N_29914);
or UO_554 (O_554,N_29948,N_29973);
and UO_555 (O_555,N_29882,N_29864);
xnor UO_556 (O_556,N_29873,N_29956);
nor UO_557 (O_557,N_29913,N_29887);
and UO_558 (O_558,N_29841,N_29831);
xor UO_559 (O_559,N_29896,N_29821);
xor UO_560 (O_560,N_29963,N_29938);
xor UO_561 (O_561,N_29963,N_29872);
or UO_562 (O_562,N_29859,N_29823);
nor UO_563 (O_563,N_29869,N_29845);
nor UO_564 (O_564,N_29968,N_29964);
nor UO_565 (O_565,N_29993,N_29890);
xor UO_566 (O_566,N_29863,N_29825);
nor UO_567 (O_567,N_29909,N_29850);
and UO_568 (O_568,N_29912,N_29813);
nor UO_569 (O_569,N_29959,N_29885);
nor UO_570 (O_570,N_29811,N_29961);
nand UO_571 (O_571,N_29949,N_29824);
or UO_572 (O_572,N_29897,N_29816);
xor UO_573 (O_573,N_29932,N_29909);
nor UO_574 (O_574,N_29805,N_29960);
xnor UO_575 (O_575,N_29959,N_29802);
nand UO_576 (O_576,N_29860,N_29808);
xnor UO_577 (O_577,N_29887,N_29870);
xor UO_578 (O_578,N_29863,N_29824);
nand UO_579 (O_579,N_29989,N_29993);
xnor UO_580 (O_580,N_29915,N_29911);
xnor UO_581 (O_581,N_29855,N_29889);
nand UO_582 (O_582,N_29888,N_29945);
xor UO_583 (O_583,N_29856,N_29824);
or UO_584 (O_584,N_29875,N_29953);
nand UO_585 (O_585,N_29995,N_29860);
nand UO_586 (O_586,N_29954,N_29879);
nor UO_587 (O_587,N_29967,N_29978);
nor UO_588 (O_588,N_29986,N_29952);
xnor UO_589 (O_589,N_29955,N_29935);
or UO_590 (O_590,N_29833,N_29998);
nor UO_591 (O_591,N_29938,N_29923);
nor UO_592 (O_592,N_29926,N_29835);
nand UO_593 (O_593,N_29812,N_29979);
nand UO_594 (O_594,N_29960,N_29940);
xnor UO_595 (O_595,N_29820,N_29841);
or UO_596 (O_596,N_29894,N_29835);
and UO_597 (O_597,N_29821,N_29827);
xnor UO_598 (O_598,N_29932,N_29872);
nor UO_599 (O_599,N_29886,N_29929);
or UO_600 (O_600,N_29881,N_29930);
or UO_601 (O_601,N_29890,N_29876);
nand UO_602 (O_602,N_29969,N_29885);
nand UO_603 (O_603,N_29930,N_29907);
nand UO_604 (O_604,N_29940,N_29901);
nand UO_605 (O_605,N_29862,N_29938);
nand UO_606 (O_606,N_29954,N_29909);
xor UO_607 (O_607,N_29965,N_29868);
nand UO_608 (O_608,N_29958,N_29819);
nand UO_609 (O_609,N_29955,N_29938);
nor UO_610 (O_610,N_29952,N_29963);
nor UO_611 (O_611,N_29855,N_29929);
nor UO_612 (O_612,N_29809,N_29876);
or UO_613 (O_613,N_29803,N_29896);
nand UO_614 (O_614,N_29879,N_29894);
or UO_615 (O_615,N_29823,N_29874);
nor UO_616 (O_616,N_29891,N_29938);
xnor UO_617 (O_617,N_29817,N_29918);
or UO_618 (O_618,N_29883,N_29916);
nor UO_619 (O_619,N_29864,N_29813);
nand UO_620 (O_620,N_29958,N_29951);
and UO_621 (O_621,N_29950,N_29997);
nor UO_622 (O_622,N_29884,N_29885);
and UO_623 (O_623,N_29916,N_29958);
and UO_624 (O_624,N_29954,N_29864);
and UO_625 (O_625,N_29925,N_29876);
and UO_626 (O_626,N_29933,N_29891);
xor UO_627 (O_627,N_29925,N_29909);
xnor UO_628 (O_628,N_29999,N_29990);
nand UO_629 (O_629,N_29980,N_29987);
xnor UO_630 (O_630,N_29985,N_29974);
and UO_631 (O_631,N_29906,N_29966);
nand UO_632 (O_632,N_29973,N_29805);
nor UO_633 (O_633,N_29926,N_29868);
nand UO_634 (O_634,N_29913,N_29843);
or UO_635 (O_635,N_29925,N_29974);
nand UO_636 (O_636,N_29858,N_29987);
nand UO_637 (O_637,N_29899,N_29911);
and UO_638 (O_638,N_29930,N_29898);
xor UO_639 (O_639,N_29851,N_29968);
and UO_640 (O_640,N_29984,N_29803);
and UO_641 (O_641,N_29895,N_29996);
nand UO_642 (O_642,N_29985,N_29825);
and UO_643 (O_643,N_29806,N_29891);
xor UO_644 (O_644,N_29946,N_29820);
nand UO_645 (O_645,N_29880,N_29859);
xnor UO_646 (O_646,N_29816,N_29831);
or UO_647 (O_647,N_29804,N_29899);
xnor UO_648 (O_648,N_29889,N_29827);
and UO_649 (O_649,N_29867,N_29952);
nor UO_650 (O_650,N_29832,N_29835);
xnor UO_651 (O_651,N_29869,N_29965);
nand UO_652 (O_652,N_29811,N_29954);
and UO_653 (O_653,N_29849,N_29983);
nor UO_654 (O_654,N_29846,N_29966);
and UO_655 (O_655,N_29846,N_29878);
xnor UO_656 (O_656,N_29929,N_29968);
nor UO_657 (O_657,N_29979,N_29870);
nand UO_658 (O_658,N_29831,N_29887);
and UO_659 (O_659,N_29988,N_29932);
nor UO_660 (O_660,N_29877,N_29950);
or UO_661 (O_661,N_29936,N_29918);
and UO_662 (O_662,N_29951,N_29943);
and UO_663 (O_663,N_29930,N_29852);
or UO_664 (O_664,N_29909,N_29821);
xor UO_665 (O_665,N_29833,N_29884);
or UO_666 (O_666,N_29861,N_29965);
xnor UO_667 (O_667,N_29933,N_29846);
nand UO_668 (O_668,N_29925,N_29995);
and UO_669 (O_669,N_29963,N_29851);
or UO_670 (O_670,N_29822,N_29959);
and UO_671 (O_671,N_29932,N_29966);
xnor UO_672 (O_672,N_29834,N_29870);
and UO_673 (O_673,N_29953,N_29947);
nand UO_674 (O_674,N_29804,N_29989);
nor UO_675 (O_675,N_29983,N_29932);
nand UO_676 (O_676,N_29895,N_29811);
nand UO_677 (O_677,N_29909,N_29995);
xnor UO_678 (O_678,N_29847,N_29900);
or UO_679 (O_679,N_29805,N_29964);
xnor UO_680 (O_680,N_29892,N_29916);
and UO_681 (O_681,N_29915,N_29816);
or UO_682 (O_682,N_29863,N_29980);
and UO_683 (O_683,N_29994,N_29855);
and UO_684 (O_684,N_29967,N_29830);
or UO_685 (O_685,N_29890,N_29988);
nand UO_686 (O_686,N_29993,N_29803);
or UO_687 (O_687,N_29995,N_29914);
and UO_688 (O_688,N_29937,N_29938);
or UO_689 (O_689,N_29807,N_29894);
xor UO_690 (O_690,N_29986,N_29812);
nand UO_691 (O_691,N_29871,N_29890);
xor UO_692 (O_692,N_29839,N_29829);
xnor UO_693 (O_693,N_29920,N_29939);
or UO_694 (O_694,N_29836,N_29881);
nor UO_695 (O_695,N_29995,N_29963);
xnor UO_696 (O_696,N_29989,N_29985);
and UO_697 (O_697,N_29820,N_29844);
and UO_698 (O_698,N_29816,N_29829);
xnor UO_699 (O_699,N_29950,N_29929);
nor UO_700 (O_700,N_29807,N_29828);
and UO_701 (O_701,N_29832,N_29817);
nor UO_702 (O_702,N_29803,N_29883);
and UO_703 (O_703,N_29993,N_29962);
nand UO_704 (O_704,N_29904,N_29801);
nand UO_705 (O_705,N_29879,N_29838);
xor UO_706 (O_706,N_29827,N_29971);
xnor UO_707 (O_707,N_29813,N_29992);
nand UO_708 (O_708,N_29807,N_29986);
nand UO_709 (O_709,N_29854,N_29968);
nor UO_710 (O_710,N_29976,N_29812);
nand UO_711 (O_711,N_29858,N_29805);
or UO_712 (O_712,N_29996,N_29811);
xnor UO_713 (O_713,N_29870,N_29821);
nand UO_714 (O_714,N_29837,N_29892);
nor UO_715 (O_715,N_29891,N_29929);
and UO_716 (O_716,N_29924,N_29969);
and UO_717 (O_717,N_29915,N_29825);
nor UO_718 (O_718,N_29937,N_29955);
xnor UO_719 (O_719,N_29871,N_29934);
nor UO_720 (O_720,N_29974,N_29952);
xor UO_721 (O_721,N_29831,N_29871);
nor UO_722 (O_722,N_29836,N_29985);
nor UO_723 (O_723,N_29958,N_29806);
nand UO_724 (O_724,N_29929,N_29853);
nand UO_725 (O_725,N_29989,N_29971);
nand UO_726 (O_726,N_29905,N_29969);
xor UO_727 (O_727,N_29877,N_29919);
xor UO_728 (O_728,N_29897,N_29827);
and UO_729 (O_729,N_29990,N_29806);
nand UO_730 (O_730,N_29912,N_29819);
or UO_731 (O_731,N_29991,N_29987);
xor UO_732 (O_732,N_29917,N_29987);
or UO_733 (O_733,N_29897,N_29887);
nor UO_734 (O_734,N_29993,N_29953);
nor UO_735 (O_735,N_29992,N_29936);
nand UO_736 (O_736,N_29927,N_29991);
nand UO_737 (O_737,N_29938,N_29858);
xor UO_738 (O_738,N_29969,N_29904);
nor UO_739 (O_739,N_29918,N_29807);
or UO_740 (O_740,N_29907,N_29832);
xor UO_741 (O_741,N_29825,N_29847);
and UO_742 (O_742,N_29903,N_29873);
nor UO_743 (O_743,N_29905,N_29877);
and UO_744 (O_744,N_29859,N_29887);
nor UO_745 (O_745,N_29827,N_29961);
or UO_746 (O_746,N_29842,N_29821);
or UO_747 (O_747,N_29922,N_29860);
nand UO_748 (O_748,N_29889,N_29873);
or UO_749 (O_749,N_29841,N_29930);
or UO_750 (O_750,N_29828,N_29831);
or UO_751 (O_751,N_29970,N_29977);
xnor UO_752 (O_752,N_29934,N_29834);
and UO_753 (O_753,N_29912,N_29994);
and UO_754 (O_754,N_29989,N_29839);
nand UO_755 (O_755,N_29826,N_29974);
or UO_756 (O_756,N_29918,N_29808);
xor UO_757 (O_757,N_29927,N_29844);
and UO_758 (O_758,N_29813,N_29928);
nand UO_759 (O_759,N_29870,N_29990);
or UO_760 (O_760,N_29964,N_29801);
xnor UO_761 (O_761,N_29954,N_29833);
or UO_762 (O_762,N_29820,N_29938);
nor UO_763 (O_763,N_29844,N_29825);
and UO_764 (O_764,N_29863,N_29974);
nor UO_765 (O_765,N_29860,N_29940);
xor UO_766 (O_766,N_29992,N_29877);
nand UO_767 (O_767,N_29959,N_29919);
or UO_768 (O_768,N_29887,N_29854);
and UO_769 (O_769,N_29801,N_29906);
nor UO_770 (O_770,N_29899,N_29937);
or UO_771 (O_771,N_29942,N_29893);
nand UO_772 (O_772,N_29965,N_29834);
nand UO_773 (O_773,N_29877,N_29851);
xnor UO_774 (O_774,N_29886,N_29834);
and UO_775 (O_775,N_29852,N_29897);
nor UO_776 (O_776,N_29929,N_29861);
nor UO_777 (O_777,N_29831,N_29900);
xor UO_778 (O_778,N_29801,N_29827);
nor UO_779 (O_779,N_29873,N_29987);
or UO_780 (O_780,N_29847,N_29868);
nand UO_781 (O_781,N_29979,N_29864);
nor UO_782 (O_782,N_29809,N_29861);
or UO_783 (O_783,N_29968,N_29897);
nor UO_784 (O_784,N_29872,N_29871);
or UO_785 (O_785,N_29869,N_29895);
nand UO_786 (O_786,N_29957,N_29932);
and UO_787 (O_787,N_29911,N_29975);
nor UO_788 (O_788,N_29880,N_29888);
and UO_789 (O_789,N_29946,N_29983);
nor UO_790 (O_790,N_29890,N_29814);
and UO_791 (O_791,N_29990,N_29836);
nand UO_792 (O_792,N_29948,N_29858);
xnor UO_793 (O_793,N_29957,N_29967);
nor UO_794 (O_794,N_29982,N_29915);
nand UO_795 (O_795,N_29940,N_29853);
xnor UO_796 (O_796,N_29977,N_29995);
xor UO_797 (O_797,N_29966,N_29996);
or UO_798 (O_798,N_29871,N_29850);
and UO_799 (O_799,N_29808,N_29960);
nand UO_800 (O_800,N_29982,N_29865);
nor UO_801 (O_801,N_29929,N_29942);
and UO_802 (O_802,N_29855,N_29859);
or UO_803 (O_803,N_29807,N_29849);
nand UO_804 (O_804,N_29841,N_29911);
nor UO_805 (O_805,N_29880,N_29856);
xor UO_806 (O_806,N_29818,N_29880);
or UO_807 (O_807,N_29988,N_29937);
nor UO_808 (O_808,N_29964,N_29847);
or UO_809 (O_809,N_29987,N_29927);
nand UO_810 (O_810,N_29822,N_29879);
and UO_811 (O_811,N_29929,N_29893);
or UO_812 (O_812,N_29827,N_29908);
nand UO_813 (O_813,N_29842,N_29800);
xnor UO_814 (O_814,N_29846,N_29970);
or UO_815 (O_815,N_29851,N_29954);
or UO_816 (O_816,N_29907,N_29973);
nor UO_817 (O_817,N_29976,N_29843);
nor UO_818 (O_818,N_29925,N_29802);
xor UO_819 (O_819,N_29988,N_29856);
and UO_820 (O_820,N_29887,N_29829);
nand UO_821 (O_821,N_29911,N_29976);
nor UO_822 (O_822,N_29972,N_29801);
nand UO_823 (O_823,N_29941,N_29971);
and UO_824 (O_824,N_29832,N_29983);
xnor UO_825 (O_825,N_29899,N_29888);
xnor UO_826 (O_826,N_29835,N_29804);
nand UO_827 (O_827,N_29895,N_29843);
and UO_828 (O_828,N_29878,N_29962);
nor UO_829 (O_829,N_29936,N_29961);
and UO_830 (O_830,N_29818,N_29933);
or UO_831 (O_831,N_29999,N_29915);
nand UO_832 (O_832,N_29891,N_29852);
or UO_833 (O_833,N_29906,N_29900);
or UO_834 (O_834,N_29863,N_29817);
xor UO_835 (O_835,N_29800,N_29993);
nand UO_836 (O_836,N_29916,N_29934);
or UO_837 (O_837,N_29919,N_29932);
and UO_838 (O_838,N_29901,N_29927);
nor UO_839 (O_839,N_29921,N_29831);
xor UO_840 (O_840,N_29983,N_29968);
nand UO_841 (O_841,N_29835,N_29831);
nor UO_842 (O_842,N_29974,N_29929);
nand UO_843 (O_843,N_29975,N_29982);
nand UO_844 (O_844,N_29842,N_29960);
and UO_845 (O_845,N_29875,N_29998);
nand UO_846 (O_846,N_29821,N_29894);
nor UO_847 (O_847,N_29841,N_29918);
xor UO_848 (O_848,N_29867,N_29986);
and UO_849 (O_849,N_29899,N_29978);
or UO_850 (O_850,N_29808,N_29810);
or UO_851 (O_851,N_29925,N_29881);
or UO_852 (O_852,N_29920,N_29800);
nor UO_853 (O_853,N_29811,N_29863);
and UO_854 (O_854,N_29875,N_29810);
nor UO_855 (O_855,N_29960,N_29817);
or UO_856 (O_856,N_29859,N_29976);
xnor UO_857 (O_857,N_29812,N_29980);
xnor UO_858 (O_858,N_29872,N_29805);
nor UO_859 (O_859,N_29857,N_29804);
nand UO_860 (O_860,N_29901,N_29928);
xnor UO_861 (O_861,N_29889,N_29846);
and UO_862 (O_862,N_29876,N_29947);
nand UO_863 (O_863,N_29871,N_29968);
nand UO_864 (O_864,N_29889,N_29867);
or UO_865 (O_865,N_29965,N_29839);
nor UO_866 (O_866,N_29924,N_29869);
nor UO_867 (O_867,N_29862,N_29963);
xnor UO_868 (O_868,N_29969,N_29834);
and UO_869 (O_869,N_29882,N_29839);
nor UO_870 (O_870,N_29859,N_29870);
nor UO_871 (O_871,N_29988,N_29829);
nor UO_872 (O_872,N_29868,N_29921);
xor UO_873 (O_873,N_29997,N_29885);
xnor UO_874 (O_874,N_29904,N_29853);
nor UO_875 (O_875,N_29929,N_29993);
or UO_876 (O_876,N_29931,N_29957);
nor UO_877 (O_877,N_29972,N_29804);
and UO_878 (O_878,N_29905,N_29824);
nor UO_879 (O_879,N_29878,N_29819);
and UO_880 (O_880,N_29822,N_29923);
nand UO_881 (O_881,N_29826,N_29973);
and UO_882 (O_882,N_29965,N_29818);
nand UO_883 (O_883,N_29814,N_29898);
xnor UO_884 (O_884,N_29949,N_29885);
or UO_885 (O_885,N_29885,N_29882);
nand UO_886 (O_886,N_29965,N_29949);
xor UO_887 (O_887,N_29882,N_29934);
and UO_888 (O_888,N_29909,N_29899);
nor UO_889 (O_889,N_29990,N_29983);
and UO_890 (O_890,N_29847,N_29850);
and UO_891 (O_891,N_29993,N_29914);
nor UO_892 (O_892,N_29984,N_29839);
nand UO_893 (O_893,N_29915,N_29837);
nand UO_894 (O_894,N_29850,N_29836);
nor UO_895 (O_895,N_29927,N_29971);
xnor UO_896 (O_896,N_29811,N_29963);
nand UO_897 (O_897,N_29828,N_29999);
nor UO_898 (O_898,N_29835,N_29946);
nor UO_899 (O_899,N_29875,N_29871);
or UO_900 (O_900,N_29864,N_29930);
or UO_901 (O_901,N_29834,N_29998);
and UO_902 (O_902,N_29984,N_29993);
xor UO_903 (O_903,N_29820,N_29809);
xnor UO_904 (O_904,N_29849,N_29851);
nor UO_905 (O_905,N_29999,N_29837);
or UO_906 (O_906,N_29979,N_29946);
and UO_907 (O_907,N_29872,N_29839);
nor UO_908 (O_908,N_29928,N_29810);
and UO_909 (O_909,N_29986,N_29961);
and UO_910 (O_910,N_29845,N_29947);
or UO_911 (O_911,N_29891,N_29819);
or UO_912 (O_912,N_29899,N_29979);
nand UO_913 (O_913,N_29962,N_29802);
and UO_914 (O_914,N_29807,N_29859);
and UO_915 (O_915,N_29854,N_29857);
nor UO_916 (O_916,N_29827,N_29873);
xnor UO_917 (O_917,N_29923,N_29898);
nand UO_918 (O_918,N_29802,N_29840);
and UO_919 (O_919,N_29981,N_29959);
nor UO_920 (O_920,N_29824,N_29965);
and UO_921 (O_921,N_29951,N_29814);
or UO_922 (O_922,N_29969,N_29944);
or UO_923 (O_923,N_29996,N_29893);
and UO_924 (O_924,N_29865,N_29885);
or UO_925 (O_925,N_29878,N_29830);
nor UO_926 (O_926,N_29865,N_29940);
and UO_927 (O_927,N_29832,N_29864);
and UO_928 (O_928,N_29869,N_29915);
and UO_929 (O_929,N_29913,N_29960);
nand UO_930 (O_930,N_29861,N_29825);
or UO_931 (O_931,N_29998,N_29869);
xnor UO_932 (O_932,N_29999,N_29849);
and UO_933 (O_933,N_29896,N_29959);
nor UO_934 (O_934,N_29856,N_29933);
or UO_935 (O_935,N_29908,N_29890);
nor UO_936 (O_936,N_29869,N_29898);
and UO_937 (O_937,N_29943,N_29958);
nor UO_938 (O_938,N_29897,N_29883);
nor UO_939 (O_939,N_29977,N_29941);
nand UO_940 (O_940,N_29881,N_29974);
nor UO_941 (O_941,N_29837,N_29900);
nand UO_942 (O_942,N_29940,N_29816);
nor UO_943 (O_943,N_29815,N_29950);
xor UO_944 (O_944,N_29973,N_29980);
nor UO_945 (O_945,N_29907,N_29977);
or UO_946 (O_946,N_29947,N_29960);
nand UO_947 (O_947,N_29936,N_29957);
nand UO_948 (O_948,N_29926,N_29932);
or UO_949 (O_949,N_29909,N_29822);
and UO_950 (O_950,N_29986,N_29848);
xor UO_951 (O_951,N_29877,N_29861);
nand UO_952 (O_952,N_29858,N_29943);
or UO_953 (O_953,N_29820,N_29857);
nand UO_954 (O_954,N_29924,N_29967);
or UO_955 (O_955,N_29845,N_29965);
nand UO_956 (O_956,N_29858,N_29956);
xor UO_957 (O_957,N_29910,N_29965);
xor UO_958 (O_958,N_29862,N_29944);
and UO_959 (O_959,N_29921,N_29979);
and UO_960 (O_960,N_29996,N_29937);
nor UO_961 (O_961,N_29931,N_29882);
and UO_962 (O_962,N_29877,N_29821);
xnor UO_963 (O_963,N_29869,N_29881);
and UO_964 (O_964,N_29976,N_29955);
or UO_965 (O_965,N_29930,N_29899);
xor UO_966 (O_966,N_29810,N_29900);
nand UO_967 (O_967,N_29919,N_29987);
nor UO_968 (O_968,N_29931,N_29918);
and UO_969 (O_969,N_29838,N_29877);
and UO_970 (O_970,N_29800,N_29823);
nor UO_971 (O_971,N_29871,N_29997);
or UO_972 (O_972,N_29818,N_29989);
nand UO_973 (O_973,N_29826,N_29919);
or UO_974 (O_974,N_29940,N_29999);
nand UO_975 (O_975,N_29857,N_29803);
or UO_976 (O_976,N_29887,N_29862);
nor UO_977 (O_977,N_29885,N_29901);
nand UO_978 (O_978,N_29887,N_29925);
nand UO_979 (O_979,N_29846,N_29893);
nor UO_980 (O_980,N_29888,N_29889);
and UO_981 (O_981,N_29970,N_29971);
xnor UO_982 (O_982,N_29809,N_29824);
nor UO_983 (O_983,N_29924,N_29825);
nand UO_984 (O_984,N_29905,N_29945);
nor UO_985 (O_985,N_29806,N_29932);
nor UO_986 (O_986,N_29899,N_29957);
and UO_987 (O_987,N_29804,N_29978);
nand UO_988 (O_988,N_29934,N_29823);
or UO_989 (O_989,N_29800,N_29869);
nand UO_990 (O_990,N_29813,N_29860);
xnor UO_991 (O_991,N_29888,N_29893);
nand UO_992 (O_992,N_29864,N_29833);
nand UO_993 (O_993,N_29900,N_29893);
nand UO_994 (O_994,N_29836,N_29868);
or UO_995 (O_995,N_29971,N_29900);
nor UO_996 (O_996,N_29827,N_29951);
nand UO_997 (O_997,N_29857,N_29953);
nor UO_998 (O_998,N_29819,N_29817);
or UO_999 (O_999,N_29845,N_29907);
xnor UO_1000 (O_1000,N_29961,N_29998);
and UO_1001 (O_1001,N_29861,N_29906);
xnor UO_1002 (O_1002,N_29897,N_29917);
or UO_1003 (O_1003,N_29997,N_29906);
nand UO_1004 (O_1004,N_29861,N_29894);
and UO_1005 (O_1005,N_29902,N_29814);
nand UO_1006 (O_1006,N_29980,N_29830);
nand UO_1007 (O_1007,N_29840,N_29878);
or UO_1008 (O_1008,N_29933,N_29950);
or UO_1009 (O_1009,N_29994,N_29917);
xnor UO_1010 (O_1010,N_29990,N_29940);
xnor UO_1011 (O_1011,N_29956,N_29867);
nor UO_1012 (O_1012,N_29917,N_29841);
or UO_1013 (O_1013,N_29997,N_29828);
nor UO_1014 (O_1014,N_29968,N_29915);
nand UO_1015 (O_1015,N_29922,N_29887);
nor UO_1016 (O_1016,N_29889,N_29884);
or UO_1017 (O_1017,N_29837,N_29978);
nor UO_1018 (O_1018,N_29919,N_29910);
or UO_1019 (O_1019,N_29879,N_29858);
or UO_1020 (O_1020,N_29954,N_29927);
and UO_1021 (O_1021,N_29910,N_29911);
and UO_1022 (O_1022,N_29863,N_29985);
nand UO_1023 (O_1023,N_29947,N_29867);
or UO_1024 (O_1024,N_29850,N_29967);
or UO_1025 (O_1025,N_29824,N_29834);
xnor UO_1026 (O_1026,N_29967,N_29853);
nor UO_1027 (O_1027,N_29996,N_29946);
nand UO_1028 (O_1028,N_29991,N_29814);
and UO_1029 (O_1029,N_29837,N_29931);
nor UO_1030 (O_1030,N_29941,N_29891);
nor UO_1031 (O_1031,N_29934,N_29827);
nor UO_1032 (O_1032,N_29993,N_29877);
or UO_1033 (O_1033,N_29962,N_29959);
xnor UO_1034 (O_1034,N_29827,N_29875);
and UO_1035 (O_1035,N_29973,N_29900);
nor UO_1036 (O_1036,N_29840,N_29942);
and UO_1037 (O_1037,N_29873,N_29904);
nand UO_1038 (O_1038,N_29894,N_29816);
nor UO_1039 (O_1039,N_29834,N_29957);
nor UO_1040 (O_1040,N_29978,N_29968);
nand UO_1041 (O_1041,N_29936,N_29857);
or UO_1042 (O_1042,N_29997,N_29815);
and UO_1043 (O_1043,N_29931,N_29973);
nand UO_1044 (O_1044,N_29935,N_29932);
and UO_1045 (O_1045,N_29926,N_29867);
nand UO_1046 (O_1046,N_29893,N_29815);
xnor UO_1047 (O_1047,N_29927,N_29919);
nand UO_1048 (O_1048,N_29974,N_29827);
nor UO_1049 (O_1049,N_29902,N_29820);
and UO_1050 (O_1050,N_29850,N_29999);
and UO_1051 (O_1051,N_29975,N_29918);
and UO_1052 (O_1052,N_29961,N_29836);
or UO_1053 (O_1053,N_29937,N_29823);
or UO_1054 (O_1054,N_29807,N_29996);
xnor UO_1055 (O_1055,N_29842,N_29969);
xor UO_1056 (O_1056,N_29851,N_29996);
nor UO_1057 (O_1057,N_29884,N_29839);
or UO_1058 (O_1058,N_29819,N_29896);
nor UO_1059 (O_1059,N_29970,N_29980);
xnor UO_1060 (O_1060,N_29914,N_29979);
and UO_1061 (O_1061,N_29993,N_29821);
nor UO_1062 (O_1062,N_29817,N_29875);
nand UO_1063 (O_1063,N_29994,N_29913);
nor UO_1064 (O_1064,N_29809,N_29878);
xnor UO_1065 (O_1065,N_29809,N_29946);
or UO_1066 (O_1066,N_29886,N_29935);
and UO_1067 (O_1067,N_29865,N_29985);
or UO_1068 (O_1068,N_29878,N_29807);
nor UO_1069 (O_1069,N_29807,N_29944);
or UO_1070 (O_1070,N_29993,N_29828);
or UO_1071 (O_1071,N_29842,N_29895);
nor UO_1072 (O_1072,N_29812,N_29863);
nand UO_1073 (O_1073,N_29854,N_29804);
or UO_1074 (O_1074,N_29976,N_29983);
nand UO_1075 (O_1075,N_29983,N_29998);
xor UO_1076 (O_1076,N_29950,N_29873);
and UO_1077 (O_1077,N_29830,N_29993);
nand UO_1078 (O_1078,N_29817,N_29876);
nand UO_1079 (O_1079,N_29995,N_29845);
and UO_1080 (O_1080,N_29904,N_29909);
and UO_1081 (O_1081,N_29935,N_29848);
nor UO_1082 (O_1082,N_29995,N_29906);
and UO_1083 (O_1083,N_29991,N_29864);
nand UO_1084 (O_1084,N_29942,N_29902);
or UO_1085 (O_1085,N_29894,N_29829);
and UO_1086 (O_1086,N_29949,N_29991);
nor UO_1087 (O_1087,N_29850,N_29919);
and UO_1088 (O_1088,N_29857,N_29893);
nor UO_1089 (O_1089,N_29821,N_29980);
and UO_1090 (O_1090,N_29821,N_29959);
and UO_1091 (O_1091,N_29884,N_29901);
nand UO_1092 (O_1092,N_29874,N_29924);
or UO_1093 (O_1093,N_29801,N_29868);
nor UO_1094 (O_1094,N_29950,N_29941);
nor UO_1095 (O_1095,N_29828,N_29920);
nand UO_1096 (O_1096,N_29972,N_29965);
and UO_1097 (O_1097,N_29813,N_29826);
or UO_1098 (O_1098,N_29983,N_29893);
xnor UO_1099 (O_1099,N_29805,N_29878);
nand UO_1100 (O_1100,N_29809,N_29885);
nor UO_1101 (O_1101,N_29966,N_29865);
nand UO_1102 (O_1102,N_29877,N_29943);
and UO_1103 (O_1103,N_29800,N_29924);
and UO_1104 (O_1104,N_29902,N_29888);
and UO_1105 (O_1105,N_29816,N_29896);
nand UO_1106 (O_1106,N_29974,N_29949);
nand UO_1107 (O_1107,N_29941,N_29962);
nand UO_1108 (O_1108,N_29920,N_29915);
and UO_1109 (O_1109,N_29837,N_29879);
and UO_1110 (O_1110,N_29991,N_29845);
or UO_1111 (O_1111,N_29841,N_29806);
and UO_1112 (O_1112,N_29942,N_29894);
nand UO_1113 (O_1113,N_29873,N_29995);
or UO_1114 (O_1114,N_29864,N_29939);
nand UO_1115 (O_1115,N_29858,N_29910);
or UO_1116 (O_1116,N_29950,N_29979);
nor UO_1117 (O_1117,N_29998,N_29910);
nor UO_1118 (O_1118,N_29997,N_29895);
and UO_1119 (O_1119,N_29887,N_29950);
nor UO_1120 (O_1120,N_29939,N_29907);
and UO_1121 (O_1121,N_29865,N_29957);
nand UO_1122 (O_1122,N_29862,N_29961);
xor UO_1123 (O_1123,N_29914,N_29818);
nor UO_1124 (O_1124,N_29821,N_29912);
xnor UO_1125 (O_1125,N_29882,N_29979);
xnor UO_1126 (O_1126,N_29976,N_29931);
nor UO_1127 (O_1127,N_29800,N_29841);
nor UO_1128 (O_1128,N_29870,N_29889);
or UO_1129 (O_1129,N_29902,N_29869);
and UO_1130 (O_1130,N_29948,N_29888);
and UO_1131 (O_1131,N_29942,N_29946);
nor UO_1132 (O_1132,N_29905,N_29847);
and UO_1133 (O_1133,N_29951,N_29997);
and UO_1134 (O_1134,N_29863,N_29946);
nor UO_1135 (O_1135,N_29999,N_29895);
nor UO_1136 (O_1136,N_29860,N_29907);
or UO_1137 (O_1137,N_29972,N_29994);
xnor UO_1138 (O_1138,N_29848,N_29851);
nor UO_1139 (O_1139,N_29955,N_29811);
and UO_1140 (O_1140,N_29861,N_29878);
or UO_1141 (O_1141,N_29859,N_29867);
or UO_1142 (O_1142,N_29940,N_29825);
nand UO_1143 (O_1143,N_29849,N_29958);
nand UO_1144 (O_1144,N_29839,N_29946);
nor UO_1145 (O_1145,N_29941,N_29978);
or UO_1146 (O_1146,N_29947,N_29965);
xnor UO_1147 (O_1147,N_29927,N_29804);
nor UO_1148 (O_1148,N_29832,N_29919);
xor UO_1149 (O_1149,N_29950,N_29939);
or UO_1150 (O_1150,N_29990,N_29897);
nor UO_1151 (O_1151,N_29877,N_29802);
xor UO_1152 (O_1152,N_29815,N_29801);
or UO_1153 (O_1153,N_29962,N_29815);
or UO_1154 (O_1154,N_29806,N_29838);
xnor UO_1155 (O_1155,N_29968,N_29836);
or UO_1156 (O_1156,N_29886,N_29989);
or UO_1157 (O_1157,N_29830,N_29829);
or UO_1158 (O_1158,N_29800,N_29840);
xnor UO_1159 (O_1159,N_29992,N_29942);
xnor UO_1160 (O_1160,N_29821,N_29996);
or UO_1161 (O_1161,N_29915,N_29873);
and UO_1162 (O_1162,N_29864,N_29905);
nor UO_1163 (O_1163,N_29803,N_29972);
nand UO_1164 (O_1164,N_29812,N_29846);
xnor UO_1165 (O_1165,N_29891,N_29907);
xor UO_1166 (O_1166,N_29854,N_29989);
or UO_1167 (O_1167,N_29810,N_29872);
and UO_1168 (O_1168,N_29956,N_29942);
and UO_1169 (O_1169,N_29842,N_29858);
nand UO_1170 (O_1170,N_29811,N_29923);
nand UO_1171 (O_1171,N_29924,N_29905);
or UO_1172 (O_1172,N_29822,N_29943);
nor UO_1173 (O_1173,N_29893,N_29915);
nand UO_1174 (O_1174,N_29813,N_29855);
nor UO_1175 (O_1175,N_29927,N_29977);
or UO_1176 (O_1176,N_29938,N_29951);
and UO_1177 (O_1177,N_29907,N_29808);
xnor UO_1178 (O_1178,N_29921,N_29889);
nor UO_1179 (O_1179,N_29826,N_29806);
and UO_1180 (O_1180,N_29987,N_29823);
xnor UO_1181 (O_1181,N_29955,N_29973);
and UO_1182 (O_1182,N_29914,N_29968);
and UO_1183 (O_1183,N_29954,N_29998);
xnor UO_1184 (O_1184,N_29912,N_29935);
and UO_1185 (O_1185,N_29836,N_29887);
or UO_1186 (O_1186,N_29895,N_29998);
and UO_1187 (O_1187,N_29823,N_29838);
and UO_1188 (O_1188,N_29893,N_29858);
nor UO_1189 (O_1189,N_29911,N_29848);
xor UO_1190 (O_1190,N_29885,N_29955);
or UO_1191 (O_1191,N_29932,N_29965);
and UO_1192 (O_1192,N_29896,N_29844);
xnor UO_1193 (O_1193,N_29899,N_29908);
or UO_1194 (O_1194,N_29826,N_29939);
nand UO_1195 (O_1195,N_29889,N_29903);
and UO_1196 (O_1196,N_29981,N_29865);
and UO_1197 (O_1197,N_29925,N_29999);
or UO_1198 (O_1198,N_29912,N_29913);
or UO_1199 (O_1199,N_29979,N_29819);
nor UO_1200 (O_1200,N_29861,N_29807);
nand UO_1201 (O_1201,N_29878,N_29816);
nor UO_1202 (O_1202,N_29877,N_29904);
and UO_1203 (O_1203,N_29983,N_29802);
xor UO_1204 (O_1204,N_29949,N_29985);
or UO_1205 (O_1205,N_29988,N_29843);
nor UO_1206 (O_1206,N_29995,N_29986);
nand UO_1207 (O_1207,N_29831,N_29965);
nor UO_1208 (O_1208,N_29981,N_29870);
and UO_1209 (O_1209,N_29864,N_29956);
nor UO_1210 (O_1210,N_29959,N_29828);
xor UO_1211 (O_1211,N_29917,N_29839);
nand UO_1212 (O_1212,N_29828,N_29971);
or UO_1213 (O_1213,N_29854,N_29837);
nor UO_1214 (O_1214,N_29854,N_29891);
and UO_1215 (O_1215,N_29993,N_29933);
nand UO_1216 (O_1216,N_29975,N_29999);
nor UO_1217 (O_1217,N_29870,N_29914);
nor UO_1218 (O_1218,N_29909,N_29859);
nand UO_1219 (O_1219,N_29975,N_29810);
nor UO_1220 (O_1220,N_29889,N_29822);
nor UO_1221 (O_1221,N_29819,N_29971);
and UO_1222 (O_1222,N_29916,N_29996);
and UO_1223 (O_1223,N_29827,N_29843);
nor UO_1224 (O_1224,N_29857,N_29994);
nor UO_1225 (O_1225,N_29810,N_29960);
and UO_1226 (O_1226,N_29852,N_29806);
or UO_1227 (O_1227,N_29825,N_29968);
or UO_1228 (O_1228,N_29888,N_29936);
xnor UO_1229 (O_1229,N_29891,N_29877);
and UO_1230 (O_1230,N_29846,N_29899);
xnor UO_1231 (O_1231,N_29832,N_29935);
nand UO_1232 (O_1232,N_29858,N_29869);
nand UO_1233 (O_1233,N_29835,N_29930);
xnor UO_1234 (O_1234,N_29969,N_29918);
nand UO_1235 (O_1235,N_29905,N_29858);
xor UO_1236 (O_1236,N_29922,N_29858);
xor UO_1237 (O_1237,N_29939,N_29989);
nand UO_1238 (O_1238,N_29903,N_29920);
nand UO_1239 (O_1239,N_29911,N_29805);
nand UO_1240 (O_1240,N_29967,N_29836);
nor UO_1241 (O_1241,N_29824,N_29929);
nand UO_1242 (O_1242,N_29960,N_29828);
or UO_1243 (O_1243,N_29973,N_29930);
and UO_1244 (O_1244,N_29880,N_29930);
or UO_1245 (O_1245,N_29877,N_29885);
or UO_1246 (O_1246,N_29897,N_29817);
xnor UO_1247 (O_1247,N_29808,N_29944);
and UO_1248 (O_1248,N_29966,N_29859);
xnor UO_1249 (O_1249,N_29873,N_29918);
and UO_1250 (O_1250,N_29923,N_29931);
or UO_1251 (O_1251,N_29879,N_29803);
nand UO_1252 (O_1252,N_29945,N_29866);
and UO_1253 (O_1253,N_29803,N_29951);
nand UO_1254 (O_1254,N_29936,N_29823);
and UO_1255 (O_1255,N_29890,N_29816);
or UO_1256 (O_1256,N_29848,N_29975);
and UO_1257 (O_1257,N_29974,N_29850);
nand UO_1258 (O_1258,N_29916,N_29914);
nand UO_1259 (O_1259,N_29982,N_29867);
nor UO_1260 (O_1260,N_29868,N_29880);
xor UO_1261 (O_1261,N_29832,N_29968);
nand UO_1262 (O_1262,N_29994,N_29940);
nand UO_1263 (O_1263,N_29944,N_29867);
nand UO_1264 (O_1264,N_29878,N_29968);
xor UO_1265 (O_1265,N_29852,N_29841);
nand UO_1266 (O_1266,N_29993,N_29834);
or UO_1267 (O_1267,N_29970,N_29885);
or UO_1268 (O_1268,N_29932,N_29897);
xnor UO_1269 (O_1269,N_29810,N_29924);
or UO_1270 (O_1270,N_29953,N_29997);
and UO_1271 (O_1271,N_29803,N_29954);
xnor UO_1272 (O_1272,N_29986,N_29907);
nand UO_1273 (O_1273,N_29921,N_29956);
or UO_1274 (O_1274,N_29899,N_29834);
and UO_1275 (O_1275,N_29847,N_29889);
nand UO_1276 (O_1276,N_29969,N_29837);
xor UO_1277 (O_1277,N_29849,N_29864);
or UO_1278 (O_1278,N_29848,N_29959);
or UO_1279 (O_1279,N_29995,N_29822);
xnor UO_1280 (O_1280,N_29899,N_29844);
nor UO_1281 (O_1281,N_29950,N_29964);
and UO_1282 (O_1282,N_29962,N_29950);
nand UO_1283 (O_1283,N_29871,N_29955);
nand UO_1284 (O_1284,N_29935,N_29901);
or UO_1285 (O_1285,N_29882,N_29872);
nor UO_1286 (O_1286,N_29979,N_29886);
nand UO_1287 (O_1287,N_29810,N_29833);
and UO_1288 (O_1288,N_29917,N_29803);
and UO_1289 (O_1289,N_29881,N_29939);
nand UO_1290 (O_1290,N_29827,N_29900);
nor UO_1291 (O_1291,N_29861,N_29887);
or UO_1292 (O_1292,N_29905,N_29853);
xnor UO_1293 (O_1293,N_29984,N_29958);
nor UO_1294 (O_1294,N_29920,N_29978);
xnor UO_1295 (O_1295,N_29844,N_29965);
nand UO_1296 (O_1296,N_29863,N_29803);
nor UO_1297 (O_1297,N_29970,N_29925);
and UO_1298 (O_1298,N_29955,N_29895);
and UO_1299 (O_1299,N_29965,N_29948);
or UO_1300 (O_1300,N_29801,N_29823);
xnor UO_1301 (O_1301,N_29822,N_29827);
nand UO_1302 (O_1302,N_29866,N_29904);
nor UO_1303 (O_1303,N_29985,N_29818);
nor UO_1304 (O_1304,N_29945,N_29848);
nor UO_1305 (O_1305,N_29951,N_29847);
xor UO_1306 (O_1306,N_29957,N_29813);
and UO_1307 (O_1307,N_29891,N_29801);
nand UO_1308 (O_1308,N_29835,N_29917);
and UO_1309 (O_1309,N_29976,N_29830);
and UO_1310 (O_1310,N_29938,N_29931);
and UO_1311 (O_1311,N_29890,N_29840);
and UO_1312 (O_1312,N_29805,N_29959);
nand UO_1313 (O_1313,N_29888,N_29827);
nand UO_1314 (O_1314,N_29831,N_29844);
or UO_1315 (O_1315,N_29975,N_29913);
xnor UO_1316 (O_1316,N_29912,N_29961);
xor UO_1317 (O_1317,N_29857,N_29926);
and UO_1318 (O_1318,N_29841,N_29937);
nand UO_1319 (O_1319,N_29859,N_29851);
nand UO_1320 (O_1320,N_29972,N_29824);
nor UO_1321 (O_1321,N_29865,N_29991);
xor UO_1322 (O_1322,N_29923,N_29925);
and UO_1323 (O_1323,N_29978,N_29900);
xnor UO_1324 (O_1324,N_29952,N_29878);
xor UO_1325 (O_1325,N_29949,N_29891);
nor UO_1326 (O_1326,N_29910,N_29862);
or UO_1327 (O_1327,N_29974,N_29910);
xor UO_1328 (O_1328,N_29916,N_29920);
nand UO_1329 (O_1329,N_29965,N_29887);
nor UO_1330 (O_1330,N_29923,N_29928);
and UO_1331 (O_1331,N_29813,N_29889);
xor UO_1332 (O_1332,N_29854,N_29955);
xor UO_1333 (O_1333,N_29940,N_29932);
nor UO_1334 (O_1334,N_29838,N_29922);
and UO_1335 (O_1335,N_29976,N_29963);
and UO_1336 (O_1336,N_29846,N_29940);
nor UO_1337 (O_1337,N_29872,N_29964);
nand UO_1338 (O_1338,N_29959,N_29940);
or UO_1339 (O_1339,N_29995,N_29807);
xnor UO_1340 (O_1340,N_29882,N_29972);
or UO_1341 (O_1341,N_29897,N_29913);
xnor UO_1342 (O_1342,N_29920,N_29973);
and UO_1343 (O_1343,N_29998,N_29861);
and UO_1344 (O_1344,N_29962,N_29990);
xor UO_1345 (O_1345,N_29915,N_29927);
nor UO_1346 (O_1346,N_29943,N_29934);
and UO_1347 (O_1347,N_29863,N_29953);
nor UO_1348 (O_1348,N_29934,N_29931);
nor UO_1349 (O_1349,N_29800,N_29966);
xnor UO_1350 (O_1350,N_29823,N_29922);
nor UO_1351 (O_1351,N_29813,N_29829);
nand UO_1352 (O_1352,N_29850,N_29902);
nand UO_1353 (O_1353,N_29991,N_29976);
nor UO_1354 (O_1354,N_29864,N_29993);
and UO_1355 (O_1355,N_29819,N_29811);
nand UO_1356 (O_1356,N_29974,N_29828);
xor UO_1357 (O_1357,N_29805,N_29933);
and UO_1358 (O_1358,N_29967,N_29862);
nand UO_1359 (O_1359,N_29993,N_29918);
or UO_1360 (O_1360,N_29982,N_29935);
xnor UO_1361 (O_1361,N_29956,N_29820);
xor UO_1362 (O_1362,N_29930,N_29943);
xnor UO_1363 (O_1363,N_29908,N_29850);
nand UO_1364 (O_1364,N_29801,N_29988);
xnor UO_1365 (O_1365,N_29854,N_29822);
or UO_1366 (O_1366,N_29935,N_29928);
nor UO_1367 (O_1367,N_29980,N_29891);
xor UO_1368 (O_1368,N_29840,N_29914);
or UO_1369 (O_1369,N_29937,N_29924);
nand UO_1370 (O_1370,N_29967,N_29973);
and UO_1371 (O_1371,N_29954,N_29881);
and UO_1372 (O_1372,N_29988,N_29879);
xor UO_1373 (O_1373,N_29800,N_29893);
nor UO_1374 (O_1374,N_29917,N_29810);
or UO_1375 (O_1375,N_29877,N_29858);
xor UO_1376 (O_1376,N_29901,N_29983);
xnor UO_1377 (O_1377,N_29816,N_29895);
nor UO_1378 (O_1378,N_29899,N_29840);
or UO_1379 (O_1379,N_29807,N_29905);
nor UO_1380 (O_1380,N_29818,N_29835);
or UO_1381 (O_1381,N_29903,N_29964);
nor UO_1382 (O_1382,N_29927,N_29983);
or UO_1383 (O_1383,N_29819,N_29832);
nand UO_1384 (O_1384,N_29801,N_29987);
or UO_1385 (O_1385,N_29811,N_29836);
or UO_1386 (O_1386,N_29887,N_29906);
nand UO_1387 (O_1387,N_29888,N_29933);
or UO_1388 (O_1388,N_29811,N_29956);
nor UO_1389 (O_1389,N_29966,N_29887);
or UO_1390 (O_1390,N_29908,N_29917);
nand UO_1391 (O_1391,N_29869,N_29941);
xnor UO_1392 (O_1392,N_29893,N_29847);
xor UO_1393 (O_1393,N_29929,N_29868);
nor UO_1394 (O_1394,N_29873,N_29894);
xnor UO_1395 (O_1395,N_29948,N_29845);
or UO_1396 (O_1396,N_29945,N_29958);
and UO_1397 (O_1397,N_29961,N_29838);
nor UO_1398 (O_1398,N_29859,N_29939);
and UO_1399 (O_1399,N_29850,N_29966);
nand UO_1400 (O_1400,N_29987,N_29902);
xor UO_1401 (O_1401,N_29852,N_29953);
or UO_1402 (O_1402,N_29892,N_29885);
xnor UO_1403 (O_1403,N_29897,N_29896);
xor UO_1404 (O_1404,N_29908,N_29918);
or UO_1405 (O_1405,N_29861,N_29971);
nand UO_1406 (O_1406,N_29824,N_29845);
nand UO_1407 (O_1407,N_29801,N_29841);
or UO_1408 (O_1408,N_29845,N_29867);
and UO_1409 (O_1409,N_29851,N_29897);
xor UO_1410 (O_1410,N_29986,N_29901);
or UO_1411 (O_1411,N_29945,N_29852);
nor UO_1412 (O_1412,N_29983,N_29826);
nor UO_1413 (O_1413,N_29899,N_29971);
nand UO_1414 (O_1414,N_29957,N_29812);
nor UO_1415 (O_1415,N_29874,N_29913);
and UO_1416 (O_1416,N_29885,N_29967);
nor UO_1417 (O_1417,N_29888,N_29955);
xnor UO_1418 (O_1418,N_29846,N_29851);
and UO_1419 (O_1419,N_29888,N_29809);
xnor UO_1420 (O_1420,N_29990,N_29957);
nand UO_1421 (O_1421,N_29817,N_29855);
and UO_1422 (O_1422,N_29810,N_29904);
or UO_1423 (O_1423,N_29893,N_29810);
nor UO_1424 (O_1424,N_29936,N_29965);
nand UO_1425 (O_1425,N_29955,N_29860);
nand UO_1426 (O_1426,N_29997,N_29919);
nand UO_1427 (O_1427,N_29968,N_29962);
nor UO_1428 (O_1428,N_29927,N_29860);
or UO_1429 (O_1429,N_29920,N_29930);
nor UO_1430 (O_1430,N_29909,N_29901);
nand UO_1431 (O_1431,N_29922,N_29828);
and UO_1432 (O_1432,N_29840,N_29862);
and UO_1433 (O_1433,N_29852,N_29962);
or UO_1434 (O_1434,N_29975,N_29985);
nand UO_1435 (O_1435,N_29958,N_29999);
nor UO_1436 (O_1436,N_29976,N_29820);
nor UO_1437 (O_1437,N_29959,N_29869);
xnor UO_1438 (O_1438,N_29876,N_29933);
and UO_1439 (O_1439,N_29852,N_29935);
and UO_1440 (O_1440,N_29960,N_29991);
nand UO_1441 (O_1441,N_29998,N_29993);
and UO_1442 (O_1442,N_29924,N_29836);
nor UO_1443 (O_1443,N_29874,N_29901);
or UO_1444 (O_1444,N_29817,N_29830);
nor UO_1445 (O_1445,N_29920,N_29960);
nor UO_1446 (O_1446,N_29842,N_29886);
and UO_1447 (O_1447,N_29801,N_29956);
xnor UO_1448 (O_1448,N_29887,N_29990);
and UO_1449 (O_1449,N_29959,N_29927);
or UO_1450 (O_1450,N_29925,N_29874);
xor UO_1451 (O_1451,N_29895,N_29971);
nor UO_1452 (O_1452,N_29912,N_29899);
and UO_1453 (O_1453,N_29991,N_29965);
xnor UO_1454 (O_1454,N_29898,N_29844);
and UO_1455 (O_1455,N_29942,N_29977);
or UO_1456 (O_1456,N_29866,N_29855);
and UO_1457 (O_1457,N_29986,N_29927);
and UO_1458 (O_1458,N_29928,N_29855);
nor UO_1459 (O_1459,N_29872,N_29951);
nand UO_1460 (O_1460,N_29985,N_29844);
nand UO_1461 (O_1461,N_29999,N_29882);
nor UO_1462 (O_1462,N_29919,N_29822);
xor UO_1463 (O_1463,N_29871,N_29941);
or UO_1464 (O_1464,N_29981,N_29908);
xor UO_1465 (O_1465,N_29835,N_29851);
xnor UO_1466 (O_1466,N_29964,N_29908);
or UO_1467 (O_1467,N_29873,N_29839);
xnor UO_1468 (O_1468,N_29821,N_29865);
xnor UO_1469 (O_1469,N_29867,N_29997);
xor UO_1470 (O_1470,N_29824,N_29950);
and UO_1471 (O_1471,N_29857,N_29951);
nor UO_1472 (O_1472,N_29935,N_29941);
xnor UO_1473 (O_1473,N_29910,N_29847);
or UO_1474 (O_1474,N_29968,N_29973);
or UO_1475 (O_1475,N_29937,N_29821);
and UO_1476 (O_1476,N_29923,N_29842);
xor UO_1477 (O_1477,N_29945,N_29938);
nor UO_1478 (O_1478,N_29976,N_29953);
nor UO_1479 (O_1479,N_29888,N_29916);
nor UO_1480 (O_1480,N_29895,N_29844);
nor UO_1481 (O_1481,N_29858,N_29840);
xnor UO_1482 (O_1482,N_29878,N_29899);
or UO_1483 (O_1483,N_29811,N_29894);
or UO_1484 (O_1484,N_29896,N_29806);
or UO_1485 (O_1485,N_29842,N_29852);
and UO_1486 (O_1486,N_29981,N_29920);
nand UO_1487 (O_1487,N_29888,N_29921);
xor UO_1488 (O_1488,N_29824,N_29846);
nand UO_1489 (O_1489,N_29921,N_29926);
xor UO_1490 (O_1490,N_29999,N_29981);
and UO_1491 (O_1491,N_29976,N_29926);
nand UO_1492 (O_1492,N_29870,N_29835);
or UO_1493 (O_1493,N_29875,N_29940);
xor UO_1494 (O_1494,N_29950,N_29963);
or UO_1495 (O_1495,N_29901,N_29806);
xnor UO_1496 (O_1496,N_29861,N_29839);
and UO_1497 (O_1497,N_29800,N_29892);
nor UO_1498 (O_1498,N_29994,N_29979);
nand UO_1499 (O_1499,N_29824,N_29925);
or UO_1500 (O_1500,N_29888,N_29946);
and UO_1501 (O_1501,N_29905,N_29889);
nand UO_1502 (O_1502,N_29895,N_29854);
xor UO_1503 (O_1503,N_29992,N_29893);
or UO_1504 (O_1504,N_29835,N_29986);
or UO_1505 (O_1505,N_29972,N_29955);
xor UO_1506 (O_1506,N_29973,N_29834);
and UO_1507 (O_1507,N_29887,N_29956);
and UO_1508 (O_1508,N_29868,N_29994);
or UO_1509 (O_1509,N_29821,N_29906);
nor UO_1510 (O_1510,N_29843,N_29936);
xnor UO_1511 (O_1511,N_29869,N_29990);
xor UO_1512 (O_1512,N_29913,N_29867);
or UO_1513 (O_1513,N_29901,N_29817);
nor UO_1514 (O_1514,N_29821,N_29946);
nand UO_1515 (O_1515,N_29978,N_29867);
or UO_1516 (O_1516,N_29945,N_29910);
and UO_1517 (O_1517,N_29969,N_29954);
or UO_1518 (O_1518,N_29985,N_29902);
xor UO_1519 (O_1519,N_29968,N_29834);
nor UO_1520 (O_1520,N_29964,N_29865);
xor UO_1521 (O_1521,N_29985,N_29924);
or UO_1522 (O_1522,N_29880,N_29841);
or UO_1523 (O_1523,N_29862,N_29945);
and UO_1524 (O_1524,N_29858,N_29903);
and UO_1525 (O_1525,N_29866,N_29986);
xor UO_1526 (O_1526,N_29861,N_29896);
and UO_1527 (O_1527,N_29825,N_29918);
or UO_1528 (O_1528,N_29944,N_29905);
nand UO_1529 (O_1529,N_29873,N_29848);
nor UO_1530 (O_1530,N_29946,N_29981);
xor UO_1531 (O_1531,N_29825,N_29973);
xnor UO_1532 (O_1532,N_29951,N_29864);
and UO_1533 (O_1533,N_29860,N_29987);
nand UO_1534 (O_1534,N_29845,N_29870);
xnor UO_1535 (O_1535,N_29978,N_29998);
or UO_1536 (O_1536,N_29994,N_29845);
and UO_1537 (O_1537,N_29938,N_29936);
nor UO_1538 (O_1538,N_29911,N_29815);
and UO_1539 (O_1539,N_29832,N_29936);
xor UO_1540 (O_1540,N_29832,N_29888);
or UO_1541 (O_1541,N_29892,N_29923);
nand UO_1542 (O_1542,N_29964,N_29941);
nor UO_1543 (O_1543,N_29842,N_29938);
and UO_1544 (O_1544,N_29859,N_29970);
nor UO_1545 (O_1545,N_29907,N_29882);
nor UO_1546 (O_1546,N_29984,N_29826);
or UO_1547 (O_1547,N_29895,N_29908);
or UO_1548 (O_1548,N_29866,N_29910);
nor UO_1549 (O_1549,N_29808,N_29850);
or UO_1550 (O_1550,N_29829,N_29944);
and UO_1551 (O_1551,N_29942,N_29908);
and UO_1552 (O_1552,N_29900,N_29999);
nor UO_1553 (O_1553,N_29912,N_29852);
nand UO_1554 (O_1554,N_29932,N_29984);
and UO_1555 (O_1555,N_29972,N_29812);
nand UO_1556 (O_1556,N_29861,N_29811);
nand UO_1557 (O_1557,N_29936,N_29968);
nand UO_1558 (O_1558,N_29817,N_29831);
or UO_1559 (O_1559,N_29842,N_29971);
nand UO_1560 (O_1560,N_29950,N_29812);
and UO_1561 (O_1561,N_29980,N_29995);
nor UO_1562 (O_1562,N_29812,N_29855);
nor UO_1563 (O_1563,N_29967,N_29988);
nand UO_1564 (O_1564,N_29841,N_29965);
xnor UO_1565 (O_1565,N_29955,N_29870);
and UO_1566 (O_1566,N_29948,N_29841);
nor UO_1567 (O_1567,N_29869,N_29962);
nor UO_1568 (O_1568,N_29835,N_29941);
or UO_1569 (O_1569,N_29943,N_29966);
and UO_1570 (O_1570,N_29803,N_29908);
nand UO_1571 (O_1571,N_29933,N_29845);
and UO_1572 (O_1572,N_29858,N_29856);
or UO_1573 (O_1573,N_29957,N_29862);
and UO_1574 (O_1574,N_29919,N_29802);
and UO_1575 (O_1575,N_29855,N_29842);
and UO_1576 (O_1576,N_29954,N_29839);
nand UO_1577 (O_1577,N_29855,N_29914);
or UO_1578 (O_1578,N_29962,N_29888);
xor UO_1579 (O_1579,N_29843,N_29998);
nor UO_1580 (O_1580,N_29897,N_29800);
or UO_1581 (O_1581,N_29912,N_29955);
or UO_1582 (O_1582,N_29843,N_29929);
xor UO_1583 (O_1583,N_29833,N_29905);
xor UO_1584 (O_1584,N_29831,N_29949);
and UO_1585 (O_1585,N_29864,N_29997);
or UO_1586 (O_1586,N_29883,N_29956);
nor UO_1587 (O_1587,N_29914,N_29883);
nor UO_1588 (O_1588,N_29933,N_29852);
xnor UO_1589 (O_1589,N_29815,N_29894);
nand UO_1590 (O_1590,N_29913,N_29902);
nor UO_1591 (O_1591,N_29964,N_29990);
nand UO_1592 (O_1592,N_29972,N_29876);
xor UO_1593 (O_1593,N_29928,N_29849);
and UO_1594 (O_1594,N_29906,N_29803);
or UO_1595 (O_1595,N_29903,N_29961);
xnor UO_1596 (O_1596,N_29855,N_29869);
xor UO_1597 (O_1597,N_29857,N_29842);
xnor UO_1598 (O_1598,N_29836,N_29820);
nor UO_1599 (O_1599,N_29986,N_29815);
and UO_1600 (O_1600,N_29959,N_29887);
and UO_1601 (O_1601,N_29912,N_29917);
nor UO_1602 (O_1602,N_29829,N_29801);
or UO_1603 (O_1603,N_29864,N_29975);
nor UO_1604 (O_1604,N_29961,N_29867);
xnor UO_1605 (O_1605,N_29979,N_29800);
xor UO_1606 (O_1606,N_29995,N_29890);
or UO_1607 (O_1607,N_29854,N_29920);
nor UO_1608 (O_1608,N_29876,N_29952);
nand UO_1609 (O_1609,N_29958,N_29974);
nand UO_1610 (O_1610,N_29916,N_29918);
and UO_1611 (O_1611,N_29960,N_29909);
and UO_1612 (O_1612,N_29969,N_29839);
and UO_1613 (O_1613,N_29841,N_29979);
nor UO_1614 (O_1614,N_29814,N_29865);
nor UO_1615 (O_1615,N_29859,N_29989);
nand UO_1616 (O_1616,N_29842,N_29959);
xor UO_1617 (O_1617,N_29884,N_29980);
and UO_1618 (O_1618,N_29935,N_29960);
and UO_1619 (O_1619,N_29987,N_29806);
nand UO_1620 (O_1620,N_29849,N_29843);
nor UO_1621 (O_1621,N_29888,N_29892);
nand UO_1622 (O_1622,N_29965,N_29857);
and UO_1623 (O_1623,N_29878,N_29961);
or UO_1624 (O_1624,N_29807,N_29958);
or UO_1625 (O_1625,N_29907,N_29963);
and UO_1626 (O_1626,N_29985,N_29920);
nor UO_1627 (O_1627,N_29818,N_29934);
xor UO_1628 (O_1628,N_29929,N_29937);
and UO_1629 (O_1629,N_29991,N_29871);
and UO_1630 (O_1630,N_29992,N_29818);
or UO_1631 (O_1631,N_29928,N_29809);
and UO_1632 (O_1632,N_29828,N_29869);
nor UO_1633 (O_1633,N_29962,N_29805);
nor UO_1634 (O_1634,N_29819,N_29812);
xnor UO_1635 (O_1635,N_29868,N_29845);
and UO_1636 (O_1636,N_29898,N_29828);
and UO_1637 (O_1637,N_29862,N_29836);
or UO_1638 (O_1638,N_29942,N_29802);
nand UO_1639 (O_1639,N_29998,N_29814);
nor UO_1640 (O_1640,N_29882,N_29800);
nand UO_1641 (O_1641,N_29840,N_29990);
and UO_1642 (O_1642,N_29832,N_29979);
nand UO_1643 (O_1643,N_29899,N_29832);
nor UO_1644 (O_1644,N_29941,N_29879);
or UO_1645 (O_1645,N_29983,N_29885);
xor UO_1646 (O_1646,N_29816,N_29872);
or UO_1647 (O_1647,N_29835,N_29954);
xor UO_1648 (O_1648,N_29931,N_29869);
and UO_1649 (O_1649,N_29936,N_29811);
or UO_1650 (O_1650,N_29984,N_29929);
and UO_1651 (O_1651,N_29823,N_29879);
and UO_1652 (O_1652,N_29802,N_29990);
or UO_1653 (O_1653,N_29941,N_29850);
nand UO_1654 (O_1654,N_29964,N_29831);
or UO_1655 (O_1655,N_29828,N_29948);
nor UO_1656 (O_1656,N_29828,N_29849);
and UO_1657 (O_1657,N_29800,N_29999);
or UO_1658 (O_1658,N_29857,N_29941);
and UO_1659 (O_1659,N_29814,N_29855);
nand UO_1660 (O_1660,N_29978,N_29973);
or UO_1661 (O_1661,N_29988,N_29994);
nand UO_1662 (O_1662,N_29845,N_29895);
and UO_1663 (O_1663,N_29823,N_29802);
nand UO_1664 (O_1664,N_29927,N_29888);
xnor UO_1665 (O_1665,N_29997,N_29829);
xor UO_1666 (O_1666,N_29819,N_29897);
and UO_1667 (O_1667,N_29982,N_29872);
and UO_1668 (O_1668,N_29924,N_29946);
or UO_1669 (O_1669,N_29810,N_29942);
or UO_1670 (O_1670,N_29807,N_29966);
or UO_1671 (O_1671,N_29800,N_29848);
or UO_1672 (O_1672,N_29810,N_29947);
xor UO_1673 (O_1673,N_29829,N_29921);
nand UO_1674 (O_1674,N_29985,N_29961);
xor UO_1675 (O_1675,N_29997,N_29976);
or UO_1676 (O_1676,N_29982,N_29948);
nor UO_1677 (O_1677,N_29893,N_29935);
and UO_1678 (O_1678,N_29983,N_29941);
nor UO_1679 (O_1679,N_29875,N_29826);
nor UO_1680 (O_1680,N_29807,N_29889);
nand UO_1681 (O_1681,N_29883,N_29866);
nor UO_1682 (O_1682,N_29833,N_29899);
and UO_1683 (O_1683,N_29810,N_29867);
nand UO_1684 (O_1684,N_29916,N_29856);
or UO_1685 (O_1685,N_29987,N_29846);
nand UO_1686 (O_1686,N_29943,N_29809);
nor UO_1687 (O_1687,N_29922,N_29866);
or UO_1688 (O_1688,N_29939,N_29911);
and UO_1689 (O_1689,N_29819,N_29857);
or UO_1690 (O_1690,N_29941,N_29910);
nand UO_1691 (O_1691,N_29966,N_29963);
nor UO_1692 (O_1692,N_29810,N_29987);
nor UO_1693 (O_1693,N_29957,N_29894);
nor UO_1694 (O_1694,N_29810,N_29926);
nor UO_1695 (O_1695,N_29934,N_29966);
and UO_1696 (O_1696,N_29803,N_29994);
nor UO_1697 (O_1697,N_29854,N_29950);
and UO_1698 (O_1698,N_29991,N_29876);
nor UO_1699 (O_1699,N_29906,N_29949);
nand UO_1700 (O_1700,N_29934,N_29831);
nand UO_1701 (O_1701,N_29986,N_29810);
nand UO_1702 (O_1702,N_29950,N_29906);
xnor UO_1703 (O_1703,N_29947,N_29929);
nand UO_1704 (O_1704,N_29888,N_29971);
and UO_1705 (O_1705,N_29985,N_29941);
or UO_1706 (O_1706,N_29822,N_29869);
or UO_1707 (O_1707,N_29907,N_29867);
and UO_1708 (O_1708,N_29920,N_29996);
nor UO_1709 (O_1709,N_29846,N_29939);
or UO_1710 (O_1710,N_29928,N_29990);
and UO_1711 (O_1711,N_29845,N_29969);
or UO_1712 (O_1712,N_29831,N_29946);
nand UO_1713 (O_1713,N_29854,N_29954);
nor UO_1714 (O_1714,N_29912,N_29835);
nand UO_1715 (O_1715,N_29800,N_29960);
xor UO_1716 (O_1716,N_29825,N_29882);
xor UO_1717 (O_1717,N_29809,N_29960);
and UO_1718 (O_1718,N_29908,N_29809);
nand UO_1719 (O_1719,N_29832,N_29831);
xnor UO_1720 (O_1720,N_29869,N_29945);
xor UO_1721 (O_1721,N_29926,N_29903);
nor UO_1722 (O_1722,N_29856,N_29878);
nor UO_1723 (O_1723,N_29934,N_29962);
and UO_1724 (O_1724,N_29983,N_29815);
and UO_1725 (O_1725,N_29926,N_29951);
nand UO_1726 (O_1726,N_29807,N_29848);
xnor UO_1727 (O_1727,N_29829,N_29891);
nor UO_1728 (O_1728,N_29901,N_29894);
and UO_1729 (O_1729,N_29806,N_29969);
nand UO_1730 (O_1730,N_29888,N_29922);
or UO_1731 (O_1731,N_29818,N_29908);
or UO_1732 (O_1732,N_29926,N_29993);
nand UO_1733 (O_1733,N_29984,N_29919);
and UO_1734 (O_1734,N_29819,N_29890);
xnor UO_1735 (O_1735,N_29970,N_29945);
and UO_1736 (O_1736,N_29820,N_29806);
and UO_1737 (O_1737,N_29944,N_29864);
or UO_1738 (O_1738,N_29862,N_29915);
and UO_1739 (O_1739,N_29863,N_29992);
nand UO_1740 (O_1740,N_29908,N_29975);
or UO_1741 (O_1741,N_29827,N_29800);
or UO_1742 (O_1742,N_29809,N_29901);
xnor UO_1743 (O_1743,N_29982,N_29844);
nor UO_1744 (O_1744,N_29915,N_29812);
nand UO_1745 (O_1745,N_29859,N_29975);
nor UO_1746 (O_1746,N_29865,N_29911);
nand UO_1747 (O_1747,N_29991,N_29866);
nor UO_1748 (O_1748,N_29917,N_29930);
nor UO_1749 (O_1749,N_29900,N_29931);
xor UO_1750 (O_1750,N_29856,N_29991);
and UO_1751 (O_1751,N_29872,N_29849);
nor UO_1752 (O_1752,N_29970,N_29887);
nor UO_1753 (O_1753,N_29853,N_29932);
nand UO_1754 (O_1754,N_29920,N_29969);
xor UO_1755 (O_1755,N_29879,N_29877);
nor UO_1756 (O_1756,N_29977,N_29950);
xor UO_1757 (O_1757,N_29949,N_29859);
nor UO_1758 (O_1758,N_29954,N_29923);
or UO_1759 (O_1759,N_29934,N_29999);
or UO_1760 (O_1760,N_29916,N_29978);
xor UO_1761 (O_1761,N_29841,N_29980);
and UO_1762 (O_1762,N_29860,N_29992);
nor UO_1763 (O_1763,N_29955,N_29882);
nand UO_1764 (O_1764,N_29936,N_29901);
nand UO_1765 (O_1765,N_29966,N_29944);
and UO_1766 (O_1766,N_29905,N_29930);
nor UO_1767 (O_1767,N_29936,N_29994);
and UO_1768 (O_1768,N_29971,N_29807);
and UO_1769 (O_1769,N_29947,N_29809);
or UO_1770 (O_1770,N_29977,N_29890);
xnor UO_1771 (O_1771,N_29954,N_29865);
xnor UO_1772 (O_1772,N_29969,N_29897);
or UO_1773 (O_1773,N_29890,N_29932);
and UO_1774 (O_1774,N_29917,N_29914);
or UO_1775 (O_1775,N_29898,N_29806);
xnor UO_1776 (O_1776,N_29898,N_29891);
nand UO_1777 (O_1777,N_29803,N_29982);
or UO_1778 (O_1778,N_29950,N_29841);
nor UO_1779 (O_1779,N_29921,N_29876);
xnor UO_1780 (O_1780,N_29897,N_29905);
nor UO_1781 (O_1781,N_29905,N_29946);
and UO_1782 (O_1782,N_29816,N_29833);
xor UO_1783 (O_1783,N_29958,N_29858);
and UO_1784 (O_1784,N_29998,N_29969);
nand UO_1785 (O_1785,N_29853,N_29979);
nand UO_1786 (O_1786,N_29900,N_29858);
or UO_1787 (O_1787,N_29807,N_29899);
nand UO_1788 (O_1788,N_29845,N_29955);
nor UO_1789 (O_1789,N_29888,N_29830);
xor UO_1790 (O_1790,N_29982,N_29997);
and UO_1791 (O_1791,N_29870,N_29840);
or UO_1792 (O_1792,N_29916,N_29994);
nand UO_1793 (O_1793,N_29817,N_29926);
nand UO_1794 (O_1794,N_29870,N_29943);
nor UO_1795 (O_1795,N_29861,N_29989);
nand UO_1796 (O_1796,N_29848,N_29914);
nand UO_1797 (O_1797,N_29805,N_29919);
and UO_1798 (O_1798,N_29894,N_29859);
nor UO_1799 (O_1799,N_29973,N_29974);
nand UO_1800 (O_1800,N_29809,N_29860);
or UO_1801 (O_1801,N_29918,N_29846);
and UO_1802 (O_1802,N_29885,N_29828);
or UO_1803 (O_1803,N_29922,N_29910);
or UO_1804 (O_1804,N_29900,N_29996);
xnor UO_1805 (O_1805,N_29801,N_29910);
nor UO_1806 (O_1806,N_29869,N_29884);
nand UO_1807 (O_1807,N_29849,N_29899);
xnor UO_1808 (O_1808,N_29950,N_29937);
or UO_1809 (O_1809,N_29862,N_29864);
or UO_1810 (O_1810,N_29944,N_29865);
xor UO_1811 (O_1811,N_29922,N_29882);
or UO_1812 (O_1812,N_29921,N_29960);
xnor UO_1813 (O_1813,N_29818,N_29879);
nor UO_1814 (O_1814,N_29955,N_29983);
or UO_1815 (O_1815,N_29992,N_29951);
nand UO_1816 (O_1816,N_29994,N_29809);
nand UO_1817 (O_1817,N_29897,N_29965);
xnor UO_1818 (O_1818,N_29817,N_29881);
nand UO_1819 (O_1819,N_29898,N_29977);
xor UO_1820 (O_1820,N_29973,N_29914);
or UO_1821 (O_1821,N_29954,N_29812);
xor UO_1822 (O_1822,N_29946,N_29999);
nand UO_1823 (O_1823,N_29857,N_29915);
nor UO_1824 (O_1824,N_29829,N_29971);
and UO_1825 (O_1825,N_29987,N_29992);
nor UO_1826 (O_1826,N_29921,N_29966);
or UO_1827 (O_1827,N_29826,N_29997);
or UO_1828 (O_1828,N_29924,N_29912);
or UO_1829 (O_1829,N_29925,N_29993);
or UO_1830 (O_1830,N_29999,N_29979);
nor UO_1831 (O_1831,N_29953,N_29918);
or UO_1832 (O_1832,N_29878,N_29860);
and UO_1833 (O_1833,N_29933,N_29997);
or UO_1834 (O_1834,N_29943,N_29937);
or UO_1835 (O_1835,N_29923,N_29877);
xnor UO_1836 (O_1836,N_29954,N_29875);
nor UO_1837 (O_1837,N_29997,N_29820);
or UO_1838 (O_1838,N_29936,N_29865);
and UO_1839 (O_1839,N_29940,N_29961);
nand UO_1840 (O_1840,N_29882,N_29841);
and UO_1841 (O_1841,N_29808,N_29928);
nand UO_1842 (O_1842,N_29940,N_29905);
and UO_1843 (O_1843,N_29925,N_29944);
or UO_1844 (O_1844,N_29831,N_29925);
or UO_1845 (O_1845,N_29885,N_29805);
xnor UO_1846 (O_1846,N_29980,N_29954);
xnor UO_1847 (O_1847,N_29864,N_29899);
nand UO_1848 (O_1848,N_29844,N_29926);
and UO_1849 (O_1849,N_29915,N_29804);
nor UO_1850 (O_1850,N_29914,N_29857);
nand UO_1851 (O_1851,N_29941,N_29981);
xor UO_1852 (O_1852,N_29923,N_29958);
xnor UO_1853 (O_1853,N_29967,N_29946);
xor UO_1854 (O_1854,N_29802,N_29815);
xnor UO_1855 (O_1855,N_29897,N_29890);
or UO_1856 (O_1856,N_29956,N_29893);
nor UO_1857 (O_1857,N_29979,N_29801);
or UO_1858 (O_1858,N_29982,N_29969);
or UO_1859 (O_1859,N_29895,N_29968);
xnor UO_1860 (O_1860,N_29865,N_29826);
or UO_1861 (O_1861,N_29848,N_29925);
xnor UO_1862 (O_1862,N_29905,N_29838);
xor UO_1863 (O_1863,N_29853,N_29906);
nor UO_1864 (O_1864,N_29845,N_29982);
nand UO_1865 (O_1865,N_29813,N_29913);
or UO_1866 (O_1866,N_29910,N_29885);
and UO_1867 (O_1867,N_29876,N_29857);
nor UO_1868 (O_1868,N_29856,N_29870);
xnor UO_1869 (O_1869,N_29972,N_29969);
nand UO_1870 (O_1870,N_29977,N_29943);
and UO_1871 (O_1871,N_29958,N_29938);
xnor UO_1872 (O_1872,N_29876,N_29966);
or UO_1873 (O_1873,N_29963,N_29810);
and UO_1874 (O_1874,N_29911,N_29801);
and UO_1875 (O_1875,N_29829,N_29967);
or UO_1876 (O_1876,N_29942,N_29892);
or UO_1877 (O_1877,N_29956,N_29969);
and UO_1878 (O_1878,N_29969,N_29922);
or UO_1879 (O_1879,N_29981,N_29802);
nand UO_1880 (O_1880,N_29947,N_29932);
or UO_1881 (O_1881,N_29964,N_29851);
or UO_1882 (O_1882,N_29916,N_29828);
and UO_1883 (O_1883,N_29940,N_29852);
xor UO_1884 (O_1884,N_29952,N_29954);
and UO_1885 (O_1885,N_29956,N_29851);
nor UO_1886 (O_1886,N_29938,N_29994);
or UO_1887 (O_1887,N_29932,N_29991);
nor UO_1888 (O_1888,N_29951,N_29976);
or UO_1889 (O_1889,N_29835,N_29959);
and UO_1890 (O_1890,N_29923,N_29883);
and UO_1891 (O_1891,N_29823,N_29847);
and UO_1892 (O_1892,N_29846,N_29915);
nand UO_1893 (O_1893,N_29888,N_29810);
and UO_1894 (O_1894,N_29887,N_29802);
and UO_1895 (O_1895,N_29915,N_29840);
nor UO_1896 (O_1896,N_29894,N_29808);
or UO_1897 (O_1897,N_29829,N_29892);
xnor UO_1898 (O_1898,N_29990,N_29895);
xnor UO_1899 (O_1899,N_29996,N_29885);
xor UO_1900 (O_1900,N_29991,N_29875);
xor UO_1901 (O_1901,N_29891,N_29808);
nand UO_1902 (O_1902,N_29966,N_29802);
nand UO_1903 (O_1903,N_29987,N_29866);
xor UO_1904 (O_1904,N_29980,N_29848);
and UO_1905 (O_1905,N_29938,N_29902);
or UO_1906 (O_1906,N_29859,N_29809);
nand UO_1907 (O_1907,N_29993,N_29831);
xor UO_1908 (O_1908,N_29807,N_29840);
nand UO_1909 (O_1909,N_29847,N_29970);
nor UO_1910 (O_1910,N_29820,N_29980);
xnor UO_1911 (O_1911,N_29951,N_29821);
xor UO_1912 (O_1912,N_29956,N_29987);
xor UO_1913 (O_1913,N_29970,N_29921);
xor UO_1914 (O_1914,N_29924,N_29842);
nand UO_1915 (O_1915,N_29806,N_29978);
nor UO_1916 (O_1916,N_29898,N_29933);
and UO_1917 (O_1917,N_29951,N_29983);
nor UO_1918 (O_1918,N_29845,N_29855);
and UO_1919 (O_1919,N_29983,N_29888);
xor UO_1920 (O_1920,N_29818,N_29839);
or UO_1921 (O_1921,N_29942,N_29958);
and UO_1922 (O_1922,N_29965,N_29864);
xnor UO_1923 (O_1923,N_29940,N_29827);
or UO_1924 (O_1924,N_29968,N_29833);
nand UO_1925 (O_1925,N_29921,N_29825);
and UO_1926 (O_1926,N_29988,N_29935);
or UO_1927 (O_1927,N_29853,N_29867);
or UO_1928 (O_1928,N_29808,N_29811);
nand UO_1929 (O_1929,N_29843,N_29818);
nand UO_1930 (O_1930,N_29898,N_29967);
xnor UO_1931 (O_1931,N_29946,N_29972);
or UO_1932 (O_1932,N_29965,N_29974);
nor UO_1933 (O_1933,N_29929,N_29811);
nand UO_1934 (O_1934,N_29866,N_29998);
nor UO_1935 (O_1935,N_29893,N_29880);
or UO_1936 (O_1936,N_29854,N_29897);
nand UO_1937 (O_1937,N_29845,N_29996);
nor UO_1938 (O_1938,N_29976,N_29846);
or UO_1939 (O_1939,N_29915,N_29983);
nor UO_1940 (O_1940,N_29822,N_29887);
or UO_1941 (O_1941,N_29876,N_29894);
and UO_1942 (O_1942,N_29939,N_29822);
nor UO_1943 (O_1943,N_29961,N_29927);
nand UO_1944 (O_1944,N_29916,N_29906);
nor UO_1945 (O_1945,N_29962,N_29897);
and UO_1946 (O_1946,N_29865,N_29965);
nor UO_1947 (O_1947,N_29843,N_29908);
and UO_1948 (O_1948,N_29922,N_29848);
xnor UO_1949 (O_1949,N_29989,N_29822);
and UO_1950 (O_1950,N_29808,N_29939);
nand UO_1951 (O_1951,N_29810,N_29948);
and UO_1952 (O_1952,N_29858,N_29831);
xnor UO_1953 (O_1953,N_29984,N_29938);
xor UO_1954 (O_1954,N_29814,N_29808);
nor UO_1955 (O_1955,N_29890,N_29919);
xnor UO_1956 (O_1956,N_29921,N_29850);
and UO_1957 (O_1957,N_29813,N_29983);
nor UO_1958 (O_1958,N_29838,N_29957);
nand UO_1959 (O_1959,N_29870,N_29993);
nand UO_1960 (O_1960,N_29994,N_29852);
nand UO_1961 (O_1961,N_29950,N_29814);
and UO_1962 (O_1962,N_29809,N_29839);
or UO_1963 (O_1963,N_29885,N_29819);
and UO_1964 (O_1964,N_29899,N_29973);
nand UO_1965 (O_1965,N_29942,N_29944);
nor UO_1966 (O_1966,N_29948,N_29825);
xnor UO_1967 (O_1967,N_29973,N_29814);
xor UO_1968 (O_1968,N_29867,N_29983);
and UO_1969 (O_1969,N_29826,N_29817);
nand UO_1970 (O_1970,N_29832,N_29946);
xor UO_1971 (O_1971,N_29813,N_29859);
nand UO_1972 (O_1972,N_29872,N_29899);
or UO_1973 (O_1973,N_29950,N_29916);
nand UO_1974 (O_1974,N_29836,N_29976);
or UO_1975 (O_1975,N_29887,N_29833);
nand UO_1976 (O_1976,N_29852,N_29981);
or UO_1977 (O_1977,N_29922,N_29992);
nor UO_1978 (O_1978,N_29963,N_29875);
nand UO_1979 (O_1979,N_29872,N_29905);
xor UO_1980 (O_1980,N_29846,N_29994);
or UO_1981 (O_1981,N_29929,N_29879);
xor UO_1982 (O_1982,N_29885,N_29896);
nor UO_1983 (O_1983,N_29838,N_29913);
nand UO_1984 (O_1984,N_29902,N_29963);
nor UO_1985 (O_1985,N_29897,N_29828);
or UO_1986 (O_1986,N_29919,N_29824);
nand UO_1987 (O_1987,N_29962,N_29942);
or UO_1988 (O_1988,N_29916,N_29904);
nor UO_1989 (O_1989,N_29819,N_29831);
and UO_1990 (O_1990,N_29831,N_29801);
and UO_1991 (O_1991,N_29841,N_29969);
or UO_1992 (O_1992,N_29888,N_29843);
or UO_1993 (O_1993,N_29893,N_29821);
or UO_1994 (O_1994,N_29921,N_29917);
nand UO_1995 (O_1995,N_29847,N_29941);
and UO_1996 (O_1996,N_29838,N_29919);
nor UO_1997 (O_1997,N_29818,N_29851);
and UO_1998 (O_1998,N_29872,N_29959);
and UO_1999 (O_1999,N_29863,N_29872);
or UO_2000 (O_2000,N_29826,N_29998);
xor UO_2001 (O_2001,N_29814,N_29825);
xor UO_2002 (O_2002,N_29827,N_29893);
nand UO_2003 (O_2003,N_29997,N_29967);
nor UO_2004 (O_2004,N_29842,N_29827);
nor UO_2005 (O_2005,N_29960,N_29915);
nor UO_2006 (O_2006,N_29930,N_29887);
xnor UO_2007 (O_2007,N_29859,N_29865);
nand UO_2008 (O_2008,N_29864,N_29898);
or UO_2009 (O_2009,N_29844,N_29854);
xor UO_2010 (O_2010,N_29972,N_29850);
xor UO_2011 (O_2011,N_29848,N_29871);
or UO_2012 (O_2012,N_29910,N_29816);
nor UO_2013 (O_2013,N_29942,N_29833);
and UO_2014 (O_2014,N_29933,N_29821);
nor UO_2015 (O_2015,N_29863,N_29883);
and UO_2016 (O_2016,N_29939,N_29987);
or UO_2017 (O_2017,N_29936,N_29959);
nor UO_2018 (O_2018,N_29927,N_29843);
nor UO_2019 (O_2019,N_29888,N_29811);
xor UO_2020 (O_2020,N_29816,N_29853);
xnor UO_2021 (O_2021,N_29963,N_29989);
nand UO_2022 (O_2022,N_29839,N_29805);
nand UO_2023 (O_2023,N_29920,N_29814);
nor UO_2024 (O_2024,N_29808,N_29856);
or UO_2025 (O_2025,N_29862,N_29865);
nor UO_2026 (O_2026,N_29990,N_29845);
or UO_2027 (O_2027,N_29914,N_29841);
xor UO_2028 (O_2028,N_29814,N_29888);
nand UO_2029 (O_2029,N_29857,N_29939);
nand UO_2030 (O_2030,N_29968,N_29821);
or UO_2031 (O_2031,N_29809,N_29962);
nor UO_2032 (O_2032,N_29878,N_29822);
nor UO_2033 (O_2033,N_29804,N_29946);
nand UO_2034 (O_2034,N_29830,N_29902);
nor UO_2035 (O_2035,N_29955,N_29823);
nor UO_2036 (O_2036,N_29941,N_29819);
nor UO_2037 (O_2037,N_29917,N_29875);
nand UO_2038 (O_2038,N_29888,N_29968);
nand UO_2039 (O_2039,N_29872,N_29886);
nor UO_2040 (O_2040,N_29927,N_29874);
nor UO_2041 (O_2041,N_29820,N_29947);
xor UO_2042 (O_2042,N_29832,N_29821);
or UO_2043 (O_2043,N_29972,N_29918);
nand UO_2044 (O_2044,N_29992,N_29991);
and UO_2045 (O_2045,N_29887,N_29820);
nor UO_2046 (O_2046,N_29988,N_29837);
and UO_2047 (O_2047,N_29800,N_29814);
nand UO_2048 (O_2048,N_29828,N_29876);
xor UO_2049 (O_2049,N_29948,N_29972);
or UO_2050 (O_2050,N_29856,N_29898);
xnor UO_2051 (O_2051,N_29905,N_29978);
xnor UO_2052 (O_2052,N_29946,N_29846);
xnor UO_2053 (O_2053,N_29839,N_29856);
or UO_2054 (O_2054,N_29941,N_29997);
or UO_2055 (O_2055,N_29807,N_29885);
nor UO_2056 (O_2056,N_29999,N_29815);
or UO_2057 (O_2057,N_29833,N_29902);
xnor UO_2058 (O_2058,N_29872,N_29834);
nor UO_2059 (O_2059,N_29822,N_29853);
and UO_2060 (O_2060,N_29953,N_29842);
and UO_2061 (O_2061,N_29867,N_29953);
or UO_2062 (O_2062,N_29839,N_29801);
and UO_2063 (O_2063,N_29864,N_29869);
xnor UO_2064 (O_2064,N_29929,N_29998);
and UO_2065 (O_2065,N_29808,N_29825);
nor UO_2066 (O_2066,N_29814,N_29832);
xor UO_2067 (O_2067,N_29955,N_29927);
xnor UO_2068 (O_2068,N_29971,N_29961);
xnor UO_2069 (O_2069,N_29981,N_29996);
nand UO_2070 (O_2070,N_29842,N_29919);
xor UO_2071 (O_2071,N_29970,N_29842);
and UO_2072 (O_2072,N_29882,N_29815);
xnor UO_2073 (O_2073,N_29957,N_29930);
nand UO_2074 (O_2074,N_29820,N_29813);
or UO_2075 (O_2075,N_29932,N_29907);
nor UO_2076 (O_2076,N_29935,N_29933);
and UO_2077 (O_2077,N_29810,N_29932);
nand UO_2078 (O_2078,N_29820,N_29925);
nor UO_2079 (O_2079,N_29871,N_29833);
or UO_2080 (O_2080,N_29886,N_29875);
or UO_2081 (O_2081,N_29899,N_29857);
nor UO_2082 (O_2082,N_29811,N_29972);
xor UO_2083 (O_2083,N_29891,N_29943);
or UO_2084 (O_2084,N_29819,N_29874);
xor UO_2085 (O_2085,N_29871,N_29902);
xnor UO_2086 (O_2086,N_29903,N_29834);
xnor UO_2087 (O_2087,N_29890,N_29800);
nor UO_2088 (O_2088,N_29853,N_29980);
nor UO_2089 (O_2089,N_29963,N_29850);
nor UO_2090 (O_2090,N_29872,N_29975);
nand UO_2091 (O_2091,N_29959,N_29818);
nor UO_2092 (O_2092,N_29966,N_29917);
and UO_2093 (O_2093,N_29945,N_29878);
nand UO_2094 (O_2094,N_29811,N_29859);
nand UO_2095 (O_2095,N_29861,N_29922);
nor UO_2096 (O_2096,N_29835,N_29950);
nand UO_2097 (O_2097,N_29802,N_29860);
or UO_2098 (O_2098,N_29854,N_29880);
nand UO_2099 (O_2099,N_29811,N_29911);
nor UO_2100 (O_2100,N_29846,N_29843);
or UO_2101 (O_2101,N_29857,N_29828);
or UO_2102 (O_2102,N_29858,N_29951);
or UO_2103 (O_2103,N_29908,N_29829);
nand UO_2104 (O_2104,N_29850,N_29896);
nor UO_2105 (O_2105,N_29849,N_29948);
nor UO_2106 (O_2106,N_29945,N_29941);
and UO_2107 (O_2107,N_29858,N_29801);
nor UO_2108 (O_2108,N_29829,N_29946);
xor UO_2109 (O_2109,N_29900,N_29924);
or UO_2110 (O_2110,N_29975,N_29876);
or UO_2111 (O_2111,N_29976,N_29941);
or UO_2112 (O_2112,N_29969,N_29816);
nand UO_2113 (O_2113,N_29862,N_29822);
xor UO_2114 (O_2114,N_29924,N_29878);
or UO_2115 (O_2115,N_29893,N_29872);
nor UO_2116 (O_2116,N_29995,N_29841);
and UO_2117 (O_2117,N_29837,N_29800);
or UO_2118 (O_2118,N_29890,N_29900);
or UO_2119 (O_2119,N_29960,N_29979);
or UO_2120 (O_2120,N_29895,N_29917);
or UO_2121 (O_2121,N_29824,N_29974);
xor UO_2122 (O_2122,N_29868,N_29816);
nand UO_2123 (O_2123,N_29845,N_29946);
nand UO_2124 (O_2124,N_29808,N_29961);
nand UO_2125 (O_2125,N_29820,N_29837);
or UO_2126 (O_2126,N_29828,N_29911);
and UO_2127 (O_2127,N_29966,N_29941);
nand UO_2128 (O_2128,N_29994,N_29824);
nor UO_2129 (O_2129,N_29986,N_29836);
nand UO_2130 (O_2130,N_29960,N_29899);
and UO_2131 (O_2131,N_29935,N_29846);
nor UO_2132 (O_2132,N_29875,N_29914);
xor UO_2133 (O_2133,N_29995,N_29940);
xor UO_2134 (O_2134,N_29953,N_29995);
nor UO_2135 (O_2135,N_29863,N_29830);
nor UO_2136 (O_2136,N_29908,N_29815);
nand UO_2137 (O_2137,N_29933,N_29963);
or UO_2138 (O_2138,N_29906,N_29910);
nand UO_2139 (O_2139,N_29902,N_29964);
xor UO_2140 (O_2140,N_29877,N_29917);
nand UO_2141 (O_2141,N_29932,N_29840);
and UO_2142 (O_2142,N_29916,N_29838);
or UO_2143 (O_2143,N_29991,N_29869);
xor UO_2144 (O_2144,N_29899,N_29867);
or UO_2145 (O_2145,N_29893,N_29972);
and UO_2146 (O_2146,N_29941,N_29969);
or UO_2147 (O_2147,N_29971,N_29896);
or UO_2148 (O_2148,N_29936,N_29831);
nor UO_2149 (O_2149,N_29920,N_29891);
xnor UO_2150 (O_2150,N_29901,N_29896);
xor UO_2151 (O_2151,N_29912,N_29990);
nand UO_2152 (O_2152,N_29929,N_29800);
nor UO_2153 (O_2153,N_29895,N_29927);
and UO_2154 (O_2154,N_29826,N_29903);
nor UO_2155 (O_2155,N_29882,N_29829);
xnor UO_2156 (O_2156,N_29854,N_29834);
or UO_2157 (O_2157,N_29820,N_29920);
nor UO_2158 (O_2158,N_29829,N_29896);
nand UO_2159 (O_2159,N_29960,N_29898);
nand UO_2160 (O_2160,N_29968,N_29816);
nand UO_2161 (O_2161,N_29855,N_29919);
and UO_2162 (O_2162,N_29914,N_29939);
xor UO_2163 (O_2163,N_29935,N_29958);
or UO_2164 (O_2164,N_29870,N_29844);
or UO_2165 (O_2165,N_29800,N_29846);
and UO_2166 (O_2166,N_29898,N_29971);
xnor UO_2167 (O_2167,N_29818,N_29866);
and UO_2168 (O_2168,N_29829,N_29863);
nand UO_2169 (O_2169,N_29866,N_29861);
or UO_2170 (O_2170,N_29983,N_29881);
or UO_2171 (O_2171,N_29832,N_29851);
xor UO_2172 (O_2172,N_29883,N_29920);
nand UO_2173 (O_2173,N_29868,N_29834);
xor UO_2174 (O_2174,N_29941,N_29938);
and UO_2175 (O_2175,N_29959,N_29878);
nor UO_2176 (O_2176,N_29892,N_29840);
nor UO_2177 (O_2177,N_29823,N_29894);
xor UO_2178 (O_2178,N_29859,N_29941);
or UO_2179 (O_2179,N_29952,N_29814);
and UO_2180 (O_2180,N_29895,N_29918);
and UO_2181 (O_2181,N_29857,N_29980);
xnor UO_2182 (O_2182,N_29988,N_29958);
xnor UO_2183 (O_2183,N_29977,N_29940);
nand UO_2184 (O_2184,N_29960,N_29818);
xor UO_2185 (O_2185,N_29830,N_29912);
or UO_2186 (O_2186,N_29934,N_29923);
xor UO_2187 (O_2187,N_29815,N_29852);
or UO_2188 (O_2188,N_29831,N_29991);
and UO_2189 (O_2189,N_29829,N_29819);
nor UO_2190 (O_2190,N_29935,N_29864);
xnor UO_2191 (O_2191,N_29986,N_29937);
or UO_2192 (O_2192,N_29955,N_29843);
nand UO_2193 (O_2193,N_29879,N_29915);
nand UO_2194 (O_2194,N_29819,N_29865);
xor UO_2195 (O_2195,N_29920,N_29881);
or UO_2196 (O_2196,N_29805,N_29974);
nand UO_2197 (O_2197,N_29956,N_29814);
xor UO_2198 (O_2198,N_29873,N_29929);
xor UO_2199 (O_2199,N_29902,N_29947);
and UO_2200 (O_2200,N_29922,N_29995);
and UO_2201 (O_2201,N_29994,N_29821);
nand UO_2202 (O_2202,N_29978,N_29832);
xnor UO_2203 (O_2203,N_29925,N_29962);
or UO_2204 (O_2204,N_29940,N_29896);
or UO_2205 (O_2205,N_29931,N_29849);
xnor UO_2206 (O_2206,N_29957,N_29964);
or UO_2207 (O_2207,N_29827,N_29975);
nor UO_2208 (O_2208,N_29859,N_29973);
nor UO_2209 (O_2209,N_29806,N_29811);
and UO_2210 (O_2210,N_29901,N_29887);
nand UO_2211 (O_2211,N_29861,N_29801);
nor UO_2212 (O_2212,N_29932,N_29985);
nor UO_2213 (O_2213,N_29948,N_29970);
or UO_2214 (O_2214,N_29828,N_29800);
and UO_2215 (O_2215,N_29819,N_29855);
nand UO_2216 (O_2216,N_29817,N_29958);
and UO_2217 (O_2217,N_29927,N_29803);
and UO_2218 (O_2218,N_29933,N_29945);
nor UO_2219 (O_2219,N_29894,N_29912);
or UO_2220 (O_2220,N_29928,N_29964);
or UO_2221 (O_2221,N_29947,N_29998);
nor UO_2222 (O_2222,N_29925,N_29915);
and UO_2223 (O_2223,N_29833,N_29862);
nor UO_2224 (O_2224,N_29892,N_29965);
xnor UO_2225 (O_2225,N_29837,N_29840);
and UO_2226 (O_2226,N_29909,N_29916);
or UO_2227 (O_2227,N_29994,N_29874);
or UO_2228 (O_2228,N_29813,N_29830);
nor UO_2229 (O_2229,N_29900,N_29853);
nor UO_2230 (O_2230,N_29859,N_29871);
xor UO_2231 (O_2231,N_29823,N_29953);
and UO_2232 (O_2232,N_29846,N_29884);
nor UO_2233 (O_2233,N_29990,N_29860);
nand UO_2234 (O_2234,N_29913,N_29899);
xor UO_2235 (O_2235,N_29820,N_29934);
or UO_2236 (O_2236,N_29919,N_29954);
nor UO_2237 (O_2237,N_29856,N_29968);
nand UO_2238 (O_2238,N_29900,N_29860);
nand UO_2239 (O_2239,N_29909,N_29912);
nand UO_2240 (O_2240,N_29899,N_29977);
or UO_2241 (O_2241,N_29927,N_29970);
nand UO_2242 (O_2242,N_29955,N_29897);
nor UO_2243 (O_2243,N_29985,N_29933);
nand UO_2244 (O_2244,N_29961,N_29890);
and UO_2245 (O_2245,N_29887,N_29996);
and UO_2246 (O_2246,N_29926,N_29838);
or UO_2247 (O_2247,N_29922,N_29916);
xnor UO_2248 (O_2248,N_29910,N_29824);
nand UO_2249 (O_2249,N_29870,N_29852);
and UO_2250 (O_2250,N_29912,N_29831);
xnor UO_2251 (O_2251,N_29889,N_29925);
nor UO_2252 (O_2252,N_29938,N_29970);
or UO_2253 (O_2253,N_29930,N_29953);
nor UO_2254 (O_2254,N_29885,N_29878);
nand UO_2255 (O_2255,N_29961,N_29941);
nand UO_2256 (O_2256,N_29877,N_29810);
nor UO_2257 (O_2257,N_29970,N_29870);
nor UO_2258 (O_2258,N_29974,N_29819);
nand UO_2259 (O_2259,N_29963,N_29848);
nor UO_2260 (O_2260,N_29841,N_29927);
or UO_2261 (O_2261,N_29925,N_29869);
or UO_2262 (O_2262,N_29844,N_29878);
and UO_2263 (O_2263,N_29985,N_29947);
or UO_2264 (O_2264,N_29899,N_29875);
and UO_2265 (O_2265,N_29976,N_29865);
and UO_2266 (O_2266,N_29878,N_29893);
xor UO_2267 (O_2267,N_29868,N_29906);
or UO_2268 (O_2268,N_29981,N_29987);
xnor UO_2269 (O_2269,N_29915,N_29908);
xnor UO_2270 (O_2270,N_29922,N_29968);
nand UO_2271 (O_2271,N_29961,N_29960);
xnor UO_2272 (O_2272,N_29868,N_29809);
or UO_2273 (O_2273,N_29924,N_29826);
nor UO_2274 (O_2274,N_29933,N_29989);
nor UO_2275 (O_2275,N_29884,N_29850);
xor UO_2276 (O_2276,N_29871,N_29816);
xnor UO_2277 (O_2277,N_29812,N_29965);
and UO_2278 (O_2278,N_29941,N_29948);
and UO_2279 (O_2279,N_29802,N_29888);
xor UO_2280 (O_2280,N_29928,N_29916);
nor UO_2281 (O_2281,N_29893,N_29985);
nand UO_2282 (O_2282,N_29934,N_29894);
and UO_2283 (O_2283,N_29896,N_29873);
and UO_2284 (O_2284,N_29851,N_29949);
xnor UO_2285 (O_2285,N_29964,N_29806);
xnor UO_2286 (O_2286,N_29982,N_29850);
xnor UO_2287 (O_2287,N_29968,N_29889);
and UO_2288 (O_2288,N_29911,N_29827);
nand UO_2289 (O_2289,N_29833,N_29801);
and UO_2290 (O_2290,N_29993,N_29859);
or UO_2291 (O_2291,N_29860,N_29805);
nand UO_2292 (O_2292,N_29958,N_29852);
xor UO_2293 (O_2293,N_29941,N_29955);
nand UO_2294 (O_2294,N_29983,N_29863);
and UO_2295 (O_2295,N_29944,N_29913);
nor UO_2296 (O_2296,N_29884,N_29845);
or UO_2297 (O_2297,N_29891,N_29925);
and UO_2298 (O_2298,N_29856,N_29926);
or UO_2299 (O_2299,N_29888,N_29974);
or UO_2300 (O_2300,N_29816,N_29869);
and UO_2301 (O_2301,N_29807,N_29993);
nand UO_2302 (O_2302,N_29965,N_29848);
or UO_2303 (O_2303,N_29883,N_29993);
or UO_2304 (O_2304,N_29898,N_29917);
or UO_2305 (O_2305,N_29924,N_29875);
and UO_2306 (O_2306,N_29943,N_29895);
and UO_2307 (O_2307,N_29987,N_29979);
nor UO_2308 (O_2308,N_29830,N_29998);
nor UO_2309 (O_2309,N_29981,N_29828);
nor UO_2310 (O_2310,N_29860,N_29924);
xnor UO_2311 (O_2311,N_29931,N_29817);
nand UO_2312 (O_2312,N_29925,N_29919);
xnor UO_2313 (O_2313,N_29840,N_29956);
or UO_2314 (O_2314,N_29957,N_29819);
and UO_2315 (O_2315,N_29838,N_29814);
xnor UO_2316 (O_2316,N_29842,N_29891);
xnor UO_2317 (O_2317,N_29977,N_29891);
nand UO_2318 (O_2318,N_29858,N_29844);
nand UO_2319 (O_2319,N_29966,N_29908);
and UO_2320 (O_2320,N_29853,N_29869);
nand UO_2321 (O_2321,N_29963,N_29853);
and UO_2322 (O_2322,N_29923,N_29967);
or UO_2323 (O_2323,N_29955,N_29945);
or UO_2324 (O_2324,N_29950,N_29840);
or UO_2325 (O_2325,N_29987,N_29969);
or UO_2326 (O_2326,N_29816,N_29984);
nand UO_2327 (O_2327,N_29818,N_29935);
nor UO_2328 (O_2328,N_29945,N_29953);
or UO_2329 (O_2329,N_29841,N_29945);
xor UO_2330 (O_2330,N_29918,N_29814);
xor UO_2331 (O_2331,N_29996,N_29803);
or UO_2332 (O_2332,N_29963,N_29914);
nand UO_2333 (O_2333,N_29853,N_29961);
xor UO_2334 (O_2334,N_29910,N_29902);
nor UO_2335 (O_2335,N_29998,N_29860);
nor UO_2336 (O_2336,N_29979,N_29846);
or UO_2337 (O_2337,N_29925,N_29822);
nor UO_2338 (O_2338,N_29807,N_29831);
and UO_2339 (O_2339,N_29976,N_29855);
xnor UO_2340 (O_2340,N_29908,N_29819);
or UO_2341 (O_2341,N_29870,N_29968);
or UO_2342 (O_2342,N_29879,N_29839);
or UO_2343 (O_2343,N_29964,N_29976);
xnor UO_2344 (O_2344,N_29816,N_29832);
nand UO_2345 (O_2345,N_29998,N_29831);
nor UO_2346 (O_2346,N_29841,N_29886);
nor UO_2347 (O_2347,N_29800,N_29941);
or UO_2348 (O_2348,N_29866,N_29893);
and UO_2349 (O_2349,N_29925,N_29886);
nand UO_2350 (O_2350,N_29842,N_29860);
xnor UO_2351 (O_2351,N_29993,N_29981);
and UO_2352 (O_2352,N_29825,N_29826);
xnor UO_2353 (O_2353,N_29825,N_29898);
or UO_2354 (O_2354,N_29906,N_29872);
xor UO_2355 (O_2355,N_29944,N_29811);
nor UO_2356 (O_2356,N_29940,N_29803);
xor UO_2357 (O_2357,N_29961,N_29919);
nor UO_2358 (O_2358,N_29970,N_29902);
xnor UO_2359 (O_2359,N_29955,N_29846);
xnor UO_2360 (O_2360,N_29911,N_29904);
nor UO_2361 (O_2361,N_29827,N_29815);
nor UO_2362 (O_2362,N_29887,N_29980);
xnor UO_2363 (O_2363,N_29961,N_29885);
nor UO_2364 (O_2364,N_29995,N_29852);
nor UO_2365 (O_2365,N_29873,N_29838);
nand UO_2366 (O_2366,N_29946,N_29973);
or UO_2367 (O_2367,N_29915,N_29956);
or UO_2368 (O_2368,N_29949,N_29897);
and UO_2369 (O_2369,N_29970,N_29918);
xor UO_2370 (O_2370,N_29889,N_29833);
or UO_2371 (O_2371,N_29926,N_29963);
and UO_2372 (O_2372,N_29900,N_29935);
or UO_2373 (O_2373,N_29954,N_29953);
and UO_2374 (O_2374,N_29827,N_29997);
nor UO_2375 (O_2375,N_29867,N_29991);
nand UO_2376 (O_2376,N_29936,N_29858);
or UO_2377 (O_2377,N_29978,N_29970);
nand UO_2378 (O_2378,N_29956,N_29827);
or UO_2379 (O_2379,N_29859,N_29843);
or UO_2380 (O_2380,N_29887,N_29895);
nand UO_2381 (O_2381,N_29936,N_29890);
or UO_2382 (O_2382,N_29801,N_29943);
and UO_2383 (O_2383,N_29832,N_29951);
xnor UO_2384 (O_2384,N_29931,N_29822);
xnor UO_2385 (O_2385,N_29969,N_29831);
nand UO_2386 (O_2386,N_29969,N_29871);
and UO_2387 (O_2387,N_29973,N_29818);
nor UO_2388 (O_2388,N_29913,N_29892);
or UO_2389 (O_2389,N_29981,N_29975);
nor UO_2390 (O_2390,N_29917,N_29997);
and UO_2391 (O_2391,N_29945,N_29881);
nor UO_2392 (O_2392,N_29914,N_29965);
xnor UO_2393 (O_2393,N_29842,N_29873);
or UO_2394 (O_2394,N_29963,N_29808);
nor UO_2395 (O_2395,N_29878,N_29965);
nor UO_2396 (O_2396,N_29897,N_29967);
or UO_2397 (O_2397,N_29905,N_29990);
nand UO_2398 (O_2398,N_29994,N_29920);
nor UO_2399 (O_2399,N_29826,N_29890);
and UO_2400 (O_2400,N_29898,N_29857);
nand UO_2401 (O_2401,N_29965,N_29819);
nand UO_2402 (O_2402,N_29959,N_29855);
and UO_2403 (O_2403,N_29870,N_29865);
nor UO_2404 (O_2404,N_29886,N_29946);
xor UO_2405 (O_2405,N_29807,N_29866);
and UO_2406 (O_2406,N_29819,N_29981);
nor UO_2407 (O_2407,N_29863,N_29965);
nor UO_2408 (O_2408,N_29874,N_29804);
or UO_2409 (O_2409,N_29881,N_29804);
nand UO_2410 (O_2410,N_29835,N_29869);
or UO_2411 (O_2411,N_29907,N_29840);
nor UO_2412 (O_2412,N_29902,N_29958);
nand UO_2413 (O_2413,N_29949,N_29958);
nand UO_2414 (O_2414,N_29905,N_29863);
nand UO_2415 (O_2415,N_29859,N_29812);
and UO_2416 (O_2416,N_29823,N_29881);
nand UO_2417 (O_2417,N_29895,N_29830);
xnor UO_2418 (O_2418,N_29865,N_29955);
nand UO_2419 (O_2419,N_29833,N_29935);
or UO_2420 (O_2420,N_29968,N_29931);
and UO_2421 (O_2421,N_29944,N_29974);
and UO_2422 (O_2422,N_29823,N_29951);
xnor UO_2423 (O_2423,N_29959,N_29888);
xor UO_2424 (O_2424,N_29818,N_29849);
nand UO_2425 (O_2425,N_29861,N_29910);
nor UO_2426 (O_2426,N_29835,N_29803);
or UO_2427 (O_2427,N_29823,N_29995);
or UO_2428 (O_2428,N_29996,N_29961);
nor UO_2429 (O_2429,N_29887,N_29923);
and UO_2430 (O_2430,N_29964,N_29885);
or UO_2431 (O_2431,N_29906,N_29956);
xnor UO_2432 (O_2432,N_29905,N_29805);
or UO_2433 (O_2433,N_29938,N_29889);
nand UO_2434 (O_2434,N_29955,N_29886);
nor UO_2435 (O_2435,N_29851,N_29806);
xnor UO_2436 (O_2436,N_29902,N_29975);
and UO_2437 (O_2437,N_29900,N_29894);
nand UO_2438 (O_2438,N_29936,N_29869);
nor UO_2439 (O_2439,N_29854,N_29948);
xnor UO_2440 (O_2440,N_29884,N_29856);
nand UO_2441 (O_2441,N_29890,N_29845);
and UO_2442 (O_2442,N_29907,N_29919);
xor UO_2443 (O_2443,N_29908,N_29814);
nand UO_2444 (O_2444,N_29868,N_29806);
nand UO_2445 (O_2445,N_29827,N_29932);
or UO_2446 (O_2446,N_29912,N_29941);
xnor UO_2447 (O_2447,N_29927,N_29892);
xor UO_2448 (O_2448,N_29973,N_29957);
or UO_2449 (O_2449,N_29809,N_29953);
xnor UO_2450 (O_2450,N_29809,N_29939);
nor UO_2451 (O_2451,N_29941,N_29954);
xnor UO_2452 (O_2452,N_29901,N_29855);
nand UO_2453 (O_2453,N_29851,N_29936);
and UO_2454 (O_2454,N_29834,N_29991);
nor UO_2455 (O_2455,N_29894,N_29898);
xnor UO_2456 (O_2456,N_29953,N_29946);
nor UO_2457 (O_2457,N_29891,N_29805);
or UO_2458 (O_2458,N_29985,N_29927);
and UO_2459 (O_2459,N_29870,N_29986);
or UO_2460 (O_2460,N_29949,N_29953);
xor UO_2461 (O_2461,N_29810,N_29800);
nand UO_2462 (O_2462,N_29842,N_29823);
nor UO_2463 (O_2463,N_29962,N_29948);
nand UO_2464 (O_2464,N_29812,N_29925);
nor UO_2465 (O_2465,N_29850,N_29992);
or UO_2466 (O_2466,N_29978,N_29993);
xnor UO_2467 (O_2467,N_29879,N_29921);
and UO_2468 (O_2468,N_29812,N_29875);
or UO_2469 (O_2469,N_29893,N_29836);
or UO_2470 (O_2470,N_29819,N_29948);
and UO_2471 (O_2471,N_29974,N_29969);
nand UO_2472 (O_2472,N_29838,N_29822);
nand UO_2473 (O_2473,N_29917,N_29986);
nand UO_2474 (O_2474,N_29821,N_29857);
nand UO_2475 (O_2475,N_29852,N_29820);
and UO_2476 (O_2476,N_29937,N_29958);
and UO_2477 (O_2477,N_29978,N_29831);
nor UO_2478 (O_2478,N_29876,N_29837);
or UO_2479 (O_2479,N_29984,N_29843);
nand UO_2480 (O_2480,N_29803,N_29827);
xor UO_2481 (O_2481,N_29819,N_29922);
xor UO_2482 (O_2482,N_29985,N_29973);
or UO_2483 (O_2483,N_29947,N_29871);
nand UO_2484 (O_2484,N_29933,N_29905);
nor UO_2485 (O_2485,N_29959,N_29905);
and UO_2486 (O_2486,N_29918,N_29848);
or UO_2487 (O_2487,N_29966,N_29852);
and UO_2488 (O_2488,N_29913,N_29942);
nand UO_2489 (O_2489,N_29964,N_29921);
xnor UO_2490 (O_2490,N_29804,N_29923);
nor UO_2491 (O_2491,N_29947,N_29975);
nor UO_2492 (O_2492,N_29880,N_29987);
or UO_2493 (O_2493,N_29906,N_29965);
nand UO_2494 (O_2494,N_29926,N_29887);
nor UO_2495 (O_2495,N_29914,N_29921);
and UO_2496 (O_2496,N_29999,N_29842);
nand UO_2497 (O_2497,N_29997,N_29898);
xor UO_2498 (O_2498,N_29830,N_29962);
or UO_2499 (O_2499,N_29958,N_29967);
nor UO_2500 (O_2500,N_29932,N_29809);
nor UO_2501 (O_2501,N_29864,N_29888);
or UO_2502 (O_2502,N_29893,N_29962);
and UO_2503 (O_2503,N_29919,N_29813);
nand UO_2504 (O_2504,N_29830,N_29951);
xor UO_2505 (O_2505,N_29822,N_29990);
nor UO_2506 (O_2506,N_29848,N_29826);
nand UO_2507 (O_2507,N_29942,N_29820);
or UO_2508 (O_2508,N_29812,N_29918);
xnor UO_2509 (O_2509,N_29800,N_29894);
nor UO_2510 (O_2510,N_29993,N_29894);
or UO_2511 (O_2511,N_29807,N_29969);
nor UO_2512 (O_2512,N_29839,N_29817);
or UO_2513 (O_2513,N_29815,N_29939);
or UO_2514 (O_2514,N_29802,N_29881);
and UO_2515 (O_2515,N_29806,N_29927);
nand UO_2516 (O_2516,N_29993,N_29988);
nor UO_2517 (O_2517,N_29852,N_29967);
nor UO_2518 (O_2518,N_29921,N_29806);
nand UO_2519 (O_2519,N_29852,N_29909);
or UO_2520 (O_2520,N_29963,N_29821);
nand UO_2521 (O_2521,N_29890,N_29850);
and UO_2522 (O_2522,N_29903,N_29864);
nand UO_2523 (O_2523,N_29902,N_29859);
or UO_2524 (O_2524,N_29905,N_29874);
and UO_2525 (O_2525,N_29957,N_29950);
nand UO_2526 (O_2526,N_29985,N_29875);
nand UO_2527 (O_2527,N_29948,N_29907);
and UO_2528 (O_2528,N_29963,N_29958);
or UO_2529 (O_2529,N_29888,N_29853);
or UO_2530 (O_2530,N_29803,N_29912);
or UO_2531 (O_2531,N_29864,N_29800);
xnor UO_2532 (O_2532,N_29866,N_29862);
xnor UO_2533 (O_2533,N_29891,N_29857);
nor UO_2534 (O_2534,N_29901,N_29820);
xor UO_2535 (O_2535,N_29816,N_29806);
and UO_2536 (O_2536,N_29831,N_29839);
xnor UO_2537 (O_2537,N_29934,N_29908);
and UO_2538 (O_2538,N_29959,N_29918);
or UO_2539 (O_2539,N_29999,N_29885);
nor UO_2540 (O_2540,N_29990,N_29986);
nand UO_2541 (O_2541,N_29945,N_29853);
or UO_2542 (O_2542,N_29802,N_29862);
nand UO_2543 (O_2543,N_29858,N_29941);
xnor UO_2544 (O_2544,N_29881,N_29842);
or UO_2545 (O_2545,N_29985,N_29870);
nor UO_2546 (O_2546,N_29921,N_29887);
xnor UO_2547 (O_2547,N_29939,N_29821);
or UO_2548 (O_2548,N_29947,N_29813);
xor UO_2549 (O_2549,N_29859,N_29826);
and UO_2550 (O_2550,N_29846,N_29859);
and UO_2551 (O_2551,N_29994,N_29975);
nor UO_2552 (O_2552,N_29800,N_29847);
or UO_2553 (O_2553,N_29940,N_29863);
nor UO_2554 (O_2554,N_29822,N_29948);
nor UO_2555 (O_2555,N_29803,N_29856);
nand UO_2556 (O_2556,N_29865,N_29992);
nor UO_2557 (O_2557,N_29999,N_29963);
nor UO_2558 (O_2558,N_29808,N_29893);
xor UO_2559 (O_2559,N_29983,N_29895);
nor UO_2560 (O_2560,N_29876,N_29936);
and UO_2561 (O_2561,N_29884,N_29899);
nand UO_2562 (O_2562,N_29809,N_29847);
nand UO_2563 (O_2563,N_29822,N_29852);
nand UO_2564 (O_2564,N_29971,N_29983);
and UO_2565 (O_2565,N_29886,N_29873);
xnor UO_2566 (O_2566,N_29995,N_29951);
and UO_2567 (O_2567,N_29826,N_29921);
and UO_2568 (O_2568,N_29949,N_29812);
and UO_2569 (O_2569,N_29945,N_29949);
and UO_2570 (O_2570,N_29842,N_29937);
and UO_2571 (O_2571,N_29974,N_29982);
and UO_2572 (O_2572,N_29825,N_29936);
nand UO_2573 (O_2573,N_29860,N_29816);
or UO_2574 (O_2574,N_29955,N_29856);
nand UO_2575 (O_2575,N_29874,N_29811);
nand UO_2576 (O_2576,N_29976,N_29921);
xor UO_2577 (O_2577,N_29885,N_29816);
xor UO_2578 (O_2578,N_29850,N_29922);
nor UO_2579 (O_2579,N_29956,N_29830);
nand UO_2580 (O_2580,N_29935,N_29992);
or UO_2581 (O_2581,N_29889,N_29932);
or UO_2582 (O_2582,N_29841,N_29855);
xor UO_2583 (O_2583,N_29847,N_29828);
nand UO_2584 (O_2584,N_29899,N_29939);
nor UO_2585 (O_2585,N_29905,N_29837);
and UO_2586 (O_2586,N_29953,N_29964);
nor UO_2587 (O_2587,N_29888,N_29988);
or UO_2588 (O_2588,N_29877,N_29893);
nor UO_2589 (O_2589,N_29863,N_29888);
or UO_2590 (O_2590,N_29861,N_29852);
and UO_2591 (O_2591,N_29826,N_29918);
nor UO_2592 (O_2592,N_29950,N_29813);
and UO_2593 (O_2593,N_29895,N_29977);
xnor UO_2594 (O_2594,N_29925,N_29989);
or UO_2595 (O_2595,N_29820,N_29927);
or UO_2596 (O_2596,N_29906,N_29859);
xor UO_2597 (O_2597,N_29880,N_29892);
nor UO_2598 (O_2598,N_29892,N_29870);
nor UO_2599 (O_2599,N_29960,N_29957);
or UO_2600 (O_2600,N_29930,N_29890);
nand UO_2601 (O_2601,N_29860,N_29836);
and UO_2602 (O_2602,N_29872,N_29817);
nand UO_2603 (O_2603,N_29982,N_29890);
nand UO_2604 (O_2604,N_29985,N_29858);
and UO_2605 (O_2605,N_29879,N_29999);
nor UO_2606 (O_2606,N_29952,N_29905);
nor UO_2607 (O_2607,N_29874,N_29963);
nor UO_2608 (O_2608,N_29950,N_29817);
nand UO_2609 (O_2609,N_29960,N_29945);
xor UO_2610 (O_2610,N_29860,N_29985);
xor UO_2611 (O_2611,N_29953,N_29984);
xor UO_2612 (O_2612,N_29804,N_29818);
and UO_2613 (O_2613,N_29951,N_29891);
or UO_2614 (O_2614,N_29986,N_29932);
xnor UO_2615 (O_2615,N_29846,N_29822);
nand UO_2616 (O_2616,N_29981,N_29848);
and UO_2617 (O_2617,N_29850,N_29960);
and UO_2618 (O_2618,N_29831,N_29955);
and UO_2619 (O_2619,N_29978,N_29988);
xor UO_2620 (O_2620,N_29981,N_29994);
xnor UO_2621 (O_2621,N_29945,N_29915);
nand UO_2622 (O_2622,N_29952,N_29951);
xor UO_2623 (O_2623,N_29840,N_29806);
and UO_2624 (O_2624,N_29968,N_29933);
xor UO_2625 (O_2625,N_29817,N_29986);
nor UO_2626 (O_2626,N_29834,N_29896);
xor UO_2627 (O_2627,N_29971,N_29930);
and UO_2628 (O_2628,N_29865,N_29956);
nor UO_2629 (O_2629,N_29805,N_29846);
xnor UO_2630 (O_2630,N_29868,N_29995);
or UO_2631 (O_2631,N_29833,N_29876);
nand UO_2632 (O_2632,N_29940,N_29835);
nor UO_2633 (O_2633,N_29831,N_29863);
or UO_2634 (O_2634,N_29943,N_29810);
and UO_2635 (O_2635,N_29966,N_29914);
xor UO_2636 (O_2636,N_29877,N_29803);
or UO_2637 (O_2637,N_29879,N_29875);
nor UO_2638 (O_2638,N_29889,N_29810);
nor UO_2639 (O_2639,N_29884,N_29926);
nand UO_2640 (O_2640,N_29955,N_29934);
and UO_2641 (O_2641,N_29983,N_29839);
and UO_2642 (O_2642,N_29858,N_29959);
nor UO_2643 (O_2643,N_29926,N_29823);
and UO_2644 (O_2644,N_29844,N_29883);
xor UO_2645 (O_2645,N_29878,N_29972);
nand UO_2646 (O_2646,N_29815,N_29969);
or UO_2647 (O_2647,N_29918,N_29827);
xnor UO_2648 (O_2648,N_29977,N_29896);
xnor UO_2649 (O_2649,N_29863,N_29855);
nor UO_2650 (O_2650,N_29809,N_29846);
and UO_2651 (O_2651,N_29841,N_29915);
and UO_2652 (O_2652,N_29930,N_29946);
nand UO_2653 (O_2653,N_29804,N_29926);
nand UO_2654 (O_2654,N_29863,N_29998);
nand UO_2655 (O_2655,N_29842,N_29956);
and UO_2656 (O_2656,N_29910,N_29971);
nand UO_2657 (O_2657,N_29879,N_29989);
xor UO_2658 (O_2658,N_29957,N_29944);
nor UO_2659 (O_2659,N_29947,N_29990);
or UO_2660 (O_2660,N_29873,N_29891);
or UO_2661 (O_2661,N_29801,N_29967);
and UO_2662 (O_2662,N_29867,N_29822);
nor UO_2663 (O_2663,N_29814,N_29845);
or UO_2664 (O_2664,N_29989,N_29992);
nand UO_2665 (O_2665,N_29903,N_29803);
and UO_2666 (O_2666,N_29895,N_29989);
nor UO_2667 (O_2667,N_29942,N_29927);
and UO_2668 (O_2668,N_29852,N_29929);
nor UO_2669 (O_2669,N_29885,N_29804);
or UO_2670 (O_2670,N_29972,N_29991);
nor UO_2671 (O_2671,N_29951,N_29800);
nor UO_2672 (O_2672,N_29943,N_29815);
nand UO_2673 (O_2673,N_29923,N_29897);
nor UO_2674 (O_2674,N_29922,N_29982);
or UO_2675 (O_2675,N_29945,N_29817);
nand UO_2676 (O_2676,N_29943,N_29828);
and UO_2677 (O_2677,N_29995,N_29821);
xor UO_2678 (O_2678,N_29829,N_29818);
xor UO_2679 (O_2679,N_29807,N_29914);
and UO_2680 (O_2680,N_29975,N_29991);
nand UO_2681 (O_2681,N_29927,N_29947);
nand UO_2682 (O_2682,N_29945,N_29886);
or UO_2683 (O_2683,N_29818,N_29834);
nor UO_2684 (O_2684,N_29842,N_29980);
and UO_2685 (O_2685,N_29962,N_29854);
nor UO_2686 (O_2686,N_29921,N_29860);
or UO_2687 (O_2687,N_29880,N_29824);
nand UO_2688 (O_2688,N_29914,N_29902);
nor UO_2689 (O_2689,N_29923,N_29919);
and UO_2690 (O_2690,N_29873,N_29937);
and UO_2691 (O_2691,N_29858,N_29963);
or UO_2692 (O_2692,N_29880,N_29980);
xor UO_2693 (O_2693,N_29862,N_29948);
xor UO_2694 (O_2694,N_29945,N_29931);
nand UO_2695 (O_2695,N_29958,N_29898);
xor UO_2696 (O_2696,N_29944,N_29985);
and UO_2697 (O_2697,N_29914,N_29865);
or UO_2698 (O_2698,N_29879,N_29971);
nand UO_2699 (O_2699,N_29897,N_29986);
nand UO_2700 (O_2700,N_29829,N_29915);
and UO_2701 (O_2701,N_29878,N_29875);
xnor UO_2702 (O_2702,N_29977,N_29881);
and UO_2703 (O_2703,N_29856,N_29865);
and UO_2704 (O_2704,N_29933,N_29903);
xor UO_2705 (O_2705,N_29893,N_29830);
xor UO_2706 (O_2706,N_29830,N_29972);
or UO_2707 (O_2707,N_29854,N_29960);
xor UO_2708 (O_2708,N_29918,N_29903);
and UO_2709 (O_2709,N_29871,N_29923);
and UO_2710 (O_2710,N_29855,N_29911);
nand UO_2711 (O_2711,N_29934,N_29865);
xor UO_2712 (O_2712,N_29940,N_29993);
nor UO_2713 (O_2713,N_29930,N_29848);
or UO_2714 (O_2714,N_29802,N_29806);
xor UO_2715 (O_2715,N_29917,N_29836);
nand UO_2716 (O_2716,N_29961,N_29920);
nor UO_2717 (O_2717,N_29925,N_29994);
or UO_2718 (O_2718,N_29902,N_29977);
nand UO_2719 (O_2719,N_29812,N_29838);
nand UO_2720 (O_2720,N_29856,N_29961);
and UO_2721 (O_2721,N_29945,N_29926);
or UO_2722 (O_2722,N_29991,N_29921);
xnor UO_2723 (O_2723,N_29917,N_29855);
and UO_2724 (O_2724,N_29959,N_29984);
xnor UO_2725 (O_2725,N_29912,N_29956);
nand UO_2726 (O_2726,N_29995,N_29911);
and UO_2727 (O_2727,N_29927,N_29966);
nand UO_2728 (O_2728,N_29832,N_29963);
and UO_2729 (O_2729,N_29891,N_29802);
nand UO_2730 (O_2730,N_29843,N_29970);
nand UO_2731 (O_2731,N_29904,N_29912);
nor UO_2732 (O_2732,N_29971,N_29868);
nor UO_2733 (O_2733,N_29972,N_29832);
nor UO_2734 (O_2734,N_29923,N_29838);
nand UO_2735 (O_2735,N_29886,N_29931);
nor UO_2736 (O_2736,N_29940,N_29996);
or UO_2737 (O_2737,N_29905,N_29891);
or UO_2738 (O_2738,N_29824,N_29954);
or UO_2739 (O_2739,N_29991,N_29946);
and UO_2740 (O_2740,N_29825,N_29843);
xor UO_2741 (O_2741,N_29937,N_29874);
xor UO_2742 (O_2742,N_29833,N_29866);
xnor UO_2743 (O_2743,N_29858,N_29830);
and UO_2744 (O_2744,N_29827,N_29906);
or UO_2745 (O_2745,N_29988,N_29836);
xor UO_2746 (O_2746,N_29898,N_29979);
and UO_2747 (O_2747,N_29922,N_29846);
or UO_2748 (O_2748,N_29984,N_29842);
nand UO_2749 (O_2749,N_29852,N_29817);
and UO_2750 (O_2750,N_29871,N_29944);
xor UO_2751 (O_2751,N_29843,N_29809);
and UO_2752 (O_2752,N_29891,N_29999);
xnor UO_2753 (O_2753,N_29958,N_29913);
or UO_2754 (O_2754,N_29934,N_29970);
and UO_2755 (O_2755,N_29996,N_29988);
nand UO_2756 (O_2756,N_29938,N_29928);
nand UO_2757 (O_2757,N_29847,N_29877);
nor UO_2758 (O_2758,N_29992,N_29816);
nor UO_2759 (O_2759,N_29953,N_29958);
nor UO_2760 (O_2760,N_29827,N_29833);
nor UO_2761 (O_2761,N_29853,N_29831);
nand UO_2762 (O_2762,N_29982,N_29947);
xnor UO_2763 (O_2763,N_29854,N_29841);
and UO_2764 (O_2764,N_29836,N_29901);
and UO_2765 (O_2765,N_29928,N_29976);
and UO_2766 (O_2766,N_29829,N_29804);
nand UO_2767 (O_2767,N_29980,N_29990);
xnor UO_2768 (O_2768,N_29845,N_29956);
nand UO_2769 (O_2769,N_29872,N_29804);
or UO_2770 (O_2770,N_29825,N_29830);
nand UO_2771 (O_2771,N_29930,N_29950);
nor UO_2772 (O_2772,N_29916,N_29965);
and UO_2773 (O_2773,N_29955,N_29872);
nand UO_2774 (O_2774,N_29901,N_29841);
xnor UO_2775 (O_2775,N_29879,N_29948);
nand UO_2776 (O_2776,N_29925,N_29966);
or UO_2777 (O_2777,N_29813,N_29933);
nand UO_2778 (O_2778,N_29926,N_29922);
nand UO_2779 (O_2779,N_29965,N_29852);
or UO_2780 (O_2780,N_29871,N_29843);
xor UO_2781 (O_2781,N_29996,N_29970);
xnor UO_2782 (O_2782,N_29996,N_29855);
or UO_2783 (O_2783,N_29808,N_29829);
or UO_2784 (O_2784,N_29928,N_29948);
nand UO_2785 (O_2785,N_29993,N_29846);
and UO_2786 (O_2786,N_29861,N_29999);
xor UO_2787 (O_2787,N_29932,N_29915);
and UO_2788 (O_2788,N_29829,N_29852);
or UO_2789 (O_2789,N_29976,N_29960);
or UO_2790 (O_2790,N_29879,N_29906);
xor UO_2791 (O_2791,N_29814,N_29953);
and UO_2792 (O_2792,N_29857,N_29948);
nand UO_2793 (O_2793,N_29801,N_29862);
and UO_2794 (O_2794,N_29952,N_29877);
or UO_2795 (O_2795,N_29899,N_29829);
xnor UO_2796 (O_2796,N_29874,N_29911);
nor UO_2797 (O_2797,N_29856,N_29848);
and UO_2798 (O_2798,N_29938,N_29950);
or UO_2799 (O_2799,N_29892,N_29962);
nand UO_2800 (O_2800,N_29917,N_29909);
nor UO_2801 (O_2801,N_29867,N_29848);
and UO_2802 (O_2802,N_29830,N_29803);
xnor UO_2803 (O_2803,N_29996,N_29847);
nor UO_2804 (O_2804,N_29884,N_29879);
xor UO_2805 (O_2805,N_29895,N_29906);
or UO_2806 (O_2806,N_29872,N_29820);
nand UO_2807 (O_2807,N_29842,N_29935);
xnor UO_2808 (O_2808,N_29998,N_29825);
xnor UO_2809 (O_2809,N_29872,N_29917);
nand UO_2810 (O_2810,N_29955,N_29847);
xor UO_2811 (O_2811,N_29829,N_29841);
nor UO_2812 (O_2812,N_29845,N_29812);
xnor UO_2813 (O_2813,N_29957,N_29907);
or UO_2814 (O_2814,N_29900,N_29933);
and UO_2815 (O_2815,N_29903,N_29897);
nand UO_2816 (O_2816,N_29889,N_29914);
nand UO_2817 (O_2817,N_29982,N_29875);
nor UO_2818 (O_2818,N_29848,N_29822);
nand UO_2819 (O_2819,N_29844,N_29819);
and UO_2820 (O_2820,N_29864,N_29836);
or UO_2821 (O_2821,N_29865,N_29937);
or UO_2822 (O_2822,N_29804,N_29807);
or UO_2823 (O_2823,N_29977,N_29814);
nand UO_2824 (O_2824,N_29874,N_29978);
xor UO_2825 (O_2825,N_29949,N_29978);
nand UO_2826 (O_2826,N_29944,N_29834);
nor UO_2827 (O_2827,N_29939,N_29931);
nor UO_2828 (O_2828,N_29946,N_29938);
or UO_2829 (O_2829,N_29916,N_29837);
nor UO_2830 (O_2830,N_29909,N_29834);
nor UO_2831 (O_2831,N_29916,N_29852);
xnor UO_2832 (O_2832,N_29935,N_29802);
and UO_2833 (O_2833,N_29931,N_29907);
nor UO_2834 (O_2834,N_29900,N_29910);
nand UO_2835 (O_2835,N_29970,N_29850);
nor UO_2836 (O_2836,N_29982,N_29950);
or UO_2837 (O_2837,N_29838,N_29907);
nor UO_2838 (O_2838,N_29838,N_29950);
nand UO_2839 (O_2839,N_29851,N_29955);
nand UO_2840 (O_2840,N_29934,N_29806);
nor UO_2841 (O_2841,N_29967,N_29994);
nor UO_2842 (O_2842,N_29889,N_29895);
nor UO_2843 (O_2843,N_29861,N_29936);
or UO_2844 (O_2844,N_29992,N_29886);
or UO_2845 (O_2845,N_29943,N_29956);
or UO_2846 (O_2846,N_29881,N_29917);
xor UO_2847 (O_2847,N_29976,N_29901);
nor UO_2848 (O_2848,N_29960,N_29820);
and UO_2849 (O_2849,N_29891,N_29824);
or UO_2850 (O_2850,N_29891,N_29940);
nor UO_2851 (O_2851,N_29880,N_29998);
nand UO_2852 (O_2852,N_29955,N_29991);
or UO_2853 (O_2853,N_29949,N_29934);
nor UO_2854 (O_2854,N_29901,N_29995);
nand UO_2855 (O_2855,N_29855,N_29921);
and UO_2856 (O_2856,N_29956,N_29881);
xnor UO_2857 (O_2857,N_29883,N_29985);
nor UO_2858 (O_2858,N_29921,N_29932);
and UO_2859 (O_2859,N_29989,N_29844);
or UO_2860 (O_2860,N_29810,N_29969);
xor UO_2861 (O_2861,N_29941,N_29944);
xor UO_2862 (O_2862,N_29855,N_29990);
nand UO_2863 (O_2863,N_29842,N_29910);
xor UO_2864 (O_2864,N_29885,N_29832);
nand UO_2865 (O_2865,N_29945,N_29836);
xor UO_2866 (O_2866,N_29978,N_29895);
and UO_2867 (O_2867,N_29913,N_29977);
nand UO_2868 (O_2868,N_29990,N_29883);
or UO_2869 (O_2869,N_29872,N_29866);
or UO_2870 (O_2870,N_29867,N_29976);
xnor UO_2871 (O_2871,N_29934,N_29939);
nor UO_2872 (O_2872,N_29807,N_29890);
and UO_2873 (O_2873,N_29980,N_29835);
and UO_2874 (O_2874,N_29825,N_29981);
xor UO_2875 (O_2875,N_29874,N_29985);
or UO_2876 (O_2876,N_29882,N_29868);
and UO_2877 (O_2877,N_29968,N_29930);
nor UO_2878 (O_2878,N_29858,N_29843);
and UO_2879 (O_2879,N_29959,N_29967);
or UO_2880 (O_2880,N_29968,N_29982);
nor UO_2881 (O_2881,N_29922,N_29998);
nor UO_2882 (O_2882,N_29952,N_29942);
nand UO_2883 (O_2883,N_29904,N_29839);
nand UO_2884 (O_2884,N_29819,N_29973);
xnor UO_2885 (O_2885,N_29973,N_29873);
nor UO_2886 (O_2886,N_29818,N_29868);
or UO_2887 (O_2887,N_29846,N_29947);
nor UO_2888 (O_2888,N_29866,N_29871);
nand UO_2889 (O_2889,N_29810,N_29840);
nand UO_2890 (O_2890,N_29923,N_29848);
xnor UO_2891 (O_2891,N_29887,N_29958);
xor UO_2892 (O_2892,N_29853,N_29931);
or UO_2893 (O_2893,N_29809,N_29982);
nand UO_2894 (O_2894,N_29927,N_29862);
nor UO_2895 (O_2895,N_29906,N_29944);
nor UO_2896 (O_2896,N_29917,N_29960);
xnor UO_2897 (O_2897,N_29805,N_29848);
xor UO_2898 (O_2898,N_29964,N_29922);
nand UO_2899 (O_2899,N_29834,N_29947);
and UO_2900 (O_2900,N_29949,N_29957);
xor UO_2901 (O_2901,N_29958,N_29964);
or UO_2902 (O_2902,N_29848,N_29885);
or UO_2903 (O_2903,N_29873,N_29920);
or UO_2904 (O_2904,N_29848,N_29862);
or UO_2905 (O_2905,N_29891,N_29814);
and UO_2906 (O_2906,N_29974,N_29894);
and UO_2907 (O_2907,N_29911,N_29964);
nor UO_2908 (O_2908,N_29854,N_29973);
nor UO_2909 (O_2909,N_29846,N_29876);
and UO_2910 (O_2910,N_29935,N_29993);
and UO_2911 (O_2911,N_29868,N_29946);
nor UO_2912 (O_2912,N_29936,N_29940);
nor UO_2913 (O_2913,N_29894,N_29866);
xnor UO_2914 (O_2914,N_29805,N_29994);
xnor UO_2915 (O_2915,N_29985,N_29826);
xnor UO_2916 (O_2916,N_29862,N_29881);
and UO_2917 (O_2917,N_29985,N_29872);
nor UO_2918 (O_2918,N_29828,N_29982);
xor UO_2919 (O_2919,N_29851,N_29878);
xor UO_2920 (O_2920,N_29880,N_29959);
xor UO_2921 (O_2921,N_29830,N_29948);
xnor UO_2922 (O_2922,N_29861,N_29990);
and UO_2923 (O_2923,N_29826,N_29836);
and UO_2924 (O_2924,N_29957,N_29835);
and UO_2925 (O_2925,N_29897,N_29825);
xor UO_2926 (O_2926,N_29940,N_29991);
and UO_2927 (O_2927,N_29948,N_29947);
and UO_2928 (O_2928,N_29804,N_29898);
and UO_2929 (O_2929,N_29978,N_29992);
xnor UO_2930 (O_2930,N_29864,N_29861);
and UO_2931 (O_2931,N_29944,N_29924);
and UO_2932 (O_2932,N_29965,N_29930);
xor UO_2933 (O_2933,N_29995,N_29858);
and UO_2934 (O_2934,N_29887,N_29954);
nand UO_2935 (O_2935,N_29835,N_29987);
nand UO_2936 (O_2936,N_29816,N_29809);
nor UO_2937 (O_2937,N_29837,N_29806);
nor UO_2938 (O_2938,N_29857,N_29880);
nor UO_2939 (O_2939,N_29940,N_29970);
nand UO_2940 (O_2940,N_29900,N_29917);
xnor UO_2941 (O_2941,N_29894,N_29843);
nor UO_2942 (O_2942,N_29862,N_29939);
nor UO_2943 (O_2943,N_29841,N_29939);
or UO_2944 (O_2944,N_29973,N_29932);
nor UO_2945 (O_2945,N_29845,N_29834);
xnor UO_2946 (O_2946,N_29847,N_29995);
nor UO_2947 (O_2947,N_29977,N_29804);
and UO_2948 (O_2948,N_29941,N_29878);
xor UO_2949 (O_2949,N_29894,N_29838);
nand UO_2950 (O_2950,N_29882,N_29809);
nor UO_2951 (O_2951,N_29840,N_29919);
and UO_2952 (O_2952,N_29885,N_29826);
xor UO_2953 (O_2953,N_29874,N_29987);
nand UO_2954 (O_2954,N_29843,N_29962);
nor UO_2955 (O_2955,N_29947,N_29807);
nor UO_2956 (O_2956,N_29828,N_29842);
nand UO_2957 (O_2957,N_29922,N_29859);
xor UO_2958 (O_2958,N_29994,N_29833);
or UO_2959 (O_2959,N_29853,N_29826);
nand UO_2960 (O_2960,N_29825,N_29960);
nand UO_2961 (O_2961,N_29802,N_29870);
nor UO_2962 (O_2962,N_29856,N_29879);
nand UO_2963 (O_2963,N_29906,N_29914);
nor UO_2964 (O_2964,N_29858,N_29898);
or UO_2965 (O_2965,N_29922,N_29812);
or UO_2966 (O_2966,N_29982,N_29853);
xnor UO_2967 (O_2967,N_29856,N_29860);
nand UO_2968 (O_2968,N_29808,N_29990);
nand UO_2969 (O_2969,N_29955,N_29978);
xor UO_2970 (O_2970,N_29801,N_29928);
nand UO_2971 (O_2971,N_29884,N_29943);
and UO_2972 (O_2972,N_29951,N_29893);
or UO_2973 (O_2973,N_29942,N_29869);
and UO_2974 (O_2974,N_29845,N_29964);
or UO_2975 (O_2975,N_29973,N_29959);
or UO_2976 (O_2976,N_29975,N_29912);
nand UO_2977 (O_2977,N_29979,N_29969);
nand UO_2978 (O_2978,N_29903,N_29981);
nand UO_2979 (O_2979,N_29860,N_29966);
and UO_2980 (O_2980,N_29835,N_29907);
and UO_2981 (O_2981,N_29957,N_29884);
and UO_2982 (O_2982,N_29823,N_29832);
xnor UO_2983 (O_2983,N_29939,N_29925);
nor UO_2984 (O_2984,N_29844,N_29843);
xnor UO_2985 (O_2985,N_29870,N_29992);
xnor UO_2986 (O_2986,N_29885,N_29898);
nor UO_2987 (O_2987,N_29878,N_29902);
or UO_2988 (O_2988,N_29970,N_29919);
and UO_2989 (O_2989,N_29841,N_29867);
nor UO_2990 (O_2990,N_29964,N_29900);
xor UO_2991 (O_2991,N_29861,N_29840);
and UO_2992 (O_2992,N_29812,N_29902);
nand UO_2993 (O_2993,N_29817,N_29829);
or UO_2994 (O_2994,N_29873,N_29941);
nor UO_2995 (O_2995,N_29927,N_29883);
nor UO_2996 (O_2996,N_29951,N_29896);
xor UO_2997 (O_2997,N_29951,N_29886);
nand UO_2998 (O_2998,N_29850,N_29832);
nand UO_2999 (O_2999,N_29810,N_29819);
nand UO_3000 (O_3000,N_29837,N_29819);
or UO_3001 (O_3001,N_29994,N_29993);
and UO_3002 (O_3002,N_29923,N_29949);
nor UO_3003 (O_3003,N_29913,N_29967);
nand UO_3004 (O_3004,N_29928,N_29998);
nand UO_3005 (O_3005,N_29953,N_29817);
nor UO_3006 (O_3006,N_29863,N_29864);
nor UO_3007 (O_3007,N_29822,N_29896);
nor UO_3008 (O_3008,N_29934,N_29807);
nand UO_3009 (O_3009,N_29881,N_29926);
nor UO_3010 (O_3010,N_29935,N_29902);
nand UO_3011 (O_3011,N_29813,N_29902);
nand UO_3012 (O_3012,N_29910,N_29916);
nor UO_3013 (O_3013,N_29978,N_29983);
xnor UO_3014 (O_3014,N_29984,N_29971);
nor UO_3015 (O_3015,N_29931,N_29979);
and UO_3016 (O_3016,N_29960,N_29803);
and UO_3017 (O_3017,N_29988,N_29921);
and UO_3018 (O_3018,N_29838,N_29833);
nand UO_3019 (O_3019,N_29821,N_29929);
nor UO_3020 (O_3020,N_29861,N_29982);
and UO_3021 (O_3021,N_29907,N_29900);
nor UO_3022 (O_3022,N_29811,N_29973);
or UO_3023 (O_3023,N_29911,N_29847);
or UO_3024 (O_3024,N_29968,N_29970);
nand UO_3025 (O_3025,N_29825,N_29842);
nand UO_3026 (O_3026,N_29800,N_29872);
nand UO_3027 (O_3027,N_29906,N_29989);
and UO_3028 (O_3028,N_29924,N_29936);
nand UO_3029 (O_3029,N_29930,N_29940);
nor UO_3030 (O_3030,N_29809,N_29837);
or UO_3031 (O_3031,N_29942,N_29932);
or UO_3032 (O_3032,N_29894,N_29970);
nand UO_3033 (O_3033,N_29877,N_29931);
nor UO_3034 (O_3034,N_29847,N_29904);
nor UO_3035 (O_3035,N_29897,N_29976);
xor UO_3036 (O_3036,N_29819,N_29935);
nor UO_3037 (O_3037,N_29810,N_29863);
or UO_3038 (O_3038,N_29830,N_29923);
nor UO_3039 (O_3039,N_29832,N_29839);
nor UO_3040 (O_3040,N_29911,N_29851);
and UO_3041 (O_3041,N_29978,N_29862);
nor UO_3042 (O_3042,N_29930,N_29933);
and UO_3043 (O_3043,N_29960,N_29994);
nand UO_3044 (O_3044,N_29812,N_29888);
nor UO_3045 (O_3045,N_29829,N_29917);
xor UO_3046 (O_3046,N_29976,N_29981);
xnor UO_3047 (O_3047,N_29983,N_29923);
or UO_3048 (O_3048,N_29978,N_29817);
nor UO_3049 (O_3049,N_29993,N_29961);
nand UO_3050 (O_3050,N_29914,N_29908);
nand UO_3051 (O_3051,N_29955,N_29913);
nor UO_3052 (O_3052,N_29939,N_29810);
and UO_3053 (O_3053,N_29932,N_29888);
or UO_3054 (O_3054,N_29911,N_29934);
or UO_3055 (O_3055,N_29835,N_29858);
nand UO_3056 (O_3056,N_29953,N_29830);
and UO_3057 (O_3057,N_29933,N_29965);
nand UO_3058 (O_3058,N_29829,N_29827);
or UO_3059 (O_3059,N_29814,N_29944);
or UO_3060 (O_3060,N_29970,N_29802);
nor UO_3061 (O_3061,N_29888,N_29976);
xnor UO_3062 (O_3062,N_29890,N_29952);
nand UO_3063 (O_3063,N_29947,N_29916);
xnor UO_3064 (O_3064,N_29850,N_29814);
or UO_3065 (O_3065,N_29872,N_29870);
xnor UO_3066 (O_3066,N_29884,N_29835);
and UO_3067 (O_3067,N_29815,N_29973);
and UO_3068 (O_3068,N_29823,N_29928);
xor UO_3069 (O_3069,N_29897,N_29812);
or UO_3070 (O_3070,N_29821,N_29828);
nand UO_3071 (O_3071,N_29952,N_29819);
nor UO_3072 (O_3072,N_29961,N_29995);
nor UO_3073 (O_3073,N_29976,N_29858);
nand UO_3074 (O_3074,N_29999,N_29839);
nor UO_3075 (O_3075,N_29947,N_29987);
or UO_3076 (O_3076,N_29879,N_29848);
and UO_3077 (O_3077,N_29954,N_29892);
nand UO_3078 (O_3078,N_29812,N_29827);
and UO_3079 (O_3079,N_29945,N_29842);
nor UO_3080 (O_3080,N_29837,N_29901);
or UO_3081 (O_3081,N_29809,N_29984);
nand UO_3082 (O_3082,N_29847,N_29830);
nand UO_3083 (O_3083,N_29970,N_29853);
and UO_3084 (O_3084,N_29902,N_29934);
nand UO_3085 (O_3085,N_29995,N_29965);
nand UO_3086 (O_3086,N_29967,N_29948);
or UO_3087 (O_3087,N_29878,N_29937);
and UO_3088 (O_3088,N_29887,N_29815);
nor UO_3089 (O_3089,N_29841,N_29905);
xor UO_3090 (O_3090,N_29861,N_29888);
xor UO_3091 (O_3091,N_29926,N_29816);
nor UO_3092 (O_3092,N_29815,N_29910);
xor UO_3093 (O_3093,N_29997,N_29937);
xor UO_3094 (O_3094,N_29921,N_29984);
and UO_3095 (O_3095,N_29831,N_29827);
nor UO_3096 (O_3096,N_29869,N_29885);
nor UO_3097 (O_3097,N_29898,N_29991);
nor UO_3098 (O_3098,N_29824,N_29818);
or UO_3099 (O_3099,N_29979,N_29992);
and UO_3100 (O_3100,N_29949,N_29846);
xor UO_3101 (O_3101,N_29908,N_29822);
nand UO_3102 (O_3102,N_29936,N_29947);
and UO_3103 (O_3103,N_29936,N_29979);
and UO_3104 (O_3104,N_29935,N_29858);
xor UO_3105 (O_3105,N_29982,N_29852);
or UO_3106 (O_3106,N_29857,N_29937);
nand UO_3107 (O_3107,N_29842,N_29811);
xor UO_3108 (O_3108,N_29917,N_29879);
nor UO_3109 (O_3109,N_29839,N_29958);
and UO_3110 (O_3110,N_29874,N_29847);
xor UO_3111 (O_3111,N_29880,N_29958);
nor UO_3112 (O_3112,N_29820,N_29873);
nor UO_3113 (O_3113,N_29979,N_29952);
and UO_3114 (O_3114,N_29804,N_29878);
xor UO_3115 (O_3115,N_29987,N_29818);
nor UO_3116 (O_3116,N_29994,N_29908);
and UO_3117 (O_3117,N_29997,N_29949);
and UO_3118 (O_3118,N_29941,N_29929);
nand UO_3119 (O_3119,N_29933,N_29961);
nor UO_3120 (O_3120,N_29867,N_29972);
or UO_3121 (O_3121,N_29940,N_29984);
or UO_3122 (O_3122,N_29880,N_29807);
and UO_3123 (O_3123,N_29873,N_29909);
and UO_3124 (O_3124,N_29996,N_29907);
or UO_3125 (O_3125,N_29806,N_29900);
and UO_3126 (O_3126,N_29809,N_29823);
nor UO_3127 (O_3127,N_29878,N_29917);
nand UO_3128 (O_3128,N_29847,N_29806);
and UO_3129 (O_3129,N_29866,N_29895);
or UO_3130 (O_3130,N_29885,N_29864);
nor UO_3131 (O_3131,N_29821,N_29880);
xnor UO_3132 (O_3132,N_29973,N_29988);
and UO_3133 (O_3133,N_29984,N_29920);
nor UO_3134 (O_3134,N_29861,N_29919);
or UO_3135 (O_3135,N_29974,N_29996);
nand UO_3136 (O_3136,N_29889,N_29987);
and UO_3137 (O_3137,N_29881,N_29953);
nor UO_3138 (O_3138,N_29936,N_29923);
nand UO_3139 (O_3139,N_29843,N_29914);
xor UO_3140 (O_3140,N_29836,N_29884);
nor UO_3141 (O_3141,N_29851,N_29843);
nor UO_3142 (O_3142,N_29830,N_29809);
nor UO_3143 (O_3143,N_29921,N_29849);
xnor UO_3144 (O_3144,N_29915,N_29834);
or UO_3145 (O_3145,N_29844,N_29865);
xor UO_3146 (O_3146,N_29881,N_29807);
and UO_3147 (O_3147,N_29990,N_29970);
or UO_3148 (O_3148,N_29894,N_29819);
or UO_3149 (O_3149,N_29849,N_29982);
nand UO_3150 (O_3150,N_29832,N_29957);
nand UO_3151 (O_3151,N_29815,N_29880);
and UO_3152 (O_3152,N_29863,N_29937);
or UO_3153 (O_3153,N_29854,N_29892);
or UO_3154 (O_3154,N_29826,N_29810);
and UO_3155 (O_3155,N_29994,N_29939);
and UO_3156 (O_3156,N_29867,N_29843);
nand UO_3157 (O_3157,N_29809,N_29922);
or UO_3158 (O_3158,N_29937,N_29854);
and UO_3159 (O_3159,N_29895,N_29826);
and UO_3160 (O_3160,N_29927,N_29938);
or UO_3161 (O_3161,N_29822,N_29857);
or UO_3162 (O_3162,N_29900,N_29920);
and UO_3163 (O_3163,N_29826,N_29909);
or UO_3164 (O_3164,N_29898,N_29808);
xnor UO_3165 (O_3165,N_29908,N_29971);
and UO_3166 (O_3166,N_29917,N_29804);
nand UO_3167 (O_3167,N_29805,N_29951);
xnor UO_3168 (O_3168,N_29865,N_29882);
nand UO_3169 (O_3169,N_29985,N_29978);
nor UO_3170 (O_3170,N_29967,N_29941);
xnor UO_3171 (O_3171,N_29818,N_29915);
nor UO_3172 (O_3172,N_29848,N_29883);
nand UO_3173 (O_3173,N_29848,N_29939);
or UO_3174 (O_3174,N_29894,N_29806);
or UO_3175 (O_3175,N_29909,N_29967);
or UO_3176 (O_3176,N_29904,N_29988);
xor UO_3177 (O_3177,N_29872,N_29878);
nor UO_3178 (O_3178,N_29850,N_29940);
nand UO_3179 (O_3179,N_29887,N_29806);
nor UO_3180 (O_3180,N_29938,N_29892);
nor UO_3181 (O_3181,N_29818,N_29863);
nor UO_3182 (O_3182,N_29878,N_29865);
xnor UO_3183 (O_3183,N_29905,N_29862);
nand UO_3184 (O_3184,N_29904,N_29996);
nand UO_3185 (O_3185,N_29982,N_29937);
nand UO_3186 (O_3186,N_29993,N_29851);
nand UO_3187 (O_3187,N_29999,N_29912);
nand UO_3188 (O_3188,N_29818,N_29822);
or UO_3189 (O_3189,N_29801,N_29929);
or UO_3190 (O_3190,N_29983,N_29887);
xnor UO_3191 (O_3191,N_29821,N_29966);
nor UO_3192 (O_3192,N_29930,N_29925);
xor UO_3193 (O_3193,N_29979,N_29971);
or UO_3194 (O_3194,N_29866,N_29926);
and UO_3195 (O_3195,N_29987,N_29851);
and UO_3196 (O_3196,N_29949,N_29977);
or UO_3197 (O_3197,N_29942,N_29824);
xnor UO_3198 (O_3198,N_29848,N_29992);
and UO_3199 (O_3199,N_29878,N_29881);
nor UO_3200 (O_3200,N_29955,N_29997);
and UO_3201 (O_3201,N_29806,N_29813);
nor UO_3202 (O_3202,N_29895,N_29881);
and UO_3203 (O_3203,N_29899,N_29859);
xor UO_3204 (O_3204,N_29882,N_29973);
and UO_3205 (O_3205,N_29821,N_29973);
or UO_3206 (O_3206,N_29802,N_29949);
xnor UO_3207 (O_3207,N_29866,N_29911);
xnor UO_3208 (O_3208,N_29819,N_29915);
and UO_3209 (O_3209,N_29895,N_29934);
xor UO_3210 (O_3210,N_29960,N_29885);
or UO_3211 (O_3211,N_29884,N_29940);
or UO_3212 (O_3212,N_29888,N_29833);
nor UO_3213 (O_3213,N_29899,N_29842);
xnor UO_3214 (O_3214,N_29855,N_29972);
xor UO_3215 (O_3215,N_29804,N_29938);
or UO_3216 (O_3216,N_29964,N_29898);
nand UO_3217 (O_3217,N_29816,N_29801);
xor UO_3218 (O_3218,N_29976,N_29959);
nand UO_3219 (O_3219,N_29881,N_29982);
or UO_3220 (O_3220,N_29973,N_29944);
nand UO_3221 (O_3221,N_29840,N_29991);
nand UO_3222 (O_3222,N_29968,N_29891);
xor UO_3223 (O_3223,N_29897,N_29836);
nor UO_3224 (O_3224,N_29934,N_29809);
nor UO_3225 (O_3225,N_29912,N_29860);
and UO_3226 (O_3226,N_29860,N_29974);
nor UO_3227 (O_3227,N_29899,N_29860);
nor UO_3228 (O_3228,N_29955,N_29815);
and UO_3229 (O_3229,N_29890,N_29946);
xnor UO_3230 (O_3230,N_29864,N_29921);
nand UO_3231 (O_3231,N_29899,N_29818);
xnor UO_3232 (O_3232,N_29989,N_29926);
and UO_3233 (O_3233,N_29919,N_29872);
nand UO_3234 (O_3234,N_29844,N_29905);
xnor UO_3235 (O_3235,N_29825,N_29804);
nor UO_3236 (O_3236,N_29967,N_29939);
and UO_3237 (O_3237,N_29851,N_29884);
nor UO_3238 (O_3238,N_29870,N_29958);
nor UO_3239 (O_3239,N_29833,N_29892);
nand UO_3240 (O_3240,N_29832,N_29847);
nor UO_3241 (O_3241,N_29954,N_29964);
nor UO_3242 (O_3242,N_29853,N_29861);
nor UO_3243 (O_3243,N_29848,N_29947);
nand UO_3244 (O_3244,N_29975,N_29887);
xor UO_3245 (O_3245,N_29946,N_29803);
nand UO_3246 (O_3246,N_29901,N_29860);
nor UO_3247 (O_3247,N_29867,N_29920);
xnor UO_3248 (O_3248,N_29860,N_29979);
or UO_3249 (O_3249,N_29891,N_29847);
xnor UO_3250 (O_3250,N_29842,N_29905);
xnor UO_3251 (O_3251,N_29881,N_29955);
nand UO_3252 (O_3252,N_29864,N_29866);
nor UO_3253 (O_3253,N_29896,N_29956);
or UO_3254 (O_3254,N_29846,N_29823);
nor UO_3255 (O_3255,N_29895,N_29933);
or UO_3256 (O_3256,N_29909,N_29983);
nand UO_3257 (O_3257,N_29848,N_29874);
xnor UO_3258 (O_3258,N_29872,N_29858);
or UO_3259 (O_3259,N_29891,N_29822);
nor UO_3260 (O_3260,N_29875,N_29870);
xor UO_3261 (O_3261,N_29921,N_29815);
nor UO_3262 (O_3262,N_29887,N_29993);
nor UO_3263 (O_3263,N_29822,N_29839);
and UO_3264 (O_3264,N_29929,N_29922);
xor UO_3265 (O_3265,N_29871,N_29962);
nand UO_3266 (O_3266,N_29996,N_29831);
nor UO_3267 (O_3267,N_29831,N_29958);
and UO_3268 (O_3268,N_29817,N_29903);
nor UO_3269 (O_3269,N_29832,N_29932);
nand UO_3270 (O_3270,N_29944,N_29800);
nand UO_3271 (O_3271,N_29844,N_29978);
xor UO_3272 (O_3272,N_29899,N_29902);
nand UO_3273 (O_3273,N_29804,N_29842);
and UO_3274 (O_3274,N_29920,N_29860);
or UO_3275 (O_3275,N_29813,N_29884);
nand UO_3276 (O_3276,N_29867,N_29831);
and UO_3277 (O_3277,N_29982,N_29926);
or UO_3278 (O_3278,N_29912,N_29946);
or UO_3279 (O_3279,N_29986,N_29979);
nor UO_3280 (O_3280,N_29808,N_29950);
nand UO_3281 (O_3281,N_29881,N_29938);
xnor UO_3282 (O_3282,N_29956,N_29937);
nor UO_3283 (O_3283,N_29934,N_29826);
and UO_3284 (O_3284,N_29817,N_29808);
or UO_3285 (O_3285,N_29996,N_29865);
nor UO_3286 (O_3286,N_29998,N_29942);
nand UO_3287 (O_3287,N_29828,N_29883);
xor UO_3288 (O_3288,N_29819,N_29845);
and UO_3289 (O_3289,N_29829,N_29859);
nor UO_3290 (O_3290,N_29870,N_29829);
and UO_3291 (O_3291,N_29893,N_29940);
nor UO_3292 (O_3292,N_29912,N_29855);
nand UO_3293 (O_3293,N_29835,N_29890);
nand UO_3294 (O_3294,N_29870,N_29952);
or UO_3295 (O_3295,N_29810,N_29813);
nor UO_3296 (O_3296,N_29866,N_29831);
nand UO_3297 (O_3297,N_29881,N_29850);
xor UO_3298 (O_3298,N_29877,N_29845);
xor UO_3299 (O_3299,N_29946,N_29813);
xor UO_3300 (O_3300,N_29898,N_29878);
nor UO_3301 (O_3301,N_29915,N_29971);
and UO_3302 (O_3302,N_29990,N_29831);
and UO_3303 (O_3303,N_29897,N_29928);
and UO_3304 (O_3304,N_29988,N_29807);
or UO_3305 (O_3305,N_29832,N_29940);
nor UO_3306 (O_3306,N_29956,N_29990);
or UO_3307 (O_3307,N_29847,N_29963);
nor UO_3308 (O_3308,N_29883,N_29851);
xor UO_3309 (O_3309,N_29982,N_29962);
and UO_3310 (O_3310,N_29911,N_29918);
and UO_3311 (O_3311,N_29845,N_29809);
and UO_3312 (O_3312,N_29910,N_29932);
and UO_3313 (O_3313,N_29922,N_29825);
or UO_3314 (O_3314,N_29860,N_29840);
nor UO_3315 (O_3315,N_29852,N_29849);
nand UO_3316 (O_3316,N_29859,N_29948);
nand UO_3317 (O_3317,N_29915,N_29917);
nor UO_3318 (O_3318,N_29937,N_29849);
or UO_3319 (O_3319,N_29984,N_29866);
xor UO_3320 (O_3320,N_29901,N_29958);
and UO_3321 (O_3321,N_29986,N_29865);
or UO_3322 (O_3322,N_29925,N_29884);
or UO_3323 (O_3323,N_29920,N_29974);
and UO_3324 (O_3324,N_29830,N_29960);
or UO_3325 (O_3325,N_29917,N_29971);
and UO_3326 (O_3326,N_29979,N_29940);
nor UO_3327 (O_3327,N_29883,N_29838);
and UO_3328 (O_3328,N_29884,N_29945);
nand UO_3329 (O_3329,N_29825,N_29892);
xnor UO_3330 (O_3330,N_29817,N_29833);
nand UO_3331 (O_3331,N_29802,N_29828);
and UO_3332 (O_3332,N_29880,N_29940);
nor UO_3333 (O_3333,N_29951,N_29813);
nor UO_3334 (O_3334,N_29817,N_29853);
xor UO_3335 (O_3335,N_29851,N_29894);
and UO_3336 (O_3336,N_29834,N_29997);
or UO_3337 (O_3337,N_29837,N_29950);
or UO_3338 (O_3338,N_29803,N_29971);
and UO_3339 (O_3339,N_29903,N_29839);
and UO_3340 (O_3340,N_29818,N_29901);
and UO_3341 (O_3341,N_29975,N_29907);
and UO_3342 (O_3342,N_29889,N_29940);
or UO_3343 (O_3343,N_29877,N_29971);
nand UO_3344 (O_3344,N_29946,N_29875);
xor UO_3345 (O_3345,N_29991,N_29874);
nor UO_3346 (O_3346,N_29959,N_29957);
nor UO_3347 (O_3347,N_29893,N_29863);
and UO_3348 (O_3348,N_29831,N_29855);
xor UO_3349 (O_3349,N_29910,N_29929);
and UO_3350 (O_3350,N_29882,N_29941);
xnor UO_3351 (O_3351,N_29880,N_29825);
and UO_3352 (O_3352,N_29821,N_29861);
and UO_3353 (O_3353,N_29876,N_29815);
or UO_3354 (O_3354,N_29886,N_29854);
nand UO_3355 (O_3355,N_29927,N_29856);
and UO_3356 (O_3356,N_29977,N_29968);
nor UO_3357 (O_3357,N_29910,N_29845);
nor UO_3358 (O_3358,N_29975,N_29866);
nor UO_3359 (O_3359,N_29978,N_29959);
or UO_3360 (O_3360,N_29854,N_29945);
nand UO_3361 (O_3361,N_29807,N_29808);
and UO_3362 (O_3362,N_29839,N_29812);
and UO_3363 (O_3363,N_29870,N_29991);
xnor UO_3364 (O_3364,N_29853,N_29898);
xnor UO_3365 (O_3365,N_29998,N_29924);
nor UO_3366 (O_3366,N_29891,N_29901);
and UO_3367 (O_3367,N_29827,N_29948);
and UO_3368 (O_3368,N_29972,N_29848);
nand UO_3369 (O_3369,N_29927,N_29923);
nand UO_3370 (O_3370,N_29805,N_29831);
or UO_3371 (O_3371,N_29980,N_29929);
or UO_3372 (O_3372,N_29841,N_29998);
nor UO_3373 (O_3373,N_29898,N_29970);
nand UO_3374 (O_3374,N_29831,N_29876);
nor UO_3375 (O_3375,N_29891,N_29948);
nor UO_3376 (O_3376,N_29968,N_29809);
and UO_3377 (O_3377,N_29868,N_29993);
xor UO_3378 (O_3378,N_29924,N_29881);
nand UO_3379 (O_3379,N_29945,N_29863);
xor UO_3380 (O_3380,N_29920,N_29906);
xor UO_3381 (O_3381,N_29958,N_29966);
nand UO_3382 (O_3382,N_29887,N_29838);
xnor UO_3383 (O_3383,N_29977,N_29828);
xor UO_3384 (O_3384,N_29940,N_29987);
nor UO_3385 (O_3385,N_29971,N_29800);
or UO_3386 (O_3386,N_29886,N_29850);
xnor UO_3387 (O_3387,N_29816,N_29859);
xnor UO_3388 (O_3388,N_29864,N_29914);
xor UO_3389 (O_3389,N_29830,N_29874);
xnor UO_3390 (O_3390,N_29837,N_29882);
nor UO_3391 (O_3391,N_29884,N_29822);
or UO_3392 (O_3392,N_29891,N_29884);
nor UO_3393 (O_3393,N_29988,N_29848);
and UO_3394 (O_3394,N_29864,N_29893);
xor UO_3395 (O_3395,N_29933,N_29910);
xnor UO_3396 (O_3396,N_29828,N_29894);
nor UO_3397 (O_3397,N_29981,N_29872);
nor UO_3398 (O_3398,N_29887,N_29968);
and UO_3399 (O_3399,N_29835,N_29821);
and UO_3400 (O_3400,N_29831,N_29952);
nand UO_3401 (O_3401,N_29939,N_29926);
nor UO_3402 (O_3402,N_29966,N_29891);
nor UO_3403 (O_3403,N_29908,N_29976);
nor UO_3404 (O_3404,N_29838,N_29936);
nor UO_3405 (O_3405,N_29920,N_29857);
xnor UO_3406 (O_3406,N_29889,N_29859);
xor UO_3407 (O_3407,N_29908,N_29830);
or UO_3408 (O_3408,N_29923,N_29921);
nor UO_3409 (O_3409,N_29906,N_29815);
nor UO_3410 (O_3410,N_29802,N_29811);
nor UO_3411 (O_3411,N_29969,N_29889);
xnor UO_3412 (O_3412,N_29839,N_29961);
or UO_3413 (O_3413,N_29863,N_29814);
nor UO_3414 (O_3414,N_29809,N_29895);
nor UO_3415 (O_3415,N_29867,N_29860);
or UO_3416 (O_3416,N_29817,N_29895);
or UO_3417 (O_3417,N_29982,N_29961);
nor UO_3418 (O_3418,N_29879,N_29998);
xnor UO_3419 (O_3419,N_29815,N_29873);
and UO_3420 (O_3420,N_29945,N_29857);
nor UO_3421 (O_3421,N_29901,N_29870);
and UO_3422 (O_3422,N_29802,N_29968);
nand UO_3423 (O_3423,N_29842,N_29916);
nand UO_3424 (O_3424,N_29874,N_29838);
nand UO_3425 (O_3425,N_29999,N_29930);
or UO_3426 (O_3426,N_29944,N_29931);
or UO_3427 (O_3427,N_29885,N_29984);
and UO_3428 (O_3428,N_29991,N_29934);
xor UO_3429 (O_3429,N_29804,N_29817);
nand UO_3430 (O_3430,N_29955,N_29998);
xnor UO_3431 (O_3431,N_29894,N_29880);
xor UO_3432 (O_3432,N_29895,N_29911);
and UO_3433 (O_3433,N_29876,N_29935);
and UO_3434 (O_3434,N_29901,N_29889);
xnor UO_3435 (O_3435,N_29901,N_29879);
nand UO_3436 (O_3436,N_29856,N_29995);
or UO_3437 (O_3437,N_29963,N_29881);
nand UO_3438 (O_3438,N_29907,N_29805);
or UO_3439 (O_3439,N_29868,N_29942);
xnor UO_3440 (O_3440,N_29896,N_29854);
nor UO_3441 (O_3441,N_29958,N_29939);
xor UO_3442 (O_3442,N_29975,N_29811);
or UO_3443 (O_3443,N_29804,N_29996);
nor UO_3444 (O_3444,N_29928,N_29840);
or UO_3445 (O_3445,N_29918,N_29811);
and UO_3446 (O_3446,N_29849,N_29817);
xnor UO_3447 (O_3447,N_29911,N_29963);
xor UO_3448 (O_3448,N_29996,N_29975);
nand UO_3449 (O_3449,N_29844,N_29849);
or UO_3450 (O_3450,N_29811,N_29942);
or UO_3451 (O_3451,N_29836,N_29992);
xor UO_3452 (O_3452,N_29890,N_29974);
nor UO_3453 (O_3453,N_29824,N_29802);
or UO_3454 (O_3454,N_29992,N_29828);
nand UO_3455 (O_3455,N_29922,N_29960);
and UO_3456 (O_3456,N_29867,N_29834);
nor UO_3457 (O_3457,N_29902,N_29906);
xnor UO_3458 (O_3458,N_29928,N_29910);
nor UO_3459 (O_3459,N_29830,N_29846);
nand UO_3460 (O_3460,N_29836,N_29800);
or UO_3461 (O_3461,N_29802,N_29810);
and UO_3462 (O_3462,N_29894,N_29820);
xnor UO_3463 (O_3463,N_29920,N_29898);
or UO_3464 (O_3464,N_29874,N_29967);
and UO_3465 (O_3465,N_29985,N_29840);
nand UO_3466 (O_3466,N_29852,N_29905);
and UO_3467 (O_3467,N_29850,N_29987);
xor UO_3468 (O_3468,N_29865,N_29998);
nand UO_3469 (O_3469,N_29978,N_29962);
or UO_3470 (O_3470,N_29857,N_29940);
and UO_3471 (O_3471,N_29873,N_29882);
or UO_3472 (O_3472,N_29959,N_29935);
nor UO_3473 (O_3473,N_29883,N_29967);
xnor UO_3474 (O_3474,N_29865,N_29900);
and UO_3475 (O_3475,N_29801,N_29807);
or UO_3476 (O_3476,N_29878,N_29850);
xnor UO_3477 (O_3477,N_29870,N_29848);
xnor UO_3478 (O_3478,N_29904,N_29946);
nand UO_3479 (O_3479,N_29950,N_29999);
nor UO_3480 (O_3480,N_29813,N_29965);
and UO_3481 (O_3481,N_29835,N_29887);
xor UO_3482 (O_3482,N_29863,N_29865);
and UO_3483 (O_3483,N_29811,N_29892);
or UO_3484 (O_3484,N_29865,N_29994);
xnor UO_3485 (O_3485,N_29938,N_29801);
nor UO_3486 (O_3486,N_29968,N_29847);
xnor UO_3487 (O_3487,N_29890,N_29820);
xnor UO_3488 (O_3488,N_29927,N_29816);
or UO_3489 (O_3489,N_29943,N_29955);
and UO_3490 (O_3490,N_29968,N_29941);
xor UO_3491 (O_3491,N_29943,N_29941);
nand UO_3492 (O_3492,N_29996,N_29873);
nand UO_3493 (O_3493,N_29885,N_29839);
xnor UO_3494 (O_3494,N_29897,N_29929);
nand UO_3495 (O_3495,N_29852,N_29836);
nor UO_3496 (O_3496,N_29950,N_29899);
nand UO_3497 (O_3497,N_29876,N_29814);
or UO_3498 (O_3498,N_29840,N_29848);
xor UO_3499 (O_3499,N_29989,N_29832);
endmodule