module basic_2500_25000_3000_4_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18844,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18872,N_18873,N_18874,N_18875,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18930,N_18931,N_18932,N_18934,N_18935,N_18936,N_18937,N_18939,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19136,N_19137,N_19138,N_19139,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19192,N_19193,N_19194,N_19196,N_19197,N_19198,N_19199,N_19200,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19328,N_19329,N_19330,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19384,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19472,N_19473,N_19474,N_19475,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19672,N_19673,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20045,N_20046,N_20047,N_20048,N_20049,N_20051,N_20052,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20092,N_20093,N_20094,N_20096,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20346,N_20347,N_20349,N_20350,N_20351,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20629,N_20630,N_20631,N_20632,N_20633,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20858,N_20859,N_20860,N_20861,N_20862,N_20864,N_20865,N_20866,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20900,N_20901,N_20902,N_20903,N_20904,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21066,N_21067,N_21068,N_21069,N_21070,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21605,N_21606,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21833,N_21834,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22164,N_22165,N_22166,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22242,N_22243,N_22244,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22398,N_22399,N_22400,N_22401,N_22402,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22495,N_22496,N_22499,N_22500,N_22501,N_22502,N_22503,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22670,N_22671,N_22672,N_22673,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22877,N_22879,N_22880,N_22881,N_22882,N_22883,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22957,N_22958,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23408,N_23409,N_23410,N_23411,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23467,N_23468,N_23469,N_23470,N_23471,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23504,N_23505,N_23506,N_23507,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23577,N_23578,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23593,N_23594,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23637,N_23639,N_23640,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23819,N_23821,N_23822,N_23823,N_23824,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23911,N_23912,N_23913,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24171,N_24172,N_24173,N_24174,N_24175,N_24177,N_24178,N_24179,N_24180,N_24181,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24630,N_24631,N_24632,N_24634,N_24635,N_24636,N_24637,N_24638,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24868,N_24869,N_24870,N_24872,N_24873,N_24874,N_24875,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24928,N_24929,N_24930,N_24931,N_24932,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24999;
and U0 (N_0,In_2061,In_774);
nand U1 (N_1,In_1148,In_1835);
xnor U2 (N_2,In_717,In_1744);
and U3 (N_3,In_1796,In_1528);
xnor U4 (N_4,In_1572,In_670);
xnor U5 (N_5,In_140,In_2136);
and U6 (N_6,In_1998,In_2451);
or U7 (N_7,In_46,In_898);
xor U8 (N_8,In_302,In_1280);
nand U9 (N_9,In_1075,In_1548);
nor U10 (N_10,In_1306,In_1353);
and U11 (N_11,In_1347,In_835);
or U12 (N_12,In_1982,In_840);
nor U13 (N_13,In_674,In_690);
and U14 (N_14,In_1498,In_1650);
or U15 (N_15,In_2268,In_1319);
xor U16 (N_16,In_2360,In_2241);
nand U17 (N_17,In_938,In_130);
and U18 (N_18,In_267,In_2312);
nor U19 (N_19,In_1077,In_374);
xnor U20 (N_20,In_1341,In_2368);
xor U21 (N_21,In_2327,In_1657);
nor U22 (N_22,In_671,In_1905);
and U23 (N_23,In_752,In_26);
or U24 (N_24,In_413,In_2149);
nand U25 (N_25,In_1120,In_2191);
or U26 (N_26,In_2169,In_380);
xor U27 (N_27,In_494,In_458);
and U28 (N_28,In_1575,In_197);
and U29 (N_29,In_609,In_724);
xnor U30 (N_30,In_764,In_355);
nor U31 (N_31,In_1547,In_1252);
or U32 (N_32,In_820,In_1539);
xor U33 (N_33,In_1298,In_143);
or U34 (N_34,In_1625,In_2117);
and U35 (N_35,In_1587,In_1179);
nor U36 (N_36,In_836,In_2197);
or U37 (N_37,In_1397,In_842);
xnor U38 (N_38,In_1832,In_940);
or U39 (N_39,In_613,In_1065);
xor U40 (N_40,In_366,In_367);
nor U41 (N_41,In_1047,In_926);
and U42 (N_42,In_2185,In_877);
xor U43 (N_43,In_470,In_971);
nor U44 (N_44,In_1508,In_1874);
xnor U45 (N_45,In_1748,In_1914);
nand U46 (N_46,In_610,In_2464);
or U47 (N_47,In_2220,In_45);
and U48 (N_48,In_1685,In_1597);
nand U49 (N_49,In_727,In_2199);
and U50 (N_50,In_863,In_648);
nand U51 (N_51,In_2407,In_2218);
nand U52 (N_52,In_529,In_1787);
nand U53 (N_53,In_2290,In_2303);
nor U54 (N_54,In_386,In_1195);
and U55 (N_55,In_371,In_2144);
and U56 (N_56,In_340,In_2329);
and U57 (N_57,In_397,In_914);
and U58 (N_58,In_2043,In_281);
nand U59 (N_59,In_1724,In_2397);
nor U60 (N_60,In_2284,In_684);
and U61 (N_61,In_1689,In_291);
and U62 (N_62,In_1191,In_1901);
or U63 (N_63,In_1963,In_1576);
and U64 (N_64,In_362,In_1741);
and U65 (N_65,In_51,In_1590);
and U66 (N_66,In_1884,In_1023);
nor U67 (N_67,In_1115,In_1454);
or U68 (N_68,In_1544,In_1500);
nand U69 (N_69,In_521,In_955);
nor U70 (N_70,In_778,In_1612);
and U71 (N_71,In_1536,In_2016);
and U72 (N_72,In_704,In_672);
xor U73 (N_73,In_2021,In_813);
xnor U74 (N_74,In_1162,In_791);
nor U75 (N_75,In_663,In_2343);
nand U76 (N_76,In_777,In_358);
or U77 (N_77,In_2387,In_1947);
xnor U78 (N_78,In_2010,In_1211);
or U79 (N_79,In_447,In_1303);
nor U80 (N_80,In_731,In_2308);
nor U81 (N_81,In_2419,In_2210);
or U82 (N_82,In_608,In_1696);
or U83 (N_83,In_288,In_449);
and U84 (N_84,In_72,In_541);
nand U85 (N_85,In_584,In_80);
nor U86 (N_86,In_409,In_1531);
xor U87 (N_87,In_1763,In_153);
nor U88 (N_88,In_621,In_1903);
nor U89 (N_89,In_1995,In_2075);
and U90 (N_90,In_1395,In_2354);
nand U91 (N_91,In_878,In_210);
nand U92 (N_92,In_1526,In_2480);
nor U93 (N_93,In_1794,In_2055);
or U94 (N_94,In_796,In_2279);
and U95 (N_95,In_207,In_1402);
nor U96 (N_96,In_296,In_766);
and U97 (N_97,In_1878,In_1631);
nor U98 (N_98,In_1555,In_536);
nand U99 (N_99,In_1076,In_2215);
nor U100 (N_100,In_2007,In_351);
xor U101 (N_101,In_1557,In_1036);
or U102 (N_102,In_639,In_201);
nor U103 (N_103,In_199,In_1435);
or U104 (N_104,In_68,In_948);
or U105 (N_105,In_1061,In_2282);
nor U106 (N_106,In_2053,In_1579);
and U107 (N_107,In_2017,In_1320);
or U108 (N_108,In_1089,In_238);
xor U109 (N_109,In_991,In_1213);
nor U110 (N_110,In_1223,In_850);
nor U111 (N_111,In_559,In_1734);
xnor U112 (N_112,In_1289,In_248);
xor U113 (N_113,In_275,In_2320);
nor U114 (N_114,In_1846,In_178);
xnor U115 (N_115,In_2306,In_280);
nor U116 (N_116,In_183,In_2214);
nand U117 (N_117,In_1139,In_285);
or U118 (N_118,In_2334,In_533);
and U119 (N_119,In_1296,In_861);
and U120 (N_120,In_1387,In_925);
nand U121 (N_121,In_537,In_173);
nand U122 (N_122,In_693,In_718);
or U123 (N_123,In_93,In_1038);
or U124 (N_124,In_688,In_1189);
nand U125 (N_125,In_893,In_1552);
and U126 (N_126,In_2231,In_139);
nor U127 (N_127,In_1329,In_2233);
xor U128 (N_128,In_2195,In_1183);
or U129 (N_129,In_544,In_1440);
nor U130 (N_130,In_636,In_1840);
and U131 (N_131,In_947,In_1750);
and U132 (N_132,In_645,In_1591);
xnor U133 (N_133,In_901,In_2375);
nor U134 (N_134,In_401,In_792);
xor U135 (N_135,In_538,In_12);
or U136 (N_136,In_1181,In_982);
and U137 (N_137,In_120,In_799);
and U138 (N_138,In_1244,In_2478);
or U139 (N_139,In_431,In_1661);
xnor U140 (N_140,In_2009,In_1717);
or U141 (N_141,In_325,In_492);
nor U142 (N_142,In_370,In_763);
and U143 (N_143,In_307,In_1966);
nand U144 (N_144,In_1399,In_1375);
nand U145 (N_145,In_416,In_2158);
xnor U146 (N_146,In_2413,In_1735);
xor U147 (N_147,In_49,In_125);
xor U148 (N_148,In_1083,In_2322);
nand U149 (N_149,In_1326,In_475);
or U150 (N_150,In_1628,In_1176);
xor U151 (N_151,In_993,In_2270);
and U152 (N_152,In_700,In_1239);
nand U153 (N_153,In_1136,In_1423);
nor U154 (N_154,In_360,In_1324);
nand U155 (N_155,In_1865,In_2423);
nand U156 (N_156,In_719,In_174);
nor U157 (N_157,In_1825,In_776);
nor U158 (N_158,In_2065,In_2458);
nand U159 (N_159,In_463,In_558);
or U160 (N_160,In_2147,In_229);
nor U161 (N_161,In_1565,In_624);
and U162 (N_162,In_2484,In_865);
and U163 (N_163,In_341,In_977);
or U164 (N_164,In_1322,In_2159);
xnor U165 (N_165,In_1644,In_2142);
or U166 (N_166,In_2316,In_240);
and U167 (N_167,In_761,In_313);
xnor U168 (N_168,In_1664,In_2255);
nand U169 (N_169,In_958,In_1706);
xor U170 (N_170,In_1824,In_2091);
or U171 (N_171,In_2425,In_1566);
and U172 (N_172,In_1798,In_188);
nor U173 (N_173,In_2477,In_354);
xnor U174 (N_174,In_2467,In_1908);
nor U175 (N_175,In_802,In_1785);
or U176 (N_176,In_368,In_1659);
and U177 (N_177,In_2096,In_1809);
and U178 (N_178,In_2088,In_904);
nor U179 (N_179,In_954,In_819);
nor U180 (N_180,In_1906,In_9);
and U181 (N_181,In_377,In_1417);
and U182 (N_182,In_2294,In_650);
or U183 (N_183,In_1721,In_2223);
nand U184 (N_184,In_841,In_2039);
xor U185 (N_185,In_2276,In_641);
nand U186 (N_186,In_450,In_205);
nand U187 (N_187,In_448,In_1455);
xnor U188 (N_188,In_2200,In_1014);
and U189 (N_189,In_1126,In_398);
and U190 (N_190,In_432,In_582);
xor U191 (N_191,In_1935,In_1974);
nor U192 (N_192,In_2325,In_257);
nand U193 (N_193,In_344,In_2167);
nand U194 (N_194,In_960,In_2352);
or U195 (N_195,In_2066,In_1946);
nor U196 (N_196,In_716,In_1822);
and U197 (N_197,In_1524,In_2350);
and U198 (N_198,In_1254,In_1704);
or U199 (N_199,In_963,In_949);
nand U200 (N_200,In_1771,In_299);
xnor U201 (N_201,In_1215,In_177);
nor U202 (N_202,In_1134,In_1419);
xor U203 (N_203,In_1509,In_1339);
xor U204 (N_204,In_2495,In_381);
nand U205 (N_205,In_2379,In_666);
xor U206 (N_206,In_736,In_1499);
xnor U207 (N_207,In_874,In_2042);
nand U208 (N_208,In_200,In_2172);
or U209 (N_209,In_2374,In_456);
and U210 (N_210,In_1066,In_806);
or U211 (N_211,In_808,In_2309);
nand U212 (N_212,In_2445,In_1686);
xnor U213 (N_213,In_1662,In_198);
nor U214 (N_214,In_998,In_562);
nand U215 (N_215,In_1920,In_987);
nand U216 (N_216,In_1604,In_1198);
and U217 (N_217,In_618,In_1523);
xnor U218 (N_218,In_2001,In_437);
or U219 (N_219,In_1217,In_1068);
or U220 (N_220,In_1346,In_1609);
or U221 (N_221,In_742,In_1043);
or U222 (N_222,In_965,In_1106);
and U223 (N_223,In_647,In_1487);
nor U224 (N_224,In_1638,In_224);
nand U225 (N_225,In_2222,In_108);
nor U226 (N_226,In_2205,In_2110);
xnor U227 (N_227,In_1677,In_311);
xor U228 (N_228,In_2333,In_287);
nor U229 (N_229,In_654,In_91);
nor U230 (N_230,In_263,In_2485);
or U231 (N_231,In_899,In_543);
and U232 (N_232,In_1485,In_1277);
or U233 (N_233,In_968,In_896);
nand U234 (N_234,In_53,In_1328);
and U235 (N_235,In_260,In_894);
or U236 (N_236,In_662,In_1848);
or U237 (N_237,In_2038,In_1979);
and U238 (N_238,In_2119,In_2362);
and U239 (N_239,In_921,In_997);
and U240 (N_240,In_204,In_2137);
xor U241 (N_241,In_2494,In_1983);
or U242 (N_242,In_1196,In_1891);
nor U243 (N_243,In_1772,In_1535);
or U244 (N_244,In_1505,In_2217);
and U245 (N_245,In_1969,In_726);
nand U246 (N_246,In_2019,In_219);
xor U247 (N_247,In_709,In_1551);
or U248 (N_248,In_2126,In_103);
or U249 (N_249,In_811,In_1984);
or U250 (N_250,In_834,In_4);
and U251 (N_251,In_1960,In_873);
or U252 (N_252,In_887,In_637);
nor U253 (N_253,In_585,In_110);
or U254 (N_254,In_376,In_2022);
nor U255 (N_255,In_1538,In_1570);
nand U256 (N_256,In_597,In_713);
nor U257 (N_257,In_1224,In_234);
and U258 (N_258,In_314,In_326);
nor U259 (N_259,In_32,In_434);
nand U260 (N_260,In_509,In_56);
xnor U261 (N_261,In_950,In_1086);
and U262 (N_262,In_815,In_772);
or U263 (N_263,In_83,In_1948);
nor U264 (N_264,In_1517,In_746);
and U265 (N_265,In_1275,In_885);
nor U266 (N_266,In_1046,In_1085);
and U267 (N_267,In_990,In_321);
nand U268 (N_268,In_1924,In_1005);
and U269 (N_269,In_61,In_757);
or U270 (N_270,In_2174,In_1405);
xnor U271 (N_271,In_2092,In_906);
and U272 (N_272,In_943,In_105);
nand U273 (N_273,In_37,In_186);
nand U274 (N_274,In_383,In_1764);
nor U275 (N_275,In_145,In_1934);
xor U276 (N_276,In_312,In_620);
nor U277 (N_277,In_1063,In_1645);
and U278 (N_278,In_2184,In_102);
or U279 (N_279,In_821,In_1117);
nor U280 (N_280,In_817,In_1016);
and U281 (N_281,In_816,In_2435);
nand U282 (N_282,In_1710,In_635);
nand U283 (N_283,In_916,In_1917);
nand U284 (N_284,In_1774,In_1507);
nand U285 (N_285,In_452,In_1127);
or U286 (N_286,In_2086,In_1679);
xor U287 (N_287,In_106,In_1550);
nand U288 (N_288,In_436,In_747);
or U289 (N_289,In_1055,In_328);
nor U290 (N_290,In_85,In_1128);
or U291 (N_291,In_1406,In_1009);
xnor U292 (N_292,In_357,In_1894);
and U293 (N_293,In_631,In_13);
or U294 (N_294,In_823,In_41);
and U295 (N_295,In_1462,In_1413);
and U296 (N_296,In_1605,In_2121);
xor U297 (N_297,In_305,In_2289);
nand U298 (N_298,In_259,In_150);
and U299 (N_299,In_493,In_484);
nand U300 (N_300,In_441,In_593);
and U301 (N_301,In_1981,In_503);
xnor U302 (N_302,In_854,In_1335);
or U303 (N_303,In_1311,In_1541);
nand U304 (N_304,In_879,In_2351);
and U305 (N_305,In_1461,In_1242);
nand U306 (N_306,In_2094,In_504);
nor U307 (N_307,In_428,In_1390);
xnor U308 (N_308,In_162,In_1201);
or U309 (N_309,In_97,In_973);
xnor U310 (N_310,In_1173,In_782);
or U311 (N_311,In_208,In_369);
nand U312 (N_312,In_552,In_1453);
or U313 (N_313,In_2390,In_1119);
xor U314 (N_314,In_1997,In_1820);
nand U315 (N_315,In_1624,In_1877);
and U316 (N_316,In_525,In_828);
nor U317 (N_317,In_1409,In_395);
xor U318 (N_318,In_2287,In_333);
nor U319 (N_319,In_2421,In_384);
nand U320 (N_320,In_1141,In_2024);
and U321 (N_321,In_1931,In_1457);
nor U322 (N_322,In_2188,In_1048);
nand U323 (N_323,In_118,In_168);
nand U324 (N_324,In_625,In_1032);
nor U325 (N_325,In_510,In_20);
and U326 (N_326,In_1850,In_159);
xor U327 (N_327,In_1308,In_1826);
nor U328 (N_328,In_1837,In_2156);
nand U329 (N_329,In_2489,In_1815);
nand U330 (N_330,In_1022,In_1013);
nor U331 (N_331,In_2130,In_283);
or U332 (N_332,In_1806,In_2353);
or U333 (N_333,In_1937,In_1999);
or U334 (N_334,In_251,In_402);
and U335 (N_335,In_738,In_1779);
nand U336 (N_336,In_1688,In_1632);
nor U337 (N_337,In_485,In_890);
or U338 (N_338,In_2050,In_1245);
and U339 (N_339,In_1342,In_1648);
xor U340 (N_340,In_2426,In_1915);
and U341 (N_341,In_1200,In_2405);
nor U342 (N_342,In_771,In_535);
nor U343 (N_343,In_1610,In_107);
nor U344 (N_344,In_867,In_1425);
nor U345 (N_345,In_2078,In_19);
and U346 (N_346,In_419,In_2392);
xor U347 (N_347,In_1377,In_190);
or U348 (N_348,In_1232,In_2103);
or U349 (N_349,In_615,In_1113);
nand U350 (N_350,In_1116,In_2409);
and U351 (N_351,In_1384,In_710);
xor U352 (N_352,In_2030,In_414);
nand U353 (N_353,In_216,In_167);
xnor U354 (N_354,In_352,In_2492);
nand U355 (N_355,In_147,In_630);
xor U356 (N_356,In_981,In_1955);
nor U357 (N_357,In_1545,In_266);
or U358 (N_358,In_406,In_2240);
nand U359 (N_359,In_1140,In_1909);
or U360 (N_360,In_2356,In_1182);
nand U361 (N_361,In_427,In_1433);
nor U362 (N_362,In_1283,In_2281);
xor U363 (N_363,In_770,In_1554);
and U364 (N_364,In_524,In_520);
or U365 (N_365,In_683,In_1694);
nand U366 (N_366,In_2166,In_30);
nand U367 (N_367,In_545,In_1170);
xnor U368 (N_368,In_1705,In_2273);
nand U369 (N_369,In_780,In_286);
nor U370 (N_370,In_2148,In_1203);
xor U371 (N_371,In_98,In_274);
xnor U372 (N_372,In_182,In_2193);
xnor U373 (N_373,In_1081,In_1668);
nand U374 (N_374,In_2288,In_669);
xnor U375 (N_375,In_64,In_1615);
or U376 (N_376,In_391,In_1144);
nor U377 (N_377,In_2064,In_2278);
nand U378 (N_378,In_923,In_574);
nor U379 (N_379,In_195,In_1373);
xnor U380 (N_380,In_1887,In_268);
and U381 (N_381,In_750,In_1365);
xor U382 (N_382,In_1082,In_2162);
or U383 (N_383,In_2432,In_623);
or U384 (N_384,In_1775,In_1976);
or U385 (N_385,In_1760,In_203);
nand U386 (N_386,In_2378,In_1432);
xor U387 (N_387,In_1071,In_1466);
xor U388 (N_388,In_721,In_653);
nand U389 (N_389,In_1354,In_1227);
nor U390 (N_390,In_184,In_1060);
xnor U391 (N_391,In_1219,In_473);
nor U392 (N_392,In_556,In_1431);
nor U393 (N_393,In_497,In_304);
and U394 (N_394,In_1002,In_1284);
nor U395 (N_395,In_1749,In_711);
or U396 (N_396,In_569,In_1092);
nand U397 (N_397,In_1584,In_1852);
or U398 (N_398,In_1026,In_2109);
or U399 (N_399,In_660,In_1621);
xnor U400 (N_400,In_1029,In_759);
nand U401 (N_401,In_1681,In_228);
nand U402 (N_402,In_814,In_2328);
or U403 (N_403,In_1646,In_1330);
or U404 (N_404,In_443,In_1768);
nand U405 (N_405,In_2084,In_909);
xnor U406 (N_406,In_1429,In_1159);
nand U407 (N_407,In_586,In_1372);
xnor U408 (N_408,In_2439,In_855);
nand U409 (N_409,In_2283,In_1105);
nor U410 (N_410,In_1165,In_2443);
and U411 (N_411,In_2310,In_363);
and U412 (N_412,In_276,In_212);
and U413 (N_413,In_236,In_967);
or U414 (N_414,In_945,In_349);
nor U415 (N_415,In_629,In_364);
nor U416 (N_416,In_2372,In_1715);
and U417 (N_417,In_1147,In_2194);
xor U418 (N_418,In_476,In_2302);
xnor U419 (N_419,In_578,In_853);
nand U420 (N_420,In_1349,In_246);
and U421 (N_421,In_1109,In_1481);
xnor U422 (N_422,In_1701,In_423);
nand U423 (N_423,In_2450,In_644);
or U424 (N_424,In_90,In_712);
nor U425 (N_425,In_1961,In_918);
xnor U426 (N_426,In_58,In_1011);
nand U427 (N_427,In_194,In_471);
xor U428 (N_428,In_24,In_1965);
nor U429 (N_429,In_310,In_2151);
xor U430 (N_430,In_845,In_1758);
and U431 (N_431,In_1828,In_454);
and U432 (N_432,In_1589,In_2253);
nor U433 (N_433,In_913,In_1129);
xnor U434 (N_434,In_1504,In_353);
or U435 (N_435,In_540,In_2361);
or U436 (N_436,In_1844,In_622);
nor U437 (N_437,In_2460,In_2262);
xnor U438 (N_438,In_1279,In_1782);
or U439 (N_439,In_1344,In_1006);
nand U440 (N_440,In_1132,In_271);
xor U441 (N_441,In_2168,In_1593);
xor U442 (N_442,In_82,In_999);
nor U443 (N_443,In_1666,In_883);
or U444 (N_444,In_527,In_2326);
nand U445 (N_445,In_2072,In_1237);
xor U446 (N_446,In_2059,In_832);
or U447 (N_447,In_1178,In_1492);
nor U448 (N_448,In_289,In_1807);
and U449 (N_449,In_1996,In_1278);
and U450 (N_450,In_129,In_1040);
xor U451 (N_451,In_1292,In_465);
or U452 (N_452,In_786,In_2323);
and U453 (N_453,In_1110,In_679);
nor U454 (N_454,In_77,In_372);
nand U455 (N_455,In_1293,In_2422);
nand U456 (N_456,In_133,In_2363);
or U457 (N_457,In_705,In_2012);
xor U458 (N_458,In_1516,In_1441);
xnor U459 (N_459,In_2087,In_1230);
xor U460 (N_460,In_986,In_1450);
xnor U461 (N_461,In_1859,In_1167);
or U462 (N_462,In_849,In_1728);
and U463 (N_463,In_3,In_969);
nand U464 (N_464,In_1871,In_460);
or U465 (N_465,In_2002,In_1663);
nor U466 (N_466,In_1830,In_469);
and U467 (N_467,In_2133,In_563);
or U468 (N_468,In_1875,In_546);
or U469 (N_469,In_2277,In_1261);
nor U470 (N_470,In_348,In_160);
or U471 (N_471,In_2369,In_323);
and U472 (N_472,In_2348,In_1333);
nand U473 (N_473,In_1755,In_903);
and U474 (N_474,In_1379,In_2020);
nand U475 (N_475,In_1559,In_1357);
and U476 (N_476,In_646,In_2411);
nor U477 (N_477,In_1773,In_1037);
and U478 (N_478,In_1053,In_784);
or U479 (N_479,In_1345,In_1428);
nor U480 (N_480,In_1939,In_330);
nand U481 (N_481,In_1953,In_2018);
or U482 (N_482,In_466,In_831);
and U483 (N_483,In_1879,In_1912);
or U484 (N_484,In_1514,In_250);
and U485 (N_485,In_332,In_104);
xnor U486 (N_486,In_222,In_785);
or U487 (N_487,In_2376,In_175);
nor U488 (N_488,In_1582,In_233);
or U489 (N_489,In_2234,In_1988);
nand U490 (N_490,In_1421,In_2111);
or U491 (N_491,In_2101,In_1392);
nor U492 (N_492,In_607,In_665);
or U493 (N_493,In_1031,In_1367);
nand U494 (N_494,In_2139,In_2127);
and U495 (N_495,In_875,In_576);
and U496 (N_496,In_1904,In_1494);
nor U497 (N_497,In_435,In_2332);
xor U498 (N_498,In_935,In_788);
and U499 (N_499,In_642,In_1805);
nand U500 (N_500,In_775,In_375);
or U501 (N_501,In_1474,In_499);
or U502 (N_502,In_342,In_602);
nor U503 (N_503,In_300,In_1951);
nand U504 (N_504,In_189,In_1197);
or U505 (N_505,In_2377,In_2499);
and U506 (N_506,In_478,In_2123);
or U507 (N_507,In_753,In_63);
and U508 (N_508,In_2385,In_2206);
nor U509 (N_509,In_881,In_708);
and U510 (N_510,In_2083,In_2189);
or U511 (N_511,In_1751,In_1745);
and U512 (N_512,In_2260,In_40);
or U513 (N_513,In_185,In_1967);
and U514 (N_514,In_908,In_837);
nor U515 (N_515,In_1596,In_512);
nand U516 (N_516,In_2098,In_1056);
or U517 (N_517,In_508,In_2330);
and U518 (N_518,In_1332,In_2247);
xor U519 (N_519,In_1620,In_668);
nor U520 (N_520,In_1585,In_1427);
nand U521 (N_521,In_62,In_592);
and U522 (N_522,In_1381,In_1725);
xnor U523 (N_523,In_1549,In_421);
and U524 (N_524,In_2331,In_846);
and U525 (N_525,In_822,In_1674);
xor U526 (N_526,In_2453,In_729);
nor U527 (N_527,In_2227,In_826);
or U528 (N_528,In_633,In_1784);
or U529 (N_529,In_2099,In_1388);
xor U530 (N_530,In_343,In_1021);
nand U531 (N_531,In_1560,In_171);
nor U532 (N_532,In_1880,In_1723);
and U533 (N_533,In_1102,In_117);
or U534 (N_534,In_1972,In_1711);
xor U535 (N_535,In_1163,In_1430);
or U536 (N_536,In_2412,In_838);
or U537 (N_537,In_793,In_253);
or U538 (N_538,In_1030,In_2358);
nand U539 (N_539,In_1108,In_2297);
and U540 (N_540,In_1600,In_23);
nor U541 (N_541,In_1743,In_76);
and U542 (N_542,In_2498,In_1290);
nand U543 (N_543,In_567,In_1571);
or U544 (N_544,In_2080,In_1099);
or U545 (N_545,In_1893,In_1472);
nor U546 (N_546,In_65,In_8);
and U547 (N_547,In_1135,In_498);
or U548 (N_548,In_2182,In_1713);
nor U549 (N_549,In_480,In_2496);
xor U550 (N_550,In_420,In_561);
nor U551 (N_551,In_2011,In_1731);
and U552 (N_552,In_1697,In_1114);
and U553 (N_553,In_180,In_2389);
xnor U554 (N_554,In_1295,In_265);
nor U555 (N_555,In_564,In_844);
or U556 (N_556,In_1769,In_1118);
xor U557 (N_557,In_1358,In_2128);
nor U558 (N_558,In_571,In_1187);
nor U559 (N_559,In_590,In_2271);
and U560 (N_560,In_2198,In_1892);
nor U561 (N_561,In_803,In_2141);
xnor U562 (N_562,In_787,In_1511);
and U563 (N_563,In_1465,In_1288);
nand U564 (N_564,In_550,In_70);
nor U565 (N_565,In_1291,In_1540);
nand U566 (N_566,In_596,In_34);
nor U567 (N_567,In_396,In_329);
and U568 (N_568,In_1954,In_1351);
and U569 (N_569,In_1578,In_2077);
or U570 (N_570,In_2221,In_1000);
nand U571 (N_571,In_100,In_1321);
nand U572 (N_572,In_2132,In_2482);
nor U573 (N_573,In_1276,In_939);
xor U574 (N_574,In_1799,In_1817);
nand U575 (N_575,In_256,In_2429);
and U576 (N_576,In_526,In_941);
nand U577 (N_577,In_390,In_779);
and U578 (N_578,In_277,In_1452);
xor U579 (N_579,In_1336,In_1088);
xnor U580 (N_580,In_1226,In_2164);
nor U581 (N_581,In_467,In_2466);
or U582 (N_582,In_161,In_2497);
and U583 (N_583,In_1952,In_239);
xnor U584 (N_584,In_1352,In_1157);
nor U585 (N_585,In_1194,In_2176);
and U586 (N_586,In_39,In_2371);
nand U587 (N_587,In_18,In_1639);
nand U588 (N_588,In_1103,In_942);
nand U589 (N_589,In_1175,In_2062);
xnor U590 (N_590,In_2415,In_1757);
xnor U591 (N_591,In_2236,In_560);
xor U592 (N_592,In_1263,In_966);
and U593 (N_593,In_601,In_254);
nor U594 (N_594,In_2406,In_2140);
nand U595 (N_595,In_1980,In_851);
nor U596 (N_596,In_804,In_1155);
xnor U597 (N_597,In_1949,In_1338);
xor U598 (N_598,In_864,In_1193);
or U599 (N_599,In_2388,In_1315);
xor U600 (N_600,In_482,In_407);
nand U601 (N_601,In_1727,In_1041);
or U602 (N_602,In_1889,In_2380);
and U603 (N_603,In_163,In_1855);
xnor U604 (N_604,In_137,In_519);
xor U605 (N_605,In_1484,In_1302);
nand U606 (N_606,In_611,In_1537);
nor U607 (N_607,In_1285,In_897);
or U608 (N_608,In_2259,In_2447);
or U609 (N_609,In_2417,In_1897);
nand U610 (N_610,In_1172,In_627);
and U611 (N_611,In_1250,In_2357);
nor U612 (N_612,In_1216,In_440);
nor U613 (N_613,In_1309,In_856);
nor U614 (N_614,In_479,In_1255);
xnor U615 (N_615,In_1154,In_1190);
or U616 (N_616,In_1823,In_2051);
or U617 (N_617,In_292,In_511);
nand U618 (N_618,In_1438,In_359);
nand U619 (N_619,In_1121,In_2393);
and U620 (N_620,In_211,In_1527);
nand U621 (N_621,In_1045,In_1622);
xnor U622 (N_622,In_1218,In_483);
xor U623 (N_623,In_116,In_2396);
nand U624 (N_624,In_2023,In_1693);
nand U625 (N_625,In_697,In_2037);
nand U626 (N_626,In_1316,In_2367);
and U627 (N_627,In_2265,In_55);
nor U628 (N_628,In_1104,In_1810);
and U629 (N_629,In_1652,In_2232);
or U630 (N_630,In_1936,In_2252);
or U631 (N_631,In_2463,In_1364);
and U632 (N_632,In_1918,In_247);
nand U633 (N_633,In_1467,In_1214);
and U634 (N_634,In_2449,In_953);
nor U635 (N_635,In_1458,In_1883);
xnor U636 (N_636,In_1376,In_2455);
or U637 (N_637,In_1690,In_2317);
nor U638 (N_638,In_2044,In_1786);
nand U639 (N_639,In_1902,In_2454);
xor U640 (N_640,In_215,In_2448);
nand U641 (N_641,In_970,In_2060);
xor U642 (N_642,In_294,In_2324);
nand U643 (N_643,In_2301,In_1287);
nor U644 (N_644,In_1732,In_1495);
nand U645 (N_645,In_1112,In_551);
and U646 (N_646,In_1658,In_1923);
xor U647 (N_647,In_308,In_868);
xnor U648 (N_648,In_2031,In_565);
xor U649 (N_649,In_334,In_866);
nand U650 (N_650,In_1864,In_1530);
xor U651 (N_651,In_113,In_1192);
and U652 (N_652,In_1637,In_2089);
nand U653 (N_653,In_1862,In_47);
and U654 (N_654,In_1486,In_2486);
xor U655 (N_655,In_2428,In_566);
and U656 (N_656,In_2338,In_767);
or U657 (N_657,In_1256,In_2211);
and U658 (N_658,In_1094,In_11);
or U659 (N_659,In_2076,In_619);
nand U660 (N_660,In_715,In_2000);
xnor U661 (N_661,In_1304,In_2212);
or U662 (N_662,In_1678,In_1583);
or U663 (N_663,In_1635,In_144);
and U664 (N_664,In_762,In_1653);
xnor U665 (N_665,In_1074,In_1445);
or U666 (N_666,In_335,In_489);
xnor U667 (N_667,In_1122,In_2);
xnor U668 (N_668,In_1143,In_1456);
xnor U669 (N_669,In_394,In_2224);
nand U670 (N_670,In_884,In_1107);
nor U671 (N_671,In_1096,In_2095);
nand U672 (N_672,In_1222,In_1414);
or U673 (N_673,In_575,In_1137);
nand U674 (N_674,In_151,In_1739);
xor U675 (N_675,In_591,In_1133);
nand U676 (N_676,In_1070,In_242);
xor U677 (N_677,In_1707,In_983);
and U678 (N_678,In_154,In_732);
nor U679 (N_679,In_2135,In_972);
or U680 (N_680,In_317,In_1534);
xor U681 (N_681,In_825,In_14);
or U682 (N_682,In_739,In_1708);
or U683 (N_683,In_1776,In_1922);
nor U684 (N_684,In_1101,In_930);
nor U685 (N_685,In_1543,In_1919);
and U686 (N_686,In_2452,In_1851);
and U687 (N_687,In_453,In_2203);
xor U688 (N_688,In_1034,In_123);
nor U689 (N_689,In_1673,In_1647);
nand U690 (N_690,In_2264,In_149);
and U691 (N_691,In_2033,In_1401);
xor U692 (N_692,In_142,In_301);
nor U693 (N_693,In_2472,In_192);
nand U694 (N_694,In_1795,In_255);
nor U695 (N_695,In_1649,In_1595);
or U696 (N_696,In_1881,In_2219);
xor U697 (N_697,In_264,In_1091);
or U698 (N_698,In_221,In_1362);
or U699 (N_699,In_2090,In_2171);
nor U700 (N_700,In_1766,In_232);
nor U701 (N_701,In_2364,In_933);
or U702 (N_702,In_87,In_2237);
or U703 (N_703,In_272,In_1443);
xor U704 (N_704,In_2335,In_1420);
xnor U705 (N_705,In_1271,In_1503);
xnor U706 (N_706,In_694,In_67);
or U707 (N_707,In_2049,In_2468);
xor U708 (N_708,In_1793,In_681);
nand U709 (N_709,In_1310,In_1861);
nor U710 (N_710,In_2398,In_600);
xor U711 (N_711,In_2471,In_1380);
nor U712 (N_712,In_322,In_1863);
nand U713 (N_713,In_1248,In_319);
or U714 (N_714,In_809,In_410);
or U715 (N_715,In_985,In_2441);
nand U716 (N_716,In_1238,In_2008);
nor U717 (N_717,In_1940,In_661);
xnor U718 (N_718,In_862,In_807);
nor U719 (N_719,In_2216,In_298);
nand U720 (N_720,In_2298,In_976);
or U721 (N_721,In_438,In_500);
xnor U722 (N_722,In_2226,In_2456);
nand U723 (N_723,In_2355,In_1158);
or U724 (N_724,In_911,In_439);
or U725 (N_725,In_1594,In_517);
nand U726 (N_726,In_2267,In_1383);
nand U727 (N_727,In_2105,In_706);
and U728 (N_728,In_614,In_1761);
xnor U729 (N_729,In_269,In_403);
xor U730 (N_730,In_572,In_880);
or U731 (N_731,In_895,In_1281);
nand U732 (N_732,In_2120,In_111);
nand U733 (N_733,In_1833,In_1259);
nand U734 (N_734,In_1636,In_425);
or U735 (N_735,In_338,In_632);
nor U736 (N_736,In_1424,In_946);
or U737 (N_737,In_1251,In_1506);
and U738 (N_738,In_783,In_931);
nand U739 (N_739,In_1973,In_33);
or U740 (N_740,In_1003,In_1777);
nand U741 (N_741,In_2160,In_2438);
xnor U742 (N_742,In_1149,In_2183);
xor U743 (N_743,In_2444,In_1619);
nor U744 (N_744,In_1225,In_1001);
or U745 (N_745,In_22,In_1925);
and U746 (N_746,In_1231,In_800);
nand U747 (N_747,In_1437,In_975);
xnor U748 (N_748,In_548,In_889);
and U749 (N_749,In_2483,In_2479);
nand U750 (N_750,In_801,In_699);
xnor U751 (N_751,In_1359,In_345);
xor U752 (N_752,In_213,In_2314);
xor U753 (N_753,In_664,In_978);
and U754 (N_754,In_1482,In_743);
xor U755 (N_755,In_2437,In_1228);
nor U756 (N_756,In_1403,In_6);
xnor U757 (N_757,In_659,In_2112);
and U758 (N_758,In_2440,In_2047);
nand U759 (N_759,In_0,In_1956);
nor U760 (N_760,In_1651,In_2246);
and U761 (N_761,In_1235,In_1928);
nand U762 (N_762,In_790,In_1627);
or U763 (N_763,In_860,In_1601);
xor U764 (N_764,In_2280,In_1186);
xor U765 (N_765,In_1802,In_824);
xnor U766 (N_766,In_496,In_48);
nor U767 (N_767,In_399,In_1490);
xor U768 (N_768,In_872,In_749);
or U769 (N_769,In_1518,In_733);
and U770 (N_770,In_2243,In_1598);
nand U771 (N_771,In_974,In_744);
nor U772 (N_772,In_2373,In_871);
and U773 (N_773,In_134,In_1067);
nor U774 (N_774,In_1209,In_922);
and U775 (N_775,In_1035,In_1702);
nor U776 (N_776,In_1130,In_2143);
and U777 (N_777,In_1028,In_2175);
nor U778 (N_778,In_626,In_1297);
xor U779 (N_779,In_680,In_1860);
xor U780 (N_780,In_1546,In_2349);
and U781 (N_781,In_2213,In_1356);
and U782 (N_782,In_1991,In_2269);
nand U783 (N_783,In_2015,In_2005);
nor U784 (N_784,In_1910,In_1899);
nand U785 (N_785,In_331,In_758);
and U786 (N_786,In_1145,In_2116);
nor U787 (N_787,In_598,In_1079);
or U788 (N_788,In_472,In_382);
nand U789 (N_789,In_385,In_2296);
nand U790 (N_790,In_2311,In_1558);
nand U791 (N_791,In_2266,In_89);
nand U792 (N_792,In_658,In_121);
or U793 (N_793,In_293,In_1470);
nand U794 (N_794,In_2465,In_2074);
nand U795 (N_795,In_964,In_555);
and U796 (N_796,In_994,In_686);
xor U797 (N_797,In_1404,In_523);
and U798 (N_798,In_1845,In_2319);
nor U799 (N_799,In_2244,In_1361);
nand U800 (N_800,In_1312,In_1475);
and U801 (N_801,In_1854,In_1412);
nand U802 (N_802,In_2258,In_870);
xnor U803 (N_803,In_696,In_888);
nand U804 (N_804,In_2336,In_1781);
xor U805 (N_805,In_1703,In_278);
nand U806 (N_806,In_1941,In_2152);
and U807 (N_807,In_2082,In_1174);
xnor U808 (N_808,In_1207,In_1989);
and U809 (N_809,In_714,In_1561);
xor U810 (N_810,In_2416,In_1268);
and U811 (N_811,In_2370,In_373);
xor U812 (N_812,In_1184,In_603);
nor U813 (N_813,In_442,In_1229);
or U814 (N_814,In_52,In_491);
xor U815 (N_815,In_2125,In_1);
nand U816 (N_816,In_1801,In_1348);
and U817 (N_817,In_2207,In_2414);
nor U818 (N_818,In_464,In_17);
nor U819 (N_819,In_379,In_1718);
nor U820 (N_820,In_2034,In_95);
nor U821 (N_821,In_769,In_2180);
and U822 (N_822,In_1900,In_751);
nor U823 (N_823,In_1586,In_1095);
nor U824 (N_824,In_1847,In_1987);
nand U825 (N_825,In_1426,In_490);
nor U826 (N_826,In_1930,In_1202);
or U827 (N_827,In_1747,In_1943);
nand U828 (N_828,In_1234,In_1762);
nand U829 (N_829,In_461,In_1978);
nand U830 (N_830,In_1273,In_912);
nand U831 (N_831,In_2069,In_1355);
nor U832 (N_832,In_1299,In_187);
xor U833 (N_833,In_531,In_2071);
xor U834 (N_834,In_446,In_1410);
or U835 (N_835,In_1926,In_1574);
xnor U836 (N_836,In_638,In_318);
nand U837 (N_837,In_996,In_1340);
or U838 (N_838,In_2402,In_2124);
nand U839 (N_839,In_2481,In_1123);
or U840 (N_840,In_655,In_430);
xnor U841 (N_841,In_1675,In_1240);
nor U842 (N_842,In_75,In_339);
nor U843 (N_843,In_361,In_2347);
or U844 (N_844,In_936,In_910);
nand U845 (N_845,In_1479,In_667);
and U846 (N_846,In_1233,In_2304);
nor U847 (N_847,In_1460,In_900);
xnor U848 (N_848,In_1501,In_2134);
nor U849 (N_849,In_1640,In_2004);
or U850 (N_850,In_1606,In_1712);
or U851 (N_851,In_2431,In_2261);
and U852 (N_852,In_230,In_1366);
xor U853 (N_853,In_346,In_995);
and U854 (N_854,In_1567,In_588);
nand U855 (N_855,In_60,In_1876);
xnor U856 (N_856,In_2190,In_1532);
xor U857 (N_857,In_905,In_859);
nand U858 (N_858,In_2473,In_634);
and U859 (N_859,In_1641,In_2313);
and U860 (N_860,In_2115,In_2300);
nor U861 (N_861,In_412,In_1722);
xor U862 (N_862,In_225,In_1266);
nor U863 (N_863,In_35,In_2491);
and U864 (N_864,In_1436,In_959);
xor U865 (N_865,In_2291,In_417);
or U866 (N_866,In_115,In_723);
nor U867 (N_867,In_1272,In_1971);
nor U868 (N_868,In_1788,In_141);
nor U869 (N_869,In_243,In_43);
and U870 (N_870,In_1665,In_692);
or U871 (N_871,In_1746,In_2196);
or U872 (N_872,In_1607,In_2490);
and U873 (N_873,In_2046,In_1869);
xor U874 (N_874,In_71,In_164);
nand U875 (N_875,In_57,In_2251);
nor U876 (N_876,In_852,In_1151);
and U877 (N_877,In_2436,In_2365);
or U878 (N_878,In_2238,In_1736);
xor U879 (N_879,In_701,In_1726);
or U880 (N_880,In_1890,In_2394);
xor U881 (N_881,In_1882,In_745);
and U882 (N_882,In_1740,In_1039);
and U883 (N_883,In_984,In_415);
xor U884 (N_884,In_583,In_928);
xor U885 (N_885,In_128,In_2165);
or U886 (N_886,In_1834,In_1733);
xor U887 (N_887,In_2150,In_337);
and U888 (N_888,In_2003,In_1098);
and U889 (N_889,In_2225,In_1059);
nor U890 (N_890,In_2461,In_768);
xnor U891 (N_891,In_829,In_5);
or U892 (N_892,In_2056,In_1153);
xor U893 (N_893,In_1838,In_1400);
and U894 (N_894,In_929,In_577);
nor U895 (N_895,In_1208,In_2462);
xnor U896 (N_896,In_156,In_1054);
and U897 (N_897,In_2118,In_324);
nor U898 (N_898,In_1888,In_2107);
or U899 (N_899,In_245,In_2321);
xor U900 (N_900,In_934,In_1626);
nand U901 (N_901,In_1780,In_1958);
or U902 (N_902,In_1325,In_2305);
nand U903 (N_903,In_1730,In_481);
and U904 (N_904,In_2208,In_1811);
and U905 (N_905,In_1792,In_534);
xor U906 (N_906,In_2025,In_42);
nor U907 (N_907,In_515,In_1913);
or U908 (N_908,In_961,In_176);
nor U909 (N_909,In_741,In_1737);
xor U910 (N_910,In_29,In_1778);
nand U911 (N_911,In_765,In_702);
xor U912 (N_912,In_1568,In_1642);
or U913 (N_913,In_1993,In_2057);
and U914 (N_914,In_2249,In_1687);
and U915 (N_915,In_748,In_1857);
nand U916 (N_916,In_1282,In_2292);
nand U917 (N_917,In_295,In_1269);
xnor U918 (N_918,In_193,In_1073);
xnor U919 (N_919,In_756,In_798);
nor U920 (N_920,In_857,In_1267);
and U921 (N_921,In_389,In_2032);
nand U922 (N_922,In_1634,In_1617);
and U923 (N_923,In_528,In_547);
xnor U924 (N_924,In_262,In_226);
or U925 (N_925,In_1301,In_2173);
and U926 (N_926,In_781,In_249);
nor U927 (N_927,In_1418,In_573);
or U928 (N_928,In_1742,In_2408);
xor U929 (N_929,In_2131,In_2476);
nand U930 (N_930,In_920,In_992);
or U931 (N_931,In_172,In_1152);
nand U932 (N_932,In_1142,In_1012);
or U933 (N_933,In_1394,In_1770);
or U934 (N_934,In_2028,In_1819);
or U935 (N_935,In_2493,In_1015);
nor U936 (N_936,In_1611,In_1699);
xor U937 (N_937,In_2400,In_1253);
and U938 (N_938,In_1416,In_2399);
nor U939 (N_939,In_594,In_728);
xor U940 (N_940,In_1078,In_2192);
and U941 (N_941,In_2488,In_495);
nand U942 (N_942,In_689,In_218);
and U943 (N_943,In_1468,In_1483);
nand U944 (N_944,In_698,In_400);
or U945 (N_945,In_2386,In_886);
nor U946 (N_946,In_1258,In_1633);
or U947 (N_947,In_932,In_2097);
xnor U948 (N_948,In_649,In_505);
and U949 (N_949,In_1448,In_252);
or U950 (N_950,In_1790,In_73);
nor U951 (N_951,In_36,In_408);
nor U952 (N_952,In_2433,In_1100);
nand U953 (N_953,In_2154,In_2344);
nor U954 (N_954,In_1221,In_2146);
nand U955 (N_955,In_1274,In_1867);
or U956 (N_956,In_2138,In_1169);
nand U957 (N_957,In_1700,In_773);
nand U958 (N_958,In_206,In_2187);
nor U959 (N_959,In_1754,In_99);
xnor U960 (N_960,In_1262,In_1049);
or U961 (N_961,In_2401,In_2469);
and U962 (N_962,In_2040,In_1895);
nand U963 (N_963,In_1812,In_1446);
or U964 (N_964,In_1360,In_1449);
and U965 (N_965,In_1950,In_988);
nand U966 (N_966,In_1313,In_606);
nor U967 (N_967,In_1856,In_1719);
and U968 (N_968,In_797,In_1247);
xnor U969 (N_969,In_2446,In_1317);
and U970 (N_970,In_2250,In_1886);
and U971 (N_971,In_1602,In_1921);
nand U972 (N_972,In_1672,In_1024);
or U973 (N_973,In_1964,In_88);
xnor U974 (N_974,In_2285,In_2228);
or U975 (N_975,In_1323,In_2014);
nor U976 (N_976,In_1185,In_1393);
or U977 (N_977,In_2181,In_2245);
xor U978 (N_978,In_170,In_2155);
or U979 (N_979,In_273,In_2340);
or U980 (N_980,In_2286,In_1525);
and U981 (N_981,In_1522,In_1471);
and U982 (N_982,In_1025,In_818);
nor U983 (N_983,In_81,In_1827);
and U984 (N_984,In_1408,In_237);
and U985 (N_985,In_1415,In_2346);
and U986 (N_986,In_1767,In_122);
xnor U987 (N_987,In_1469,In_138);
xor U988 (N_988,In_16,In_445);
xor U989 (N_989,In_2315,In_707);
xnor U990 (N_990,In_2081,In_1087);
xnor U991 (N_991,In_2179,In_157);
and U992 (N_992,In_241,In_1050);
nor U993 (N_993,In_1146,In_1260);
nor U994 (N_994,In_1180,In_915);
xor U995 (N_995,In_109,In_979);
and U996 (N_996,In_2239,In_956);
and U997 (N_997,In_1220,In_2235);
nor U998 (N_998,In_1870,In_135);
or U999 (N_999,In_131,In_651);
or U1000 (N_1000,In_1716,In_2299);
or U1001 (N_1001,In_2383,In_315);
nand U1002 (N_1002,In_2427,In_2341);
and U1003 (N_1003,In_1808,In_794);
xnor U1004 (N_1004,In_1007,In_1350);
nand U1005 (N_1005,In_919,In_1300);
nand U1006 (N_1006,In_1804,In_1439);
xnor U1007 (N_1007,In_1569,In_1434);
or U1008 (N_1008,In_2384,In_1519);
nand U1009 (N_1009,In_1156,In_2178);
nand U1010 (N_1010,In_1872,In_1752);
nor U1011 (N_1011,In_1588,In_1111);
and U1012 (N_1012,In_1473,In_387);
nor U1013 (N_1013,In_1520,In_1051);
or U1014 (N_1014,In_297,In_2263);
and U1015 (N_1015,In_1343,In_2201);
or U1016 (N_1016,In_1853,In_1843);
or U1017 (N_1017,In_1660,In_640);
or U1018 (N_1018,In_136,In_1010);
xor U1019 (N_1019,In_2366,In_2307);
nor U1020 (N_1020,In_1676,In_839);
and U1021 (N_1021,In_418,In_1797);
nor U1022 (N_1022,In_1382,In_2006);
nor U1023 (N_1023,In_581,In_1680);
or U1024 (N_1024,In_2070,In_2248);
or U1025 (N_1025,In_2202,In_687);
and U1026 (N_1026,In_2170,In_1985);
nor U1027 (N_1027,In_557,In_1422);
nor U1028 (N_1028,In_94,In_1667);
and U1029 (N_1029,In_506,In_2345);
or U1030 (N_1030,In_501,In_2403);
nand U1031 (N_1031,In_1533,In_2382);
or U1032 (N_1032,In_1821,In_1264);
nor U1033 (N_1033,In_1171,In_1932);
or U1034 (N_1034,In_1800,In_725);
nor U1035 (N_1035,In_1698,In_1265);
or U1036 (N_1036,In_1057,In_119);
nor U1037 (N_1037,In_2106,In_468);
and U1038 (N_1038,In_1803,In_1097);
nor U1039 (N_1039,In_158,In_1368);
xor U1040 (N_1040,In_1161,In_1166);
xor U1041 (N_1041,In_2391,In_1205);
nand U1042 (N_1042,In_223,In_2153);
or U1043 (N_1043,In_1643,In_451);
and U1044 (N_1044,In_502,In_2256);
xnor U1045 (N_1045,In_132,In_1616);
and U1046 (N_1046,In_847,In_740);
or U1047 (N_1047,In_539,In_1305);
and U1048 (N_1048,In_907,In_166);
nand U1049 (N_1049,In_589,In_695);
and U1050 (N_1050,In_1942,In_1370);
nand U1051 (N_1051,In_1072,In_869);
or U1052 (N_1052,In_1916,In_84);
or U1053 (N_1053,In_1818,In_2475);
nand U1054 (N_1054,In_1389,In_1873);
and U1055 (N_1055,In_1695,In_1849);
and U1056 (N_1056,In_554,In_1959);
nor U1057 (N_1057,In_2418,In_2145);
or U1058 (N_1058,In_1896,In_2474);
nand U1059 (N_1059,In_682,In_1246);
nor U1060 (N_1060,In_2063,In_1670);
xor U1061 (N_1061,In_579,In_1020);
nand U1062 (N_1062,In_1911,In_2430);
xor U1063 (N_1063,In_1188,In_2073);
xor U1064 (N_1064,In_282,In_902);
nand U1065 (N_1065,In_1337,In_1396);
nand U1066 (N_1066,In_2257,In_810);
or U1067 (N_1067,In_848,In_79);
xnor U1068 (N_1068,In_1019,In_2293);
or U1069 (N_1069,In_1783,In_7);
and U1070 (N_1070,In_179,In_1720);
or U1071 (N_1071,In_1150,In_830);
and U1072 (N_1072,In_2100,In_1199);
nor U1073 (N_1073,In_1378,In_1044);
nor U1074 (N_1074,In_2104,In_1374);
or U1075 (N_1075,In_15,In_2085);
or U1076 (N_1076,In_2186,In_1841);
and U1077 (N_1077,In_320,In_1477);
and U1078 (N_1078,In_38,In_196);
or U1079 (N_1079,In_2442,In_487);
or U1080 (N_1080,In_514,In_927);
or U1081 (N_1081,In_1709,In_27);
or U1082 (N_1082,In_1564,In_2029);
nor U1083 (N_1083,In_486,In_1407);
or U1084 (N_1084,In_522,In_843);
xor U1085 (N_1085,In_2163,In_2058);
xor U1086 (N_1086,In_530,In_513);
and U1087 (N_1087,In_1411,In_2242);
nand U1088 (N_1088,In_2420,In_1459);
or U1089 (N_1089,In_457,In_675);
nand U1090 (N_1090,In_734,In_1385);
or U1091 (N_1091,In_944,In_1371);
xnor U1092 (N_1092,In_1614,In_2036);
nor U1093 (N_1093,In_59,In_617);
xnor U1094 (N_1094,In_1866,In_1270);
xnor U1095 (N_1095,In_1618,In_1691);
xor U1096 (N_1096,In_1608,In_258);
and U1097 (N_1097,In_1008,In_2457);
and U1098 (N_1098,In_1553,In_227);
nor U1099 (N_1099,In_429,In_2067);
and U1100 (N_1100,In_25,In_411);
nand U1101 (N_1101,In_1491,In_316);
xor U1102 (N_1102,In_44,In_1463);
or U1103 (N_1103,In_2470,In_444);
and U1104 (N_1104,In_604,In_1629);
xnor U1105 (N_1105,In_1164,In_126);
xor U1106 (N_1106,In_261,In_703);
and U1107 (N_1107,In_1603,In_1938);
xnor U1108 (N_1108,In_2318,In_1968);
or U1109 (N_1109,In_1580,In_2129);
or U1110 (N_1110,In_952,In_336);
xor U1111 (N_1111,In_2229,In_549);
nor U1112 (N_1112,In_1529,In_306);
or U1113 (N_1113,In_279,In_1369);
nor U1114 (N_1114,In_1513,In_1975);
nor U1115 (N_1115,In_676,In_691);
and U1116 (N_1116,In_1521,In_1017);
or U1117 (N_1117,In_673,In_1478);
or U1118 (N_1118,In_404,In_2013);
and U1119 (N_1119,In_1630,In_1160);
nand U1120 (N_1120,In_169,In_1334);
nor U1121 (N_1121,In_1868,In_152);
nor U1122 (N_1122,In_209,In_1033);
nand U1123 (N_1123,In_92,In_722);
xor U1124 (N_1124,In_1684,In_1496);
nand U1125 (N_1125,In_155,In_1168);
or U1126 (N_1126,In_1476,In_1756);
xnor U1127 (N_1127,In_220,In_1813);
or U1128 (N_1128,In_891,In_2204);
and U1129 (N_1129,In_477,In_1125);
and U1130 (N_1130,In_393,In_1493);
nor U1131 (N_1131,In_962,In_1398);
or U1132 (N_1132,In_2048,In_217);
and U1133 (N_1133,In_678,In_1018);
xor U1134 (N_1134,In_1502,In_2424);
xnor U1135 (N_1135,In_833,In_2381);
nand U1136 (N_1136,In_1080,In_365);
nor U1137 (N_1137,In_730,In_2295);
or U1138 (N_1138,In_2041,In_21);
or U1139 (N_1139,In_532,In_735);
and U1140 (N_1140,In_112,In_2254);
nor U1141 (N_1141,In_231,In_1990);
nand U1142 (N_1142,In_378,In_2337);
and U1143 (N_1143,In_2054,In_2052);
and U1144 (N_1144,In_424,In_812);
nor U1145 (N_1145,In_1042,In_1655);
nor U1146 (N_1146,In_1004,In_146);
xnor U1147 (N_1147,In_392,In_270);
or U1148 (N_1148,In_474,In_1957);
or U1149 (N_1149,In_1515,In_2122);
or U1150 (N_1150,In_917,In_1992);
or U1151 (N_1151,In_643,In_1692);
nand U1152 (N_1152,In_2161,In_1789);
or U1153 (N_1153,In_1177,In_1489);
nand U1154 (N_1154,In_685,In_181);
and U1155 (N_1155,In_1212,In_1986);
nand U1156 (N_1156,In_1831,In_1654);
nand U1157 (N_1157,In_1656,In_507);
nor U1158 (N_1158,In_2026,In_605);
xnor U1159 (N_1159,In_1962,In_1442);
nor U1160 (N_1160,In_2157,In_1836);
xor U1161 (N_1161,In_124,In_1907);
nor U1162 (N_1162,In_760,In_1842);
nand U1163 (N_1163,In_2108,In_426);
nor U1164 (N_1164,In_327,In_580);
nand U1165 (N_1165,In_1977,In_1765);
xor U1166 (N_1166,In_542,In_2102);
or U1167 (N_1167,In_876,In_2114);
nor U1168 (N_1168,In_924,In_96);
or U1169 (N_1169,In_980,In_1241);
or U1170 (N_1170,In_1249,In_1327);
and U1171 (N_1171,In_1447,In_1753);
and U1172 (N_1172,In_2035,In_754);
or U1173 (N_1173,In_1994,In_737);
nor U1174 (N_1174,In_1480,In_462);
or U1175 (N_1175,In_2404,In_2093);
and U1176 (N_1176,In_2487,In_1236);
or U1177 (N_1177,In_612,In_1204);
nor U1178 (N_1178,In_54,In_1577);
or U1179 (N_1179,In_1759,In_1444);
xor U1180 (N_1180,In_1391,In_516);
and U1181 (N_1181,In_1581,In_101);
or U1182 (N_1182,In_892,In_284);
or U1183 (N_1183,In_214,In_1131);
xnor U1184 (N_1184,In_31,In_1451);
or U1185 (N_1185,In_1138,In_347);
nand U1186 (N_1186,In_356,In_235);
nor U1187 (N_1187,In_2113,In_805);
nor U1188 (N_1188,In_244,In_1898);
or U1189 (N_1189,In_1562,In_127);
nand U1190 (N_1190,In_2230,In_1363);
or U1191 (N_1191,In_1318,In_455);
xor U1192 (N_1192,In_2339,In_2459);
or U1193 (N_1193,In_1839,In_2410);
and U1194 (N_1194,In_1669,In_2079);
nor U1195 (N_1195,In_1858,In_1682);
and U1196 (N_1196,In_1090,In_1592);
or U1197 (N_1197,In_587,In_1512);
nor U1198 (N_1198,In_720,In_1314);
nand U1199 (N_1199,In_518,In_652);
nor U1200 (N_1200,In_459,In_1497);
and U1201 (N_1201,In_599,In_1944);
nand U1202 (N_1202,In_165,In_488);
nor U1203 (N_1203,In_1563,In_309);
xor U1204 (N_1204,In_568,In_148);
nor U1205 (N_1205,In_789,In_957);
nand U1206 (N_1206,In_290,In_2272);
and U1207 (N_1207,In_1052,In_795);
and U1208 (N_1208,In_2068,In_628);
or U1209 (N_1209,In_1599,In_1464);
nor U1210 (N_1210,In_69,In_1064);
nand U1211 (N_1211,In_422,In_1386);
and U1212 (N_1212,In_989,In_1510);
nor U1213 (N_1213,In_1556,In_1573);
nand U1214 (N_1214,In_405,In_1093);
xnor U1215 (N_1215,In_1069,In_656);
nand U1216 (N_1216,In_827,In_951);
or U1217 (N_1217,In_858,In_1058);
and U1218 (N_1218,In_1623,In_1729);
nand U1219 (N_1219,In_616,In_1613);
or U1220 (N_1220,In_1814,In_1027);
nor U1221 (N_1221,In_1542,In_1885);
nand U1222 (N_1222,In_433,In_1243);
xor U1223 (N_1223,In_595,In_2434);
and U1224 (N_1224,In_1738,In_1829);
and U1225 (N_1225,In_350,In_1084);
or U1226 (N_1226,In_657,In_1816);
xor U1227 (N_1227,In_1331,In_10);
and U1228 (N_1228,In_2395,In_1929);
nor U1229 (N_1229,In_2359,In_74);
nand U1230 (N_1230,In_191,In_2275);
and U1231 (N_1231,In_78,In_1206);
and U1232 (N_1232,In_50,In_114);
or U1233 (N_1233,In_1062,In_1945);
xnor U1234 (N_1234,In_1671,In_2027);
and U1235 (N_1235,In_755,In_66);
xor U1236 (N_1236,In_1286,In_1488);
nand U1237 (N_1237,In_1210,In_2177);
nor U1238 (N_1238,In_1683,In_677);
xnor U1239 (N_1239,In_388,In_1933);
xor U1240 (N_1240,In_1257,In_1927);
nor U1241 (N_1241,In_202,In_2274);
or U1242 (N_1242,In_1970,In_553);
or U1243 (N_1243,In_1714,In_303);
nand U1244 (N_1244,In_570,In_1294);
or U1245 (N_1245,In_937,In_2209);
xnor U1246 (N_1246,In_1791,In_86);
nor U1247 (N_1247,In_2342,In_28);
and U1248 (N_1248,In_1307,In_882);
nor U1249 (N_1249,In_1124,In_2045);
nor U1250 (N_1250,In_926,In_2436);
or U1251 (N_1251,In_2019,In_1848);
or U1252 (N_1252,In_390,In_130);
nand U1253 (N_1253,In_1003,In_830);
nand U1254 (N_1254,In_1014,In_2150);
nor U1255 (N_1255,In_616,In_585);
nor U1256 (N_1256,In_2069,In_120);
nor U1257 (N_1257,In_1729,In_303);
nor U1258 (N_1258,In_1471,In_1287);
xor U1259 (N_1259,In_903,In_1597);
nor U1260 (N_1260,In_26,In_653);
and U1261 (N_1261,In_1627,In_1001);
nor U1262 (N_1262,In_654,In_453);
xor U1263 (N_1263,In_117,In_1369);
xor U1264 (N_1264,In_344,In_2360);
xor U1265 (N_1265,In_1114,In_574);
and U1266 (N_1266,In_40,In_2161);
or U1267 (N_1267,In_899,In_1447);
xnor U1268 (N_1268,In_2064,In_1915);
nor U1269 (N_1269,In_599,In_1647);
xnor U1270 (N_1270,In_426,In_202);
xor U1271 (N_1271,In_1872,In_1346);
xnor U1272 (N_1272,In_28,In_2261);
xnor U1273 (N_1273,In_2247,In_715);
nand U1274 (N_1274,In_1226,In_2277);
nor U1275 (N_1275,In_1106,In_702);
nor U1276 (N_1276,In_55,In_159);
and U1277 (N_1277,In_1228,In_1173);
xor U1278 (N_1278,In_1315,In_2355);
and U1279 (N_1279,In_1588,In_2493);
and U1280 (N_1280,In_2391,In_666);
nand U1281 (N_1281,In_236,In_2097);
and U1282 (N_1282,In_1416,In_1056);
nand U1283 (N_1283,In_867,In_1789);
nor U1284 (N_1284,In_1396,In_2163);
and U1285 (N_1285,In_2493,In_2270);
and U1286 (N_1286,In_1818,In_1683);
nor U1287 (N_1287,In_15,In_1337);
and U1288 (N_1288,In_1922,In_1597);
nor U1289 (N_1289,In_2026,In_320);
nand U1290 (N_1290,In_2069,In_1060);
and U1291 (N_1291,In_1645,In_1223);
or U1292 (N_1292,In_754,In_1805);
and U1293 (N_1293,In_1222,In_352);
or U1294 (N_1294,In_73,In_343);
or U1295 (N_1295,In_2007,In_1291);
or U1296 (N_1296,In_949,In_266);
and U1297 (N_1297,In_526,In_567);
or U1298 (N_1298,In_1166,In_2437);
or U1299 (N_1299,In_586,In_643);
and U1300 (N_1300,In_1266,In_1372);
nand U1301 (N_1301,In_2100,In_2014);
and U1302 (N_1302,In_1161,In_1324);
or U1303 (N_1303,In_2084,In_1585);
xnor U1304 (N_1304,In_1421,In_112);
nand U1305 (N_1305,In_1140,In_8);
xnor U1306 (N_1306,In_77,In_1688);
nor U1307 (N_1307,In_188,In_2089);
nor U1308 (N_1308,In_2285,In_700);
nor U1309 (N_1309,In_2039,In_296);
nand U1310 (N_1310,In_2447,In_628);
and U1311 (N_1311,In_1547,In_1153);
nand U1312 (N_1312,In_198,In_766);
nand U1313 (N_1313,In_2401,In_2033);
and U1314 (N_1314,In_1456,In_359);
and U1315 (N_1315,In_13,In_1191);
or U1316 (N_1316,In_1438,In_1642);
or U1317 (N_1317,In_1384,In_1514);
nand U1318 (N_1318,In_830,In_1101);
or U1319 (N_1319,In_217,In_2125);
nor U1320 (N_1320,In_2032,In_1870);
nor U1321 (N_1321,In_2414,In_150);
nand U1322 (N_1322,In_738,In_1379);
nand U1323 (N_1323,In_1175,In_1517);
xnor U1324 (N_1324,In_1405,In_37);
or U1325 (N_1325,In_1413,In_2389);
or U1326 (N_1326,In_2337,In_1733);
xor U1327 (N_1327,In_956,In_977);
nor U1328 (N_1328,In_974,In_2385);
nand U1329 (N_1329,In_195,In_816);
nand U1330 (N_1330,In_1042,In_619);
and U1331 (N_1331,In_1902,In_1103);
xor U1332 (N_1332,In_320,In_465);
nor U1333 (N_1333,In_2029,In_1721);
and U1334 (N_1334,In_2122,In_812);
nand U1335 (N_1335,In_1884,In_1415);
or U1336 (N_1336,In_303,In_826);
nand U1337 (N_1337,In_1179,In_2199);
and U1338 (N_1338,In_146,In_1753);
and U1339 (N_1339,In_2197,In_1128);
xor U1340 (N_1340,In_900,In_885);
xnor U1341 (N_1341,In_832,In_1413);
xnor U1342 (N_1342,In_550,In_536);
nand U1343 (N_1343,In_2343,In_14);
and U1344 (N_1344,In_2332,In_1556);
xor U1345 (N_1345,In_2329,In_2341);
or U1346 (N_1346,In_1779,In_714);
nor U1347 (N_1347,In_2118,In_2162);
nor U1348 (N_1348,In_2006,In_2300);
nor U1349 (N_1349,In_399,In_1188);
nand U1350 (N_1350,In_2276,In_1705);
and U1351 (N_1351,In_2189,In_272);
and U1352 (N_1352,In_844,In_2310);
and U1353 (N_1353,In_1211,In_45);
and U1354 (N_1354,In_1109,In_2435);
xor U1355 (N_1355,In_2376,In_1313);
nand U1356 (N_1356,In_2124,In_1135);
nand U1357 (N_1357,In_203,In_542);
nand U1358 (N_1358,In_2133,In_1772);
nand U1359 (N_1359,In_1377,In_803);
nand U1360 (N_1360,In_440,In_2330);
and U1361 (N_1361,In_1123,In_2338);
or U1362 (N_1362,In_28,In_2023);
nor U1363 (N_1363,In_2485,In_512);
xor U1364 (N_1364,In_976,In_230);
or U1365 (N_1365,In_1368,In_1632);
xor U1366 (N_1366,In_2375,In_785);
and U1367 (N_1367,In_1913,In_2042);
or U1368 (N_1368,In_1046,In_1619);
or U1369 (N_1369,In_1147,In_175);
and U1370 (N_1370,In_1744,In_20);
xor U1371 (N_1371,In_886,In_2238);
nand U1372 (N_1372,In_1776,In_1110);
or U1373 (N_1373,In_1849,In_2084);
xnor U1374 (N_1374,In_1782,In_2496);
nand U1375 (N_1375,In_2379,In_2023);
nand U1376 (N_1376,In_1781,In_2059);
or U1377 (N_1377,In_356,In_1614);
and U1378 (N_1378,In_779,In_1960);
nand U1379 (N_1379,In_2421,In_2492);
nor U1380 (N_1380,In_2486,In_630);
and U1381 (N_1381,In_1857,In_540);
and U1382 (N_1382,In_1206,In_1164);
nand U1383 (N_1383,In_1966,In_1608);
nand U1384 (N_1384,In_2436,In_961);
xor U1385 (N_1385,In_259,In_816);
nor U1386 (N_1386,In_870,In_1077);
nor U1387 (N_1387,In_2390,In_1199);
nand U1388 (N_1388,In_1791,In_1492);
and U1389 (N_1389,In_963,In_1888);
xor U1390 (N_1390,In_195,In_2358);
nor U1391 (N_1391,In_1884,In_856);
xor U1392 (N_1392,In_826,In_1801);
or U1393 (N_1393,In_906,In_2393);
or U1394 (N_1394,In_206,In_1148);
xor U1395 (N_1395,In_1111,In_1947);
or U1396 (N_1396,In_2134,In_622);
nor U1397 (N_1397,In_840,In_1369);
and U1398 (N_1398,In_1069,In_665);
and U1399 (N_1399,In_2409,In_19);
nor U1400 (N_1400,In_2424,In_2293);
nor U1401 (N_1401,In_199,In_129);
nor U1402 (N_1402,In_894,In_1039);
nor U1403 (N_1403,In_729,In_130);
nand U1404 (N_1404,In_570,In_1379);
or U1405 (N_1405,In_985,In_2248);
and U1406 (N_1406,In_1445,In_52);
nor U1407 (N_1407,In_1839,In_786);
nor U1408 (N_1408,In_482,In_1548);
or U1409 (N_1409,In_2498,In_1724);
xnor U1410 (N_1410,In_1542,In_573);
xnor U1411 (N_1411,In_139,In_1176);
or U1412 (N_1412,In_1275,In_1007);
nor U1413 (N_1413,In_2284,In_254);
or U1414 (N_1414,In_1949,In_1074);
or U1415 (N_1415,In_623,In_1461);
xor U1416 (N_1416,In_1479,In_2358);
or U1417 (N_1417,In_134,In_598);
xor U1418 (N_1418,In_512,In_1308);
nand U1419 (N_1419,In_1189,In_1709);
nand U1420 (N_1420,In_2011,In_332);
nor U1421 (N_1421,In_674,In_1861);
nand U1422 (N_1422,In_2281,In_2171);
or U1423 (N_1423,In_779,In_1348);
and U1424 (N_1424,In_822,In_631);
nor U1425 (N_1425,In_2451,In_607);
or U1426 (N_1426,In_916,In_1987);
nor U1427 (N_1427,In_844,In_478);
and U1428 (N_1428,In_1392,In_595);
or U1429 (N_1429,In_897,In_1149);
xnor U1430 (N_1430,In_111,In_230);
or U1431 (N_1431,In_970,In_1021);
and U1432 (N_1432,In_863,In_84);
or U1433 (N_1433,In_2433,In_1729);
and U1434 (N_1434,In_1091,In_664);
or U1435 (N_1435,In_1338,In_373);
nand U1436 (N_1436,In_1177,In_1337);
and U1437 (N_1437,In_1049,In_584);
nor U1438 (N_1438,In_1809,In_1795);
xor U1439 (N_1439,In_1430,In_2005);
or U1440 (N_1440,In_510,In_656);
xor U1441 (N_1441,In_1548,In_240);
nand U1442 (N_1442,In_1152,In_77);
and U1443 (N_1443,In_239,In_1468);
and U1444 (N_1444,In_1179,In_235);
xor U1445 (N_1445,In_1019,In_474);
nand U1446 (N_1446,In_20,In_13);
xnor U1447 (N_1447,In_1097,In_1851);
nor U1448 (N_1448,In_556,In_1528);
and U1449 (N_1449,In_520,In_903);
or U1450 (N_1450,In_849,In_671);
nand U1451 (N_1451,In_1315,In_1755);
nor U1452 (N_1452,In_2451,In_804);
and U1453 (N_1453,In_760,In_57);
nor U1454 (N_1454,In_1074,In_1480);
nand U1455 (N_1455,In_1218,In_2327);
nor U1456 (N_1456,In_2041,In_729);
nand U1457 (N_1457,In_1844,In_617);
or U1458 (N_1458,In_1034,In_1363);
xnor U1459 (N_1459,In_577,In_970);
nor U1460 (N_1460,In_1477,In_2458);
and U1461 (N_1461,In_1569,In_1296);
and U1462 (N_1462,In_2028,In_727);
and U1463 (N_1463,In_712,In_106);
xor U1464 (N_1464,In_68,In_1025);
and U1465 (N_1465,In_1056,In_467);
and U1466 (N_1466,In_2084,In_2012);
or U1467 (N_1467,In_2108,In_2338);
xnor U1468 (N_1468,In_708,In_1806);
and U1469 (N_1469,In_43,In_1378);
nor U1470 (N_1470,In_734,In_1530);
nor U1471 (N_1471,In_914,In_1630);
nor U1472 (N_1472,In_1000,In_2486);
xnor U1473 (N_1473,In_586,In_1769);
xnor U1474 (N_1474,In_661,In_379);
nand U1475 (N_1475,In_638,In_1726);
and U1476 (N_1476,In_1408,In_78);
xnor U1477 (N_1477,In_2106,In_135);
xnor U1478 (N_1478,In_2182,In_799);
nor U1479 (N_1479,In_329,In_782);
nand U1480 (N_1480,In_473,In_1682);
or U1481 (N_1481,In_552,In_103);
nand U1482 (N_1482,In_1894,In_1922);
nand U1483 (N_1483,In_729,In_2223);
xnor U1484 (N_1484,In_1744,In_1428);
nor U1485 (N_1485,In_2026,In_2204);
and U1486 (N_1486,In_1927,In_1444);
xnor U1487 (N_1487,In_2326,In_1546);
and U1488 (N_1488,In_1590,In_1317);
or U1489 (N_1489,In_1166,In_2079);
and U1490 (N_1490,In_2139,In_207);
and U1491 (N_1491,In_1440,In_884);
or U1492 (N_1492,In_2364,In_1860);
xnor U1493 (N_1493,In_242,In_1272);
and U1494 (N_1494,In_1523,In_1762);
or U1495 (N_1495,In_2492,In_134);
nand U1496 (N_1496,In_2033,In_472);
nand U1497 (N_1497,In_1360,In_1442);
nor U1498 (N_1498,In_677,In_966);
nor U1499 (N_1499,In_491,In_138);
xor U1500 (N_1500,In_138,In_175);
nor U1501 (N_1501,In_28,In_855);
and U1502 (N_1502,In_1649,In_1177);
and U1503 (N_1503,In_1627,In_1636);
xor U1504 (N_1504,In_1199,In_1315);
xor U1505 (N_1505,In_1611,In_1381);
or U1506 (N_1506,In_1644,In_1215);
nor U1507 (N_1507,In_715,In_1880);
or U1508 (N_1508,In_1668,In_465);
nor U1509 (N_1509,In_318,In_298);
nor U1510 (N_1510,In_1184,In_896);
nor U1511 (N_1511,In_864,In_673);
and U1512 (N_1512,In_553,In_1435);
nand U1513 (N_1513,In_2171,In_1765);
nor U1514 (N_1514,In_1183,In_428);
or U1515 (N_1515,In_2270,In_2184);
and U1516 (N_1516,In_1579,In_539);
or U1517 (N_1517,In_139,In_879);
nand U1518 (N_1518,In_1509,In_1446);
nand U1519 (N_1519,In_356,In_1676);
nor U1520 (N_1520,In_2307,In_1849);
nor U1521 (N_1521,In_1325,In_1802);
and U1522 (N_1522,In_983,In_1868);
xor U1523 (N_1523,In_696,In_839);
or U1524 (N_1524,In_701,In_1655);
xnor U1525 (N_1525,In_1922,In_1039);
nor U1526 (N_1526,In_512,In_2063);
and U1527 (N_1527,In_237,In_1055);
or U1528 (N_1528,In_1675,In_2486);
nor U1529 (N_1529,In_2492,In_83);
xnor U1530 (N_1530,In_381,In_121);
xor U1531 (N_1531,In_379,In_976);
xnor U1532 (N_1532,In_2260,In_2419);
nand U1533 (N_1533,In_2094,In_2085);
nand U1534 (N_1534,In_378,In_491);
nand U1535 (N_1535,In_2201,In_2096);
nor U1536 (N_1536,In_1327,In_2152);
xnor U1537 (N_1537,In_1684,In_1031);
or U1538 (N_1538,In_192,In_1026);
nor U1539 (N_1539,In_820,In_241);
xnor U1540 (N_1540,In_1137,In_1812);
and U1541 (N_1541,In_1758,In_1733);
nor U1542 (N_1542,In_611,In_296);
nor U1543 (N_1543,In_1392,In_81);
nor U1544 (N_1544,In_2005,In_203);
xor U1545 (N_1545,In_1261,In_1913);
nand U1546 (N_1546,In_2259,In_2367);
nand U1547 (N_1547,In_96,In_1216);
or U1548 (N_1548,In_237,In_844);
and U1549 (N_1549,In_279,In_1623);
or U1550 (N_1550,In_331,In_1248);
or U1551 (N_1551,In_40,In_66);
or U1552 (N_1552,In_2034,In_1482);
or U1553 (N_1553,In_1747,In_1476);
xor U1554 (N_1554,In_2213,In_1927);
xnor U1555 (N_1555,In_1352,In_761);
or U1556 (N_1556,In_1781,In_1111);
nor U1557 (N_1557,In_2059,In_292);
and U1558 (N_1558,In_139,In_993);
or U1559 (N_1559,In_2375,In_1628);
nand U1560 (N_1560,In_1838,In_152);
and U1561 (N_1561,In_1410,In_1891);
nand U1562 (N_1562,In_1176,In_773);
nor U1563 (N_1563,In_1393,In_1896);
or U1564 (N_1564,In_216,In_1941);
and U1565 (N_1565,In_232,In_887);
and U1566 (N_1566,In_1977,In_437);
and U1567 (N_1567,In_1678,In_1166);
or U1568 (N_1568,In_1634,In_1930);
xnor U1569 (N_1569,In_1353,In_2115);
and U1570 (N_1570,In_425,In_990);
nor U1571 (N_1571,In_1097,In_1744);
and U1572 (N_1572,In_1487,In_393);
and U1573 (N_1573,In_1368,In_895);
nor U1574 (N_1574,In_2012,In_1646);
xnor U1575 (N_1575,In_130,In_1241);
or U1576 (N_1576,In_874,In_130);
nor U1577 (N_1577,In_1965,In_1835);
xor U1578 (N_1578,In_104,In_373);
or U1579 (N_1579,In_1285,In_1364);
nor U1580 (N_1580,In_2473,In_1066);
nor U1581 (N_1581,In_1744,In_2145);
nor U1582 (N_1582,In_212,In_2325);
and U1583 (N_1583,In_392,In_2117);
nand U1584 (N_1584,In_366,In_1521);
or U1585 (N_1585,In_132,In_869);
and U1586 (N_1586,In_2441,In_723);
and U1587 (N_1587,In_1611,In_1153);
nor U1588 (N_1588,In_935,In_1939);
and U1589 (N_1589,In_1804,In_404);
xor U1590 (N_1590,In_1218,In_750);
or U1591 (N_1591,In_786,In_757);
and U1592 (N_1592,In_2179,In_1731);
or U1593 (N_1593,In_2383,In_334);
and U1594 (N_1594,In_1239,In_1203);
xnor U1595 (N_1595,In_2018,In_1992);
or U1596 (N_1596,In_1127,In_1575);
nand U1597 (N_1597,In_374,In_1317);
xor U1598 (N_1598,In_2435,In_2445);
or U1599 (N_1599,In_100,In_362);
or U1600 (N_1600,In_70,In_799);
or U1601 (N_1601,In_2114,In_1810);
or U1602 (N_1602,In_1650,In_1557);
and U1603 (N_1603,In_1987,In_1089);
nand U1604 (N_1604,In_1531,In_1381);
nand U1605 (N_1605,In_1310,In_1222);
nor U1606 (N_1606,In_1429,In_1755);
nand U1607 (N_1607,In_1,In_1617);
or U1608 (N_1608,In_1835,In_264);
or U1609 (N_1609,In_1833,In_2330);
or U1610 (N_1610,In_2368,In_660);
and U1611 (N_1611,In_128,In_2329);
and U1612 (N_1612,In_548,In_2314);
or U1613 (N_1613,In_61,In_1747);
nand U1614 (N_1614,In_457,In_1153);
nand U1615 (N_1615,In_1836,In_473);
nor U1616 (N_1616,In_2288,In_1765);
nand U1617 (N_1617,In_72,In_2394);
and U1618 (N_1618,In_1605,In_1458);
or U1619 (N_1619,In_400,In_1002);
or U1620 (N_1620,In_554,In_2191);
or U1621 (N_1621,In_729,In_775);
and U1622 (N_1622,In_385,In_1347);
and U1623 (N_1623,In_493,In_2251);
or U1624 (N_1624,In_2265,In_966);
or U1625 (N_1625,In_400,In_675);
or U1626 (N_1626,In_834,In_2109);
nor U1627 (N_1627,In_1808,In_717);
and U1628 (N_1628,In_2403,In_593);
and U1629 (N_1629,In_311,In_1750);
nand U1630 (N_1630,In_1527,In_385);
nor U1631 (N_1631,In_871,In_838);
or U1632 (N_1632,In_2394,In_0);
and U1633 (N_1633,In_2203,In_1974);
xnor U1634 (N_1634,In_681,In_1892);
or U1635 (N_1635,In_2107,In_955);
or U1636 (N_1636,In_1021,In_2010);
nand U1637 (N_1637,In_347,In_2411);
or U1638 (N_1638,In_1298,In_1743);
or U1639 (N_1639,In_1853,In_380);
nand U1640 (N_1640,In_1494,In_1698);
or U1641 (N_1641,In_1505,In_238);
nand U1642 (N_1642,In_1729,In_2000);
xnor U1643 (N_1643,In_1233,In_2299);
nor U1644 (N_1644,In_1902,In_1329);
and U1645 (N_1645,In_821,In_992);
or U1646 (N_1646,In_1831,In_1697);
and U1647 (N_1647,In_2481,In_1056);
or U1648 (N_1648,In_989,In_705);
nor U1649 (N_1649,In_2006,In_1593);
xor U1650 (N_1650,In_947,In_146);
xor U1651 (N_1651,In_1303,In_533);
and U1652 (N_1652,In_646,In_116);
or U1653 (N_1653,In_199,In_111);
xnor U1654 (N_1654,In_2288,In_442);
nand U1655 (N_1655,In_52,In_1186);
and U1656 (N_1656,In_1039,In_63);
xnor U1657 (N_1657,In_1682,In_1599);
nor U1658 (N_1658,In_1285,In_662);
and U1659 (N_1659,In_1801,In_1510);
nand U1660 (N_1660,In_932,In_1126);
and U1661 (N_1661,In_387,In_1960);
nand U1662 (N_1662,In_1997,In_2204);
or U1663 (N_1663,In_1497,In_471);
xnor U1664 (N_1664,In_817,In_39);
and U1665 (N_1665,In_1216,In_2221);
and U1666 (N_1666,In_795,In_1887);
nor U1667 (N_1667,In_305,In_519);
and U1668 (N_1668,In_134,In_1479);
or U1669 (N_1669,In_505,In_437);
or U1670 (N_1670,In_2429,In_1852);
nand U1671 (N_1671,In_133,In_317);
or U1672 (N_1672,In_723,In_970);
nor U1673 (N_1673,In_1653,In_2282);
xnor U1674 (N_1674,In_367,In_994);
and U1675 (N_1675,In_1041,In_1197);
xor U1676 (N_1676,In_569,In_626);
nor U1677 (N_1677,In_2037,In_299);
and U1678 (N_1678,In_1135,In_1350);
nand U1679 (N_1679,In_298,In_1784);
nor U1680 (N_1680,In_129,In_1083);
xnor U1681 (N_1681,In_147,In_663);
nor U1682 (N_1682,In_1193,In_1662);
xor U1683 (N_1683,In_298,In_2485);
or U1684 (N_1684,In_2082,In_2210);
or U1685 (N_1685,In_559,In_242);
nor U1686 (N_1686,In_734,In_300);
nand U1687 (N_1687,In_133,In_252);
and U1688 (N_1688,In_1252,In_995);
and U1689 (N_1689,In_1654,In_2461);
xor U1690 (N_1690,In_1825,In_1714);
and U1691 (N_1691,In_285,In_2022);
nand U1692 (N_1692,In_382,In_1427);
or U1693 (N_1693,In_1497,In_568);
or U1694 (N_1694,In_841,In_1383);
nor U1695 (N_1695,In_1037,In_692);
and U1696 (N_1696,In_1077,In_1574);
and U1697 (N_1697,In_677,In_661);
nand U1698 (N_1698,In_1374,In_2120);
nor U1699 (N_1699,In_2168,In_2017);
xor U1700 (N_1700,In_392,In_134);
or U1701 (N_1701,In_2148,In_696);
nand U1702 (N_1702,In_480,In_1384);
nand U1703 (N_1703,In_76,In_623);
nor U1704 (N_1704,In_2011,In_1503);
nand U1705 (N_1705,In_69,In_868);
nand U1706 (N_1706,In_1278,In_1617);
and U1707 (N_1707,In_1191,In_1028);
or U1708 (N_1708,In_1935,In_1704);
xor U1709 (N_1709,In_2402,In_2165);
nand U1710 (N_1710,In_1133,In_1168);
xnor U1711 (N_1711,In_2054,In_1334);
and U1712 (N_1712,In_1578,In_173);
nor U1713 (N_1713,In_850,In_1803);
nor U1714 (N_1714,In_1399,In_1449);
or U1715 (N_1715,In_1649,In_379);
or U1716 (N_1716,In_482,In_2497);
nor U1717 (N_1717,In_563,In_1592);
and U1718 (N_1718,In_419,In_2194);
nand U1719 (N_1719,In_368,In_579);
nand U1720 (N_1720,In_750,In_453);
nand U1721 (N_1721,In_957,In_1422);
and U1722 (N_1722,In_1958,In_301);
or U1723 (N_1723,In_2458,In_1929);
xnor U1724 (N_1724,In_1728,In_275);
and U1725 (N_1725,In_390,In_1162);
nand U1726 (N_1726,In_1392,In_901);
nor U1727 (N_1727,In_402,In_2183);
or U1728 (N_1728,In_560,In_1210);
nand U1729 (N_1729,In_269,In_39);
xnor U1730 (N_1730,In_786,In_589);
nand U1731 (N_1731,In_243,In_900);
nor U1732 (N_1732,In_163,In_1859);
nand U1733 (N_1733,In_2313,In_667);
nor U1734 (N_1734,In_391,In_776);
or U1735 (N_1735,In_2027,In_395);
xnor U1736 (N_1736,In_1241,In_226);
or U1737 (N_1737,In_567,In_1985);
xor U1738 (N_1738,In_1601,In_2008);
or U1739 (N_1739,In_1426,In_2189);
and U1740 (N_1740,In_133,In_388);
nand U1741 (N_1741,In_122,In_1617);
or U1742 (N_1742,In_1425,In_2229);
or U1743 (N_1743,In_2134,In_2090);
nor U1744 (N_1744,In_1152,In_190);
nor U1745 (N_1745,In_2084,In_1851);
xor U1746 (N_1746,In_1823,In_2281);
xor U1747 (N_1747,In_1448,In_703);
nand U1748 (N_1748,In_764,In_280);
or U1749 (N_1749,In_1540,In_1188);
and U1750 (N_1750,In_1269,In_1953);
xor U1751 (N_1751,In_1825,In_1380);
nor U1752 (N_1752,In_275,In_50);
nor U1753 (N_1753,In_488,In_981);
nor U1754 (N_1754,In_438,In_31);
and U1755 (N_1755,In_1205,In_2186);
nor U1756 (N_1756,In_1235,In_2145);
or U1757 (N_1757,In_1284,In_1373);
nor U1758 (N_1758,In_2103,In_2027);
xor U1759 (N_1759,In_534,In_2439);
xnor U1760 (N_1760,In_475,In_2198);
or U1761 (N_1761,In_1881,In_2032);
or U1762 (N_1762,In_1817,In_1830);
xor U1763 (N_1763,In_2424,In_1899);
xor U1764 (N_1764,In_1253,In_508);
and U1765 (N_1765,In_1355,In_1694);
nand U1766 (N_1766,In_859,In_2113);
and U1767 (N_1767,In_2226,In_1460);
nor U1768 (N_1768,In_1770,In_1347);
and U1769 (N_1769,In_292,In_77);
and U1770 (N_1770,In_896,In_766);
nand U1771 (N_1771,In_2406,In_240);
nand U1772 (N_1772,In_664,In_1315);
nor U1773 (N_1773,In_512,In_1840);
and U1774 (N_1774,In_1339,In_1205);
or U1775 (N_1775,In_1843,In_1181);
nand U1776 (N_1776,In_778,In_109);
nand U1777 (N_1777,In_1120,In_706);
xor U1778 (N_1778,In_2292,In_1416);
xor U1779 (N_1779,In_2392,In_969);
nor U1780 (N_1780,In_2313,In_984);
xor U1781 (N_1781,In_2069,In_1455);
or U1782 (N_1782,In_33,In_1237);
and U1783 (N_1783,In_1344,In_1809);
xor U1784 (N_1784,In_2431,In_1893);
nor U1785 (N_1785,In_595,In_1550);
xnor U1786 (N_1786,In_72,In_2169);
and U1787 (N_1787,In_2443,In_325);
and U1788 (N_1788,In_2496,In_2019);
and U1789 (N_1789,In_221,In_2415);
nor U1790 (N_1790,In_303,In_946);
or U1791 (N_1791,In_2024,In_1547);
nor U1792 (N_1792,In_1755,In_2344);
or U1793 (N_1793,In_847,In_397);
or U1794 (N_1794,In_2374,In_1495);
xor U1795 (N_1795,In_1248,In_1855);
xnor U1796 (N_1796,In_2337,In_1955);
nand U1797 (N_1797,In_1674,In_1164);
and U1798 (N_1798,In_956,In_1356);
nor U1799 (N_1799,In_135,In_1287);
or U1800 (N_1800,In_477,In_2243);
nand U1801 (N_1801,In_85,In_1476);
nor U1802 (N_1802,In_2233,In_2467);
or U1803 (N_1803,In_360,In_1463);
nand U1804 (N_1804,In_1986,In_462);
nand U1805 (N_1805,In_2096,In_2103);
or U1806 (N_1806,In_2018,In_1506);
nor U1807 (N_1807,In_2479,In_1931);
and U1808 (N_1808,In_2311,In_160);
and U1809 (N_1809,In_2060,In_63);
nand U1810 (N_1810,In_836,In_2282);
nor U1811 (N_1811,In_890,In_46);
nand U1812 (N_1812,In_646,In_323);
nand U1813 (N_1813,In_1306,In_750);
nand U1814 (N_1814,In_1829,In_1608);
xnor U1815 (N_1815,In_544,In_1538);
nor U1816 (N_1816,In_260,In_85);
and U1817 (N_1817,In_2377,In_424);
nand U1818 (N_1818,In_1914,In_1746);
xor U1819 (N_1819,In_97,In_1025);
nand U1820 (N_1820,In_55,In_2226);
or U1821 (N_1821,In_2227,In_1677);
or U1822 (N_1822,In_1307,In_1746);
or U1823 (N_1823,In_1922,In_2096);
or U1824 (N_1824,In_1836,In_2178);
nor U1825 (N_1825,In_2042,In_291);
xnor U1826 (N_1826,In_2076,In_1433);
nand U1827 (N_1827,In_1261,In_124);
or U1828 (N_1828,In_1579,In_1486);
and U1829 (N_1829,In_1673,In_925);
and U1830 (N_1830,In_744,In_2149);
and U1831 (N_1831,In_307,In_1463);
nand U1832 (N_1832,In_2392,In_181);
nand U1833 (N_1833,In_1175,In_1305);
nor U1834 (N_1834,In_548,In_1825);
or U1835 (N_1835,In_449,In_1956);
or U1836 (N_1836,In_1998,In_234);
or U1837 (N_1837,In_555,In_127);
xnor U1838 (N_1838,In_1915,In_435);
nand U1839 (N_1839,In_156,In_599);
xnor U1840 (N_1840,In_202,In_1464);
or U1841 (N_1841,In_2043,In_581);
nand U1842 (N_1842,In_1555,In_2391);
and U1843 (N_1843,In_1373,In_1547);
nand U1844 (N_1844,In_1586,In_1673);
nor U1845 (N_1845,In_213,In_2118);
and U1846 (N_1846,In_1865,In_1629);
nor U1847 (N_1847,In_670,In_2223);
xor U1848 (N_1848,In_221,In_118);
or U1849 (N_1849,In_1251,In_1076);
nor U1850 (N_1850,In_646,In_1697);
and U1851 (N_1851,In_310,In_2391);
or U1852 (N_1852,In_1298,In_1379);
nor U1853 (N_1853,In_1137,In_262);
nor U1854 (N_1854,In_1213,In_1283);
and U1855 (N_1855,In_1282,In_2342);
or U1856 (N_1856,In_1964,In_824);
nand U1857 (N_1857,In_2458,In_2342);
nor U1858 (N_1858,In_506,In_193);
or U1859 (N_1859,In_317,In_594);
xnor U1860 (N_1860,In_100,In_823);
or U1861 (N_1861,In_2204,In_758);
nor U1862 (N_1862,In_2053,In_302);
nand U1863 (N_1863,In_858,In_1861);
or U1864 (N_1864,In_1546,In_1380);
and U1865 (N_1865,In_333,In_1587);
xor U1866 (N_1866,In_1251,In_1020);
and U1867 (N_1867,In_500,In_56);
nand U1868 (N_1868,In_169,In_156);
or U1869 (N_1869,In_1379,In_2076);
xnor U1870 (N_1870,In_976,In_176);
or U1871 (N_1871,In_426,In_772);
and U1872 (N_1872,In_2350,In_2111);
nor U1873 (N_1873,In_1006,In_1740);
or U1874 (N_1874,In_227,In_924);
or U1875 (N_1875,In_751,In_1499);
or U1876 (N_1876,In_1078,In_1936);
and U1877 (N_1877,In_692,In_1385);
and U1878 (N_1878,In_270,In_1682);
or U1879 (N_1879,In_170,In_1583);
nand U1880 (N_1880,In_1450,In_1025);
nand U1881 (N_1881,In_102,In_790);
and U1882 (N_1882,In_2265,In_2497);
or U1883 (N_1883,In_1245,In_1379);
and U1884 (N_1884,In_360,In_1184);
or U1885 (N_1885,In_2264,In_1162);
nand U1886 (N_1886,In_875,In_730);
nand U1887 (N_1887,In_1856,In_2402);
or U1888 (N_1888,In_2364,In_1810);
and U1889 (N_1889,In_1524,In_212);
xnor U1890 (N_1890,In_1155,In_1719);
or U1891 (N_1891,In_1132,In_1297);
or U1892 (N_1892,In_2385,In_1162);
nand U1893 (N_1893,In_115,In_795);
nor U1894 (N_1894,In_375,In_1722);
nand U1895 (N_1895,In_936,In_2133);
nand U1896 (N_1896,In_2419,In_949);
nor U1897 (N_1897,In_1352,In_748);
nor U1898 (N_1898,In_2072,In_2461);
nand U1899 (N_1899,In_53,In_151);
xnor U1900 (N_1900,In_71,In_473);
nand U1901 (N_1901,In_1752,In_252);
xor U1902 (N_1902,In_2472,In_2338);
or U1903 (N_1903,In_2135,In_2152);
or U1904 (N_1904,In_523,In_1822);
xnor U1905 (N_1905,In_186,In_2146);
and U1906 (N_1906,In_2246,In_716);
nor U1907 (N_1907,In_1472,In_113);
xnor U1908 (N_1908,In_2102,In_1360);
nor U1909 (N_1909,In_1657,In_2110);
xor U1910 (N_1910,In_811,In_400);
nor U1911 (N_1911,In_2412,In_1852);
xor U1912 (N_1912,In_274,In_2206);
or U1913 (N_1913,In_2055,In_289);
or U1914 (N_1914,In_189,In_2424);
nand U1915 (N_1915,In_1959,In_1134);
xor U1916 (N_1916,In_137,In_298);
nand U1917 (N_1917,In_1193,In_1943);
nor U1918 (N_1918,In_1288,In_1786);
or U1919 (N_1919,In_1761,In_2233);
and U1920 (N_1920,In_2336,In_1038);
xor U1921 (N_1921,In_1289,In_1368);
nand U1922 (N_1922,In_2009,In_2106);
and U1923 (N_1923,In_1212,In_1997);
nand U1924 (N_1924,In_40,In_1387);
and U1925 (N_1925,In_2267,In_1118);
nand U1926 (N_1926,In_1785,In_658);
or U1927 (N_1927,In_692,In_2339);
or U1928 (N_1928,In_1495,In_2220);
and U1929 (N_1929,In_619,In_2351);
nor U1930 (N_1930,In_240,In_2);
or U1931 (N_1931,In_186,In_1684);
nand U1932 (N_1932,In_2164,In_1505);
or U1933 (N_1933,In_550,In_1966);
and U1934 (N_1934,In_1988,In_2391);
nor U1935 (N_1935,In_1356,In_336);
or U1936 (N_1936,In_2260,In_1702);
nor U1937 (N_1937,In_1467,In_2423);
nor U1938 (N_1938,In_120,In_234);
or U1939 (N_1939,In_1891,In_1914);
nor U1940 (N_1940,In_1839,In_1740);
and U1941 (N_1941,In_248,In_875);
and U1942 (N_1942,In_809,In_1148);
nand U1943 (N_1943,In_1292,In_1488);
or U1944 (N_1944,In_705,In_92);
xor U1945 (N_1945,In_2176,In_828);
and U1946 (N_1946,In_1181,In_2151);
nand U1947 (N_1947,In_2324,In_630);
xor U1948 (N_1948,In_211,In_734);
or U1949 (N_1949,In_2001,In_2400);
or U1950 (N_1950,In_1882,In_2308);
and U1951 (N_1951,In_368,In_2379);
xor U1952 (N_1952,In_628,In_1359);
nand U1953 (N_1953,In_1081,In_1747);
nor U1954 (N_1954,In_2071,In_2086);
and U1955 (N_1955,In_105,In_1123);
or U1956 (N_1956,In_122,In_1394);
or U1957 (N_1957,In_380,In_1897);
and U1958 (N_1958,In_31,In_1306);
nor U1959 (N_1959,In_1380,In_338);
nand U1960 (N_1960,In_382,In_320);
xnor U1961 (N_1961,In_1648,In_813);
nor U1962 (N_1962,In_546,In_2214);
or U1963 (N_1963,In_412,In_2106);
nand U1964 (N_1964,In_485,In_1036);
or U1965 (N_1965,In_2172,In_2446);
or U1966 (N_1966,In_2478,In_74);
nor U1967 (N_1967,In_1853,In_596);
nand U1968 (N_1968,In_2000,In_2080);
nand U1969 (N_1969,In_1389,In_1691);
nor U1970 (N_1970,In_2209,In_1105);
and U1971 (N_1971,In_1436,In_505);
nand U1972 (N_1972,In_1372,In_1343);
and U1973 (N_1973,In_2358,In_1580);
and U1974 (N_1974,In_626,In_1898);
and U1975 (N_1975,In_1453,In_2195);
nand U1976 (N_1976,In_1786,In_2031);
or U1977 (N_1977,In_1381,In_36);
or U1978 (N_1978,In_616,In_2411);
and U1979 (N_1979,In_563,In_1485);
or U1980 (N_1980,In_40,In_888);
or U1981 (N_1981,In_1431,In_1947);
nand U1982 (N_1982,In_2243,In_849);
nand U1983 (N_1983,In_491,In_1787);
nand U1984 (N_1984,In_1043,In_1657);
and U1985 (N_1985,In_278,In_1498);
or U1986 (N_1986,In_1129,In_1052);
and U1987 (N_1987,In_66,In_1745);
nor U1988 (N_1988,In_2290,In_1818);
nand U1989 (N_1989,In_1622,In_802);
nor U1990 (N_1990,In_1088,In_1770);
and U1991 (N_1991,In_2349,In_457);
nand U1992 (N_1992,In_383,In_2387);
xor U1993 (N_1993,In_2075,In_2337);
or U1994 (N_1994,In_1567,In_2130);
or U1995 (N_1995,In_1148,In_507);
xnor U1996 (N_1996,In_1811,In_348);
nand U1997 (N_1997,In_2306,In_719);
nand U1998 (N_1998,In_1730,In_1843);
and U1999 (N_1999,In_1725,In_1403);
or U2000 (N_2000,In_621,In_2169);
and U2001 (N_2001,In_685,In_193);
and U2002 (N_2002,In_315,In_592);
and U2003 (N_2003,In_1593,In_568);
nand U2004 (N_2004,In_1490,In_431);
or U2005 (N_2005,In_2249,In_981);
and U2006 (N_2006,In_605,In_2114);
or U2007 (N_2007,In_2115,In_1958);
or U2008 (N_2008,In_2278,In_1530);
or U2009 (N_2009,In_1228,In_1934);
nor U2010 (N_2010,In_1998,In_509);
nor U2011 (N_2011,In_1936,In_2151);
xnor U2012 (N_2012,In_1281,In_240);
or U2013 (N_2013,In_1091,In_2235);
or U2014 (N_2014,In_31,In_1935);
and U2015 (N_2015,In_448,In_1921);
xnor U2016 (N_2016,In_919,In_1585);
xnor U2017 (N_2017,In_1357,In_2461);
and U2018 (N_2018,In_2248,In_715);
or U2019 (N_2019,In_386,In_1706);
and U2020 (N_2020,In_1541,In_1327);
or U2021 (N_2021,In_1884,In_1671);
xor U2022 (N_2022,In_1518,In_1402);
or U2023 (N_2023,In_2043,In_1866);
or U2024 (N_2024,In_2484,In_399);
xnor U2025 (N_2025,In_649,In_1900);
or U2026 (N_2026,In_1939,In_477);
nor U2027 (N_2027,In_573,In_1456);
xor U2028 (N_2028,In_1592,In_544);
nand U2029 (N_2029,In_658,In_366);
nand U2030 (N_2030,In_1871,In_1417);
nor U2031 (N_2031,In_42,In_1666);
nor U2032 (N_2032,In_626,In_136);
or U2033 (N_2033,In_2400,In_381);
nand U2034 (N_2034,In_1823,In_248);
xor U2035 (N_2035,In_1893,In_223);
xor U2036 (N_2036,In_1674,In_1396);
xnor U2037 (N_2037,In_92,In_2075);
nor U2038 (N_2038,In_946,In_630);
xor U2039 (N_2039,In_618,In_1227);
or U2040 (N_2040,In_733,In_0);
nor U2041 (N_2041,In_1904,In_1000);
xnor U2042 (N_2042,In_1821,In_1557);
nand U2043 (N_2043,In_90,In_2246);
or U2044 (N_2044,In_255,In_1095);
nor U2045 (N_2045,In_1890,In_2279);
xor U2046 (N_2046,In_777,In_121);
nor U2047 (N_2047,In_1922,In_291);
nand U2048 (N_2048,In_2423,In_464);
nand U2049 (N_2049,In_1509,In_120);
nor U2050 (N_2050,In_1709,In_1289);
xnor U2051 (N_2051,In_1972,In_214);
or U2052 (N_2052,In_1161,In_1848);
nor U2053 (N_2053,In_1995,In_2012);
and U2054 (N_2054,In_1952,In_514);
nor U2055 (N_2055,In_1907,In_1640);
xor U2056 (N_2056,In_966,In_2277);
nand U2057 (N_2057,In_568,In_576);
nand U2058 (N_2058,In_1478,In_452);
or U2059 (N_2059,In_2357,In_560);
and U2060 (N_2060,In_947,In_945);
nor U2061 (N_2061,In_229,In_1846);
nand U2062 (N_2062,In_611,In_364);
or U2063 (N_2063,In_245,In_612);
nand U2064 (N_2064,In_368,In_2302);
or U2065 (N_2065,In_982,In_214);
and U2066 (N_2066,In_1218,In_371);
nand U2067 (N_2067,In_988,In_1569);
nor U2068 (N_2068,In_2436,In_1461);
xnor U2069 (N_2069,In_872,In_1965);
or U2070 (N_2070,In_1503,In_2405);
nand U2071 (N_2071,In_154,In_723);
and U2072 (N_2072,In_1307,In_2356);
nor U2073 (N_2073,In_1551,In_1459);
xor U2074 (N_2074,In_2182,In_1106);
nor U2075 (N_2075,In_1483,In_236);
xnor U2076 (N_2076,In_2245,In_627);
xnor U2077 (N_2077,In_197,In_1002);
and U2078 (N_2078,In_428,In_2057);
nor U2079 (N_2079,In_809,In_96);
nor U2080 (N_2080,In_845,In_98);
or U2081 (N_2081,In_376,In_631);
xor U2082 (N_2082,In_93,In_689);
or U2083 (N_2083,In_1893,In_735);
nand U2084 (N_2084,In_2299,In_854);
and U2085 (N_2085,In_2051,In_811);
nor U2086 (N_2086,In_2198,In_2147);
nand U2087 (N_2087,In_1708,In_1859);
or U2088 (N_2088,In_3,In_1764);
nor U2089 (N_2089,In_1554,In_1743);
or U2090 (N_2090,In_535,In_2393);
and U2091 (N_2091,In_1622,In_182);
or U2092 (N_2092,In_1975,In_814);
nand U2093 (N_2093,In_941,In_2436);
nand U2094 (N_2094,In_1094,In_1163);
nand U2095 (N_2095,In_415,In_668);
or U2096 (N_2096,In_1501,In_1316);
and U2097 (N_2097,In_47,In_1556);
nand U2098 (N_2098,In_2418,In_1521);
nor U2099 (N_2099,In_954,In_440);
and U2100 (N_2100,In_882,In_1143);
nor U2101 (N_2101,In_300,In_117);
or U2102 (N_2102,In_1764,In_2170);
or U2103 (N_2103,In_2018,In_1971);
and U2104 (N_2104,In_2073,In_1840);
or U2105 (N_2105,In_521,In_2130);
nand U2106 (N_2106,In_2429,In_1692);
xnor U2107 (N_2107,In_680,In_2012);
nand U2108 (N_2108,In_1446,In_2166);
nand U2109 (N_2109,In_1647,In_547);
xor U2110 (N_2110,In_56,In_928);
xnor U2111 (N_2111,In_2394,In_1168);
xor U2112 (N_2112,In_471,In_2397);
xnor U2113 (N_2113,In_840,In_965);
xnor U2114 (N_2114,In_1383,In_767);
and U2115 (N_2115,In_2228,In_691);
nor U2116 (N_2116,In_2087,In_1314);
nor U2117 (N_2117,In_1013,In_1502);
or U2118 (N_2118,In_2212,In_2492);
or U2119 (N_2119,In_815,In_1785);
or U2120 (N_2120,In_247,In_86);
xnor U2121 (N_2121,In_1479,In_1473);
xnor U2122 (N_2122,In_1340,In_1899);
nand U2123 (N_2123,In_1087,In_427);
or U2124 (N_2124,In_1514,In_2352);
nor U2125 (N_2125,In_1407,In_919);
xnor U2126 (N_2126,In_292,In_609);
nand U2127 (N_2127,In_1981,In_1071);
nand U2128 (N_2128,In_1308,In_330);
nor U2129 (N_2129,In_455,In_2038);
xnor U2130 (N_2130,In_1208,In_2425);
xor U2131 (N_2131,In_538,In_971);
nand U2132 (N_2132,In_2153,In_680);
and U2133 (N_2133,In_851,In_1185);
nand U2134 (N_2134,In_1565,In_1131);
nor U2135 (N_2135,In_2285,In_1625);
xor U2136 (N_2136,In_868,In_2071);
nand U2137 (N_2137,In_80,In_2150);
nand U2138 (N_2138,In_186,In_529);
nand U2139 (N_2139,In_721,In_275);
and U2140 (N_2140,In_2184,In_836);
nand U2141 (N_2141,In_1834,In_125);
or U2142 (N_2142,In_2438,In_1473);
nor U2143 (N_2143,In_1978,In_1410);
xnor U2144 (N_2144,In_2209,In_902);
and U2145 (N_2145,In_1200,In_526);
and U2146 (N_2146,In_288,In_303);
and U2147 (N_2147,In_2322,In_588);
nor U2148 (N_2148,In_2092,In_1427);
or U2149 (N_2149,In_1109,In_440);
nor U2150 (N_2150,In_2245,In_362);
xor U2151 (N_2151,In_252,In_89);
nor U2152 (N_2152,In_1567,In_1603);
and U2153 (N_2153,In_119,In_1806);
or U2154 (N_2154,In_537,In_1827);
nor U2155 (N_2155,In_1116,In_155);
and U2156 (N_2156,In_103,In_2484);
nor U2157 (N_2157,In_122,In_2033);
or U2158 (N_2158,In_1659,In_554);
nor U2159 (N_2159,In_1721,In_2044);
and U2160 (N_2160,In_690,In_607);
nand U2161 (N_2161,In_1588,In_903);
nor U2162 (N_2162,In_1376,In_1175);
nand U2163 (N_2163,In_2397,In_400);
or U2164 (N_2164,In_1743,In_2103);
or U2165 (N_2165,In_398,In_1962);
and U2166 (N_2166,In_1744,In_2441);
nor U2167 (N_2167,In_5,In_567);
xnor U2168 (N_2168,In_74,In_1465);
nor U2169 (N_2169,In_2067,In_1941);
xnor U2170 (N_2170,In_719,In_1840);
and U2171 (N_2171,In_206,In_925);
or U2172 (N_2172,In_1718,In_355);
or U2173 (N_2173,In_2467,In_2447);
and U2174 (N_2174,In_1986,In_409);
xor U2175 (N_2175,In_2376,In_248);
or U2176 (N_2176,In_2452,In_2074);
xor U2177 (N_2177,In_62,In_1956);
and U2178 (N_2178,In_827,In_2032);
nor U2179 (N_2179,In_1233,In_1215);
nor U2180 (N_2180,In_1664,In_755);
nor U2181 (N_2181,In_72,In_1180);
or U2182 (N_2182,In_306,In_1334);
xnor U2183 (N_2183,In_2284,In_1927);
or U2184 (N_2184,In_241,In_2002);
nand U2185 (N_2185,In_394,In_592);
nand U2186 (N_2186,In_1223,In_2355);
and U2187 (N_2187,In_449,In_2238);
xor U2188 (N_2188,In_1648,In_1640);
and U2189 (N_2189,In_2421,In_199);
xnor U2190 (N_2190,In_313,In_2266);
and U2191 (N_2191,In_563,In_2316);
nor U2192 (N_2192,In_204,In_189);
xor U2193 (N_2193,In_2386,In_1374);
and U2194 (N_2194,In_1452,In_522);
nand U2195 (N_2195,In_879,In_930);
nor U2196 (N_2196,In_2146,In_682);
nor U2197 (N_2197,In_1955,In_2257);
nor U2198 (N_2198,In_1938,In_1548);
xnor U2199 (N_2199,In_1571,In_856);
nand U2200 (N_2200,In_494,In_101);
nor U2201 (N_2201,In_829,In_1855);
and U2202 (N_2202,In_856,In_2035);
or U2203 (N_2203,In_968,In_514);
nand U2204 (N_2204,In_2374,In_869);
and U2205 (N_2205,In_2495,In_1970);
and U2206 (N_2206,In_2387,In_442);
xnor U2207 (N_2207,In_2461,In_191);
or U2208 (N_2208,In_1882,In_769);
nand U2209 (N_2209,In_1137,In_147);
nor U2210 (N_2210,In_1547,In_119);
xnor U2211 (N_2211,In_2113,In_2272);
nor U2212 (N_2212,In_977,In_1986);
xor U2213 (N_2213,In_2364,In_23);
or U2214 (N_2214,In_2168,In_1137);
nor U2215 (N_2215,In_2420,In_291);
xnor U2216 (N_2216,In_2486,In_466);
nor U2217 (N_2217,In_25,In_1337);
xor U2218 (N_2218,In_1893,In_1074);
nand U2219 (N_2219,In_985,In_777);
and U2220 (N_2220,In_1661,In_1268);
nor U2221 (N_2221,In_1478,In_1569);
nand U2222 (N_2222,In_1254,In_588);
xnor U2223 (N_2223,In_827,In_855);
and U2224 (N_2224,In_1662,In_1579);
and U2225 (N_2225,In_2018,In_1647);
nand U2226 (N_2226,In_2372,In_1749);
nor U2227 (N_2227,In_1205,In_1024);
xor U2228 (N_2228,In_215,In_1277);
xor U2229 (N_2229,In_2062,In_490);
nand U2230 (N_2230,In_170,In_865);
or U2231 (N_2231,In_845,In_395);
nor U2232 (N_2232,In_2345,In_891);
and U2233 (N_2233,In_1684,In_152);
xnor U2234 (N_2234,In_2070,In_2);
or U2235 (N_2235,In_1317,In_538);
nand U2236 (N_2236,In_242,In_2039);
nand U2237 (N_2237,In_1283,In_518);
nor U2238 (N_2238,In_2115,In_1927);
nand U2239 (N_2239,In_1549,In_831);
and U2240 (N_2240,In_1180,In_2365);
or U2241 (N_2241,In_1070,In_1186);
xor U2242 (N_2242,In_1622,In_1265);
nor U2243 (N_2243,In_0,In_962);
and U2244 (N_2244,In_2263,In_652);
nor U2245 (N_2245,In_1301,In_2236);
xor U2246 (N_2246,In_2069,In_1910);
nor U2247 (N_2247,In_2398,In_496);
nand U2248 (N_2248,In_975,In_1067);
or U2249 (N_2249,In_2476,In_1784);
xnor U2250 (N_2250,In_998,In_1894);
or U2251 (N_2251,In_2191,In_555);
or U2252 (N_2252,In_761,In_192);
nor U2253 (N_2253,In_1932,In_2066);
and U2254 (N_2254,In_575,In_827);
or U2255 (N_2255,In_2369,In_1070);
or U2256 (N_2256,In_2267,In_1208);
nor U2257 (N_2257,In_1165,In_1135);
or U2258 (N_2258,In_1553,In_1231);
and U2259 (N_2259,In_259,In_166);
nand U2260 (N_2260,In_718,In_958);
and U2261 (N_2261,In_147,In_1966);
xnor U2262 (N_2262,In_108,In_2171);
nor U2263 (N_2263,In_793,In_874);
xnor U2264 (N_2264,In_1044,In_1579);
and U2265 (N_2265,In_1051,In_582);
and U2266 (N_2266,In_994,In_1284);
nor U2267 (N_2267,In_2113,In_2087);
nor U2268 (N_2268,In_1210,In_2240);
or U2269 (N_2269,In_1035,In_495);
and U2270 (N_2270,In_2025,In_1273);
nand U2271 (N_2271,In_1384,In_56);
nor U2272 (N_2272,In_841,In_2057);
or U2273 (N_2273,In_1626,In_1283);
or U2274 (N_2274,In_1149,In_1781);
nor U2275 (N_2275,In_1154,In_2021);
xor U2276 (N_2276,In_758,In_526);
and U2277 (N_2277,In_811,In_2383);
and U2278 (N_2278,In_1558,In_137);
or U2279 (N_2279,In_371,In_1977);
nand U2280 (N_2280,In_1841,In_801);
nor U2281 (N_2281,In_1556,In_1165);
and U2282 (N_2282,In_1712,In_1135);
nor U2283 (N_2283,In_1343,In_52);
and U2284 (N_2284,In_1440,In_220);
nor U2285 (N_2285,In_59,In_2442);
xnor U2286 (N_2286,In_1149,In_1709);
xor U2287 (N_2287,In_539,In_425);
and U2288 (N_2288,In_1106,In_692);
nor U2289 (N_2289,In_1167,In_12);
nor U2290 (N_2290,In_1212,In_1503);
and U2291 (N_2291,In_171,In_985);
xnor U2292 (N_2292,In_584,In_653);
and U2293 (N_2293,In_2110,In_1110);
nor U2294 (N_2294,In_2239,In_697);
and U2295 (N_2295,In_893,In_1004);
and U2296 (N_2296,In_2303,In_911);
nor U2297 (N_2297,In_2051,In_662);
or U2298 (N_2298,In_1221,In_383);
xnor U2299 (N_2299,In_941,In_1297);
nand U2300 (N_2300,In_93,In_965);
and U2301 (N_2301,In_2388,In_1590);
or U2302 (N_2302,In_1348,In_1804);
and U2303 (N_2303,In_1715,In_959);
and U2304 (N_2304,In_318,In_1049);
and U2305 (N_2305,In_2434,In_654);
nand U2306 (N_2306,In_2061,In_1282);
xnor U2307 (N_2307,In_2239,In_1095);
or U2308 (N_2308,In_293,In_1326);
nand U2309 (N_2309,In_2429,In_178);
or U2310 (N_2310,In_2468,In_943);
nor U2311 (N_2311,In_2133,In_1198);
nand U2312 (N_2312,In_1849,In_1551);
or U2313 (N_2313,In_775,In_423);
nor U2314 (N_2314,In_988,In_1318);
nor U2315 (N_2315,In_862,In_1348);
xor U2316 (N_2316,In_1972,In_1062);
nand U2317 (N_2317,In_1023,In_1866);
nand U2318 (N_2318,In_1335,In_1573);
xnor U2319 (N_2319,In_1684,In_1427);
nand U2320 (N_2320,In_1983,In_436);
or U2321 (N_2321,In_1413,In_187);
and U2322 (N_2322,In_1850,In_1622);
nor U2323 (N_2323,In_1760,In_1387);
and U2324 (N_2324,In_711,In_1361);
nand U2325 (N_2325,In_1219,In_2413);
nor U2326 (N_2326,In_2212,In_2457);
or U2327 (N_2327,In_1976,In_1183);
nand U2328 (N_2328,In_284,In_1653);
nand U2329 (N_2329,In_2176,In_376);
or U2330 (N_2330,In_1721,In_266);
nand U2331 (N_2331,In_2376,In_1459);
and U2332 (N_2332,In_376,In_2449);
nor U2333 (N_2333,In_776,In_375);
nor U2334 (N_2334,In_1433,In_1825);
nor U2335 (N_2335,In_1240,In_1434);
or U2336 (N_2336,In_2428,In_1842);
xor U2337 (N_2337,In_739,In_1896);
xor U2338 (N_2338,In_2073,In_614);
nor U2339 (N_2339,In_2010,In_627);
nor U2340 (N_2340,In_995,In_2328);
or U2341 (N_2341,In_160,In_615);
xor U2342 (N_2342,In_1666,In_1188);
xor U2343 (N_2343,In_1168,In_617);
nand U2344 (N_2344,In_569,In_2353);
or U2345 (N_2345,In_1359,In_27);
and U2346 (N_2346,In_2261,In_2225);
xnor U2347 (N_2347,In_2094,In_248);
or U2348 (N_2348,In_2298,In_96);
nand U2349 (N_2349,In_2116,In_1312);
nand U2350 (N_2350,In_296,In_1623);
and U2351 (N_2351,In_1305,In_1121);
nand U2352 (N_2352,In_909,In_1897);
nor U2353 (N_2353,In_844,In_2214);
or U2354 (N_2354,In_367,In_752);
or U2355 (N_2355,In_658,In_1534);
nor U2356 (N_2356,In_426,In_693);
nand U2357 (N_2357,In_1319,In_1239);
xnor U2358 (N_2358,In_2051,In_137);
xor U2359 (N_2359,In_708,In_1546);
and U2360 (N_2360,In_1342,In_1206);
nand U2361 (N_2361,In_50,In_1368);
or U2362 (N_2362,In_1774,In_1196);
xor U2363 (N_2363,In_2278,In_1500);
nor U2364 (N_2364,In_22,In_2108);
nor U2365 (N_2365,In_155,In_1700);
and U2366 (N_2366,In_1148,In_224);
nand U2367 (N_2367,In_334,In_612);
nor U2368 (N_2368,In_898,In_2156);
or U2369 (N_2369,In_1705,In_1172);
and U2370 (N_2370,In_2183,In_2059);
xor U2371 (N_2371,In_2435,In_2124);
nand U2372 (N_2372,In_1948,In_208);
xor U2373 (N_2373,In_1425,In_405);
nand U2374 (N_2374,In_953,In_1174);
or U2375 (N_2375,In_2296,In_1557);
nor U2376 (N_2376,In_1410,In_683);
xor U2377 (N_2377,In_1576,In_407);
and U2378 (N_2378,In_1780,In_1701);
and U2379 (N_2379,In_1778,In_501);
nor U2380 (N_2380,In_885,In_224);
or U2381 (N_2381,In_1609,In_1359);
and U2382 (N_2382,In_2031,In_2008);
nor U2383 (N_2383,In_148,In_755);
nand U2384 (N_2384,In_2286,In_1780);
nand U2385 (N_2385,In_1444,In_69);
xor U2386 (N_2386,In_2495,In_1299);
or U2387 (N_2387,In_1504,In_1344);
nor U2388 (N_2388,In_1294,In_1493);
nor U2389 (N_2389,In_42,In_526);
nor U2390 (N_2390,In_729,In_1374);
xnor U2391 (N_2391,In_545,In_640);
and U2392 (N_2392,In_1436,In_1149);
and U2393 (N_2393,In_769,In_63);
nand U2394 (N_2394,In_312,In_1911);
and U2395 (N_2395,In_1004,In_896);
nand U2396 (N_2396,In_1732,In_1957);
nand U2397 (N_2397,In_1071,In_1866);
nand U2398 (N_2398,In_8,In_2067);
nor U2399 (N_2399,In_815,In_464);
xor U2400 (N_2400,In_1799,In_267);
nor U2401 (N_2401,In_1087,In_2193);
nand U2402 (N_2402,In_686,In_1535);
or U2403 (N_2403,In_643,In_105);
xor U2404 (N_2404,In_211,In_554);
xnor U2405 (N_2405,In_1727,In_897);
nor U2406 (N_2406,In_39,In_892);
and U2407 (N_2407,In_2116,In_521);
and U2408 (N_2408,In_209,In_854);
and U2409 (N_2409,In_1001,In_1448);
or U2410 (N_2410,In_130,In_1679);
xnor U2411 (N_2411,In_1982,In_1232);
or U2412 (N_2412,In_2277,In_2179);
and U2413 (N_2413,In_357,In_620);
xor U2414 (N_2414,In_780,In_2423);
nand U2415 (N_2415,In_2428,In_499);
xor U2416 (N_2416,In_416,In_1147);
nor U2417 (N_2417,In_1411,In_1866);
nand U2418 (N_2418,In_430,In_2209);
or U2419 (N_2419,In_772,In_543);
or U2420 (N_2420,In_1106,In_2112);
nand U2421 (N_2421,In_1111,In_697);
xnor U2422 (N_2422,In_733,In_74);
and U2423 (N_2423,In_256,In_1046);
xor U2424 (N_2424,In_71,In_450);
nand U2425 (N_2425,In_1460,In_1178);
xnor U2426 (N_2426,In_433,In_1705);
nand U2427 (N_2427,In_739,In_1768);
nand U2428 (N_2428,In_1399,In_1769);
xnor U2429 (N_2429,In_1792,In_389);
xnor U2430 (N_2430,In_1575,In_2415);
xnor U2431 (N_2431,In_1395,In_1107);
nand U2432 (N_2432,In_2304,In_1240);
or U2433 (N_2433,In_855,In_1482);
or U2434 (N_2434,In_2485,In_1292);
xnor U2435 (N_2435,In_1616,In_451);
and U2436 (N_2436,In_1504,In_1172);
xnor U2437 (N_2437,In_1503,In_1425);
xor U2438 (N_2438,In_883,In_2294);
or U2439 (N_2439,In_406,In_401);
and U2440 (N_2440,In_1766,In_1432);
xnor U2441 (N_2441,In_483,In_2473);
nand U2442 (N_2442,In_2495,In_2214);
xnor U2443 (N_2443,In_78,In_1319);
xor U2444 (N_2444,In_974,In_254);
and U2445 (N_2445,In_223,In_1688);
nor U2446 (N_2446,In_1324,In_1989);
and U2447 (N_2447,In_799,In_1456);
nor U2448 (N_2448,In_1090,In_2264);
nand U2449 (N_2449,In_738,In_653);
and U2450 (N_2450,In_222,In_921);
and U2451 (N_2451,In_951,In_2410);
and U2452 (N_2452,In_471,In_1155);
xor U2453 (N_2453,In_2,In_741);
and U2454 (N_2454,In_243,In_627);
or U2455 (N_2455,In_1693,In_1240);
or U2456 (N_2456,In_633,In_615);
or U2457 (N_2457,In_1768,In_1434);
and U2458 (N_2458,In_362,In_537);
nand U2459 (N_2459,In_1718,In_956);
and U2460 (N_2460,In_1038,In_438);
xnor U2461 (N_2461,In_309,In_501);
and U2462 (N_2462,In_2215,In_464);
xor U2463 (N_2463,In_157,In_940);
nand U2464 (N_2464,In_1287,In_713);
or U2465 (N_2465,In_330,In_1964);
xor U2466 (N_2466,In_673,In_1429);
and U2467 (N_2467,In_2310,In_1486);
or U2468 (N_2468,In_234,In_1812);
or U2469 (N_2469,In_1358,In_905);
and U2470 (N_2470,In_1445,In_1739);
nor U2471 (N_2471,In_167,In_900);
nand U2472 (N_2472,In_512,In_2083);
xnor U2473 (N_2473,In_129,In_1222);
and U2474 (N_2474,In_1848,In_733);
nand U2475 (N_2475,In_532,In_317);
and U2476 (N_2476,In_1487,In_887);
nor U2477 (N_2477,In_2380,In_444);
or U2478 (N_2478,In_449,In_378);
and U2479 (N_2479,In_347,In_1663);
and U2480 (N_2480,In_2313,In_1196);
xor U2481 (N_2481,In_1545,In_1558);
nand U2482 (N_2482,In_1129,In_741);
or U2483 (N_2483,In_1992,In_66);
nand U2484 (N_2484,In_1336,In_1000);
and U2485 (N_2485,In_1881,In_2420);
nor U2486 (N_2486,In_1536,In_221);
xnor U2487 (N_2487,In_678,In_1732);
nor U2488 (N_2488,In_113,In_883);
nor U2489 (N_2489,In_1416,In_1456);
or U2490 (N_2490,In_410,In_669);
nand U2491 (N_2491,In_1523,In_181);
and U2492 (N_2492,In_2253,In_904);
nand U2493 (N_2493,In_1016,In_1422);
nand U2494 (N_2494,In_382,In_1100);
xor U2495 (N_2495,In_2282,In_551);
nor U2496 (N_2496,In_1296,In_1903);
or U2497 (N_2497,In_77,In_1274);
nor U2498 (N_2498,In_181,In_646);
and U2499 (N_2499,In_2109,In_1791);
nor U2500 (N_2500,In_172,In_1648);
and U2501 (N_2501,In_915,In_2337);
nor U2502 (N_2502,In_1126,In_1533);
xor U2503 (N_2503,In_1206,In_1151);
nor U2504 (N_2504,In_458,In_2359);
and U2505 (N_2505,In_807,In_1548);
nor U2506 (N_2506,In_708,In_700);
xor U2507 (N_2507,In_2131,In_2170);
or U2508 (N_2508,In_1366,In_1219);
nor U2509 (N_2509,In_89,In_1333);
and U2510 (N_2510,In_2397,In_816);
xnor U2511 (N_2511,In_1669,In_1051);
nand U2512 (N_2512,In_747,In_353);
xnor U2513 (N_2513,In_812,In_1682);
nand U2514 (N_2514,In_2210,In_2357);
xnor U2515 (N_2515,In_146,In_1875);
or U2516 (N_2516,In_1916,In_1761);
and U2517 (N_2517,In_2183,In_874);
and U2518 (N_2518,In_923,In_1201);
or U2519 (N_2519,In_1710,In_1197);
and U2520 (N_2520,In_1300,In_643);
xor U2521 (N_2521,In_1298,In_280);
xor U2522 (N_2522,In_1072,In_139);
nor U2523 (N_2523,In_2378,In_1155);
nor U2524 (N_2524,In_1225,In_283);
nand U2525 (N_2525,In_2433,In_1303);
nor U2526 (N_2526,In_1631,In_259);
nor U2527 (N_2527,In_1793,In_874);
nand U2528 (N_2528,In_1014,In_2460);
and U2529 (N_2529,In_1305,In_1843);
xnor U2530 (N_2530,In_6,In_177);
nor U2531 (N_2531,In_198,In_506);
nor U2532 (N_2532,In_990,In_1486);
nand U2533 (N_2533,In_306,In_2412);
and U2534 (N_2534,In_1691,In_2335);
nand U2535 (N_2535,In_2213,In_49);
xor U2536 (N_2536,In_990,In_2165);
and U2537 (N_2537,In_2122,In_2434);
xor U2538 (N_2538,In_693,In_901);
xnor U2539 (N_2539,In_667,In_1693);
or U2540 (N_2540,In_1281,In_432);
and U2541 (N_2541,In_94,In_1384);
or U2542 (N_2542,In_422,In_2019);
xnor U2543 (N_2543,In_1113,In_424);
nor U2544 (N_2544,In_1342,In_1476);
xor U2545 (N_2545,In_1224,In_1834);
or U2546 (N_2546,In_1616,In_971);
and U2547 (N_2547,In_1965,In_428);
nand U2548 (N_2548,In_267,In_1101);
nor U2549 (N_2549,In_2157,In_815);
or U2550 (N_2550,In_1210,In_1875);
nand U2551 (N_2551,In_2112,In_1158);
nor U2552 (N_2552,In_789,In_916);
nand U2553 (N_2553,In_1479,In_2328);
nor U2554 (N_2554,In_2487,In_1856);
nand U2555 (N_2555,In_615,In_385);
nor U2556 (N_2556,In_381,In_1615);
nor U2557 (N_2557,In_1900,In_1807);
nor U2558 (N_2558,In_851,In_196);
or U2559 (N_2559,In_1747,In_1509);
and U2560 (N_2560,In_175,In_1578);
or U2561 (N_2561,In_16,In_706);
nor U2562 (N_2562,In_658,In_59);
or U2563 (N_2563,In_944,In_937);
xnor U2564 (N_2564,In_1330,In_1951);
nor U2565 (N_2565,In_1841,In_704);
nand U2566 (N_2566,In_1479,In_620);
nand U2567 (N_2567,In_1153,In_2483);
nor U2568 (N_2568,In_513,In_1002);
nand U2569 (N_2569,In_2315,In_153);
xnor U2570 (N_2570,In_1609,In_2249);
nor U2571 (N_2571,In_2064,In_2220);
nor U2572 (N_2572,In_1413,In_1279);
nor U2573 (N_2573,In_567,In_2367);
and U2574 (N_2574,In_2442,In_1255);
and U2575 (N_2575,In_686,In_527);
nand U2576 (N_2576,In_1999,In_90);
or U2577 (N_2577,In_2339,In_1361);
nand U2578 (N_2578,In_2315,In_959);
nor U2579 (N_2579,In_663,In_2120);
nor U2580 (N_2580,In_1351,In_1229);
nor U2581 (N_2581,In_2414,In_1568);
nand U2582 (N_2582,In_1065,In_1497);
or U2583 (N_2583,In_1126,In_1281);
or U2584 (N_2584,In_1160,In_1013);
and U2585 (N_2585,In_301,In_2412);
nand U2586 (N_2586,In_2396,In_2337);
nand U2587 (N_2587,In_1194,In_1811);
xnor U2588 (N_2588,In_1126,In_1188);
and U2589 (N_2589,In_2003,In_410);
nor U2590 (N_2590,In_589,In_554);
and U2591 (N_2591,In_2310,In_1913);
nand U2592 (N_2592,In_2103,In_753);
or U2593 (N_2593,In_2129,In_1578);
and U2594 (N_2594,In_1233,In_834);
and U2595 (N_2595,In_197,In_95);
xor U2596 (N_2596,In_100,In_557);
xor U2597 (N_2597,In_520,In_2224);
nor U2598 (N_2598,In_2057,In_1704);
nor U2599 (N_2599,In_91,In_662);
or U2600 (N_2600,In_2022,In_1949);
and U2601 (N_2601,In_81,In_1763);
xor U2602 (N_2602,In_1433,In_2318);
nor U2603 (N_2603,In_978,In_1906);
and U2604 (N_2604,In_2471,In_2227);
or U2605 (N_2605,In_1714,In_1786);
xor U2606 (N_2606,In_2261,In_2346);
nor U2607 (N_2607,In_2472,In_501);
or U2608 (N_2608,In_1879,In_1064);
xor U2609 (N_2609,In_1913,In_1880);
nor U2610 (N_2610,In_1736,In_1171);
nand U2611 (N_2611,In_383,In_1797);
and U2612 (N_2612,In_2486,In_436);
and U2613 (N_2613,In_415,In_1869);
and U2614 (N_2614,In_2421,In_2064);
nand U2615 (N_2615,In_2396,In_1638);
nand U2616 (N_2616,In_943,In_360);
or U2617 (N_2617,In_709,In_2008);
and U2618 (N_2618,In_1782,In_2337);
nor U2619 (N_2619,In_2209,In_1593);
xor U2620 (N_2620,In_1366,In_1585);
nand U2621 (N_2621,In_905,In_705);
or U2622 (N_2622,In_1751,In_596);
xor U2623 (N_2623,In_1953,In_180);
or U2624 (N_2624,In_1115,In_415);
xor U2625 (N_2625,In_581,In_1719);
nor U2626 (N_2626,In_2332,In_2007);
xor U2627 (N_2627,In_2145,In_1686);
and U2628 (N_2628,In_1961,In_1830);
or U2629 (N_2629,In_1454,In_137);
nand U2630 (N_2630,In_738,In_2088);
xnor U2631 (N_2631,In_184,In_1961);
nand U2632 (N_2632,In_1357,In_907);
xor U2633 (N_2633,In_1845,In_373);
xor U2634 (N_2634,In_608,In_536);
and U2635 (N_2635,In_2189,In_1409);
and U2636 (N_2636,In_480,In_814);
xor U2637 (N_2637,In_2399,In_2387);
or U2638 (N_2638,In_73,In_260);
nand U2639 (N_2639,In_1265,In_1530);
xor U2640 (N_2640,In_1963,In_1880);
nor U2641 (N_2641,In_1086,In_1780);
and U2642 (N_2642,In_894,In_1009);
nor U2643 (N_2643,In_2247,In_2401);
nor U2644 (N_2644,In_1650,In_2183);
xor U2645 (N_2645,In_875,In_1761);
nand U2646 (N_2646,In_1990,In_1492);
or U2647 (N_2647,In_1137,In_52);
or U2648 (N_2648,In_159,In_762);
xnor U2649 (N_2649,In_405,In_930);
xor U2650 (N_2650,In_918,In_1231);
nand U2651 (N_2651,In_406,In_613);
nor U2652 (N_2652,In_225,In_1906);
or U2653 (N_2653,In_444,In_1966);
nor U2654 (N_2654,In_814,In_1435);
xnor U2655 (N_2655,In_2231,In_1646);
nor U2656 (N_2656,In_628,In_1190);
or U2657 (N_2657,In_2307,In_1228);
nor U2658 (N_2658,In_1156,In_89);
nand U2659 (N_2659,In_729,In_370);
xnor U2660 (N_2660,In_2392,In_2297);
or U2661 (N_2661,In_640,In_1810);
and U2662 (N_2662,In_1178,In_908);
nand U2663 (N_2663,In_45,In_2433);
nand U2664 (N_2664,In_442,In_1111);
and U2665 (N_2665,In_1430,In_1123);
or U2666 (N_2666,In_1645,In_2271);
nor U2667 (N_2667,In_1610,In_1258);
nor U2668 (N_2668,In_1382,In_2220);
xor U2669 (N_2669,In_1218,In_1630);
xnor U2670 (N_2670,In_752,In_1109);
or U2671 (N_2671,In_2336,In_1678);
or U2672 (N_2672,In_50,In_1281);
or U2673 (N_2673,In_298,In_2259);
or U2674 (N_2674,In_672,In_1924);
or U2675 (N_2675,In_1853,In_2225);
nor U2676 (N_2676,In_1603,In_995);
xor U2677 (N_2677,In_642,In_1080);
and U2678 (N_2678,In_1037,In_1886);
xnor U2679 (N_2679,In_2427,In_2410);
xnor U2680 (N_2680,In_809,In_1442);
or U2681 (N_2681,In_2467,In_491);
nor U2682 (N_2682,In_2430,In_960);
xnor U2683 (N_2683,In_1638,In_16);
nor U2684 (N_2684,In_1173,In_977);
xnor U2685 (N_2685,In_1253,In_1781);
and U2686 (N_2686,In_1819,In_1986);
or U2687 (N_2687,In_1459,In_1376);
xnor U2688 (N_2688,In_482,In_1187);
and U2689 (N_2689,In_509,In_16);
xor U2690 (N_2690,In_3,In_1610);
and U2691 (N_2691,In_97,In_2060);
nand U2692 (N_2692,In_1475,In_1897);
nand U2693 (N_2693,In_1610,In_1750);
nor U2694 (N_2694,In_668,In_1835);
nor U2695 (N_2695,In_2276,In_1538);
or U2696 (N_2696,In_1713,In_1070);
nand U2697 (N_2697,In_1550,In_2093);
xnor U2698 (N_2698,In_1025,In_378);
nor U2699 (N_2699,In_1672,In_1579);
xor U2700 (N_2700,In_729,In_1775);
nor U2701 (N_2701,In_571,In_2456);
and U2702 (N_2702,In_133,In_433);
nor U2703 (N_2703,In_2407,In_1429);
or U2704 (N_2704,In_1338,In_1060);
nor U2705 (N_2705,In_2036,In_873);
or U2706 (N_2706,In_633,In_207);
nand U2707 (N_2707,In_1256,In_1751);
nor U2708 (N_2708,In_1054,In_71);
nor U2709 (N_2709,In_576,In_2198);
or U2710 (N_2710,In_678,In_166);
nor U2711 (N_2711,In_456,In_2406);
nand U2712 (N_2712,In_2452,In_877);
and U2713 (N_2713,In_2095,In_872);
or U2714 (N_2714,In_2047,In_751);
xnor U2715 (N_2715,In_87,In_1493);
nor U2716 (N_2716,In_788,In_1160);
xor U2717 (N_2717,In_1269,In_2118);
nand U2718 (N_2718,In_544,In_1026);
xnor U2719 (N_2719,In_1930,In_483);
xor U2720 (N_2720,In_1589,In_612);
and U2721 (N_2721,In_393,In_1359);
xor U2722 (N_2722,In_1273,In_2258);
and U2723 (N_2723,In_1792,In_1498);
nand U2724 (N_2724,In_741,In_1255);
nand U2725 (N_2725,In_1595,In_123);
nor U2726 (N_2726,In_214,In_1463);
nor U2727 (N_2727,In_2249,In_1235);
and U2728 (N_2728,In_325,In_2273);
nor U2729 (N_2729,In_304,In_311);
nor U2730 (N_2730,In_2214,In_901);
nand U2731 (N_2731,In_2211,In_2147);
xor U2732 (N_2732,In_1804,In_1979);
and U2733 (N_2733,In_673,In_2045);
or U2734 (N_2734,In_849,In_2031);
nand U2735 (N_2735,In_1051,In_2485);
and U2736 (N_2736,In_2246,In_328);
or U2737 (N_2737,In_1295,In_377);
nor U2738 (N_2738,In_222,In_158);
nand U2739 (N_2739,In_1009,In_1281);
and U2740 (N_2740,In_1716,In_1484);
and U2741 (N_2741,In_1390,In_1923);
nand U2742 (N_2742,In_1183,In_562);
nand U2743 (N_2743,In_2441,In_67);
xor U2744 (N_2744,In_33,In_1560);
nor U2745 (N_2745,In_1817,In_1666);
nor U2746 (N_2746,In_1642,In_1534);
xnor U2747 (N_2747,In_1439,In_530);
nor U2748 (N_2748,In_1787,In_1367);
and U2749 (N_2749,In_2198,In_2139);
nand U2750 (N_2750,In_1655,In_477);
nand U2751 (N_2751,In_145,In_1409);
nand U2752 (N_2752,In_110,In_1359);
xor U2753 (N_2753,In_1005,In_1962);
nand U2754 (N_2754,In_1967,In_272);
nor U2755 (N_2755,In_1640,In_1592);
and U2756 (N_2756,In_362,In_71);
nand U2757 (N_2757,In_2011,In_863);
nor U2758 (N_2758,In_423,In_1602);
or U2759 (N_2759,In_546,In_913);
or U2760 (N_2760,In_1227,In_1643);
nor U2761 (N_2761,In_2482,In_337);
nand U2762 (N_2762,In_1911,In_2457);
or U2763 (N_2763,In_5,In_1894);
xor U2764 (N_2764,In_2340,In_171);
nand U2765 (N_2765,In_1446,In_1078);
or U2766 (N_2766,In_1738,In_401);
and U2767 (N_2767,In_28,In_1161);
and U2768 (N_2768,In_2239,In_312);
xor U2769 (N_2769,In_2258,In_2024);
and U2770 (N_2770,In_240,In_1761);
and U2771 (N_2771,In_2337,In_2354);
and U2772 (N_2772,In_1540,In_613);
nor U2773 (N_2773,In_1261,In_683);
nand U2774 (N_2774,In_2037,In_342);
nor U2775 (N_2775,In_1961,In_1306);
nand U2776 (N_2776,In_228,In_1015);
xnor U2777 (N_2777,In_1945,In_747);
nor U2778 (N_2778,In_1149,In_2345);
nor U2779 (N_2779,In_44,In_2294);
xnor U2780 (N_2780,In_2380,In_2336);
xnor U2781 (N_2781,In_106,In_2196);
and U2782 (N_2782,In_749,In_1912);
nor U2783 (N_2783,In_653,In_1637);
or U2784 (N_2784,In_1007,In_1500);
or U2785 (N_2785,In_500,In_686);
nand U2786 (N_2786,In_2349,In_515);
xor U2787 (N_2787,In_2200,In_356);
or U2788 (N_2788,In_155,In_461);
or U2789 (N_2789,In_965,In_1644);
and U2790 (N_2790,In_1450,In_1141);
nor U2791 (N_2791,In_1539,In_1768);
and U2792 (N_2792,In_2148,In_831);
xnor U2793 (N_2793,In_148,In_2006);
nand U2794 (N_2794,In_476,In_1434);
xnor U2795 (N_2795,In_311,In_774);
xnor U2796 (N_2796,In_809,In_1007);
and U2797 (N_2797,In_1160,In_233);
nand U2798 (N_2798,In_1000,In_328);
or U2799 (N_2799,In_1320,In_785);
and U2800 (N_2800,In_2212,In_252);
and U2801 (N_2801,In_2202,In_1557);
nand U2802 (N_2802,In_1425,In_2494);
nor U2803 (N_2803,In_710,In_278);
xnor U2804 (N_2804,In_340,In_1038);
xnor U2805 (N_2805,In_1324,In_706);
or U2806 (N_2806,In_1712,In_1934);
or U2807 (N_2807,In_42,In_1845);
or U2808 (N_2808,In_2328,In_1910);
or U2809 (N_2809,In_2409,In_1285);
nand U2810 (N_2810,In_2492,In_1235);
nand U2811 (N_2811,In_1819,In_1548);
or U2812 (N_2812,In_275,In_2468);
nor U2813 (N_2813,In_1913,In_1893);
or U2814 (N_2814,In_2073,In_209);
nor U2815 (N_2815,In_360,In_634);
nand U2816 (N_2816,In_2135,In_2328);
or U2817 (N_2817,In_2435,In_509);
xor U2818 (N_2818,In_2333,In_1806);
nor U2819 (N_2819,In_999,In_1976);
and U2820 (N_2820,In_2472,In_790);
and U2821 (N_2821,In_955,In_604);
xnor U2822 (N_2822,In_580,In_1236);
and U2823 (N_2823,In_551,In_754);
and U2824 (N_2824,In_1220,In_1717);
nor U2825 (N_2825,In_1517,In_309);
nand U2826 (N_2826,In_1341,In_580);
nor U2827 (N_2827,In_616,In_1237);
and U2828 (N_2828,In_2373,In_1267);
nand U2829 (N_2829,In_430,In_628);
nor U2830 (N_2830,In_1909,In_251);
and U2831 (N_2831,In_1694,In_1674);
and U2832 (N_2832,In_1240,In_1322);
or U2833 (N_2833,In_1609,In_2402);
nand U2834 (N_2834,In_827,In_2244);
nor U2835 (N_2835,In_367,In_2402);
nor U2836 (N_2836,In_1421,In_833);
and U2837 (N_2837,In_1058,In_2420);
nand U2838 (N_2838,In_2118,In_450);
nand U2839 (N_2839,In_2096,In_1187);
nor U2840 (N_2840,In_591,In_545);
and U2841 (N_2841,In_1344,In_611);
nor U2842 (N_2842,In_268,In_30);
nor U2843 (N_2843,In_1040,In_183);
xnor U2844 (N_2844,In_2434,In_715);
and U2845 (N_2845,In_224,In_1063);
nand U2846 (N_2846,In_1016,In_1641);
or U2847 (N_2847,In_1728,In_1467);
nand U2848 (N_2848,In_2031,In_1817);
or U2849 (N_2849,In_603,In_1715);
xor U2850 (N_2850,In_934,In_675);
xor U2851 (N_2851,In_1844,In_1726);
xnor U2852 (N_2852,In_846,In_1743);
and U2853 (N_2853,In_93,In_1325);
xnor U2854 (N_2854,In_490,In_1506);
or U2855 (N_2855,In_814,In_66);
or U2856 (N_2856,In_2060,In_61);
or U2857 (N_2857,In_2438,In_1565);
or U2858 (N_2858,In_55,In_680);
and U2859 (N_2859,In_560,In_1002);
nand U2860 (N_2860,In_360,In_1309);
xor U2861 (N_2861,In_774,In_1168);
nand U2862 (N_2862,In_465,In_1257);
nor U2863 (N_2863,In_1622,In_714);
nor U2864 (N_2864,In_137,In_1912);
or U2865 (N_2865,In_35,In_1056);
nand U2866 (N_2866,In_304,In_1189);
nand U2867 (N_2867,In_2340,In_2019);
nor U2868 (N_2868,In_1791,In_1964);
xor U2869 (N_2869,In_43,In_1774);
xor U2870 (N_2870,In_1312,In_997);
and U2871 (N_2871,In_848,In_1958);
nor U2872 (N_2872,In_438,In_1421);
nor U2873 (N_2873,In_1694,In_467);
nor U2874 (N_2874,In_402,In_1511);
nor U2875 (N_2875,In_1096,In_1282);
xnor U2876 (N_2876,In_2396,In_676);
xnor U2877 (N_2877,In_199,In_1446);
nor U2878 (N_2878,In_1066,In_1915);
nand U2879 (N_2879,In_254,In_1294);
nand U2880 (N_2880,In_567,In_971);
nor U2881 (N_2881,In_846,In_1527);
nor U2882 (N_2882,In_2304,In_1327);
and U2883 (N_2883,In_2047,In_884);
xnor U2884 (N_2884,In_1072,In_2445);
and U2885 (N_2885,In_1973,In_224);
or U2886 (N_2886,In_2017,In_545);
and U2887 (N_2887,In_1717,In_88);
nor U2888 (N_2888,In_1708,In_733);
nand U2889 (N_2889,In_1048,In_523);
nand U2890 (N_2890,In_1700,In_1550);
and U2891 (N_2891,In_2428,In_1140);
or U2892 (N_2892,In_420,In_1243);
nor U2893 (N_2893,In_2398,In_709);
or U2894 (N_2894,In_441,In_1230);
and U2895 (N_2895,In_1428,In_2097);
nor U2896 (N_2896,In_2378,In_1469);
and U2897 (N_2897,In_2290,In_2482);
nand U2898 (N_2898,In_508,In_2307);
nor U2899 (N_2899,In_572,In_857);
and U2900 (N_2900,In_2059,In_1);
xnor U2901 (N_2901,In_1022,In_2323);
and U2902 (N_2902,In_914,In_1570);
nand U2903 (N_2903,In_825,In_1473);
and U2904 (N_2904,In_1525,In_1987);
nand U2905 (N_2905,In_2215,In_214);
and U2906 (N_2906,In_150,In_1863);
nand U2907 (N_2907,In_1236,In_2056);
and U2908 (N_2908,In_140,In_2123);
nor U2909 (N_2909,In_685,In_670);
and U2910 (N_2910,In_317,In_1357);
nor U2911 (N_2911,In_1983,In_2375);
nor U2912 (N_2912,In_1555,In_1408);
and U2913 (N_2913,In_198,In_1348);
xnor U2914 (N_2914,In_1678,In_485);
nand U2915 (N_2915,In_1267,In_1123);
nand U2916 (N_2916,In_934,In_1126);
nor U2917 (N_2917,In_529,In_463);
xor U2918 (N_2918,In_1734,In_805);
and U2919 (N_2919,In_2118,In_2274);
and U2920 (N_2920,In_2145,In_1303);
and U2921 (N_2921,In_1110,In_53);
or U2922 (N_2922,In_1931,In_1239);
xnor U2923 (N_2923,In_443,In_1351);
and U2924 (N_2924,In_1746,In_1881);
xnor U2925 (N_2925,In_1984,In_2021);
or U2926 (N_2926,In_2363,In_1349);
xnor U2927 (N_2927,In_1888,In_438);
and U2928 (N_2928,In_2410,In_2436);
nand U2929 (N_2929,In_1877,In_1362);
nand U2930 (N_2930,In_228,In_2313);
and U2931 (N_2931,In_10,In_2353);
nor U2932 (N_2932,In_725,In_997);
nand U2933 (N_2933,In_2276,In_1083);
xnor U2934 (N_2934,In_1325,In_1263);
or U2935 (N_2935,In_124,In_863);
nor U2936 (N_2936,In_460,In_2454);
or U2937 (N_2937,In_1541,In_2424);
and U2938 (N_2938,In_604,In_818);
and U2939 (N_2939,In_1884,In_2009);
or U2940 (N_2940,In_1751,In_1841);
or U2941 (N_2941,In_1721,In_65);
xor U2942 (N_2942,In_1917,In_648);
or U2943 (N_2943,In_1942,In_632);
xor U2944 (N_2944,In_2496,In_1509);
and U2945 (N_2945,In_703,In_1944);
or U2946 (N_2946,In_765,In_1940);
or U2947 (N_2947,In_716,In_2352);
and U2948 (N_2948,In_409,In_2052);
xnor U2949 (N_2949,In_1129,In_936);
nor U2950 (N_2950,In_1732,In_677);
or U2951 (N_2951,In_399,In_230);
nand U2952 (N_2952,In_301,In_572);
nor U2953 (N_2953,In_1531,In_1960);
nor U2954 (N_2954,In_724,In_1690);
nor U2955 (N_2955,In_2007,In_623);
nand U2956 (N_2956,In_683,In_2174);
xor U2957 (N_2957,In_115,In_2269);
and U2958 (N_2958,In_577,In_2213);
nor U2959 (N_2959,In_1393,In_1364);
and U2960 (N_2960,In_1259,In_1691);
or U2961 (N_2961,In_695,In_177);
nand U2962 (N_2962,In_441,In_2274);
or U2963 (N_2963,In_2127,In_2399);
nor U2964 (N_2964,In_2081,In_1903);
nand U2965 (N_2965,In_97,In_1549);
or U2966 (N_2966,In_440,In_669);
nand U2967 (N_2967,In_2399,In_1624);
and U2968 (N_2968,In_1562,In_725);
and U2969 (N_2969,In_2352,In_473);
nor U2970 (N_2970,In_1935,In_467);
nand U2971 (N_2971,In_371,In_13);
and U2972 (N_2972,In_1591,In_508);
nand U2973 (N_2973,In_1535,In_1325);
and U2974 (N_2974,In_407,In_518);
nor U2975 (N_2975,In_1966,In_1122);
and U2976 (N_2976,In_776,In_198);
and U2977 (N_2977,In_1830,In_996);
nor U2978 (N_2978,In_1124,In_1929);
and U2979 (N_2979,In_1742,In_765);
and U2980 (N_2980,In_2048,In_2365);
or U2981 (N_2981,In_2242,In_1652);
or U2982 (N_2982,In_2494,In_915);
and U2983 (N_2983,In_50,In_1095);
and U2984 (N_2984,In_761,In_231);
nor U2985 (N_2985,In_1489,In_1640);
nor U2986 (N_2986,In_654,In_1067);
nor U2987 (N_2987,In_732,In_568);
and U2988 (N_2988,In_1029,In_901);
and U2989 (N_2989,In_1649,In_1188);
nand U2990 (N_2990,In_1040,In_1694);
or U2991 (N_2991,In_1675,In_2430);
or U2992 (N_2992,In_1704,In_1383);
and U2993 (N_2993,In_609,In_317);
xnor U2994 (N_2994,In_1470,In_1417);
xor U2995 (N_2995,In_341,In_1709);
xor U2996 (N_2996,In_93,In_583);
nand U2997 (N_2997,In_428,In_1983);
or U2998 (N_2998,In_876,In_2040);
and U2999 (N_2999,In_1607,In_1556);
or U3000 (N_3000,In_1382,In_2419);
and U3001 (N_3001,In_2332,In_1359);
or U3002 (N_3002,In_1515,In_1365);
nand U3003 (N_3003,In_1742,In_2427);
nor U3004 (N_3004,In_701,In_2493);
xnor U3005 (N_3005,In_1220,In_1237);
or U3006 (N_3006,In_1663,In_1787);
nand U3007 (N_3007,In_492,In_460);
and U3008 (N_3008,In_1015,In_1085);
xnor U3009 (N_3009,In_146,In_502);
xnor U3010 (N_3010,In_2296,In_985);
or U3011 (N_3011,In_399,In_1421);
or U3012 (N_3012,In_1960,In_2264);
nor U3013 (N_3013,In_2327,In_694);
nand U3014 (N_3014,In_1587,In_1639);
xor U3015 (N_3015,In_221,In_1462);
or U3016 (N_3016,In_347,In_1600);
or U3017 (N_3017,In_205,In_2229);
nand U3018 (N_3018,In_112,In_2409);
and U3019 (N_3019,In_624,In_1529);
nor U3020 (N_3020,In_2294,In_795);
xnor U3021 (N_3021,In_1519,In_411);
xor U3022 (N_3022,In_971,In_1920);
nand U3023 (N_3023,In_704,In_671);
and U3024 (N_3024,In_2157,In_1519);
and U3025 (N_3025,In_2093,In_870);
xnor U3026 (N_3026,In_728,In_1686);
xor U3027 (N_3027,In_1593,In_1802);
nand U3028 (N_3028,In_2045,In_372);
and U3029 (N_3029,In_941,In_2094);
or U3030 (N_3030,In_185,In_2403);
and U3031 (N_3031,In_1590,In_1120);
and U3032 (N_3032,In_1882,In_758);
nor U3033 (N_3033,In_218,In_326);
nand U3034 (N_3034,In_1495,In_1728);
or U3035 (N_3035,In_1376,In_913);
or U3036 (N_3036,In_2413,In_519);
nor U3037 (N_3037,In_1430,In_589);
nand U3038 (N_3038,In_791,In_215);
xnor U3039 (N_3039,In_2235,In_760);
or U3040 (N_3040,In_1339,In_581);
nand U3041 (N_3041,In_695,In_2187);
nand U3042 (N_3042,In_2262,In_2328);
or U3043 (N_3043,In_2241,In_32);
xnor U3044 (N_3044,In_799,In_626);
and U3045 (N_3045,In_371,In_1451);
and U3046 (N_3046,In_2488,In_2393);
xor U3047 (N_3047,In_1007,In_877);
and U3048 (N_3048,In_914,In_497);
nand U3049 (N_3049,In_923,In_1884);
and U3050 (N_3050,In_409,In_51);
and U3051 (N_3051,In_1866,In_1783);
or U3052 (N_3052,In_1345,In_489);
nand U3053 (N_3053,In_163,In_1951);
and U3054 (N_3054,In_1126,In_923);
nand U3055 (N_3055,In_1288,In_2063);
or U3056 (N_3056,In_762,In_2422);
and U3057 (N_3057,In_1805,In_2136);
nand U3058 (N_3058,In_973,In_826);
xor U3059 (N_3059,In_814,In_940);
nor U3060 (N_3060,In_2269,In_2428);
nand U3061 (N_3061,In_1438,In_782);
xnor U3062 (N_3062,In_1429,In_559);
nor U3063 (N_3063,In_2194,In_840);
nand U3064 (N_3064,In_700,In_2470);
xnor U3065 (N_3065,In_2034,In_1389);
and U3066 (N_3066,In_929,In_1068);
nand U3067 (N_3067,In_2261,In_2318);
nand U3068 (N_3068,In_773,In_85);
and U3069 (N_3069,In_1604,In_2211);
xnor U3070 (N_3070,In_1136,In_1863);
nor U3071 (N_3071,In_795,In_2160);
nor U3072 (N_3072,In_2455,In_2042);
or U3073 (N_3073,In_2008,In_20);
nor U3074 (N_3074,In_400,In_202);
or U3075 (N_3075,In_1978,In_1818);
or U3076 (N_3076,In_2452,In_632);
nor U3077 (N_3077,In_232,In_1635);
nand U3078 (N_3078,In_415,In_434);
nor U3079 (N_3079,In_938,In_978);
xnor U3080 (N_3080,In_678,In_2279);
nand U3081 (N_3081,In_2246,In_562);
xor U3082 (N_3082,In_2259,In_1896);
or U3083 (N_3083,In_1183,In_2464);
nor U3084 (N_3084,In_1551,In_538);
nand U3085 (N_3085,In_80,In_2145);
xor U3086 (N_3086,In_1166,In_1973);
xnor U3087 (N_3087,In_1843,In_508);
xor U3088 (N_3088,In_1448,In_1695);
nand U3089 (N_3089,In_1647,In_2482);
or U3090 (N_3090,In_302,In_449);
nor U3091 (N_3091,In_1112,In_1697);
xnor U3092 (N_3092,In_1317,In_2230);
nor U3093 (N_3093,In_1004,In_2056);
and U3094 (N_3094,In_269,In_2287);
or U3095 (N_3095,In_1458,In_1015);
nor U3096 (N_3096,In_2464,In_443);
nand U3097 (N_3097,In_1517,In_2270);
and U3098 (N_3098,In_1926,In_2367);
and U3099 (N_3099,In_2385,In_1891);
and U3100 (N_3100,In_2118,In_2349);
or U3101 (N_3101,In_2046,In_2274);
nand U3102 (N_3102,In_2229,In_86);
nor U3103 (N_3103,In_281,In_1530);
or U3104 (N_3104,In_1056,In_1786);
nor U3105 (N_3105,In_1141,In_2324);
nand U3106 (N_3106,In_516,In_1922);
and U3107 (N_3107,In_2108,In_1514);
and U3108 (N_3108,In_686,In_846);
nor U3109 (N_3109,In_826,In_8);
xor U3110 (N_3110,In_482,In_263);
or U3111 (N_3111,In_1029,In_1939);
nand U3112 (N_3112,In_281,In_2394);
nor U3113 (N_3113,In_2388,In_128);
or U3114 (N_3114,In_852,In_1885);
nand U3115 (N_3115,In_2222,In_1594);
xnor U3116 (N_3116,In_1026,In_1547);
or U3117 (N_3117,In_558,In_1465);
or U3118 (N_3118,In_1412,In_237);
and U3119 (N_3119,In_2100,In_1060);
and U3120 (N_3120,In_512,In_2131);
nand U3121 (N_3121,In_780,In_1329);
and U3122 (N_3122,In_763,In_1076);
xor U3123 (N_3123,In_494,In_945);
xnor U3124 (N_3124,In_2368,In_20);
nand U3125 (N_3125,In_1674,In_504);
and U3126 (N_3126,In_1377,In_1077);
or U3127 (N_3127,In_2144,In_1376);
or U3128 (N_3128,In_959,In_2408);
xnor U3129 (N_3129,In_112,In_1087);
and U3130 (N_3130,In_1125,In_1274);
and U3131 (N_3131,In_2386,In_1403);
xnor U3132 (N_3132,In_767,In_177);
nor U3133 (N_3133,In_508,In_1928);
xor U3134 (N_3134,In_893,In_2145);
nor U3135 (N_3135,In_1452,In_1010);
and U3136 (N_3136,In_1776,In_1619);
and U3137 (N_3137,In_28,In_2313);
nand U3138 (N_3138,In_1890,In_219);
nand U3139 (N_3139,In_845,In_274);
or U3140 (N_3140,In_2253,In_2462);
and U3141 (N_3141,In_2398,In_927);
nor U3142 (N_3142,In_366,In_259);
nor U3143 (N_3143,In_1671,In_2498);
and U3144 (N_3144,In_1230,In_2048);
nand U3145 (N_3145,In_1173,In_1785);
nor U3146 (N_3146,In_723,In_768);
xor U3147 (N_3147,In_2439,In_2320);
and U3148 (N_3148,In_1587,In_2130);
and U3149 (N_3149,In_672,In_1270);
and U3150 (N_3150,In_654,In_2259);
xor U3151 (N_3151,In_245,In_1062);
nand U3152 (N_3152,In_2466,In_760);
and U3153 (N_3153,In_1070,In_186);
xor U3154 (N_3154,In_738,In_279);
nand U3155 (N_3155,In_886,In_454);
nor U3156 (N_3156,In_1473,In_1845);
xnor U3157 (N_3157,In_161,In_1494);
nor U3158 (N_3158,In_2338,In_1438);
and U3159 (N_3159,In_2239,In_975);
nand U3160 (N_3160,In_1077,In_1603);
xor U3161 (N_3161,In_780,In_1596);
and U3162 (N_3162,In_1714,In_865);
or U3163 (N_3163,In_1563,In_1002);
or U3164 (N_3164,In_860,In_2137);
or U3165 (N_3165,In_2346,In_1254);
or U3166 (N_3166,In_2483,In_554);
nand U3167 (N_3167,In_1474,In_1277);
or U3168 (N_3168,In_65,In_167);
or U3169 (N_3169,In_2152,In_1776);
nor U3170 (N_3170,In_2199,In_2499);
and U3171 (N_3171,In_1475,In_2329);
and U3172 (N_3172,In_2149,In_1605);
nor U3173 (N_3173,In_2235,In_717);
xor U3174 (N_3174,In_318,In_1830);
nand U3175 (N_3175,In_2351,In_1493);
xor U3176 (N_3176,In_134,In_220);
or U3177 (N_3177,In_751,In_1997);
or U3178 (N_3178,In_1593,In_369);
or U3179 (N_3179,In_353,In_961);
or U3180 (N_3180,In_1899,In_850);
nand U3181 (N_3181,In_1732,In_1821);
or U3182 (N_3182,In_921,In_881);
nand U3183 (N_3183,In_1970,In_1044);
and U3184 (N_3184,In_1852,In_917);
or U3185 (N_3185,In_1337,In_1715);
nor U3186 (N_3186,In_1710,In_204);
nor U3187 (N_3187,In_448,In_1945);
nor U3188 (N_3188,In_78,In_79);
or U3189 (N_3189,In_2134,In_128);
xor U3190 (N_3190,In_1803,In_1646);
and U3191 (N_3191,In_648,In_798);
xnor U3192 (N_3192,In_2036,In_1484);
nand U3193 (N_3193,In_1877,In_421);
nor U3194 (N_3194,In_1059,In_487);
nand U3195 (N_3195,In_763,In_2355);
xnor U3196 (N_3196,In_146,In_760);
and U3197 (N_3197,In_1435,In_414);
nor U3198 (N_3198,In_1449,In_1125);
nor U3199 (N_3199,In_790,In_222);
xnor U3200 (N_3200,In_832,In_284);
nor U3201 (N_3201,In_1357,In_610);
nor U3202 (N_3202,In_1659,In_206);
and U3203 (N_3203,In_289,In_2326);
and U3204 (N_3204,In_569,In_371);
and U3205 (N_3205,In_2358,In_855);
and U3206 (N_3206,In_89,In_1997);
nand U3207 (N_3207,In_2052,In_696);
or U3208 (N_3208,In_618,In_521);
nor U3209 (N_3209,In_475,In_480);
and U3210 (N_3210,In_1305,In_248);
and U3211 (N_3211,In_1918,In_1303);
and U3212 (N_3212,In_1583,In_2425);
nand U3213 (N_3213,In_1257,In_625);
and U3214 (N_3214,In_1865,In_828);
and U3215 (N_3215,In_745,In_354);
and U3216 (N_3216,In_1140,In_2035);
nand U3217 (N_3217,In_480,In_0);
and U3218 (N_3218,In_138,In_502);
or U3219 (N_3219,In_527,In_1137);
and U3220 (N_3220,In_665,In_822);
xor U3221 (N_3221,In_1588,In_621);
nand U3222 (N_3222,In_2073,In_2235);
and U3223 (N_3223,In_204,In_1111);
nor U3224 (N_3224,In_830,In_969);
nor U3225 (N_3225,In_2346,In_1308);
or U3226 (N_3226,In_1028,In_1959);
nor U3227 (N_3227,In_233,In_2276);
nor U3228 (N_3228,In_1969,In_383);
and U3229 (N_3229,In_428,In_969);
nand U3230 (N_3230,In_1869,In_411);
nor U3231 (N_3231,In_1514,In_2469);
nor U3232 (N_3232,In_1445,In_983);
nor U3233 (N_3233,In_126,In_2056);
and U3234 (N_3234,In_1943,In_2053);
nor U3235 (N_3235,In_1582,In_261);
and U3236 (N_3236,In_1818,In_2102);
nand U3237 (N_3237,In_2481,In_513);
nand U3238 (N_3238,In_2211,In_1217);
or U3239 (N_3239,In_395,In_2320);
and U3240 (N_3240,In_1414,In_2024);
nor U3241 (N_3241,In_2247,In_2327);
xnor U3242 (N_3242,In_794,In_1677);
or U3243 (N_3243,In_2279,In_1978);
and U3244 (N_3244,In_779,In_2069);
nor U3245 (N_3245,In_601,In_226);
nand U3246 (N_3246,In_2244,In_1158);
or U3247 (N_3247,In_935,In_919);
nor U3248 (N_3248,In_1530,In_501);
or U3249 (N_3249,In_1675,In_1137);
or U3250 (N_3250,In_1261,In_46);
and U3251 (N_3251,In_272,In_1480);
xnor U3252 (N_3252,In_774,In_1334);
xnor U3253 (N_3253,In_1516,In_820);
nor U3254 (N_3254,In_16,In_1372);
xnor U3255 (N_3255,In_96,In_1581);
xor U3256 (N_3256,In_1938,In_2150);
or U3257 (N_3257,In_1084,In_367);
nand U3258 (N_3258,In_373,In_1153);
or U3259 (N_3259,In_2208,In_2321);
or U3260 (N_3260,In_1288,In_553);
nor U3261 (N_3261,In_435,In_1443);
nor U3262 (N_3262,In_676,In_1255);
or U3263 (N_3263,In_726,In_2450);
or U3264 (N_3264,In_1331,In_1308);
and U3265 (N_3265,In_678,In_1526);
nand U3266 (N_3266,In_370,In_1708);
and U3267 (N_3267,In_1657,In_659);
and U3268 (N_3268,In_664,In_38);
and U3269 (N_3269,In_1901,In_935);
nor U3270 (N_3270,In_838,In_1255);
xor U3271 (N_3271,In_1081,In_2066);
and U3272 (N_3272,In_1673,In_292);
xor U3273 (N_3273,In_1336,In_2439);
or U3274 (N_3274,In_1826,In_1057);
and U3275 (N_3275,In_2130,In_777);
or U3276 (N_3276,In_1898,In_505);
xor U3277 (N_3277,In_722,In_1611);
or U3278 (N_3278,In_913,In_2296);
and U3279 (N_3279,In_813,In_330);
xor U3280 (N_3280,In_1805,In_998);
nor U3281 (N_3281,In_328,In_306);
nand U3282 (N_3282,In_660,In_1711);
or U3283 (N_3283,In_938,In_761);
and U3284 (N_3284,In_2059,In_940);
or U3285 (N_3285,In_1514,In_5);
or U3286 (N_3286,In_1497,In_961);
nand U3287 (N_3287,In_1143,In_2049);
nor U3288 (N_3288,In_354,In_1099);
and U3289 (N_3289,In_1716,In_538);
and U3290 (N_3290,In_267,In_114);
or U3291 (N_3291,In_1184,In_1685);
and U3292 (N_3292,In_1140,In_1221);
nor U3293 (N_3293,In_1118,In_263);
nor U3294 (N_3294,In_1815,In_2448);
nor U3295 (N_3295,In_2352,In_1358);
nand U3296 (N_3296,In_1108,In_1393);
or U3297 (N_3297,In_294,In_2488);
xnor U3298 (N_3298,In_622,In_1350);
and U3299 (N_3299,In_2122,In_2443);
xor U3300 (N_3300,In_1844,In_2148);
or U3301 (N_3301,In_2195,In_1508);
nand U3302 (N_3302,In_874,In_1486);
or U3303 (N_3303,In_285,In_1597);
nand U3304 (N_3304,In_2369,In_918);
and U3305 (N_3305,In_811,In_801);
and U3306 (N_3306,In_2448,In_2076);
or U3307 (N_3307,In_878,In_40);
xor U3308 (N_3308,In_2087,In_2497);
xnor U3309 (N_3309,In_1112,In_863);
xnor U3310 (N_3310,In_602,In_2);
nand U3311 (N_3311,In_564,In_1216);
nand U3312 (N_3312,In_1747,In_2257);
or U3313 (N_3313,In_403,In_12);
and U3314 (N_3314,In_2294,In_2262);
nor U3315 (N_3315,In_2263,In_310);
nor U3316 (N_3316,In_1984,In_1349);
nand U3317 (N_3317,In_1944,In_1417);
and U3318 (N_3318,In_1815,In_693);
nor U3319 (N_3319,In_1739,In_1734);
nand U3320 (N_3320,In_1759,In_2455);
nor U3321 (N_3321,In_2070,In_305);
nand U3322 (N_3322,In_485,In_205);
and U3323 (N_3323,In_1758,In_1493);
nand U3324 (N_3324,In_640,In_1691);
nand U3325 (N_3325,In_1890,In_2460);
xor U3326 (N_3326,In_1636,In_267);
and U3327 (N_3327,In_763,In_336);
or U3328 (N_3328,In_103,In_2260);
or U3329 (N_3329,In_1749,In_2336);
and U3330 (N_3330,In_2064,In_165);
nor U3331 (N_3331,In_284,In_1806);
or U3332 (N_3332,In_2237,In_1221);
nor U3333 (N_3333,In_1907,In_1600);
xor U3334 (N_3334,In_202,In_1695);
or U3335 (N_3335,In_829,In_2034);
nand U3336 (N_3336,In_504,In_2439);
xnor U3337 (N_3337,In_401,In_914);
nand U3338 (N_3338,In_1180,In_779);
and U3339 (N_3339,In_1546,In_437);
or U3340 (N_3340,In_835,In_408);
nor U3341 (N_3341,In_933,In_1057);
xnor U3342 (N_3342,In_2150,In_886);
xor U3343 (N_3343,In_76,In_1071);
xnor U3344 (N_3344,In_1262,In_199);
nand U3345 (N_3345,In_2259,In_1293);
and U3346 (N_3346,In_2212,In_547);
nor U3347 (N_3347,In_265,In_1160);
nand U3348 (N_3348,In_1261,In_2319);
xnor U3349 (N_3349,In_16,In_903);
xnor U3350 (N_3350,In_1637,In_137);
nor U3351 (N_3351,In_1313,In_2087);
or U3352 (N_3352,In_34,In_2378);
nor U3353 (N_3353,In_2000,In_127);
nor U3354 (N_3354,In_1254,In_2436);
or U3355 (N_3355,In_1894,In_89);
and U3356 (N_3356,In_1082,In_1425);
nor U3357 (N_3357,In_482,In_925);
nor U3358 (N_3358,In_543,In_1226);
and U3359 (N_3359,In_2023,In_176);
xnor U3360 (N_3360,In_366,In_1368);
or U3361 (N_3361,In_285,In_1516);
and U3362 (N_3362,In_986,In_510);
and U3363 (N_3363,In_225,In_1408);
xnor U3364 (N_3364,In_2392,In_2406);
xor U3365 (N_3365,In_322,In_307);
or U3366 (N_3366,In_967,In_819);
and U3367 (N_3367,In_1471,In_1225);
or U3368 (N_3368,In_1025,In_2375);
or U3369 (N_3369,In_2314,In_755);
xor U3370 (N_3370,In_1964,In_1923);
nand U3371 (N_3371,In_1594,In_1798);
nor U3372 (N_3372,In_1198,In_1893);
xnor U3373 (N_3373,In_1297,In_1107);
nand U3374 (N_3374,In_2009,In_2121);
and U3375 (N_3375,In_373,In_1805);
xnor U3376 (N_3376,In_1822,In_280);
nand U3377 (N_3377,In_522,In_1241);
xor U3378 (N_3378,In_1520,In_599);
nand U3379 (N_3379,In_963,In_303);
and U3380 (N_3380,In_858,In_892);
or U3381 (N_3381,In_556,In_1707);
and U3382 (N_3382,In_2096,In_2455);
and U3383 (N_3383,In_1166,In_2252);
and U3384 (N_3384,In_814,In_1660);
nor U3385 (N_3385,In_651,In_561);
and U3386 (N_3386,In_2384,In_215);
or U3387 (N_3387,In_445,In_1603);
nand U3388 (N_3388,In_1756,In_874);
xnor U3389 (N_3389,In_1790,In_2310);
nand U3390 (N_3390,In_631,In_137);
nor U3391 (N_3391,In_1229,In_1922);
nand U3392 (N_3392,In_40,In_2250);
nor U3393 (N_3393,In_2301,In_1899);
nand U3394 (N_3394,In_1492,In_1859);
nor U3395 (N_3395,In_1111,In_1024);
nor U3396 (N_3396,In_2386,In_497);
nand U3397 (N_3397,In_1069,In_282);
nor U3398 (N_3398,In_1236,In_2168);
and U3399 (N_3399,In_1734,In_661);
or U3400 (N_3400,In_117,In_1737);
xnor U3401 (N_3401,In_632,In_73);
nor U3402 (N_3402,In_14,In_858);
nand U3403 (N_3403,In_921,In_1640);
nand U3404 (N_3404,In_2440,In_1008);
xor U3405 (N_3405,In_2218,In_1268);
or U3406 (N_3406,In_465,In_150);
or U3407 (N_3407,In_2492,In_1163);
and U3408 (N_3408,In_1109,In_633);
nand U3409 (N_3409,In_2184,In_306);
or U3410 (N_3410,In_423,In_1525);
nand U3411 (N_3411,In_2054,In_1312);
or U3412 (N_3412,In_301,In_1825);
nand U3413 (N_3413,In_238,In_1774);
or U3414 (N_3414,In_1961,In_310);
or U3415 (N_3415,In_364,In_1589);
or U3416 (N_3416,In_1201,In_488);
nor U3417 (N_3417,In_1302,In_142);
nor U3418 (N_3418,In_317,In_1786);
xnor U3419 (N_3419,In_2379,In_791);
nand U3420 (N_3420,In_1656,In_1455);
nand U3421 (N_3421,In_2332,In_1819);
or U3422 (N_3422,In_451,In_1645);
nand U3423 (N_3423,In_779,In_264);
or U3424 (N_3424,In_361,In_1722);
xnor U3425 (N_3425,In_606,In_2068);
or U3426 (N_3426,In_1066,In_615);
or U3427 (N_3427,In_432,In_1213);
xor U3428 (N_3428,In_1603,In_664);
or U3429 (N_3429,In_1470,In_82);
or U3430 (N_3430,In_2220,In_368);
nor U3431 (N_3431,In_439,In_1236);
or U3432 (N_3432,In_781,In_298);
nand U3433 (N_3433,In_545,In_115);
nor U3434 (N_3434,In_2387,In_1800);
xor U3435 (N_3435,In_1372,In_1096);
nand U3436 (N_3436,In_604,In_352);
nand U3437 (N_3437,In_1962,In_74);
nand U3438 (N_3438,In_1980,In_2498);
nand U3439 (N_3439,In_436,In_2264);
nor U3440 (N_3440,In_1613,In_2183);
or U3441 (N_3441,In_606,In_1822);
or U3442 (N_3442,In_1936,In_264);
nor U3443 (N_3443,In_2270,In_1915);
xnor U3444 (N_3444,In_94,In_263);
nand U3445 (N_3445,In_909,In_2320);
nor U3446 (N_3446,In_1210,In_897);
nand U3447 (N_3447,In_1475,In_942);
xor U3448 (N_3448,In_2113,In_1892);
or U3449 (N_3449,In_281,In_1597);
or U3450 (N_3450,In_2042,In_1754);
or U3451 (N_3451,In_88,In_2483);
xnor U3452 (N_3452,In_501,In_23);
xor U3453 (N_3453,In_2118,In_1756);
and U3454 (N_3454,In_2094,In_1368);
xor U3455 (N_3455,In_632,In_327);
and U3456 (N_3456,In_1883,In_1867);
nor U3457 (N_3457,In_1513,In_1610);
nand U3458 (N_3458,In_888,In_824);
nor U3459 (N_3459,In_2061,In_1670);
nor U3460 (N_3460,In_1886,In_1127);
and U3461 (N_3461,In_1552,In_513);
nand U3462 (N_3462,In_130,In_630);
nor U3463 (N_3463,In_2340,In_2350);
or U3464 (N_3464,In_2449,In_40);
nor U3465 (N_3465,In_496,In_1066);
nor U3466 (N_3466,In_2249,In_2162);
xnor U3467 (N_3467,In_1386,In_44);
or U3468 (N_3468,In_1977,In_2464);
and U3469 (N_3469,In_523,In_2353);
xor U3470 (N_3470,In_504,In_1588);
nor U3471 (N_3471,In_1546,In_1427);
or U3472 (N_3472,In_2114,In_1789);
or U3473 (N_3473,In_915,In_331);
xnor U3474 (N_3474,In_2201,In_889);
nor U3475 (N_3475,In_989,In_1559);
xnor U3476 (N_3476,In_1084,In_2183);
or U3477 (N_3477,In_2067,In_1087);
nand U3478 (N_3478,In_606,In_2003);
xor U3479 (N_3479,In_2206,In_1067);
and U3480 (N_3480,In_1594,In_431);
and U3481 (N_3481,In_883,In_1651);
and U3482 (N_3482,In_2390,In_1197);
nand U3483 (N_3483,In_756,In_2179);
xnor U3484 (N_3484,In_505,In_288);
nand U3485 (N_3485,In_11,In_1311);
nor U3486 (N_3486,In_643,In_160);
nor U3487 (N_3487,In_1531,In_1200);
nor U3488 (N_3488,In_259,In_2220);
or U3489 (N_3489,In_397,In_2272);
and U3490 (N_3490,In_117,In_1083);
xor U3491 (N_3491,In_2248,In_1467);
nor U3492 (N_3492,In_591,In_37);
or U3493 (N_3493,In_1419,In_1249);
xnor U3494 (N_3494,In_968,In_1487);
nor U3495 (N_3495,In_2200,In_162);
or U3496 (N_3496,In_1506,In_1807);
and U3497 (N_3497,In_1739,In_212);
xnor U3498 (N_3498,In_1293,In_2109);
nor U3499 (N_3499,In_182,In_2325);
xor U3500 (N_3500,In_2076,In_669);
xor U3501 (N_3501,In_2429,In_2113);
and U3502 (N_3502,In_330,In_770);
or U3503 (N_3503,In_862,In_962);
nor U3504 (N_3504,In_1179,In_1084);
or U3505 (N_3505,In_835,In_2490);
nor U3506 (N_3506,In_964,In_2373);
or U3507 (N_3507,In_2242,In_226);
and U3508 (N_3508,In_64,In_2086);
nand U3509 (N_3509,In_442,In_216);
nor U3510 (N_3510,In_540,In_1419);
or U3511 (N_3511,In_1937,In_2181);
or U3512 (N_3512,In_1624,In_233);
xor U3513 (N_3513,In_1644,In_130);
or U3514 (N_3514,In_1456,In_1358);
nand U3515 (N_3515,In_865,In_279);
nand U3516 (N_3516,In_858,In_842);
nor U3517 (N_3517,In_20,In_1585);
nor U3518 (N_3518,In_1976,In_585);
xor U3519 (N_3519,In_1125,In_2041);
nor U3520 (N_3520,In_504,In_754);
and U3521 (N_3521,In_2378,In_2026);
xnor U3522 (N_3522,In_2490,In_657);
and U3523 (N_3523,In_2185,In_2273);
nor U3524 (N_3524,In_27,In_744);
nor U3525 (N_3525,In_1786,In_1465);
and U3526 (N_3526,In_1092,In_936);
nand U3527 (N_3527,In_2102,In_644);
or U3528 (N_3528,In_1665,In_1807);
nand U3529 (N_3529,In_1199,In_1542);
xor U3530 (N_3530,In_1995,In_914);
nand U3531 (N_3531,In_1529,In_1544);
or U3532 (N_3532,In_442,In_2396);
nand U3533 (N_3533,In_6,In_490);
nor U3534 (N_3534,In_1598,In_686);
xnor U3535 (N_3535,In_563,In_1245);
xnor U3536 (N_3536,In_395,In_1577);
nand U3537 (N_3537,In_1654,In_449);
nor U3538 (N_3538,In_258,In_290);
and U3539 (N_3539,In_1341,In_2310);
xor U3540 (N_3540,In_184,In_1061);
xnor U3541 (N_3541,In_472,In_1219);
and U3542 (N_3542,In_951,In_1959);
or U3543 (N_3543,In_30,In_1799);
nand U3544 (N_3544,In_1174,In_1147);
nand U3545 (N_3545,In_568,In_1188);
xnor U3546 (N_3546,In_1081,In_1027);
or U3547 (N_3547,In_1071,In_462);
and U3548 (N_3548,In_2021,In_735);
nand U3549 (N_3549,In_897,In_938);
or U3550 (N_3550,In_754,In_131);
nand U3551 (N_3551,In_1060,In_2438);
or U3552 (N_3552,In_2098,In_706);
or U3553 (N_3553,In_2036,In_1354);
nor U3554 (N_3554,In_38,In_397);
or U3555 (N_3555,In_25,In_618);
or U3556 (N_3556,In_75,In_39);
and U3557 (N_3557,In_1707,In_2442);
nor U3558 (N_3558,In_858,In_945);
and U3559 (N_3559,In_481,In_2318);
xnor U3560 (N_3560,In_627,In_1663);
and U3561 (N_3561,In_1498,In_376);
xnor U3562 (N_3562,In_732,In_1817);
nor U3563 (N_3563,In_215,In_2215);
xor U3564 (N_3564,In_2005,In_295);
and U3565 (N_3565,In_1159,In_2345);
nor U3566 (N_3566,In_1351,In_554);
nand U3567 (N_3567,In_1823,In_1503);
nand U3568 (N_3568,In_1629,In_1196);
nor U3569 (N_3569,In_690,In_1505);
nor U3570 (N_3570,In_846,In_423);
xor U3571 (N_3571,In_2455,In_1696);
xnor U3572 (N_3572,In_1465,In_781);
and U3573 (N_3573,In_1603,In_1888);
nor U3574 (N_3574,In_1921,In_659);
nor U3575 (N_3575,In_2365,In_2269);
xor U3576 (N_3576,In_2114,In_1587);
nor U3577 (N_3577,In_333,In_496);
xor U3578 (N_3578,In_1944,In_967);
and U3579 (N_3579,In_883,In_2366);
or U3580 (N_3580,In_1075,In_114);
xnor U3581 (N_3581,In_211,In_329);
nor U3582 (N_3582,In_524,In_2372);
and U3583 (N_3583,In_389,In_2074);
nand U3584 (N_3584,In_1084,In_442);
xnor U3585 (N_3585,In_1065,In_886);
xnor U3586 (N_3586,In_1881,In_1524);
xnor U3587 (N_3587,In_2006,In_1577);
or U3588 (N_3588,In_1952,In_2126);
and U3589 (N_3589,In_1671,In_1281);
nor U3590 (N_3590,In_180,In_2458);
xnor U3591 (N_3591,In_1419,In_1173);
xnor U3592 (N_3592,In_2014,In_1354);
xor U3593 (N_3593,In_982,In_1457);
xnor U3594 (N_3594,In_436,In_1184);
nor U3595 (N_3595,In_577,In_1966);
nor U3596 (N_3596,In_1404,In_330);
nor U3597 (N_3597,In_126,In_494);
and U3598 (N_3598,In_583,In_1384);
nor U3599 (N_3599,In_550,In_1473);
and U3600 (N_3600,In_2473,In_1115);
or U3601 (N_3601,In_1443,In_2393);
nor U3602 (N_3602,In_713,In_363);
nor U3603 (N_3603,In_2452,In_190);
or U3604 (N_3604,In_1305,In_518);
or U3605 (N_3605,In_1267,In_64);
xnor U3606 (N_3606,In_1818,In_1909);
and U3607 (N_3607,In_2385,In_700);
or U3608 (N_3608,In_655,In_1430);
nand U3609 (N_3609,In_471,In_496);
nor U3610 (N_3610,In_2271,In_724);
nand U3611 (N_3611,In_0,In_2307);
xnor U3612 (N_3612,In_2455,In_1628);
and U3613 (N_3613,In_2432,In_1421);
and U3614 (N_3614,In_598,In_2449);
or U3615 (N_3615,In_319,In_1766);
nor U3616 (N_3616,In_1546,In_1850);
and U3617 (N_3617,In_2393,In_1754);
or U3618 (N_3618,In_63,In_2171);
nor U3619 (N_3619,In_286,In_2295);
nand U3620 (N_3620,In_2352,In_1396);
and U3621 (N_3621,In_373,In_1182);
and U3622 (N_3622,In_832,In_1094);
nand U3623 (N_3623,In_1964,In_913);
and U3624 (N_3624,In_1051,In_1146);
and U3625 (N_3625,In_2164,In_2158);
xor U3626 (N_3626,In_852,In_1491);
xor U3627 (N_3627,In_477,In_216);
nor U3628 (N_3628,In_998,In_271);
and U3629 (N_3629,In_2283,In_200);
nor U3630 (N_3630,In_1450,In_189);
or U3631 (N_3631,In_188,In_2393);
and U3632 (N_3632,In_1661,In_1764);
xor U3633 (N_3633,In_2259,In_1030);
or U3634 (N_3634,In_1293,In_1905);
and U3635 (N_3635,In_2036,In_645);
nor U3636 (N_3636,In_2204,In_1599);
and U3637 (N_3637,In_1354,In_1042);
nand U3638 (N_3638,In_148,In_162);
or U3639 (N_3639,In_1294,In_574);
xor U3640 (N_3640,In_476,In_1975);
or U3641 (N_3641,In_286,In_2490);
and U3642 (N_3642,In_2408,In_2416);
xor U3643 (N_3643,In_1680,In_797);
nor U3644 (N_3644,In_407,In_1741);
nor U3645 (N_3645,In_450,In_2072);
nor U3646 (N_3646,In_1599,In_1633);
or U3647 (N_3647,In_1872,In_591);
nor U3648 (N_3648,In_2245,In_1384);
nand U3649 (N_3649,In_1394,In_1204);
nand U3650 (N_3650,In_2423,In_1142);
and U3651 (N_3651,In_1377,In_259);
nor U3652 (N_3652,In_1348,In_1120);
and U3653 (N_3653,In_1237,In_603);
xor U3654 (N_3654,In_46,In_1897);
or U3655 (N_3655,In_976,In_55);
or U3656 (N_3656,In_1599,In_691);
and U3657 (N_3657,In_419,In_2181);
xor U3658 (N_3658,In_1994,In_1473);
and U3659 (N_3659,In_482,In_205);
or U3660 (N_3660,In_1136,In_1452);
xnor U3661 (N_3661,In_2237,In_702);
xor U3662 (N_3662,In_1880,In_394);
nor U3663 (N_3663,In_979,In_1879);
nor U3664 (N_3664,In_14,In_2170);
xor U3665 (N_3665,In_164,In_959);
xor U3666 (N_3666,In_460,In_1854);
nor U3667 (N_3667,In_1700,In_135);
nand U3668 (N_3668,In_961,In_1431);
xor U3669 (N_3669,In_34,In_2046);
nor U3670 (N_3670,In_1130,In_131);
nand U3671 (N_3671,In_1952,In_2008);
or U3672 (N_3672,In_2119,In_1337);
xor U3673 (N_3673,In_325,In_1091);
or U3674 (N_3674,In_435,In_1);
xnor U3675 (N_3675,In_1565,In_477);
and U3676 (N_3676,In_1987,In_1574);
nand U3677 (N_3677,In_1613,In_1039);
xor U3678 (N_3678,In_2273,In_1693);
nand U3679 (N_3679,In_1644,In_2240);
nor U3680 (N_3680,In_901,In_1042);
and U3681 (N_3681,In_1038,In_781);
nand U3682 (N_3682,In_432,In_2475);
and U3683 (N_3683,In_1011,In_1507);
and U3684 (N_3684,In_1044,In_2268);
or U3685 (N_3685,In_113,In_1196);
and U3686 (N_3686,In_1667,In_952);
nor U3687 (N_3687,In_1564,In_513);
xnor U3688 (N_3688,In_2328,In_1547);
or U3689 (N_3689,In_2100,In_1222);
nor U3690 (N_3690,In_303,In_361);
nor U3691 (N_3691,In_1047,In_945);
and U3692 (N_3692,In_301,In_150);
or U3693 (N_3693,In_1809,In_420);
nand U3694 (N_3694,In_431,In_1129);
nand U3695 (N_3695,In_376,In_597);
nand U3696 (N_3696,In_974,In_1915);
nand U3697 (N_3697,In_1549,In_829);
and U3698 (N_3698,In_1064,In_2437);
or U3699 (N_3699,In_648,In_644);
and U3700 (N_3700,In_2006,In_629);
or U3701 (N_3701,In_1892,In_139);
xor U3702 (N_3702,In_2251,In_1185);
nor U3703 (N_3703,In_1105,In_693);
and U3704 (N_3704,In_1254,In_1728);
or U3705 (N_3705,In_492,In_466);
and U3706 (N_3706,In_1106,In_2470);
and U3707 (N_3707,In_2380,In_462);
or U3708 (N_3708,In_1064,In_448);
and U3709 (N_3709,In_1188,In_1566);
xor U3710 (N_3710,In_1570,In_920);
or U3711 (N_3711,In_204,In_692);
xnor U3712 (N_3712,In_1619,In_723);
nand U3713 (N_3713,In_1677,In_711);
xor U3714 (N_3714,In_360,In_569);
nor U3715 (N_3715,In_1050,In_2163);
nand U3716 (N_3716,In_2061,In_1130);
and U3717 (N_3717,In_400,In_408);
and U3718 (N_3718,In_2488,In_2053);
nand U3719 (N_3719,In_108,In_1761);
nand U3720 (N_3720,In_667,In_2146);
and U3721 (N_3721,In_26,In_352);
and U3722 (N_3722,In_857,In_166);
nand U3723 (N_3723,In_2355,In_2093);
nand U3724 (N_3724,In_2293,In_2429);
nand U3725 (N_3725,In_783,In_1667);
xnor U3726 (N_3726,In_36,In_305);
nor U3727 (N_3727,In_708,In_767);
xor U3728 (N_3728,In_2050,In_500);
xnor U3729 (N_3729,In_914,In_1803);
nand U3730 (N_3730,In_1539,In_2368);
nor U3731 (N_3731,In_2479,In_456);
and U3732 (N_3732,In_32,In_2108);
nand U3733 (N_3733,In_2391,In_65);
or U3734 (N_3734,In_1730,In_77);
nor U3735 (N_3735,In_1631,In_1328);
or U3736 (N_3736,In_994,In_128);
and U3737 (N_3737,In_455,In_1233);
nand U3738 (N_3738,In_653,In_560);
xnor U3739 (N_3739,In_1138,In_410);
nor U3740 (N_3740,In_69,In_660);
nor U3741 (N_3741,In_2100,In_778);
xnor U3742 (N_3742,In_817,In_1355);
nor U3743 (N_3743,In_1183,In_2331);
nand U3744 (N_3744,In_823,In_196);
xnor U3745 (N_3745,In_450,In_1726);
xor U3746 (N_3746,In_1710,In_400);
xor U3747 (N_3747,In_1409,In_2225);
or U3748 (N_3748,In_546,In_491);
or U3749 (N_3749,In_138,In_1891);
and U3750 (N_3750,In_1945,In_1075);
nor U3751 (N_3751,In_41,In_1148);
xnor U3752 (N_3752,In_826,In_889);
xnor U3753 (N_3753,In_2003,In_501);
nand U3754 (N_3754,In_1633,In_811);
xnor U3755 (N_3755,In_1895,In_2361);
or U3756 (N_3756,In_864,In_1937);
nand U3757 (N_3757,In_148,In_133);
xor U3758 (N_3758,In_2292,In_448);
nor U3759 (N_3759,In_735,In_1767);
or U3760 (N_3760,In_1280,In_430);
nor U3761 (N_3761,In_2159,In_157);
nand U3762 (N_3762,In_2148,In_1804);
and U3763 (N_3763,In_904,In_2107);
and U3764 (N_3764,In_528,In_1331);
or U3765 (N_3765,In_2251,In_1906);
nand U3766 (N_3766,In_916,In_2471);
nand U3767 (N_3767,In_1182,In_845);
or U3768 (N_3768,In_1179,In_1789);
and U3769 (N_3769,In_887,In_2080);
xor U3770 (N_3770,In_1680,In_2264);
xor U3771 (N_3771,In_2252,In_512);
xnor U3772 (N_3772,In_562,In_2087);
xnor U3773 (N_3773,In_2068,In_1484);
and U3774 (N_3774,In_1954,In_2426);
nor U3775 (N_3775,In_2480,In_1836);
nand U3776 (N_3776,In_481,In_1990);
nor U3777 (N_3777,In_1630,In_2172);
and U3778 (N_3778,In_705,In_1734);
or U3779 (N_3779,In_425,In_7);
or U3780 (N_3780,In_1936,In_375);
nor U3781 (N_3781,In_100,In_1045);
xnor U3782 (N_3782,In_954,In_1414);
nor U3783 (N_3783,In_1923,In_1494);
nor U3784 (N_3784,In_2274,In_1840);
nor U3785 (N_3785,In_1934,In_1208);
nand U3786 (N_3786,In_764,In_296);
and U3787 (N_3787,In_1336,In_1112);
and U3788 (N_3788,In_2032,In_2178);
nor U3789 (N_3789,In_1395,In_1937);
nand U3790 (N_3790,In_718,In_32);
and U3791 (N_3791,In_79,In_1629);
nor U3792 (N_3792,In_133,In_2016);
nand U3793 (N_3793,In_1933,In_571);
or U3794 (N_3794,In_803,In_2405);
or U3795 (N_3795,In_1869,In_1120);
xnor U3796 (N_3796,In_601,In_707);
nand U3797 (N_3797,In_1046,In_2283);
xnor U3798 (N_3798,In_1564,In_1735);
or U3799 (N_3799,In_808,In_646);
nor U3800 (N_3800,In_1558,In_843);
nor U3801 (N_3801,In_379,In_795);
xnor U3802 (N_3802,In_998,In_1266);
nand U3803 (N_3803,In_186,In_301);
nor U3804 (N_3804,In_781,In_156);
or U3805 (N_3805,In_907,In_1946);
and U3806 (N_3806,In_441,In_2058);
nor U3807 (N_3807,In_1272,In_434);
or U3808 (N_3808,In_1201,In_1700);
nor U3809 (N_3809,In_1407,In_1948);
nand U3810 (N_3810,In_2429,In_1972);
nand U3811 (N_3811,In_469,In_1232);
xnor U3812 (N_3812,In_1994,In_753);
xor U3813 (N_3813,In_1645,In_259);
xor U3814 (N_3814,In_81,In_179);
nor U3815 (N_3815,In_1530,In_1320);
and U3816 (N_3816,In_1066,In_1052);
xor U3817 (N_3817,In_1480,In_2264);
or U3818 (N_3818,In_1587,In_1500);
nor U3819 (N_3819,In_1639,In_2339);
nor U3820 (N_3820,In_984,In_1712);
and U3821 (N_3821,In_617,In_1097);
and U3822 (N_3822,In_1200,In_1762);
xnor U3823 (N_3823,In_2206,In_1137);
or U3824 (N_3824,In_2017,In_361);
xor U3825 (N_3825,In_1178,In_1054);
or U3826 (N_3826,In_2123,In_1265);
and U3827 (N_3827,In_1231,In_1458);
or U3828 (N_3828,In_2311,In_595);
xor U3829 (N_3829,In_1057,In_951);
or U3830 (N_3830,In_1555,In_2363);
and U3831 (N_3831,In_424,In_1298);
xnor U3832 (N_3832,In_2300,In_2422);
and U3833 (N_3833,In_360,In_971);
nand U3834 (N_3834,In_8,In_1803);
and U3835 (N_3835,In_855,In_1446);
xor U3836 (N_3836,In_1591,In_44);
nand U3837 (N_3837,In_60,In_1169);
and U3838 (N_3838,In_1463,In_397);
or U3839 (N_3839,In_246,In_729);
and U3840 (N_3840,In_836,In_145);
nor U3841 (N_3841,In_1379,In_958);
nand U3842 (N_3842,In_1254,In_2267);
nor U3843 (N_3843,In_1201,In_2456);
xnor U3844 (N_3844,In_449,In_750);
and U3845 (N_3845,In_1836,In_1742);
nor U3846 (N_3846,In_685,In_1451);
and U3847 (N_3847,In_164,In_1983);
nand U3848 (N_3848,In_1079,In_1546);
and U3849 (N_3849,In_213,In_1997);
and U3850 (N_3850,In_139,In_2173);
nor U3851 (N_3851,In_1803,In_782);
nand U3852 (N_3852,In_846,In_1025);
xor U3853 (N_3853,In_196,In_793);
nor U3854 (N_3854,In_1273,In_1902);
xor U3855 (N_3855,In_455,In_746);
xor U3856 (N_3856,In_364,In_2373);
nand U3857 (N_3857,In_1937,In_2322);
xor U3858 (N_3858,In_1100,In_388);
and U3859 (N_3859,In_1858,In_1378);
nor U3860 (N_3860,In_842,In_2024);
xor U3861 (N_3861,In_1269,In_1330);
and U3862 (N_3862,In_2189,In_1938);
xor U3863 (N_3863,In_732,In_2497);
nor U3864 (N_3864,In_252,In_373);
xor U3865 (N_3865,In_1870,In_1919);
nand U3866 (N_3866,In_2293,In_2071);
and U3867 (N_3867,In_657,In_1910);
and U3868 (N_3868,In_789,In_1095);
and U3869 (N_3869,In_1427,In_225);
or U3870 (N_3870,In_31,In_2263);
nand U3871 (N_3871,In_1443,In_431);
or U3872 (N_3872,In_2253,In_663);
or U3873 (N_3873,In_8,In_784);
or U3874 (N_3874,In_2061,In_1367);
or U3875 (N_3875,In_1698,In_1618);
or U3876 (N_3876,In_649,In_270);
nand U3877 (N_3877,In_383,In_2326);
nand U3878 (N_3878,In_1905,In_893);
nor U3879 (N_3879,In_2273,In_1602);
and U3880 (N_3880,In_1678,In_1267);
nor U3881 (N_3881,In_1520,In_1281);
and U3882 (N_3882,In_1592,In_960);
nor U3883 (N_3883,In_2123,In_2071);
or U3884 (N_3884,In_542,In_477);
and U3885 (N_3885,In_338,In_1229);
nand U3886 (N_3886,In_1954,In_1117);
and U3887 (N_3887,In_1964,In_1911);
nor U3888 (N_3888,In_1784,In_1072);
xor U3889 (N_3889,In_1423,In_562);
xnor U3890 (N_3890,In_2155,In_1199);
nand U3891 (N_3891,In_2479,In_1618);
xor U3892 (N_3892,In_1267,In_1459);
or U3893 (N_3893,In_775,In_37);
and U3894 (N_3894,In_462,In_1714);
nor U3895 (N_3895,In_1913,In_1357);
and U3896 (N_3896,In_2291,In_1432);
and U3897 (N_3897,In_1079,In_1599);
and U3898 (N_3898,In_1864,In_421);
xnor U3899 (N_3899,In_2352,In_1592);
xnor U3900 (N_3900,In_1261,In_973);
nand U3901 (N_3901,In_2473,In_1634);
xor U3902 (N_3902,In_1153,In_2436);
or U3903 (N_3903,In_1098,In_2255);
nor U3904 (N_3904,In_1293,In_168);
xor U3905 (N_3905,In_2379,In_854);
or U3906 (N_3906,In_2355,In_705);
and U3907 (N_3907,In_2486,In_1704);
and U3908 (N_3908,In_2053,In_322);
xor U3909 (N_3909,In_332,In_1711);
xor U3910 (N_3910,In_1139,In_1637);
xor U3911 (N_3911,In_201,In_1442);
or U3912 (N_3912,In_1009,In_532);
and U3913 (N_3913,In_2301,In_851);
or U3914 (N_3914,In_1470,In_170);
nand U3915 (N_3915,In_966,In_2185);
nor U3916 (N_3916,In_1369,In_1487);
nor U3917 (N_3917,In_1469,In_1);
or U3918 (N_3918,In_2290,In_1642);
nor U3919 (N_3919,In_924,In_2168);
xor U3920 (N_3920,In_985,In_519);
nor U3921 (N_3921,In_1416,In_150);
and U3922 (N_3922,In_744,In_684);
xnor U3923 (N_3923,In_1484,In_828);
or U3924 (N_3924,In_601,In_1138);
nand U3925 (N_3925,In_108,In_2012);
and U3926 (N_3926,In_95,In_438);
or U3927 (N_3927,In_603,In_1627);
nor U3928 (N_3928,In_1084,In_1491);
xor U3929 (N_3929,In_343,In_472);
or U3930 (N_3930,In_1386,In_2164);
nor U3931 (N_3931,In_917,In_717);
nand U3932 (N_3932,In_1867,In_1600);
nor U3933 (N_3933,In_1938,In_2001);
xnor U3934 (N_3934,In_1099,In_826);
xnor U3935 (N_3935,In_677,In_1963);
and U3936 (N_3936,In_243,In_2008);
xnor U3937 (N_3937,In_1515,In_1171);
nor U3938 (N_3938,In_777,In_1635);
or U3939 (N_3939,In_1674,In_2076);
and U3940 (N_3940,In_1575,In_486);
xnor U3941 (N_3941,In_1282,In_1142);
and U3942 (N_3942,In_499,In_2370);
nor U3943 (N_3943,In_965,In_217);
xor U3944 (N_3944,In_369,In_674);
nor U3945 (N_3945,In_1708,In_164);
or U3946 (N_3946,In_14,In_808);
nor U3947 (N_3947,In_983,In_92);
nand U3948 (N_3948,In_2257,In_622);
nor U3949 (N_3949,In_2404,In_433);
xor U3950 (N_3950,In_1014,In_752);
or U3951 (N_3951,In_1769,In_201);
nand U3952 (N_3952,In_1087,In_353);
nor U3953 (N_3953,In_261,In_71);
nor U3954 (N_3954,In_1913,In_1186);
and U3955 (N_3955,In_357,In_1807);
nor U3956 (N_3956,In_505,In_1229);
or U3957 (N_3957,In_1936,In_2154);
nand U3958 (N_3958,In_2093,In_471);
nor U3959 (N_3959,In_145,In_1496);
or U3960 (N_3960,In_2232,In_137);
nand U3961 (N_3961,In_1240,In_636);
and U3962 (N_3962,In_1500,In_1959);
xor U3963 (N_3963,In_2155,In_2399);
nor U3964 (N_3964,In_560,In_635);
nor U3965 (N_3965,In_1840,In_1023);
nand U3966 (N_3966,In_622,In_547);
nor U3967 (N_3967,In_2031,In_2345);
nand U3968 (N_3968,In_691,In_812);
and U3969 (N_3969,In_1130,In_1410);
xnor U3970 (N_3970,In_476,In_2397);
nor U3971 (N_3971,In_32,In_2344);
nor U3972 (N_3972,In_2050,In_80);
nor U3973 (N_3973,In_1929,In_1115);
and U3974 (N_3974,In_1475,In_438);
or U3975 (N_3975,In_690,In_767);
or U3976 (N_3976,In_932,In_825);
and U3977 (N_3977,In_1966,In_676);
or U3978 (N_3978,In_479,In_2393);
or U3979 (N_3979,In_1181,In_1243);
xor U3980 (N_3980,In_444,In_1806);
or U3981 (N_3981,In_2428,In_1677);
or U3982 (N_3982,In_918,In_2087);
nand U3983 (N_3983,In_2250,In_2079);
and U3984 (N_3984,In_497,In_164);
nor U3985 (N_3985,In_497,In_375);
or U3986 (N_3986,In_1462,In_1079);
xnor U3987 (N_3987,In_1748,In_2265);
and U3988 (N_3988,In_349,In_2453);
nor U3989 (N_3989,In_2100,In_89);
and U3990 (N_3990,In_66,In_787);
nor U3991 (N_3991,In_1780,In_2497);
and U3992 (N_3992,In_205,In_2323);
and U3993 (N_3993,In_357,In_2087);
xnor U3994 (N_3994,In_2362,In_1170);
nand U3995 (N_3995,In_174,In_2159);
or U3996 (N_3996,In_1265,In_1353);
and U3997 (N_3997,In_34,In_629);
nand U3998 (N_3998,In_2489,In_1828);
and U3999 (N_3999,In_1424,In_2465);
nor U4000 (N_4000,In_2289,In_2477);
and U4001 (N_4001,In_1595,In_602);
nand U4002 (N_4002,In_1774,In_281);
and U4003 (N_4003,In_1333,In_819);
and U4004 (N_4004,In_453,In_1929);
and U4005 (N_4005,In_856,In_2170);
nand U4006 (N_4006,In_2239,In_1731);
nand U4007 (N_4007,In_1139,In_2088);
and U4008 (N_4008,In_265,In_1371);
nor U4009 (N_4009,In_2454,In_1052);
xnor U4010 (N_4010,In_212,In_1760);
or U4011 (N_4011,In_648,In_1853);
or U4012 (N_4012,In_2391,In_2030);
and U4013 (N_4013,In_557,In_158);
nor U4014 (N_4014,In_1330,In_314);
xor U4015 (N_4015,In_1920,In_2252);
and U4016 (N_4016,In_1688,In_2032);
or U4017 (N_4017,In_2114,In_1082);
xor U4018 (N_4018,In_1163,In_1369);
xnor U4019 (N_4019,In_150,In_767);
xor U4020 (N_4020,In_741,In_422);
nand U4021 (N_4021,In_681,In_27);
or U4022 (N_4022,In_125,In_2407);
and U4023 (N_4023,In_251,In_2469);
and U4024 (N_4024,In_1913,In_890);
or U4025 (N_4025,In_1537,In_89);
and U4026 (N_4026,In_1135,In_1073);
nor U4027 (N_4027,In_1559,In_205);
nand U4028 (N_4028,In_399,In_291);
nand U4029 (N_4029,In_2435,In_1035);
and U4030 (N_4030,In_889,In_619);
nor U4031 (N_4031,In_893,In_929);
xor U4032 (N_4032,In_857,In_2158);
nor U4033 (N_4033,In_2076,In_2001);
or U4034 (N_4034,In_330,In_9);
and U4035 (N_4035,In_1249,In_2391);
nand U4036 (N_4036,In_67,In_1838);
xor U4037 (N_4037,In_1037,In_111);
nor U4038 (N_4038,In_1902,In_523);
xnor U4039 (N_4039,In_2429,In_1444);
and U4040 (N_4040,In_2316,In_188);
or U4041 (N_4041,In_498,In_2358);
nand U4042 (N_4042,In_497,In_1240);
nand U4043 (N_4043,In_1053,In_158);
and U4044 (N_4044,In_1705,In_478);
nand U4045 (N_4045,In_2330,In_1457);
and U4046 (N_4046,In_171,In_1763);
nand U4047 (N_4047,In_1445,In_208);
and U4048 (N_4048,In_636,In_1593);
xnor U4049 (N_4049,In_1738,In_4);
or U4050 (N_4050,In_1406,In_939);
or U4051 (N_4051,In_479,In_781);
nor U4052 (N_4052,In_636,In_1850);
nor U4053 (N_4053,In_586,In_2110);
nand U4054 (N_4054,In_1039,In_1079);
and U4055 (N_4055,In_108,In_2486);
or U4056 (N_4056,In_75,In_460);
and U4057 (N_4057,In_1231,In_1900);
or U4058 (N_4058,In_1101,In_1031);
nand U4059 (N_4059,In_1057,In_2474);
nand U4060 (N_4060,In_243,In_1581);
nand U4061 (N_4061,In_1681,In_2430);
and U4062 (N_4062,In_380,In_1376);
nand U4063 (N_4063,In_1856,In_121);
or U4064 (N_4064,In_381,In_1397);
xnor U4065 (N_4065,In_1983,In_1414);
or U4066 (N_4066,In_152,In_2080);
nand U4067 (N_4067,In_1828,In_819);
nand U4068 (N_4068,In_1644,In_925);
and U4069 (N_4069,In_1241,In_487);
xnor U4070 (N_4070,In_2104,In_2316);
or U4071 (N_4071,In_2219,In_1897);
or U4072 (N_4072,In_1293,In_7);
and U4073 (N_4073,In_1667,In_1228);
or U4074 (N_4074,In_509,In_441);
nor U4075 (N_4075,In_912,In_1828);
nand U4076 (N_4076,In_454,In_2055);
and U4077 (N_4077,In_905,In_1991);
xnor U4078 (N_4078,In_1114,In_1252);
nor U4079 (N_4079,In_1004,In_635);
xor U4080 (N_4080,In_1742,In_1057);
or U4081 (N_4081,In_1735,In_2046);
and U4082 (N_4082,In_62,In_1758);
nor U4083 (N_4083,In_850,In_1449);
nand U4084 (N_4084,In_727,In_2146);
nor U4085 (N_4085,In_2411,In_356);
nor U4086 (N_4086,In_806,In_977);
or U4087 (N_4087,In_1825,In_177);
or U4088 (N_4088,In_2276,In_2032);
nand U4089 (N_4089,In_242,In_392);
or U4090 (N_4090,In_1591,In_1071);
nor U4091 (N_4091,In_1986,In_109);
nor U4092 (N_4092,In_1149,In_572);
nor U4093 (N_4093,In_1307,In_2);
xor U4094 (N_4094,In_2199,In_762);
or U4095 (N_4095,In_2008,In_1516);
nor U4096 (N_4096,In_225,In_2066);
nand U4097 (N_4097,In_997,In_1715);
and U4098 (N_4098,In_339,In_2138);
nand U4099 (N_4099,In_1006,In_2343);
or U4100 (N_4100,In_1004,In_256);
xor U4101 (N_4101,In_1857,In_646);
xor U4102 (N_4102,In_177,In_782);
xor U4103 (N_4103,In_1072,In_1881);
nor U4104 (N_4104,In_99,In_1009);
nor U4105 (N_4105,In_1043,In_907);
and U4106 (N_4106,In_272,In_582);
or U4107 (N_4107,In_1683,In_1015);
and U4108 (N_4108,In_437,In_2181);
or U4109 (N_4109,In_1269,In_512);
nor U4110 (N_4110,In_2098,In_2285);
nand U4111 (N_4111,In_1990,In_941);
nand U4112 (N_4112,In_2043,In_58);
nand U4113 (N_4113,In_869,In_2206);
xnor U4114 (N_4114,In_96,In_275);
or U4115 (N_4115,In_370,In_1897);
or U4116 (N_4116,In_296,In_1691);
nor U4117 (N_4117,In_1995,In_2328);
and U4118 (N_4118,In_1543,In_1937);
nor U4119 (N_4119,In_165,In_2454);
nor U4120 (N_4120,In_1285,In_2232);
xnor U4121 (N_4121,In_1678,In_266);
nand U4122 (N_4122,In_1854,In_1252);
xor U4123 (N_4123,In_175,In_488);
or U4124 (N_4124,In_1150,In_741);
or U4125 (N_4125,In_1835,In_997);
xnor U4126 (N_4126,In_1746,In_173);
xnor U4127 (N_4127,In_2056,In_782);
and U4128 (N_4128,In_778,In_1156);
nor U4129 (N_4129,In_1549,In_449);
or U4130 (N_4130,In_2369,In_890);
xnor U4131 (N_4131,In_1898,In_1995);
nand U4132 (N_4132,In_33,In_1251);
nor U4133 (N_4133,In_1887,In_119);
nor U4134 (N_4134,In_2173,In_1826);
xnor U4135 (N_4135,In_488,In_1180);
nor U4136 (N_4136,In_1630,In_95);
nand U4137 (N_4137,In_1793,In_953);
xnor U4138 (N_4138,In_897,In_2077);
and U4139 (N_4139,In_1829,In_1113);
or U4140 (N_4140,In_143,In_1005);
xnor U4141 (N_4141,In_1175,In_210);
or U4142 (N_4142,In_110,In_937);
nor U4143 (N_4143,In_2438,In_2429);
xnor U4144 (N_4144,In_2115,In_1839);
nand U4145 (N_4145,In_863,In_245);
xnor U4146 (N_4146,In_1874,In_1897);
xnor U4147 (N_4147,In_1978,In_1943);
or U4148 (N_4148,In_1775,In_1917);
and U4149 (N_4149,In_2297,In_1402);
xor U4150 (N_4150,In_637,In_1944);
and U4151 (N_4151,In_2316,In_2390);
nand U4152 (N_4152,In_1502,In_2332);
xor U4153 (N_4153,In_1185,In_2435);
nand U4154 (N_4154,In_161,In_1357);
and U4155 (N_4155,In_802,In_2131);
nor U4156 (N_4156,In_1896,In_2277);
nand U4157 (N_4157,In_194,In_2202);
xnor U4158 (N_4158,In_1510,In_2108);
and U4159 (N_4159,In_857,In_789);
or U4160 (N_4160,In_1808,In_1468);
xor U4161 (N_4161,In_757,In_2362);
xor U4162 (N_4162,In_488,In_391);
nand U4163 (N_4163,In_2014,In_2238);
and U4164 (N_4164,In_337,In_1927);
xnor U4165 (N_4165,In_1529,In_112);
and U4166 (N_4166,In_2260,In_938);
nand U4167 (N_4167,In_677,In_1991);
nand U4168 (N_4168,In_1797,In_1643);
nor U4169 (N_4169,In_410,In_1708);
and U4170 (N_4170,In_2364,In_2167);
or U4171 (N_4171,In_1249,In_1985);
nand U4172 (N_4172,In_1737,In_959);
nand U4173 (N_4173,In_1349,In_495);
nand U4174 (N_4174,In_2218,In_1228);
nor U4175 (N_4175,In_2372,In_647);
nand U4176 (N_4176,In_754,In_12);
or U4177 (N_4177,In_0,In_1797);
nor U4178 (N_4178,In_1242,In_1111);
nor U4179 (N_4179,In_2295,In_1522);
nor U4180 (N_4180,In_1924,In_409);
and U4181 (N_4181,In_183,In_1957);
or U4182 (N_4182,In_839,In_412);
nor U4183 (N_4183,In_363,In_826);
or U4184 (N_4184,In_1692,In_1694);
and U4185 (N_4185,In_755,In_776);
xnor U4186 (N_4186,In_808,In_1297);
xnor U4187 (N_4187,In_1013,In_1822);
and U4188 (N_4188,In_969,In_2018);
and U4189 (N_4189,In_748,In_822);
nand U4190 (N_4190,In_1952,In_2025);
nor U4191 (N_4191,In_312,In_1163);
and U4192 (N_4192,In_105,In_2305);
nand U4193 (N_4193,In_1724,In_132);
nand U4194 (N_4194,In_1373,In_733);
or U4195 (N_4195,In_1990,In_329);
nand U4196 (N_4196,In_1397,In_1038);
xnor U4197 (N_4197,In_727,In_1673);
nor U4198 (N_4198,In_318,In_272);
or U4199 (N_4199,In_2354,In_762);
xor U4200 (N_4200,In_735,In_2255);
nand U4201 (N_4201,In_903,In_499);
or U4202 (N_4202,In_1999,In_959);
and U4203 (N_4203,In_587,In_812);
or U4204 (N_4204,In_1550,In_2256);
nor U4205 (N_4205,In_1345,In_2265);
nand U4206 (N_4206,In_2407,In_2220);
and U4207 (N_4207,In_1358,In_705);
or U4208 (N_4208,In_2417,In_60);
nand U4209 (N_4209,In_2472,In_1205);
nand U4210 (N_4210,In_1803,In_741);
nor U4211 (N_4211,In_2294,In_264);
nand U4212 (N_4212,In_1853,In_1123);
nand U4213 (N_4213,In_2162,In_647);
or U4214 (N_4214,In_2400,In_756);
or U4215 (N_4215,In_2330,In_54);
or U4216 (N_4216,In_2359,In_2053);
nand U4217 (N_4217,In_52,In_1264);
and U4218 (N_4218,In_1825,In_1593);
xor U4219 (N_4219,In_778,In_453);
or U4220 (N_4220,In_2348,In_1663);
and U4221 (N_4221,In_78,In_156);
and U4222 (N_4222,In_2239,In_1223);
and U4223 (N_4223,In_109,In_1659);
and U4224 (N_4224,In_272,In_118);
xor U4225 (N_4225,In_2490,In_2431);
or U4226 (N_4226,In_2100,In_295);
xnor U4227 (N_4227,In_196,In_636);
nand U4228 (N_4228,In_1812,In_2029);
or U4229 (N_4229,In_2024,In_708);
nand U4230 (N_4230,In_1401,In_1630);
nor U4231 (N_4231,In_532,In_438);
xnor U4232 (N_4232,In_752,In_2149);
and U4233 (N_4233,In_2368,In_2273);
or U4234 (N_4234,In_1085,In_1031);
xnor U4235 (N_4235,In_1399,In_1960);
and U4236 (N_4236,In_1817,In_419);
xor U4237 (N_4237,In_654,In_2015);
nor U4238 (N_4238,In_899,In_1242);
and U4239 (N_4239,In_1606,In_812);
xnor U4240 (N_4240,In_2092,In_659);
and U4241 (N_4241,In_2161,In_1117);
and U4242 (N_4242,In_1151,In_1970);
xor U4243 (N_4243,In_743,In_1037);
nor U4244 (N_4244,In_1932,In_1578);
xor U4245 (N_4245,In_562,In_522);
xnor U4246 (N_4246,In_1145,In_603);
and U4247 (N_4247,In_1326,In_2181);
xor U4248 (N_4248,In_2299,In_1709);
or U4249 (N_4249,In_1223,In_1665);
or U4250 (N_4250,In_2077,In_385);
nor U4251 (N_4251,In_810,In_1501);
xor U4252 (N_4252,In_416,In_1425);
nand U4253 (N_4253,In_689,In_1149);
nand U4254 (N_4254,In_428,In_831);
nor U4255 (N_4255,In_2234,In_1513);
nand U4256 (N_4256,In_2320,In_1385);
nand U4257 (N_4257,In_259,In_1044);
xor U4258 (N_4258,In_2424,In_896);
xnor U4259 (N_4259,In_2007,In_216);
and U4260 (N_4260,In_1491,In_1100);
nand U4261 (N_4261,In_50,In_212);
and U4262 (N_4262,In_664,In_778);
nor U4263 (N_4263,In_758,In_839);
nor U4264 (N_4264,In_753,In_918);
and U4265 (N_4265,In_1383,In_1527);
nand U4266 (N_4266,In_2190,In_1957);
xnor U4267 (N_4267,In_1795,In_2070);
nand U4268 (N_4268,In_1350,In_180);
or U4269 (N_4269,In_27,In_1984);
and U4270 (N_4270,In_417,In_1556);
nand U4271 (N_4271,In_1582,In_718);
and U4272 (N_4272,In_1152,In_283);
nor U4273 (N_4273,In_1811,In_806);
xor U4274 (N_4274,In_202,In_2296);
and U4275 (N_4275,In_1438,In_258);
nand U4276 (N_4276,In_2147,In_840);
or U4277 (N_4277,In_994,In_1103);
or U4278 (N_4278,In_727,In_2243);
nand U4279 (N_4279,In_1150,In_678);
and U4280 (N_4280,In_1352,In_41);
and U4281 (N_4281,In_1197,In_473);
and U4282 (N_4282,In_1653,In_1902);
and U4283 (N_4283,In_1368,In_180);
nor U4284 (N_4284,In_1626,In_2291);
or U4285 (N_4285,In_497,In_849);
or U4286 (N_4286,In_559,In_1587);
or U4287 (N_4287,In_1388,In_1723);
nand U4288 (N_4288,In_1121,In_1720);
or U4289 (N_4289,In_1225,In_2063);
nor U4290 (N_4290,In_2255,In_2273);
xor U4291 (N_4291,In_1677,In_583);
or U4292 (N_4292,In_900,In_54);
and U4293 (N_4293,In_918,In_248);
and U4294 (N_4294,In_2097,In_1413);
nor U4295 (N_4295,In_1886,In_45);
xor U4296 (N_4296,In_1857,In_1239);
xor U4297 (N_4297,In_120,In_2327);
and U4298 (N_4298,In_516,In_1379);
xnor U4299 (N_4299,In_524,In_363);
xnor U4300 (N_4300,In_18,In_396);
and U4301 (N_4301,In_1377,In_1119);
or U4302 (N_4302,In_412,In_2475);
or U4303 (N_4303,In_781,In_2106);
xor U4304 (N_4304,In_217,In_1790);
nor U4305 (N_4305,In_1307,In_1845);
or U4306 (N_4306,In_2335,In_576);
or U4307 (N_4307,In_322,In_680);
xor U4308 (N_4308,In_1474,In_2146);
and U4309 (N_4309,In_1928,In_759);
nand U4310 (N_4310,In_308,In_1926);
nand U4311 (N_4311,In_1822,In_2201);
nor U4312 (N_4312,In_1472,In_1525);
nand U4313 (N_4313,In_720,In_424);
or U4314 (N_4314,In_2391,In_1837);
nor U4315 (N_4315,In_154,In_1912);
nand U4316 (N_4316,In_2173,In_120);
nand U4317 (N_4317,In_2108,In_556);
or U4318 (N_4318,In_808,In_1286);
or U4319 (N_4319,In_1021,In_1555);
or U4320 (N_4320,In_1007,In_2254);
nand U4321 (N_4321,In_2020,In_2492);
xnor U4322 (N_4322,In_2090,In_515);
or U4323 (N_4323,In_1692,In_1458);
nand U4324 (N_4324,In_74,In_748);
nor U4325 (N_4325,In_1697,In_574);
nor U4326 (N_4326,In_165,In_282);
nand U4327 (N_4327,In_1372,In_329);
nand U4328 (N_4328,In_172,In_1943);
xor U4329 (N_4329,In_605,In_1700);
nand U4330 (N_4330,In_1597,In_2081);
nor U4331 (N_4331,In_1191,In_2350);
xor U4332 (N_4332,In_556,In_1288);
or U4333 (N_4333,In_2052,In_726);
nand U4334 (N_4334,In_265,In_2236);
xor U4335 (N_4335,In_1442,In_1724);
and U4336 (N_4336,In_2392,In_1706);
xor U4337 (N_4337,In_1313,In_2295);
nor U4338 (N_4338,In_1078,In_852);
nor U4339 (N_4339,In_1133,In_510);
nand U4340 (N_4340,In_960,In_2418);
nor U4341 (N_4341,In_805,In_920);
nor U4342 (N_4342,In_2105,In_2005);
nor U4343 (N_4343,In_480,In_843);
and U4344 (N_4344,In_773,In_364);
nand U4345 (N_4345,In_318,In_2008);
xnor U4346 (N_4346,In_1843,In_1660);
nand U4347 (N_4347,In_2053,In_2162);
and U4348 (N_4348,In_1022,In_1168);
nor U4349 (N_4349,In_1321,In_1843);
nor U4350 (N_4350,In_246,In_1767);
nor U4351 (N_4351,In_1415,In_149);
nor U4352 (N_4352,In_2315,In_1933);
and U4353 (N_4353,In_1892,In_290);
nand U4354 (N_4354,In_2077,In_2171);
nor U4355 (N_4355,In_1098,In_739);
xnor U4356 (N_4356,In_2119,In_943);
or U4357 (N_4357,In_1750,In_909);
or U4358 (N_4358,In_959,In_1843);
nor U4359 (N_4359,In_2395,In_589);
nand U4360 (N_4360,In_1252,In_1623);
and U4361 (N_4361,In_1664,In_1066);
nand U4362 (N_4362,In_32,In_1378);
nand U4363 (N_4363,In_1065,In_1715);
xnor U4364 (N_4364,In_1568,In_1762);
nor U4365 (N_4365,In_1556,In_352);
or U4366 (N_4366,In_33,In_248);
and U4367 (N_4367,In_1202,In_272);
or U4368 (N_4368,In_1246,In_1814);
and U4369 (N_4369,In_1516,In_784);
and U4370 (N_4370,In_1122,In_732);
or U4371 (N_4371,In_2398,In_1630);
nand U4372 (N_4372,In_2476,In_94);
xor U4373 (N_4373,In_34,In_911);
nand U4374 (N_4374,In_1209,In_1656);
nor U4375 (N_4375,In_2473,In_25);
or U4376 (N_4376,In_2064,In_128);
and U4377 (N_4377,In_934,In_1662);
xor U4378 (N_4378,In_76,In_1341);
nor U4379 (N_4379,In_1230,In_1277);
xnor U4380 (N_4380,In_2257,In_689);
nand U4381 (N_4381,In_1839,In_1860);
xor U4382 (N_4382,In_251,In_1030);
xnor U4383 (N_4383,In_1009,In_1984);
and U4384 (N_4384,In_166,In_691);
nand U4385 (N_4385,In_2318,In_723);
or U4386 (N_4386,In_650,In_2030);
or U4387 (N_4387,In_1197,In_36);
xor U4388 (N_4388,In_917,In_1808);
or U4389 (N_4389,In_2283,In_1348);
and U4390 (N_4390,In_229,In_1431);
or U4391 (N_4391,In_1936,In_513);
or U4392 (N_4392,In_957,In_1701);
or U4393 (N_4393,In_2231,In_1463);
nand U4394 (N_4394,In_2045,In_1232);
xnor U4395 (N_4395,In_2485,In_1571);
xnor U4396 (N_4396,In_1303,In_154);
or U4397 (N_4397,In_1949,In_366);
xnor U4398 (N_4398,In_106,In_393);
and U4399 (N_4399,In_518,In_2403);
or U4400 (N_4400,In_1610,In_2067);
xor U4401 (N_4401,In_1746,In_233);
xor U4402 (N_4402,In_938,In_808);
nor U4403 (N_4403,In_1396,In_204);
xnor U4404 (N_4404,In_2444,In_1636);
or U4405 (N_4405,In_113,In_2005);
nor U4406 (N_4406,In_1190,In_70);
xnor U4407 (N_4407,In_737,In_2202);
and U4408 (N_4408,In_2446,In_2109);
nand U4409 (N_4409,In_336,In_2322);
nand U4410 (N_4410,In_120,In_2293);
nand U4411 (N_4411,In_1239,In_1969);
nor U4412 (N_4412,In_1854,In_2160);
and U4413 (N_4413,In_644,In_2438);
and U4414 (N_4414,In_1942,In_373);
or U4415 (N_4415,In_1526,In_610);
nor U4416 (N_4416,In_604,In_926);
nand U4417 (N_4417,In_2157,In_1906);
nor U4418 (N_4418,In_2337,In_761);
xnor U4419 (N_4419,In_6,In_1923);
nor U4420 (N_4420,In_2041,In_2005);
xnor U4421 (N_4421,In_875,In_727);
xor U4422 (N_4422,In_1204,In_2351);
or U4423 (N_4423,In_2404,In_379);
or U4424 (N_4424,In_197,In_709);
xnor U4425 (N_4425,In_2406,In_1095);
xnor U4426 (N_4426,In_1900,In_1464);
and U4427 (N_4427,In_97,In_1929);
nor U4428 (N_4428,In_1129,In_1363);
nand U4429 (N_4429,In_1600,In_2222);
nand U4430 (N_4430,In_1108,In_1556);
nand U4431 (N_4431,In_1925,In_571);
xnor U4432 (N_4432,In_748,In_1594);
and U4433 (N_4433,In_405,In_1964);
and U4434 (N_4434,In_2406,In_1468);
nand U4435 (N_4435,In_1372,In_2139);
nand U4436 (N_4436,In_1427,In_2175);
nand U4437 (N_4437,In_1855,In_1358);
xor U4438 (N_4438,In_1653,In_339);
or U4439 (N_4439,In_507,In_1766);
and U4440 (N_4440,In_344,In_531);
nand U4441 (N_4441,In_2320,In_2111);
nand U4442 (N_4442,In_2234,In_2113);
or U4443 (N_4443,In_687,In_1322);
and U4444 (N_4444,In_935,In_1992);
nor U4445 (N_4445,In_1494,In_1505);
and U4446 (N_4446,In_1522,In_57);
nor U4447 (N_4447,In_1212,In_304);
nand U4448 (N_4448,In_887,In_2131);
xor U4449 (N_4449,In_696,In_618);
nand U4450 (N_4450,In_44,In_2426);
and U4451 (N_4451,In_544,In_572);
or U4452 (N_4452,In_644,In_2346);
and U4453 (N_4453,In_241,In_2132);
nand U4454 (N_4454,In_2023,In_840);
or U4455 (N_4455,In_321,In_740);
and U4456 (N_4456,In_2328,In_2370);
or U4457 (N_4457,In_288,In_2058);
xor U4458 (N_4458,In_2384,In_550);
nor U4459 (N_4459,In_1792,In_2280);
and U4460 (N_4460,In_1489,In_123);
or U4461 (N_4461,In_2337,In_1151);
nand U4462 (N_4462,In_488,In_955);
and U4463 (N_4463,In_412,In_135);
nand U4464 (N_4464,In_604,In_2000);
nor U4465 (N_4465,In_240,In_534);
nand U4466 (N_4466,In_390,In_773);
or U4467 (N_4467,In_20,In_540);
xnor U4468 (N_4468,In_800,In_2349);
xor U4469 (N_4469,In_1153,In_2191);
and U4470 (N_4470,In_1714,In_411);
xor U4471 (N_4471,In_362,In_2161);
xnor U4472 (N_4472,In_186,In_1563);
and U4473 (N_4473,In_397,In_1001);
nor U4474 (N_4474,In_370,In_1117);
nor U4475 (N_4475,In_238,In_2422);
xor U4476 (N_4476,In_1692,In_923);
nand U4477 (N_4477,In_1717,In_1245);
or U4478 (N_4478,In_291,In_1766);
and U4479 (N_4479,In_754,In_1498);
nand U4480 (N_4480,In_467,In_432);
and U4481 (N_4481,In_334,In_801);
nand U4482 (N_4482,In_615,In_846);
or U4483 (N_4483,In_2224,In_1497);
or U4484 (N_4484,In_632,In_1501);
xor U4485 (N_4485,In_1462,In_1020);
or U4486 (N_4486,In_2060,In_1218);
nor U4487 (N_4487,In_2130,In_2260);
nor U4488 (N_4488,In_63,In_534);
nand U4489 (N_4489,In_1859,In_1286);
and U4490 (N_4490,In_2072,In_1590);
xor U4491 (N_4491,In_1253,In_2137);
nor U4492 (N_4492,In_90,In_264);
xnor U4493 (N_4493,In_1968,In_2197);
or U4494 (N_4494,In_37,In_1494);
nor U4495 (N_4495,In_831,In_976);
nor U4496 (N_4496,In_1265,In_421);
nor U4497 (N_4497,In_2495,In_54);
xnor U4498 (N_4498,In_1623,In_1292);
nor U4499 (N_4499,In_1895,In_1802);
xor U4500 (N_4500,In_1243,In_642);
or U4501 (N_4501,In_1815,In_346);
nand U4502 (N_4502,In_1360,In_2229);
or U4503 (N_4503,In_2020,In_2244);
or U4504 (N_4504,In_159,In_894);
and U4505 (N_4505,In_1417,In_477);
or U4506 (N_4506,In_603,In_925);
nor U4507 (N_4507,In_308,In_152);
xnor U4508 (N_4508,In_544,In_512);
and U4509 (N_4509,In_2323,In_1213);
and U4510 (N_4510,In_1018,In_1157);
nand U4511 (N_4511,In_1979,In_2209);
or U4512 (N_4512,In_1898,In_1839);
and U4513 (N_4513,In_199,In_1619);
nand U4514 (N_4514,In_1651,In_30);
xor U4515 (N_4515,In_479,In_257);
or U4516 (N_4516,In_1533,In_1264);
nor U4517 (N_4517,In_853,In_1646);
or U4518 (N_4518,In_1779,In_586);
and U4519 (N_4519,In_1822,In_2137);
and U4520 (N_4520,In_2229,In_818);
or U4521 (N_4521,In_2366,In_1331);
nand U4522 (N_4522,In_1654,In_2285);
or U4523 (N_4523,In_65,In_2472);
and U4524 (N_4524,In_2266,In_744);
and U4525 (N_4525,In_650,In_579);
nand U4526 (N_4526,In_1637,In_712);
or U4527 (N_4527,In_1133,In_2195);
or U4528 (N_4528,In_1526,In_769);
nor U4529 (N_4529,In_2255,In_1522);
or U4530 (N_4530,In_1992,In_944);
or U4531 (N_4531,In_701,In_2219);
xnor U4532 (N_4532,In_511,In_592);
nand U4533 (N_4533,In_505,In_2113);
nor U4534 (N_4534,In_1686,In_1168);
xor U4535 (N_4535,In_1606,In_842);
or U4536 (N_4536,In_2273,In_182);
or U4537 (N_4537,In_2124,In_420);
nor U4538 (N_4538,In_473,In_1762);
and U4539 (N_4539,In_2281,In_77);
and U4540 (N_4540,In_853,In_2218);
xnor U4541 (N_4541,In_680,In_1317);
or U4542 (N_4542,In_843,In_1266);
and U4543 (N_4543,In_67,In_329);
xor U4544 (N_4544,In_2001,In_1578);
nor U4545 (N_4545,In_1538,In_746);
and U4546 (N_4546,In_362,In_755);
and U4547 (N_4547,In_207,In_1069);
nand U4548 (N_4548,In_1888,In_2091);
nor U4549 (N_4549,In_17,In_1549);
and U4550 (N_4550,In_765,In_1631);
xor U4551 (N_4551,In_464,In_1705);
nand U4552 (N_4552,In_1649,In_2047);
and U4553 (N_4553,In_701,In_2008);
nand U4554 (N_4554,In_1334,In_1250);
and U4555 (N_4555,In_1038,In_342);
xnor U4556 (N_4556,In_951,In_1080);
or U4557 (N_4557,In_684,In_1054);
nand U4558 (N_4558,In_683,In_1274);
or U4559 (N_4559,In_935,In_1579);
xnor U4560 (N_4560,In_521,In_1130);
nand U4561 (N_4561,In_1353,In_1066);
and U4562 (N_4562,In_428,In_1500);
xnor U4563 (N_4563,In_572,In_596);
nand U4564 (N_4564,In_1106,In_2157);
xnor U4565 (N_4565,In_1892,In_677);
xnor U4566 (N_4566,In_2233,In_575);
and U4567 (N_4567,In_1121,In_2134);
xnor U4568 (N_4568,In_498,In_2139);
or U4569 (N_4569,In_1714,In_391);
nand U4570 (N_4570,In_1792,In_2165);
and U4571 (N_4571,In_1838,In_1980);
nor U4572 (N_4572,In_662,In_411);
nand U4573 (N_4573,In_252,In_610);
xnor U4574 (N_4574,In_850,In_671);
or U4575 (N_4575,In_946,In_629);
nor U4576 (N_4576,In_1845,In_1674);
or U4577 (N_4577,In_910,In_1970);
nor U4578 (N_4578,In_846,In_1508);
and U4579 (N_4579,In_1898,In_84);
or U4580 (N_4580,In_1051,In_1693);
or U4581 (N_4581,In_891,In_2237);
and U4582 (N_4582,In_1533,In_1471);
nor U4583 (N_4583,In_1632,In_1179);
nor U4584 (N_4584,In_1654,In_749);
or U4585 (N_4585,In_903,In_1259);
and U4586 (N_4586,In_675,In_1610);
nand U4587 (N_4587,In_376,In_1478);
xnor U4588 (N_4588,In_1105,In_668);
or U4589 (N_4589,In_985,In_201);
xor U4590 (N_4590,In_1963,In_1060);
and U4591 (N_4591,In_1492,In_794);
nand U4592 (N_4592,In_817,In_763);
nor U4593 (N_4593,In_1785,In_1042);
nor U4594 (N_4594,In_1461,In_230);
and U4595 (N_4595,In_710,In_1778);
nand U4596 (N_4596,In_1893,In_1755);
nand U4597 (N_4597,In_1189,In_1595);
or U4598 (N_4598,In_1382,In_1747);
xor U4599 (N_4599,In_208,In_1374);
and U4600 (N_4600,In_2436,In_1507);
nor U4601 (N_4601,In_1486,In_316);
and U4602 (N_4602,In_1814,In_1293);
xor U4603 (N_4603,In_120,In_590);
or U4604 (N_4604,In_543,In_722);
and U4605 (N_4605,In_503,In_22);
nor U4606 (N_4606,In_682,In_1158);
nor U4607 (N_4607,In_771,In_920);
xor U4608 (N_4608,In_1744,In_2182);
nor U4609 (N_4609,In_1182,In_2126);
nor U4610 (N_4610,In_455,In_1553);
and U4611 (N_4611,In_2214,In_2431);
xor U4612 (N_4612,In_997,In_2063);
and U4613 (N_4613,In_478,In_41);
and U4614 (N_4614,In_412,In_1846);
or U4615 (N_4615,In_773,In_1341);
nand U4616 (N_4616,In_320,In_1491);
and U4617 (N_4617,In_1612,In_2133);
nand U4618 (N_4618,In_2172,In_839);
xnor U4619 (N_4619,In_591,In_2258);
nor U4620 (N_4620,In_526,In_1997);
nand U4621 (N_4621,In_2038,In_918);
and U4622 (N_4622,In_2185,In_1248);
and U4623 (N_4623,In_1139,In_927);
and U4624 (N_4624,In_986,In_266);
or U4625 (N_4625,In_1600,In_835);
and U4626 (N_4626,In_1540,In_874);
or U4627 (N_4627,In_776,In_675);
or U4628 (N_4628,In_2444,In_1059);
xnor U4629 (N_4629,In_1098,In_1704);
and U4630 (N_4630,In_848,In_2445);
or U4631 (N_4631,In_592,In_1514);
and U4632 (N_4632,In_1005,In_1724);
nor U4633 (N_4633,In_1248,In_1808);
xor U4634 (N_4634,In_2304,In_1986);
nor U4635 (N_4635,In_1042,In_2152);
nor U4636 (N_4636,In_1192,In_1105);
xnor U4637 (N_4637,In_579,In_2275);
nand U4638 (N_4638,In_1974,In_335);
and U4639 (N_4639,In_1938,In_2095);
xnor U4640 (N_4640,In_2202,In_1444);
nor U4641 (N_4641,In_1652,In_257);
xnor U4642 (N_4642,In_2313,In_2222);
xor U4643 (N_4643,In_685,In_1751);
xnor U4644 (N_4644,In_683,In_2199);
xnor U4645 (N_4645,In_1470,In_1359);
nor U4646 (N_4646,In_281,In_2494);
xnor U4647 (N_4647,In_404,In_399);
nand U4648 (N_4648,In_1748,In_855);
nand U4649 (N_4649,In_1996,In_1263);
nor U4650 (N_4650,In_634,In_1624);
nor U4651 (N_4651,In_448,In_759);
or U4652 (N_4652,In_1995,In_117);
nand U4653 (N_4653,In_1150,In_1814);
and U4654 (N_4654,In_1019,In_1565);
and U4655 (N_4655,In_36,In_824);
nor U4656 (N_4656,In_306,In_2076);
and U4657 (N_4657,In_197,In_691);
xor U4658 (N_4658,In_826,In_235);
nor U4659 (N_4659,In_645,In_2035);
and U4660 (N_4660,In_629,In_960);
nor U4661 (N_4661,In_1214,In_256);
nand U4662 (N_4662,In_1430,In_1282);
nand U4663 (N_4663,In_1275,In_1175);
and U4664 (N_4664,In_1096,In_2166);
xnor U4665 (N_4665,In_1922,In_1332);
nor U4666 (N_4666,In_1018,In_251);
nor U4667 (N_4667,In_30,In_209);
or U4668 (N_4668,In_663,In_2328);
xor U4669 (N_4669,In_1556,In_1954);
xor U4670 (N_4670,In_1822,In_1101);
nor U4671 (N_4671,In_430,In_1282);
xnor U4672 (N_4672,In_1582,In_1064);
xnor U4673 (N_4673,In_704,In_1381);
or U4674 (N_4674,In_1359,In_508);
or U4675 (N_4675,In_585,In_114);
or U4676 (N_4676,In_1740,In_2094);
nand U4677 (N_4677,In_845,In_584);
and U4678 (N_4678,In_187,In_183);
and U4679 (N_4679,In_1863,In_440);
or U4680 (N_4680,In_1696,In_1327);
nand U4681 (N_4681,In_665,In_2083);
nor U4682 (N_4682,In_1155,In_857);
nand U4683 (N_4683,In_1161,In_583);
or U4684 (N_4684,In_1259,In_139);
or U4685 (N_4685,In_2036,In_2248);
xnor U4686 (N_4686,In_590,In_305);
xor U4687 (N_4687,In_2,In_2239);
or U4688 (N_4688,In_2284,In_1153);
nor U4689 (N_4689,In_791,In_1083);
or U4690 (N_4690,In_208,In_2083);
nor U4691 (N_4691,In_1798,In_270);
or U4692 (N_4692,In_1198,In_2012);
xor U4693 (N_4693,In_139,In_589);
xor U4694 (N_4694,In_644,In_347);
or U4695 (N_4695,In_2265,In_2120);
xnor U4696 (N_4696,In_646,In_1701);
and U4697 (N_4697,In_240,In_308);
or U4698 (N_4698,In_415,In_1152);
and U4699 (N_4699,In_175,In_1376);
xnor U4700 (N_4700,In_1072,In_243);
nor U4701 (N_4701,In_989,In_159);
nor U4702 (N_4702,In_465,In_473);
xor U4703 (N_4703,In_2001,In_1615);
or U4704 (N_4704,In_2133,In_1738);
or U4705 (N_4705,In_983,In_242);
or U4706 (N_4706,In_2176,In_657);
or U4707 (N_4707,In_2149,In_1339);
or U4708 (N_4708,In_958,In_623);
nand U4709 (N_4709,In_1516,In_2458);
and U4710 (N_4710,In_1224,In_1515);
xnor U4711 (N_4711,In_1819,In_1958);
nand U4712 (N_4712,In_1761,In_2195);
and U4713 (N_4713,In_1113,In_927);
and U4714 (N_4714,In_1168,In_441);
nand U4715 (N_4715,In_1938,In_1511);
nand U4716 (N_4716,In_714,In_198);
nand U4717 (N_4717,In_1583,In_0);
and U4718 (N_4718,In_2213,In_2344);
and U4719 (N_4719,In_1469,In_784);
or U4720 (N_4720,In_1058,In_964);
nand U4721 (N_4721,In_1212,In_1542);
nand U4722 (N_4722,In_2333,In_417);
nor U4723 (N_4723,In_2044,In_1527);
nand U4724 (N_4724,In_1787,In_1752);
nor U4725 (N_4725,In_1279,In_1905);
nor U4726 (N_4726,In_2316,In_816);
xor U4727 (N_4727,In_2472,In_29);
xor U4728 (N_4728,In_2235,In_286);
or U4729 (N_4729,In_1415,In_1806);
and U4730 (N_4730,In_2191,In_1909);
or U4731 (N_4731,In_235,In_225);
nand U4732 (N_4732,In_2310,In_1224);
xnor U4733 (N_4733,In_2106,In_798);
or U4734 (N_4734,In_2,In_2333);
nor U4735 (N_4735,In_2150,In_794);
xnor U4736 (N_4736,In_125,In_1738);
and U4737 (N_4737,In_2402,In_1122);
and U4738 (N_4738,In_1762,In_966);
nand U4739 (N_4739,In_614,In_1983);
xnor U4740 (N_4740,In_1962,In_1118);
or U4741 (N_4741,In_2208,In_1281);
xnor U4742 (N_4742,In_984,In_148);
and U4743 (N_4743,In_954,In_1220);
and U4744 (N_4744,In_2235,In_1233);
xnor U4745 (N_4745,In_2204,In_1827);
nor U4746 (N_4746,In_2009,In_1318);
nand U4747 (N_4747,In_705,In_274);
or U4748 (N_4748,In_2466,In_2082);
nor U4749 (N_4749,In_1541,In_485);
nand U4750 (N_4750,In_2348,In_2006);
nand U4751 (N_4751,In_1768,In_2005);
nand U4752 (N_4752,In_368,In_1164);
or U4753 (N_4753,In_746,In_468);
and U4754 (N_4754,In_945,In_164);
and U4755 (N_4755,In_173,In_913);
nand U4756 (N_4756,In_2153,In_554);
xor U4757 (N_4757,In_1409,In_1910);
and U4758 (N_4758,In_1516,In_1450);
or U4759 (N_4759,In_1837,In_683);
nor U4760 (N_4760,In_478,In_1247);
and U4761 (N_4761,In_1311,In_601);
and U4762 (N_4762,In_208,In_1138);
xnor U4763 (N_4763,In_2184,In_1802);
xnor U4764 (N_4764,In_2229,In_1790);
nor U4765 (N_4765,In_2266,In_2315);
xnor U4766 (N_4766,In_694,In_1071);
nor U4767 (N_4767,In_186,In_1540);
nor U4768 (N_4768,In_1846,In_758);
nand U4769 (N_4769,In_2426,In_1100);
nand U4770 (N_4770,In_1613,In_113);
and U4771 (N_4771,In_1235,In_2480);
nor U4772 (N_4772,In_2346,In_1049);
xor U4773 (N_4773,In_522,In_1337);
or U4774 (N_4774,In_2486,In_1397);
nand U4775 (N_4775,In_1497,In_673);
nor U4776 (N_4776,In_792,In_744);
xor U4777 (N_4777,In_125,In_379);
xor U4778 (N_4778,In_1553,In_2049);
and U4779 (N_4779,In_137,In_1079);
and U4780 (N_4780,In_344,In_854);
nor U4781 (N_4781,In_1873,In_1761);
nor U4782 (N_4782,In_2456,In_1156);
xor U4783 (N_4783,In_2046,In_1424);
nand U4784 (N_4784,In_2393,In_2378);
and U4785 (N_4785,In_1967,In_1832);
and U4786 (N_4786,In_2397,In_1602);
or U4787 (N_4787,In_1837,In_2187);
xor U4788 (N_4788,In_938,In_44);
nand U4789 (N_4789,In_2079,In_1117);
and U4790 (N_4790,In_1894,In_181);
xnor U4791 (N_4791,In_1465,In_2124);
nand U4792 (N_4792,In_2016,In_2188);
nor U4793 (N_4793,In_500,In_2364);
and U4794 (N_4794,In_1275,In_1064);
nand U4795 (N_4795,In_1092,In_856);
or U4796 (N_4796,In_1115,In_281);
and U4797 (N_4797,In_423,In_2371);
xnor U4798 (N_4798,In_108,In_1152);
nand U4799 (N_4799,In_55,In_2233);
nand U4800 (N_4800,In_1968,In_25);
xor U4801 (N_4801,In_817,In_489);
and U4802 (N_4802,In_141,In_1832);
nor U4803 (N_4803,In_2306,In_2120);
xor U4804 (N_4804,In_815,In_480);
or U4805 (N_4805,In_1427,In_2453);
nand U4806 (N_4806,In_1087,In_2022);
or U4807 (N_4807,In_769,In_2154);
and U4808 (N_4808,In_1512,In_1681);
or U4809 (N_4809,In_568,In_1576);
or U4810 (N_4810,In_2293,In_388);
or U4811 (N_4811,In_1693,In_30);
nand U4812 (N_4812,In_385,In_1169);
nand U4813 (N_4813,In_1281,In_872);
or U4814 (N_4814,In_1926,In_930);
xnor U4815 (N_4815,In_330,In_438);
and U4816 (N_4816,In_1306,In_1979);
xor U4817 (N_4817,In_166,In_285);
or U4818 (N_4818,In_2197,In_1704);
or U4819 (N_4819,In_1403,In_2156);
nor U4820 (N_4820,In_736,In_1024);
or U4821 (N_4821,In_1152,In_1212);
nor U4822 (N_4822,In_1936,In_1347);
nand U4823 (N_4823,In_1564,In_1783);
and U4824 (N_4824,In_1968,In_1711);
and U4825 (N_4825,In_2158,In_1255);
and U4826 (N_4826,In_2452,In_343);
and U4827 (N_4827,In_616,In_2307);
or U4828 (N_4828,In_1360,In_182);
and U4829 (N_4829,In_1459,In_479);
xnor U4830 (N_4830,In_1928,In_1198);
xor U4831 (N_4831,In_73,In_1409);
xor U4832 (N_4832,In_2478,In_969);
and U4833 (N_4833,In_2025,In_5);
and U4834 (N_4834,In_317,In_139);
nand U4835 (N_4835,In_123,In_1308);
or U4836 (N_4836,In_950,In_1891);
or U4837 (N_4837,In_877,In_247);
and U4838 (N_4838,In_1586,In_2356);
nand U4839 (N_4839,In_679,In_1109);
or U4840 (N_4840,In_236,In_2301);
nand U4841 (N_4841,In_46,In_2131);
and U4842 (N_4842,In_1321,In_2165);
nand U4843 (N_4843,In_785,In_929);
xnor U4844 (N_4844,In_1990,In_136);
nand U4845 (N_4845,In_2409,In_1994);
xor U4846 (N_4846,In_765,In_1163);
nand U4847 (N_4847,In_1898,In_348);
or U4848 (N_4848,In_209,In_2174);
nor U4849 (N_4849,In_1484,In_1138);
nor U4850 (N_4850,In_1468,In_320);
nor U4851 (N_4851,In_765,In_171);
and U4852 (N_4852,In_2400,In_573);
and U4853 (N_4853,In_1710,In_379);
or U4854 (N_4854,In_2326,In_1444);
xor U4855 (N_4855,In_189,In_478);
and U4856 (N_4856,In_889,In_1183);
nor U4857 (N_4857,In_1152,In_691);
and U4858 (N_4858,In_74,In_648);
and U4859 (N_4859,In_928,In_398);
or U4860 (N_4860,In_692,In_2097);
nand U4861 (N_4861,In_485,In_2370);
or U4862 (N_4862,In_1078,In_1848);
or U4863 (N_4863,In_1262,In_2265);
xnor U4864 (N_4864,In_543,In_1867);
nor U4865 (N_4865,In_317,In_1523);
nor U4866 (N_4866,In_672,In_878);
nand U4867 (N_4867,In_257,In_17);
xor U4868 (N_4868,In_2226,In_596);
or U4869 (N_4869,In_596,In_26);
nand U4870 (N_4870,In_1109,In_849);
or U4871 (N_4871,In_232,In_1685);
nor U4872 (N_4872,In_2313,In_2256);
nor U4873 (N_4873,In_2206,In_1443);
or U4874 (N_4874,In_1673,In_1106);
xnor U4875 (N_4875,In_2370,In_2235);
or U4876 (N_4876,In_254,In_449);
nand U4877 (N_4877,In_1317,In_2150);
nor U4878 (N_4878,In_2323,In_428);
nand U4879 (N_4879,In_993,In_427);
or U4880 (N_4880,In_1922,In_341);
xnor U4881 (N_4881,In_2334,In_1518);
and U4882 (N_4882,In_940,In_155);
or U4883 (N_4883,In_1574,In_2461);
nor U4884 (N_4884,In_618,In_2494);
nor U4885 (N_4885,In_1205,In_72);
or U4886 (N_4886,In_1102,In_691);
nor U4887 (N_4887,In_317,In_1051);
or U4888 (N_4888,In_2093,In_1245);
and U4889 (N_4889,In_402,In_596);
or U4890 (N_4890,In_1319,In_2137);
or U4891 (N_4891,In_1073,In_1917);
nand U4892 (N_4892,In_1490,In_506);
nand U4893 (N_4893,In_2440,In_1472);
or U4894 (N_4894,In_1068,In_1052);
xor U4895 (N_4895,In_646,In_1562);
nand U4896 (N_4896,In_1043,In_1718);
or U4897 (N_4897,In_1780,In_155);
or U4898 (N_4898,In_1707,In_959);
and U4899 (N_4899,In_2373,In_1680);
or U4900 (N_4900,In_215,In_431);
or U4901 (N_4901,In_1339,In_1592);
nor U4902 (N_4902,In_985,In_1452);
or U4903 (N_4903,In_907,In_1007);
and U4904 (N_4904,In_1675,In_29);
nand U4905 (N_4905,In_1569,In_817);
nor U4906 (N_4906,In_218,In_2393);
xor U4907 (N_4907,In_2076,In_443);
and U4908 (N_4908,In_298,In_604);
or U4909 (N_4909,In_451,In_741);
xnor U4910 (N_4910,In_1506,In_1488);
xnor U4911 (N_4911,In_1541,In_2473);
nor U4912 (N_4912,In_1583,In_516);
xnor U4913 (N_4913,In_962,In_681);
nand U4914 (N_4914,In_838,In_2395);
and U4915 (N_4915,In_1009,In_1079);
or U4916 (N_4916,In_147,In_1758);
or U4917 (N_4917,In_1591,In_20);
nor U4918 (N_4918,In_1267,In_1198);
nor U4919 (N_4919,In_1250,In_2037);
nand U4920 (N_4920,In_97,In_25);
or U4921 (N_4921,In_1863,In_2281);
or U4922 (N_4922,In_1521,In_2012);
and U4923 (N_4923,In_2406,In_66);
or U4924 (N_4924,In_1381,In_1823);
or U4925 (N_4925,In_1131,In_110);
or U4926 (N_4926,In_2301,In_1791);
or U4927 (N_4927,In_2178,In_34);
xnor U4928 (N_4928,In_1373,In_415);
or U4929 (N_4929,In_1112,In_1660);
nor U4930 (N_4930,In_892,In_2333);
nor U4931 (N_4931,In_199,In_555);
or U4932 (N_4932,In_919,In_1803);
nand U4933 (N_4933,In_2268,In_287);
nand U4934 (N_4934,In_57,In_933);
xnor U4935 (N_4935,In_1378,In_48);
nand U4936 (N_4936,In_2317,In_2495);
xor U4937 (N_4937,In_1174,In_906);
nor U4938 (N_4938,In_2260,In_714);
and U4939 (N_4939,In_2081,In_592);
nor U4940 (N_4940,In_1268,In_512);
and U4941 (N_4941,In_255,In_1654);
xnor U4942 (N_4942,In_622,In_861);
nand U4943 (N_4943,In_815,In_827);
and U4944 (N_4944,In_2335,In_2211);
or U4945 (N_4945,In_2028,In_1996);
or U4946 (N_4946,In_1397,In_2411);
and U4947 (N_4947,In_2467,In_987);
nand U4948 (N_4948,In_2438,In_1344);
or U4949 (N_4949,In_2173,In_917);
nand U4950 (N_4950,In_729,In_1588);
nor U4951 (N_4951,In_2432,In_738);
or U4952 (N_4952,In_1611,In_11);
or U4953 (N_4953,In_950,In_277);
or U4954 (N_4954,In_2312,In_2248);
xor U4955 (N_4955,In_260,In_754);
nand U4956 (N_4956,In_1079,In_535);
nor U4957 (N_4957,In_2336,In_1113);
and U4958 (N_4958,In_1166,In_1402);
or U4959 (N_4959,In_197,In_2292);
or U4960 (N_4960,In_2456,In_1049);
nand U4961 (N_4961,In_2209,In_223);
or U4962 (N_4962,In_804,In_1359);
xor U4963 (N_4963,In_1593,In_1117);
xnor U4964 (N_4964,In_154,In_1632);
nor U4965 (N_4965,In_1117,In_1490);
nand U4966 (N_4966,In_2399,In_1584);
nand U4967 (N_4967,In_2044,In_556);
and U4968 (N_4968,In_162,In_581);
and U4969 (N_4969,In_786,In_1381);
nand U4970 (N_4970,In_209,In_225);
nand U4971 (N_4971,In_662,In_1859);
nor U4972 (N_4972,In_416,In_2415);
nor U4973 (N_4973,In_1014,In_1232);
nor U4974 (N_4974,In_1435,In_2364);
nand U4975 (N_4975,In_2082,In_1092);
or U4976 (N_4976,In_260,In_292);
or U4977 (N_4977,In_1440,In_1618);
and U4978 (N_4978,In_1945,In_1629);
or U4979 (N_4979,In_1048,In_1307);
nor U4980 (N_4980,In_1339,In_2447);
xor U4981 (N_4981,In_1472,In_1877);
xor U4982 (N_4982,In_2237,In_1947);
and U4983 (N_4983,In_678,In_831);
nand U4984 (N_4984,In_1781,In_1981);
nand U4985 (N_4985,In_275,In_832);
nor U4986 (N_4986,In_2355,In_2180);
xnor U4987 (N_4987,In_1334,In_1940);
and U4988 (N_4988,In_1539,In_23);
or U4989 (N_4989,In_1866,In_854);
nand U4990 (N_4990,In_933,In_2444);
or U4991 (N_4991,In_557,In_1205);
and U4992 (N_4992,In_1336,In_1191);
nor U4993 (N_4993,In_1614,In_993);
nand U4994 (N_4994,In_569,In_1059);
xnor U4995 (N_4995,In_388,In_672);
or U4996 (N_4996,In_102,In_1391);
xnor U4997 (N_4997,In_1932,In_1525);
xnor U4998 (N_4998,In_1513,In_2003);
nand U4999 (N_4999,In_1954,In_2442);
xor U5000 (N_5000,In_1293,In_1813);
nand U5001 (N_5001,In_1338,In_1642);
nor U5002 (N_5002,In_1143,In_1099);
or U5003 (N_5003,In_2166,In_376);
or U5004 (N_5004,In_354,In_149);
and U5005 (N_5005,In_1528,In_1749);
nand U5006 (N_5006,In_1356,In_861);
nor U5007 (N_5007,In_1050,In_209);
nand U5008 (N_5008,In_788,In_1226);
xnor U5009 (N_5009,In_1953,In_1144);
and U5010 (N_5010,In_499,In_2116);
nand U5011 (N_5011,In_243,In_346);
xor U5012 (N_5012,In_391,In_606);
and U5013 (N_5013,In_443,In_882);
and U5014 (N_5014,In_1779,In_792);
and U5015 (N_5015,In_1087,In_1600);
nand U5016 (N_5016,In_444,In_2163);
xor U5017 (N_5017,In_254,In_813);
nor U5018 (N_5018,In_929,In_2081);
or U5019 (N_5019,In_2411,In_1470);
xnor U5020 (N_5020,In_1516,In_365);
nand U5021 (N_5021,In_173,In_780);
nand U5022 (N_5022,In_1082,In_487);
and U5023 (N_5023,In_993,In_1870);
nor U5024 (N_5024,In_810,In_1787);
nor U5025 (N_5025,In_458,In_625);
nand U5026 (N_5026,In_2241,In_1429);
nand U5027 (N_5027,In_806,In_1572);
xnor U5028 (N_5028,In_2110,In_2185);
or U5029 (N_5029,In_717,In_819);
and U5030 (N_5030,In_2014,In_884);
xnor U5031 (N_5031,In_1245,In_1030);
or U5032 (N_5032,In_209,In_806);
xor U5033 (N_5033,In_1743,In_1992);
or U5034 (N_5034,In_1551,In_1604);
xor U5035 (N_5035,In_1221,In_1235);
xor U5036 (N_5036,In_16,In_2487);
nand U5037 (N_5037,In_1483,In_263);
nor U5038 (N_5038,In_472,In_1446);
xor U5039 (N_5039,In_2053,In_1086);
nor U5040 (N_5040,In_595,In_624);
nor U5041 (N_5041,In_1417,In_1315);
and U5042 (N_5042,In_1212,In_1507);
or U5043 (N_5043,In_380,In_1792);
and U5044 (N_5044,In_1142,In_1055);
or U5045 (N_5045,In_1063,In_1340);
and U5046 (N_5046,In_883,In_369);
nand U5047 (N_5047,In_1614,In_300);
nor U5048 (N_5048,In_595,In_2055);
nor U5049 (N_5049,In_2048,In_711);
xor U5050 (N_5050,In_601,In_1928);
nor U5051 (N_5051,In_870,In_1516);
nand U5052 (N_5052,In_1459,In_823);
or U5053 (N_5053,In_2351,In_1715);
xnor U5054 (N_5054,In_1427,In_1267);
or U5055 (N_5055,In_1144,In_988);
nand U5056 (N_5056,In_1272,In_365);
nand U5057 (N_5057,In_627,In_724);
or U5058 (N_5058,In_32,In_2494);
nor U5059 (N_5059,In_1502,In_1636);
nor U5060 (N_5060,In_2027,In_1651);
and U5061 (N_5061,In_1713,In_1535);
and U5062 (N_5062,In_1844,In_1776);
xnor U5063 (N_5063,In_2376,In_204);
xor U5064 (N_5064,In_1671,In_1778);
nand U5065 (N_5065,In_1000,In_1672);
or U5066 (N_5066,In_47,In_1647);
nand U5067 (N_5067,In_945,In_2255);
nor U5068 (N_5068,In_1827,In_1488);
and U5069 (N_5069,In_2245,In_332);
or U5070 (N_5070,In_236,In_722);
or U5071 (N_5071,In_2442,In_2340);
nor U5072 (N_5072,In_1437,In_2024);
xnor U5073 (N_5073,In_1810,In_2371);
xnor U5074 (N_5074,In_1931,In_741);
or U5075 (N_5075,In_1759,In_2350);
or U5076 (N_5076,In_1843,In_505);
xor U5077 (N_5077,In_319,In_1075);
or U5078 (N_5078,In_721,In_1016);
xnor U5079 (N_5079,In_119,In_1869);
or U5080 (N_5080,In_1411,In_1838);
and U5081 (N_5081,In_31,In_1058);
and U5082 (N_5082,In_2183,In_1672);
nor U5083 (N_5083,In_1954,In_1824);
xor U5084 (N_5084,In_299,In_729);
and U5085 (N_5085,In_754,In_193);
nand U5086 (N_5086,In_583,In_2090);
xnor U5087 (N_5087,In_119,In_747);
nor U5088 (N_5088,In_1583,In_1961);
or U5089 (N_5089,In_1365,In_254);
nor U5090 (N_5090,In_383,In_1132);
or U5091 (N_5091,In_2151,In_2466);
xnor U5092 (N_5092,In_1967,In_2388);
nor U5093 (N_5093,In_1763,In_755);
nor U5094 (N_5094,In_1676,In_277);
or U5095 (N_5095,In_1002,In_178);
and U5096 (N_5096,In_1281,In_128);
nor U5097 (N_5097,In_2393,In_659);
and U5098 (N_5098,In_1503,In_252);
or U5099 (N_5099,In_228,In_979);
nor U5100 (N_5100,In_935,In_1667);
or U5101 (N_5101,In_1730,In_1575);
nand U5102 (N_5102,In_1413,In_757);
xor U5103 (N_5103,In_651,In_765);
or U5104 (N_5104,In_1743,In_137);
nand U5105 (N_5105,In_1704,In_71);
xor U5106 (N_5106,In_1307,In_1691);
nand U5107 (N_5107,In_1788,In_1729);
nor U5108 (N_5108,In_1375,In_1463);
nand U5109 (N_5109,In_2018,In_223);
and U5110 (N_5110,In_1763,In_836);
or U5111 (N_5111,In_848,In_1982);
or U5112 (N_5112,In_1551,In_1451);
and U5113 (N_5113,In_509,In_826);
and U5114 (N_5114,In_1745,In_873);
xor U5115 (N_5115,In_2254,In_1044);
or U5116 (N_5116,In_808,In_513);
nand U5117 (N_5117,In_2458,In_902);
and U5118 (N_5118,In_1488,In_987);
nor U5119 (N_5119,In_79,In_2150);
xor U5120 (N_5120,In_699,In_2267);
and U5121 (N_5121,In_2470,In_1600);
xor U5122 (N_5122,In_438,In_115);
xor U5123 (N_5123,In_1978,In_138);
xor U5124 (N_5124,In_448,In_2002);
xnor U5125 (N_5125,In_853,In_1326);
nor U5126 (N_5126,In_1251,In_460);
xnor U5127 (N_5127,In_1228,In_1603);
nor U5128 (N_5128,In_1606,In_1629);
xnor U5129 (N_5129,In_1983,In_1565);
and U5130 (N_5130,In_1067,In_1814);
nand U5131 (N_5131,In_2236,In_2262);
or U5132 (N_5132,In_899,In_968);
nor U5133 (N_5133,In_1329,In_648);
or U5134 (N_5134,In_2400,In_1846);
nand U5135 (N_5135,In_955,In_816);
nor U5136 (N_5136,In_2419,In_719);
nand U5137 (N_5137,In_1413,In_981);
nand U5138 (N_5138,In_610,In_2018);
or U5139 (N_5139,In_2463,In_1386);
xnor U5140 (N_5140,In_1981,In_367);
nor U5141 (N_5141,In_2427,In_821);
and U5142 (N_5142,In_416,In_1376);
and U5143 (N_5143,In_1135,In_151);
xnor U5144 (N_5144,In_1145,In_1708);
nand U5145 (N_5145,In_1505,In_2202);
and U5146 (N_5146,In_1943,In_493);
or U5147 (N_5147,In_1971,In_1838);
and U5148 (N_5148,In_1002,In_1838);
nand U5149 (N_5149,In_671,In_636);
and U5150 (N_5150,In_1022,In_300);
and U5151 (N_5151,In_598,In_73);
xor U5152 (N_5152,In_1163,In_1262);
nand U5153 (N_5153,In_2461,In_881);
xnor U5154 (N_5154,In_947,In_70);
and U5155 (N_5155,In_1780,In_389);
or U5156 (N_5156,In_1404,In_609);
nand U5157 (N_5157,In_1280,In_1474);
and U5158 (N_5158,In_843,In_1407);
xor U5159 (N_5159,In_2178,In_80);
and U5160 (N_5160,In_2429,In_1651);
or U5161 (N_5161,In_1530,In_574);
or U5162 (N_5162,In_2466,In_1295);
nand U5163 (N_5163,In_388,In_1865);
and U5164 (N_5164,In_1159,In_2338);
and U5165 (N_5165,In_359,In_659);
nor U5166 (N_5166,In_2016,In_407);
or U5167 (N_5167,In_1983,In_1750);
xor U5168 (N_5168,In_1968,In_971);
and U5169 (N_5169,In_1728,In_2284);
nand U5170 (N_5170,In_371,In_95);
nand U5171 (N_5171,In_2045,In_2017);
and U5172 (N_5172,In_2025,In_341);
xnor U5173 (N_5173,In_2218,In_526);
xor U5174 (N_5174,In_2474,In_177);
nor U5175 (N_5175,In_433,In_2294);
nor U5176 (N_5176,In_842,In_1970);
and U5177 (N_5177,In_564,In_1867);
or U5178 (N_5178,In_615,In_326);
xor U5179 (N_5179,In_232,In_433);
xnor U5180 (N_5180,In_22,In_1159);
xor U5181 (N_5181,In_2350,In_2054);
and U5182 (N_5182,In_1521,In_2260);
nor U5183 (N_5183,In_123,In_2481);
or U5184 (N_5184,In_1115,In_565);
nor U5185 (N_5185,In_710,In_1133);
and U5186 (N_5186,In_1382,In_458);
nor U5187 (N_5187,In_1937,In_2448);
and U5188 (N_5188,In_2119,In_1731);
nor U5189 (N_5189,In_1338,In_1957);
or U5190 (N_5190,In_1218,In_165);
nand U5191 (N_5191,In_141,In_1541);
nor U5192 (N_5192,In_1497,In_1811);
nor U5193 (N_5193,In_2493,In_752);
and U5194 (N_5194,In_1014,In_1095);
or U5195 (N_5195,In_2234,In_494);
nand U5196 (N_5196,In_144,In_1166);
xnor U5197 (N_5197,In_1743,In_2326);
and U5198 (N_5198,In_2014,In_680);
and U5199 (N_5199,In_263,In_266);
xor U5200 (N_5200,In_2012,In_423);
nand U5201 (N_5201,In_53,In_2119);
nor U5202 (N_5202,In_1841,In_399);
or U5203 (N_5203,In_1733,In_1265);
nor U5204 (N_5204,In_2001,In_1138);
nand U5205 (N_5205,In_1622,In_1075);
and U5206 (N_5206,In_2044,In_498);
and U5207 (N_5207,In_701,In_596);
and U5208 (N_5208,In_2004,In_1463);
and U5209 (N_5209,In_1078,In_864);
nor U5210 (N_5210,In_621,In_1119);
xor U5211 (N_5211,In_1412,In_1609);
nand U5212 (N_5212,In_105,In_476);
nand U5213 (N_5213,In_1104,In_1150);
xnor U5214 (N_5214,In_1284,In_1858);
or U5215 (N_5215,In_543,In_2100);
nor U5216 (N_5216,In_216,In_1734);
xor U5217 (N_5217,In_902,In_1552);
and U5218 (N_5218,In_265,In_988);
xor U5219 (N_5219,In_737,In_1852);
nand U5220 (N_5220,In_198,In_706);
xor U5221 (N_5221,In_1271,In_1889);
nor U5222 (N_5222,In_1941,In_2074);
nor U5223 (N_5223,In_2069,In_750);
xnor U5224 (N_5224,In_2265,In_587);
and U5225 (N_5225,In_817,In_1769);
nand U5226 (N_5226,In_1907,In_482);
xor U5227 (N_5227,In_85,In_106);
xnor U5228 (N_5228,In_2146,In_1316);
or U5229 (N_5229,In_740,In_2287);
or U5230 (N_5230,In_1810,In_803);
xor U5231 (N_5231,In_1015,In_1455);
nand U5232 (N_5232,In_343,In_2135);
nand U5233 (N_5233,In_782,In_1540);
nor U5234 (N_5234,In_5,In_261);
nand U5235 (N_5235,In_324,In_1878);
nor U5236 (N_5236,In_1207,In_2381);
xnor U5237 (N_5237,In_1852,In_77);
nand U5238 (N_5238,In_719,In_1468);
xor U5239 (N_5239,In_806,In_2303);
nand U5240 (N_5240,In_2191,In_327);
or U5241 (N_5241,In_1606,In_1679);
or U5242 (N_5242,In_1692,In_456);
nand U5243 (N_5243,In_2155,In_493);
xnor U5244 (N_5244,In_1184,In_1080);
and U5245 (N_5245,In_1254,In_2171);
nor U5246 (N_5246,In_1592,In_2479);
and U5247 (N_5247,In_1478,In_651);
nor U5248 (N_5248,In_1958,In_1310);
nor U5249 (N_5249,In_748,In_474);
nand U5250 (N_5250,In_908,In_658);
and U5251 (N_5251,In_2286,In_1398);
nand U5252 (N_5252,In_2312,In_742);
nand U5253 (N_5253,In_1404,In_2163);
or U5254 (N_5254,In_2214,In_1592);
or U5255 (N_5255,In_2187,In_2259);
xnor U5256 (N_5256,In_1292,In_851);
and U5257 (N_5257,In_1447,In_933);
or U5258 (N_5258,In_1080,In_474);
nor U5259 (N_5259,In_1614,In_1477);
xnor U5260 (N_5260,In_577,In_97);
and U5261 (N_5261,In_1512,In_663);
nor U5262 (N_5262,In_142,In_241);
xnor U5263 (N_5263,In_1008,In_1211);
and U5264 (N_5264,In_1411,In_768);
and U5265 (N_5265,In_2121,In_215);
nand U5266 (N_5266,In_641,In_2054);
xor U5267 (N_5267,In_1116,In_487);
nor U5268 (N_5268,In_310,In_1125);
or U5269 (N_5269,In_534,In_437);
nand U5270 (N_5270,In_449,In_2252);
xnor U5271 (N_5271,In_2390,In_2148);
nor U5272 (N_5272,In_97,In_1952);
and U5273 (N_5273,In_2316,In_964);
or U5274 (N_5274,In_1396,In_622);
nand U5275 (N_5275,In_781,In_315);
nor U5276 (N_5276,In_2214,In_1126);
and U5277 (N_5277,In_1275,In_253);
nor U5278 (N_5278,In_297,In_1847);
nand U5279 (N_5279,In_1811,In_1007);
and U5280 (N_5280,In_966,In_2292);
or U5281 (N_5281,In_385,In_245);
nand U5282 (N_5282,In_899,In_2477);
and U5283 (N_5283,In_414,In_1815);
or U5284 (N_5284,In_860,In_1406);
nor U5285 (N_5285,In_2447,In_1299);
and U5286 (N_5286,In_1287,In_1478);
xor U5287 (N_5287,In_2163,In_1062);
or U5288 (N_5288,In_2082,In_500);
or U5289 (N_5289,In_467,In_678);
xor U5290 (N_5290,In_718,In_1121);
and U5291 (N_5291,In_1725,In_1655);
and U5292 (N_5292,In_862,In_815);
xnor U5293 (N_5293,In_273,In_1656);
nor U5294 (N_5294,In_810,In_1645);
or U5295 (N_5295,In_1405,In_2345);
nor U5296 (N_5296,In_1254,In_535);
and U5297 (N_5297,In_704,In_1469);
nand U5298 (N_5298,In_159,In_1131);
nand U5299 (N_5299,In_1733,In_942);
or U5300 (N_5300,In_1894,In_1902);
or U5301 (N_5301,In_541,In_13);
nor U5302 (N_5302,In_1496,In_1759);
and U5303 (N_5303,In_803,In_2094);
nand U5304 (N_5304,In_235,In_1464);
nor U5305 (N_5305,In_1332,In_1830);
nor U5306 (N_5306,In_1731,In_1993);
nand U5307 (N_5307,In_401,In_1397);
or U5308 (N_5308,In_388,In_828);
or U5309 (N_5309,In_2351,In_2246);
or U5310 (N_5310,In_1415,In_1873);
xor U5311 (N_5311,In_1080,In_1166);
or U5312 (N_5312,In_2204,In_1679);
xor U5313 (N_5313,In_135,In_1014);
xnor U5314 (N_5314,In_833,In_251);
nand U5315 (N_5315,In_1823,In_110);
or U5316 (N_5316,In_1248,In_1412);
xnor U5317 (N_5317,In_963,In_1422);
or U5318 (N_5318,In_525,In_2303);
xor U5319 (N_5319,In_2188,In_1324);
nand U5320 (N_5320,In_1026,In_1360);
nor U5321 (N_5321,In_388,In_584);
nand U5322 (N_5322,In_2253,In_927);
xor U5323 (N_5323,In_2430,In_546);
or U5324 (N_5324,In_2047,In_528);
and U5325 (N_5325,In_656,In_1963);
nor U5326 (N_5326,In_1221,In_846);
xnor U5327 (N_5327,In_335,In_701);
nand U5328 (N_5328,In_2358,In_2172);
or U5329 (N_5329,In_2385,In_926);
nor U5330 (N_5330,In_755,In_1954);
or U5331 (N_5331,In_2431,In_573);
or U5332 (N_5332,In_1545,In_2221);
or U5333 (N_5333,In_628,In_2451);
nor U5334 (N_5334,In_498,In_1811);
and U5335 (N_5335,In_1678,In_1504);
or U5336 (N_5336,In_493,In_1762);
and U5337 (N_5337,In_2139,In_2362);
and U5338 (N_5338,In_547,In_1517);
nor U5339 (N_5339,In_1541,In_1141);
nand U5340 (N_5340,In_145,In_2307);
nor U5341 (N_5341,In_595,In_1294);
nor U5342 (N_5342,In_248,In_873);
or U5343 (N_5343,In_1399,In_2420);
and U5344 (N_5344,In_913,In_1346);
nand U5345 (N_5345,In_2181,In_1603);
or U5346 (N_5346,In_1869,In_1017);
nor U5347 (N_5347,In_795,In_358);
nand U5348 (N_5348,In_451,In_221);
and U5349 (N_5349,In_1699,In_1776);
xor U5350 (N_5350,In_1877,In_2276);
xor U5351 (N_5351,In_338,In_1825);
nand U5352 (N_5352,In_2259,In_2273);
xnor U5353 (N_5353,In_1336,In_1237);
nand U5354 (N_5354,In_728,In_1144);
or U5355 (N_5355,In_851,In_1829);
and U5356 (N_5356,In_934,In_2230);
and U5357 (N_5357,In_809,In_1285);
and U5358 (N_5358,In_784,In_61);
xnor U5359 (N_5359,In_997,In_792);
or U5360 (N_5360,In_541,In_1154);
or U5361 (N_5361,In_1306,In_2435);
nand U5362 (N_5362,In_861,In_345);
xnor U5363 (N_5363,In_1967,In_1485);
xor U5364 (N_5364,In_2249,In_348);
xor U5365 (N_5365,In_1310,In_1553);
nor U5366 (N_5366,In_155,In_1263);
and U5367 (N_5367,In_2051,In_2084);
nor U5368 (N_5368,In_1625,In_1337);
nor U5369 (N_5369,In_1137,In_2239);
xnor U5370 (N_5370,In_1026,In_1837);
and U5371 (N_5371,In_967,In_2473);
or U5372 (N_5372,In_1701,In_2414);
or U5373 (N_5373,In_1979,In_1179);
nor U5374 (N_5374,In_27,In_949);
nor U5375 (N_5375,In_303,In_1826);
and U5376 (N_5376,In_1550,In_2490);
and U5377 (N_5377,In_2092,In_2019);
nor U5378 (N_5378,In_711,In_653);
nand U5379 (N_5379,In_1287,In_1102);
and U5380 (N_5380,In_2250,In_881);
and U5381 (N_5381,In_78,In_2282);
nand U5382 (N_5382,In_1782,In_841);
or U5383 (N_5383,In_1524,In_241);
nor U5384 (N_5384,In_779,In_101);
nor U5385 (N_5385,In_271,In_1839);
and U5386 (N_5386,In_1438,In_611);
or U5387 (N_5387,In_435,In_1783);
xnor U5388 (N_5388,In_1650,In_352);
xor U5389 (N_5389,In_1200,In_400);
or U5390 (N_5390,In_871,In_1732);
nor U5391 (N_5391,In_1482,In_1690);
nor U5392 (N_5392,In_1391,In_1298);
nor U5393 (N_5393,In_751,In_1132);
nand U5394 (N_5394,In_2239,In_1036);
nor U5395 (N_5395,In_1394,In_1583);
nand U5396 (N_5396,In_308,In_2444);
nor U5397 (N_5397,In_1585,In_1049);
nor U5398 (N_5398,In_354,In_734);
xor U5399 (N_5399,In_849,In_318);
nand U5400 (N_5400,In_240,In_1973);
or U5401 (N_5401,In_587,In_1664);
and U5402 (N_5402,In_2070,In_558);
xnor U5403 (N_5403,In_769,In_851);
xor U5404 (N_5404,In_234,In_132);
or U5405 (N_5405,In_319,In_529);
or U5406 (N_5406,In_1619,In_1223);
and U5407 (N_5407,In_1302,In_2099);
xnor U5408 (N_5408,In_2131,In_192);
and U5409 (N_5409,In_122,In_1264);
nand U5410 (N_5410,In_161,In_2374);
or U5411 (N_5411,In_500,In_1279);
nor U5412 (N_5412,In_831,In_1063);
nor U5413 (N_5413,In_1994,In_2042);
and U5414 (N_5414,In_157,In_787);
or U5415 (N_5415,In_713,In_1417);
or U5416 (N_5416,In_1798,In_2001);
xor U5417 (N_5417,In_2172,In_1258);
nand U5418 (N_5418,In_690,In_1958);
nand U5419 (N_5419,In_2426,In_1769);
or U5420 (N_5420,In_1961,In_2154);
xnor U5421 (N_5421,In_1625,In_1760);
and U5422 (N_5422,In_1446,In_2449);
or U5423 (N_5423,In_1910,In_1811);
nand U5424 (N_5424,In_41,In_1757);
nor U5425 (N_5425,In_993,In_2226);
xor U5426 (N_5426,In_383,In_1383);
and U5427 (N_5427,In_1318,In_2385);
xor U5428 (N_5428,In_853,In_950);
nor U5429 (N_5429,In_1469,In_623);
nand U5430 (N_5430,In_10,In_1305);
nor U5431 (N_5431,In_387,In_2092);
nor U5432 (N_5432,In_884,In_1670);
and U5433 (N_5433,In_318,In_435);
nand U5434 (N_5434,In_2073,In_1213);
or U5435 (N_5435,In_870,In_837);
nand U5436 (N_5436,In_1232,In_1871);
nand U5437 (N_5437,In_522,In_1713);
and U5438 (N_5438,In_136,In_700);
and U5439 (N_5439,In_2177,In_1884);
nor U5440 (N_5440,In_1725,In_1439);
nor U5441 (N_5441,In_1514,In_120);
and U5442 (N_5442,In_1938,In_1978);
and U5443 (N_5443,In_2472,In_373);
xnor U5444 (N_5444,In_1711,In_462);
nor U5445 (N_5445,In_710,In_913);
and U5446 (N_5446,In_2246,In_129);
and U5447 (N_5447,In_1465,In_1670);
xnor U5448 (N_5448,In_1363,In_956);
nor U5449 (N_5449,In_1603,In_1708);
or U5450 (N_5450,In_2344,In_1762);
nor U5451 (N_5451,In_1930,In_754);
xnor U5452 (N_5452,In_2246,In_1557);
nand U5453 (N_5453,In_1889,In_475);
and U5454 (N_5454,In_390,In_473);
nor U5455 (N_5455,In_1528,In_2053);
nand U5456 (N_5456,In_1008,In_1343);
xor U5457 (N_5457,In_850,In_1366);
or U5458 (N_5458,In_830,In_960);
or U5459 (N_5459,In_755,In_2413);
nand U5460 (N_5460,In_218,In_718);
and U5461 (N_5461,In_219,In_2081);
and U5462 (N_5462,In_466,In_1548);
nand U5463 (N_5463,In_148,In_97);
nor U5464 (N_5464,In_912,In_1581);
or U5465 (N_5465,In_896,In_1565);
xor U5466 (N_5466,In_745,In_1699);
and U5467 (N_5467,In_750,In_1966);
or U5468 (N_5468,In_2094,In_554);
nor U5469 (N_5469,In_2204,In_1358);
or U5470 (N_5470,In_2028,In_1064);
nand U5471 (N_5471,In_1990,In_1475);
nand U5472 (N_5472,In_659,In_365);
or U5473 (N_5473,In_1629,In_758);
or U5474 (N_5474,In_504,In_1158);
xor U5475 (N_5475,In_165,In_986);
and U5476 (N_5476,In_2021,In_1214);
or U5477 (N_5477,In_1399,In_2299);
nand U5478 (N_5478,In_1258,In_1971);
nand U5479 (N_5479,In_1951,In_1957);
or U5480 (N_5480,In_1909,In_1230);
and U5481 (N_5481,In_2191,In_1260);
and U5482 (N_5482,In_1061,In_331);
xor U5483 (N_5483,In_1490,In_1523);
nor U5484 (N_5484,In_1124,In_1840);
nand U5485 (N_5485,In_2176,In_1347);
and U5486 (N_5486,In_1010,In_1340);
nand U5487 (N_5487,In_2411,In_1442);
xnor U5488 (N_5488,In_296,In_2470);
nand U5489 (N_5489,In_1313,In_590);
nand U5490 (N_5490,In_2289,In_1205);
or U5491 (N_5491,In_1396,In_2169);
and U5492 (N_5492,In_1147,In_2087);
nand U5493 (N_5493,In_1197,In_2302);
xor U5494 (N_5494,In_1644,In_1954);
nand U5495 (N_5495,In_1274,In_348);
nor U5496 (N_5496,In_1442,In_115);
nand U5497 (N_5497,In_1779,In_441);
nor U5498 (N_5498,In_383,In_1146);
nor U5499 (N_5499,In_856,In_2407);
nor U5500 (N_5500,In_146,In_1262);
xor U5501 (N_5501,In_78,In_1262);
and U5502 (N_5502,In_1268,In_384);
or U5503 (N_5503,In_1693,In_759);
nand U5504 (N_5504,In_391,In_1322);
nand U5505 (N_5505,In_1890,In_1369);
or U5506 (N_5506,In_484,In_937);
nor U5507 (N_5507,In_2211,In_1778);
and U5508 (N_5508,In_707,In_83);
nor U5509 (N_5509,In_1749,In_1907);
nor U5510 (N_5510,In_2049,In_456);
nand U5511 (N_5511,In_2415,In_127);
xnor U5512 (N_5512,In_603,In_784);
or U5513 (N_5513,In_1303,In_2384);
xor U5514 (N_5514,In_1627,In_486);
or U5515 (N_5515,In_404,In_1657);
nand U5516 (N_5516,In_481,In_2490);
nand U5517 (N_5517,In_413,In_1682);
nand U5518 (N_5518,In_2375,In_397);
or U5519 (N_5519,In_680,In_225);
nand U5520 (N_5520,In_1076,In_2206);
nor U5521 (N_5521,In_591,In_2089);
or U5522 (N_5522,In_2324,In_104);
and U5523 (N_5523,In_2476,In_563);
or U5524 (N_5524,In_1230,In_879);
xnor U5525 (N_5525,In_532,In_2355);
xor U5526 (N_5526,In_570,In_2395);
nor U5527 (N_5527,In_496,In_1253);
xnor U5528 (N_5528,In_1475,In_1482);
and U5529 (N_5529,In_1327,In_2098);
nand U5530 (N_5530,In_370,In_2228);
xnor U5531 (N_5531,In_836,In_363);
xnor U5532 (N_5532,In_127,In_935);
and U5533 (N_5533,In_1203,In_919);
xor U5534 (N_5534,In_1352,In_1426);
nand U5535 (N_5535,In_2251,In_2204);
and U5536 (N_5536,In_1591,In_2109);
xnor U5537 (N_5537,In_1239,In_4);
and U5538 (N_5538,In_267,In_163);
nand U5539 (N_5539,In_2167,In_885);
xor U5540 (N_5540,In_1634,In_1729);
nand U5541 (N_5541,In_1400,In_2209);
xor U5542 (N_5542,In_1877,In_1035);
nand U5543 (N_5543,In_78,In_94);
xor U5544 (N_5544,In_1345,In_2278);
nand U5545 (N_5545,In_2010,In_1112);
and U5546 (N_5546,In_1701,In_493);
nor U5547 (N_5547,In_1312,In_2329);
xor U5548 (N_5548,In_1689,In_1041);
and U5549 (N_5549,In_686,In_1211);
and U5550 (N_5550,In_2466,In_163);
nand U5551 (N_5551,In_274,In_1306);
and U5552 (N_5552,In_1845,In_2297);
nor U5553 (N_5553,In_723,In_56);
nor U5554 (N_5554,In_621,In_37);
or U5555 (N_5555,In_1126,In_1795);
or U5556 (N_5556,In_1599,In_861);
xor U5557 (N_5557,In_77,In_675);
nor U5558 (N_5558,In_1577,In_1912);
or U5559 (N_5559,In_1055,In_2103);
or U5560 (N_5560,In_741,In_1804);
nand U5561 (N_5561,In_1847,In_1257);
and U5562 (N_5562,In_931,In_1592);
xnor U5563 (N_5563,In_2223,In_736);
xnor U5564 (N_5564,In_462,In_1612);
nor U5565 (N_5565,In_1503,In_1315);
and U5566 (N_5566,In_1909,In_2265);
or U5567 (N_5567,In_1513,In_1847);
and U5568 (N_5568,In_1945,In_950);
xor U5569 (N_5569,In_1248,In_49);
nor U5570 (N_5570,In_710,In_222);
or U5571 (N_5571,In_134,In_654);
and U5572 (N_5572,In_1715,In_91);
and U5573 (N_5573,In_1334,In_217);
nand U5574 (N_5574,In_2476,In_225);
and U5575 (N_5575,In_2423,In_65);
nor U5576 (N_5576,In_1476,In_1593);
nand U5577 (N_5577,In_1510,In_1456);
nand U5578 (N_5578,In_1046,In_948);
nand U5579 (N_5579,In_1240,In_2462);
nand U5580 (N_5580,In_2150,In_913);
and U5581 (N_5581,In_982,In_527);
nand U5582 (N_5582,In_652,In_567);
and U5583 (N_5583,In_1339,In_625);
nand U5584 (N_5584,In_494,In_1475);
nand U5585 (N_5585,In_1112,In_1444);
and U5586 (N_5586,In_326,In_1043);
xnor U5587 (N_5587,In_1892,In_268);
nand U5588 (N_5588,In_703,In_1331);
or U5589 (N_5589,In_322,In_223);
xnor U5590 (N_5590,In_518,In_1687);
nand U5591 (N_5591,In_2462,In_1168);
and U5592 (N_5592,In_2232,In_1234);
nand U5593 (N_5593,In_310,In_1541);
nand U5594 (N_5594,In_1245,In_2251);
or U5595 (N_5595,In_601,In_952);
nand U5596 (N_5596,In_274,In_2450);
or U5597 (N_5597,In_1540,In_2309);
or U5598 (N_5598,In_2264,In_1164);
and U5599 (N_5599,In_785,In_2099);
nor U5600 (N_5600,In_504,In_1376);
or U5601 (N_5601,In_701,In_339);
or U5602 (N_5602,In_1727,In_1403);
or U5603 (N_5603,In_56,In_403);
and U5604 (N_5604,In_1704,In_1837);
nor U5605 (N_5605,In_455,In_1527);
xnor U5606 (N_5606,In_1910,In_465);
or U5607 (N_5607,In_2340,In_2093);
nor U5608 (N_5608,In_1695,In_2227);
xor U5609 (N_5609,In_1503,In_643);
nand U5610 (N_5610,In_824,In_961);
and U5611 (N_5611,In_945,In_2205);
nor U5612 (N_5612,In_1372,In_461);
xor U5613 (N_5613,In_48,In_272);
and U5614 (N_5614,In_101,In_2410);
and U5615 (N_5615,In_396,In_2352);
and U5616 (N_5616,In_107,In_372);
xor U5617 (N_5617,In_1923,In_1122);
or U5618 (N_5618,In_1267,In_152);
nand U5619 (N_5619,In_1308,In_1599);
nand U5620 (N_5620,In_867,In_2128);
or U5621 (N_5621,In_1101,In_1571);
and U5622 (N_5622,In_482,In_373);
and U5623 (N_5623,In_867,In_82);
and U5624 (N_5624,In_2042,In_654);
or U5625 (N_5625,In_1103,In_410);
xnor U5626 (N_5626,In_549,In_405);
and U5627 (N_5627,In_1351,In_1363);
or U5628 (N_5628,In_1404,In_1071);
xor U5629 (N_5629,In_1020,In_375);
nor U5630 (N_5630,In_1776,In_1891);
or U5631 (N_5631,In_1778,In_1780);
or U5632 (N_5632,In_1635,In_2297);
nand U5633 (N_5633,In_2147,In_488);
nor U5634 (N_5634,In_714,In_653);
or U5635 (N_5635,In_353,In_528);
xnor U5636 (N_5636,In_1261,In_1738);
nor U5637 (N_5637,In_967,In_2461);
and U5638 (N_5638,In_9,In_224);
nand U5639 (N_5639,In_428,In_1665);
or U5640 (N_5640,In_329,In_1542);
nor U5641 (N_5641,In_6,In_2152);
and U5642 (N_5642,In_2396,In_742);
nand U5643 (N_5643,In_128,In_2238);
or U5644 (N_5644,In_1193,In_1741);
nand U5645 (N_5645,In_2120,In_2435);
and U5646 (N_5646,In_622,In_2492);
or U5647 (N_5647,In_1171,In_109);
xor U5648 (N_5648,In_111,In_202);
nor U5649 (N_5649,In_2454,In_270);
nand U5650 (N_5650,In_358,In_1489);
nand U5651 (N_5651,In_1891,In_1040);
nand U5652 (N_5652,In_2424,In_419);
nor U5653 (N_5653,In_2069,In_517);
or U5654 (N_5654,In_1122,In_715);
and U5655 (N_5655,In_60,In_2106);
nor U5656 (N_5656,In_6,In_2038);
xor U5657 (N_5657,In_915,In_1945);
xnor U5658 (N_5658,In_1428,In_436);
xor U5659 (N_5659,In_2499,In_2073);
or U5660 (N_5660,In_1670,In_1349);
xor U5661 (N_5661,In_2420,In_1803);
nand U5662 (N_5662,In_1849,In_376);
or U5663 (N_5663,In_1148,In_2037);
nor U5664 (N_5664,In_2437,In_1080);
nand U5665 (N_5665,In_420,In_1240);
xnor U5666 (N_5666,In_666,In_888);
nand U5667 (N_5667,In_2184,In_529);
xnor U5668 (N_5668,In_396,In_2291);
and U5669 (N_5669,In_955,In_1470);
xor U5670 (N_5670,In_1271,In_2160);
nand U5671 (N_5671,In_406,In_2432);
xor U5672 (N_5672,In_1707,In_1229);
nand U5673 (N_5673,In_1551,In_31);
nor U5674 (N_5674,In_2088,In_793);
or U5675 (N_5675,In_1231,In_1606);
nor U5676 (N_5676,In_419,In_295);
nor U5677 (N_5677,In_1265,In_862);
or U5678 (N_5678,In_2196,In_968);
nand U5679 (N_5679,In_898,In_2147);
or U5680 (N_5680,In_404,In_1621);
or U5681 (N_5681,In_330,In_2402);
nand U5682 (N_5682,In_224,In_2027);
nor U5683 (N_5683,In_2264,In_1312);
xnor U5684 (N_5684,In_1792,In_2273);
and U5685 (N_5685,In_409,In_167);
or U5686 (N_5686,In_1883,In_92);
xnor U5687 (N_5687,In_2182,In_1953);
and U5688 (N_5688,In_1165,In_1979);
or U5689 (N_5689,In_183,In_2006);
xor U5690 (N_5690,In_580,In_2139);
xnor U5691 (N_5691,In_1762,In_2244);
nand U5692 (N_5692,In_398,In_167);
or U5693 (N_5693,In_2370,In_170);
nor U5694 (N_5694,In_2236,In_2127);
xnor U5695 (N_5695,In_427,In_2266);
nor U5696 (N_5696,In_1021,In_2418);
nor U5697 (N_5697,In_1089,In_52);
nand U5698 (N_5698,In_1548,In_478);
or U5699 (N_5699,In_147,In_2436);
xnor U5700 (N_5700,In_2372,In_359);
nor U5701 (N_5701,In_1821,In_1846);
and U5702 (N_5702,In_1092,In_589);
nor U5703 (N_5703,In_1573,In_2131);
or U5704 (N_5704,In_463,In_1323);
and U5705 (N_5705,In_302,In_231);
and U5706 (N_5706,In_2120,In_739);
or U5707 (N_5707,In_2383,In_2320);
or U5708 (N_5708,In_2113,In_2473);
xor U5709 (N_5709,In_1128,In_1959);
or U5710 (N_5710,In_1997,In_1295);
nor U5711 (N_5711,In_1618,In_2348);
nor U5712 (N_5712,In_75,In_232);
and U5713 (N_5713,In_962,In_1244);
xor U5714 (N_5714,In_2435,In_1639);
nor U5715 (N_5715,In_1938,In_333);
nand U5716 (N_5716,In_44,In_1137);
xor U5717 (N_5717,In_1610,In_856);
or U5718 (N_5718,In_2456,In_1350);
or U5719 (N_5719,In_2047,In_2290);
nor U5720 (N_5720,In_549,In_1712);
or U5721 (N_5721,In_547,In_1683);
nand U5722 (N_5722,In_1492,In_1419);
or U5723 (N_5723,In_2281,In_662);
nand U5724 (N_5724,In_1559,In_1699);
nor U5725 (N_5725,In_1260,In_1665);
xor U5726 (N_5726,In_1881,In_1381);
or U5727 (N_5727,In_2156,In_1098);
nand U5728 (N_5728,In_735,In_864);
xor U5729 (N_5729,In_1740,In_390);
nor U5730 (N_5730,In_1400,In_82);
and U5731 (N_5731,In_2382,In_253);
nand U5732 (N_5732,In_2012,In_919);
xor U5733 (N_5733,In_1062,In_1743);
xor U5734 (N_5734,In_1732,In_397);
and U5735 (N_5735,In_2431,In_2097);
and U5736 (N_5736,In_2002,In_911);
and U5737 (N_5737,In_772,In_667);
and U5738 (N_5738,In_2275,In_2472);
nor U5739 (N_5739,In_1236,In_193);
nor U5740 (N_5740,In_2124,In_1265);
xor U5741 (N_5741,In_24,In_1408);
nand U5742 (N_5742,In_907,In_870);
or U5743 (N_5743,In_1182,In_270);
nor U5744 (N_5744,In_1228,In_2149);
nor U5745 (N_5745,In_1135,In_2435);
nand U5746 (N_5746,In_513,In_286);
xor U5747 (N_5747,In_716,In_1411);
nor U5748 (N_5748,In_1761,In_1365);
xnor U5749 (N_5749,In_2314,In_2015);
or U5750 (N_5750,In_1002,In_2422);
nor U5751 (N_5751,In_491,In_1375);
nand U5752 (N_5752,In_1988,In_894);
and U5753 (N_5753,In_875,In_2129);
xor U5754 (N_5754,In_1498,In_1493);
and U5755 (N_5755,In_1843,In_722);
nand U5756 (N_5756,In_2136,In_2417);
and U5757 (N_5757,In_721,In_2467);
or U5758 (N_5758,In_1272,In_2477);
or U5759 (N_5759,In_23,In_2073);
xor U5760 (N_5760,In_4,In_20);
nand U5761 (N_5761,In_931,In_1266);
and U5762 (N_5762,In_1628,In_877);
nand U5763 (N_5763,In_2065,In_273);
nor U5764 (N_5764,In_1187,In_32);
nor U5765 (N_5765,In_2209,In_1448);
nor U5766 (N_5766,In_1506,In_2290);
or U5767 (N_5767,In_682,In_753);
xor U5768 (N_5768,In_505,In_2427);
nor U5769 (N_5769,In_1677,In_1382);
nor U5770 (N_5770,In_1906,In_2395);
and U5771 (N_5771,In_1125,In_984);
nand U5772 (N_5772,In_424,In_993);
nand U5773 (N_5773,In_527,In_2474);
or U5774 (N_5774,In_2172,In_1352);
nand U5775 (N_5775,In_1808,In_850);
nor U5776 (N_5776,In_1103,In_801);
or U5777 (N_5777,In_2376,In_441);
nand U5778 (N_5778,In_2433,In_654);
xnor U5779 (N_5779,In_1370,In_717);
xor U5780 (N_5780,In_1138,In_579);
nand U5781 (N_5781,In_1621,In_385);
and U5782 (N_5782,In_1209,In_2038);
and U5783 (N_5783,In_1033,In_2360);
or U5784 (N_5784,In_381,In_221);
nand U5785 (N_5785,In_427,In_2);
xor U5786 (N_5786,In_2060,In_660);
or U5787 (N_5787,In_1490,In_1434);
xnor U5788 (N_5788,In_1887,In_11);
nor U5789 (N_5789,In_582,In_626);
or U5790 (N_5790,In_1881,In_1766);
xor U5791 (N_5791,In_910,In_2190);
and U5792 (N_5792,In_2303,In_1276);
and U5793 (N_5793,In_775,In_1287);
xor U5794 (N_5794,In_73,In_492);
xor U5795 (N_5795,In_1308,In_601);
nand U5796 (N_5796,In_1852,In_534);
or U5797 (N_5797,In_1828,In_1878);
or U5798 (N_5798,In_811,In_516);
or U5799 (N_5799,In_444,In_1869);
nand U5800 (N_5800,In_118,In_1633);
and U5801 (N_5801,In_1727,In_1388);
nand U5802 (N_5802,In_47,In_1692);
nor U5803 (N_5803,In_1521,In_147);
nor U5804 (N_5804,In_1231,In_873);
or U5805 (N_5805,In_1743,In_702);
nor U5806 (N_5806,In_487,In_915);
nand U5807 (N_5807,In_1338,In_1801);
xnor U5808 (N_5808,In_658,In_1242);
nand U5809 (N_5809,In_302,In_1352);
nand U5810 (N_5810,In_923,In_1638);
nand U5811 (N_5811,In_1242,In_895);
nand U5812 (N_5812,In_2078,In_2247);
xnor U5813 (N_5813,In_688,In_1631);
xnor U5814 (N_5814,In_1818,In_2244);
xnor U5815 (N_5815,In_1234,In_279);
xnor U5816 (N_5816,In_2091,In_457);
and U5817 (N_5817,In_1354,In_546);
nand U5818 (N_5818,In_252,In_907);
nand U5819 (N_5819,In_2456,In_1110);
or U5820 (N_5820,In_46,In_1157);
or U5821 (N_5821,In_1374,In_29);
xor U5822 (N_5822,In_1299,In_645);
xnor U5823 (N_5823,In_793,In_314);
xor U5824 (N_5824,In_2321,In_1527);
or U5825 (N_5825,In_504,In_2374);
xnor U5826 (N_5826,In_1944,In_79);
or U5827 (N_5827,In_2401,In_1630);
or U5828 (N_5828,In_1284,In_1401);
nor U5829 (N_5829,In_646,In_1024);
and U5830 (N_5830,In_1397,In_2);
or U5831 (N_5831,In_1384,In_106);
and U5832 (N_5832,In_184,In_1413);
or U5833 (N_5833,In_1503,In_2067);
or U5834 (N_5834,In_439,In_1465);
and U5835 (N_5835,In_646,In_545);
nor U5836 (N_5836,In_2003,In_1035);
xnor U5837 (N_5837,In_2240,In_1333);
xor U5838 (N_5838,In_844,In_1160);
and U5839 (N_5839,In_207,In_588);
nor U5840 (N_5840,In_2,In_1508);
and U5841 (N_5841,In_939,In_1046);
nand U5842 (N_5842,In_529,In_1606);
nand U5843 (N_5843,In_1997,In_649);
nor U5844 (N_5844,In_39,In_1013);
or U5845 (N_5845,In_1466,In_2293);
and U5846 (N_5846,In_1746,In_1158);
and U5847 (N_5847,In_1557,In_2245);
or U5848 (N_5848,In_2111,In_305);
xor U5849 (N_5849,In_313,In_1728);
nor U5850 (N_5850,In_127,In_2171);
xor U5851 (N_5851,In_2016,In_682);
xnor U5852 (N_5852,In_429,In_126);
and U5853 (N_5853,In_2162,In_1714);
or U5854 (N_5854,In_558,In_1585);
xor U5855 (N_5855,In_2158,In_251);
nand U5856 (N_5856,In_1373,In_522);
or U5857 (N_5857,In_17,In_1243);
xnor U5858 (N_5858,In_1843,In_289);
and U5859 (N_5859,In_1590,In_302);
nand U5860 (N_5860,In_1853,In_585);
nor U5861 (N_5861,In_993,In_127);
xor U5862 (N_5862,In_1956,In_1166);
xnor U5863 (N_5863,In_1095,In_1294);
nor U5864 (N_5864,In_1106,In_1178);
nand U5865 (N_5865,In_1009,In_401);
nor U5866 (N_5866,In_1880,In_547);
or U5867 (N_5867,In_2398,In_219);
xor U5868 (N_5868,In_1938,In_1220);
nor U5869 (N_5869,In_1146,In_2260);
nor U5870 (N_5870,In_0,In_751);
or U5871 (N_5871,In_1811,In_1525);
xor U5872 (N_5872,In_2278,In_1871);
nor U5873 (N_5873,In_508,In_2282);
nor U5874 (N_5874,In_223,In_360);
and U5875 (N_5875,In_904,In_651);
and U5876 (N_5876,In_328,In_1651);
nor U5877 (N_5877,In_1653,In_499);
and U5878 (N_5878,In_2034,In_2106);
nand U5879 (N_5879,In_77,In_84);
nand U5880 (N_5880,In_1140,In_637);
xor U5881 (N_5881,In_2223,In_2249);
nand U5882 (N_5882,In_2134,In_1576);
and U5883 (N_5883,In_1984,In_1903);
nand U5884 (N_5884,In_563,In_757);
xnor U5885 (N_5885,In_1888,In_2305);
or U5886 (N_5886,In_1942,In_556);
nand U5887 (N_5887,In_178,In_2069);
or U5888 (N_5888,In_1547,In_440);
and U5889 (N_5889,In_1062,In_1105);
nand U5890 (N_5890,In_830,In_1854);
xnor U5891 (N_5891,In_23,In_1886);
or U5892 (N_5892,In_2494,In_1531);
xor U5893 (N_5893,In_1926,In_209);
xnor U5894 (N_5894,In_612,In_682);
nor U5895 (N_5895,In_2062,In_1244);
and U5896 (N_5896,In_955,In_1940);
xor U5897 (N_5897,In_1719,In_1246);
and U5898 (N_5898,In_13,In_842);
nand U5899 (N_5899,In_2450,In_1822);
or U5900 (N_5900,In_1204,In_922);
and U5901 (N_5901,In_204,In_1621);
nand U5902 (N_5902,In_1277,In_1903);
xnor U5903 (N_5903,In_472,In_2208);
xor U5904 (N_5904,In_986,In_2291);
nand U5905 (N_5905,In_1157,In_1121);
nor U5906 (N_5906,In_966,In_499);
and U5907 (N_5907,In_1665,In_2314);
nor U5908 (N_5908,In_1267,In_82);
xnor U5909 (N_5909,In_735,In_2421);
nor U5910 (N_5910,In_2284,In_2069);
nor U5911 (N_5911,In_1414,In_2115);
nor U5912 (N_5912,In_312,In_2170);
nor U5913 (N_5913,In_1090,In_1136);
xnor U5914 (N_5914,In_2433,In_2243);
xnor U5915 (N_5915,In_1125,In_586);
xnor U5916 (N_5916,In_22,In_1832);
and U5917 (N_5917,In_252,In_1981);
or U5918 (N_5918,In_574,In_1049);
nand U5919 (N_5919,In_1738,In_942);
or U5920 (N_5920,In_2367,In_1145);
nor U5921 (N_5921,In_610,In_1610);
nor U5922 (N_5922,In_1713,In_1491);
xor U5923 (N_5923,In_214,In_251);
or U5924 (N_5924,In_2007,In_1994);
and U5925 (N_5925,In_596,In_842);
nor U5926 (N_5926,In_169,In_1002);
nor U5927 (N_5927,In_1138,In_2411);
and U5928 (N_5928,In_2007,In_714);
and U5929 (N_5929,In_1029,In_1557);
nand U5930 (N_5930,In_6,In_2024);
or U5931 (N_5931,In_1152,In_1697);
or U5932 (N_5932,In_2089,In_2079);
nor U5933 (N_5933,In_944,In_1120);
or U5934 (N_5934,In_1566,In_1047);
xnor U5935 (N_5935,In_938,In_1624);
and U5936 (N_5936,In_2435,In_2346);
nor U5937 (N_5937,In_695,In_904);
nor U5938 (N_5938,In_1008,In_650);
nor U5939 (N_5939,In_1403,In_485);
xor U5940 (N_5940,In_1062,In_1091);
and U5941 (N_5941,In_2355,In_1660);
nand U5942 (N_5942,In_348,In_2242);
xnor U5943 (N_5943,In_7,In_365);
and U5944 (N_5944,In_1470,In_190);
xor U5945 (N_5945,In_2099,In_1542);
nand U5946 (N_5946,In_1618,In_2423);
nor U5947 (N_5947,In_192,In_1073);
nand U5948 (N_5948,In_1894,In_1090);
nor U5949 (N_5949,In_256,In_1271);
or U5950 (N_5950,In_691,In_1017);
nor U5951 (N_5951,In_2252,In_261);
nand U5952 (N_5952,In_1793,In_1273);
xor U5953 (N_5953,In_465,In_1452);
xnor U5954 (N_5954,In_2036,In_1984);
nor U5955 (N_5955,In_256,In_795);
or U5956 (N_5956,In_1285,In_172);
nand U5957 (N_5957,In_2389,In_2019);
and U5958 (N_5958,In_1078,In_1938);
nor U5959 (N_5959,In_308,In_2216);
and U5960 (N_5960,In_1285,In_2273);
nand U5961 (N_5961,In_1362,In_1312);
xnor U5962 (N_5962,In_575,In_2214);
and U5963 (N_5963,In_959,In_800);
and U5964 (N_5964,In_224,In_707);
or U5965 (N_5965,In_153,In_1754);
or U5966 (N_5966,In_2305,In_65);
or U5967 (N_5967,In_2133,In_1190);
and U5968 (N_5968,In_515,In_126);
xnor U5969 (N_5969,In_2279,In_1667);
and U5970 (N_5970,In_312,In_2387);
or U5971 (N_5971,In_2157,In_1173);
or U5972 (N_5972,In_2468,In_1076);
xnor U5973 (N_5973,In_1538,In_112);
or U5974 (N_5974,In_509,In_730);
xnor U5975 (N_5975,In_1576,In_367);
and U5976 (N_5976,In_1165,In_1578);
or U5977 (N_5977,In_1129,In_2256);
and U5978 (N_5978,In_1731,In_287);
nand U5979 (N_5979,In_915,In_2306);
nor U5980 (N_5980,In_1653,In_1709);
nor U5981 (N_5981,In_2158,In_2450);
and U5982 (N_5982,In_2348,In_1442);
and U5983 (N_5983,In_2093,In_1720);
or U5984 (N_5984,In_1301,In_2267);
and U5985 (N_5985,In_486,In_1893);
and U5986 (N_5986,In_1049,In_571);
xnor U5987 (N_5987,In_1752,In_2060);
nor U5988 (N_5988,In_1858,In_123);
nor U5989 (N_5989,In_351,In_387);
xor U5990 (N_5990,In_763,In_249);
xnor U5991 (N_5991,In_1412,In_719);
nand U5992 (N_5992,In_2469,In_339);
and U5993 (N_5993,In_198,In_1335);
or U5994 (N_5994,In_1177,In_345);
or U5995 (N_5995,In_1117,In_194);
and U5996 (N_5996,In_1210,In_1023);
or U5997 (N_5997,In_1116,In_1320);
or U5998 (N_5998,In_321,In_665);
xor U5999 (N_5999,In_1705,In_529);
and U6000 (N_6000,In_2058,In_1687);
and U6001 (N_6001,In_1907,In_1551);
xor U6002 (N_6002,In_1100,In_2035);
and U6003 (N_6003,In_1105,In_2005);
xor U6004 (N_6004,In_1267,In_2228);
nor U6005 (N_6005,In_862,In_1916);
nor U6006 (N_6006,In_65,In_1708);
nand U6007 (N_6007,In_2224,In_683);
xor U6008 (N_6008,In_2220,In_1423);
nand U6009 (N_6009,In_417,In_98);
and U6010 (N_6010,In_1332,In_2457);
nor U6011 (N_6011,In_1315,In_2131);
or U6012 (N_6012,In_1160,In_603);
nand U6013 (N_6013,In_1664,In_1567);
nand U6014 (N_6014,In_713,In_1180);
xnor U6015 (N_6015,In_33,In_1847);
nor U6016 (N_6016,In_403,In_556);
nor U6017 (N_6017,In_1290,In_312);
xor U6018 (N_6018,In_1758,In_1315);
or U6019 (N_6019,In_762,In_2024);
nor U6020 (N_6020,In_1702,In_488);
and U6021 (N_6021,In_922,In_617);
and U6022 (N_6022,In_1192,In_948);
and U6023 (N_6023,In_459,In_299);
nor U6024 (N_6024,In_825,In_1087);
nor U6025 (N_6025,In_45,In_2255);
xor U6026 (N_6026,In_804,In_1772);
or U6027 (N_6027,In_979,In_422);
nor U6028 (N_6028,In_2462,In_2218);
or U6029 (N_6029,In_1043,In_2365);
or U6030 (N_6030,In_55,In_1158);
nor U6031 (N_6031,In_1437,In_1026);
or U6032 (N_6032,In_831,In_29);
or U6033 (N_6033,In_2190,In_44);
and U6034 (N_6034,In_1705,In_1914);
or U6035 (N_6035,In_216,In_567);
and U6036 (N_6036,In_541,In_1033);
xnor U6037 (N_6037,In_2083,In_2342);
nand U6038 (N_6038,In_2341,In_1330);
xnor U6039 (N_6039,In_2134,In_1802);
nor U6040 (N_6040,In_1504,In_2415);
nor U6041 (N_6041,In_1106,In_2119);
nand U6042 (N_6042,In_135,In_789);
xor U6043 (N_6043,In_847,In_1417);
nand U6044 (N_6044,In_599,In_522);
nand U6045 (N_6045,In_1658,In_841);
nor U6046 (N_6046,In_1941,In_550);
nor U6047 (N_6047,In_1619,In_968);
xor U6048 (N_6048,In_1023,In_607);
and U6049 (N_6049,In_1002,In_1154);
nand U6050 (N_6050,In_1403,In_1303);
nand U6051 (N_6051,In_1944,In_1931);
xor U6052 (N_6052,In_1623,In_604);
nor U6053 (N_6053,In_1515,In_73);
nor U6054 (N_6054,In_619,In_562);
xor U6055 (N_6055,In_1340,In_2293);
and U6056 (N_6056,In_387,In_2303);
and U6057 (N_6057,In_157,In_1005);
xnor U6058 (N_6058,In_1263,In_534);
nor U6059 (N_6059,In_27,In_1739);
nor U6060 (N_6060,In_496,In_1088);
or U6061 (N_6061,In_1614,In_2077);
xor U6062 (N_6062,In_1521,In_1700);
xnor U6063 (N_6063,In_1646,In_1642);
and U6064 (N_6064,In_1997,In_1785);
or U6065 (N_6065,In_1341,In_1516);
xnor U6066 (N_6066,In_1622,In_2233);
nor U6067 (N_6067,In_628,In_418);
or U6068 (N_6068,In_1962,In_1292);
or U6069 (N_6069,In_738,In_1316);
nand U6070 (N_6070,In_672,In_576);
nor U6071 (N_6071,In_1331,In_871);
nand U6072 (N_6072,In_2060,In_105);
nand U6073 (N_6073,In_1349,In_92);
and U6074 (N_6074,In_1484,In_127);
nand U6075 (N_6075,In_1867,In_1860);
xor U6076 (N_6076,In_1109,In_568);
or U6077 (N_6077,In_1848,In_2406);
or U6078 (N_6078,In_70,In_2023);
nand U6079 (N_6079,In_460,In_2435);
or U6080 (N_6080,In_1881,In_1201);
nor U6081 (N_6081,In_828,In_2432);
nand U6082 (N_6082,In_1944,In_1339);
nand U6083 (N_6083,In_215,In_1488);
or U6084 (N_6084,In_1336,In_1108);
nor U6085 (N_6085,In_342,In_2457);
nand U6086 (N_6086,In_1504,In_1323);
nand U6087 (N_6087,In_872,In_1303);
nand U6088 (N_6088,In_1229,In_1571);
or U6089 (N_6089,In_2429,In_1020);
and U6090 (N_6090,In_58,In_2027);
or U6091 (N_6091,In_1699,In_2419);
xor U6092 (N_6092,In_1147,In_2040);
or U6093 (N_6093,In_1449,In_1304);
nand U6094 (N_6094,In_1904,In_2387);
and U6095 (N_6095,In_406,In_1468);
and U6096 (N_6096,In_1962,In_2179);
and U6097 (N_6097,In_2338,In_1781);
xor U6098 (N_6098,In_1579,In_979);
xnor U6099 (N_6099,In_762,In_1193);
nor U6100 (N_6100,In_2485,In_1902);
or U6101 (N_6101,In_1189,In_1237);
xor U6102 (N_6102,In_1825,In_348);
nor U6103 (N_6103,In_498,In_274);
and U6104 (N_6104,In_2452,In_399);
nand U6105 (N_6105,In_1494,In_288);
nand U6106 (N_6106,In_885,In_3);
nor U6107 (N_6107,In_104,In_2345);
nand U6108 (N_6108,In_2118,In_304);
nor U6109 (N_6109,In_54,In_1942);
and U6110 (N_6110,In_2398,In_1765);
nand U6111 (N_6111,In_417,In_1457);
nand U6112 (N_6112,In_1203,In_763);
nand U6113 (N_6113,In_2325,In_638);
or U6114 (N_6114,In_371,In_119);
xor U6115 (N_6115,In_2310,In_634);
and U6116 (N_6116,In_57,In_77);
or U6117 (N_6117,In_326,In_912);
nand U6118 (N_6118,In_1555,In_1106);
nor U6119 (N_6119,In_44,In_1025);
xor U6120 (N_6120,In_436,In_697);
and U6121 (N_6121,In_2429,In_1272);
nor U6122 (N_6122,In_1391,In_944);
and U6123 (N_6123,In_1042,In_496);
nor U6124 (N_6124,In_898,In_1699);
or U6125 (N_6125,In_713,In_2043);
xnor U6126 (N_6126,In_1642,In_565);
and U6127 (N_6127,In_392,In_49);
nand U6128 (N_6128,In_1141,In_841);
and U6129 (N_6129,In_1671,In_1026);
or U6130 (N_6130,In_2313,In_1367);
nand U6131 (N_6131,In_146,In_734);
or U6132 (N_6132,In_383,In_682);
nand U6133 (N_6133,In_2391,In_1133);
or U6134 (N_6134,In_986,In_1980);
xnor U6135 (N_6135,In_238,In_1609);
or U6136 (N_6136,In_1793,In_1691);
and U6137 (N_6137,In_1657,In_1835);
nand U6138 (N_6138,In_1910,In_1376);
xor U6139 (N_6139,In_1965,In_408);
or U6140 (N_6140,In_1073,In_78);
nand U6141 (N_6141,In_1757,In_1135);
and U6142 (N_6142,In_932,In_1987);
or U6143 (N_6143,In_2201,In_1702);
xor U6144 (N_6144,In_1020,In_2028);
xor U6145 (N_6145,In_785,In_2339);
nor U6146 (N_6146,In_1376,In_442);
and U6147 (N_6147,In_459,In_1677);
xnor U6148 (N_6148,In_726,In_2225);
or U6149 (N_6149,In_1813,In_937);
or U6150 (N_6150,In_33,In_1686);
nor U6151 (N_6151,In_534,In_2323);
xnor U6152 (N_6152,In_1548,In_1815);
xor U6153 (N_6153,In_2217,In_430);
nand U6154 (N_6154,In_680,In_1377);
nand U6155 (N_6155,In_521,In_2139);
nor U6156 (N_6156,In_2073,In_380);
and U6157 (N_6157,In_1055,In_2065);
xnor U6158 (N_6158,In_1650,In_847);
nand U6159 (N_6159,In_654,In_2079);
or U6160 (N_6160,In_1743,In_546);
or U6161 (N_6161,In_866,In_699);
or U6162 (N_6162,In_417,In_2322);
or U6163 (N_6163,In_523,In_1610);
or U6164 (N_6164,In_2438,In_258);
or U6165 (N_6165,In_343,In_1732);
xor U6166 (N_6166,In_1584,In_637);
nand U6167 (N_6167,In_1999,In_1910);
and U6168 (N_6168,In_922,In_249);
and U6169 (N_6169,In_394,In_1494);
xor U6170 (N_6170,In_1284,In_962);
nand U6171 (N_6171,In_1180,In_1480);
nor U6172 (N_6172,In_2073,In_1997);
or U6173 (N_6173,In_271,In_2499);
or U6174 (N_6174,In_2370,In_1290);
xnor U6175 (N_6175,In_2284,In_435);
nor U6176 (N_6176,In_754,In_973);
and U6177 (N_6177,In_2375,In_788);
nor U6178 (N_6178,In_610,In_581);
or U6179 (N_6179,In_1612,In_671);
and U6180 (N_6180,In_728,In_1388);
and U6181 (N_6181,In_2059,In_1459);
nand U6182 (N_6182,In_1211,In_1351);
and U6183 (N_6183,In_177,In_2409);
nand U6184 (N_6184,In_445,In_1394);
and U6185 (N_6185,In_1511,In_2338);
nor U6186 (N_6186,In_1512,In_2328);
nand U6187 (N_6187,In_2294,In_1931);
nand U6188 (N_6188,In_2328,In_1365);
or U6189 (N_6189,In_66,In_615);
nor U6190 (N_6190,In_168,In_1672);
xnor U6191 (N_6191,In_60,In_2025);
xnor U6192 (N_6192,In_2169,In_2360);
xnor U6193 (N_6193,In_58,In_59);
and U6194 (N_6194,In_1829,In_828);
nand U6195 (N_6195,In_927,In_503);
xor U6196 (N_6196,In_1536,In_2180);
nor U6197 (N_6197,In_384,In_2217);
nor U6198 (N_6198,In_2378,In_2439);
and U6199 (N_6199,In_2320,In_1033);
and U6200 (N_6200,In_1096,In_1825);
nor U6201 (N_6201,In_2330,In_1888);
nand U6202 (N_6202,In_2090,In_445);
and U6203 (N_6203,In_649,In_501);
nand U6204 (N_6204,In_1830,In_1532);
or U6205 (N_6205,In_2135,In_452);
xor U6206 (N_6206,In_2244,In_2482);
and U6207 (N_6207,In_307,In_1905);
nor U6208 (N_6208,In_523,In_51);
nor U6209 (N_6209,In_2076,In_1181);
or U6210 (N_6210,In_867,In_1180);
nand U6211 (N_6211,In_1542,In_2052);
nand U6212 (N_6212,In_1977,In_995);
nor U6213 (N_6213,In_2186,In_1561);
xor U6214 (N_6214,In_298,In_516);
or U6215 (N_6215,In_1705,In_731);
xor U6216 (N_6216,In_1097,In_692);
xor U6217 (N_6217,In_1770,In_2495);
and U6218 (N_6218,In_1807,In_1358);
xnor U6219 (N_6219,In_2086,In_37);
nor U6220 (N_6220,In_1255,In_1428);
or U6221 (N_6221,In_1328,In_750);
or U6222 (N_6222,In_642,In_347);
and U6223 (N_6223,In_2114,In_372);
nor U6224 (N_6224,In_369,In_966);
nor U6225 (N_6225,In_2027,In_1776);
xor U6226 (N_6226,In_855,In_2032);
nor U6227 (N_6227,In_1374,In_1245);
or U6228 (N_6228,In_519,In_1869);
and U6229 (N_6229,In_826,In_2187);
xor U6230 (N_6230,In_2190,In_1955);
xnor U6231 (N_6231,In_765,In_1314);
xor U6232 (N_6232,In_1665,In_1084);
nand U6233 (N_6233,In_2350,In_2177);
nand U6234 (N_6234,In_1853,In_1851);
nand U6235 (N_6235,In_1406,In_1041);
or U6236 (N_6236,In_1647,In_1959);
nand U6237 (N_6237,In_1430,In_2010);
xnor U6238 (N_6238,In_2405,In_994);
and U6239 (N_6239,In_690,In_1933);
nor U6240 (N_6240,In_1118,In_603);
nor U6241 (N_6241,In_1525,In_345);
and U6242 (N_6242,In_545,In_1911);
and U6243 (N_6243,In_1661,In_40);
nor U6244 (N_6244,In_1979,In_216);
nand U6245 (N_6245,In_449,In_1979);
nor U6246 (N_6246,In_1277,In_1368);
and U6247 (N_6247,In_1988,In_893);
and U6248 (N_6248,In_1142,In_1435);
and U6249 (N_6249,In_2173,In_92);
nor U6250 (N_6250,N_3629,N_6097);
nor U6251 (N_6251,N_4975,N_2995);
nor U6252 (N_6252,N_4786,N_3539);
xnor U6253 (N_6253,N_1158,N_768);
and U6254 (N_6254,N_771,N_2593);
or U6255 (N_6255,N_1912,N_2457);
nor U6256 (N_6256,N_3584,N_2844);
nor U6257 (N_6257,N_2701,N_2374);
or U6258 (N_6258,N_5248,N_3905);
nor U6259 (N_6259,N_703,N_4691);
nor U6260 (N_6260,N_5773,N_4366);
nor U6261 (N_6261,N_5740,N_5944);
nand U6262 (N_6262,N_4046,N_3470);
nand U6263 (N_6263,N_4248,N_2114);
nand U6264 (N_6264,N_5220,N_3908);
xnor U6265 (N_6265,N_2389,N_827);
xnor U6266 (N_6266,N_377,N_2443);
or U6267 (N_6267,N_416,N_419);
xor U6268 (N_6268,N_2221,N_4392);
or U6269 (N_6269,N_1669,N_2375);
and U6270 (N_6270,N_2670,N_2472);
and U6271 (N_6271,N_3604,N_1133);
and U6272 (N_6272,N_2352,N_4995);
xor U6273 (N_6273,N_3952,N_5455);
or U6274 (N_6274,N_3519,N_5934);
nand U6275 (N_6275,N_3988,N_1592);
nor U6276 (N_6276,N_645,N_5490);
or U6277 (N_6277,N_229,N_6152);
or U6278 (N_6278,N_4315,N_2083);
and U6279 (N_6279,N_4679,N_5257);
nand U6280 (N_6280,N_2402,N_1676);
nand U6281 (N_6281,N_2179,N_2590);
nand U6282 (N_6282,N_4860,N_2610);
or U6283 (N_6283,N_2945,N_6041);
and U6284 (N_6284,N_3244,N_4377);
nand U6285 (N_6285,N_3522,N_2511);
and U6286 (N_6286,N_1111,N_5504);
or U6287 (N_6287,N_2267,N_614);
or U6288 (N_6288,N_4038,N_1447);
xor U6289 (N_6289,N_3137,N_670);
and U6290 (N_6290,N_5725,N_5562);
and U6291 (N_6291,N_424,N_5909);
or U6292 (N_6292,N_4822,N_5601);
or U6293 (N_6293,N_3845,N_1638);
xnor U6294 (N_6294,N_249,N_2488);
or U6295 (N_6295,N_444,N_2287);
nor U6296 (N_6296,N_418,N_1875);
nor U6297 (N_6297,N_3619,N_6134);
and U6298 (N_6298,N_2621,N_2341);
xor U6299 (N_6299,N_1119,N_5958);
nand U6300 (N_6300,N_585,N_4701);
nand U6301 (N_6301,N_244,N_4967);
xnor U6302 (N_6302,N_886,N_4211);
nand U6303 (N_6303,N_2058,N_1361);
nor U6304 (N_6304,N_185,N_3714);
nor U6305 (N_6305,N_4693,N_2640);
nand U6306 (N_6306,N_815,N_359);
nand U6307 (N_6307,N_564,N_3465);
nand U6308 (N_6308,N_5786,N_540);
and U6309 (N_6309,N_3931,N_1194);
nand U6310 (N_6310,N_944,N_4240);
nor U6311 (N_6311,N_4141,N_765);
xnor U6312 (N_6312,N_5249,N_4403);
xor U6313 (N_6313,N_2420,N_4996);
nand U6314 (N_6314,N_5791,N_3422);
nor U6315 (N_6315,N_5412,N_3155);
and U6316 (N_6316,N_3111,N_3225);
nand U6317 (N_6317,N_4711,N_2202);
nor U6318 (N_6318,N_3737,N_2134);
xor U6319 (N_6319,N_3428,N_84);
and U6320 (N_6320,N_5263,N_998);
nor U6321 (N_6321,N_3708,N_5867);
or U6322 (N_6322,N_2490,N_1419);
xnor U6323 (N_6323,N_6157,N_4533);
and U6324 (N_6324,N_2576,N_3805);
nor U6325 (N_6325,N_1320,N_480);
and U6326 (N_6326,N_989,N_3408);
nor U6327 (N_6327,N_5034,N_1177);
xnor U6328 (N_6328,N_5957,N_3592);
xnor U6329 (N_6329,N_145,N_4184);
or U6330 (N_6330,N_3031,N_3828);
and U6331 (N_6331,N_1706,N_6091);
and U6332 (N_6332,N_1748,N_3966);
xnor U6333 (N_6333,N_3199,N_5981);
nand U6334 (N_6334,N_710,N_3792);
xnor U6335 (N_6335,N_6086,N_2695);
xor U6336 (N_6336,N_1917,N_3882);
and U6337 (N_6337,N_3634,N_2192);
nand U6338 (N_6338,N_1034,N_3261);
xor U6339 (N_6339,N_4775,N_1244);
or U6340 (N_6340,N_3733,N_3844);
nand U6341 (N_6341,N_5564,N_652);
or U6342 (N_6342,N_2525,N_5092);
nor U6343 (N_6343,N_2999,N_1427);
nand U6344 (N_6344,N_182,N_4953);
nor U6345 (N_6345,N_2749,N_2926);
and U6346 (N_6346,N_2757,N_3383);
nor U6347 (N_6347,N_1303,N_4472);
and U6348 (N_6348,N_3223,N_5202);
xnor U6349 (N_6349,N_758,N_5319);
and U6350 (N_6350,N_516,N_48);
and U6351 (N_6351,N_5609,N_5528);
or U6352 (N_6352,N_3872,N_5965);
and U6353 (N_6353,N_5332,N_3332);
nor U6354 (N_6354,N_931,N_4842);
nand U6355 (N_6355,N_5394,N_5181);
and U6356 (N_6356,N_2030,N_4872);
or U6357 (N_6357,N_3684,N_657);
nand U6358 (N_6358,N_1659,N_512);
xor U6359 (N_6359,N_4130,N_2264);
nor U6360 (N_6360,N_5897,N_3846);
nand U6361 (N_6361,N_4567,N_4494);
xor U6362 (N_6362,N_1124,N_150);
xnor U6363 (N_6363,N_1752,N_1157);
xnor U6364 (N_6364,N_4960,N_1895);
nand U6365 (N_6365,N_3642,N_1190);
nor U6366 (N_6366,N_1742,N_35);
nand U6367 (N_6367,N_2155,N_1134);
xor U6368 (N_6368,N_5076,N_4944);
nand U6369 (N_6369,N_4600,N_6104);
and U6370 (N_6370,N_4294,N_3163);
and U6371 (N_6371,N_4964,N_4192);
xor U6372 (N_6372,N_180,N_690);
or U6373 (N_6373,N_3214,N_173);
or U6374 (N_6374,N_4805,N_3541);
nor U6375 (N_6375,N_2406,N_5375);
xor U6376 (N_6376,N_3655,N_5453);
nand U6377 (N_6377,N_1822,N_2300);
or U6378 (N_6378,N_2778,N_4004);
or U6379 (N_6379,N_5531,N_5086);
and U6380 (N_6380,N_1193,N_3531);
or U6381 (N_6381,N_1670,N_1282);
xnor U6382 (N_6382,N_2400,N_3020);
and U6383 (N_6383,N_3812,N_3994);
nand U6384 (N_6384,N_3645,N_591);
xnor U6385 (N_6385,N_4589,N_1746);
nand U6386 (N_6386,N_628,N_5150);
or U6387 (N_6387,N_4512,N_295);
xor U6388 (N_6388,N_5733,N_874);
xnor U6389 (N_6389,N_4927,N_5316);
nand U6390 (N_6390,N_2917,N_2512);
nand U6391 (N_6391,N_5955,N_2830);
xnor U6392 (N_6392,N_6095,N_3780);
nand U6393 (N_6393,N_3478,N_4994);
nor U6394 (N_6394,N_3766,N_3011);
and U6395 (N_6395,N_2685,N_2183);
xnor U6396 (N_6396,N_4848,N_2542);
nand U6397 (N_6397,N_2851,N_1508);
or U6398 (N_6398,N_1088,N_2760);
or U6399 (N_6399,N_544,N_2766);
xor U6400 (N_6400,N_5060,N_2638);
or U6401 (N_6401,N_3398,N_4478);
or U6402 (N_6402,N_4982,N_2803);
xor U6403 (N_6403,N_2022,N_4083);
or U6404 (N_6404,N_3987,N_918);
and U6405 (N_6405,N_2820,N_6121);
and U6406 (N_6406,N_1653,N_3929);
and U6407 (N_6407,N_2632,N_5831);
nand U6408 (N_6408,N_1780,N_5515);
nand U6409 (N_6409,N_4210,N_2273);
or U6410 (N_6410,N_3120,N_5828);
and U6411 (N_6411,N_5846,N_2816);
or U6412 (N_6412,N_4262,N_2673);
nor U6413 (N_6413,N_1403,N_5424);
and U6414 (N_6414,N_1219,N_5629);
or U6415 (N_6415,N_5172,N_5517);
nand U6416 (N_6416,N_1665,N_4666);
xnor U6417 (N_6417,N_3041,N_5621);
or U6418 (N_6418,N_3884,N_5117);
xnor U6419 (N_6419,N_707,N_1646);
or U6420 (N_6420,N_2852,N_5167);
xor U6421 (N_6421,N_1835,N_624);
nor U6422 (N_6422,N_4115,N_2465);
nand U6423 (N_6423,N_3087,N_2990);
nand U6424 (N_6424,N_1873,N_3823);
or U6425 (N_6425,N_3509,N_2002);
nor U6426 (N_6426,N_967,N_2763);
or U6427 (N_6427,N_3854,N_5668);
nor U6428 (N_6428,N_5112,N_5323);
and U6429 (N_6429,N_4131,N_3969);
xnor U6430 (N_6430,N_233,N_5469);
xnor U6431 (N_6431,N_2100,N_4959);
nand U6432 (N_6432,N_4214,N_5447);
xor U6433 (N_6433,N_341,N_1591);
or U6434 (N_6434,N_1285,N_1781);
nor U6435 (N_6435,N_3382,N_5577);
and U6436 (N_6436,N_5251,N_3360);
and U6437 (N_6437,N_5523,N_1518);
nand U6438 (N_6438,N_2009,N_620);
xnor U6439 (N_6439,N_307,N_4002);
xor U6440 (N_6440,N_423,N_1817);
xnor U6441 (N_6441,N_2158,N_5492);
nand U6442 (N_6442,N_6160,N_5479);
and U6443 (N_6443,N_3207,N_1496);
nor U6444 (N_6444,N_4317,N_4109);
and U6445 (N_6445,N_629,N_3633);
or U6446 (N_6446,N_700,N_1547);
nor U6447 (N_6447,N_4560,N_2679);
or U6448 (N_6448,N_3935,N_3082);
xnor U6449 (N_6449,N_5992,N_4074);
xnor U6450 (N_6450,N_4970,N_1245);
xnor U6451 (N_6451,N_2654,N_6026);
or U6452 (N_6452,N_841,N_2359);
and U6453 (N_6453,N_4321,N_77);
or U6454 (N_6454,N_1163,N_3683);
nand U6455 (N_6455,N_531,N_6228);
xnor U6456 (N_6456,N_636,N_2107);
xnor U6457 (N_6457,N_5315,N_1605);
xnor U6458 (N_6458,N_747,N_5380);
nor U6459 (N_6459,N_2552,N_4837);
and U6460 (N_6460,N_470,N_3387);
or U6461 (N_6461,N_5575,N_1604);
and U6462 (N_6462,N_1795,N_2655);
or U6463 (N_6463,N_6237,N_6223);
nor U6464 (N_6464,N_3896,N_3572);
and U6465 (N_6465,N_308,N_828);
nor U6466 (N_6466,N_253,N_2631);
nand U6467 (N_6467,N_4823,N_2815);
nand U6468 (N_6468,N_3279,N_5038);
xnor U6469 (N_6469,N_607,N_5074);
nor U6470 (N_6470,N_5713,N_4370);
nor U6471 (N_6471,N_2825,N_872);
and U6472 (N_6472,N_1899,N_1929);
xnor U6473 (N_6473,N_1626,N_1637);
or U6474 (N_6474,N_1035,N_817);
xor U6475 (N_6475,N_2506,N_5650);
nand U6476 (N_6476,N_2156,N_2170);
nor U6477 (N_6477,N_6094,N_1750);
or U6478 (N_6478,N_4182,N_5374);
and U6479 (N_6479,N_5694,N_4509);
nand U6480 (N_6480,N_1350,N_306);
or U6481 (N_6481,N_4120,N_1504);
nor U6482 (N_6482,N_5090,N_1732);
xnor U6483 (N_6483,N_1559,N_1054);
or U6484 (N_6484,N_4898,N_274);
xor U6485 (N_6485,N_5945,N_2249);
xnor U6486 (N_6486,N_4025,N_5045);
and U6487 (N_6487,N_4851,N_4892);
or U6488 (N_6488,N_2897,N_1624);
or U6489 (N_6489,N_1884,N_2424);
xnor U6490 (N_6490,N_3260,N_4780);
xor U6491 (N_6491,N_315,N_67);
and U6492 (N_6492,N_4980,N_5085);
xnor U6493 (N_6493,N_3299,N_3363);
and U6494 (N_6494,N_38,N_2948);
or U6495 (N_6495,N_1718,N_3088);
xnor U6496 (N_6496,N_1384,N_17);
nand U6497 (N_6497,N_2203,N_1411);
or U6498 (N_6498,N_366,N_3991);
nor U6499 (N_6499,N_973,N_3038);
nand U6500 (N_6500,N_3226,N_5704);
xor U6501 (N_6501,N_99,N_1811);
nand U6502 (N_6502,N_5298,N_954);
nand U6503 (N_6503,N_1114,N_1315);
nor U6504 (N_6504,N_280,N_5735);
xor U6505 (N_6505,N_4066,N_1333);
nand U6506 (N_6506,N_999,N_1269);
nand U6507 (N_6507,N_488,N_4069);
xor U6508 (N_6508,N_4625,N_2000);
xor U6509 (N_6509,N_126,N_1443);
and U6510 (N_6510,N_3526,N_5377);
nor U6511 (N_6511,N_165,N_5480);
xnor U6512 (N_6512,N_2079,N_3463);
and U6513 (N_6513,N_3400,N_5819);
nand U6514 (N_6514,N_4636,N_5578);
or U6515 (N_6515,N_3173,N_662);
nor U6516 (N_6516,N_5497,N_1429);
and U6517 (N_6517,N_1844,N_81);
or U6518 (N_6518,N_1627,N_291);
or U6519 (N_6519,N_3649,N_5751);
and U6520 (N_6520,N_5947,N_1451);
and U6521 (N_6521,N_1914,N_4945);
nand U6522 (N_6522,N_2435,N_316);
nor U6523 (N_6523,N_2061,N_3471);
and U6524 (N_6524,N_934,N_4225);
and U6525 (N_6525,N_5916,N_1023);
or U6526 (N_6526,N_2832,N_1513);
nand U6527 (N_6527,N_692,N_3103);
and U6528 (N_6528,N_4414,N_3089);
nand U6529 (N_6529,N_2343,N_4782);
or U6530 (N_6530,N_5581,N_2565);
or U6531 (N_6531,N_3608,N_2937);
nor U6532 (N_6532,N_2947,N_264);
and U6533 (N_6533,N_689,N_2703);
xnor U6534 (N_6534,N_176,N_5130);
nor U6535 (N_6535,N_500,N_4270);
and U6536 (N_6536,N_3615,N_674);
or U6537 (N_6537,N_2024,N_169);
nand U6538 (N_6538,N_243,N_2605);
nand U6539 (N_6539,N_4882,N_0);
xor U6540 (N_6540,N_2821,N_4511);
nand U6541 (N_6541,N_2784,N_503);
xnor U6542 (N_6542,N_902,N_4457);
and U6543 (N_6543,N_957,N_1127);
or U6544 (N_6544,N_5120,N_221);
nor U6545 (N_6545,N_935,N_2041);
nor U6546 (N_6546,N_457,N_5418);
or U6547 (N_6547,N_4889,N_3004);
or U6548 (N_6548,N_1,N_5776);
xor U6549 (N_6549,N_2016,N_580);
nand U6550 (N_6550,N_310,N_873);
or U6551 (N_6551,N_5718,N_2120);
or U6552 (N_6552,N_3467,N_4737);
nand U6553 (N_6553,N_3488,N_1717);
and U6554 (N_6554,N_1967,N_2275);
nand U6555 (N_6555,N_3962,N_5977);
and U6556 (N_6556,N_1985,N_1568);
nor U6557 (N_6557,N_2053,N_4274);
nand U6558 (N_6558,N_5851,N_3959);
or U6559 (N_6559,N_2042,N_3493);
xnor U6560 (N_6560,N_5449,N_2925);
or U6561 (N_6561,N_4904,N_1255);
xnor U6562 (N_6562,N_1038,N_3809);
nand U6563 (N_6563,N_5296,N_3536);
xnor U6564 (N_6564,N_5863,N_5306);
nor U6565 (N_6565,N_1691,N_5078);
or U6566 (N_6566,N_2367,N_5547);
xor U6567 (N_6567,N_2276,N_4900);
nand U6568 (N_6568,N_5289,N_5844);
xor U6569 (N_6569,N_3913,N_583);
nor U6570 (N_6570,N_3549,N_3009);
nand U6571 (N_6571,N_753,N_2860);
nor U6572 (N_6572,N_1342,N_120);
and U6573 (N_6573,N_393,N_3235);
nand U6574 (N_6574,N_677,N_6061);
nand U6575 (N_6575,N_5646,N_24);
nand U6576 (N_6576,N_2785,N_4932);
or U6577 (N_6577,N_701,N_5813);
nand U6578 (N_6578,N_349,N_2034);
nor U6579 (N_6579,N_3601,N_3118);
and U6580 (N_6580,N_5665,N_560);
and U6581 (N_6581,N_2805,N_1402);
and U6582 (N_6582,N_6052,N_494);
xnor U6583 (N_6583,N_992,N_6105);
nand U6584 (N_6584,N_1457,N_25);
nand U6585 (N_6585,N_4316,N_491);
xnor U6586 (N_6586,N_2991,N_5989);
nor U6587 (N_6587,N_4217,N_2697);
and U6588 (N_6588,N_1128,N_3753);
or U6589 (N_6589,N_5333,N_2672);
nand U6590 (N_6590,N_4971,N_4745);
or U6591 (N_6591,N_3600,N_2021);
nor U6592 (N_6592,N_776,N_402);
xnor U6593 (N_6593,N_1071,N_3015);
nand U6594 (N_6594,N_5829,N_4330);
or U6595 (N_6595,N_4553,N_2123);
or U6596 (N_6596,N_960,N_4524);
nor U6597 (N_6597,N_4830,N_2004);
and U6598 (N_6598,N_5104,N_4716);
nand U6599 (N_6599,N_2329,N_2770);
nand U6600 (N_6600,N_927,N_4452);
and U6601 (N_6601,N_806,N_3256);
and U6602 (N_6602,N_6078,N_2719);
and U6603 (N_6603,N_2879,N_6166);
xor U6604 (N_6604,N_5197,N_1357);
nor U6605 (N_6605,N_4643,N_345);
nand U6606 (N_6606,N_413,N_2536);
xnor U6607 (N_6607,N_4529,N_5689);
xnor U6608 (N_6608,N_526,N_1955);
or U6609 (N_6609,N_822,N_2228);
or U6610 (N_6610,N_5710,N_3414);
or U6611 (N_6611,N_2121,N_2417);
nand U6612 (N_6612,N_4163,N_2464);
or U6613 (N_6613,N_1837,N_472);
nor U6614 (N_6614,N_4514,N_2366);
or U6615 (N_6615,N_1058,N_581);
and U6616 (N_6616,N_338,N_2445);
nand U6617 (N_6617,N_3175,N_3501);
nor U6618 (N_6618,N_1956,N_460);
xnor U6619 (N_6619,N_610,N_4307);
and U6620 (N_6620,N_157,N_5613);
nand U6621 (N_6621,N_4078,N_5189);
xnor U6622 (N_6622,N_2976,N_5586);
or U6623 (N_6623,N_625,N_3293);
nand U6624 (N_6624,N_4912,N_1861);
or U6625 (N_6625,N_602,N_1405);
and U6626 (N_6626,N_368,N_4474);
xor U6627 (N_6627,N_3930,N_3210);
or U6628 (N_6628,N_4629,N_752);
or U6629 (N_6629,N_1398,N_6096);
nor U6630 (N_6630,N_3919,N_3984);
xor U6631 (N_6631,N_4869,N_816);
and U6632 (N_6632,N_4049,N_4379);
xor U6633 (N_6633,N_1919,N_1898);
nor U6634 (N_6634,N_1032,N_592);
nand U6635 (N_6635,N_777,N_2476);
nor U6636 (N_6636,N_5529,N_497);
nor U6637 (N_6637,N_5914,N_6010);
or U6638 (N_6638,N_1329,N_3694);
or U6639 (N_6639,N_2164,N_2579);
and U6640 (N_6640,N_722,N_3081);
and U6641 (N_6641,N_972,N_2358);
xor U6642 (N_6642,N_807,N_4776);
nor U6643 (N_6643,N_74,N_3142);
xor U6644 (N_6644,N_5643,N_496);
xnor U6645 (N_6645,N_6247,N_2858);
xor U6646 (N_6646,N_5759,N_2639);
nor U6647 (N_6647,N_3850,N_5638);
and U6648 (N_6648,N_5278,N_5177);
or U6649 (N_6649,N_4208,N_5388);
nand U6650 (N_6650,N_5381,N_2233);
and U6651 (N_6651,N_4827,N_5505);
and U6652 (N_6652,N_2798,N_1102);
and U6653 (N_6653,N_5135,N_5576);
nand U6654 (N_6654,N_2483,N_5911);
or U6655 (N_6655,N_3911,N_6133);
xor U6656 (N_6656,N_2152,N_54);
nor U6657 (N_6657,N_3014,N_5420);
xor U6658 (N_6658,N_5811,N_2014);
nand U6659 (N_6659,N_3889,N_299);
nor U6660 (N_6660,N_1227,N_4221);
nand U6661 (N_6661,N_3401,N_2978);
or U6662 (N_6662,N_3076,N_5703);
and U6663 (N_6663,N_4997,N_3329);
xor U6664 (N_6664,N_917,N_1876);
xnor U6665 (N_6665,N_46,N_204);
and U6666 (N_6666,N_1546,N_4481);
or U6667 (N_6667,N_2438,N_5138);
nand U6668 (N_6668,N_880,N_518);
or U6669 (N_6669,N_321,N_114);
or U6670 (N_6670,N_4581,N_5818);
or U6671 (N_6671,N_759,N_991);
xnor U6672 (N_6672,N_864,N_2508);
nor U6673 (N_6673,N_857,N_3603);
nor U6674 (N_6674,N_4770,N_705);
nand U6675 (N_6675,N_4467,N_1011);
or U6676 (N_6676,N_4697,N_3143);
and U6677 (N_6677,N_4398,N_4267);
and U6678 (N_6678,N_1075,N_4537);
xor U6679 (N_6679,N_5917,N_4611);
nand U6680 (N_6680,N_1891,N_2437);
xor U6681 (N_6681,N_3295,N_5254);
xor U6682 (N_6682,N_2268,N_5148);
or U6683 (N_6683,N_3628,N_2663);
nand U6684 (N_6684,N_4369,N_5218);
nand U6685 (N_6685,N_1712,N_5842);
nand U6686 (N_6686,N_3134,N_2133);
nor U6687 (N_6687,N_2169,N_3373);
and U6688 (N_6688,N_2109,N_6051);
or U6689 (N_6689,N_1213,N_4495);
nand U6690 (N_6690,N_2773,N_4979);
or U6691 (N_6691,N_2001,N_869);
xor U6692 (N_6692,N_1186,N_2197);
xnor U6693 (N_6693,N_866,N_2873);
xor U6694 (N_6694,N_4844,N_735);
nand U6695 (N_6695,N_1341,N_6098);
or U6696 (N_6696,N_4488,N_2376);
nand U6697 (N_6697,N_5737,N_527);
nand U6698 (N_6698,N_6170,N_5877);
nand U6699 (N_6699,N_4672,N_5003);
nand U6700 (N_6700,N_2979,N_4929);
nor U6701 (N_6701,N_669,N_1662);
nand U6702 (N_6702,N_3249,N_1330);
xor U6703 (N_6703,N_4277,N_837);
and U6704 (N_6704,N_4862,N_4309);
xnor U6705 (N_6705,N_2215,N_3877);
and U6706 (N_6706,N_3754,N_1561);
nor U6707 (N_6707,N_5262,N_5727);
and U6708 (N_6708,N_4358,N_4520);
and U6709 (N_6709,N_5188,N_951);
nand U6710 (N_6710,N_2449,N_4938);
or U6711 (N_6711,N_2835,N_2587);
or U6712 (N_6712,N_6154,N_133);
xnor U6713 (N_6713,N_2236,N_164);
xor U6714 (N_6714,N_4203,N_5013);
nor U6715 (N_6715,N_351,N_1367);
nor U6716 (N_6716,N_49,N_2814);
xnor U6717 (N_6717,N_1521,N_1253);
xnor U6718 (N_6718,N_1866,N_139);
nand U6719 (N_6719,N_5072,N_2140);
or U6720 (N_6720,N_2921,N_1577);
or U6721 (N_6721,N_4329,N_6130);
xnor U6722 (N_6722,N_2531,N_2889);
and U6723 (N_6723,N_3888,N_3231);
nor U6724 (N_6724,N_2505,N_4655);
nor U6725 (N_6725,N_5775,N_2912);
and U6726 (N_6726,N_794,N_3827);
or U6727 (N_6727,N_1503,N_3266);
nand U6728 (N_6728,N_1710,N_4966);
and U6729 (N_6729,N_5935,N_3472);
nand U6730 (N_6730,N_4390,N_5937);
xnor U6731 (N_6731,N_2391,N_5596);
or U6732 (N_6732,N_4350,N_63);
or U6733 (N_6733,N_406,N_958);
nand U6734 (N_6734,N_211,N_3668);
xor U6735 (N_6735,N_5448,N_4947);
or U6736 (N_6736,N_2853,N_1558);
and U6737 (N_6737,N_2931,N_2);
xnor U6738 (N_6738,N_867,N_2727);
nor U6739 (N_6739,N_1160,N_4918);
nand U6740 (N_6740,N_5890,N_3862);
nand U6741 (N_6741,N_1000,N_1142);
and U6742 (N_6742,N_4915,N_1312);
and U6743 (N_6743,N_66,N_4371);
nand U6744 (N_6744,N_597,N_5966);
xor U6745 (N_6745,N_5618,N_4942);
nand U6746 (N_6746,N_4630,N_5275);
nor U6747 (N_6747,N_5606,N_2751);
or U6748 (N_6748,N_4784,N_4489);
nand U6749 (N_6749,N_1409,N_803);
or U6750 (N_6750,N_2077,N_3079);
nand U6751 (N_6751,N_5560,N_622);
nor U6752 (N_6752,N_3561,N_513);
or U6753 (N_6753,N_547,N_4584);
nor U6754 (N_6754,N_5572,N_3334);
nand U6755 (N_6755,N_1355,N_4029);
and U6756 (N_6756,N_5114,N_1430);
and U6757 (N_6757,N_1882,N_5373);
or U6758 (N_6758,N_6171,N_5335);
nand U6759 (N_6759,N_1250,N_1731);
or U6760 (N_6760,N_5053,N_2491);
nor U6761 (N_6761,N_3866,N_4186);
xnor U6762 (N_6762,N_3188,N_2175);
and U6763 (N_6763,N_4470,N_5724);
and U6764 (N_6764,N_4665,N_575);
or U6765 (N_6765,N_4156,N_3578);
nand U6766 (N_6766,N_4508,N_4496);
nor U6767 (N_6767,N_5682,N_1562);
xor U6768 (N_6768,N_852,N_1144);
nor U6769 (N_6769,N_4740,N_708);
nor U6770 (N_6770,N_2298,N_738);
xnor U6771 (N_6771,N_3899,N_906);
nand U6772 (N_6772,N_5294,N_3185);
or U6773 (N_6773,N_5305,N_5978);
nand U6774 (N_6774,N_6201,N_4499);
xor U6775 (N_6775,N_5597,N_5125);
nand U6776 (N_6776,N_5421,N_5998);
and U6777 (N_6777,N_5454,N_4709);
nor U6778 (N_6778,N_5075,N_3777);
or U6779 (N_6779,N_3238,N_4620);
nand U6780 (N_6780,N_3255,N_5018);
and U6781 (N_6781,N_3570,N_3820);
or U6782 (N_6782,N_370,N_3903);
nor U6783 (N_6783,N_3605,N_2429);
or U6784 (N_6784,N_1793,N_3598);
nand U6785 (N_6785,N_273,N_1366);
nand U6786 (N_6786,N_490,N_2081);
xnor U6787 (N_6787,N_681,N_1517);
or U6788 (N_6788,N_421,N_4808);
nand U6789 (N_6789,N_2916,N_6065);
xor U6790 (N_6790,N_1628,N_2934);
nor U6791 (N_6791,N_2005,N_4647);
nor U6792 (N_6792,N_4613,N_2068);
xor U6793 (N_6793,N_3302,N_317);
xnor U6794 (N_6794,N_910,N_161);
nor U6795 (N_6795,N_2230,N_1836);
nor U6796 (N_6796,N_2553,N_2224);
xnor U6797 (N_6797,N_154,N_6174);
or U6798 (N_6798,N_5110,N_2208);
xor U6799 (N_6799,N_6022,N_1608);
or U6800 (N_6800,N_5159,N_5939);
nand U6801 (N_6801,N_3404,N_2759);
xor U6802 (N_6802,N_3721,N_847);
and U6803 (N_6803,N_5359,N_3985);
and U6804 (N_6804,N_4659,N_799);
xnor U6805 (N_6805,N_5519,N_3625);
and U6806 (N_6806,N_510,N_4877);
and U6807 (N_6807,N_1962,N_4464);
or U6808 (N_6808,N_947,N_3791);
and U6809 (N_6809,N_4746,N_635);
nor U6810 (N_6810,N_5127,N_5526);
nor U6811 (N_6811,N_1211,N_1084);
nand U6812 (N_6812,N_1880,N_408);
nand U6813 (N_6813,N_1853,N_1009);
and U6814 (N_6814,N_1946,N_5814);
xnor U6815 (N_6815,N_2390,N_2983);
xnor U6816 (N_6816,N_5956,N_5620);
nand U6817 (N_6817,N_5845,N_1380);
and U6818 (N_6818,N_1617,N_4884);
nand U6819 (N_6819,N_3682,N_2072);
nand U6820 (N_6820,N_3530,N_2495);
nand U6821 (N_6821,N_2755,N_3498);
or U6822 (N_6822,N_1018,N_6085);
or U6823 (N_6823,N_773,N_68);
nor U6824 (N_6824,N_3133,N_2317);
or U6825 (N_6825,N_2761,N_4634);
nor U6826 (N_6826,N_301,N_4532);
nor U6827 (N_6827,N_2589,N_667);
nor U6828 (N_6828,N_5321,N_5513);
nand U6829 (N_6829,N_778,N_5593);
nand U6830 (N_6830,N_5182,N_5044);
xor U6831 (N_6831,N_4673,N_750);
nand U6832 (N_6832,N_619,N_697);
or U6833 (N_6833,N_3431,N_3476);
xnor U6834 (N_6834,N_5088,N_4310);
nand U6835 (N_6835,N_1815,N_4466);
nand U6836 (N_6836,N_3356,N_2848);
nand U6837 (N_6837,N_1902,N_3271);
or U6838 (N_6838,N_1590,N_325);
nor U6839 (N_6839,N_766,N_4710);
xnor U6840 (N_6840,N_2199,N_1894);
xor U6841 (N_6841,N_2650,N_6006);
nand U6842 (N_6842,N_4670,N_515);
or U6843 (N_6843,N_4723,N_638);
nor U6844 (N_6844,N_3413,N_4955);
nand U6845 (N_6845,N_5477,N_3863);
nand U6846 (N_6846,N_604,N_1143);
nand U6847 (N_6847,N_4642,N_3965);
or U6848 (N_6848,N_4133,N_3189);
nor U6849 (N_6849,N_3316,N_5452);
xor U6850 (N_6850,N_428,N_1074);
and U6851 (N_6851,N_1401,N_4327);
or U6852 (N_6852,N_5036,N_3046);
xnor U6853 (N_6853,N_4593,N_4216);
nand U6854 (N_6854,N_4684,N_5731);
or U6855 (N_6855,N_1246,N_3113);
or U6856 (N_6856,N_1943,N_447);
nand U6857 (N_6857,N_883,N_2907);
and U6858 (N_6858,N_414,N_4626);
xnor U6859 (N_6859,N_2144,N_5602);
or U6860 (N_6860,N_5860,N_4170);
nor U6861 (N_6861,N_4047,N_1295);
nand U6862 (N_6862,N_474,N_2052);
nand U6863 (N_6863,N_149,N_3542);
nor U6864 (N_6864,N_4158,N_4282);
or U6865 (N_6865,N_1770,N_5200);
and U6866 (N_6866,N_2797,N_2623);
xnor U6867 (N_6867,N_850,N_1007);
nand U6868 (N_6868,N_3150,N_1916);
nand U6869 (N_6869,N_4252,N_1549);
nor U6870 (N_6870,N_4289,N_623);
nand U6871 (N_6871,N_36,N_3698);
nor U6872 (N_6872,N_1222,N_5551);
and U6873 (N_6873,N_4084,N_4656);
nand U6874 (N_6874,N_764,N_1774);
and U6875 (N_6875,N_2694,N_4086);
or U6876 (N_6876,N_1540,N_1498);
xnor U6877 (N_6877,N_1393,N_1528);
or U6878 (N_6878,N_922,N_696);
and U6879 (N_6879,N_1204,N_2257);
nand U6880 (N_6880,N_6210,N_889);
xnor U6881 (N_6881,N_5758,N_6080);
and U6882 (N_6882,N_6072,N_4424);
nand U6883 (N_6883,N_1480,N_3583);
and U6884 (N_6884,N_4867,N_5194);
and U6885 (N_6885,N_507,N_200);
xnor U6886 (N_6886,N_6173,N_2993);
and U6887 (N_6887,N_1030,N_1452);
nand U6888 (N_6888,N_579,N_342);
xor U6889 (N_6889,N_2709,N_2582);
or U6890 (N_6890,N_2841,N_1039);
xnor U6891 (N_6891,N_3912,N_1846);
and U6892 (N_6892,N_3939,N_3366);
nand U6893 (N_6893,N_332,N_1543);
nand U6894 (N_6894,N_6033,N_1953);
nand U6895 (N_6895,N_1324,N_5478);
xor U6896 (N_6896,N_286,N_2362);
nor U6897 (N_6897,N_4394,N_6158);
nor U6898 (N_6898,N_3246,N_2020);
and U6899 (N_6899,N_3824,N_5241);
and U6900 (N_6900,N_1941,N_3538);
xnor U6901 (N_6901,N_2188,N_3184);
and U6902 (N_6902,N_569,N_4183);
xnor U6903 (N_6903,N_3068,N_1416);
xnor U6904 (N_6904,N_3585,N_5588);
xnor U6905 (N_6905,N_5483,N_2791);
xnor U6906 (N_6906,N_4102,N_4008);
or U6907 (N_6907,N_3801,N_3974);
and U6908 (N_6908,N_138,N_1215);
or U6909 (N_6909,N_4501,N_473);
nor U6910 (N_6910,N_5915,N_1391);
nor U6911 (N_6911,N_4138,N_1635);
nand U6912 (N_6912,N_572,N_1200);
xnor U6913 (N_6913,N_1816,N_4941);
nand U6914 (N_6914,N_4845,N_1286);
or U6915 (N_6915,N_3636,N_4569);
nor U6916 (N_6916,N_6211,N_2309);
xnor U6917 (N_6917,N_2484,N_6189);
and U6918 (N_6918,N_5023,N_1004);
nor U6919 (N_6919,N_3953,N_4858);
xor U6920 (N_6920,N_646,N_5026);
and U6921 (N_6921,N_3126,N_4881);
nand U6922 (N_6922,N_4652,N_361);
nor U6923 (N_6923,N_1070,N_1197);
and U6924 (N_6924,N_2347,N_4423);
nor U6925 (N_6925,N_3632,N_3156);
nand U6926 (N_6926,N_4195,N_4136);
nor U6927 (N_6927,N_4564,N_5111);
or U6928 (N_6928,N_5287,N_4907);
nor U6929 (N_6929,N_5648,N_1799);
nor U6930 (N_6930,N_3552,N_5151);
nor U6931 (N_6931,N_4972,N_6137);
and U6932 (N_6932,N_2369,N_3751);
or U6933 (N_6933,N_4126,N_4384);
nand U6934 (N_6934,N_3095,N_4497);
xnor U6935 (N_6935,N_1552,N_3781);
nor U6936 (N_6936,N_5557,N_2094);
and U6937 (N_6937,N_3234,N_1618);
xor U6938 (N_6938,N_4991,N_1545);
or U6939 (N_6939,N_4108,N_6124);
nand U6940 (N_6940,N_1810,N_1867);
nand U6941 (N_6941,N_5010,N_4759);
nand U6942 (N_6942,N_5397,N_1386);
nor U6943 (N_6943,N_4859,N_2413);
or U6944 (N_6944,N_5196,N_5796);
xor U6945 (N_6945,N_2147,N_443);
or U6946 (N_6946,N_2657,N_2739);
and U6947 (N_6947,N_4246,N_5579);
nor U6948 (N_6948,N_88,N_893);
nand U6949 (N_6949,N_20,N_5163);
xnor U6950 (N_6950,N_2771,N_1003);
nand U6951 (N_6951,N_3327,N_2132);
nand U6952 (N_6952,N_2478,N_1614);
nand U6953 (N_6953,N_4205,N_3917);
nand U6954 (N_6954,N_4492,N_3417);
nand U6955 (N_6955,N_6209,N_3343);
and U6956 (N_6956,N_3607,N_797);
nor U6957 (N_6957,N_3517,N_1365);
xor U6958 (N_6958,N_2452,N_3686);
nor U6959 (N_6959,N_1818,N_1455);
xor U6960 (N_6960,N_4787,N_5536);
and U6961 (N_6961,N_5970,N_767);
nand U6962 (N_6962,N_333,N_5506);
or U6963 (N_6963,N_405,N_1505);
nand U6964 (N_6964,N_699,N_968);
or U6965 (N_6965,N_6002,N_1153);
nand U6966 (N_6966,N_2870,N_2425);
nor U6967 (N_6967,N_4436,N_1871);
xnor U6968 (N_6968,N_4791,N_1611);
nand U6969 (N_6969,N_1068,N_4810);
nand U6970 (N_6970,N_5510,N_4660);
nand U6971 (N_6971,N_4155,N_1660);
xor U6972 (N_6972,N_1744,N_3445);
nand U6973 (N_6973,N_3136,N_5198);
nand U6974 (N_6974,N_6245,N_5175);
and U6975 (N_6975,N_2141,N_4241);
nor U6976 (N_6976,N_1047,N_1716);
or U6977 (N_6977,N_5678,N_3993);
or U6978 (N_6978,N_2282,N_3581);
nor U6979 (N_6979,N_2783,N_451);
or U6980 (N_6980,N_2702,N_990);
and U6981 (N_6981,N_511,N_1692);
xor U6982 (N_6982,N_5607,N_2740);
nor U6983 (N_6983,N_4050,N_1497);
and U6984 (N_6984,N_2033,N_4568);
and U6985 (N_6985,N_2651,N_5191);
nor U6986 (N_6986,N_1796,N_3706);
or U6987 (N_6987,N_4068,N_5903);
nand U6988 (N_6988,N_481,N_1438);
xnor U6989 (N_6989,N_364,N_4432);
and U6990 (N_6990,N_2346,N_5195);
or U6991 (N_6991,N_5962,N_2327);
or U6992 (N_6992,N_6183,N_1462);
xor U6993 (N_6993,N_2383,N_2125);
and U6994 (N_6994,N_1668,N_1002);
xor U6995 (N_6995,N_795,N_1336);
nand U6996 (N_6996,N_5039,N_1535);
nor U6997 (N_6997,N_5530,N_247);
nor U6998 (N_6998,N_964,N_4961);
xor U6999 (N_6999,N_6066,N_1714);
nand U7000 (N_7000,N_2274,N_4169);
nand U7001 (N_7001,N_788,N_6017);
xnor U7002 (N_7002,N_586,N_2754);
or U7003 (N_7003,N_1856,N_4344);
and U7004 (N_7004,N_162,N_1298);
and U7005 (N_7005,N_5960,N_5610);
or U7006 (N_7006,N_5290,N_1878);
or U7007 (N_7007,N_4341,N_5614);
xnor U7008 (N_7008,N_745,N_4256);
xor U7009 (N_7009,N_4261,N_5068);
nand U7010 (N_7010,N_5,N_6135);
nand U7011 (N_7011,N_6241,N_2913);
xnor U7012 (N_7012,N_4001,N_3527);
nor U7013 (N_7013,N_1828,N_5012);
nor U7014 (N_7014,N_4381,N_3715);
or U7015 (N_7015,N_5462,N_2729);
nand U7016 (N_7016,N_5556,N_3100);
nand U7017 (N_7017,N_1814,N_174);
nand U7018 (N_7018,N_617,N_5124);
xor U7019 (N_7019,N_3614,N_3717);
nor U7020 (N_7020,N_5803,N_3442);
nor U7021 (N_7021,N_4437,N_1469);
nor U7022 (N_7022,N_4286,N_2370);
nor U7023 (N_7023,N_2725,N_1809);
nor U7024 (N_7024,N_1299,N_4798);
nor U7025 (N_7025,N_3712,N_1076);
or U7026 (N_7026,N_3322,N_2035);
nor U7027 (N_7027,N_1383,N_1369);
nand U7028 (N_7028,N_4257,N_2361);
nand U7029 (N_7029,N_4958,N_3742);
nand U7030 (N_7030,N_2302,N_2028);
nand U7031 (N_7031,N_5749,N_5304);
or U7032 (N_7032,N_1173,N_3811);
or U7033 (N_7033,N_6208,N_14);
nand U7034 (N_7034,N_15,N_1584);
nor U7035 (N_7035,N_4678,N_3145);
nand U7036 (N_7036,N_2371,N_5670);
or U7037 (N_7037,N_5310,N_3723);
or U7038 (N_7038,N_3219,N_1771);
nor U7039 (N_7039,N_2613,N_440);
nor U7040 (N_7040,N_5825,N_85);
xnor U7041 (N_7041,N_5383,N_3595);
and U7042 (N_7042,N_2758,N_4616);
xor U7043 (N_7043,N_835,N_4132);
or U7044 (N_7044,N_4431,N_588);
and U7045 (N_7045,N_438,N_292);
nor U7046 (N_7046,N_5570,N_6187);
nand U7047 (N_7047,N_913,N_4728);
nor U7048 (N_7048,N_137,N_2288);
nand U7049 (N_7049,N_5784,N_2229);
and U7050 (N_7050,N_5767,N_6031);
nand U7051 (N_7051,N_5655,N_2251);
nor U7052 (N_7052,N_128,N_1446);
or U7053 (N_7053,N_4937,N_3101);
nand U7054 (N_7054,N_994,N_5561);
nand U7055 (N_7055,N_975,N_1101);
or U7056 (N_7056,N_5208,N_5184);
nand U7057 (N_7057,N_3013,N_5491);
xor U7058 (N_7058,N_6030,N_4114);
nor U7059 (N_7059,N_4631,N_2543);
or U7060 (N_7060,N_1980,N_4348);
or U7061 (N_7061,N_3693,N_3032);
xnor U7062 (N_7062,N_1235,N_3840);
nand U7063 (N_7063,N_2875,N_519);
nor U7064 (N_7064,N_965,N_2305);
xnor U7065 (N_7065,N_2297,N_4543);
nand U7066 (N_7066,N_4931,N_1798);
nor U7067 (N_7067,N_3,N_5153);
nor U7068 (N_7068,N_1042,N_1896);
nand U7069 (N_7069,N_4895,N_6039);
or U7070 (N_7070,N_1857,N_391);
nor U7071 (N_7071,N_881,N_1512);
or U7072 (N_7072,N_27,N_1595);
and U7073 (N_7073,N_567,N_4648);
and U7074 (N_7074,N_1465,N_3834);
nor U7075 (N_7075,N_729,N_4747);
nor U7076 (N_7076,N_1489,N_3066);
nand U7077 (N_7077,N_4228,N_23);
nor U7078 (N_7078,N_1787,N_5899);
or U7079 (N_7079,N_2753,N_1031);
and U7080 (N_7080,N_4352,N_1524);
and U7081 (N_7081,N_1937,N_4159);
or U7082 (N_7082,N_4541,N_3772);
nand U7083 (N_7083,N_1399,N_6015);
xnor U7084 (N_7084,N_2547,N_5371);
xnor U7085 (N_7085,N_3301,N_5719);
nor U7086 (N_7086,N_740,N_1593);
nor U7087 (N_7087,N_4556,N_5269);
nand U7088 (N_7088,N_4592,N_6142);
or U7089 (N_7089,N_3423,N_303);
nor U7090 (N_7090,N_318,N_4288);
and U7091 (N_7091,N_445,N_4802);
xnor U7092 (N_7092,N_3251,N_4632);
nor U7093 (N_7093,N_5711,N_1208);
nand U7094 (N_7094,N_1340,N_5360);
xor U7095 (N_7095,N_6219,N_4326);
and U7096 (N_7096,N_1749,N_5457);
and U7097 (N_7097,N_1170,N_132);
or U7098 (N_7098,N_4160,N_2940);
nor U7099 (N_7099,N_5280,N_1527);
or U7100 (N_7100,N_2198,N_1978);
and U7101 (N_7101,N_3354,N_5600);
or U7102 (N_7102,N_1897,N_1064);
nor U7103 (N_7103,N_26,N_525);
nand U7104 (N_7104,N_898,N_1585);
and U7105 (N_7105,N_96,N_4099);
nor U7106 (N_7106,N_2323,N_294);
or U7107 (N_7107,N_5985,N_4668);
nand U7108 (N_7108,N_555,N_5865);
and U7109 (N_7109,N_127,N_5134);
and U7110 (N_7110,N_3856,N_5862);
nor U7111 (N_7111,N_2157,N_5340);
nand U7112 (N_7112,N_5855,N_5544);
nor U7113 (N_7113,N_4220,N_2239);
or U7114 (N_7114,N_1351,N_5214);
and U7115 (N_7115,N_5129,N_986);
nand U7116 (N_7116,N_2382,N_5015);
or U7117 (N_7117,N_5174,N_501);
or U7118 (N_7118,N_2643,N_6176);
and U7119 (N_7119,N_2063,N_1790);
or U7120 (N_7120,N_1141,N_5625);
nor U7121 (N_7121,N_870,N_4298);
nor U7122 (N_7122,N_130,N_4588);
nor U7123 (N_7123,N_4254,N_1531);
xor U7124 (N_7124,N_259,N_468);
or U7125 (N_7125,N_4380,N_4333);
xor U7126 (N_7126,N_4193,N_3793);
nor U7127 (N_7127,N_2258,N_932);
nand U7128 (N_7128,N_2683,N_4285);
and U7129 (N_7129,N_4916,N_2550);
nand U7130 (N_7130,N_2546,N_2447);
and U7131 (N_7131,N_2624,N_5265);
and U7132 (N_7132,N_1083,N_1413);
and U7133 (N_7133,N_4044,N_6100);
nand U7134 (N_7134,N_4447,N_1556);
nand U7135 (N_7135,N_5599,N_4119);
and U7136 (N_7136,N_2585,N_3818);
nand U7137 (N_7137,N_5499,N_1907);
nand U7138 (N_7138,N_3894,N_2102);
or U7139 (N_7139,N_3124,N_5794);
or U7140 (N_7140,N_4396,N_1346);
xor U7141 (N_7141,N_1777,N_454);
and U7142 (N_7142,N_4913,N_1936);
and U7143 (N_7143,N_5930,N_226);
xnor U7144 (N_7144,N_1428,N_4296);
or U7145 (N_7145,N_5539,N_1768);
xor U7146 (N_7146,N_5730,N_4070);
or U7147 (N_7147,N_3787,N_2113);
or U7148 (N_7148,N_4518,N_1478);
nand U7149 (N_7149,N_441,N_4768);
xnor U7150 (N_7150,N_3617,N_420);
and U7151 (N_7151,N_4319,N_5239);
or U7152 (N_7152,N_5387,N_4871);
nand U7153 (N_7153,N_5035,N_5021);
nand U7154 (N_7154,N_1942,N_2630);
and U7155 (N_7155,N_1283,N_2308);
nand U7156 (N_7156,N_721,N_483);
nand U7157 (N_7157,N_1765,N_3277);
nor U7158 (N_7158,N_1107,N_5395);
nand U7159 (N_7159,N_1248,N_812);
xnor U7160 (N_7160,N_4674,N_1868);
or U7161 (N_7161,N_682,N_1747);
nand U7162 (N_7162,N_1406,N_5386);
and U7163 (N_7163,N_3989,N_337);
xnor U7164 (N_7164,N_2903,N_51);
nand U7165 (N_7165,N_3187,N_4763);
nand U7166 (N_7166,N_4772,N_3665);
nand U7167 (N_7167,N_340,N_1014);
or U7168 (N_7168,N_5476,N_5057);
and U7169 (N_7169,N_2177,N_3395);
or U7170 (N_7170,N_92,N_3351);
and U7171 (N_7171,N_1602,N_5894);
nor U7172 (N_7172,N_2289,N_2340);
xor U7173 (N_7173,N_1236,N_3602);
nor U7174 (N_7174,N_4173,N_4405);
nand U7175 (N_7175,N_6087,N_1597);
xnor U7176 (N_7176,N_4342,N_1723);
and U7177 (N_7177,N_524,N_5696);
xor U7178 (N_7178,N_2874,N_4018);
xor U7179 (N_7179,N_1743,N_2064);
xnor U7180 (N_7180,N_6067,N_2946);
and U7181 (N_7181,N_1495,N_4795);
nand U7182 (N_7182,N_819,N_2241);
and U7183 (N_7183,N_5404,N_5299);
nor U7184 (N_7184,N_5094,N_4677);
or U7185 (N_7185,N_5399,N_4713);
or U7186 (N_7186,N_1782,N_1539);
and U7187 (N_7187,N_1112,N_3168);
or U7188 (N_7188,N_6204,N_4914);
xnor U7189 (N_7189,N_2818,N_2539);
nor U7190 (N_7190,N_374,N_395);
or U7191 (N_7191,N_4559,N_3898);
nand U7192 (N_7192,N_4105,N_1870);
or U7193 (N_7193,N_3724,N_5559);
nor U7194 (N_7194,N_5876,N_2118);
nor U7195 (N_7195,N_2721,N_5518);
xor U7196 (N_7196,N_2043,N_2159);
or U7197 (N_7197,N_2796,N_5815);
nor U7198 (N_7198,N_4928,N_5245);
xnor U7199 (N_7199,N_5712,N_5961);
or U7200 (N_7200,N_4011,N_1025);
nor U7201 (N_7201,N_4535,N_383);
xor U7202 (N_7202,N_3785,N_2356);
nand U7203 (N_7203,N_1767,N_5640);
or U7204 (N_7204,N_4179,N_32);
nand U7205 (N_7205,N_5770,N_3242);
and U7206 (N_7206,N_205,N_5866);
nor U7207 (N_7207,N_6144,N_955);
nand U7208 (N_7208,N_4265,N_4428);
nand U7209 (N_7209,N_22,N_3026);
or U7210 (N_7210,N_1609,N_2250);
nor U7211 (N_7211,N_3537,N_4395);
or U7212 (N_7212,N_1892,N_5924);
nand U7213 (N_7213,N_3761,N_879);
and U7214 (N_7214,N_5659,N_95);
and U7215 (N_7215,N_3901,N_6055);
xnor U7216 (N_7216,N_2649,N_4989);
xnor U7217 (N_7217,N_2410,N_1314);
xnor U7218 (N_7218,N_4849,N_160);
or U7219 (N_7219,N_2187,N_608);
or U7220 (N_7220,N_4052,N_5830);
nor U7221 (N_7221,N_5885,N_3003);
or U7222 (N_7222,N_5656,N_1672);
xnor U7223 (N_7223,N_2817,N_2191);
xnor U7224 (N_7224,N_4500,N_2833);
and U7225 (N_7225,N_3756,N_4059);
xnor U7226 (N_7226,N_4734,N_2558);
or U7227 (N_7227,N_600,N_2938);
xnor U7228 (N_7228,N_290,N_4204);
or U7229 (N_7229,N_3409,N_6131);
nor U7230 (N_7230,N_2088,N_3995);
nand U7231 (N_7231,N_1108,N_5409);
or U7232 (N_7232,N_915,N_4181);
nand U7233 (N_7233,N_3587,N_1012);
or U7234 (N_7234,N_4530,N_5363);
or U7235 (N_7235,N_3298,N_93);
nor U7236 (N_7236,N_3483,N_5954);
and U7237 (N_7237,N_549,N_2217);
xnor U7238 (N_7238,N_4549,N_1317);
nor U7239 (N_7239,N_3310,N_2419);
xnor U7240 (N_7240,N_2232,N_3631);
or U7241 (N_7241,N_3575,N_1769);
xnor U7242 (N_7242,N_1165,N_1982);
and U7243 (N_7243,N_938,N_551);
xor U7244 (N_7244,N_5225,N_3482);
nor U7245 (N_7245,N_4063,N_1251);
or U7246 (N_7246,N_4843,N_706);
or U7247 (N_7247,N_5158,N_3025);
nor U7248 (N_7248,N_4399,N_1993);
nor U7249 (N_7249,N_1589,N_4293);
xnor U7250 (N_7250,N_4411,N_5888);
nor U7251 (N_7251,N_2059,N_5230);
xnor U7252 (N_7252,N_3192,N_3873);
nand U7253 (N_7253,N_3759,N_4426);
xor U7254 (N_7254,N_2213,N_6139);
nand U7255 (N_7255,N_1069,N_2884);
or U7256 (N_7256,N_4493,N_477);
nor U7257 (N_7257,N_3368,N_4528);
and U7258 (N_7258,N_4312,N_2065);
xnor U7259 (N_7259,N_5698,N_5141);
xor U7260 (N_7260,N_2855,N_1625);
xnor U7261 (N_7261,N_1945,N_2286);
xor U7262 (N_7262,N_3627,N_3885);
and U7263 (N_7263,N_1933,N_2403);
and U7264 (N_7264,N_5887,N_3336);
nand U7265 (N_7265,N_4586,N_5810);
nand U7266 (N_7266,N_2615,N_1467);
nand U7267 (N_7267,N_4582,N_4685);
and U7268 (N_7268,N_1347,N_5201);
and U7269 (N_7269,N_3324,N_3563);
xor U7270 (N_7270,N_1719,N_2354);
xor U7271 (N_7271,N_2075,N_2635);
xnor U7272 (N_7272,N_235,N_5928);
xnor U7273 (N_7273,N_76,N_4993);
and U7274 (N_7274,N_4071,N_5276);
and U7275 (N_7275,N_6020,N_2900);
xor U7276 (N_7276,N_1491,N_4504);
and U7277 (N_7277,N_1449,N_5905);
and U7278 (N_7278,N_1261,N_2661);
or U7279 (N_7279,N_6123,N_4885);
xnor U7280 (N_7280,N_5651,N_912);
xnor U7281 (N_7281,N_4936,N_6025);
nor U7282 (N_7282,N_3593,N_3813);
and U7283 (N_7283,N_2089,N_4570);
nor U7284 (N_7284,N_3853,N_5362);
and U7285 (N_7285,N_858,N_3317);
xor U7286 (N_7286,N_6090,N_4963);
or U7287 (N_7287,N_749,N_843);
or U7288 (N_7288,N_327,N_5755);
or U7289 (N_7289,N_3944,N_4754);
or U7290 (N_7290,N_3677,N_3857);
and U7291 (N_7291,N_2279,N_3544);
xnor U7292 (N_7292,N_3800,N_5797);
xnor U7293 (N_7293,N_2569,N_2280);
xnor U7294 (N_7294,N_1951,N_5766);
or U7295 (N_7295,N_3342,N_1424);
and U7296 (N_7296,N_5674,N_257);
or U7297 (N_7297,N_5984,N_2600);
xor U7298 (N_7298,N_5707,N_6054);
or U7299 (N_7299,N_458,N_2314);
or U7300 (N_7300,N_230,N_3622);
or U7301 (N_7301,N_1740,N_4601);
nor U7302 (N_7302,N_2955,N_3457);
nand U7303 (N_7303,N_3577,N_1051);
or U7304 (N_7304,N_4646,N_2019);
xnor U7305 (N_7305,N_4188,N_2793);
nor U7306 (N_7306,N_3127,N_4525);
or U7307 (N_7307,N_5617,N_1095);
and U7308 (N_7308,N_832,N_4608);
xor U7309 (N_7309,N_3661,N_2322);
and U7310 (N_7310,N_3523,N_4276);
nor U7311 (N_7311,N_3829,N_5032);
nor U7312 (N_7312,N_5389,N_4299);
xnor U7313 (N_7313,N_3051,N_1091);
or U7314 (N_7314,N_1010,N_2996);
nor U7315 (N_7315,N_3144,N_1506);
nand U7316 (N_7316,N_2328,N_2284);
xnor U7317 (N_7317,N_4940,N_4873);
nand U7318 (N_7318,N_3217,N_3000);
xnor U7319 (N_7319,N_3325,N_4375);
and U7320 (N_7320,N_2137,N_4255);
xnor U7321 (N_7321,N_5309,N_948);
or U7322 (N_7322,N_2893,N_436);
or U7323 (N_7323,N_1359,N_2190);
nand U7324 (N_7324,N_378,N_5516);
and U7325 (N_7325,N_2145,N_4382);
and U7326 (N_7326,N_1062,N_3008);
xnor U7327 (N_7327,N_4401,N_2501);
and U7328 (N_7328,N_2482,N_245);
and U7329 (N_7329,N_1854,N_587);
nor U7330 (N_7330,N_576,N_4349);
xor U7331 (N_7331,N_1110,N_781);
nand U7332 (N_7332,N_2392,N_6003);
xnor U7333 (N_7333,N_1045,N_343);
nand U7334 (N_7334,N_5986,N_946);
or U7335 (N_7335,N_3253,N_3730);
xnor U7336 (N_7336,N_121,N_2548);
nand U7337 (N_7337,N_1313,N_3250);
nand U7338 (N_7338,N_5503,N_730);
nor U7339 (N_7339,N_1460,N_4328);
xnor U7340 (N_7340,N_3049,N_5252);
xor U7341 (N_7341,N_1872,N_2430);
and U7342 (N_7342,N_360,N_1490);
nand U7343 (N_7343,N_4019,N_1225);
xnor U7344 (N_7344,N_2222,N_2253);
and U7345 (N_7345,N_4896,N_4978);
xnor U7346 (N_7346,N_3180,N_4804);
xnor U7347 (N_7347,N_3762,N_4888);
or U7348 (N_7348,N_2227,N_4056);
nand U7349 (N_7349,N_4368,N_1422);
xor U7350 (N_7350,N_2652,N_4128);
and U7351 (N_7351,N_533,N_4834);
or U7352 (N_7352,N_2986,N_903);
nand U7353 (N_7353,N_2311,N_3909);
or U7354 (N_7354,N_723,N_2245);
xor U7355 (N_7355,N_1106,N_2628);
nor U7356 (N_7356,N_5524,N_5922);
xnor U7357 (N_7357,N_6107,N_73);
or U7358 (N_7358,N_5820,N_5662);
or U7359 (N_7359,N_2149,N_1813);
xor U7360 (N_7360,N_535,N_1574);
nand U7361 (N_7361,N_4127,N_4408);
xor U7362 (N_7362,N_1974,N_2333);
or U7363 (N_7363,N_3390,N_1601);
nand U7364 (N_7364,N_4406,N_725);
nand U7365 (N_7365,N_4743,N_5001);
or U7366 (N_7366,N_5017,N_4527);
nor U7367 (N_7367,N_3411,N_3646);
nor U7368 (N_7368,N_1570,N_6012);
or U7369 (N_7369,N_5693,N_4855);
nand U7370 (N_7370,N_5792,N_4354);
nand U7371 (N_7371,N_3073,N_5795);
or U7372 (N_7372,N_1538,N_2598);
and U7373 (N_7373,N_1772,N_320);
nor U7374 (N_7374,N_5259,N_839);
nand U7375 (N_7375,N_4219,N_5827);
xor U7376 (N_7376,N_2235,N_4562);
or U7377 (N_7377,N_3347,N_1499);
or U7378 (N_7378,N_3941,N_3286);
and U7379 (N_7379,N_5522,N_4835);
nand U7380 (N_7380,N_2161,N_2567);
nand U7381 (N_7381,N_5594,N_5949);
xor U7382 (N_7382,N_844,N_3515);
and U7383 (N_7383,N_2416,N_3594);
xor U7384 (N_7384,N_3494,N_5615);
and U7385 (N_7385,N_3503,N_216);
and U7386 (N_7386,N_1550,N_3330);
nor U7387 (N_7387,N_287,N_5619);
or U7388 (N_7388,N_802,N_6138);
xnor U7389 (N_7389,N_4283,N_1530);
nor U7390 (N_7390,N_4857,N_4628);
xnor U7391 (N_7391,N_5893,N_3852);
or U7392 (N_7392,N_4548,N_4946);
nand U7393 (N_7393,N_5369,N_5508);
or U7394 (N_7394,N_2723,N_2659);
nor U7395 (N_7395,N_464,N_484);
or U7396 (N_7396,N_1214,N_4813);
nand U7397 (N_7397,N_4151,N_452);
nor U7398 (N_7398,N_5722,N_2130);
and U7399 (N_7399,N_5227,N_3027);
or U7400 (N_7400,N_5987,N_1258);
xnor U7401 (N_7401,N_4230,N_2339);
nor U7402 (N_7402,N_3741,N_5019);
nand U7403 (N_7403,N_456,N_2474);
nand U7404 (N_7404,N_3590,N_2471);
and U7405 (N_7405,N_1109,N_3652);
nand U7406 (N_7406,N_4547,N_3364);
nor U7407 (N_7407,N_4641,N_4774);
or U7408 (N_7408,N_1845,N_3380);
and U7409 (N_7409,N_4313,N_4698);
or U7410 (N_7410,N_208,N_3553);
or U7411 (N_7411,N_5641,N_231);
nand U7412 (N_7412,N_5128,N_988);
nor U7413 (N_7413,N_2399,N_3620);
nand U7414 (N_7414,N_1191,N_5558);
xor U7415 (N_7415,N_5878,N_4682);
xnor U7416 (N_7416,N_1238,N_4992);
and U7417 (N_7417,N_4323,N_3140);
and U7418 (N_7418,N_2828,N_285);
nor U7419 (N_7419,N_3568,N_920);
and U7420 (N_7420,N_5709,N_5463);
nand U7421 (N_7421,N_4197,N_2706);
nor U7422 (N_7422,N_1130,N_4998);
nand U7423 (N_7423,N_2260,N_3203);
nor U7424 (N_7424,N_1651,N_119);
nor U7425 (N_7425,N_1218,N_5300);
xor U7426 (N_7426,N_1579,N_4612);
and U7427 (N_7427,N_4836,N_5066);
or U7428 (N_7428,N_2060,N_3182);
nand U7429 (N_7429,N_3112,N_4705);
or U7430 (N_7430,N_5405,N_2678);
xnor U7431 (N_7431,N_937,N_1848);
xnor U7432 (N_7432,N_6083,N_4676);
and U7433 (N_7433,N_4650,N_613);
xor U7434 (N_7434,N_4891,N_2070);
and U7435 (N_7435,N_190,N_2176);
or U7436 (N_7436,N_680,N_1507);
and U7437 (N_7437,N_4079,N_5097);
or U7438 (N_7438,N_2952,N_1823);
and U7439 (N_7439,N_1862,N_901);
xor U7440 (N_7440,N_552,N_5365);
xor U7441 (N_7441,N_3934,N_1630);
nor U7442 (N_7442,N_3022,N_6200);
or U7443 (N_7443,N_2746,N_2756);
nor U7444 (N_7444,N_5281,N_1382);
nor U7445 (N_7445,N_2696,N_1118);
or U7446 (N_7446,N_3157,N_3550);
and U7447 (N_7447,N_1778,N_210);
nand U7448 (N_7448,N_5902,N_2026);
or U7449 (N_7449,N_1137,N_2195);
or U7450 (N_7450,N_5133,N_485);
nand U7451 (N_7451,N_1526,N_5132);
or U7452 (N_7452,N_3375,N_2332);
nor U7453 (N_7453,N_1027,N_5990);
nor U7454 (N_7454,N_1022,N_3070);
xnor U7455 (N_7455,N_1721,N_19);
nor U7456 (N_7456,N_2811,N_3814);
and U7457 (N_7457,N_1827,N_4597);
xor U7458 (N_7458,N_2570,N_3750);
nor U7459 (N_7459,N_539,N_5553);
or U7460 (N_7460,N_936,N_953);
or U7461 (N_7461,N_2563,N_5571);
xnor U7462 (N_7462,N_5765,N_4781);
xor U7463 (N_7463,N_5715,N_5868);
and U7464 (N_7464,N_4118,N_5762);
nand U7465 (N_7465,N_1453,N_3321);
and U7466 (N_7466,N_6141,N_1544);
nand U7467 (N_7467,N_5343,N_3285);
nor U7468 (N_7468,N_3358,N_1825);
nor U7469 (N_7469,N_4386,N_151);
and U7470 (N_7470,N_3102,N_3452);
nand U7471 (N_7471,N_5183,N_4430);
nand U7472 (N_7472,N_272,N_1237);
or U7473 (N_7473,N_2032,N_929);
nand U7474 (N_7474,N_1674,N_3290);
xnor U7475 (N_7475,N_6092,N_5331);
xnor U7476 (N_7476,N_314,N_3861);
xnor U7477 (N_7477,N_775,N_3589);
nor U7478 (N_7478,N_2384,N_1709);
and U7479 (N_7479,N_328,N_1180);
or U7480 (N_7480,N_853,N_5509);
or U7481 (N_7481,N_4206,N_59);
nor U7482 (N_7482,N_3397,N_4622);
and U7483 (N_7483,N_3461,N_5881);
xor U7484 (N_7484,N_3331,N_3034);
nand U7485 (N_7485,N_4165,N_1203);
and U7486 (N_7486,N_2541,N_1802);
xnor U7487 (N_7487,N_1580,N_55);
nor U7488 (N_7488,N_6036,N_2182);
nand U7489 (N_7489,N_2883,N_97);
xnor U7490 (N_7490,N_5507,N_4680);
xnor U7491 (N_7491,N_5353,N_3826);
nand U7492 (N_7492,N_156,N_2415);
xnor U7493 (N_7493,N_5266,N_5757);
nand U7494 (N_7494,N_5203,N_2960);
and U7495 (N_7495,N_3481,N_2270);
nand U7496 (N_7496,N_352,N_2324);
xor U7497 (N_7497,N_1607,N_2768);
nand U7498 (N_7498,N_4345,N_1209);
nand U7499 (N_7499,N_3296,N_4243);
or U7500 (N_7500,N_2902,N_5357);
nor U7501 (N_7501,N_2504,N_434);
xnor U7502 (N_7502,N_4765,N_4794);
xnor U7503 (N_7503,N_5157,N_2029);
xor U7504 (N_7504,N_5475,N_2572);
and U7505 (N_7505,N_5679,N_217);
xnor U7506 (N_7506,N_5799,N_2171);
and U7507 (N_7507,N_4400,N_478);
nand U7508 (N_7508,N_6042,N_6213);
nor U7509 (N_7509,N_945,N_1833);
or U7510 (N_7510,N_5009,N_5500);
xnor U7511 (N_7511,N_86,N_4517);
and U7512 (N_7512,N_4686,N_209);
or U7513 (N_7513,N_4538,N_2614);
nand U7514 (N_7514,N_207,N_1308);
or U7515 (N_7515,N_2982,N_330);
nand U7516 (N_7516,N_6069,N_505);
xor U7517 (N_7517,N_6018,N_981);
or U7518 (N_7518,N_2012,N_2126);
nand U7519 (N_7519,N_3345,N_5372);
nor U7520 (N_7520,N_6214,N_2313);
nand U7521 (N_7521,N_2054,N_4191);
and U7522 (N_7522,N_4140,N_2423);
or U7523 (N_7523,N_3487,N_5040);
nand U7524 (N_7524,N_4692,N_626);
xnor U7525 (N_7525,N_1915,N_5901);
and U7526 (N_7526,N_5952,N_5234);
nor U7527 (N_7527,N_4605,N_1860);
xnor U7528 (N_7528,N_3104,N_6034);
or U7529 (N_7529,N_1753,N_4391);
nor U7530 (N_7530,N_2494,N_2644);
xor U7531 (N_7531,N_3775,N_1016);
nand U7532 (N_7532,N_6203,N_1318);
nor U7533 (N_7533,N_1356,N_1758);
or U7534 (N_7534,N_4112,N_4957);
nand U7535 (N_7535,N_4061,N_5816);
xor U7536 (N_7536,N_2071,N_2124);
and U7537 (N_7537,N_4999,N_648);
or U7538 (N_7538,N_578,N_5288);
nand U7539 (N_7539,N_5031,N_2008);
nor U7540 (N_7540,N_1541,N_2837);
nor U7541 (N_7541,N_1210,N_3558);
and U7542 (N_7542,N_4215,N_3412);
nand U7543 (N_7543,N_4014,N_5277);
nand U7544 (N_7544,N_4272,N_4832);
and U7545 (N_7545,N_793,N_168);
nand U7546 (N_7546,N_2487,N_1598);
nor U7547 (N_7547,N_12,N_5964);
and U7548 (N_7548,N_6249,N_1594);
nand U7549 (N_7549,N_3815,N_1307);
xnor U7550 (N_7550,N_4135,N_1481);
nor U7551 (N_7551,N_548,N_1729);
or U7552 (N_7552,N_3647,N_4758);
or U7553 (N_7553,N_3640,N_2151);
or U7554 (N_7554,N_4921,N_5432);
xnor U7555 (N_7555,N_5000,N_5637);
nor U7556 (N_7556,N_809,N_6119);
or U7557 (N_7557,N_5550,N_1789);
xor U7558 (N_7558,N_3513,N_398);
xor U7559 (N_7559,N_3370,N_5144);
or U7560 (N_7560,N_5573,N_3547);
xnor U7561 (N_7561,N_5714,N_3107);
nor U7562 (N_7562,N_5974,N_5089);
or U7563 (N_7563,N_694,N_3821);
nand U7564 (N_7564,N_5282,N_1696);
nand U7565 (N_7565,N_1493,N_2062);
or U7566 (N_7566,N_565,N_3942);
xnor U7567 (N_7567,N_1479,N_4269);
nor U7568 (N_7568,N_6172,N_5062);
and U7569 (N_7569,N_1368,N_4681);
nand U7570 (N_7570,N_1969,N_2335);
or U7571 (N_7571,N_3516,N_498);
xnor U7572 (N_7572,N_4977,N_4949);
and U7573 (N_7573,N_2411,N_4055);
nand U7574 (N_7574,N_4565,N_1162);
xnor U7575 (N_7575,N_2351,N_1600);
nand U7576 (N_7576,N_4819,N_6198);
xor U7577 (N_7577,N_2728,N_3116);
or U7578 (N_7578,N_1344,N_3990);
xnor U7579 (N_7579,N_3058,N_506);
nand U7580 (N_7580,N_4526,N_5470);
xnor U7581 (N_7581,N_2680,N_2326);
nor U7582 (N_7582,N_3664,N_4245);
nor U7583 (N_7583,N_3115,N_1960);
nor U7584 (N_7584,N_2966,N_2812);
xnor U7585 (N_7585,N_5774,N_4258);
or U7586 (N_7586,N_6073,N_4189);
nand U7587 (N_7587,N_5493,N_2067);
nor U7588 (N_7588,N_5080,N_397);
xnor U7589 (N_7589,N_5988,N_2730);
xnor U7590 (N_7590,N_334,N_672);
or U7591 (N_7591,N_4783,N_6235);
or U7592 (N_7592,N_225,N_4663);
and U7593 (N_7593,N_3288,N_3524);
and U7594 (N_7594,N_5474,N_3928);
and U7595 (N_7595,N_2675,N_3224);
or U7596 (N_7596,N_2910,N_2899);
and U7597 (N_7597,N_4000,N_1290);
nand U7598 (N_7598,N_4161,N_4073);
or U7599 (N_7599,N_4594,N_3795);
xor U7600 (N_7600,N_5798,N_5417);
or U7601 (N_7601,N_2011,N_21);
xnor U7602 (N_7602,N_3096,N_3094);
and U7603 (N_7603,N_4235,N_60);
nor U7604 (N_7604,N_2379,N_1487);
nor U7605 (N_7605,N_554,N_5410);
nor U7606 (N_7606,N_192,N_595);
nand U7607 (N_7607,N_3673,N_5054);
nand U7608 (N_7608,N_5686,N_3462);
xnor U7609 (N_7609,N_5734,N_1705);
or U7610 (N_7610,N_5839,N_5568);
nor U7611 (N_7611,N_3833,N_401);
or U7612 (N_7612,N_475,N_4719);
xnor U7613 (N_7613,N_6236,N_716);
and U7614 (N_7614,N_3313,N_6113);
nor U7615 (N_7615,N_3228,N_1737);
or U7616 (N_7616,N_6243,N_1321);
nand U7617 (N_7617,N_201,N_4699);
nand U7618 (N_7618,N_3446,N_762);
nand U7619 (N_7619,N_4353,N_313);
nand U7620 (N_7620,N_5109,N_2665);
or U7621 (N_7621,N_6044,N_2688);
nor U7622 (N_7622,N_2802,N_3747);
nor U7623 (N_7623,N_6089,N_1041);
xor U7624 (N_7624,N_1964,N_2143);
nor U7625 (N_7625,N_4150,N_4355);
or U7626 (N_7626,N_4082,N_3114);
xnor U7627 (N_7627,N_2393,N_2997);
xnor U7628 (N_7628,N_2752,N_2554);
and U7629 (N_7629,N_1224,N_5243);
and U7630 (N_7630,N_821,N_1963);
nand U7631 (N_7631,N_3802,N_2507);
xnor U7632 (N_7632,N_949,N_309);
xor U7633 (N_7633,N_6008,N_4824);
nor U7634 (N_7634,N_1720,N_4534);
nor U7635 (N_7635,N_508,N_5900);
or U7636 (N_7636,N_5953,N_5929);
nor U7637 (N_7637,N_774,N_2193);
or U7638 (N_7638,N_4148,N_594);
xnor U7639 (N_7639,N_2691,N_1328);
xnor U7640 (N_7640,N_100,N_5832);
nand U7641 (N_7641,N_5817,N_2888);
xor U7642 (N_7642,N_6048,N_2583);
or U7643 (N_7643,N_5427,N_3871);
nor U7644 (N_7644,N_1971,N_772);
nor U7645 (N_7645,N_1201,N_184);
and U7646 (N_7646,N_4034,N_884);
nor U7647 (N_7647,N_3123,N_3954);
nor U7648 (N_7648,N_1728,N_1156);
or U7649 (N_7649,N_5396,N_463);
nand U7650 (N_7650,N_3270,N_3241);
and U7651 (N_7651,N_1046,N_353);
xor U7652 (N_7652,N_2401,N_1006);
nor U7653 (N_7653,N_6077,N_6082);
xnor U7654 (N_7654,N_399,N_5456);
or U7655 (N_7655,N_1738,N_3320);
xnor U7656 (N_7656,N_4480,N_4733);
or U7657 (N_7657,N_517,N_5489);
or U7658 (N_7658,N_2266,N_3021);
xnor U7659 (N_7659,N_813,N_3012);
xnor U7660 (N_7660,N_4878,N_3788);
nand U7661 (N_7661,N_2781,N_3725);
nor U7662 (N_7662,N_1800,N_30);
xor U7663 (N_7663,N_3480,N_5994);
or U7664 (N_7664,N_2765,N_4818);
nand U7665 (N_7665,N_4336,N_855);
or U7666 (N_7666,N_3160,N_2647);
nand U7667 (N_7667,N_1736,N_787);
nor U7668 (N_7668,N_3205,N_1697);
nand U7669 (N_7669,N_5279,N_5423);
nor U7670 (N_7670,N_2929,N_2218);
xnor U7671 (N_7671,N_467,N_5063);
or U7672 (N_7672,N_2532,N_388);
nand U7673 (N_7673,N_4180,N_2240);
and U7674 (N_7674,N_2023,N_1925);
and U7675 (N_7675,N_2475,N_3841);
xnor U7676 (N_7676,N_2612,N_2607);
nand U7677 (N_7677,N_5973,N_3744);
or U7678 (N_7678,N_3697,N_3312);
nand U7679 (N_7679,N_2473,N_737);
or U7680 (N_7680,N_3473,N_2824);
xnor U7681 (N_7681,N_2544,N_5258);
nor U7682 (N_7682,N_5835,N_4841);
or U7683 (N_7683,N_5886,N_5271);
nor U7684 (N_7684,N_4032,N_2533);
or U7685 (N_7685,N_2538,N_3726);
or U7686 (N_7686,N_3230,N_1434);
nor U7687 (N_7687,N_2618,N_5667);
or U7688 (N_7688,N_1373,N_798);
xor U7689 (N_7689,N_2385,N_1166);
nand U7690 (N_7690,N_2444,N_5821);
or U7691 (N_7691,N_3865,N_1981);
nor U7692 (N_7692,N_2436,N_5654);
or U7693 (N_7693,N_2580,N_1990);
and U7694 (N_7694,N_2977,N_5237);
and U7695 (N_7695,N_3968,N_4250);
and U7696 (N_7696,N_4821,N_1205);
nor U7697 (N_7697,N_3056,N_3427);
or U7698 (N_7698,N_4190,N_5590);
nand U7699 (N_7699,N_1603,N_3657);
nand U7700 (N_7700,N_4487,N_2318);
xnor U7701 (N_7701,N_4920,N_3054);
xnor U7702 (N_7702,N_2368,N_1663);
nand U7703 (N_7703,N_5428,N_1021);
or U7704 (N_7704,N_2984,N_2892);
xnor U7705 (N_7705,N_5729,N_5292);
xnor U7706 (N_7706,N_6081,N_2716);
and U7707 (N_7707,N_3559,N_64);
nand U7708 (N_7708,N_756,N_2299);
nor U7709 (N_7709,N_5166,N_3407);
nor U7710 (N_7710,N_3239,N_3851);
and U7711 (N_7711,N_4442,N_5541);
and U7712 (N_7712,N_2496,N_1441);
nand U7713 (N_7713,N_887,N_183);
and U7714 (N_7714,N_3138,N_2923);
nor U7715 (N_7715,N_4065,N_2564);
nand U7716 (N_7716,N_3195,N_4714);
nand U7717 (N_7717,N_5046,N_1831);
nand U7718 (N_7718,N_3738,N_1745);
and U7719 (N_7719,N_993,N_1633);
nor U7720 (N_7720,N_2867,N_5115);
or U7721 (N_7721,N_4956,N_5336);
and U7722 (N_7722,N_4696,N_4806);
or U7723 (N_7723,N_6009,N_3691);
and U7724 (N_7724,N_5996,N_6239);
and U7725 (N_7725,N_3997,N_4607);
nand U7726 (N_7726,N_4619,N_2975);
xnor U7727 (N_7727,N_3639,N_5284);
xor U7728 (N_7728,N_5162,N_1082);
and U7729 (N_7729,N_2378,N_693);
and U7730 (N_7730,N_3743,N_2846);
xnor U7731 (N_7731,N_5750,N_3105);
xnor U7732 (N_7732,N_875,N_4137);
xor U7733 (N_7733,N_1681,N_6108);
nand U7734 (N_7734,N_1687,N_3879);
nor U7735 (N_7735,N_1703,N_5684);
xor U7736 (N_7736,N_5884,N_522);
and U7737 (N_7737,N_4455,N_763);
and U7738 (N_7738,N_3050,N_2336);
nand U7739 (N_7739,N_3318,N_5782);
xor U7740 (N_7740,N_116,N_4485);
nor U7741 (N_7741,N_1325,N_3430);
or U7742 (N_7742,N_2732,N_3533);
nor U7743 (N_7743,N_215,N_4662);
and U7744 (N_7744,N_2518,N_3340);
nand U7745 (N_7745,N_3129,N_5270);
nor U7746 (N_7746,N_4374,N_4730);
nand U7747 (N_7747,N_3703,N_1086);
and U7748 (N_7748,N_1739,N_4060);
or U7749 (N_7749,N_4100,N_289);
or U7750 (N_7750,N_1675,N_4301);
and U7751 (N_7751,N_5912,N_110);
xnor U7752 (N_7752,N_5495,N_1695);
nand U7753 (N_7753,N_4902,N_1372);
nor U7754 (N_7754,N_1256,N_6146);
and U7755 (N_7755,N_2868,N_2325);
nand U7756 (N_7756,N_3512,N_6147);
xnor U7757 (N_7757,N_2017,N_3434);
nor U7758 (N_7758,N_4801,N_562);
and U7759 (N_7759,N_3842,N_2407);
or U7760 (N_7760,N_72,N_1560);
nand U7761 (N_7761,N_2316,N_5748);
nand U7762 (N_7762,N_6049,N_2684);
xnor U7763 (N_7763,N_3106,N_2519);
nor U7764 (N_7764,N_1500,N_1741);
or U7765 (N_7765,N_124,N_348);
xnor U7766 (N_7766,N_1206,N_3338);
xor U7767 (N_7767,N_4757,N_536);
nor U7768 (N_7768,N_1277,N_8);
nor U7769 (N_7769,N_4218,N_5070);
and U7770 (N_7770,N_1694,N_2466);
and U7771 (N_7771,N_4833,N_346);
nor U7772 (N_7772,N_1418,N_3010);
or U7773 (N_7773,N_1702,N_2049);
nand U7774 (N_7774,N_1374,N_2168);
xnor U7775 (N_7775,N_3001,N_5603);
xor U7776 (N_7776,N_3378,N_2953);
and U7777 (N_7777,N_2574,N_6019);
xnor U7778 (N_7778,N_5460,N_3776);
xnor U7779 (N_7779,N_5055,N_5169);
or U7780 (N_7780,N_6182,N_4815);
nor U7781 (N_7781,N_4443,N_2363);
or U7782 (N_7782,N_5024,N_3662);
and U7783 (N_7783,N_3843,N_1178);
nand U7784 (N_7784,N_2603,N_660);
nand U7785 (N_7785,N_3918,N_4209);
nor U7786 (N_7786,N_2211,N_1097);
nand U7787 (N_7787,N_3037,N_783);
xor U7788 (N_7788,N_1909,N_4861);
xnor U7789 (N_7789,N_4393,N_553);
nor U7790 (N_7790,N_743,N_3855);
and U7791 (N_7791,N_5822,N_3782);
and U7792 (N_7792,N_4751,N_1148);
and U7793 (N_7793,N_4854,N_3450);
xnor U7794 (N_7794,N_6175,N_3825);
nor U7795 (N_7795,N_1475,N_3771);
xnor U7796 (N_7796,N_1392,N_6140);
xnor U7797 (N_7797,N_2857,N_2066);
and U7798 (N_7798,N_2951,N_911);
xor U7799 (N_7799,N_909,N_5253);
xor U7800 (N_7800,N_3979,N_5959);
or U7801 (N_7801,N_4596,N_5921);
or U7802 (N_7802,N_4017,N_1036);
and U7803 (N_7803,N_2769,N_2397);
and U7804 (N_7804,N_4577,N_2139);
xor U7805 (N_7805,N_713,N_3092);
xnor U7806 (N_7806,N_3339,N_1149);
and U7807 (N_7807,N_4735,N_4618);
nand U7808 (N_7808,N_241,N_1975);
nand U7809 (N_7809,N_329,N_3314);
xnor U7810 (N_7810,N_2885,N_2434);
xnor U7811 (N_7811,N_2658,N_5971);
xor U7812 (N_7812,N_2296,N_1948);
or U7813 (N_7813,N_1057,N_3588);
or U7814 (N_7814,N_2927,N_5226);
and U7815 (N_7815,N_6234,N_1432);
and U7816 (N_7816,N_1569,N_382);
nor U7817 (N_7817,N_3790,N_4006);
nand U7818 (N_7818,N_4281,N_1001);
nand U7819 (N_7819,N_4778,N_5415);
nor U7820 (N_7820,N_3135,N_2660);
and U7821 (N_7821,N_1226,N_50);
or U7822 (N_7822,N_5342,N_495);
or U7823 (N_7823,N_5612,N_6024);
nand U7824 (N_7824,N_4339,N_6197);
xnor U7825 (N_7825,N_2535,N_1242);
nor U7826 (N_7826,N_933,N_542);
xor U7827 (N_7827,N_3769,N_4037);
and U7828 (N_7828,N_630,N_3444);
nor U7829 (N_7829,N_5339,N_2395);
xor U7830 (N_7830,N_2698,N_5904);
nor U7831 (N_7831,N_1454,N_2595);
and U7832 (N_7832,N_1578,N_2839);
and U7833 (N_7833,N_2448,N_5743);
nand U7834 (N_7834,N_5426,N_1783);
and U7835 (N_7835,N_2057,N_2422);
xnor U7836 (N_7836,N_5880,N_3838);
and U7837 (N_7837,N_782,N_1136);
and U7838 (N_7838,N_188,N_1701);
nor U7839 (N_7839,N_4657,N_890);
xor U7840 (N_7840,N_6064,N_5808);
xor U7841 (N_7841,N_2085,N_3986);
xnor U7842 (N_7842,N_5207,N_2377);
nor U7843 (N_7843,N_3504,N_1358);
or U7844 (N_7844,N_605,N_3970);
xnor U7845 (N_7845,N_5069,N_563);
xnor U7846 (N_7846,N_1877,N_4402);
nand U7847 (N_7847,N_432,N_3490);
xnor U7848 (N_7848,N_4718,N_2338);
or U7849 (N_7849,N_5052,N_5706);
xor U7850 (N_7850,N_6014,N_5429);
and U7851 (N_7851,N_2301,N_78);
nand U7852 (N_7852,N_5756,N_5630);
xnor U7853 (N_7853,N_4717,N_4194);
xor U7854 (N_7854,N_1620,N_4554);
or U7855 (N_7855,N_5170,N_599);
nor U7856 (N_7856,N_5471,N_786);
nand U7857 (N_7857,N_928,N_2080);
or U7858 (N_7858,N_3728,N_4260);
or U7859 (N_7859,N_980,N_1396);
xor U7860 (N_7860,N_2596,N_2453);
nand U7861 (N_7861,N_1887,N_136);
xnor U7862 (N_7862,N_2006,N_41);
nand U7863 (N_7863,N_3485,N_868);
nand U7864 (N_7864,N_4419,N_2549);
and U7865 (N_7865,N_664,N_1843);
nand U7866 (N_7866,N_4089,N_1879);
xor U7867 (N_7867,N_796,N_2842);
nand U7868 (N_7868,N_1693,N_4124);
and U7869 (N_7869,N_2782,N_5657);
and U7870 (N_7870,N_3176,N_198);
nor U7871 (N_7871,N_3147,N_4305);
nand U7872 (N_7872,N_4874,N_3702);
nor U7873 (N_7873,N_4164,N_2135);
or U7874 (N_7874,N_279,N_684);
nand U7875 (N_7875,N_5920,N_668);
nand U7876 (N_7876,N_709,N_1715);
nand U7877 (N_7877,N_5414,N_4816);
nand U7878 (N_7878,N_1362,N_4793);
xnor U7879 (N_7879,N_4449,N_5468);
or U7880 (N_7880,N_4337,N_3685);
nor U7881 (N_7881,N_6161,N_1337);
nor U7882 (N_7882,N_1689,N_5807);
and U7883 (N_7883,N_3540,N_4199);
or U7884 (N_7884,N_3393,N_3699);
nand U7885 (N_7885,N_1179,N_3424);
nor U7886 (N_7886,N_2503,N_6129);
nand U7887 (N_7887,N_590,N_4645);
nand U7888 (N_7888,N_1812,N_5967);
and U7889 (N_7889,N_3658,N_2586);
nand U7890 (N_7890,N_824,N_3440);
xor U7891 (N_7891,N_4968,N_3870);
xnor U7892 (N_7892,N_3650,N_538);
and U7893 (N_7893,N_4334,N_4308);
or U7894 (N_7894,N_1059,N_1376);
or U7895 (N_7895,N_4361,N_537);
xnor U7896 (N_7896,N_5628,N_4304);
nand U7897 (N_7897,N_6240,N_1647);
and U7898 (N_7898,N_3701,N_5837);
nor U7899 (N_7899,N_639,N_1883);
nand U7900 (N_7900,N_178,N_5240);
xnor U7901 (N_7901,N_5442,N_372);
or U7902 (N_7902,N_61,N_2747);
or U7903 (N_7903,N_6224,N_6191);
nand U7904 (N_7904,N_4410,N_1407);
xor U7905 (N_7905,N_5367,N_1260);
nand U7906 (N_7906,N_3502,N_1081);
nand U7907 (N_7907,N_1207,N_4890);
xnor U7908 (N_7908,N_2743,N_3758);
nand U7909 (N_7909,N_3433,N_3274);
nand U7910 (N_7910,N_3797,N_739);
nand U7911 (N_7911,N_5099,N_1958);
nor U7912 (N_7912,N_2455,N_13);
nand U7913 (N_7913,N_2291,N_571);
xor U7914 (N_7914,N_5328,N_5854);
nor U7915 (N_7915,N_3902,N_4516);
xnor U7916 (N_7916,N_4085,N_3007);
and U7917 (N_7917,N_810,N_962);
and U7918 (N_7918,N_2184,N_4185);
or U7919 (N_7919,N_983,N_6);
and U7920 (N_7920,N_5639,N_1116);
nand U7921 (N_7921,N_2129,N_5473);
nor U7922 (N_7922,N_1511,N_189);
or U7923 (N_7923,N_3676,N_4244);
or U7924 (N_7924,N_2699,N_237);
nor U7925 (N_7925,N_1516,N_820);
nand U7926 (N_7926,N_1970,N_666);
nand U7927 (N_7927,N_897,N_3348);
xnor U7928 (N_7928,N_1122,N_2971);
and U7929 (N_7929,N_4654,N_5512);
nor U7930 (N_7930,N_3240,N_2522);
and U7931 (N_7931,N_3720,N_3071);
or U7932 (N_7932,N_4771,N_2265);
and U7933 (N_7933,N_4098,N_1886);
or U7934 (N_7934,N_2686,N_996);
nor U7935 (N_7935,N_4471,N_297);
nor U7936 (N_7936,N_2150,N_3736);
and U7937 (N_7937,N_3311,N_4483);
xor U7938 (N_7938,N_4561,N_4147);
nand U7939 (N_7939,N_3938,N_3429);
xor U7940 (N_7940,N_1996,N_5204);
xor U7941 (N_7941,N_3864,N_5537);
nor U7942 (N_7942,N_283,N_5677);
and U7943 (N_7943,N_5852,N_4475);
and U7944 (N_7944,N_4505,N_5326);
xor U7945 (N_7945,N_5058,N_437);
nor U7946 (N_7946,N_5801,N_5872);
xor U7947 (N_7947,N_5223,N_3817);
or U7948 (N_7948,N_4314,N_2431);
or U7949 (N_7949,N_3613,N_3679);
and U7950 (N_7950,N_2687,N_363);
and U7951 (N_7951,N_3557,N_2731);
nand U7952 (N_7952,N_1395,N_5548);
or U7953 (N_7953,N_2212,N_2693);
or U7954 (N_7954,N_3289,N_865);
or U7955 (N_7955,N_3035,N_1707);
nand U7956 (N_7956,N_5016,N_4441);
nor U7957 (N_7957,N_6013,N_1523);
nor U7958 (N_7958,N_1169,N_331);
and U7959 (N_7959,N_2098,N_523);
or U7960 (N_7960,N_5435,N_1154);
nor U7961 (N_7961,N_2950,N_4777);
or U7962 (N_7962,N_322,N_6084);
nand U7963 (N_7963,N_2421,N_3425);
xnor U7964 (N_7964,N_4045,N_2078);
xnor U7965 (N_7965,N_2381,N_3278);
nand U7966 (N_7966,N_5317,N_1616);
and U7967 (N_7967,N_6050,N_5692);
and U7968 (N_7968,N_106,N_1807);
xor U7969 (N_7969,N_4387,N_375);
nor U7970 (N_7970,N_123,N_3511);
or U7971 (N_7971,N_234,N_1893);
nand U7972 (N_7972,N_3353,N_6053);
nand U7973 (N_7973,N_255,N_2671);
nor U7974 (N_7974,N_5875,N_5652);
xor U7975 (N_7975,N_593,N_4335);
nor U7976 (N_7976,N_252,N_3281);
nand U7977 (N_7977,N_5401,N_5437);
nor U7978 (N_7978,N_5861,N_1661);
xor U7979 (N_7979,N_2869,N_4271);
and U7980 (N_7980,N_861,N_5549);
nor U7981 (N_7981,N_5028,N_115);
nor U7982 (N_7982,N_5095,N_1131);
and U7983 (N_7983,N_2941,N_1216);
nand U7984 (N_7984,N_4450,N_3644);
nor U7985 (N_7985,N_1587,N_4924);
or U7986 (N_7986,N_3789,N_4473);
xor U7987 (N_7987,N_4373,N_3305);
nand U7988 (N_7988,N_2200,N_3891);
and U7989 (N_7989,N_4923,N_4042);
or U7990 (N_7990,N_1377,N_6059);
nor U7991 (N_7991,N_1901,N_4720);
nor U7992 (N_7992,N_260,N_1199);
and U7993 (N_7993,N_300,N_6005);
nor U7994 (N_7994,N_4790,N_3169);
xnor U7995 (N_7995,N_3696,N_3893);
nand U7996 (N_7996,N_3876,N_4624);
and U7997 (N_7997,N_2625,N_4187);
xor U7998 (N_7998,N_4035,N_2556);
and U7999 (N_7999,N_1921,N_4590);
nand U8000 (N_8000,N_4351,N_5626);
xor U8001 (N_8001,N_1764,N_3660);
nor U8002 (N_8002,N_3910,N_2537);
nand U8003 (N_8003,N_44,N_4362);
and U8004 (N_8004,N_2944,N_1339);
nor U8005 (N_8005,N_6000,N_1900);
xnor U8006 (N_8006,N_3243,N_5061);
nand U8007 (N_8007,N_3303,N_4103);
nor U8008 (N_8008,N_925,N_3291);
nor U8009 (N_8009,N_3093,N_4850);
and U8010 (N_8010,N_4785,N_3165);
xnor U8011 (N_8011,N_5809,N_228);
and U8012 (N_8012,N_1913,N_2928);
or U8013 (N_8013,N_5847,N_1444);
nand U8014 (N_8014,N_5355,N_3016);
or U8015 (N_8015,N_6040,N_1037);
and U8016 (N_8016,N_4268,N_1100);
or U8017 (N_8017,N_1013,N_1113);
or U8018 (N_8018,N_5043,N_1773);
xor U8019 (N_8019,N_6202,N_5247);
nand U8020 (N_8020,N_5746,N_1276);
xnor U8021 (N_8021,N_4295,N_1264);
and U8022 (N_8022,N_3075,N_3023);
nor U8023 (N_8023,N_2142,N_714);
nor U8024 (N_8024,N_1164,N_589);
nor U8025 (N_8025,N_3164,N_502);
and U8026 (N_8026,N_4866,N_3384);
xnor U8027 (N_8027,N_5806,N_5754);
and U8028 (N_8028,N_661,N_3319);
nand U8029 (N_8029,N_1548,N_3847);
xnor U8030 (N_8030,N_5923,N_846);
and U8031 (N_8031,N_520,N_1622);
and U8032 (N_8032,N_5190,N_2994);
and U8033 (N_8033,N_2636,N_1049);
nor U8034 (N_8034,N_5314,N_459);
nor U8035 (N_8035,N_5764,N_4811);
nand U8036 (N_8036,N_3148,N_4153);
nor U8037 (N_8037,N_4003,N_3213);
xnor U8038 (N_8038,N_1734,N_1066);
nor U8039 (N_8039,N_2849,N_271);
and U8040 (N_8040,N_439,N_476);
or U8041 (N_8041,N_3265,N_3904);
nor U8042 (N_8042,N_3710,N_3591);
and U8043 (N_8043,N_166,N_1094);
and U8044 (N_8044,N_1159,N_2261);
or U8045 (N_8045,N_2342,N_4695);
nand U8046 (N_8046,N_5598,N_5354);
or U8047 (N_8047,N_728,N_101);
xor U8048 (N_8048,N_312,N_5826);
xor U8049 (N_8049,N_1564,N_5106);
nor U8050 (N_8050,N_5466,N_2963);
nand U8051 (N_8051,N_5768,N_3671);
nand U8052 (N_8052,N_3564,N_3525);
nand U8053 (N_8053,N_2408,N_1992);
nand U8054 (N_8054,N_4238,N_2529);
nand U8055 (N_8055,N_90,N_6056);
and U8056 (N_8056,N_4413,N_1304);
xnor U8057 (N_8057,N_4637,N_4725);
nand U8058 (N_8058,N_3282,N_4174);
and U8059 (N_8059,N_5554,N_4290);
xnor U8060 (N_8060,N_4421,N_609);
or U8061 (N_8061,N_1229,N_1212);
nand U8062 (N_8062,N_3582,N_3651);
nand U8063 (N_8063,N_1363,N_45);
and U8064 (N_8064,N_3179,N_736);
nor U8065 (N_8065,N_5772,N_3623);
and U8066 (N_8066,N_3043,N_5236);
or U8067 (N_8067,N_3162,N_5732);
nand U8068 (N_8068,N_6222,N_4435);
nor U8069 (N_8069,N_2653,N_4300);
or U8070 (N_8070,N_134,N_641);
nor U8071 (N_8071,N_5122,N_6116);
and U8072 (N_8072,N_2259,N_4062);
or U8073 (N_8073,N_2905,N_4332);
and U8074 (N_8074,N_5217,N_2117);
nor U8075 (N_8075,N_1632,N_790);
nand U8076 (N_8076,N_298,N_1167);
xnor U8077 (N_8077,N_5312,N_3300);
or U8078 (N_8078,N_3436,N_4879);
nor U8079 (N_8079,N_5025,N_3130);
xnor U8080 (N_8080,N_3972,N_3139);
nor U8081 (N_8081,N_830,N_780);
xnor U8082 (N_8082,N_2256,N_5450);
xnor U8083 (N_8083,N_5346,N_3222);
xnor U8084 (N_8084,N_4122,N_2304);
and U8085 (N_8085,N_2520,N_2872);
nand U8086 (N_8086,N_1791,N_3152);
nand U8087 (N_8087,N_2278,N_2620);
nor U8088 (N_8088,N_4653,N_3385);
nor U8089 (N_8089,N_860,N_5164);
xor U8090 (N_8090,N_1125,N_1565);
nand U8091 (N_8091,N_3132,N_3624);
xor U8092 (N_8092,N_58,N_2047);
nor U8093 (N_8093,N_5318,N_4200);
xor U8094 (N_8094,N_2509,N_5065);
nor U8095 (N_8095,N_4110,N_4675);
or U8096 (N_8096,N_4744,N_3090);
nor U8097 (N_8097,N_5451,N_6007);
xnor U8098 (N_8098,N_5645,N_1448);
nand U8099 (N_8099,N_469,N_1294);
and U8100 (N_8100,N_5219,N_1690);
and U8101 (N_8101,N_4459,N_3048);
and U8102 (N_8102,N_3344,N_2664);
and U8103 (N_8103,N_1536,N_2409);
nor U8104 (N_8104,N_5459,N_111);
nand U8105 (N_8105,N_1364,N_2292);
or U8106 (N_8106,N_907,N_4919);
or U8107 (N_8107,N_6216,N_4064);
nor U8108 (N_8108,N_6046,N_4024);
xnor U8109 (N_8109,N_4542,N_5037);
nor U8110 (N_8110,N_5297,N_969);
xnor U8111 (N_8111,N_5273,N_1072);
nand U8112 (N_8112,N_5212,N_1172);
nand U8113 (N_8113,N_4640,N_4418);
or U8114 (N_8114,N_2800,N_6232);
or U8115 (N_8115,N_3359,N_4555);
or U8116 (N_8116,N_5118,N_3267);
nand U8117 (N_8117,N_2344,N_2074);
or U8118 (N_8118,N_3975,N_5943);
and U8119 (N_8119,N_263,N_5224);
xnor U8120 (N_8120,N_4764,N_644);
or U8121 (N_8121,N_2530,N_1239);
nor U8122 (N_8122,N_2040,N_3718);
nand U8123 (N_8123,N_647,N_1220);
nor U8124 (N_8124,N_829,N_6004);
xor U8125 (N_8125,N_4731,N_3263);
nor U8126 (N_8126,N_4638,N_3122);
and U8127 (N_8127,N_5179,N_4585);
nor U8128 (N_8128,N_5215,N_1471);
or U8129 (N_8129,N_4175,N_2307);
and U8130 (N_8130,N_1078,N_4145);
and U8131 (N_8131,N_5494,N_678);
or U8132 (N_8132,N_4104,N_3976);
or U8133 (N_8133,N_1634,N_2357);
nor U8134 (N_8134,N_3880,N_6047);
xor U8135 (N_8135,N_1830,N_1494);
nor U8136 (N_8136,N_4094,N_4462);
nand U8137 (N_8137,N_5633,N_2933);
and U8138 (N_8138,N_4477,N_3453);
or U8139 (N_8139,N_2446,N_98);
nand U8140 (N_8140,N_877,N_5379);
or U8141 (N_8141,N_637,N_3500);
or U8142 (N_8142,N_2985,N_1279);
xor U8143 (N_8143,N_6132,N_1288);
nand U8144 (N_8144,N_1575,N_2456);
xnor U8145 (N_8145,N_734,N_688);
and U8146 (N_8146,N_5439,N_3555);
nand U8147 (N_8147,N_3084,N_3579);
nand U8148 (N_8148,N_427,N_2561);
and U8149 (N_8149,N_1175,N_2890);
and U8150 (N_8150,N_4639,N_2980);
xor U8151 (N_8151,N_1576,N_407);
xnor U8152 (N_8152,N_5205,N_4054);
xnor U8153 (N_8153,N_2099,N_2451);
xnor U8154 (N_8154,N_2223,N_3967);
nand U8155 (N_8155,N_1532,N_5785);
nor U8156 (N_8156,N_4875,N_3507);
nor U8157 (N_8157,N_769,N_2037);
and U8158 (N_8158,N_3468,N_2214);
nor U8159 (N_8159,N_2777,N_4397);
and U8160 (N_8160,N_4669,N_5067);
or U8161 (N_8161,N_1385,N_3653);
nand U8162 (N_8162,N_1040,N_541);
nor U8163 (N_8163,N_4649,N_826);
or U8164 (N_8164,N_532,N_3024);
nand U8165 (N_8165,N_319,N_5771);
nand U8166 (N_8166,N_34,N_1698);
and U8167 (N_8167,N_193,N_135);
or U8168 (N_8168,N_1353,N_6099);
nand U8169 (N_8169,N_5484,N_6043);
xnor U8170 (N_8170,N_5858,N_1322);
or U8171 (N_8171,N_4623,N_5653);
xor U8172 (N_8172,N_741,N_4870);
xnor U8173 (N_8173,N_4687,N_1103);
or U8174 (N_8174,N_3121,N_4088);
and U8175 (N_8175,N_2470,N_4229);
xor U8176 (N_8176,N_1501,N_3206);
nand U8177 (N_8177,N_6242,N_1757);
or U8178 (N_8178,N_1020,N_4965);
or U8179 (N_8179,N_4213,N_5672);
nand U8180 (N_8180,N_1874,N_3635);
or U8181 (N_8181,N_665,N_5763);
nor U8182 (N_8182,N_818,N_2633);
or U8183 (N_8183,N_2138,N_1063);
nand U8184 (N_8184,N_1983,N_3774);
xor U8185 (N_8185,N_3719,N_4840);
or U8186 (N_8186,N_5307,N_450);
xnor U8187 (N_8187,N_5605,N_4080);
nand U8188 (N_8188,N_5436,N_2804);
nor U8189 (N_8189,N_5222,N_4468);
nor U8190 (N_8190,N_5108,N_224);
nor U8191 (N_8191,N_4876,N_2882);
nand U8192 (N_8192,N_33,N_702);
and U8193 (N_8193,N_3705,N_3060);
and U8194 (N_8194,N_2160,N_5870);
and U8195 (N_8195,N_2920,N_282);
and U8196 (N_8196,N_1470,N_1821);
or U8197 (N_8197,N_2738,N_1664);
xor U8198 (N_8198,N_4232,N_718);
nor U8199 (N_8199,N_4595,N_3190);
nor U8200 (N_8200,N_4667,N_6230);
nor U8201 (N_8201,N_3767,N_744);
or U8202 (N_8202,N_6190,N_4092);
and U8203 (N_8203,N_1123,N_1126);
and U8204 (N_8204,N_1735,N_1145);
and U8205 (N_8205,N_1648,N_5283);
nor U8206 (N_8206,N_4917,N_1502);
xor U8207 (N_8207,N_2606,N_5527);
and U8208 (N_8208,N_4575,N_5180);
nor U8209 (N_8209,N_6148,N_2772);
nand U8210 (N_8210,N_2534,N_4905);
nand U8211 (N_8211,N_2914,N_4365);
nand U8212 (N_8212,N_4502,N_2901);
nand U8213 (N_8213,N_1468,N_5165);
and U8214 (N_8214,N_489,N_5285);
nor U8215 (N_8215,N_2594,N_952);
nand U8216 (N_8216,N_5187,N_2826);
or U8217 (N_8217,N_5444,N_4331);
and U8218 (N_8218,N_3315,N_5783);
and U8219 (N_8219,N_6195,N_1297);
nor U8220 (N_8220,N_3374,N_2018);
and U8221 (N_8221,N_3402,N_1621);
and U8222 (N_8222,N_4521,N_5320);
and U8223 (N_8223,N_6227,N_5137);
or U8224 (N_8224,N_805,N_5565);
xnor U8225 (N_8225,N_1529,N_833);
nor U8226 (N_8226,N_4340,N_11);
nand U8227 (N_8227,N_1257,N_2442);
nor U8228 (N_8228,N_4015,N_504);
xnor U8229 (N_8229,N_356,N_6115);
and U8230 (N_8230,N_4573,N_4415);
nand U8231 (N_8231,N_5805,N_2181);
or U8232 (N_8232,N_6156,N_4934);
or U8233 (N_8233,N_4484,N_4865);
nand U8234 (N_8234,N_673,N_632);
or U8235 (N_8235,N_3172,N_3496);
and U8236 (N_8236,N_4617,N_3275);
xor U8237 (N_8237,N_1230,N_4847);
and U8238 (N_8238,N_3920,N_663);
and U8239 (N_8239,N_1784,N_5742);
and U8240 (N_8240,N_5488,N_4974);
nand U8241 (N_8241,N_2206,N_2283);
xnor U8242 (N_8242,N_978,N_3745);
or U8243 (N_8243,N_871,N_1147);
nand U8244 (N_8244,N_108,N_557);
xnor U8245 (N_8245,N_5856,N_5781);
xnor U8246 (N_8246,N_3069,N_2092);
nor U8247 (N_8247,N_5891,N_2104);
and U8248 (N_8248,N_3672,N_4491);
xnor U8249 (N_8249,N_2762,N_1301);
and U8250 (N_8250,N_1904,N_5081);
nor U8251 (N_8251,N_2091,N_3403);
and U8252 (N_8252,N_1650,N_5589);
nor U8253 (N_8253,N_4149,N_1727);
nand U8254 (N_8254,N_3208,N_3982);
nand U8255 (N_8255,N_5349,N_3236);
or U8256 (N_8256,N_3479,N_5788);
nor U8257 (N_8257,N_4057,N_3688);
or U8258 (N_8258,N_5691,N_3666);
nor U8259 (N_8259,N_5345,N_4013);
xor U8260 (N_8260,N_863,N_5071);
xnor U8261 (N_8261,N_5033,N_1270);
or U8262 (N_8262,N_4704,N_3191);
nor U8263 (N_8263,N_2742,N_3532);
and U8264 (N_8264,N_1572,N_455);
and U8265 (N_8265,N_1371,N_4948);
and U8266 (N_8266,N_2807,N_3836);
nor U8267 (N_8267,N_1554,N_748);
or U8268 (N_8268,N_2566,N_107);
nor U8269 (N_8269,N_2592,N_5700);
and U8270 (N_8270,N_5337,N_755);
or U8271 (N_8271,N_4544,N_2365);
nand U8272 (N_8272,N_2294,N_1759);
and U8273 (N_8273,N_1379,N_125);
nand U8274 (N_8274,N_892,N_5787);
or U8275 (N_8275,N_2604,N_2087);
or U8276 (N_8276,N_5869,N_3599);
and U8277 (N_8277,N_2167,N_5465);
nor U8278 (N_8278,N_1008,N_3521);
or U8279 (N_8279,N_1168,N_3399);
nor U8280 (N_8280,N_1292,N_4603);
xnor U8281 (N_8281,N_5481,N_3292);
nand U8282 (N_8282,N_3018,N_5303);
nand U8283 (N_8283,N_831,N_2790);
nand U8284 (N_8284,N_908,N_2557);
nor U8285 (N_8285,N_997,N_6110);
nor U8286 (N_8286,N_199,N_5082);
nand U8287 (N_8287,N_1865,N_288);
nor U8288 (N_8288,N_1056,N_5623);
or U8289 (N_8289,N_5272,N_2493);
nor U8290 (N_8290,N_5925,N_5301);
nor U8291 (N_8291,N_1079,N_335);
nand U8292 (N_8292,N_3441,N_3835);
or U8293 (N_8293,N_5649,N_296);
or U8294 (N_8294,N_3518,N_5979);
and U8295 (N_8295,N_2204,N_2898);
nor U8296 (N_8296,N_6165,N_3822);
nand U8297 (N_8297,N_3752,N_2880);
and U8298 (N_8298,N_3763,N_2427);
or U8299 (N_8299,N_5416,N_2517);
and U8300 (N_8300,N_302,N_4727);
nand U8301 (N_8301,N_3484,N_1492);
nand U8302 (N_8302,N_6149,N_3700);
and U8303 (N_8303,N_1858,N_2485);
nand U8304 (N_8304,N_2792,N_3064);
nand U8305 (N_8305,N_2051,N_1477);
or U8306 (N_8306,N_4490,N_5334);
nor U8307 (N_8307,N_6112,N_2154);
and U8308 (N_8308,N_1686,N_3171);
nand U8309 (N_8309,N_5849,N_2895);
or U8310 (N_8310,N_1420,N_2970);
nand U8311 (N_8311,N_2481,N_5311);
and U8312 (N_8312,N_5433,N_2736);
xnor U8313 (N_8313,N_1677,N_3816);
nand U8314 (N_8314,N_6023,N_4093);
or U8315 (N_8315,N_5644,N_3198);
and U8316 (N_8316,N_3709,N_1792);
nand U8317 (N_8317,N_5892,N_5113);
and U8318 (N_8318,N_603,N_2602);
nor U8319 (N_8319,N_1704,N_1966);
or U8320 (N_8320,N_1073,N_2708);
nor U8321 (N_8321,N_462,N_742);
nor U8322 (N_8322,N_1415,N_4789);
nor U8323 (N_8323,N_3280,N_5616);
and U8324 (N_8324,N_3245,N_4752);
nor U8325 (N_8325,N_862,N_1794);
nor U8326 (N_8326,N_3221,N_3663);
and U8327 (N_8327,N_905,N_471);
nor U8328 (N_8328,N_1839,N_3477);
nor U8329 (N_8329,N_385,N_3597);
nand U8330 (N_8330,N_3562,N_4990);
and U8331 (N_8331,N_5002,N_3576);
nand U8332 (N_8332,N_3097,N_2398);
nand U8333 (N_8333,N_3459,N_400);
nand U8334 (N_8334,N_3389,N_4807);
xnor U8335 (N_8335,N_5160,N_2965);
or U8336 (N_8336,N_4930,N_6233);
xnor U8337 (N_8337,N_5804,N_2303);
and U8338 (N_8338,N_195,N_2972);
nand U8339 (N_8339,N_1281,N_3297);
xor U8340 (N_8340,N_5368,N_6136);
and U8341 (N_8341,N_435,N_268);
or U8342 (N_8342,N_4741,N_2973);
xnor U8343 (N_8343,N_1458,N_2492);
and U8344 (N_8344,N_5874,N_3681);
or U8345 (N_8345,N_1044,N_5676);
xor U8346 (N_8346,N_2601,N_1387);
nor U8347 (N_8347,N_1048,N_789);
and U8348 (N_8348,N_4984,N_5434);
or U8349 (N_8349,N_5946,N_956);
or U8350 (N_8350,N_2205,N_1930);
and U8351 (N_8351,N_573,N_3196);
nand U8352 (N_8352,N_3125,N_1551);
nor U8353 (N_8353,N_4688,N_675);
nand U8354 (N_8354,N_3956,N_726);
or U8355 (N_8355,N_1060,N_4868);
nand U8356 (N_8356,N_5385,N_1889);
or U8357 (N_8357,N_2840,N_248);
nor U8358 (N_8358,N_1296,N_102);
and U8359 (N_8359,N_3554,N_304);
nand U8360 (N_8360,N_1649,N_1666);
and U8361 (N_8361,N_4263,N_2254);
nand U8362 (N_8362,N_4284,N_5014);
nor U8363 (N_8363,N_2500,N_381);
or U8364 (N_8364,N_5918,N_3284);
nand U8365 (N_8365,N_6075,N_430);
xor U8366 (N_8366,N_770,N_2881);
or U8367 (N_8367,N_2774,N_2861);
xor U8368 (N_8368,N_2992,N_265);
xor U8369 (N_8369,N_6186,N_4756);
xor U8370 (N_8370,N_6145,N_2319);
and U8371 (N_8371,N_971,N_3916);
nand U8372 (N_8372,N_4828,N_521);
and U8373 (N_8373,N_5963,N_5139);
nand U8374 (N_8374,N_3955,N_5235);
and U8375 (N_8375,N_754,N_959);
nor U8376 (N_8376,N_3573,N_4429);
nor U8377 (N_8377,N_2637,N_4792);
nand U8378 (N_8378,N_4039,N_2712);
and U8379 (N_8379,N_2115,N_6127);
nand U8380 (N_8380,N_2877,N_4242);
xnor U8381 (N_8381,N_5501,N_6088);
nand U8382 (N_8382,N_2293,N_3945);
nor U8383 (N_8383,N_1841,N_5580);
nor U8384 (N_8384,N_731,N_5871);
nor U8385 (N_8385,N_1588,N_122);
or U8386 (N_8386,N_1274,N_985);
and U8387 (N_8387,N_717,N_1859);
nor U8388 (N_8388,N_5910,N_3881);
or U8389 (N_8389,N_1965,N_4388);
and U8390 (N_8390,N_3259,N_1228);
xor U8391 (N_8391,N_5050,N_4121);
and U8392 (N_8392,N_3768,N_1033);
nor U8393 (N_8393,N_658,N_5293);
nand U8394 (N_8394,N_1931,N_1431);
or U8395 (N_8395,N_3337,N_4664);
or U8396 (N_8396,N_656,N_2450);
nand U8397 (N_8397,N_1726,N_3451);
or U8398 (N_8398,N_1488,N_3757);
and U8399 (N_8399,N_5079,N_3371);
or U8400 (N_8400,N_465,N_1423);
or U8401 (N_8401,N_840,N_5378);
nor U8402 (N_8402,N_3421,N_751);
or U8403 (N_8403,N_2831,N_4095);
xor U8404 (N_8404,N_5566,N_3146);
and U8405 (N_8405,N_2682,N_2689);
nor U8406 (N_8406,N_2949,N_649);
and U8407 (N_8407,N_1085,N_5185);
or U8408 (N_8408,N_3369,N_4275);
and U8409 (N_8409,N_203,N_5688);
xor U8410 (N_8410,N_293,N_4633);
nand U8411 (N_8411,N_2285,N_3803);
nand U8412 (N_8412,N_4950,N_2642);
or U8413 (N_8413,N_5199,N_1138);
nor U8414 (N_8414,N_711,N_1805);
and U8415 (N_8415,N_3832,N_1642);
xnor U8416 (N_8416,N_5049,N_5622);
xnor U8417 (N_8417,N_1267,N_4760);
xnor U8418 (N_8418,N_3722,N_825);
or U8419 (N_8419,N_2799,N_3804);
nand U8420 (N_8420,N_514,N_977);
xnor U8421 (N_8421,N_5064,N_5857);
nand U8422 (N_8422,N_2069,N_3611);
or U8423 (N_8423,N_2748,N_3232);
or U8424 (N_8424,N_281,N_4324);
and U8425 (N_8425,N_4563,N_5514);
xor U8426 (N_8426,N_1077,N_94);
xnor U8427 (N_8427,N_2871,N_6035);
nand U8428 (N_8428,N_2524,N_1557);
nor U8429 (N_8429,N_1019,N_596);
or U8430 (N_8430,N_5635,N_1121);
or U8431 (N_8431,N_3571,N_2108);
nand U8432 (N_8432,N_258,N_4985);
and U8433 (N_8433,N_3304,N_2540);
xnor U8434 (N_8434,N_4453,N_4212);
nand U8435 (N_8435,N_4707,N_1132);
or U8436 (N_8436,N_4615,N_5376);
nor U8437 (N_8437,N_6102,N_574);
and U8438 (N_8438,N_2345,N_4016);
nor U8439 (N_8439,N_5105,N_1977);
and U8440 (N_8440,N_5327,N_2744);
nor U8441 (N_8441,N_3212,N_143);
and U8442 (N_8442,N_5091,N_1641);
or U8443 (N_8443,N_923,N_4903);
or U8444 (N_8444,N_6220,N_1187);
nor U8445 (N_8445,N_3197,N_598);
nor U8446 (N_8446,N_4422,N_4863);
or U8447 (N_8447,N_392,N_3362);
and U8448 (N_8448,N_5406,N_2428);
xor U8449 (N_8449,N_3294,N_3098);
xor U8450 (N_8450,N_4456,N_4292);
and U8451 (N_8451,N_3869,N_1196);
nor U8452 (N_8452,N_1202,N_2242);
nand U8453 (N_8453,N_5999,N_3167);
xnor U8454 (N_8454,N_3764,N_71);
nor U8455 (N_8455,N_5898,N_3365);
nand U8456 (N_8456,N_1906,N_43);
or U8457 (N_8457,N_2829,N_1555);
nand U8458 (N_8458,N_3346,N_4);
and U8459 (N_8459,N_4825,N_2112);
nor U8460 (N_8460,N_2097,N_4803);
nand U8461 (N_8461,N_2153,N_5738);
or U8462 (N_8462,N_144,N_3695);
or U8463 (N_8463,N_2086,N_2737);
nand U8464 (N_8464,N_4722,N_4166);
or U8465 (N_8465,N_1485,N_387);
nand U8466 (N_8466,N_3819,N_1776);
nand U8467 (N_8467,N_1483,N_181);
nor U8468 (N_8468,N_5096,N_2468);
nor U8469 (N_8469,N_2128,N_5382);
nand U8470 (N_8470,N_2194,N_404);
xor U8471 (N_8471,N_5116,N_6122);
xor U8472 (N_8472,N_3181,N_679);
or U8473 (N_8473,N_2611,N_4306);
nand U8474 (N_8474,N_2827,N_4027);
xnor U8475 (N_8475,N_4318,N_197);
nor U8476 (N_8476,N_112,N_1840);
or U8477 (N_8477,N_6248,N_3019);
nor U8478 (N_8478,N_4231,N_3367);
nor U8479 (N_8479,N_187,N_3086);
nor U8480 (N_8480,N_5780,N_2906);
and U8481 (N_8481,N_1120,N_921);
or U8482 (N_8482,N_3372,N_4962);
xor U8483 (N_8483,N_3495,N_1785);
nor U8484 (N_8484,N_5210,N_1316);
or U8485 (N_8485,N_3716,N_1247);
xor U8486 (N_8486,N_3808,N_4051);
or U8487 (N_8487,N_5569,N_3426);
and U8488 (N_8488,N_3269,N_4820);
and U8489 (N_8489,N_2513,N_1855);
or U8490 (N_8490,N_6117,N_3674);
xnor U8491 (N_8491,N_2082,N_1583);
nand U8492 (N_8492,N_5980,N_5983);
xor U8493 (N_8493,N_3174,N_1435);
xnor U8494 (N_8494,N_3868,N_4106);
or U8495 (N_8495,N_3794,N_5567);
and U8496 (N_8496,N_5535,N_3711);
and U8497 (N_8497,N_4101,N_1573);
or U8498 (N_8498,N_671,N_1849);
nor U8499 (N_8499,N_1476,N_4479);
or U8500 (N_8500,N_3257,N_2497);
nand U8501 (N_8501,N_1869,N_5407);
xor U8502 (N_8502,N_885,N_3560);
nor U8503 (N_8503,N_1903,N_1052);
nand U8504 (N_8504,N_4465,N_2750);
xnor U8505 (N_8505,N_1370,N_4273);
nor U8506 (N_8506,N_2847,N_5543);
or U8507 (N_8507,N_6192,N_2597);
nand U8508 (N_8508,N_4009,N_1293);
and U8509 (N_8509,N_4007,N_1268);
nand U8510 (N_8510,N_3248,N_1979);
or U8511 (N_8511,N_4817,N_3454);
or U8512 (N_8512,N_4546,N_4708);
nand U8513 (N_8513,N_1181,N_2641);
nand U8514 (N_8514,N_4986,N_3052);
or U8515 (N_8515,N_4498,N_1684);
nand U8516 (N_8516,N_2025,N_1425);
and U8517 (N_8517,N_5752,N_4506);
or U8518 (N_8518,N_2426,N_6163);
xnor U8519 (N_8519,N_4389,N_800);
nor U8520 (N_8520,N_10,N_3377);
nor U8521 (N_8521,N_5708,N_3641);
nor U8522 (N_8522,N_1525,N_6079);
and U8523 (N_8523,N_3437,N_1278);
xor U8524 (N_8524,N_2432,N_5683);
and U8525 (N_8525,N_2591,N_1221);
xnor U8526 (N_8526,N_4826,N_1273);
nand U8527 (N_8527,N_2767,N_5149);
nand U8528 (N_8528,N_5896,N_2609);
nand U8529 (N_8529,N_1636,N_305);
and U8530 (N_8530,N_3110,N_987);
and U8531 (N_8531,N_4864,N_5042);
and U8532 (N_8532,N_6181,N_966);
xnor U8533 (N_8533,N_2714,N_1751);
nor U8534 (N_8534,N_3875,N_5020);
nor U8535 (N_8535,N_219,N_1456);
and U8536 (N_8536,N_6188,N_2710);
nor U8537 (N_8537,N_984,N_350);
or U8538 (N_8538,N_4476,N_3276);
or U8539 (N_8539,N_2414,N_4223);
xnor U8540 (N_8540,N_2617,N_4800);
nor U8541 (N_8541,N_3890,N_3586);
nor U8542 (N_8542,N_5107,N_3964);
nand U8543 (N_8543,N_2981,N_808);
and U8544 (N_8544,N_4515,N_1826);
xnor U8545 (N_8545,N_5859,N_2523);
nand U8546 (N_8546,N_4712,N_3227);
nor U8547 (N_8547,N_618,N_5664);
and U8548 (N_8548,N_5400,N_5793);
nand U8549 (N_8549,N_4981,N_4933);
and U8550 (N_8550,N_4732,N_2467);
nand U8551 (N_8551,N_3439,N_1319);
nor U8552 (N_8552,N_232,N_5595);
or U8553 (N_8553,N_2502,N_250);
and U8554 (N_8554,N_1155,N_5178);
xor U8555 (N_8555,N_5836,N_1533);
xor U8556 (N_8556,N_5608,N_1804);
xnor U8557 (N_8557,N_4249,N_3963);
nand U8558 (N_8558,N_4773,N_2957);
xor U8559 (N_8559,N_1847,N_1612);
nand U8560 (N_8560,N_6058,N_5521);
nand U8561 (N_8561,N_3755,N_939);
and U8562 (N_8562,N_4434,N_4033);
xnor U8563 (N_8563,N_2896,N_3923);
or U8564 (N_8564,N_3565,N_695);
or U8565 (N_8565,N_493,N_2808);
xor U8566 (N_8566,N_2859,N_3933);
and U8567 (N_8567,N_1596,N_659);
nand U8568 (N_8568,N_2562,N_1519);
xor U8569 (N_8569,N_2577,N_5777);
xnor U8570 (N_8570,N_3447,N_2616);
xnor U8571 (N_8571,N_1619,N_5056);
and U8572 (N_8572,N_1885,N_5642);
and U8573 (N_8573,N_3551,N_1233);
and U8574 (N_8574,N_2364,N_5968);
or U8575 (N_8575,N_2373,N_227);
nor U8576 (N_8576,N_6194,N_1473);
nand U8577 (N_8577,N_4454,N_5171);
nand U8578 (N_8578,N_4425,N_2717);
nand U8579 (N_8579,N_1093,N_2915);
xnor U8580 (N_8580,N_1571,N_2498);
and U8581 (N_8581,N_5926,N_172);
nor U8582 (N_8582,N_1096,N_5232);
xnor U8583 (N_8583,N_2387,N_3352);
and U8584 (N_8584,N_3349,N_1394);
and U8585 (N_8585,N_5445,N_3937);
nor U8586 (N_8586,N_3119,N_2962);
nor U8587 (N_8587,N_3415,N_1834);
and U8588 (N_8588,N_1188,N_2355);
or U8589 (N_8589,N_2813,N_1005);
xor U8590 (N_8590,N_5726,N_5487);
nand U8591 (N_8591,N_3492,N_87);
nand U8592 (N_8592,N_482,N_3983);
xor U8593 (N_8593,N_2090,N_1028);
nand U8594 (N_8594,N_6037,N_1972);
and U8595 (N_8595,N_2460,N_2015);
nand U8596 (N_8596,N_5587,N_2627);
or U8597 (N_8597,N_1461,N_4539);
xnor U8598 (N_8598,N_369,N_2526);
or U8599 (N_8599,N_1926,N_449);
nor U8600 (N_8600,N_3667,N_5384);
or U8601 (N_8601,N_5228,N_1263);
or U8602 (N_8602,N_5022,N_4651);
xnor U8603 (N_8603,N_3545,N_5800);
or U8604 (N_8604,N_486,N_5408);
nor U8605 (N_8605,N_412,N_5274);
xor U8606 (N_8606,N_1080,N_2810);
xor U8607 (N_8607,N_409,N_2096);
or U8608 (N_8608,N_2178,N_6184);
nand U8609 (N_8609,N_2959,N_2904);
or U8610 (N_8610,N_900,N_4043);
xor U8611 (N_8611,N_2116,N_410);
nand U8612 (N_8612,N_5147,N_118);
xnor U8613 (N_8613,N_311,N_5850);
or U8614 (N_8614,N_1655,N_2036);
and U8615 (N_8615,N_3514,N_4207);
nand U8616 (N_8616,N_801,N_5697);
xnor U8617 (N_8617,N_6212,N_5446);
or U8618 (N_8618,N_3074,N_1397);
nand U8619 (N_8619,N_5840,N_3388);
xor U8620 (N_8620,N_3435,N_1243);
or U8621 (N_8621,N_4935,N_2185);
and U8622 (N_8622,N_2046,N_5555);
and U8623 (N_8623,N_4988,N_3678);
or U8624 (N_8624,N_355,N_785);
nor U8625 (N_8625,N_6093,N_3469);
xor U8626 (N_8626,N_2312,N_4097);
nand U8627 (N_8627,N_2095,N_1331);
nor U8628 (N_8628,N_5083,N_2486);
or U8629 (N_8629,N_3405,N_1657);
xor U8630 (N_8630,N_2038,N_2418);
nand U8631 (N_8631,N_5950,N_3059);
and U8632 (N_8632,N_3215,N_4113);
xnor U8633 (N_8633,N_655,N_4812);
and U8634 (N_8634,N_240,N_5100);
nor U8635 (N_8635,N_6021,N_2055);
or U8636 (N_8636,N_2396,N_4482);
nand U8637 (N_8637,N_621,N_3455);
nor U8638 (N_8638,N_633,N_2225);
nor U8639 (N_8639,N_2166,N_4302);
nor U8640 (N_8640,N_2441,N_1586);
nor U8641 (N_8641,N_642,N_4322);
nor U8642 (N_8642,N_3355,N_1378);
nor U8643 (N_8643,N_2581,N_529);
nor U8644 (N_8644,N_979,N_4010);
or U8645 (N_8645,N_1654,N_3406);
nand U8646 (N_8646,N_2789,N_1140);
or U8647 (N_8647,N_4604,N_6231);
nand U8648 (N_8648,N_5356,N_634);
or U8649 (N_8649,N_4721,N_2969);
xor U8650 (N_8650,N_1566,N_4226);
xor U8651 (N_8651,N_3166,N_4911);
nand U8652 (N_8652,N_1952,N_5206);
nand U8653 (N_8653,N_1280,N_390);
nor U8654 (N_8654,N_4583,N_1927);
xnor U8655 (N_8655,N_1445,N_5216);
and U8656 (N_8656,N_269,N_1146);
or U8657 (N_8657,N_6168,N_2668);
and U8658 (N_8658,N_3211,N_2084);
xor U8659 (N_8659,N_3042,N_2779);
nand U8660 (N_8660,N_239,N_3247);
nand U8661 (N_8661,N_5231,N_1117);
nor U8662 (N_8662,N_3859,N_2263);
or U8663 (N_8663,N_1017,N_1658);
nor U8664 (N_8664,N_2922,N_1161);
or U8665 (N_8665,N_3039,N_1928);
and U8666 (N_8666,N_4627,N_1390);
and U8667 (N_8667,N_5972,N_5761);
and U8668 (N_8668,N_1754,N_5841);
or U8669 (N_8669,N_5004,N_3154);
or U8670 (N_8670,N_6180,N_1881);
nand U8671 (N_8671,N_2894,N_6205);
and U8672 (N_8672,N_3420,N_6063);
nor U8673 (N_8673,N_2924,N_5295);
nand U8674 (N_8674,N_3892,N_37);
or U8675 (N_8675,N_4753,N_1417);
and U8676 (N_8676,N_3692,N_1050);
or U8677 (N_8677,N_3204,N_2734);
or U8678 (N_8678,N_222,N_3689);
nand U8679 (N_8679,N_5940,N_5997);
or U8680 (N_8680,N_4606,N_4510);
or U8681 (N_8681,N_3936,N_2956);
or U8682 (N_8682,N_950,N_6169);
and U8683 (N_8683,N_1949,N_1908);
nor U8684 (N_8684,N_2545,N_5048);
or U8685 (N_8685,N_685,N_509);
nand U8686 (N_8686,N_6150,N_1474);
or U8687 (N_8687,N_1055,N_2794);
nand U8688 (N_8688,N_2440,N_357);
xnor U8689 (N_8689,N_814,N_606);
nor U8690 (N_8690,N_4897,N_3807);
and U8691 (N_8691,N_6016,N_2622);
nor U8692 (N_8692,N_5789,N_4644);
nand U8693 (N_8693,N_5932,N_4227);
nor U8694 (N_8694,N_930,N_4143);
and U8695 (N_8695,N_5250,N_1923);
and U8696 (N_8696,N_3520,N_5155);
and U8697 (N_8697,N_1683,N_1412);
nand U8698 (N_8698,N_4020,N_1259);
or U8699 (N_8699,N_1615,N_3992);
nor U8700 (N_8700,N_4144,N_4954);
and U8701 (N_8701,N_1284,N_6143);
nand U8702 (N_8702,N_5209,N_5193);
nand U8703 (N_8703,N_2463,N_2974);
nor U8704 (N_8704,N_3141,N_3874);
and U8705 (N_8705,N_2764,N_2111);
xor U8706 (N_8706,N_1932,N_2786);
xor U8707 (N_8707,N_2645,N_1842);
xor U8708 (N_8708,N_4706,N_1938);
nand U8709 (N_8709,N_3510,N_1439);
and U8710 (N_8710,N_3328,N_4222);
or U8711 (N_8711,N_2262,N_3740);
nor U8712 (N_8712,N_1375,N_5403);
and U8713 (N_8713,N_3030,N_3323);
nor U8714 (N_8714,N_2499,N_186);
xor U8715 (N_8715,N_2629,N_2964);
and U8716 (N_8716,N_1421,N_3381);
or U8717 (N_8717,N_5647,N_16);
nand U8718 (N_8718,N_2353,N_4021);
and U8719 (N_8719,N_4658,N_3849);
nor U8720 (N_8720,N_2380,N_5344);
or U8721 (N_8721,N_5848,N_3017);
xnor U8722 (N_8722,N_140,N_2372);
nand U8723 (N_8723,N_1824,N_3361);
xnor U8724 (N_8724,N_1542,N_2180);
and U8725 (N_8725,N_82,N_5660);
and U8726 (N_8726,N_9,N_4587);
or U8727 (N_8727,N_1699,N_246);
nor U8728 (N_8728,N_3508,N_131);
or U8729 (N_8729,N_3637,N_1722);
nor U8730 (N_8730,N_3806,N_570);
and U8731 (N_8731,N_83,N_1310);
and U8732 (N_8732,N_3449,N_3233);
and U8733 (N_8733,N_5552,N_89);
nor U8734 (N_8734,N_4077,N_2776);
nor U8735 (N_8735,N_1271,N_3149);
xnor U8736 (N_8736,N_2277,N_5485);
and U8737 (N_8737,N_4253,N_6101);
or U8738 (N_8738,N_5286,N_1613);
and U8739 (N_8739,N_2231,N_1713);
and U8740 (N_8740,N_3648,N_5098);
or U8741 (N_8741,N_4829,N_3394);
and U8742 (N_8742,N_2863,N_3704);
nand U8743 (N_8743,N_4750,N_6011);
nor U8744 (N_8744,N_2469,N_5919);
xor U8745 (N_8745,N_3948,N_1924);
and U8746 (N_8746,N_4558,N_2667);
nor U8747 (N_8747,N_4557,N_5716);
and U8748 (N_8748,N_2146,N_3386);
nand U8749 (N_8749,N_1832,N_236);
nand U8750 (N_8750,N_3077,N_4886);
and U8751 (N_8751,N_5520,N_3283);
xor U8752 (N_8752,N_4404,N_3272);
and U8753 (N_8753,N_6060,N_1414);
nor U8754 (N_8754,N_5186,N_3460);
xnor U8755 (N_8755,N_3489,N_2619);
or U8756 (N_8756,N_80,N_2521);
nor U8757 (N_8757,N_2780,N_1291);
nor U8758 (N_8758,N_6185,N_4894);
nand U8759 (N_8759,N_3609,N_2010);
and U8760 (N_8760,N_4107,N_3961);
xor U8761 (N_8761,N_5812,N_5695);
xnor U8762 (N_8762,N_4910,N_1534);
xnor U8763 (N_8763,N_3151,N_2775);
xor U8764 (N_8764,N_3005,N_6029);
nor U8765 (N_8765,N_4123,N_1537);
nand U8766 (N_8766,N_1410,N_5041);
nand U8767 (N_8767,N_3783,N_941);
and U8768 (N_8768,N_1786,N_2101);
or U8769 (N_8769,N_2439,N_3810);
xor U8770 (N_8770,N_3006,N_1643);
or U8771 (N_8771,N_1463,N_3973);
nor U8772 (N_8772,N_5636,N_4438);
nor U8773 (N_8773,N_3927,N_4287);
nor U8774 (N_8774,N_3333,N_2989);
nand U8775 (N_8775,N_4463,N_213);
nor U8776 (N_8776,N_2479,N_386);
or U8777 (N_8777,N_379,N_3379);
and U8778 (N_8778,N_2459,N_5461);
and U8779 (N_8779,N_4291,N_5370);
or U8780 (N_8780,N_4899,N_4700);
nand U8781 (N_8781,N_167,N_5671);
xor U8782 (N_8782,N_5545,N_1986);
nand U8783 (N_8783,N_2608,N_1388);
xor U8784 (N_8784,N_2173,N_3072);
and U8785 (N_8785,N_2007,N_2105);
nor U8786 (N_8786,N_1400,N_367);
and U8787 (N_8787,N_6001,N_3943);
or U8788 (N_8788,N_1185,N_5244);
or U8789 (N_8789,N_3932,N_5341);
nor U8790 (N_8790,N_2891,N_1389);
nor U8791 (N_8791,N_3922,N_3229);
nand U8792 (N_8792,N_3914,N_1472);
nand U8793 (N_8793,N_6062,N_453);
xnor U8794 (N_8794,N_1311,N_5008);
xor U8795 (N_8795,N_2935,N_2584);
xor U8796 (N_8796,N_3067,N_5402);
nor U8797 (N_8797,N_1198,N_3799);
nand U8798 (N_8798,N_4239,N_4591);
nand U8799 (N_8799,N_1360,N_69);
nor U8800 (N_8800,N_3002,N_242);
and U8801 (N_8801,N_403,N_878);
nand U8802 (N_8802,N_3273,N_4171);
or U8803 (N_8803,N_326,N_2559);
nand U8804 (N_8804,N_3506,N_4376);
nor U8805 (N_8805,N_380,N_995);
nor U8806 (N_8806,N_546,N_3981);
xor U8807 (N_8807,N_3535,N_1024);
and U8808 (N_8808,N_4729,N_396);
xnor U8809 (N_8809,N_4048,N_5951);
or U8810 (N_8810,N_152,N_1922);
nand U8811 (N_8811,N_3065,N_5176);
xor U8812 (N_8812,N_1129,N_415);
and U8813 (N_8813,N_171,N_976);
or U8814 (N_8814,N_4838,N_4363);
nor U8815 (N_8815,N_5632,N_2700);
nor U8816 (N_8816,N_4030,N_2386);
or U8817 (N_8817,N_651,N_4683);
xnor U8818 (N_8818,N_5467,N_3669);
nor U8819 (N_8819,N_2290,N_6164);
nor U8820 (N_8820,N_1808,N_6028);
nand U8821 (N_8821,N_6162,N_3980);
xnor U8822 (N_8822,N_147,N_4162);
and U8823 (N_8823,N_3201,N_2809);
nand U8824 (N_8824,N_1973,N_601);
nor U8825 (N_8825,N_746,N_3858);
and U8826 (N_8826,N_1234,N_5690);
or U8827 (N_8827,N_611,N_5533);
nor U8828 (N_8828,N_2836,N_3727);
nor U8829 (N_8829,N_2801,N_582);
nand U8830 (N_8830,N_4343,N_5942);
xnor U8831 (N_8831,N_1995,N_4320);
nand U8832 (N_8832,N_256,N_2348);
xnor U8833 (N_8833,N_3410,N_4096);
xnor U8834 (N_8834,N_5975,N_4531);
or U8835 (N_8835,N_1640,N_942);
nor U8836 (N_8836,N_29,N_5933);
nand U8837 (N_8837,N_4177,N_5464);
xnor U8838 (N_8838,N_2106,N_5291);
and U8839 (N_8839,N_2551,N_1184);
xnor U8840 (N_8840,N_394,N_5728);
nor U8841 (N_8841,N_5051,N_1352);
nand U8842 (N_8842,N_5152,N_3773);
nand U8843 (N_8843,N_4012,N_6045);
nand U8844 (N_8844,N_724,N_2866);
nor U8845 (N_8845,N_1289,N_1104);
or U8846 (N_8846,N_4325,N_1959);
xor U8847 (N_8847,N_3131,N_3391);
nor U8848 (N_8848,N_3566,N_4726);
xor U8849 (N_8849,N_5047,N_3109);
and U8850 (N_8850,N_212,N_4661);
nand U8851 (N_8851,N_6153,N_267);
and U8852 (N_8852,N_3907,N_3392);
and U8853 (N_8853,N_1989,N_6238);
xnor U8854 (N_8854,N_284,N_3779);
or U8855 (N_8855,N_1265,N_1275);
nor U8856 (N_8856,N_3638,N_4076);
xnor U8857 (N_8857,N_6215,N_6109);
nor U8858 (N_8858,N_2954,N_4125);
and U8859 (N_8859,N_179,N_4026);
nor U8860 (N_8860,N_4154,N_5347);
xnor U8861 (N_8861,N_2226,N_899);
and U8862 (N_8862,N_358,N_4925);
or U8863 (N_8863,N_2219,N_5268);
xor U8864 (N_8864,N_5631,N_1026);
nor U8865 (N_8865,N_3999,N_4196);
nand U8866 (N_8866,N_2248,N_1934);
nor U8867 (N_8867,N_1087,N_760);
or U8868 (N_8868,N_1890,N_4880);
or U8869 (N_8869,N_5422,N_1440);
nor U8870 (N_8870,N_3670,N_4440);
and U8871 (N_8871,N_2733,N_5364);
or U8872 (N_8872,N_1053,N_4364);
nor U8873 (N_8873,N_3567,N_1999);
xor U8874 (N_8874,N_153,N_4767);
xnor U8875 (N_8875,N_3596,N_1309);
nor U8876 (N_8876,N_5126,N_1905);
nor U8877 (N_8877,N_75,N_686);
or U8878 (N_8878,N_5351,N_362);
xnor U8879 (N_8879,N_3063,N_3921);
nand U8880 (N_8880,N_4755,N_3091);
or U8881 (N_8881,N_170,N_4444);
xnor U8882 (N_8882,N_6218,N_2588);
xor U8883 (N_8883,N_4852,N_3085);
and U8884 (N_8884,N_2031,N_2865);
nor U8885 (N_8885,N_4237,N_1888);
or U8886 (N_8886,N_4671,N_159);
nand U8887 (N_8887,N_1486,N_791);
xor U8888 (N_8888,N_2196,N_654);
or U8889 (N_8889,N_2988,N_5213);
nand U8890 (N_8890,N_3178,N_5669);
or U8891 (N_8891,N_4507,N_2634);
nor U8892 (N_8892,N_2127,N_4448);
nor U8893 (N_8893,N_3606,N_429);
nand U8894 (N_8894,N_3061,N_1976);
and U8895 (N_8895,N_4167,N_1343);
and U8896 (N_8896,N_5634,N_584);
and U8897 (N_8897,N_856,N_4367);
xor U8898 (N_8898,N_411,N_1509);
xor U8899 (N_8899,N_448,N_1939);
nand U8900 (N_8900,N_2246,N_1610);
xor U8901 (N_8901,N_961,N_5267);
nand U8902 (N_8902,N_3580,N_5472);
nand U8903 (N_8903,N_4168,N_4458);
and U8904 (N_8904,N_5760,N_4433);
or U8905 (N_8905,N_4311,N_4572);
xnor U8906 (N_8906,N_278,N_612);
nor U8907 (N_8907,N_4234,N_2887);
or U8908 (N_8908,N_1305,N_1241);
nor U8909 (N_8909,N_4749,N_2707);
nor U8910 (N_8910,N_4427,N_40);
nand U8911 (N_8911,N_47,N_3867);
xor U8912 (N_8912,N_4856,N_5680);
or U8913 (N_8913,N_5352,N_676);
xor U8914 (N_8914,N_5073,N_1679);
and U8915 (N_8915,N_5538,N_5769);
nor U8916 (N_8916,N_4736,N_4552);
or U8917 (N_8917,N_6111,N_2930);
xor U8918 (N_8918,N_3760,N_888);
xnor U8919 (N_8919,N_155,N_4111);
or U8920 (N_8920,N_848,N_896);
nand U8921 (N_8921,N_2961,N_2073);
nor U8922 (N_8922,N_792,N_6071);
nand U8923 (N_8923,N_5322,N_433);
and U8924 (N_8924,N_1029,N_5430);
and U8925 (N_8925,N_461,N_104);
nor U8926 (N_8926,N_2238,N_2306);
and U8927 (N_8927,N_3924,N_4090);
nand U8928 (N_8928,N_3287,N_3839);
and U8929 (N_8929,N_3376,N_2247);
or U8930 (N_8930,N_1957,N_3033);
xor U8931 (N_8931,N_3878,N_4522);
xnor U8932 (N_8932,N_732,N_389);
nand U8933 (N_8933,N_5154,N_5699);
nand U8934 (N_8934,N_1354,N_1252);
xor U8935 (N_8935,N_3497,N_117);
nand U8936 (N_8936,N_2131,N_2806);
or U8937 (N_8937,N_5348,N_4976);
nand U8938 (N_8938,N_5059,N_4689);
nor U8939 (N_8939,N_4412,N_5666);
or U8940 (N_8940,N_5778,N_251);
and U8941 (N_8941,N_5030,N_3357);
xor U8942 (N_8942,N_4503,N_4091);
nor U8943 (N_8943,N_5229,N_6120);
and U8944 (N_8944,N_4922,N_1262);
nor U8945 (N_8945,N_2932,N_5721);
nor U8946 (N_8946,N_4278,N_3432);
nand U8947 (N_8947,N_3170,N_3309);
nand U8948 (N_8948,N_5161,N_1174);
xor U8949 (N_8949,N_1176,N_3680);
or U8950 (N_8950,N_5584,N_1678);
nand U8951 (N_8951,N_4445,N_4420);
xnor U8952 (N_8952,N_1733,N_5908);
xnor U8953 (N_8953,N_5246,N_1563);
xor U8954 (N_8954,N_2676,N_202);
nor U8955 (N_8955,N_492,N_1629);
nor U8956 (N_8956,N_4198,N_5745);
nor U8957 (N_8957,N_5661,N_3419);
or U8958 (N_8958,N_5313,N_3529);
xnor U8959 (N_8959,N_2350,N_5542);
and U8960 (N_8960,N_2555,N_2281);
or U8961 (N_8961,N_3307,N_5005);
nor U8962 (N_8962,N_940,N_2854);
nand U8963 (N_8963,N_2626,N_6070);
and U8964 (N_8964,N_4853,N_1089);
nand U8965 (N_8965,N_2337,N_6103);
nor U8966 (N_8966,N_417,N_4157);
nor U8967 (N_8967,N_7,N_3448);
nand U8968 (N_8968,N_5882,N_1302);
and U8969 (N_8969,N_5131,N_5398);
nand U8970 (N_8970,N_5329,N_2172);
or U8971 (N_8971,N_3209,N_779);
xnor U8972 (N_8972,N_1223,N_4416);
or U8973 (N_8973,N_220,N_1961);
or U8974 (N_8974,N_6057,N_1652);
and U8975 (N_8975,N_28,N_5604);
xor U8976 (N_8976,N_1788,N_4031);
xor U8977 (N_8977,N_1910,N_615);
nor U8978 (N_8978,N_4797,N_2575);
or U8979 (N_8979,N_276,N_5390);
nor U8980 (N_8980,N_1673,N_6226);
and U8981 (N_8981,N_845,N_5790);
and U8982 (N_8982,N_5741,N_4742);
and U8983 (N_8983,N_3418,N_2724);
or U8984 (N_8984,N_4574,N_2681);
nor U8985 (N_8985,N_1984,N_3044);
or U8986 (N_8986,N_1935,N_543);
nand U8987 (N_8987,N_4036,N_3177);
xnor U8988 (N_8988,N_5027,N_5883);
and U8989 (N_8989,N_5611,N_528);
nand U8990 (N_8990,N_1115,N_6177);
or U8991 (N_8991,N_3729,N_5324);
xor U8992 (N_8992,N_499,N_1098);
xnor U8993 (N_8993,N_882,N_5102);
or U8994 (N_8994,N_4602,N_2514);
nor U8995 (N_8995,N_3957,N_3047);
xor U8996 (N_8996,N_2578,N_5441);
nor U8997 (N_8997,N_5101,N_3548);
and U8998 (N_8998,N_6221,N_2050);
or U8999 (N_8999,N_3055,N_2271);
nor U9000 (N_9000,N_534,N_3895);
or U9001 (N_9001,N_6151,N_1232);
nor U9002 (N_9002,N_376,N_4266);
nand U9003 (N_9003,N_2987,N_4908);
nor U9004 (N_9004,N_5173,N_2704);
or U9005 (N_9005,N_1947,N_1994);
xnor U9006 (N_9006,N_566,N_1192);
nand U9007 (N_9007,N_1850,N_5143);
or U9008 (N_9008,N_5168,N_1338);
nand U9009 (N_9009,N_6032,N_5438);
nor U9010 (N_9010,N_2027,N_2110);
nor U9011 (N_9011,N_5540,N_3499);
or U9012 (N_9012,N_3029,N_2174);
xnor U9013 (N_9013,N_4846,N_2209);
nand U9014 (N_9014,N_2220,N_2201);
xnor U9015 (N_9015,N_3262,N_3475);
and U9016 (N_9016,N_5591,N_3749);
xnor U9017 (N_9017,N_4748,N_2715);
xnor U9018 (N_9018,N_1756,N_5913);
nand U9019 (N_9019,N_2690,N_4280);
xnor U9020 (N_9020,N_261,N_5853);
and U9021 (N_9021,N_196,N_3848);
and U9022 (N_9022,N_3996,N_1991);
nor U9023 (N_9023,N_191,N_5624);
or U9024 (N_9024,N_5717,N_3456);
and U9025 (N_9025,N_5938,N_1135);
and U9026 (N_9026,N_1150,N_5119);
nand U9027 (N_9027,N_894,N_974);
xnor U9028 (N_9028,N_3057,N_2334);
nand U9029 (N_9029,N_5393,N_530);
nand U9030 (N_9030,N_3053,N_1724);
nor U9031 (N_9031,N_4566,N_479);
xnor U9032 (N_9032,N_2942,N_2838);
or U9033 (N_9033,N_1105,N_1326);
nor U9034 (N_9034,N_4796,N_5496);
xor U9035 (N_9035,N_2148,N_4540);
and U9036 (N_9036,N_4738,N_1272);
and U9037 (N_9037,N_6199,N_1644);
xnor U9038 (N_9038,N_1067,N_4081);
xor U9039 (N_9039,N_1708,N_56);
nor U9040 (N_9040,N_5498,N_3612);
nor U9041 (N_9041,N_3687,N_2713);
xor U9042 (N_9042,N_3159,N_373);
and U9043 (N_9043,N_6167,N_616);
nand U9044 (N_9044,N_3786,N_2943);
and U9045 (N_9045,N_804,N_2741);
or U9046 (N_9046,N_1711,N_4550);
nor U9047 (N_9047,N_2843,N_5723);
xor U9048 (N_9048,N_3998,N_4372);
xnor U9049 (N_9049,N_5563,N_4176);
or U9050 (N_9050,N_4598,N_365);
and U9051 (N_9051,N_5720,N_4236);
or U9052 (N_9052,N_4224,N_5140);
or U9053 (N_9053,N_3416,N_2599);
xnor U9054 (N_9054,N_5084,N_5242);
and U9055 (N_9055,N_1482,N_1323);
or U9056 (N_9056,N_1287,N_4259);
xnor U9057 (N_9057,N_2862,N_6178);
xnor U9058 (N_9058,N_238,N_3618);
nand U9059 (N_9059,N_339,N_2186);
and U9060 (N_9060,N_3748,N_347);
or U9061 (N_9061,N_1656,N_4359);
xor U9062 (N_9062,N_2255,N_1090);
nor U9063 (N_9063,N_1381,N_4761);
and U9064 (N_9064,N_148,N_3534);
and U9065 (N_9065,N_2003,N_970);
nand U9066 (N_9066,N_1466,N_691);
xor U9067 (N_9067,N_1581,N_6038);
or U9068 (N_9068,N_1092,N_109);
xnor U9069 (N_9069,N_3186,N_4347);
and U9070 (N_9070,N_4519,N_2819);
and U9071 (N_9071,N_842,N_70);
xor U9072 (N_9072,N_2237,N_4579);
and U9073 (N_9073,N_5685,N_3731);
nor U9074 (N_9074,N_4117,N_5308);
xor U9075 (N_9075,N_1762,N_4201);
and U9076 (N_9076,N_3466,N_1152);
xor U9077 (N_9077,N_3158,N_3062);
and U9078 (N_9078,N_5511,N_1182);
xnor U9079 (N_9079,N_4690,N_720);
nand U9080 (N_9080,N_1775,N_904);
nor U9081 (N_9081,N_2908,N_1755);
or U9082 (N_9082,N_2939,N_175);
and U9083 (N_9083,N_2918,N_3616);
xnor U9084 (N_9084,N_2462,N_4116);
nor U9085 (N_9085,N_545,N_1631);
or U9086 (N_9086,N_3306,N_2568);
or U9087 (N_9087,N_3396,N_4067);
xor U9088 (N_9088,N_4702,N_1599);
nor U9089 (N_9089,N_1997,N_4939);
and U9090 (N_9090,N_1266,N_6206);
or U9091 (N_9091,N_146,N_1797);
nor U9092 (N_9092,N_4969,N_2405);
or U9093 (N_9093,N_2674,N_943);
nor U9094 (N_9094,N_1944,N_3977);
or U9095 (N_9095,N_2252,N_5391);
nand U9096 (N_9096,N_218,N_2122);
nor U9097 (N_9097,N_4739,N_2320);
nor U9098 (N_9098,N_4446,N_2216);
and U9099 (N_9099,N_683,N_1851);
nand U9100 (N_9100,N_5705,N_4385);
nand U9101 (N_9101,N_5702,N_4788);
and U9102 (N_9102,N_3734,N_1987);
nor U9103 (N_9103,N_556,N_129);
nand U9104 (N_9104,N_5931,N_2878);
and U9105 (N_9105,N_2958,N_18);
nand U9106 (N_9106,N_1761,N_4831);
xor U9107 (N_9107,N_627,N_2669);
xnor U9108 (N_9108,N_3438,N_1433);
xnor U9109 (N_9109,N_5592,N_4486);
nor U9110 (N_9110,N_733,N_2394);
nor U9111 (N_9111,N_3543,N_3078);
and U9112 (N_9112,N_1779,N_3505);
xnor U9113 (N_9113,N_5145,N_5546);
nor U9114 (N_9114,N_6074,N_1645);
nand U9115 (N_9115,N_3335,N_784);
nor U9116 (N_9116,N_4536,N_715);
xnor U9117 (N_9117,N_3950,N_3574);
and U9118 (N_9118,N_5350,N_1829);
nand U9119 (N_9119,N_5361,N_2573);
nand U9120 (N_9120,N_6229,N_5255);
nand U9121 (N_9121,N_3045,N_4814);
or U9122 (N_9122,N_5976,N_1231);
xor U9123 (N_9123,N_354,N_79);
nand U9124 (N_9124,N_3621,N_4769);
xor U9125 (N_9125,N_1327,N_1349);
xor U9126 (N_9126,N_1520,N_3735);
and U9127 (N_9127,N_4409,N_4578);
and U9128 (N_9128,N_1730,N_1863);
or U9129 (N_9129,N_3947,N_698);
nor U9130 (N_9130,N_1819,N_653);
xnor U9131 (N_9131,N_5824,N_2119);
xor U9132 (N_9132,N_712,N_1139);
or U9133 (N_9133,N_6125,N_2745);
or U9134 (N_9134,N_3778,N_1183);
nand U9135 (N_9135,N_1404,N_4139);
or U9136 (N_9136,N_4383,N_5739);
and U9137 (N_9137,N_3252,N_5211);
and U9138 (N_9138,N_6159,N_1806);
xor U9139 (N_9139,N_5123,N_275);
and U9140 (N_9140,N_3117,N_4357);
xnor U9141 (N_9141,N_5843,N_1334);
nor U9142 (N_9142,N_3556,N_1639);
or U9143 (N_9143,N_2315,N_2850);
nand U9144 (N_9144,N_3491,N_3675);
xor U9145 (N_9145,N_3099,N_2360);
xnor U9146 (N_9146,N_6196,N_2787);
nand U9147 (N_9147,N_1685,N_5736);
and U9148 (N_9148,N_1968,N_3220);
xnor U9149 (N_9149,N_4779,N_2076);
nor U9150 (N_9150,N_324,N_3643);
nor U9151 (N_9151,N_5302,N_442);
or U9152 (N_9152,N_5007,N_1725);
nand U9153 (N_9153,N_3915,N_838);
nand U9154 (N_9154,N_834,N_4883);
nand U9155 (N_9155,N_254,N_1998);
xor U9156 (N_9156,N_1954,N_1240);
nor U9157 (N_9157,N_2967,N_2044);
nand U9158 (N_9158,N_3308,N_1426);
xnor U9159 (N_9159,N_1195,N_2711);
or U9160 (N_9160,N_206,N_4041);
nor U9161 (N_9161,N_5502,N_2560);
nand U9162 (N_9162,N_4460,N_919);
and U9163 (N_9163,N_446,N_113);
xnor U9164 (N_9164,N_52,N_336);
or U9165 (N_9165,N_2310,N_2013);
or U9166 (N_9166,N_6207,N_4072);
or U9167 (N_9167,N_1464,N_2458);
nand U9168 (N_9168,N_4407,N_1348);
nor U9169 (N_9169,N_2163,N_3350);
nor U9170 (N_9170,N_1171,N_5330);
and U9171 (N_9171,N_3897,N_31);
nand U9172 (N_9172,N_2243,N_4609);
xor U9173 (N_9173,N_3656,N_1015);
and U9174 (N_9174,N_2856,N_757);
and U9175 (N_9175,N_105,N_6027);
and U9176 (N_9176,N_5458,N_2834);
or U9177 (N_9177,N_1766,N_4576);
nor U9178 (N_9178,N_3654,N_914);
nand U9179 (N_9179,N_5583,N_3528);
xor U9180 (N_9180,N_2656,N_5136);
or U9181 (N_9181,N_2795,N_5582);
nand U9182 (N_9182,N_2692,N_422);
nand U9183 (N_9183,N_4551,N_1567);
xnor U9184 (N_9184,N_2269,N_2886);
nand U9185 (N_9185,N_3464,N_3036);
nand U9186 (N_9186,N_2489,N_727);
or U9187 (N_9187,N_5895,N_3326);
nand U9188 (N_9188,N_1950,N_2515);
and U9189 (N_9189,N_4040,N_982);
nor U9190 (N_9190,N_1918,N_5982);
xnor U9191 (N_9191,N_1667,N_2666);
nor U9192 (N_9192,N_6246,N_2412);
nor U9193 (N_9193,N_3887,N_2528);
or U9194 (N_9194,N_163,N_5338);
nand U9195 (N_9195,N_3739,N_6128);
and U9196 (N_9196,N_1682,N_2093);
xnor U9197 (N_9197,N_3268,N_3254);
xnor U9198 (N_9198,N_1306,N_2788);
or U9199 (N_9199,N_6217,N_1151);
and U9200 (N_9200,N_3690,N_3626);
and U9201 (N_9201,N_5941,N_6106);
nand U9202 (N_9202,N_4901,N_1335);
or U9203 (N_9203,N_2207,N_39);
nor U9204 (N_9204,N_262,N_643);
nand U9205 (N_9205,N_811,N_1760);
or U9206 (N_9206,N_4134,N_4264);
nand U9207 (N_9207,N_5663,N_5256);
and U9208 (N_9208,N_2823,N_5093);
nand U9209 (N_9209,N_2039,N_4926);
xnor U9210 (N_9210,N_4303,N_3194);
and U9211 (N_9211,N_5532,N_5907);
or U9212 (N_9212,N_5687,N_4451);
or U9213 (N_9213,N_431,N_5142);
xor U9214 (N_9214,N_5574,N_1043);
xnor U9215 (N_9215,N_371,N_4360);
xor U9216 (N_9216,N_2876,N_3784);
or U9217 (N_9217,N_3083,N_3798);
xor U9218 (N_9218,N_1099,N_2735);
and U9219 (N_9219,N_65,N_5906);
or U9220 (N_9220,N_3237,N_4724);
or U9221 (N_9221,N_823,N_4028);
xnor U9222 (N_9222,N_577,N_91);
and U9223 (N_9223,N_5673,N_1606);
nand U9224 (N_9224,N_4951,N_3193);
xor U9225 (N_9225,N_2477,N_3080);
nand U9226 (N_9226,N_3341,N_2571);
xnor U9227 (N_9227,N_4279,N_2330);
nand U9228 (N_9228,N_5233,N_3707);
and U9229 (N_9229,N_1459,N_2845);
nor U9230 (N_9230,N_3837,N_141);
xnor U9231 (N_9231,N_4202,N_1940);
nor U9232 (N_9232,N_640,N_3264);
nand U9233 (N_9233,N_2461,N_4523);
nand U9234 (N_9234,N_5969,N_4887);
and U9235 (N_9235,N_4233,N_3569);
nand U9236 (N_9236,N_1300,N_3108);
xor U9237 (N_9237,N_561,N_1436);
and U9238 (N_9238,N_4703,N_5103);
and U9239 (N_9239,N_1801,N_277);
and U9240 (N_9240,N_5261,N_4635);
and U9241 (N_9241,N_4909,N_3926);
nor U9242 (N_9242,N_3486,N_5993);
nor U9243 (N_9243,N_4005,N_323);
and U9244 (N_9244,N_2648,N_3713);
nor U9245 (N_9245,N_2705,N_3659);
nor U9246 (N_9246,N_631,N_5747);
nand U9247 (N_9247,N_704,N_3830);
and U9248 (N_9248,N_2662,N_2331);
xor U9249 (N_9249,N_1838,N_5419);
or U9250 (N_9250,N_1514,N_6155);
or U9251 (N_9251,N_2998,N_6179);
xor U9252 (N_9252,N_3951,N_4417);
xnor U9253 (N_9253,N_1249,N_5486);
and U9254 (N_9254,N_194,N_2454);
nor U9255 (N_9255,N_851,N_5264);
nand U9256 (N_9256,N_4694,N_4762);
and U9257 (N_9257,N_4346,N_2677);
and U9258 (N_9258,N_3028,N_5443);
nand U9259 (N_9259,N_4378,N_4297);
nor U9260 (N_9260,N_3925,N_4799);
xnor U9261 (N_9261,N_1680,N_5889);
nand U9262 (N_9262,N_5744,N_5440);
xor U9263 (N_9263,N_550,N_5991);
nor U9264 (N_9264,N_5833,N_6225);
or U9265 (N_9265,N_4356,N_4614);
xnor U9266 (N_9266,N_1522,N_4983);
nor U9267 (N_9267,N_3746,N_3831);
nor U9268 (N_9268,N_6068,N_5838);
nand U9269 (N_9269,N_4075,N_5221);
xor U9270 (N_9270,N_3949,N_344);
xor U9271 (N_9271,N_5948,N_425);
xor U9272 (N_9272,N_4178,N_2136);
nand U9273 (N_9273,N_5753,N_2165);
or U9274 (N_9274,N_5192,N_4022);
nand U9275 (N_9275,N_4152,N_2968);
nand U9276 (N_9276,N_3200,N_270);
nor U9277 (N_9277,N_5585,N_4513);
and U9278 (N_9278,N_4058,N_3216);
and U9279 (N_9279,N_487,N_2388);
xor U9280 (N_9280,N_2210,N_214);
nand U9281 (N_9281,N_5413,N_3860);
nand U9282 (N_9282,N_1515,N_4621);
and U9283 (N_9283,N_916,N_4906);
and U9284 (N_9284,N_2433,N_158);
and U9285 (N_9285,N_687,N_568);
nand U9286 (N_9286,N_1623,N_5658);
and U9287 (N_9287,N_3960,N_5879);
xnor U9288 (N_9288,N_1988,N_1442);
and U9289 (N_9289,N_1345,N_3183);
nand U9290 (N_9290,N_4172,N_4053);
or U9291 (N_9291,N_924,N_2718);
and U9292 (N_9292,N_2103,N_3458);
xor U9293 (N_9293,N_3218,N_3770);
or U9294 (N_9294,N_2919,N_895);
nand U9295 (N_9295,N_53,N_5779);
and U9296 (N_9296,N_2646,N_426);
xor U9297 (N_9297,N_5011,N_4247);
and U9298 (N_9298,N_5146,N_761);
xor U9299 (N_9299,N_1189,N_3906);
xor U9300 (N_9300,N_5873,N_1061);
and U9301 (N_9301,N_3886,N_57);
and U9302 (N_9302,N_3978,N_4251);
and U9303 (N_9303,N_4129,N_223);
and U9304 (N_9304,N_891,N_1688);
and U9305 (N_9305,N_2936,N_1852);
nand U9306 (N_9306,N_5431,N_1450);
and U9307 (N_9307,N_559,N_3971);
nand U9308 (N_9308,N_6114,N_3958);
and U9309 (N_9309,N_4973,N_4469);
nor U9310 (N_9310,N_1820,N_4087);
or U9311 (N_9311,N_3128,N_4580);
nand U9312 (N_9312,N_5864,N_859);
nand U9313 (N_9313,N_5995,N_849);
and U9314 (N_9314,N_926,N_2244);
xor U9315 (N_9315,N_2527,N_1437);
xor U9316 (N_9316,N_266,N_4146);
nand U9317 (N_9317,N_1911,N_5534);
xor U9318 (N_9318,N_5834,N_4943);
and U9319 (N_9319,N_558,N_5482);
nand U9320 (N_9320,N_2349,N_876);
xnor U9321 (N_9321,N_6126,N_2234);
nand U9322 (N_9322,N_2864,N_5077);
nor U9323 (N_9323,N_4715,N_4023);
nand U9324 (N_9324,N_5411,N_3765);
xnor U9325 (N_9325,N_1408,N_1484);
and U9326 (N_9326,N_2048,N_2404);
nor U9327 (N_9327,N_1332,N_4952);
nor U9328 (N_9328,N_466,N_1510);
and U9329 (N_9329,N_2822,N_5675);
xnor U9330 (N_9330,N_3443,N_2162);
or U9331 (N_9331,N_5802,N_6076);
nand U9332 (N_9332,N_5121,N_4893);
and U9333 (N_9333,N_2911,N_3946);
or U9334 (N_9334,N_5156,N_836);
and U9335 (N_9335,N_5927,N_3883);
xnor U9336 (N_9336,N_5425,N_2510);
or U9337 (N_9337,N_5238,N_1065);
and U9338 (N_9338,N_5525,N_963);
xor U9339 (N_9339,N_1217,N_1920);
or U9340 (N_9340,N_5358,N_4599);
and U9341 (N_9341,N_4839,N_1582);
nand U9342 (N_9342,N_3940,N_4545);
nor U9343 (N_9343,N_4571,N_5701);
xor U9344 (N_9344,N_5936,N_4439);
or U9345 (N_9345,N_2272,N_3630);
and U9346 (N_9346,N_2909,N_650);
or U9347 (N_9347,N_2321,N_2516);
xnor U9348 (N_9348,N_3153,N_3546);
nor U9349 (N_9349,N_6118,N_1763);
and U9350 (N_9350,N_5392,N_3474);
or U9351 (N_9351,N_5325,N_2056);
xor U9352 (N_9352,N_1254,N_1864);
nor U9353 (N_9353,N_3732,N_2045);
and U9354 (N_9354,N_2726,N_854);
xor U9355 (N_9355,N_1671,N_1553);
nor U9356 (N_9356,N_3258,N_3161);
nor U9357 (N_9357,N_4461,N_384);
nand U9358 (N_9358,N_6244,N_42);
nor U9359 (N_9359,N_5366,N_5260);
xor U9360 (N_9360,N_103,N_5006);
and U9361 (N_9361,N_4809,N_1700);
or U9362 (N_9362,N_1803,N_142);
nand U9363 (N_9363,N_3796,N_3610);
xor U9364 (N_9364,N_5681,N_2295);
nand U9365 (N_9365,N_4610,N_5087);
and U9366 (N_9366,N_2189,N_5823);
nand U9367 (N_9367,N_3900,N_2720);
nor U9368 (N_9368,N_62,N_4766);
and U9369 (N_9369,N_2722,N_3040);
and U9370 (N_9370,N_2480,N_4338);
and U9371 (N_9371,N_177,N_5029);
nand U9372 (N_9372,N_4987,N_6193);
nand U9373 (N_9373,N_5627,N_3202);
xor U9374 (N_9374,N_4142,N_719);
xnor U9375 (N_9375,N_3659,N_4465);
xnor U9376 (N_9376,N_4921,N_3271);
and U9377 (N_9377,N_3067,N_1677);
xnor U9378 (N_9378,N_2877,N_4147);
or U9379 (N_9379,N_3410,N_2433);
and U9380 (N_9380,N_2476,N_1118);
xor U9381 (N_9381,N_131,N_4574);
and U9382 (N_9382,N_5352,N_1555);
and U9383 (N_9383,N_3747,N_5133);
xnor U9384 (N_9384,N_894,N_1136);
or U9385 (N_9385,N_1864,N_1880);
xor U9386 (N_9386,N_4051,N_2580);
or U9387 (N_9387,N_2329,N_1186);
and U9388 (N_9388,N_2913,N_5872);
xnor U9389 (N_9389,N_710,N_5066);
xnor U9390 (N_9390,N_4338,N_478);
and U9391 (N_9391,N_5722,N_1539);
nor U9392 (N_9392,N_3718,N_3749);
nand U9393 (N_9393,N_5515,N_3840);
xor U9394 (N_9394,N_2067,N_1315);
and U9395 (N_9395,N_5459,N_2709);
xor U9396 (N_9396,N_553,N_1748);
xnor U9397 (N_9397,N_4309,N_4591);
or U9398 (N_9398,N_1860,N_6238);
xnor U9399 (N_9399,N_2298,N_2058);
and U9400 (N_9400,N_5267,N_5369);
nor U9401 (N_9401,N_2348,N_3392);
nand U9402 (N_9402,N_3892,N_4050);
xnor U9403 (N_9403,N_4390,N_1385);
xnor U9404 (N_9404,N_5993,N_3465);
nor U9405 (N_9405,N_1868,N_6086);
nand U9406 (N_9406,N_1303,N_2084);
nor U9407 (N_9407,N_3692,N_2171);
nor U9408 (N_9408,N_4242,N_6213);
nor U9409 (N_9409,N_602,N_187);
nor U9410 (N_9410,N_2518,N_6096);
nand U9411 (N_9411,N_3482,N_251);
or U9412 (N_9412,N_3380,N_2685);
and U9413 (N_9413,N_828,N_1399);
nor U9414 (N_9414,N_1990,N_1500);
xor U9415 (N_9415,N_2327,N_3061);
nor U9416 (N_9416,N_5838,N_553);
xnor U9417 (N_9417,N_838,N_5149);
nand U9418 (N_9418,N_1249,N_754);
and U9419 (N_9419,N_5380,N_4591);
xor U9420 (N_9420,N_5702,N_4632);
xnor U9421 (N_9421,N_2766,N_3275);
xnor U9422 (N_9422,N_2132,N_4845);
nor U9423 (N_9423,N_1716,N_3382);
nor U9424 (N_9424,N_4846,N_1161);
or U9425 (N_9425,N_855,N_3932);
xor U9426 (N_9426,N_579,N_666);
and U9427 (N_9427,N_2339,N_2387);
and U9428 (N_9428,N_1699,N_3444);
and U9429 (N_9429,N_5077,N_5290);
and U9430 (N_9430,N_4144,N_4978);
nand U9431 (N_9431,N_938,N_1809);
or U9432 (N_9432,N_1464,N_2982);
and U9433 (N_9433,N_1842,N_3074);
and U9434 (N_9434,N_1071,N_4447);
and U9435 (N_9435,N_3005,N_6131);
nor U9436 (N_9436,N_4014,N_4404);
and U9437 (N_9437,N_1573,N_6046);
nand U9438 (N_9438,N_3610,N_5776);
xnor U9439 (N_9439,N_3290,N_4485);
or U9440 (N_9440,N_2778,N_1970);
nand U9441 (N_9441,N_4799,N_4299);
nand U9442 (N_9442,N_6094,N_2828);
and U9443 (N_9443,N_3763,N_818);
or U9444 (N_9444,N_662,N_4308);
nor U9445 (N_9445,N_1080,N_3804);
or U9446 (N_9446,N_5012,N_1763);
nand U9447 (N_9447,N_5194,N_6190);
nor U9448 (N_9448,N_5050,N_5072);
nor U9449 (N_9449,N_585,N_1614);
xnor U9450 (N_9450,N_1003,N_4455);
xnor U9451 (N_9451,N_4658,N_3156);
and U9452 (N_9452,N_2195,N_1902);
xnor U9453 (N_9453,N_3712,N_4657);
and U9454 (N_9454,N_974,N_5629);
nand U9455 (N_9455,N_3429,N_3139);
nor U9456 (N_9456,N_1403,N_2275);
and U9457 (N_9457,N_1341,N_5420);
nand U9458 (N_9458,N_2906,N_1173);
nor U9459 (N_9459,N_5694,N_1683);
or U9460 (N_9460,N_5267,N_5853);
nand U9461 (N_9461,N_6208,N_2358);
or U9462 (N_9462,N_5833,N_5715);
nor U9463 (N_9463,N_5564,N_4323);
or U9464 (N_9464,N_1969,N_3751);
and U9465 (N_9465,N_606,N_4989);
and U9466 (N_9466,N_1679,N_934);
and U9467 (N_9467,N_1428,N_3067);
nand U9468 (N_9468,N_6228,N_3666);
nor U9469 (N_9469,N_2283,N_5909);
nor U9470 (N_9470,N_4375,N_2060);
nor U9471 (N_9471,N_2537,N_22);
and U9472 (N_9472,N_1421,N_4170);
nor U9473 (N_9473,N_3081,N_584);
or U9474 (N_9474,N_3852,N_4720);
xnor U9475 (N_9475,N_3483,N_751);
nand U9476 (N_9476,N_4573,N_2014);
nand U9477 (N_9477,N_1726,N_4649);
or U9478 (N_9478,N_3787,N_3430);
xor U9479 (N_9479,N_5097,N_4787);
or U9480 (N_9480,N_1161,N_4887);
nor U9481 (N_9481,N_1940,N_4448);
and U9482 (N_9482,N_4788,N_1018);
xor U9483 (N_9483,N_4123,N_3256);
xnor U9484 (N_9484,N_2913,N_3479);
and U9485 (N_9485,N_2259,N_3541);
nand U9486 (N_9486,N_1952,N_3939);
nand U9487 (N_9487,N_5708,N_827);
nor U9488 (N_9488,N_1501,N_1555);
nand U9489 (N_9489,N_1719,N_4225);
nand U9490 (N_9490,N_4569,N_6244);
nand U9491 (N_9491,N_850,N_4794);
xor U9492 (N_9492,N_3045,N_3006);
nand U9493 (N_9493,N_569,N_1704);
and U9494 (N_9494,N_5478,N_1621);
or U9495 (N_9495,N_2623,N_1055);
or U9496 (N_9496,N_6187,N_75);
nor U9497 (N_9497,N_2164,N_1747);
nor U9498 (N_9498,N_1127,N_1426);
and U9499 (N_9499,N_21,N_6016);
nand U9500 (N_9500,N_2971,N_5028);
and U9501 (N_9501,N_3781,N_3740);
nand U9502 (N_9502,N_5424,N_348);
nand U9503 (N_9503,N_5166,N_4198);
nand U9504 (N_9504,N_2295,N_3152);
xnor U9505 (N_9505,N_3126,N_1754);
nand U9506 (N_9506,N_5459,N_2683);
or U9507 (N_9507,N_5975,N_4567);
and U9508 (N_9508,N_1821,N_1336);
nor U9509 (N_9509,N_60,N_768);
or U9510 (N_9510,N_5267,N_1816);
xor U9511 (N_9511,N_5281,N_2219);
and U9512 (N_9512,N_1179,N_3181);
and U9513 (N_9513,N_5701,N_4436);
or U9514 (N_9514,N_4054,N_485);
nand U9515 (N_9515,N_2829,N_4842);
or U9516 (N_9516,N_266,N_4885);
xor U9517 (N_9517,N_4515,N_4517);
or U9518 (N_9518,N_3620,N_3400);
xor U9519 (N_9519,N_3114,N_3339);
or U9520 (N_9520,N_1518,N_1789);
and U9521 (N_9521,N_1751,N_985);
or U9522 (N_9522,N_1291,N_5242);
nor U9523 (N_9523,N_2263,N_373);
or U9524 (N_9524,N_3862,N_4028);
xor U9525 (N_9525,N_6206,N_5908);
and U9526 (N_9526,N_3451,N_826);
and U9527 (N_9527,N_6210,N_3700);
nand U9528 (N_9528,N_4647,N_2153);
nor U9529 (N_9529,N_1955,N_2340);
xnor U9530 (N_9530,N_1822,N_1268);
nor U9531 (N_9531,N_1511,N_5321);
and U9532 (N_9532,N_2057,N_5602);
nand U9533 (N_9533,N_4212,N_2026);
or U9534 (N_9534,N_831,N_5217);
or U9535 (N_9535,N_2164,N_5957);
xor U9536 (N_9536,N_159,N_1027);
or U9537 (N_9537,N_3279,N_2943);
nand U9538 (N_9538,N_2275,N_4303);
nand U9539 (N_9539,N_2828,N_4680);
or U9540 (N_9540,N_5240,N_5285);
xnor U9541 (N_9541,N_4772,N_5794);
or U9542 (N_9542,N_1343,N_354);
nand U9543 (N_9543,N_2974,N_1023);
and U9544 (N_9544,N_1306,N_2955);
xor U9545 (N_9545,N_5513,N_6009);
nor U9546 (N_9546,N_924,N_2840);
nand U9547 (N_9547,N_2536,N_2045);
nor U9548 (N_9548,N_1603,N_1753);
xnor U9549 (N_9549,N_3759,N_1204);
or U9550 (N_9550,N_3304,N_5034);
xnor U9551 (N_9551,N_414,N_1162);
and U9552 (N_9552,N_1894,N_3740);
or U9553 (N_9553,N_4158,N_4859);
and U9554 (N_9554,N_573,N_3717);
or U9555 (N_9555,N_142,N_4323);
xnor U9556 (N_9556,N_5200,N_4451);
xnor U9557 (N_9557,N_1533,N_1783);
or U9558 (N_9558,N_4298,N_3393);
nor U9559 (N_9559,N_4376,N_2950);
and U9560 (N_9560,N_5369,N_923);
xnor U9561 (N_9561,N_4540,N_3092);
xor U9562 (N_9562,N_1959,N_4912);
xor U9563 (N_9563,N_2834,N_14);
nor U9564 (N_9564,N_3233,N_482);
nor U9565 (N_9565,N_4689,N_3594);
and U9566 (N_9566,N_6188,N_4158);
nor U9567 (N_9567,N_1812,N_4220);
nor U9568 (N_9568,N_2282,N_6125);
xor U9569 (N_9569,N_3886,N_3688);
or U9570 (N_9570,N_3773,N_1937);
nor U9571 (N_9571,N_5970,N_4223);
or U9572 (N_9572,N_5981,N_3147);
nand U9573 (N_9573,N_4485,N_564);
nor U9574 (N_9574,N_625,N_4668);
nand U9575 (N_9575,N_1580,N_6115);
and U9576 (N_9576,N_3389,N_3176);
xor U9577 (N_9577,N_3315,N_2222);
nand U9578 (N_9578,N_3279,N_4055);
nand U9579 (N_9579,N_2131,N_1223);
xnor U9580 (N_9580,N_4990,N_4423);
xor U9581 (N_9581,N_2274,N_5799);
nand U9582 (N_9582,N_2988,N_6094);
nor U9583 (N_9583,N_1262,N_5306);
or U9584 (N_9584,N_2347,N_1263);
or U9585 (N_9585,N_3814,N_2637);
xnor U9586 (N_9586,N_3826,N_3687);
or U9587 (N_9587,N_5158,N_3767);
nand U9588 (N_9588,N_4222,N_867);
and U9589 (N_9589,N_4633,N_17);
xor U9590 (N_9590,N_1746,N_1312);
and U9591 (N_9591,N_5435,N_4618);
nor U9592 (N_9592,N_2884,N_501);
nand U9593 (N_9593,N_2745,N_1439);
and U9594 (N_9594,N_5901,N_6177);
nand U9595 (N_9595,N_243,N_1329);
nor U9596 (N_9596,N_5597,N_2944);
nor U9597 (N_9597,N_2931,N_1765);
or U9598 (N_9598,N_3664,N_1490);
xnor U9599 (N_9599,N_5495,N_1367);
and U9600 (N_9600,N_2519,N_5978);
xor U9601 (N_9601,N_134,N_6248);
and U9602 (N_9602,N_2008,N_4762);
nand U9603 (N_9603,N_3589,N_4903);
xnor U9604 (N_9604,N_3168,N_4900);
nor U9605 (N_9605,N_1829,N_2637);
nor U9606 (N_9606,N_3646,N_1949);
or U9607 (N_9607,N_3723,N_528);
or U9608 (N_9608,N_911,N_2044);
nor U9609 (N_9609,N_835,N_2194);
xor U9610 (N_9610,N_4108,N_4167);
xnor U9611 (N_9611,N_4681,N_3661);
nand U9612 (N_9612,N_639,N_5089);
and U9613 (N_9613,N_2016,N_742);
or U9614 (N_9614,N_4623,N_1036);
nor U9615 (N_9615,N_1152,N_1609);
nand U9616 (N_9616,N_5699,N_597);
or U9617 (N_9617,N_5889,N_1782);
or U9618 (N_9618,N_5228,N_2555);
nand U9619 (N_9619,N_1809,N_5861);
and U9620 (N_9620,N_385,N_2387);
xnor U9621 (N_9621,N_6196,N_3489);
nand U9622 (N_9622,N_5902,N_4046);
and U9623 (N_9623,N_3565,N_2975);
nor U9624 (N_9624,N_4619,N_4809);
and U9625 (N_9625,N_1527,N_5377);
nor U9626 (N_9626,N_199,N_5666);
and U9627 (N_9627,N_1714,N_2875);
xor U9628 (N_9628,N_4679,N_5011);
nor U9629 (N_9629,N_5546,N_41);
nand U9630 (N_9630,N_4201,N_5508);
xor U9631 (N_9631,N_1096,N_3860);
and U9632 (N_9632,N_2781,N_5885);
or U9633 (N_9633,N_5596,N_5736);
and U9634 (N_9634,N_5678,N_1999);
nor U9635 (N_9635,N_650,N_3041);
xnor U9636 (N_9636,N_4761,N_3249);
and U9637 (N_9637,N_5707,N_5759);
nand U9638 (N_9638,N_512,N_3068);
nand U9639 (N_9639,N_399,N_4026);
and U9640 (N_9640,N_4234,N_4500);
and U9641 (N_9641,N_2078,N_5510);
nand U9642 (N_9642,N_1518,N_2171);
or U9643 (N_9643,N_5031,N_4245);
xor U9644 (N_9644,N_434,N_3416);
or U9645 (N_9645,N_1462,N_5841);
nand U9646 (N_9646,N_5122,N_411);
and U9647 (N_9647,N_2596,N_2017);
and U9648 (N_9648,N_3719,N_5788);
nand U9649 (N_9649,N_4381,N_6169);
and U9650 (N_9650,N_2075,N_2673);
or U9651 (N_9651,N_2780,N_1397);
and U9652 (N_9652,N_1781,N_5209);
nand U9653 (N_9653,N_3560,N_1449);
or U9654 (N_9654,N_132,N_2097);
nand U9655 (N_9655,N_3518,N_3388);
nand U9656 (N_9656,N_1746,N_656);
or U9657 (N_9657,N_2402,N_4237);
nor U9658 (N_9658,N_5045,N_6243);
and U9659 (N_9659,N_4904,N_3785);
nand U9660 (N_9660,N_4692,N_2576);
xnor U9661 (N_9661,N_3969,N_2076);
or U9662 (N_9662,N_2846,N_898);
and U9663 (N_9663,N_186,N_1854);
nor U9664 (N_9664,N_4258,N_1179);
or U9665 (N_9665,N_1948,N_2450);
or U9666 (N_9666,N_5681,N_1243);
nor U9667 (N_9667,N_5885,N_1200);
nand U9668 (N_9668,N_3589,N_345);
nor U9669 (N_9669,N_4968,N_5370);
and U9670 (N_9670,N_3416,N_3261);
xor U9671 (N_9671,N_5083,N_420);
and U9672 (N_9672,N_6004,N_3963);
nor U9673 (N_9673,N_2852,N_2860);
and U9674 (N_9674,N_5292,N_350);
nor U9675 (N_9675,N_3383,N_4660);
and U9676 (N_9676,N_1177,N_1167);
xnor U9677 (N_9677,N_5644,N_3203);
xnor U9678 (N_9678,N_1193,N_2666);
xor U9679 (N_9679,N_3374,N_5712);
xnor U9680 (N_9680,N_6051,N_2725);
nor U9681 (N_9681,N_4127,N_3787);
or U9682 (N_9682,N_805,N_4);
nand U9683 (N_9683,N_2838,N_4281);
xnor U9684 (N_9684,N_1829,N_4164);
nor U9685 (N_9685,N_4120,N_4646);
xnor U9686 (N_9686,N_1010,N_4424);
or U9687 (N_9687,N_1836,N_5317);
or U9688 (N_9688,N_5313,N_347);
nand U9689 (N_9689,N_996,N_1592);
or U9690 (N_9690,N_4353,N_4146);
nand U9691 (N_9691,N_1479,N_3147);
and U9692 (N_9692,N_5752,N_2758);
xnor U9693 (N_9693,N_5778,N_905);
xor U9694 (N_9694,N_2940,N_4925);
or U9695 (N_9695,N_2975,N_2730);
and U9696 (N_9696,N_725,N_4925);
nor U9697 (N_9697,N_3162,N_975);
xnor U9698 (N_9698,N_5932,N_832);
and U9699 (N_9699,N_1851,N_5789);
or U9700 (N_9700,N_614,N_4176);
nand U9701 (N_9701,N_319,N_1912);
xor U9702 (N_9702,N_4313,N_6028);
and U9703 (N_9703,N_1790,N_4964);
or U9704 (N_9704,N_2712,N_2424);
and U9705 (N_9705,N_5257,N_2045);
nor U9706 (N_9706,N_4742,N_5553);
or U9707 (N_9707,N_766,N_4082);
nor U9708 (N_9708,N_3778,N_1911);
xnor U9709 (N_9709,N_3953,N_1739);
nand U9710 (N_9710,N_3730,N_3250);
nand U9711 (N_9711,N_312,N_647);
and U9712 (N_9712,N_4141,N_3367);
and U9713 (N_9713,N_3167,N_580);
xnor U9714 (N_9714,N_5164,N_2221);
or U9715 (N_9715,N_4729,N_1026);
nand U9716 (N_9716,N_4529,N_628);
nor U9717 (N_9717,N_205,N_4652);
nor U9718 (N_9718,N_6123,N_3336);
nor U9719 (N_9719,N_1229,N_5851);
nand U9720 (N_9720,N_5293,N_5203);
xor U9721 (N_9721,N_627,N_3983);
nand U9722 (N_9722,N_478,N_3674);
xor U9723 (N_9723,N_2985,N_1002);
nor U9724 (N_9724,N_5092,N_4296);
xnor U9725 (N_9725,N_3456,N_4515);
xor U9726 (N_9726,N_4512,N_1312);
and U9727 (N_9727,N_5652,N_1524);
nand U9728 (N_9728,N_2355,N_5051);
nor U9729 (N_9729,N_2583,N_2788);
xnor U9730 (N_9730,N_5935,N_4090);
or U9731 (N_9731,N_2628,N_6138);
or U9732 (N_9732,N_5440,N_62);
nor U9733 (N_9733,N_2462,N_4417);
nand U9734 (N_9734,N_3462,N_4852);
and U9735 (N_9735,N_2619,N_2836);
nand U9736 (N_9736,N_2825,N_2593);
or U9737 (N_9737,N_2180,N_2944);
or U9738 (N_9738,N_4375,N_1049);
nand U9739 (N_9739,N_5258,N_3379);
nand U9740 (N_9740,N_4570,N_5378);
or U9741 (N_9741,N_5687,N_1080);
nor U9742 (N_9742,N_5310,N_3390);
nand U9743 (N_9743,N_4906,N_2468);
nor U9744 (N_9744,N_2092,N_4347);
or U9745 (N_9745,N_3079,N_1387);
nand U9746 (N_9746,N_5133,N_5247);
nor U9747 (N_9747,N_2403,N_4289);
nor U9748 (N_9748,N_2468,N_192);
nand U9749 (N_9749,N_6014,N_4280);
nor U9750 (N_9750,N_2575,N_1163);
nand U9751 (N_9751,N_3020,N_3310);
or U9752 (N_9752,N_2144,N_2188);
xnor U9753 (N_9753,N_2661,N_4162);
or U9754 (N_9754,N_4932,N_1321);
xnor U9755 (N_9755,N_5536,N_1078);
and U9756 (N_9756,N_2050,N_423);
nand U9757 (N_9757,N_5559,N_5963);
nand U9758 (N_9758,N_2548,N_5178);
xnor U9759 (N_9759,N_1414,N_3221);
nand U9760 (N_9760,N_530,N_13);
and U9761 (N_9761,N_4198,N_5587);
nand U9762 (N_9762,N_1592,N_3251);
xnor U9763 (N_9763,N_839,N_3737);
nand U9764 (N_9764,N_5646,N_1658);
and U9765 (N_9765,N_3343,N_2904);
or U9766 (N_9766,N_1794,N_3391);
nor U9767 (N_9767,N_818,N_686);
nor U9768 (N_9768,N_4075,N_3876);
nor U9769 (N_9769,N_2191,N_5230);
xor U9770 (N_9770,N_567,N_4805);
and U9771 (N_9771,N_1483,N_3871);
nor U9772 (N_9772,N_2292,N_3582);
nor U9773 (N_9773,N_1212,N_3150);
and U9774 (N_9774,N_498,N_2330);
and U9775 (N_9775,N_3563,N_1678);
or U9776 (N_9776,N_5109,N_3440);
and U9777 (N_9777,N_2524,N_1592);
nand U9778 (N_9778,N_107,N_3944);
xnor U9779 (N_9779,N_1276,N_1144);
or U9780 (N_9780,N_3035,N_4729);
and U9781 (N_9781,N_4738,N_2477);
xnor U9782 (N_9782,N_1819,N_1368);
xor U9783 (N_9783,N_694,N_4957);
nor U9784 (N_9784,N_4776,N_2032);
or U9785 (N_9785,N_1574,N_3999);
or U9786 (N_9786,N_1571,N_917);
nor U9787 (N_9787,N_2427,N_781);
or U9788 (N_9788,N_5852,N_1959);
nand U9789 (N_9789,N_1052,N_1419);
and U9790 (N_9790,N_5380,N_3866);
or U9791 (N_9791,N_5101,N_2784);
nand U9792 (N_9792,N_371,N_1594);
xor U9793 (N_9793,N_5504,N_1337);
and U9794 (N_9794,N_1574,N_3184);
xnor U9795 (N_9795,N_4041,N_6021);
or U9796 (N_9796,N_5434,N_644);
or U9797 (N_9797,N_6088,N_4871);
nor U9798 (N_9798,N_1435,N_5824);
nor U9799 (N_9799,N_3608,N_1355);
or U9800 (N_9800,N_2518,N_283);
or U9801 (N_9801,N_3374,N_2037);
xnor U9802 (N_9802,N_902,N_5887);
nor U9803 (N_9803,N_1693,N_1077);
xor U9804 (N_9804,N_2868,N_603);
or U9805 (N_9805,N_1563,N_1859);
nand U9806 (N_9806,N_5589,N_3837);
nor U9807 (N_9807,N_4001,N_4473);
nand U9808 (N_9808,N_1132,N_5667);
and U9809 (N_9809,N_3786,N_4682);
or U9810 (N_9810,N_3042,N_4428);
nand U9811 (N_9811,N_5921,N_6124);
or U9812 (N_9812,N_363,N_2439);
or U9813 (N_9813,N_776,N_87);
nand U9814 (N_9814,N_6077,N_5058);
nor U9815 (N_9815,N_3310,N_391);
or U9816 (N_9816,N_4240,N_5985);
xor U9817 (N_9817,N_2220,N_5693);
nand U9818 (N_9818,N_4508,N_174);
nand U9819 (N_9819,N_4460,N_4726);
and U9820 (N_9820,N_2611,N_2305);
nor U9821 (N_9821,N_2099,N_5710);
xnor U9822 (N_9822,N_1544,N_541);
nand U9823 (N_9823,N_676,N_5151);
and U9824 (N_9824,N_3905,N_5478);
nand U9825 (N_9825,N_725,N_1791);
and U9826 (N_9826,N_6022,N_3210);
or U9827 (N_9827,N_1051,N_3008);
xor U9828 (N_9828,N_1848,N_6237);
and U9829 (N_9829,N_1721,N_1204);
xor U9830 (N_9830,N_1706,N_222);
and U9831 (N_9831,N_251,N_36);
and U9832 (N_9832,N_3439,N_4335);
or U9833 (N_9833,N_1298,N_2153);
and U9834 (N_9834,N_1568,N_2153);
and U9835 (N_9835,N_2974,N_2370);
and U9836 (N_9836,N_5376,N_1672);
or U9837 (N_9837,N_3128,N_5456);
xnor U9838 (N_9838,N_1789,N_2979);
nor U9839 (N_9839,N_4518,N_5272);
nand U9840 (N_9840,N_5808,N_4609);
nand U9841 (N_9841,N_4532,N_5208);
or U9842 (N_9842,N_144,N_348);
or U9843 (N_9843,N_2262,N_4973);
nor U9844 (N_9844,N_4147,N_1690);
or U9845 (N_9845,N_1698,N_2848);
xor U9846 (N_9846,N_4148,N_2707);
and U9847 (N_9847,N_4985,N_1125);
nand U9848 (N_9848,N_2330,N_5734);
nand U9849 (N_9849,N_5571,N_2825);
nor U9850 (N_9850,N_6157,N_687);
nor U9851 (N_9851,N_6058,N_2049);
nor U9852 (N_9852,N_4894,N_1797);
nor U9853 (N_9853,N_4712,N_5607);
nand U9854 (N_9854,N_2876,N_2240);
or U9855 (N_9855,N_858,N_2058);
nor U9856 (N_9856,N_3252,N_560);
or U9857 (N_9857,N_4634,N_2199);
or U9858 (N_9858,N_313,N_2218);
nor U9859 (N_9859,N_3374,N_2036);
and U9860 (N_9860,N_2395,N_2433);
nand U9861 (N_9861,N_1501,N_5697);
and U9862 (N_9862,N_1262,N_5180);
or U9863 (N_9863,N_4510,N_5259);
nand U9864 (N_9864,N_1480,N_1329);
xnor U9865 (N_9865,N_1198,N_772);
or U9866 (N_9866,N_2489,N_3074);
nor U9867 (N_9867,N_1574,N_2516);
xnor U9868 (N_9868,N_1054,N_1296);
and U9869 (N_9869,N_3416,N_4223);
and U9870 (N_9870,N_5525,N_3968);
nor U9871 (N_9871,N_3237,N_1477);
nand U9872 (N_9872,N_1531,N_1994);
nand U9873 (N_9873,N_3900,N_3082);
nand U9874 (N_9874,N_3519,N_4411);
and U9875 (N_9875,N_548,N_3120);
and U9876 (N_9876,N_6108,N_5140);
xor U9877 (N_9877,N_3702,N_5504);
nand U9878 (N_9878,N_5226,N_5486);
or U9879 (N_9879,N_5545,N_4960);
or U9880 (N_9880,N_4399,N_1933);
and U9881 (N_9881,N_3163,N_3565);
xor U9882 (N_9882,N_3615,N_882);
or U9883 (N_9883,N_2596,N_198);
and U9884 (N_9884,N_3622,N_3880);
and U9885 (N_9885,N_4667,N_1747);
xor U9886 (N_9886,N_1669,N_2956);
nand U9887 (N_9887,N_754,N_5201);
and U9888 (N_9888,N_1760,N_6196);
xnor U9889 (N_9889,N_4627,N_4483);
xnor U9890 (N_9890,N_2787,N_4754);
xor U9891 (N_9891,N_1925,N_16);
nand U9892 (N_9892,N_583,N_4247);
or U9893 (N_9893,N_6084,N_336);
nor U9894 (N_9894,N_4312,N_1787);
nor U9895 (N_9895,N_4698,N_401);
xnor U9896 (N_9896,N_1780,N_1446);
or U9897 (N_9897,N_6191,N_3537);
xor U9898 (N_9898,N_386,N_1247);
and U9899 (N_9899,N_5150,N_3438);
xor U9900 (N_9900,N_4346,N_2480);
nor U9901 (N_9901,N_2414,N_1276);
xnor U9902 (N_9902,N_2216,N_4763);
and U9903 (N_9903,N_4165,N_2766);
nand U9904 (N_9904,N_1149,N_5291);
xnor U9905 (N_9905,N_4741,N_145);
nand U9906 (N_9906,N_3354,N_5956);
and U9907 (N_9907,N_5152,N_6030);
and U9908 (N_9908,N_5883,N_957);
and U9909 (N_9909,N_1836,N_5225);
nor U9910 (N_9910,N_2350,N_1816);
nand U9911 (N_9911,N_423,N_178);
xnor U9912 (N_9912,N_2270,N_3288);
xor U9913 (N_9913,N_1465,N_5376);
nor U9914 (N_9914,N_913,N_827);
or U9915 (N_9915,N_163,N_3911);
nor U9916 (N_9916,N_6209,N_932);
xor U9917 (N_9917,N_5755,N_117);
nor U9918 (N_9918,N_4274,N_3115);
and U9919 (N_9919,N_1499,N_1870);
or U9920 (N_9920,N_6195,N_3651);
nand U9921 (N_9921,N_3479,N_2906);
or U9922 (N_9922,N_5739,N_1407);
xor U9923 (N_9923,N_3548,N_1411);
or U9924 (N_9924,N_4410,N_5297);
and U9925 (N_9925,N_141,N_4954);
xnor U9926 (N_9926,N_5996,N_2787);
xor U9927 (N_9927,N_2271,N_3723);
xor U9928 (N_9928,N_3638,N_1294);
nor U9929 (N_9929,N_3702,N_2097);
xnor U9930 (N_9930,N_610,N_1882);
xor U9931 (N_9931,N_379,N_6214);
or U9932 (N_9932,N_5876,N_2653);
xnor U9933 (N_9933,N_5893,N_2020);
nand U9934 (N_9934,N_2082,N_4504);
xor U9935 (N_9935,N_2012,N_132);
or U9936 (N_9936,N_3604,N_1882);
xnor U9937 (N_9937,N_109,N_3980);
and U9938 (N_9938,N_517,N_6199);
nand U9939 (N_9939,N_4876,N_975);
nor U9940 (N_9940,N_4955,N_2613);
nand U9941 (N_9941,N_4864,N_5999);
and U9942 (N_9942,N_989,N_1247);
xor U9943 (N_9943,N_4402,N_6191);
or U9944 (N_9944,N_5948,N_5957);
and U9945 (N_9945,N_4487,N_2720);
xnor U9946 (N_9946,N_5508,N_5205);
or U9947 (N_9947,N_1504,N_2748);
nor U9948 (N_9948,N_5197,N_1878);
xnor U9949 (N_9949,N_6195,N_4131);
nor U9950 (N_9950,N_2250,N_5930);
nor U9951 (N_9951,N_377,N_5201);
or U9952 (N_9952,N_3762,N_3039);
or U9953 (N_9953,N_1384,N_6080);
nand U9954 (N_9954,N_3587,N_5711);
or U9955 (N_9955,N_2025,N_5412);
and U9956 (N_9956,N_3999,N_2714);
or U9957 (N_9957,N_46,N_6027);
nand U9958 (N_9958,N_1235,N_4600);
or U9959 (N_9959,N_3759,N_4036);
nand U9960 (N_9960,N_152,N_5674);
nor U9961 (N_9961,N_268,N_177);
nor U9962 (N_9962,N_4910,N_2905);
xnor U9963 (N_9963,N_1803,N_2670);
xor U9964 (N_9964,N_197,N_3813);
nand U9965 (N_9965,N_812,N_2301);
or U9966 (N_9966,N_4990,N_2671);
or U9967 (N_9967,N_3911,N_4397);
and U9968 (N_9968,N_201,N_6039);
xor U9969 (N_9969,N_715,N_2792);
xnor U9970 (N_9970,N_2962,N_0);
or U9971 (N_9971,N_3895,N_2010);
and U9972 (N_9972,N_2503,N_2954);
or U9973 (N_9973,N_6115,N_1942);
nand U9974 (N_9974,N_3504,N_3189);
xnor U9975 (N_9975,N_2133,N_3697);
nand U9976 (N_9976,N_1262,N_3462);
or U9977 (N_9977,N_3008,N_267);
or U9978 (N_9978,N_1148,N_2198);
xor U9979 (N_9979,N_4768,N_4418);
nand U9980 (N_9980,N_1547,N_5311);
xor U9981 (N_9981,N_2117,N_2055);
xor U9982 (N_9982,N_4226,N_597);
nand U9983 (N_9983,N_2151,N_5634);
xor U9984 (N_9984,N_359,N_4662);
xor U9985 (N_9985,N_5572,N_674);
or U9986 (N_9986,N_1073,N_4630);
xor U9987 (N_9987,N_1864,N_1418);
nand U9988 (N_9988,N_2226,N_3101);
xor U9989 (N_9989,N_3304,N_5124);
or U9990 (N_9990,N_264,N_1064);
and U9991 (N_9991,N_1643,N_2588);
xnor U9992 (N_9992,N_996,N_2185);
and U9993 (N_9993,N_4769,N_1122);
xor U9994 (N_9994,N_675,N_4550);
xnor U9995 (N_9995,N_2639,N_3394);
xnor U9996 (N_9996,N_2076,N_1645);
nand U9997 (N_9997,N_5853,N_1074);
and U9998 (N_9998,N_2531,N_5527);
nand U9999 (N_9999,N_4213,N_4);
or U10000 (N_10000,N_3753,N_5565);
or U10001 (N_10001,N_3159,N_5966);
xor U10002 (N_10002,N_1464,N_1226);
and U10003 (N_10003,N_2751,N_5272);
and U10004 (N_10004,N_408,N_312);
xor U10005 (N_10005,N_4109,N_5343);
xor U10006 (N_10006,N_4716,N_262);
nor U10007 (N_10007,N_1439,N_3221);
xor U10008 (N_10008,N_3812,N_2550);
nand U10009 (N_10009,N_3860,N_849);
xnor U10010 (N_10010,N_930,N_734);
and U10011 (N_10011,N_3913,N_2594);
nand U10012 (N_10012,N_3871,N_5226);
or U10013 (N_10013,N_630,N_2368);
nand U10014 (N_10014,N_3677,N_4730);
nand U10015 (N_10015,N_2628,N_578);
nor U10016 (N_10016,N_5244,N_3265);
or U10017 (N_10017,N_1354,N_4482);
nor U10018 (N_10018,N_2399,N_5596);
or U10019 (N_10019,N_4159,N_978);
nor U10020 (N_10020,N_4586,N_1687);
and U10021 (N_10021,N_5910,N_1482);
nand U10022 (N_10022,N_1983,N_4872);
nand U10023 (N_10023,N_1435,N_3458);
nor U10024 (N_10024,N_1611,N_3000);
nand U10025 (N_10025,N_265,N_567);
and U10026 (N_10026,N_4461,N_1223);
and U10027 (N_10027,N_3580,N_1819);
nor U10028 (N_10028,N_4084,N_4088);
or U10029 (N_10029,N_5448,N_4021);
nor U10030 (N_10030,N_1949,N_3740);
nand U10031 (N_10031,N_2856,N_355);
nand U10032 (N_10032,N_493,N_3611);
or U10033 (N_10033,N_3373,N_1494);
nand U10034 (N_10034,N_5393,N_1921);
and U10035 (N_10035,N_4955,N_1062);
nand U10036 (N_10036,N_4578,N_644);
nand U10037 (N_10037,N_2880,N_3178);
and U10038 (N_10038,N_6217,N_5681);
and U10039 (N_10039,N_597,N_4700);
or U10040 (N_10040,N_2072,N_6202);
nor U10041 (N_10041,N_951,N_5541);
xnor U10042 (N_10042,N_589,N_6007);
nor U10043 (N_10043,N_384,N_1837);
nand U10044 (N_10044,N_5531,N_3924);
nand U10045 (N_10045,N_3205,N_3798);
nor U10046 (N_10046,N_3398,N_4593);
and U10047 (N_10047,N_1531,N_1981);
nor U10048 (N_10048,N_2532,N_1564);
xor U10049 (N_10049,N_3105,N_1101);
nor U10050 (N_10050,N_5678,N_707);
xnor U10051 (N_10051,N_3881,N_6126);
nor U10052 (N_10052,N_1552,N_1786);
xor U10053 (N_10053,N_6165,N_2233);
nand U10054 (N_10054,N_141,N_5639);
nand U10055 (N_10055,N_2515,N_5708);
or U10056 (N_10056,N_7,N_4821);
and U10057 (N_10057,N_2306,N_4371);
or U10058 (N_10058,N_5057,N_4900);
or U10059 (N_10059,N_5061,N_3516);
and U10060 (N_10060,N_4340,N_4685);
xnor U10061 (N_10061,N_3208,N_1890);
or U10062 (N_10062,N_5119,N_4774);
nor U10063 (N_10063,N_3325,N_1453);
and U10064 (N_10064,N_6109,N_528);
or U10065 (N_10065,N_3039,N_3208);
nor U10066 (N_10066,N_3289,N_3890);
nor U10067 (N_10067,N_4063,N_2080);
nand U10068 (N_10068,N_5632,N_550);
nand U10069 (N_10069,N_1536,N_2435);
nor U10070 (N_10070,N_4989,N_1481);
nor U10071 (N_10071,N_2233,N_4936);
nor U10072 (N_10072,N_6142,N_3838);
nand U10073 (N_10073,N_4335,N_5881);
and U10074 (N_10074,N_295,N_3462);
xnor U10075 (N_10075,N_5671,N_2980);
xor U10076 (N_10076,N_927,N_3010);
nor U10077 (N_10077,N_5148,N_1190);
xnor U10078 (N_10078,N_6013,N_5729);
and U10079 (N_10079,N_5831,N_837);
nand U10080 (N_10080,N_2982,N_2129);
and U10081 (N_10081,N_699,N_4759);
nor U10082 (N_10082,N_2037,N_4093);
and U10083 (N_10083,N_1829,N_3510);
nand U10084 (N_10084,N_5136,N_6207);
and U10085 (N_10085,N_4157,N_4180);
nor U10086 (N_10086,N_1852,N_4684);
nor U10087 (N_10087,N_3629,N_6069);
and U10088 (N_10088,N_5447,N_4503);
or U10089 (N_10089,N_2014,N_6114);
and U10090 (N_10090,N_5671,N_1726);
xnor U10091 (N_10091,N_5243,N_4213);
xnor U10092 (N_10092,N_2891,N_2401);
or U10093 (N_10093,N_3595,N_2144);
and U10094 (N_10094,N_4448,N_87);
nand U10095 (N_10095,N_621,N_971);
or U10096 (N_10096,N_508,N_497);
or U10097 (N_10097,N_4135,N_5553);
nand U10098 (N_10098,N_629,N_4091);
nor U10099 (N_10099,N_1930,N_5697);
nor U10100 (N_10100,N_1525,N_3099);
or U10101 (N_10101,N_4168,N_6172);
or U10102 (N_10102,N_2359,N_2222);
nor U10103 (N_10103,N_5859,N_224);
or U10104 (N_10104,N_5614,N_3518);
nand U10105 (N_10105,N_1533,N_4930);
nor U10106 (N_10106,N_1224,N_864);
xor U10107 (N_10107,N_1875,N_240);
xor U10108 (N_10108,N_4302,N_4503);
xnor U10109 (N_10109,N_5661,N_6023);
xor U10110 (N_10110,N_3412,N_5056);
nand U10111 (N_10111,N_6220,N_846);
xor U10112 (N_10112,N_5742,N_2975);
nand U10113 (N_10113,N_2633,N_319);
xor U10114 (N_10114,N_5688,N_4974);
or U10115 (N_10115,N_455,N_5837);
nand U10116 (N_10116,N_5138,N_3792);
or U10117 (N_10117,N_2262,N_4204);
nor U10118 (N_10118,N_5828,N_2643);
and U10119 (N_10119,N_400,N_1015);
nor U10120 (N_10120,N_5694,N_2554);
or U10121 (N_10121,N_2784,N_2730);
xor U10122 (N_10122,N_417,N_2704);
nor U10123 (N_10123,N_5550,N_4875);
xnor U10124 (N_10124,N_4900,N_447);
and U10125 (N_10125,N_1868,N_3568);
nor U10126 (N_10126,N_5996,N_4320);
and U10127 (N_10127,N_4200,N_2639);
nand U10128 (N_10128,N_783,N_4084);
xnor U10129 (N_10129,N_3857,N_5046);
nor U10130 (N_10130,N_2540,N_1772);
nor U10131 (N_10131,N_751,N_5013);
nand U10132 (N_10132,N_4398,N_2381);
xor U10133 (N_10133,N_3574,N_2275);
and U10134 (N_10134,N_3602,N_3378);
nor U10135 (N_10135,N_3569,N_5371);
xnor U10136 (N_10136,N_4006,N_679);
nand U10137 (N_10137,N_887,N_4912);
nor U10138 (N_10138,N_3179,N_5822);
or U10139 (N_10139,N_2017,N_2963);
and U10140 (N_10140,N_6105,N_1562);
xnor U10141 (N_10141,N_303,N_1191);
or U10142 (N_10142,N_5707,N_5296);
nor U10143 (N_10143,N_5878,N_2437);
xnor U10144 (N_10144,N_759,N_4564);
nand U10145 (N_10145,N_4317,N_3322);
nor U10146 (N_10146,N_5585,N_4623);
and U10147 (N_10147,N_3580,N_6115);
or U10148 (N_10148,N_621,N_2802);
or U10149 (N_10149,N_3266,N_5416);
xnor U10150 (N_10150,N_2903,N_5203);
nor U10151 (N_10151,N_2808,N_1878);
and U10152 (N_10152,N_2188,N_2100);
or U10153 (N_10153,N_3462,N_6227);
nand U10154 (N_10154,N_2695,N_6205);
or U10155 (N_10155,N_1320,N_4956);
nor U10156 (N_10156,N_221,N_1249);
xnor U10157 (N_10157,N_5686,N_2811);
or U10158 (N_10158,N_625,N_5258);
nor U10159 (N_10159,N_2394,N_966);
nand U10160 (N_10160,N_5197,N_724);
or U10161 (N_10161,N_3683,N_1396);
or U10162 (N_10162,N_5420,N_2642);
nor U10163 (N_10163,N_4189,N_5534);
or U10164 (N_10164,N_142,N_2044);
nand U10165 (N_10165,N_837,N_5817);
or U10166 (N_10166,N_3522,N_2160);
nor U10167 (N_10167,N_3312,N_5590);
and U10168 (N_10168,N_2519,N_5148);
nor U10169 (N_10169,N_2841,N_556);
and U10170 (N_10170,N_5256,N_486);
xor U10171 (N_10171,N_2285,N_4255);
nand U10172 (N_10172,N_2619,N_4342);
nand U10173 (N_10173,N_5037,N_5086);
nand U10174 (N_10174,N_700,N_63);
nor U10175 (N_10175,N_4958,N_3723);
xnor U10176 (N_10176,N_3854,N_4284);
and U10177 (N_10177,N_4635,N_4950);
or U10178 (N_10178,N_2428,N_1015);
and U10179 (N_10179,N_5564,N_2662);
nand U10180 (N_10180,N_677,N_519);
and U10181 (N_10181,N_4733,N_4187);
xor U10182 (N_10182,N_5907,N_3464);
xnor U10183 (N_10183,N_2066,N_5396);
nand U10184 (N_10184,N_4245,N_2731);
or U10185 (N_10185,N_139,N_1206);
or U10186 (N_10186,N_6008,N_6081);
nand U10187 (N_10187,N_1279,N_6224);
xor U10188 (N_10188,N_1782,N_3159);
xnor U10189 (N_10189,N_2855,N_2651);
or U10190 (N_10190,N_5272,N_830);
or U10191 (N_10191,N_4227,N_31);
xnor U10192 (N_10192,N_2031,N_3272);
nor U10193 (N_10193,N_400,N_2550);
nor U10194 (N_10194,N_5961,N_1804);
or U10195 (N_10195,N_3056,N_2709);
and U10196 (N_10196,N_6127,N_870);
nand U10197 (N_10197,N_872,N_830);
or U10198 (N_10198,N_3927,N_5816);
xor U10199 (N_10199,N_795,N_4364);
or U10200 (N_10200,N_5257,N_4270);
nand U10201 (N_10201,N_5458,N_5942);
nand U10202 (N_10202,N_2743,N_5824);
and U10203 (N_10203,N_6117,N_2318);
or U10204 (N_10204,N_4424,N_5454);
nand U10205 (N_10205,N_159,N_4447);
nand U10206 (N_10206,N_4390,N_4250);
nand U10207 (N_10207,N_1867,N_6191);
nand U10208 (N_10208,N_2349,N_5781);
nand U10209 (N_10209,N_32,N_1568);
nand U10210 (N_10210,N_3259,N_4289);
or U10211 (N_10211,N_4265,N_1168);
nor U10212 (N_10212,N_5360,N_2030);
nand U10213 (N_10213,N_6123,N_5781);
or U10214 (N_10214,N_5257,N_2988);
or U10215 (N_10215,N_2797,N_5125);
nand U10216 (N_10216,N_4490,N_1769);
and U10217 (N_10217,N_482,N_6054);
nor U10218 (N_10218,N_2474,N_5542);
or U10219 (N_10219,N_4566,N_5933);
and U10220 (N_10220,N_636,N_3738);
and U10221 (N_10221,N_1439,N_4735);
nand U10222 (N_10222,N_123,N_2276);
xnor U10223 (N_10223,N_388,N_215);
and U10224 (N_10224,N_2636,N_528);
nand U10225 (N_10225,N_1581,N_5127);
and U10226 (N_10226,N_4450,N_4131);
and U10227 (N_10227,N_3436,N_6230);
and U10228 (N_10228,N_3694,N_884);
and U10229 (N_10229,N_3224,N_3017);
nor U10230 (N_10230,N_2481,N_4528);
or U10231 (N_10231,N_4293,N_6040);
xor U10232 (N_10232,N_4530,N_1764);
and U10233 (N_10233,N_324,N_2634);
nor U10234 (N_10234,N_3770,N_3815);
nor U10235 (N_10235,N_1626,N_2404);
and U10236 (N_10236,N_1865,N_1267);
nand U10237 (N_10237,N_3910,N_2781);
xnor U10238 (N_10238,N_3945,N_5409);
nor U10239 (N_10239,N_2489,N_1961);
xor U10240 (N_10240,N_1296,N_1681);
and U10241 (N_10241,N_1606,N_5181);
nand U10242 (N_10242,N_963,N_3428);
or U10243 (N_10243,N_139,N_5517);
or U10244 (N_10244,N_4440,N_5960);
or U10245 (N_10245,N_1555,N_4952);
nand U10246 (N_10246,N_378,N_5607);
or U10247 (N_10247,N_2917,N_3163);
or U10248 (N_10248,N_5750,N_4157);
xor U10249 (N_10249,N_321,N_3036);
or U10250 (N_10250,N_3409,N_148);
nor U10251 (N_10251,N_3396,N_5655);
nand U10252 (N_10252,N_4014,N_5806);
nand U10253 (N_10253,N_1140,N_1853);
nor U10254 (N_10254,N_3660,N_1759);
and U10255 (N_10255,N_5137,N_4850);
xor U10256 (N_10256,N_964,N_4987);
nand U10257 (N_10257,N_874,N_1075);
nor U10258 (N_10258,N_1134,N_445);
xor U10259 (N_10259,N_2945,N_2006);
nor U10260 (N_10260,N_1625,N_5060);
and U10261 (N_10261,N_2457,N_3958);
xor U10262 (N_10262,N_4645,N_4198);
or U10263 (N_10263,N_1352,N_2659);
xor U10264 (N_10264,N_2770,N_1357);
nor U10265 (N_10265,N_2846,N_68);
or U10266 (N_10266,N_3169,N_3465);
and U10267 (N_10267,N_4237,N_4090);
xor U10268 (N_10268,N_4258,N_866);
and U10269 (N_10269,N_4531,N_2455);
or U10270 (N_10270,N_4109,N_5235);
nor U10271 (N_10271,N_1889,N_1566);
and U10272 (N_10272,N_4085,N_1828);
or U10273 (N_10273,N_4133,N_612);
nor U10274 (N_10274,N_1566,N_4797);
xnor U10275 (N_10275,N_1302,N_2955);
nand U10276 (N_10276,N_740,N_687);
xnor U10277 (N_10277,N_3943,N_1499);
and U10278 (N_10278,N_2808,N_103);
or U10279 (N_10279,N_3096,N_5406);
nor U10280 (N_10280,N_5468,N_4116);
xnor U10281 (N_10281,N_384,N_1349);
and U10282 (N_10282,N_4600,N_5116);
or U10283 (N_10283,N_4603,N_2312);
xnor U10284 (N_10284,N_1952,N_5332);
nand U10285 (N_10285,N_842,N_3966);
and U10286 (N_10286,N_4379,N_2203);
nor U10287 (N_10287,N_1499,N_5115);
and U10288 (N_10288,N_4565,N_4778);
xnor U10289 (N_10289,N_5090,N_3296);
xnor U10290 (N_10290,N_372,N_3059);
and U10291 (N_10291,N_157,N_180);
nor U10292 (N_10292,N_4521,N_2690);
nand U10293 (N_10293,N_2160,N_2050);
and U10294 (N_10294,N_5742,N_2374);
and U10295 (N_10295,N_4422,N_5802);
and U10296 (N_10296,N_2343,N_3182);
nor U10297 (N_10297,N_1287,N_4706);
nand U10298 (N_10298,N_2594,N_149);
or U10299 (N_10299,N_5856,N_5980);
xnor U10300 (N_10300,N_4657,N_2433);
and U10301 (N_10301,N_2097,N_4122);
nor U10302 (N_10302,N_5589,N_1348);
nand U10303 (N_10303,N_566,N_4930);
nand U10304 (N_10304,N_3883,N_5510);
nor U10305 (N_10305,N_545,N_1223);
and U10306 (N_10306,N_1785,N_2389);
xnor U10307 (N_10307,N_2057,N_3109);
nand U10308 (N_10308,N_5789,N_1320);
nor U10309 (N_10309,N_1638,N_1486);
nand U10310 (N_10310,N_5489,N_2455);
xnor U10311 (N_10311,N_341,N_2035);
and U10312 (N_10312,N_958,N_2713);
nor U10313 (N_10313,N_2468,N_1578);
or U10314 (N_10314,N_4865,N_656);
or U10315 (N_10315,N_2960,N_5077);
nand U10316 (N_10316,N_4413,N_3253);
nor U10317 (N_10317,N_5231,N_582);
xor U10318 (N_10318,N_5184,N_191);
or U10319 (N_10319,N_728,N_4826);
or U10320 (N_10320,N_4672,N_5724);
or U10321 (N_10321,N_259,N_4099);
or U10322 (N_10322,N_374,N_5644);
nor U10323 (N_10323,N_5081,N_5183);
xor U10324 (N_10324,N_558,N_2305);
xnor U10325 (N_10325,N_2305,N_1337);
nor U10326 (N_10326,N_2490,N_4380);
and U10327 (N_10327,N_1268,N_2955);
and U10328 (N_10328,N_1054,N_280);
or U10329 (N_10329,N_4892,N_5094);
and U10330 (N_10330,N_5208,N_6229);
nor U10331 (N_10331,N_3162,N_3386);
nor U10332 (N_10332,N_5397,N_234);
or U10333 (N_10333,N_2348,N_1731);
nor U10334 (N_10334,N_5439,N_808);
nand U10335 (N_10335,N_2040,N_2808);
and U10336 (N_10336,N_4380,N_3791);
nor U10337 (N_10337,N_2656,N_4589);
xnor U10338 (N_10338,N_4005,N_4340);
xor U10339 (N_10339,N_3708,N_204);
nor U10340 (N_10340,N_4091,N_3010);
or U10341 (N_10341,N_1011,N_4242);
and U10342 (N_10342,N_1240,N_150);
xor U10343 (N_10343,N_4035,N_3115);
nand U10344 (N_10344,N_5523,N_4767);
or U10345 (N_10345,N_3520,N_2427);
nor U10346 (N_10346,N_4704,N_5729);
xnor U10347 (N_10347,N_347,N_620);
and U10348 (N_10348,N_2650,N_6189);
xnor U10349 (N_10349,N_5562,N_2497);
nor U10350 (N_10350,N_1235,N_5982);
nand U10351 (N_10351,N_3296,N_6171);
nor U10352 (N_10352,N_877,N_5179);
and U10353 (N_10353,N_5575,N_3145);
nand U10354 (N_10354,N_5082,N_746);
nand U10355 (N_10355,N_5156,N_1079);
xnor U10356 (N_10356,N_4921,N_1062);
nand U10357 (N_10357,N_5555,N_4058);
nor U10358 (N_10358,N_1816,N_2185);
nor U10359 (N_10359,N_2230,N_1899);
nor U10360 (N_10360,N_4515,N_4760);
xnor U10361 (N_10361,N_4973,N_4277);
or U10362 (N_10362,N_2161,N_1577);
xnor U10363 (N_10363,N_3828,N_4417);
nor U10364 (N_10364,N_5691,N_784);
or U10365 (N_10365,N_5013,N_6078);
nor U10366 (N_10366,N_3405,N_3294);
nor U10367 (N_10367,N_5809,N_208);
xnor U10368 (N_10368,N_1258,N_872);
xor U10369 (N_10369,N_413,N_319);
and U10370 (N_10370,N_4457,N_3990);
nand U10371 (N_10371,N_1007,N_2237);
xor U10372 (N_10372,N_1438,N_5186);
and U10373 (N_10373,N_4659,N_454);
nor U10374 (N_10374,N_5374,N_3955);
or U10375 (N_10375,N_982,N_5041);
nand U10376 (N_10376,N_531,N_2532);
or U10377 (N_10377,N_3430,N_463);
nor U10378 (N_10378,N_251,N_1155);
nor U10379 (N_10379,N_5334,N_4149);
xor U10380 (N_10380,N_2165,N_4464);
nand U10381 (N_10381,N_5877,N_4981);
xnor U10382 (N_10382,N_2027,N_3519);
and U10383 (N_10383,N_1220,N_4141);
nand U10384 (N_10384,N_105,N_791);
and U10385 (N_10385,N_2784,N_911);
nand U10386 (N_10386,N_48,N_6120);
nand U10387 (N_10387,N_3572,N_3770);
and U10388 (N_10388,N_1711,N_3412);
or U10389 (N_10389,N_1498,N_1774);
nor U10390 (N_10390,N_4455,N_727);
nand U10391 (N_10391,N_2328,N_407);
nand U10392 (N_10392,N_2038,N_5464);
or U10393 (N_10393,N_3282,N_294);
or U10394 (N_10394,N_4203,N_4765);
xnor U10395 (N_10395,N_2851,N_6124);
nor U10396 (N_10396,N_515,N_5919);
and U10397 (N_10397,N_2701,N_3475);
and U10398 (N_10398,N_5139,N_5443);
nor U10399 (N_10399,N_3758,N_186);
nand U10400 (N_10400,N_4221,N_3542);
and U10401 (N_10401,N_5635,N_2924);
and U10402 (N_10402,N_4917,N_3566);
or U10403 (N_10403,N_1038,N_1140);
or U10404 (N_10404,N_3098,N_5672);
xnor U10405 (N_10405,N_4832,N_1148);
nor U10406 (N_10406,N_4736,N_3929);
nand U10407 (N_10407,N_2812,N_4843);
nand U10408 (N_10408,N_5019,N_2013);
or U10409 (N_10409,N_3831,N_1276);
or U10410 (N_10410,N_4724,N_3591);
or U10411 (N_10411,N_4954,N_2702);
and U10412 (N_10412,N_3444,N_3275);
nand U10413 (N_10413,N_5527,N_2629);
xnor U10414 (N_10414,N_2602,N_1550);
nand U10415 (N_10415,N_5930,N_6176);
and U10416 (N_10416,N_93,N_165);
xor U10417 (N_10417,N_5281,N_3483);
and U10418 (N_10418,N_6228,N_2456);
xnor U10419 (N_10419,N_2932,N_4690);
and U10420 (N_10420,N_4830,N_2586);
and U10421 (N_10421,N_2451,N_85);
xnor U10422 (N_10422,N_826,N_5103);
or U10423 (N_10423,N_5431,N_2774);
nor U10424 (N_10424,N_1283,N_2746);
nand U10425 (N_10425,N_4566,N_3963);
or U10426 (N_10426,N_5011,N_4299);
nor U10427 (N_10427,N_1659,N_2224);
nor U10428 (N_10428,N_4360,N_1112);
xor U10429 (N_10429,N_6041,N_4719);
nand U10430 (N_10430,N_2538,N_553);
nand U10431 (N_10431,N_3174,N_2463);
nor U10432 (N_10432,N_3239,N_5904);
nor U10433 (N_10433,N_67,N_2279);
nand U10434 (N_10434,N_3397,N_771);
and U10435 (N_10435,N_3441,N_1402);
and U10436 (N_10436,N_5831,N_3650);
and U10437 (N_10437,N_3839,N_2271);
nor U10438 (N_10438,N_4854,N_2417);
nor U10439 (N_10439,N_5104,N_3698);
or U10440 (N_10440,N_2904,N_2493);
and U10441 (N_10441,N_1681,N_4518);
nand U10442 (N_10442,N_5585,N_2729);
or U10443 (N_10443,N_4303,N_5662);
nand U10444 (N_10444,N_1624,N_4868);
or U10445 (N_10445,N_4627,N_4994);
nand U10446 (N_10446,N_3291,N_499);
or U10447 (N_10447,N_1170,N_3604);
or U10448 (N_10448,N_2019,N_4471);
and U10449 (N_10449,N_3344,N_2729);
xor U10450 (N_10450,N_3543,N_227);
xnor U10451 (N_10451,N_2287,N_1645);
and U10452 (N_10452,N_3735,N_2448);
nand U10453 (N_10453,N_6100,N_5708);
or U10454 (N_10454,N_5183,N_5688);
or U10455 (N_10455,N_4346,N_4996);
or U10456 (N_10456,N_3154,N_3397);
nand U10457 (N_10457,N_5270,N_281);
and U10458 (N_10458,N_2080,N_1280);
xnor U10459 (N_10459,N_5671,N_5614);
and U10460 (N_10460,N_1021,N_5564);
nand U10461 (N_10461,N_1548,N_5158);
xor U10462 (N_10462,N_1780,N_1684);
or U10463 (N_10463,N_4734,N_4544);
or U10464 (N_10464,N_3401,N_3080);
or U10465 (N_10465,N_4205,N_2501);
xor U10466 (N_10466,N_5919,N_4498);
xor U10467 (N_10467,N_4797,N_5464);
nor U10468 (N_10468,N_5181,N_1083);
xnor U10469 (N_10469,N_4705,N_4891);
nor U10470 (N_10470,N_769,N_3706);
or U10471 (N_10471,N_2820,N_1365);
or U10472 (N_10472,N_1104,N_2983);
and U10473 (N_10473,N_379,N_4831);
nor U10474 (N_10474,N_4395,N_2583);
nor U10475 (N_10475,N_849,N_3197);
xor U10476 (N_10476,N_133,N_3246);
or U10477 (N_10477,N_6222,N_3506);
nand U10478 (N_10478,N_249,N_3696);
xor U10479 (N_10479,N_2440,N_4125);
or U10480 (N_10480,N_4606,N_5691);
nand U10481 (N_10481,N_5015,N_4936);
and U10482 (N_10482,N_2937,N_1968);
nor U10483 (N_10483,N_1704,N_5109);
and U10484 (N_10484,N_5066,N_6235);
and U10485 (N_10485,N_130,N_192);
nand U10486 (N_10486,N_2222,N_1627);
nor U10487 (N_10487,N_194,N_5301);
nor U10488 (N_10488,N_5506,N_4038);
xnor U10489 (N_10489,N_4017,N_2355);
nor U10490 (N_10490,N_2681,N_1196);
or U10491 (N_10491,N_1263,N_4194);
and U10492 (N_10492,N_1684,N_906);
nor U10493 (N_10493,N_5274,N_4954);
or U10494 (N_10494,N_4730,N_6094);
and U10495 (N_10495,N_3803,N_3106);
or U10496 (N_10496,N_245,N_5671);
or U10497 (N_10497,N_5511,N_2257);
or U10498 (N_10498,N_1847,N_1796);
and U10499 (N_10499,N_5472,N_3336);
or U10500 (N_10500,N_180,N_4170);
nand U10501 (N_10501,N_5794,N_2612);
xnor U10502 (N_10502,N_4877,N_4926);
nor U10503 (N_10503,N_275,N_3899);
and U10504 (N_10504,N_1856,N_2227);
or U10505 (N_10505,N_1609,N_4504);
and U10506 (N_10506,N_150,N_3098);
and U10507 (N_10507,N_566,N_1285);
nand U10508 (N_10508,N_3578,N_3654);
nand U10509 (N_10509,N_2288,N_5133);
xnor U10510 (N_10510,N_700,N_1959);
nor U10511 (N_10511,N_1266,N_3469);
and U10512 (N_10512,N_4112,N_1519);
xnor U10513 (N_10513,N_1145,N_4691);
nand U10514 (N_10514,N_427,N_6030);
or U10515 (N_10515,N_6003,N_4137);
nor U10516 (N_10516,N_1800,N_242);
nor U10517 (N_10517,N_5052,N_5352);
nor U10518 (N_10518,N_176,N_221);
nor U10519 (N_10519,N_5427,N_2050);
nor U10520 (N_10520,N_1054,N_814);
xor U10521 (N_10521,N_4900,N_79);
nor U10522 (N_10522,N_362,N_3409);
nand U10523 (N_10523,N_5549,N_2581);
xor U10524 (N_10524,N_1564,N_1527);
or U10525 (N_10525,N_1938,N_409);
and U10526 (N_10526,N_991,N_4015);
or U10527 (N_10527,N_3892,N_3745);
nor U10528 (N_10528,N_6092,N_1863);
xor U10529 (N_10529,N_2495,N_559);
nand U10530 (N_10530,N_3873,N_5369);
and U10531 (N_10531,N_4961,N_916);
nor U10532 (N_10532,N_4805,N_2678);
nor U10533 (N_10533,N_3992,N_2832);
or U10534 (N_10534,N_4759,N_5343);
or U10535 (N_10535,N_5201,N_4081);
and U10536 (N_10536,N_3747,N_1461);
and U10537 (N_10537,N_5258,N_6187);
nand U10538 (N_10538,N_1322,N_1404);
and U10539 (N_10539,N_5545,N_5732);
or U10540 (N_10540,N_2390,N_5528);
nor U10541 (N_10541,N_3421,N_4942);
nand U10542 (N_10542,N_4929,N_219);
and U10543 (N_10543,N_4767,N_5097);
nor U10544 (N_10544,N_56,N_2690);
nand U10545 (N_10545,N_1031,N_2256);
xnor U10546 (N_10546,N_4470,N_3890);
and U10547 (N_10547,N_5880,N_474);
or U10548 (N_10548,N_2815,N_1797);
or U10549 (N_10549,N_4212,N_5414);
xor U10550 (N_10550,N_5878,N_5517);
nand U10551 (N_10551,N_1452,N_2054);
and U10552 (N_10552,N_6127,N_3357);
or U10553 (N_10553,N_3627,N_4109);
and U10554 (N_10554,N_306,N_6001);
xnor U10555 (N_10555,N_3917,N_1169);
and U10556 (N_10556,N_2826,N_2240);
nand U10557 (N_10557,N_4736,N_434);
nand U10558 (N_10558,N_4830,N_3486);
xor U10559 (N_10559,N_6034,N_1019);
or U10560 (N_10560,N_1012,N_3853);
or U10561 (N_10561,N_2185,N_3169);
or U10562 (N_10562,N_5305,N_2550);
or U10563 (N_10563,N_5878,N_5559);
xnor U10564 (N_10564,N_3932,N_5423);
and U10565 (N_10565,N_3072,N_92);
or U10566 (N_10566,N_1796,N_4355);
or U10567 (N_10567,N_5056,N_3051);
and U10568 (N_10568,N_826,N_202);
nand U10569 (N_10569,N_3439,N_1542);
and U10570 (N_10570,N_4917,N_120);
nor U10571 (N_10571,N_748,N_795);
nor U10572 (N_10572,N_2453,N_5137);
xnor U10573 (N_10573,N_3837,N_5608);
or U10574 (N_10574,N_4088,N_5530);
xor U10575 (N_10575,N_4578,N_3112);
or U10576 (N_10576,N_721,N_3303);
xor U10577 (N_10577,N_3888,N_4142);
or U10578 (N_10578,N_3565,N_5529);
xor U10579 (N_10579,N_4789,N_537);
or U10580 (N_10580,N_3426,N_4927);
and U10581 (N_10581,N_5664,N_1476);
xor U10582 (N_10582,N_1611,N_5743);
nor U10583 (N_10583,N_3687,N_3591);
nand U10584 (N_10584,N_6022,N_3615);
nand U10585 (N_10585,N_1756,N_2307);
nand U10586 (N_10586,N_1073,N_1359);
or U10587 (N_10587,N_4091,N_3556);
nand U10588 (N_10588,N_3330,N_5167);
xor U10589 (N_10589,N_830,N_168);
nand U10590 (N_10590,N_3784,N_6233);
or U10591 (N_10591,N_899,N_4902);
nor U10592 (N_10592,N_3019,N_128);
and U10593 (N_10593,N_5296,N_2848);
nand U10594 (N_10594,N_29,N_1558);
and U10595 (N_10595,N_5225,N_635);
xor U10596 (N_10596,N_2701,N_1052);
or U10597 (N_10597,N_318,N_3370);
and U10598 (N_10598,N_54,N_3662);
nor U10599 (N_10599,N_1278,N_2614);
nor U10600 (N_10600,N_6013,N_4995);
xnor U10601 (N_10601,N_4082,N_4778);
or U10602 (N_10602,N_884,N_1969);
nor U10603 (N_10603,N_5955,N_3658);
and U10604 (N_10604,N_4166,N_2675);
xnor U10605 (N_10605,N_2176,N_429);
nor U10606 (N_10606,N_2029,N_1457);
xnor U10607 (N_10607,N_30,N_4882);
xnor U10608 (N_10608,N_5898,N_2414);
nand U10609 (N_10609,N_3327,N_359);
nor U10610 (N_10610,N_3630,N_2240);
xor U10611 (N_10611,N_5686,N_1263);
and U10612 (N_10612,N_1641,N_1355);
xnor U10613 (N_10613,N_391,N_2144);
xnor U10614 (N_10614,N_2517,N_4059);
or U10615 (N_10615,N_4559,N_547);
xnor U10616 (N_10616,N_2469,N_1318);
nand U10617 (N_10617,N_6005,N_204);
xor U10618 (N_10618,N_5005,N_4653);
and U10619 (N_10619,N_1474,N_638);
and U10620 (N_10620,N_750,N_1619);
nor U10621 (N_10621,N_5605,N_1325);
and U10622 (N_10622,N_3008,N_5085);
or U10623 (N_10623,N_5612,N_6094);
or U10624 (N_10624,N_2135,N_6118);
and U10625 (N_10625,N_9,N_3222);
nor U10626 (N_10626,N_2353,N_5841);
nor U10627 (N_10627,N_2045,N_1055);
nor U10628 (N_10628,N_1803,N_5505);
or U10629 (N_10629,N_1261,N_39);
xor U10630 (N_10630,N_2587,N_3288);
xor U10631 (N_10631,N_2566,N_3955);
nor U10632 (N_10632,N_1932,N_4758);
and U10633 (N_10633,N_5327,N_5296);
or U10634 (N_10634,N_91,N_3463);
or U10635 (N_10635,N_1706,N_2955);
or U10636 (N_10636,N_4006,N_4675);
nand U10637 (N_10637,N_3246,N_4912);
or U10638 (N_10638,N_2462,N_2651);
or U10639 (N_10639,N_533,N_3065);
and U10640 (N_10640,N_1377,N_4703);
and U10641 (N_10641,N_448,N_2391);
xor U10642 (N_10642,N_2170,N_5030);
and U10643 (N_10643,N_4540,N_1831);
nand U10644 (N_10644,N_2763,N_3513);
or U10645 (N_10645,N_4915,N_4364);
nand U10646 (N_10646,N_4745,N_4256);
nor U10647 (N_10647,N_315,N_5062);
or U10648 (N_10648,N_4325,N_5967);
nor U10649 (N_10649,N_5638,N_4048);
or U10650 (N_10650,N_3978,N_3315);
nand U10651 (N_10651,N_3312,N_5196);
or U10652 (N_10652,N_1894,N_1244);
nor U10653 (N_10653,N_645,N_589);
or U10654 (N_10654,N_5220,N_2724);
nand U10655 (N_10655,N_4100,N_2883);
nand U10656 (N_10656,N_4601,N_3401);
nand U10657 (N_10657,N_5529,N_2590);
xnor U10658 (N_10658,N_4851,N_1312);
or U10659 (N_10659,N_2847,N_340);
xnor U10660 (N_10660,N_441,N_332);
nand U10661 (N_10661,N_3807,N_6006);
nand U10662 (N_10662,N_172,N_2081);
xor U10663 (N_10663,N_6231,N_1321);
and U10664 (N_10664,N_904,N_956);
nor U10665 (N_10665,N_2387,N_2978);
nand U10666 (N_10666,N_5218,N_4363);
xnor U10667 (N_10667,N_4305,N_4285);
and U10668 (N_10668,N_1898,N_5899);
nand U10669 (N_10669,N_4699,N_2200);
or U10670 (N_10670,N_2046,N_1841);
nor U10671 (N_10671,N_859,N_570);
or U10672 (N_10672,N_1564,N_5530);
xor U10673 (N_10673,N_5364,N_2580);
xor U10674 (N_10674,N_5166,N_1588);
and U10675 (N_10675,N_1473,N_3007);
nand U10676 (N_10676,N_817,N_355);
nand U10677 (N_10677,N_1334,N_3193);
and U10678 (N_10678,N_296,N_6008);
and U10679 (N_10679,N_5509,N_1223);
and U10680 (N_10680,N_2804,N_4131);
or U10681 (N_10681,N_5418,N_256);
or U10682 (N_10682,N_2484,N_2737);
nand U10683 (N_10683,N_1681,N_3274);
or U10684 (N_10684,N_3052,N_1115);
or U10685 (N_10685,N_1144,N_1435);
or U10686 (N_10686,N_5980,N_105);
nand U10687 (N_10687,N_1671,N_733);
or U10688 (N_10688,N_3917,N_5296);
xor U10689 (N_10689,N_5264,N_1807);
nand U10690 (N_10690,N_3931,N_4499);
xor U10691 (N_10691,N_896,N_2215);
nand U10692 (N_10692,N_3890,N_2564);
or U10693 (N_10693,N_587,N_5882);
nand U10694 (N_10694,N_5697,N_2499);
xnor U10695 (N_10695,N_5623,N_1730);
nor U10696 (N_10696,N_768,N_1617);
xor U10697 (N_10697,N_2770,N_5376);
and U10698 (N_10698,N_1727,N_3836);
or U10699 (N_10699,N_2095,N_2168);
and U10700 (N_10700,N_3125,N_1784);
or U10701 (N_10701,N_4545,N_3256);
nor U10702 (N_10702,N_3887,N_5171);
xor U10703 (N_10703,N_700,N_84);
xor U10704 (N_10704,N_1073,N_5574);
nand U10705 (N_10705,N_3200,N_3598);
xor U10706 (N_10706,N_2680,N_837);
nor U10707 (N_10707,N_5194,N_741);
or U10708 (N_10708,N_1396,N_4751);
or U10709 (N_10709,N_2563,N_5069);
and U10710 (N_10710,N_3746,N_4227);
nand U10711 (N_10711,N_4096,N_470);
xnor U10712 (N_10712,N_178,N_5859);
xor U10713 (N_10713,N_6168,N_4297);
nand U10714 (N_10714,N_79,N_3350);
nand U10715 (N_10715,N_2311,N_1881);
and U10716 (N_10716,N_2545,N_4633);
and U10717 (N_10717,N_3384,N_1604);
nor U10718 (N_10718,N_1994,N_5030);
or U10719 (N_10719,N_2910,N_872);
and U10720 (N_10720,N_3432,N_4391);
xor U10721 (N_10721,N_4665,N_4024);
or U10722 (N_10722,N_3075,N_2815);
or U10723 (N_10723,N_3351,N_238);
xor U10724 (N_10724,N_2416,N_4162);
or U10725 (N_10725,N_6042,N_3762);
nand U10726 (N_10726,N_3979,N_547);
and U10727 (N_10727,N_1721,N_5888);
xor U10728 (N_10728,N_2863,N_3151);
xnor U10729 (N_10729,N_1461,N_2668);
and U10730 (N_10730,N_1960,N_2733);
and U10731 (N_10731,N_4206,N_881);
and U10732 (N_10732,N_5877,N_5497);
xnor U10733 (N_10733,N_4989,N_1757);
and U10734 (N_10734,N_2787,N_2961);
xor U10735 (N_10735,N_2152,N_5072);
or U10736 (N_10736,N_4725,N_2010);
xor U10737 (N_10737,N_1175,N_3095);
and U10738 (N_10738,N_1379,N_5234);
xnor U10739 (N_10739,N_4342,N_3924);
nor U10740 (N_10740,N_4966,N_6143);
nand U10741 (N_10741,N_2229,N_3188);
nand U10742 (N_10742,N_2684,N_2873);
nand U10743 (N_10743,N_4546,N_4623);
and U10744 (N_10744,N_3141,N_31);
xnor U10745 (N_10745,N_4014,N_106);
xnor U10746 (N_10746,N_3525,N_466);
xnor U10747 (N_10747,N_3969,N_841);
and U10748 (N_10748,N_1927,N_2774);
xnor U10749 (N_10749,N_5234,N_1829);
nand U10750 (N_10750,N_3841,N_1410);
nor U10751 (N_10751,N_3106,N_3291);
nor U10752 (N_10752,N_1908,N_1828);
nor U10753 (N_10753,N_2752,N_1605);
or U10754 (N_10754,N_2132,N_5467);
nand U10755 (N_10755,N_4185,N_2600);
nor U10756 (N_10756,N_3009,N_372);
nand U10757 (N_10757,N_1695,N_4135);
or U10758 (N_10758,N_87,N_1613);
nand U10759 (N_10759,N_4199,N_1228);
xor U10760 (N_10760,N_302,N_1673);
nand U10761 (N_10761,N_2329,N_180);
nor U10762 (N_10762,N_6166,N_6011);
and U10763 (N_10763,N_4412,N_5480);
xnor U10764 (N_10764,N_952,N_116);
nand U10765 (N_10765,N_1863,N_1233);
nand U10766 (N_10766,N_3341,N_665);
nor U10767 (N_10767,N_6053,N_3228);
and U10768 (N_10768,N_1566,N_285);
nand U10769 (N_10769,N_1575,N_645);
and U10770 (N_10770,N_5692,N_6187);
and U10771 (N_10771,N_2519,N_2665);
and U10772 (N_10772,N_691,N_4984);
and U10773 (N_10773,N_168,N_3554);
or U10774 (N_10774,N_6055,N_4149);
and U10775 (N_10775,N_3879,N_5800);
nor U10776 (N_10776,N_827,N_2322);
nor U10777 (N_10777,N_374,N_344);
xor U10778 (N_10778,N_2452,N_6154);
xor U10779 (N_10779,N_322,N_790);
nand U10780 (N_10780,N_3247,N_5409);
xor U10781 (N_10781,N_836,N_5237);
nor U10782 (N_10782,N_4783,N_229);
xnor U10783 (N_10783,N_3025,N_4549);
and U10784 (N_10784,N_663,N_3044);
or U10785 (N_10785,N_6175,N_2897);
and U10786 (N_10786,N_5285,N_4987);
nand U10787 (N_10787,N_1245,N_1609);
or U10788 (N_10788,N_1626,N_5609);
and U10789 (N_10789,N_351,N_986);
and U10790 (N_10790,N_1374,N_396);
and U10791 (N_10791,N_1384,N_2947);
or U10792 (N_10792,N_6213,N_5833);
xor U10793 (N_10793,N_4371,N_2018);
or U10794 (N_10794,N_855,N_3365);
nand U10795 (N_10795,N_1273,N_3132);
and U10796 (N_10796,N_1872,N_6182);
nor U10797 (N_10797,N_4188,N_4312);
xor U10798 (N_10798,N_1946,N_2210);
or U10799 (N_10799,N_5977,N_5336);
or U10800 (N_10800,N_618,N_1454);
or U10801 (N_10801,N_3580,N_2968);
or U10802 (N_10802,N_6227,N_4627);
nand U10803 (N_10803,N_6025,N_1364);
nor U10804 (N_10804,N_4728,N_4317);
nor U10805 (N_10805,N_5976,N_2036);
and U10806 (N_10806,N_5022,N_1993);
and U10807 (N_10807,N_4327,N_3616);
nor U10808 (N_10808,N_4079,N_2327);
xnor U10809 (N_10809,N_4516,N_2887);
and U10810 (N_10810,N_3676,N_3062);
or U10811 (N_10811,N_1885,N_1257);
or U10812 (N_10812,N_5003,N_3764);
nor U10813 (N_10813,N_1449,N_5376);
xor U10814 (N_10814,N_698,N_5566);
or U10815 (N_10815,N_4647,N_1369);
xor U10816 (N_10816,N_2242,N_4038);
or U10817 (N_10817,N_1181,N_2321);
and U10818 (N_10818,N_2081,N_1931);
nor U10819 (N_10819,N_3888,N_4433);
xor U10820 (N_10820,N_2226,N_3947);
nor U10821 (N_10821,N_988,N_4793);
and U10822 (N_10822,N_318,N_3294);
and U10823 (N_10823,N_3895,N_939);
xor U10824 (N_10824,N_2727,N_2253);
or U10825 (N_10825,N_2346,N_4232);
or U10826 (N_10826,N_2501,N_5478);
xor U10827 (N_10827,N_4960,N_2849);
nand U10828 (N_10828,N_2021,N_562);
or U10829 (N_10829,N_2890,N_4135);
xor U10830 (N_10830,N_5999,N_5591);
or U10831 (N_10831,N_1326,N_3807);
nor U10832 (N_10832,N_4092,N_438);
nor U10833 (N_10833,N_3682,N_4107);
and U10834 (N_10834,N_1101,N_4308);
nor U10835 (N_10835,N_4392,N_6139);
nor U10836 (N_10836,N_3758,N_1408);
or U10837 (N_10837,N_932,N_371);
nand U10838 (N_10838,N_1060,N_1041);
nand U10839 (N_10839,N_5192,N_4104);
and U10840 (N_10840,N_2545,N_963);
nor U10841 (N_10841,N_4393,N_1179);
or U10842 (N_10842,N_4818,N_3906);
nand U10843 (N_10843,N_695,N_2420);
xor U10844 (N_10844,N_5104,N_5088);
and U10845 (N_10845,N_1101,N_1589);
or U10846 (N_10846,N_3678,N_250);
nor U10847 (N_10847,N_3889,N_2631);
nand U10848 (N_10848,N_3897,N_6123);
and U10849 (N_10849,N_1703,N_4270);
xor U10850 (N_10850,N_6163,N_3095);
xor U10851 (N_10851,N_2412,N_2350);
and U10852 (N_10852,N_5289,N_230);
nor U10853 (N_10853,N_798,N_4544);
nor U10854 (N_10854,N_2539,N_2825);
and U10855 (N_10855,N_5787,N_1590);
nor U10856 (N_10856,N_3064,N_3854);
and U10857 (N_10857,N_5902,N_5162);
or U10858 (N_10858,N_101,N_4725);
xnor U10859 (N_10859,N_3833,N_4732);
or U10860 (N_10860,N_2124,N_777);
xnor U10861 (N_10861,N_2111,N_2668);
xor U10862 (N_10862,N_3806,N_3700);
nor U10863 (N_10863,N_2613,N_5719);
nand U10864 (N_10864,N_4633,N_1128);
nand U10865 (N_10865,N_3413,N_38);
nor U10866 (N_10866,N_5370,N_1349);
xor U10867 (N_10867,N_3007,N_4171);
xnor U10868 (N_10868,N_1888,N_6060);
or U10869 (N_10869,N_4485,N_936);
or U10870 (N_10870,N_1524,N_5452);
nand U10871 (N_10871,N_4918,N_3141);
xor U10872 (N_10872,N_629,N_5375);
nand U10873 (N_10873,N_1379,N_4304);
nand U10874 (N_10874,N_5557,N_5121);
nand U10875 (N_10875,N_4714,N_2528);
or U10876 (N_10876,N_2271,N_886);
and U10877 (N_10877,N_5292,N_5903);
nand U10878 (N_10878,N_251,N_3398);
or U10879 (N_10879,N_3962,N_5023);
nand U10880 (N_10880,N_2213,N_1271);
or U10881 (N_10881,N_6204,N_6114);
xnor U10882 (N_10882,N_1089,N_555);
xnor U10883 (N_10883,N_3643,N_794);
nor U10884 (N_10884,N_1715,N_2722);
nand U10885 (N_10885,N_2667,N_4689);
and U10886 (N_10886,N_4973,N_5732);
and U10887 (N_10887,N_2541,N_5347);
and U10888 (N_10888,N_5706,N_5358);
or U10889 (N_10889,N_5540,N_424);
or U10890 (N_10890,N_4361,N_4420);
and U10891 (N_10891,N_5492,N_1158);
xor U10892 (N_10892,N_1134,N_5683);
xor U10893 (N_10893,N_4779,N_3645);
nand U10894 (N_10894,N_5718,N_373);
or U10895 (N_10895,N_274,N_2928);
nor U10896 (N_10896,N_179,N_1120);
and U10897 (N_10897,N_4900,N_4918);
nand U10898 (N_10898,N_6244,N_1707);
xor U10899 (N_10899,N_6164,N_5012);
or U10900 (N_10900,N_3548,N_1895);
or U10901 (N_10901,N_5545,N_3252);
or U10902 (N_10902,N_5427,N_4816);
or U10903 (N_10903,N_2745,N_4908);
nor U10904 (N_10904,N_4375,N_3469);
nor U10905 (N_10905,N_2597,N_307);
nor U10906 (N_10906,N_1511,N_2537);
nand U10907 (N_10907,N_2550,N_3560);
nand U10908 (N_10908,N_112,N_4262);
and U10909 (N_10909,N_4925,N_5329);
nor U10910 (N_10910,N_5679,N_4854);
or U10911 (N_10911,N_1925,N_5832);
and U10912 (N_10912,N_2554,N_4400);
and U10913 (N_10913,N_4004,N_324);
xor U10914 (N_10914,N_3700,N_5197);
or U10915 (N_10915,N_5926,N_4175);
nor U10916 (N_10916,N_5046,N_636);
nand U10917 (N_10917,N_3899,N_1031);
or U10918 (N_10918,N_6243,N_4856);
nor U10919 (N_10919,N_2018,N_6074);
xnor U10920 (N_10920,N_6079,N_745);
nor U10921 (N_10921,N_5566,N_4470);
xnor U10922 (N_10922,N_5318,N_1819);
and U10923 (N_10923,N_2555,N_4212);
xor U10924 (N_10924,N_1419,N_5675);
nand U10925 (N_10925,N_4835,N_1050);
nand U10926 (N_10926,N_1748,N_2737);
and U10927 (N_10927,N_5860,N_5453);
nor U10928 (N_10928,N_4860,N_992);
and U10929 (N_10929,N_1830,N_5422);
nor U10930 (N_10930,N_4535,N_6053);
or U10931 (N_10931,N_5182,N_2322);
nand U10932 (N_10932,N_2021,N_2230);
or U10933 (N_10933,N_4394,N_5668);
nand U10934 (N_10934,N_133,N_2604);
or U10935 (N_10935,N_5969,N_3398);
nand U10936 (N_10936,N_3712,N_1807);
or U10937 (N_10937,N_3323,N_2);
or U10938 (N_10938,N_3626,N_1593);
xor U10939 (N_10939,N_2981,N_6195);
or U10940 (N_10940,N_5129,N_467);
nor U10941 (N_10941,N_2070,N_478);
nor U10942 (N_10942,N_5401,N_3495);
nor U10943 (N_10943,N_3746,N_2920);
xor U10944 (N_10944,N_4260,N_5714);
and U10945 (N_10945,N_3081,N_1180);
and U10946 (N_10946,N_6232,N_1638);
nand U10947 (N_10947,N_1675,N_121);
and U10948 (N_10948,N_4868,N_4982);
and U10949 (N_10949,N_1954,N_3866);
and U10950 (N_10950,N_5927,N_5347);
or U10951 (N_10951,N_2432,N_833);
and U10952 (N_10952,N_4692,N_4742);
nand U10953 (N_10953,N_5874,N_4812);
and U10954 (N_10954,N_2936,N_532);
nand U10955 (N_10955,N_6112,N_5360);
or U10956 (N_10956,N_700,N_1067);
nand U10957 (N_10957,N_1066,N_6128);
nand U10958 (N_10958,N_5729,N_6151);
and U10959 (N_10959,N_1441,N_3421);
nand U10960 (N_10960,N_3294,N_3130);
or U10961 (N_10961,N_5542,N_694);
and U10962 (N_10962,N_155,N_686);
xor U10963 (N_10963,N_3472,N_4694);
or U10964 (N_10964,N_3030,N_2063);
nand U10965 (N_10965,N_4268,N_2219);
nor U10966 (N_10966,N_1149,N_4782);
xnor U10967 (N_10967,N_5164,N_5997);
xor U10968 (N_10968,N_459,N_1083);
xnor U10969 (N_10969,N_3221,N_6189);
or U10970 (N_10970,N_207,N_5068);
or U10971 (N_10971,N_271,N_968);
nor U10972 (N_10972,N_2145,N_4299);
nor U10973 (N_10973,N_5119,N_2297);
and U10974 (N_10974,N_3442,N_3014);
or U10975 (N_10975,N_3490,N_132);
or U10976 (N_10976,N_3614,N_2626);
xnor U10977 (N_10977,N_2712,N_520);
nor U10978 (N_10978,N_1822,N_6006);
and U10979 (N_10979,N_413,N_3863);
and U10980 (N_10980,N_2375,N_2419);
and U10981 (N_10981,N_3958,N_5471);
or U10982 (N_10982,N_112,N_3063);
xnor U10983 (N_10983,N_2474,N_1074);
and U10984 (N_10984,N_905,N_3544);
or U10985 (N_10985,N_2443,N_5635);
xor U10986 (N_10986,N_5375,N_2124);
or U10987 (N_10987,N_918,N_5371);
nor U10988 (N_10988,N_1664,N_5908);
nand U10989 (N_10989,N_986,N_3667);
or U10990 (N_10990,N_4739,N_2953);
nor U10991 (N_10991,N_2700,N_1316);
nor U10992 (N_10992,N_3648,N_5023);
xor U10993 (N_10993,N_1342,N_3035);
and U10994 (N_10994,N_3777,N_6120);
nand U10995 (N_10995,N_1172,N_4290);
xnor U10996 (N_10996,N_4978,N_4970);
or U10997 (N_10997,N_5171,N_4823);
nand U10998 (N_10998,N_3270,N_1992);
and U10999 (N_10999,N_1189,N_3679);
nand U11000 (N_11000,N_5568,N_292);
and U11001 (N_11001,N_3321,N_3710);
and U11002 (N_11002,N_5312,N_2747);
nor U11003 (N_11003,N_1491,N_1570);
nand U11004 (N_11004,N_1287,N_5750);
or U11005 (N_11005,N_3459,N_1392);
xor U11006 (N_11006,N_3093,N_2713);
or U11007 (N_11007,N_4080,N_5514);
nor U11008 (N_11008,N_3710,N_2107);
nor U11009 (N_11009,N_2871,N_3449);
nand U11010 (N_11010,N_5660,N_700);
and U11011 (N_11011,N_1648,N_1620);
or U11012 (N_11012,N_4876,N_4719);
nor U11013 (N_11013,N_4003,N_29);
and U11014 (N_11014,N_1374,N_1537);
nor U11015 (N_11015,N_5372,N_5368);
or U11016 (N_11016,N_1097,N_296);
nor U11017 (N_11017,N_339,N_1331);
nand U11018 (N_11018,N_3400,N_5532);
nand U11019 (N_11019,N_4044,N_2229);
or U11020 (N_11020,N_454,N_4070);
xor U11021 (N_11021,N_241,N_175);
nor U11022 (N_11022,N_3782,N_4959);
nand U11023 (N_11023,N_1719,N_2175);
or U11024 (N_11024,N_5696,N_6150);
nand U11025 (N_11025,N_5778,N_2495);
and U11026 (N_11026,N_3743,N_65);
xor U11027 (N_11027,N_4055,N_3818);
nand U11028 (N_11028,N_5222,N_1218);
nor U11029 (N_11029,N_3652,N_814);
nand U11030 (N_11030,N_2887,N_1557);
or U11031 (N_11031,N_1849,N_346);
nor U11032 (N_11032,N_66,N_1761);
nor U11033 (N_11033,N_3259,N_6243);
and U11034 (N_11034,N_1700,N_3781);
nand U11035 (N_11035,N_3618,N_5344);
nand U11036 (N_11036,N_2638,N_4164);
xnor U11037 (N_11037,N_3458,N_4005);
or U11038 (N_11038,N_3956,N_1303);
nand U11039 (N_11039,N_1752,N_6136);
and U11040 (N_11040,N_2981,N_5561);
nor U11041 (N_11041,N_1034,N_960);
xnor U11042 (N_11042,N_2281,N_2674);
xnor U11043 (N_11043,N_2,N_2763);
nand U11044 (N_11044,N_1399,N_2478);
and U11045 (N_11045,N_5038,N_3196);
xnor U11046 (N_11046,N_4427,N_2017);
xor U11047 (N_11047,N_1829,N_4832);
and U11048 (N_11048,N_2693,N_3809);
nor U11049 (N_11049,N_6190,N_4635);
xor U11050 (N_11050,N_3957,N_6175);
nand U11051 (N_11051,N_4462,N_3601);
nor U11052 (N_11052,N_2770,N_1228);
xor U11053 (N_11053,N_2019,N_1116);
nand U11054 (N_11054,N_3321,N_1378);
and U11055 (N_11055,N_5236,N_3364);
nor U11056 (N_11056,N_2049,N_4698);
nor U11057 (N_11057,N_3224,N_3789);
and U11058 (N_11058,N_2646,N_5501);
and U11059 (N_11059,N_3155,N_1887);
nor U11060 (N_11060,N_4788,N_5174);
xnor U11061 (N_11061,N_4037,N_4358);
or U11062 (N_11062,N_6048,N_4672);
nand U11063 (N_11063,N_3261,N_4072);
or U11064 (N_11064,N_4394,N_600);
or U11065 (N_11065,N_4059,N_4569);
nand U11066 (N_11066,N_4096,N_4798);
nor U11067 (N_11067,N_3698,N_4706);
nand U11068 (N_11068,N_1596,N_5388);
nand U11069 (N_11069,N_1964,N_2999);
nor U11070 (N_11070,N_1847,N_759);
xnor U11071 (N_11071,N_6163,N_5635);
xor U11072 (N_11072,N_600,N_1210);
nor U11073 (N_11073,N_2310,N_1910);
xnor U11074 (N_11074,N_219,N_2655);
xor U11075 (N_11075,N_1242,N_5755);
or U11076 (N_11076,N_1470,N_5526);
xnor U11077 (N_11077,N_4673,N_5391);
xnor U11078 (N_11078,N_5810,N_3827);
nor U11079 (N_11079,N_6198,N_1393);
nor U11080 (N_11080,N_1065,N_5027);
xnor U11081 (N_11081,N_483,N_1411);
xor U11082 (N_11082,N_3504,N_6019);
nor U11083 (N_11083,N_3193,N_4438);
xnor U11084 (N_11084,N_4647,N_5740);
xnor U11085 (N_11085,N_279,N_2708);
or U11086 (N_11086,N_3327,N_5699);
or U11087 (N_11087,N_915,N_1850);
nand U11088 (N_11088,N_16,N_5899);
and U11089 (N_11089,N_5176,N_1816);
or U11090 (N_11090,N_5608,N_5340);
nand U11091 (N_11091,N_3675,N_5080);
or U11092 (N_11092,N_3190,N_1886);
nor U11093 (N_11093,N_2947,N_3603);
nor U11094 (N_11094,N_4612,N_5089);
or U11095 (N_11095,N_2578,N_5760);
and U11096 (N_11096,N_93,N_3395);
and U11097 (N_11097,N_2263,N_5535);
xnor U11098 (N_11098,N_2968,N_2924);
or U11099 (N_11099,N_5310,N_4898);
nor U11100 (N_11100,N_2256,N_1470);
and U11101 (N_11101,N_1024,N_2761);
xor U11102 (N_11102,N_440,N_1128);
nor U11103 (N_11103,N_1215,N_6215);
xnor U11104 (N_11104,N_4467,N_1991);
and U11105 (N_11105,N_4041,N_4407);
nor U11106 (N_11106,N_5221,N_5652);
or U11107 (N_11107,N_2290,N_372);
and U11108 (N_11108,N_4436,N_4872);
xor U11109 (N_11109,N_2649,N_2540);
nor U11110 (N_11110,N_3105,N_4177);
xnor U11111 (N_11111,N_2576,N_1604);
xnor U11112 (N_11112,N_2113,N_2083);
nand U11113 (N_11113,N_4933,N_1161);
xnor U11114 (N_11114,N_3670,N_295);
and U11115 (N_11115,N_6019,N_4809);
xor U11116 (N_11116,N_4966,N_4714);
and U11117 (N_11117,N_3764,N_1638);
or U11118 (N_11118,N_4729,N_5257);
or U11119 (N_11119,N_1738,N_1336);
nand U11120 (N_11120,N_585,N_417);
and U11121 (N_11121,N_5172,N_1881);
nand U11122 (N_11122,N_5385,N_1281);
xor U11123 (N_11123,N_5878,N_2289);
and U11124 (N_11124,N_3878,N_4974);
nor U11125 (N_11125,N_5657,N_2815);
or U11126 (N_11126,N_2049,N_4545);
and U11127 (N_11127,N_224,N_2634);
or U11128 (N_11128,N_2122,N_927);
or U11129 (N_11129,N_2909,N_2195);
nor U11130 (N_11130,N_2652,N_2710);
nor U11131 (N_11131,N_4998,N_4157);
nand U11132 (N_11132,N_4588,N_1307);
or U11133 (N_11133,N_5284,N_1157);
or U11134 (N_11134,N_4630,N_5204);
nor U11135 (N_11135,N_3359,N_6043);
nor U11136 (N_11136,N_5632,N_532);
nand U11137 (N_11137,N_3116,N_106);
and U11138 (N_11138,N_1707,N_3401);
xnor U11139 (N_11139,N_3950,N_6139);
nand U11140 (N_11140,N_4348,N_5569);
and U11141 (N_11141,N_4019,N_3263);
or U11142 (N_11142,N_3354,N_3);
nor U11143 (N_11143,N_4561,N_2099);
xnor U11144 (N_11144,N_1747,N_5685);
xor U11145 (N_11145,N_2452,N_2241);
nor U11146 (N_11146,N_36,N_3258);
xnor U11147 (N_11147,N_3105,N_4501);
nand U11148 (N_11148,N_5641,N_1469);
or U11149 (N_11149,N_3843,N_2070);
xnor U11150 (N_11150,N_832,N_262);
nor U11151 (N_11151,N_5438,N_2522);
xnor U11152 (N_11152,N_1462,N_2165);
nor U11153 (N_11153,N_1323,N_4358);
nor U11154 (N_11154,N_2132,N_510);
or U11155 (N_11155,N_4783,N_5049);
or U11156 (N_11156,N_2819,N_4611);
nor U11157 (N_11157,N_3026,N_3993);
nand U11158 (N_11158,N_1085,N_1609);
and U11159 (N_11159,N_4747,N_5285);
nand U11160 (N_11160,N_2256,N_405);
and U11161 (N_11161,N_150,N_927);
or U11162 (N_11162,N_1236,N_1145);
and U11163 (N_11163,N_681,N_5492);
nor U11164 (N_11164,N_2006,N_5383);
nor U11165 (N_11165,N_2286,N_2578);
nor U11166 (N_11166,N_3999,N_2735);
nand U11167 (N_11167,N_4428,N_5131);
nand U11168 (N_11168,N_3054,N_3261);
nand U11169 (N_11169,N_2163,N_5922);
nand U11170 (N_11170,N_5802,N_5813);
nand U11171 (N_11171,N_3259,N_198);
xnor U11172 (N_11172,N_3246,N_2297);
or U11173 (N_11173,N_5603,N_3114);
or U11174 (N_11174,N_2770,N_4506);
or U11175 (N_11175,N_4269,N_4164);
and U11176 (N_11176,N_746,N_5008);
or U11177 (N_11177,N_2915,N_5861);
xor U11178 (N_11178,N_4381,N_4547);
or U11179 (N_11179,N_3899,N_1930);
nor U11180 (N_11180,N_2516,N_51);
or U11181 (N_11181,N_3864,N_814);
nor U11182 (N_11182,N_2408,N_2746);
nand U11183 (N_11183,N_827,N_5351);
nor U11184 (N_11184,N_1749,N_5617);
xnor U11185 (N_11185,N_1380,N_3961);
and U11186 (N_11186,N_5734,N_91);
and U11187 (N_11187,N_4942,N_4956);
and U11188 (N_11188,N_2949,N_5551);
and U11189 (N_11189,N_3809,N_5982);
nor U11190 (N_11190,N_5435,N_4444);
nor U11191 (N_11191,N_5812,N_3126);
or U11192 (N_11192,N_4626,N_65);
nand U11193 (N_11193,N_3178,N_5337);
and U11194 (N_11194,N_993,N_3092);
nor U11195 (N_11195,N_5762,N_2948);
nor U11196 (N_11196,N_548,N_5562);
or U11197 (N_11197,N_3306,N_138);
nor U11198 (N_11198,N_28,N_3630);
xnor U11199 (N_11199,N_5616,N_1982);
xor U11200 (N_11200,N_2372,N_5730);
nand U11201 (N_11201,N_1447,N_20);
and U11202 (N_11202,N_2710,N_2334);
nand U11203 (N_11203,N_415,N_5893);
xor U11204 (N_11204,N_1557,N_4410);
nand U11205 (N_11205,N_3468,N_3254);
nor U11206 (N_11206,N_4403,N_5084);
nand U11207 (N_11207,N_1278,N_6135);
xnor U11208 (N_11208,N_3232,N_5713);
nor U11209 (N_11209,N_3099,N_4546);
nand U11210 (N_11210,N_2491,N_5432);
or U11211 (N_11211,N_2880,N_1138);
nand U11212 (N_11212,N_2856,N_5512);
or U11213 (N_11213,N_3570,N_3327);
xnor U11214 (N_11214,N_987,N_868);
xnor U11215 (N_11215,N_3882,N_3187);
or U11216 (N_11216,N_5025,N_4660);
and U11217 (N_11217,N_2738,N_480);
xnor U11218 (N_11218,N_3986,N_392);
and U11219 (N_11219,N_5249,N_5060);
and U11220 (N_11220,N_4111,N_3516);
nor U11221 (N_11221,N_3989,N_1689);
xnor U11222 (N_11222,N_1293,N_2283);
and U11223 (N_11223,N_1376,N_2370);
or U11224 (N_11224,N_4695,N_3318);
and U11225 (N_11225,N_6047,N_1085);
or U11226 (N_11226,N_2080,N_6199);
or U11227 (N_11227,N_4162,N_711);
xor U11228 (N_11228,N_160,N_1205);
nand U11229 (N_11229,N_2615,N_577);
nand U11230 (N_11230,N_2601,N_2466);
nor U11231 (N_11231,N_53,N_5459);
or U11232 (N_11232,N_493,N_3450);
or U11233 (N_11233,N_3419,N_2123);
nand U11234 (N_11234,N_3199,N_4561);
nand U11235 (N_11235,N_1369,N_6048);
and U11236 (N_11236,N_1260,N_2257);
nand U11237 (N_11237,N_1097,N_2638);
xnor U11238 (N_11238,N_3535,N_2476);
nor U11239 (N_11239,N_5934,N_1215);
xor U11240 (N_11240,N_1225,N_6046);
or U11241 (N_11241,N_3615,N_4773);
nor U11242 (N_11242,N_4003,N_4676);
nand U11243 (N_11243,N_4524,N_3706);
xor U11244 (N_11244,N_224,N_4995);
nor U11245 (N_11245,N_3227,N_5924);
or U11246 (N_11246,N_6106,N_533);
xnor U11247 (N_11247,N_2576,N_5977);
and U11248 (N_11248,N_2967,N_28);
nand U11249 (N_11249,N_116,N_1109);
nor U11250 (N_11250,N_358,N_2377);
or U11251 (N_11251,N_3973,N_55);
xnor U11252 (N_11252,N_2522,N_2454);
nor U11253 (N_11253,N_5212,N_743);
xnor U11254 (N_11254,N_3280,N_1930);
or U11255 (N_11255,N_6018,N_3496);
nand U11256 (N_11256,N_5058,N_3385);
or U11257 (N_11257,N_1391,N_2687);
nor U11258 (N_11258,N_5501,N_2833);
nand U11259 (N_11259,N_628,N_1378);
nor U11260 (N_11260,N_26,N_466);
and U11261 (N_11261,N_1224,N_6025);
xnor U11262 (N_11262,N_5592,N_4844);
nor U11263 (N_11263,N_3072,N_4645);
nand U11264 (N_11264,N_2476,N_5216);
nand U11265 (N_11265,N_3950,N_380);
nor U11266 (N_11266,N_6082,N_3481);
and U11267 (N_11267,N_328,N_5842);
and U11268 (N_11268,N_3227,N_3431);
and U11269 (N_11269,N_4593,N_1591);
or U11270 (N_11270,N_2885,N_6198);
xor U11271 (N_11271,N_4182,N_479);
nand U11272 (N_11272,N_4534,N_4414);
xor U11273 (N_11273,N_2292,N_3575);
nor U11274 (N_11274,N_5150,N_2902);
and U11275 (N_11275,N_5143,N_1075);
or U11276 (N_11276,N_5086,N_4767);
or U11277 (N_11277,N_4279,N_4183);
nor U11278 (N_11278,N_729,N_1852);
xor U11279 (N_11279,N_5962,N_4240);
and U11280 (N_11280,N_2929,N_4893);
nand U11281 (N_11281,N_39,N_4455);
xor U11282 (N_11282,N_3236,N_4474);
nand U11283 (N_11283,N_3063,N_2456);
and U11284 (N_11284,N_3503,N_1418);
and U11285 (N_11285,N_2382,N_3769);
xor U11286 (N_11286,N_463,N_204);
xor U11287 (N_11287,N_1691,N_5550);
xnor U11288 (N_11288,N_4821,N_2839);
and U11289 (N_11289,N_6090,N_2771);
and U11290 (N_11290,N_0,N_2374);
nor U11291 (N_11291,N_4741,N_5074);
and U11292 (N_11292,N_715,N_4015);
xnor U11293 (N_11293,N_1536,N_2428);
nor U11294 (N_11294,N_5570,N_2242);
nand U11295 (N_11295,N_5810,N_927);
xor U11296 (N_11296,N_3779,N_23);
xnor U11297 (N_11297,N_3643,N_1144);
and U11298 (N_11298,N_5244,N_4264);
nand U11299 (N_11299,N_6131,N_6116);
nor U11300 (N_11300,N_344,N_4720);
nor U11301 (N_11301,N_3038,N_3905);
xor U11302 (N_11302,N_2568,N_4647);
nand U11303 (N_11303,N_2,N_4452);
xnor U11304 (N_11304,N_5812,N_5538);
xor U11305 (N_11305,N_1075,N_1067);
nand U11306 (N_11306,N_3555,N_371);
nor U11307 (N_11307,N_1088,N_3592);
nor U11308 (N_11308,N_974,N_4898);
nor U11309 (N_11309,N_4857,N_3133);
or U11310 (N_11310,N_4895,N_5844);
or U11311 (N_11311,N_6216,N_2138);
nor U11312 (N_11312,N_157,N_1194);
and U11313 (N_11313,N_3932,N_2101);
or U11314 (N_11314,N_2053,N_4280);
and U11315 (N_11315,N_232,N_1676);
nand U11316 (N_11316,N_3413,N_5470);
xnor U11317 (N_11317,N_3116,N_4380);
or U11318 (N_11318,N_4545,N_4868);
nor U11319 (N_11319,N_3755,N_709);
nor U11320 (N_11320,N_2241,N_4848);
xor U11321 (N_11321,N_6174,N_590);
or U11322 (N_11322,N_2505,N_2750);
xor U11323 (N_11323,N_5125,N_4868);
or U11324 (N_11324,N_4353,N_4262);
and U11325 (N_11325,N_4589,N_3246);
xnor U11326 (N_11326,N_5861,N_3160);
or U11327 (N_11327,N_2429,N_5157);
nand U11328 (N_11328,N_3434,N_4218);
xnor U11329 (N_11329,N_5287,N_558);
and U11330 (N_11330,N_42,N_2207);
and U11331 (N_11331,N_2497,N_5136);
nor U11332 (N_11332,N_3875,N_1740);
nand U11333 (N_11333,N_5532,N_5088);
xor U11334 (N_11334,N_3205,N_261);
xor U11335 (N_11335,N_2540,N_6147);
xnor U11336 (N_11336,N_5643,N_5602);
nand U11337 (N_11337,N_1940,N_4200);
and U11338 (N_11338,N_4570,N_1094);
and U11339 (N_11339,N_206,N_4279);
nor U11340 (N_11340,N_6130,N_392);
or U11341 (N_11341,N_2623,N_6186);
and U11342 (N_11342,N_2532,N_5063);
nor U11343 (N_11343,N_4065,N_944);
and U11344 (N_11344,N_4016,N_5590);
or U11345 (N_11345,N_5820,N_972);
nand U11346 (N_11346,N_947,N_5490);
nand U11347 (N_11347,N_157,N_56);
and U11348 (N_11348,N_5390,N_377);
and U11349 (N_11349,N_3922,N_1934);
and U11350 (N_11350,N_3188,N_1316);
and U11351 (N_11351,N_1874,N_5660);
or U11352 (N_11352,N_2089,N_2505);
or U11353 (N_11353,N_1413,N_4414);
nor U11354 (N_11354,N_1583,N_1898);
nor U11355 (N_11355,N_2779,N_3970);
nor U11356 (N_11356,N_3056,N_3621);
xnor U11357 (N_11357,N_1419,N_1252);
and U11358 (N_11358,N_4683,N_2444);
xnor U11359 (N_11359,N_5041,N_5798);
and U11360 (N_11360,N_1736,N_4404);
nand U11361 (N_11361,N_2911,N_1904);
and U11362 (N_11362,N_26,N_5143);
and U11363 (N_11363,N_1619,N_5598);
and U11364 (N_11364,N_5676,N_2482);
or U11365 (N_11365,N_5959,N_5524);
and U11366 (N_11366,N_1519,N_827);
or U11367 (N_11367,N_4346,N_2421);
nor U11368 (N_11368,N_3680,N_5046);
and U11369 (N_11369,N_1826,N_5200);
xnor U11370 (N_11370,N_1418,N_4265);
nand U11371 (N_11371,N_3413,N_2352);
nor U11372 (N_11372,N_4475,N_566);
xnor U11373 (N_11373,N_529,N_2215);
and U11374 (N_11374,N_5784,N_1975);
and U11375 (N_11375,N_4722,N_2923);
or U11376 (N_11376,N_3254,N_4741);
and U11377 (N_11377,N_3041,N_1449);
and U11378 (N_11378,N_3971,N_4719);
or U11379 (N_11379,N_4664,N_3498);
xor U11380 (N_11380,N_4625,N_2184);
xnor U11381 (N_11381,N_3847,N_3536);
nor U11382 (N_11382,N_2560,N_3075);
xnor U11383 (N_11383,N_5030,N_5968);
xnor U11384 (N_11384,N_597,N_97);
nor U11385 (N_11385,N_4235,N_380);
and U11386 (N_11386,N_1250,N_189);
nand U11387 (N_11387,N_1206,N_5658);
or U11388 (N_11388,N_5181,N_4195);
or U11389 (N_11389,N_4341,N_5949);
nor U11390 (N_11390,N_227,N_4519);
and U11391 (N_11391,N_3859,N_2328);
nand U11392 (N_11392,N_5277,N_5202);
nand U11393 (N_11393,N_1471,N_6004);
nand U11394 (N_11394,N_3886,N_968);
and U11395 (N_11395,N_3751,N_3896);
or U11396 (N_11396,N_5842,N_5888);
xnor U11397 (N_11397,N_2909,N_3835);
or U11398 (N_11398,N_5183,N_5037);
xnor U11399 (N_11399,N_5729,N_5508);
nor U11400 (N_11400,N_2406,N_4295);
or U11401 (N_11401,N_3491,N_3356);
xnor U11402 (N_11402,N_4798,N_3677);
xnor U11403 (N_11403,N_2559,N_661);
nor U11404 (N_11404,N_6037,N_2473);
nor U11405 (N_11405,N_5382,N_2243);
and U11406 (N_11406,N_5532,N_4180);
nor U11407 (N_11407,N_448,N_4945);
nor U11408 (N_11408,N_4307,N_3989);
nor U11409 (N_11409,N_4168,N_2521);
xnor U11410 (N_11410,N_4746,N_944);
or U11411 (N_11411,N_1176,N_808);
and U11412 (N_11412,N_2359,N_5299);
xor U11413 (N_11413,N_2467,N_4638);
and U11414 (N_11414,N_5461,N_6005);
nand U11415 (N_11415,N_5144,N_1279);
or U11416 (N_11416,N_5262,N_5306);
nor U11417 (N_11417,N_3211,N_2238);
nor U11418 (N_11418,N_5951,N_4211);
nor U11419 (N_11419,N_3281,N_4525);
nand U11420 (N_11420,N_1587,N_5020);
nor U11421 (N_11421,N_4470,N_5799);
nand U11422 (N_11422,N_2872,N_553);
nand U11423 (N_11423,N_1723,N_1607);
or U11424 (N_11424,N_5033,N_3362);
nor U11425 (N_11425,N_5912,N_941);
nor U11426 (N_11426,N_1331,N_2026);
nor U11427 (N_11427,N_3387,N_5904);
nor U11428 (N_11428,N_840,N_4728);
and U11429 (N_11429,N_858,N_4358);
and U11430 (N_11430,N_1162,N_1283);
xnor U11431 (N_11431,N_321,N_6153);
and U11432 (N_11432,N_3515,N_6200);
nand U11433 (N_11433,N_4123,N_5668);
nand U11434 (N_11434,N_3843,N_965);
or U11435 (N_11435,N_2,N_4314);
or U11436 (N_11436,N_4877,N_2349);
or U11437 (N_11437,N_651,N_3701);
and U11438 (N_11438,N_866,N_1097);
and U11439 (N_11439,N_1906,N_6138);
nand U11440 (N_11440,N_2363,N_2478);
nand U11441 (N_11441,N_1529,N_3075);
nand U11442 (N_11442,N_583,N_5210);
nand U11443 (N_11443,N_4590,N_4139);
nand U11444 (N_11444,N_3062,N_1491);
nor U11445 (N_11445,N_2843,N_1368);
nor U11446 (N_11446,N_1040,N_312);
nor U11447 (N_11447,N_4416,N_426);
nand U11448 (N_11448,N_2239,N_5653);
nor U11449 (N_11449,N_1103,N_1979);
nand U11450 (N_11450,N_4579,N_2755);
xnor U11451 (N_11451,N_4742,N_3643);
nand U11452 (N_11452,N_462,N_2449);
xnor U11453 (N_11453,N_493,N_5201);
nor U11454 (N_11454,N_1735,N_5362);
and U11455 (N_11455,N_1453,N_674);
nand U11456 (N_11456,N_3817,N_4187);
or U11457 (N_11457,N_2144,N_1981);
nor U11458 (N_11458,N_5856,N_981);
nor U11459 (N_11459,N_4173,N_5617);
nor U11460 (N_11460,N_4866,N_1022);
nor U11461 (N_11461,N_3582,N_300);
or U11462 (N_11462,N_1888,N_2054);
or U11463 (N_11463,N_3746,N_734);
or U11464 (N_11464,N_4484,N_3589);
and U11465 (N_11465,N_1242,N_73);
xnor U11466 (N_11466,N_2851,N_3006);
nor U11467 (N_11467,N_4030,N_565);
nor U11468 (N_11468,N_5499,N_4962);
nand U11469 (N_11469,N_2170,N_2210);
xnor U11470 (N_11470,N_6059,N_5326);
or U11471 (N_11471,N_800,N_2011);
xor U11472 (N_11472,N_2950,N_4401);
and U11473 (N_11473,N_2905,N_4237);
or U11474 (N_11474,N_1580,N_3290);
or U11475 (N_11475,N_744,N_4064);
or U11476 (N_11476,N_2437,N_1338);
or U11477 (N_11477,N_1068,N_6084);
nor U11478 (N_11478,N_3274,N_349);
and U11479 (N_11479,N_5855,N_2451);
nor U11480 (N_11480,N_358,N_5666);
and U11481 (N_11481,N_2431,N_2099);
xnor U11482 (N_11482,N_3624,N_1129);
or U11483 (N_11483,N_3696,N_558);
xnor U11484 (N_11484,N_5443,N_1032);
or U11485 (N_11485,N_4897,N_2909);
or U11486 (N_11486,N_4897,N_834);
or U11487 (N_11487,N_2776,N_89);
nand U11488 (N_11488,N_2339,N_4905);
nand U11489 (N_11489,N_2054,N_2925);
and U11490 (N_11490,N_5927,N_3195);
or U11491 (N_11491,N_6049,N_4184);
and U11492 (N_11492,N_4974,N_2191);
or U11493 (N_11493,N_3789,N_5301);
nand U11494 (N_11494,N_2488,N_4133);
or U11495 (N_11495,N_190,N_5725);
or U11496 (N_11496,N_1717,N_737);
nand U11497 (N_11497,N_498,N_450);
nor U11498 (N_11498,N_5028,N_6);
nand U11499 (N_11499,N_5143,N_25);
xor U11500 (N_11500,N_6186,N_867);
and U11501 (N_11501,N_6016,N_2287);
xnor U11502 (N_11502,N_614,N_3780);
or U11503 (N_11503,N_169,N_4814);
xnor U11504 (N_11504,N_1833,N_3922);
nor U11505 (N_11505,N_1863,N_2054);
nor U11506 (N_11506,N_6097,N_4192);
nor U11507 (N_11507,N_5909,N_454);
nand U11508 (N_11508,N_1369,N_3433);
or U11509 (N_11509,N_640,N_429);
xnor U11510 (N_11510,N_624,N_2551);
nand U11511 (N_11511,N_3678,N_5767);
xor U11512 (N_11512,N_6153,N_225);
nor U11513 (N_11513,N_3963,N_3678);
and U11514 (N_11514,N_1841,N_3560);
or U11515 (N_11515,N_3028,N_2502);
or U11516 (N_11516,N_760,N_2203);
nand U11517 (N_11517,N_2784,N_1711);
and U11518 (N_11518,N_3705,N_5326);
or U11519 (N_11519,N_3475,N_1588);
or U11520 (N_11520,N_5651,N_6171);
and U11521 (N_11521,N_2579,N_3697);
and U11522 (N_11522,N_5668,N_441);
and U11523 (N_11523,N_3364,N_23);
nor U11524 (N_11524,N_2559,N_4226);
xor U11525 (N_11525,N_2963,N_2680);
nand U11526 (N_11526,N_4606,N_2389);
and U11527 (N_11527,N_1718,N_1867);
nor U11528 (N_11528,N_4582,N_389);
nand U11529 (N_11529,N_3411,N_5833);
nor U11530 (N_11530,N_4312,N_2853);
or U11531 (N_11531,N_1943,N_4599);
xor U11532 (N_11532,N_5299,N_4224);
xor U11533 (N_11533,N_5222,N_783);
xnor U11534 (N_11534,N_2446,N_2857);
and U11535 (N_11535,N_6148,N_446);
and U11536 (N_11536,N_1112,N_6222);
or U11537 (N_11537,N_3047,N_5086);
or U11538 (N_11538,N_3091,N_4732);
or U11539 (N_11539,N_1414,N_2721);
nand U11540 (N_11540,N_942,N_5080);
xnor U11541 (N_11541,N_4572,N_429);
xnor U11542 (N_11542,N_4786,N_885);
nand U11543 (N_11543,N_2402,N_4930);
or U11544 (N_11544,N_4426,N_2049);
xnor U11545 (N_11545,N_939,N_5472);
xor U11546 (N_11546,N_878,N_3078);
and U11547 (N_11547,N_1425,N_539);
nor U11548 (N_11548,N_3944,N_359);
or U11549 (N_11549,N_2468,N_377);
or U11550 (N_11550,N_4979,N_1263);
nor U11551 (N_11551,N_4337,N_1270);
nand U11552 (N_11552,N_1973,N_4290);
nand U11553 (N_11553,N_2969,N_3045);
xor U11554 (N_11554,N_2195,N_3247);
and U11555 (N_11555,N_362,N_310);
nand U11556 (N_11556,N_5517,N_2667);
or U11557 (N_11557,N_4873,N_1444);
xnor U11558 (N_11558,N_5440,N_3735);
or U11559 (N_11559,N_4140,N_2416);
or U11560 (N_11560,N_4975,N_4264);
xnor U11561 (N_11561,N_258,N_2595);
or U11562 (N_11562,N_5997,N_1039);
nand U11563 (N_11563,N_664,N_4597);
xor U11564 (N_11564,N_4912,N_4909);
and U11565 (N_11565,N_2725,N_4481);
nor U11566 (N_11566,N_584,N_5166);
xor U11567 (N_11567,N_3216,N_3258);
or U11568 (N_11568,N_1132,N_1556);
and U11569 (N_11569,N_1091,N_3316);
and U11570 (N_11570,N_5158,N_2501);
and U11571 (N_11571,N_2710,N_3451);
nor U11572 (N_11572,N_1031,N_3477);
nand U11573 (N_11573,N_2897,N_5902);
and U11574 (N_11574,N_420,N_4127);
and U11575 (N_11575,N_2791,N_2026);
and U11576 (N_11576,N_4915,N_4144);
and U11577 (N_11577,N_1242,N_4658);
or U11578 (N_11578,N_2940,N_5391);
nand U11579 (N_11579,N_648,N_6118);
or U11580 (N_11580,N_1671,N_1097);
nor U11581 (N_11581,N_4586,N_478);
nor U11582 (N_11582,N_5929,N_531);
and U11583 (N_11583,N_5335,N_2731);
nand U11584 (N_11584,N_1743,N_2593);
nor U11585 (N_11585,N_4005,N_1994);
and U11586 (N_11586,N_2511,N_5576);
nand U11587 (N_11587,N_5635,N_160);
nand U11588 (N_11588,N_5061,N_5400);
nor U11589 (N_11589,N_1191,N_208);
nor U11590 (N_11590,N_4460,N_4038);
or U11591 (N_11591,N_1559,N_1414);
nand U11592 (N_11592,N_5894,N_0);
or U11593 (N_11593,N_3917,N_1199);
nor U11594 (N_11594,N_6062,N_329);
nand U11595 (N_11595,N_5015,N_4578);
xnor U11596 (N_11596,N_5021,N_1237);
and U11597 (N_11597,N_1478,N_1654);
nor U11598 (N_11598,N_5359,N_1233);
or U11599 (N_11599,N_4445,N_3687);
xor U11600 (N_11600,N_3694,N_3490);
nand U11601 (N_11601,N_3021,N_3856);
and U11602 (N_11602,N_1732,N_3317);
nand U11603 (N_11603,N_3763,N_3023);
nor U11604 (N_11604,N_4760,N_1176);
nor U11605 (N_11605,N_4186,N_4543);
or U11606 (N_11606,N_2943,N_3089);
or U11607 (N_11607,N_822,N_4135);
nand U11608 (N_11608,N_3575,N_4212);
xor U11609 (N_11609,N_2503,N_66);
nor U11610 (N_11610,N_413,N_330);
nand U11611 (N_11611,N_2142,N_2796);
nand U11612 (N_11612,N_5964,N_884);
and U11613 (N_11613,N_6109,N_3123);
or U11614 (N_11614,N_3967,N_1184);
and U11615 (N_11615,N_298,N_4558);
and U11616 (N_11616,N_5092,N_439);
or U11617 (N_11617,N_6185,N_1832);
nand U11618 (N_11618,N_1230,N_1186);
and U11619 (N_11619,N_3208,N_4126);
or U11620 (N_11620,N_4232,N_138);
or U11621 (N_11621,N_5495,N_5945);
nor U11622 (N_11622,N_3684,N_1625);
and U11623 (N_11623,N_239,N_5961);
nand U11624 (N_11624,N_3904,N_1932);
nand U11625 (N_11625,N_812,N_3198);
and U11626 (N_11626,N_1847,N_1617);
and U11627 (N_11627,N_5727,N_6172);
or U11628 (N_11628,N_590,N_3029);
nand U11629 (N_11629,N_5418,N_3128);
nand U11630 (N_11630,N_5866,N_4903);
nand U11631 (N_11631,N_3873,N_2324);
and U11632 (N_11632,N_57,N_115);
or U11633 (N_11633,N_4046,N_1942);
xor U11634 (N_11634,N_1513,N_4194);
and U11635 (N_11635,N_5526,N_3811);
xor U11636 (N_11636,N_1233,N_4275);
xnor U11637 (N_11637,N_4117,N_3460);
and U11638 (N_11638,N_6066,N_5500);
nand U11639 (N_11639,N_1269,N_4445);
nand U11640 (N_11640,N_2538,N_1803);
nand U11641 (N_11641,N_4991,N_1194);
nor U11642 (N_11642,N_1261,N_5792);
xor U11643 (N_11643,N_2886,N_691);
nand U11644 (N_11644,N_667,N_1347);
or U11645 (N_11645,N_4329,N_3981);
or U11646 (N_11646,N_4133,N_230);
nor U11647 (N_11647,N_3487,N_5988);
nand U11648 (N_11648,N_2285,N_572);
or U11649 (N_11649,N_3961,N_4461);
nor U11650 (N_11650,N_3406,N_1430);
nor U11651 (N_11651,N_2964,N_5078);
nand U11652 (N_11652,N_2898,N_89);
and U11653 (N_11653,N_523,N_4816);
xor U11654 (N_11654,N_3323,N_2712);
nor U11655 (N_11655,N_3762,N_178);
or U11656 (N_11656,N_2939,N_3517);
nand U11657 (N_11657,N_1816,N_821);
nor U11658 (N_11658,N_5915,N_105);
nand U11659 (N_11659,N_3719,N_1517);
or U11660 (N_11660,N_2941,N_4808);
and U11661 (N_11661,N_6152,N_2684);
and U11662 (N_11662,N_4206,N_774);
nand U11663 (N_11663,N_3086,N_5119);
nand U11664 (N_11664,N_4789,N_3310);
nor U11665 (N_11665,N_250,N_5474);
xor U11666 (N_11666,N_6012,N_2934);
or U11667 (N_11667,N_3955,N_3716);
nor U11668 (N_11668,N_5013,N_4682);
and U11669 (N_11669,N_4675,N_3822);
nor U11670 (N_11670,N_959,N_5954);
xor U11671 (N_11671,N_2727,N_575);
and U11672 (N_11672,N_4076,N_3857);
nor U11673 (N_11673,N_3079,N_5759);
nor U11674 (N_11674,N_5052,N_399);
xnor U11675 (N_11675,N_4981,N_6176);
xor U11676 (N_11676,N_5194,N_6244);
nor U11677 (N_11677,N_2870,N_5098);
xor U11678 (N_11678,N_436,N_4623);
and U11679 (N_11679,N_1228,N_2737);
xnor U11680 (N_11680,N_5287,N_2777);
nand U11681 (N_11681,N_1480,N_1261);
nand U11682 (N_11682,N_2019,N_2439);
or U11683 (N_11683,N_1164,N_2628);
and U11684 (N_11684,N_3345,N_3885);
nand U11685 (N_11685,N_2792,N_532);
nor U11686 (N_11686,N_1968,N_2903);
nand U11687 (N_11687,N_38,N_3460);
and U11688 (N_11688,N_2143,N_6037);
nor U11689 (N_11689,N_4038,N_3319);
and U11690 (N_11690,N_5623,N_2794);
or U11691 (N_11691,N_3119,N_4440);
and U11692 (N_11692,N_2299,N_2759);
xor U11693 (N_11693,N_2360,N_4576);
nand U11694 (N_11694,N_2517,N_1854);
and U11695 (N_11695,N_2374,N_1020);
xor U11696 (N_11696,N_3718,N_965);
or U11697 (N_11697,N_4613,N_1151);
nand U11698 (N_11698,N_4422,N_4327);
nor U11699 (N_11699,N_863,N_1389);
nor U11700 (N_11700,N_3369,N_765);
nor U11701 (N_11701,N_4353,N_3516);
or U11702 (N_11702,N_3406,N_2583);
nand U11703 (N_11703,N_3857,N_155);
or U11704 (N_11704,N_5609,N_5739);
nor U11705 (N_11705,N_272,N_3235);
and U11706 (N_11706,N_3030,N_3373);
or U11707 (N_11707,N_2944,N_3260);
nand U11708 (N_11708,N_3163,N_601);
xor U11709 (N_11709,N_1816,N_3249);
xor U11710 (N_11710,N_345,N_4145);
nand U11711 (N_11711,N_6229,N_1811);
or U11712 (N_11712,N_2640,N_378);
xnor U11713 (N_11713,N_3528,N_2334);
nor U11714 (N_11714,N_2699,N_3958);
xor U11715 (N_11715,N_338,N_6227);
nand U11716 (N_11716,N_3913,N_4603);
and U11717 (N_11717,N_2953,N_3678);
and U11718 (N_11718,N_624,N_3384);
or U11719 (N_11719,N_1949,N_1450);
nand U11720 (N_11720,N_3103,N_2006);
and U11721 (N_11721,N_3690,N_3197);
and U11722 (N_11722,N_6245,N_1133);
nor U11723 (N_11723,N_3874,N_704);
xnor U11724 (N_11724,N_5907,N_3204);
or U11725 (N_11725,N_294,N_40);
xnor U11726 (N_11726,N_9,N_2536);
nand U11727 (N_11727,N_517,N_4787);
xnor U11728 (N_11728,N_2298,N_4240);
or U11729 (N_11729,N_1205,N_4801);
and U11730 (N_11730,N_5903,N_5708);
or U11731 (N_11731,N_1428,N_3481);
nand U11732 (N_11732,N_1646,N_3885);
nand U11733 (N_11733,N_5434,N_5101);
and U11734 (N_11734,N_5040,N_3572);
or U11735 (N_11735,N_6158,N_5324);
nand U11736 (N_11736,N_5820,N_5373);
xnor U11737 (N_11737,N_4405,N_6063);
and U11738 (N_11738,N_3957,N_5527);
nand U11739 (N_11739,N_1049,N_3437);
nand U11740 (N_11740,N_3311,N_241);
xnor U11741 (N_11741,N_3763,N_3401);
and U11742 (N_11742,N_2149,N_1495);
or U11743 (N_11743,N_5617,N_1577);
nand U11744 (N_11744,N_2004,N_4782);
xor U11745 (N_11745,N_4107,N_5941);
nor U11746 (N_11746,N_1227,N_2595);
nand U11747 (N_11747,N_131,N_3586);
nor U11748 (N_11748,N_606,N_3803);
xnor U11749 (N_11749,N_3540,N_2366);
nand U11750 (N_11750,N_2668,N_2967);
nand U11751 (N_11751,N_4803,N_3927);
or U11752 (N_11752,N_4148,N_2648);
xor U11753 (N_11753,N_809,N_4412);
nand U11754 (N_11754,N_4395,N_1773);
and U11755 (N_11755,N_2209,N_4617);
xor U11756 (N_11756,N_2346,N_1931);
nor U11757 (N_11757,N_1592,N_995);
and U11758 (N_11758,N_5602,N_5579);
and U11759 (N_11759,N_663,N_6047);
xnor U11760 (N_11760,N_3872,N_3827);
nand U11761 (N_11761,N_36,N_1737);
xor U11762 (N_11762,N_471,N_4072);
xor U11763 (N_11763,N_5075,N_3730);
xor U11764 (N_11764,N_4072,N_1818);
xnor U11765 (N_11765,N_5134,N_2198);
nand U11766 (N_11766,N_443,N_3746);
nor U11767 (N_11767,N_4546,N_773);
xor U11768 (N_11768,N_701,N_1494);
nor U11769 (N_11769,N_5912,N_713);
nor U11770 (N_11770,N_3924,N_5890);
nand U11771 (N_11771,N_1936,N_2281);
nand U11772 (N_11772,N_4047,N_5415);
nand U11773 (N_11773,N_4070,N_1678);
nor U11774 (N_11774,N_4371,N_5968);
and U11775 (N_11775,N_369,N_4991);
or U11776 (N_11776,N_2998,N_6046);
nand U11777 (N_11777,N_1211,N_307);
xnor U11778 (N_11778,N_4004,N_4486);
nand U11779 (N_11779,N_4829,N_5759);
nor U11780 (N_11780,N_4296,N_4093);
xor U11781 (N_11781,N_5945,N_5295);
and U11782 (N_11782,N_2117,N_3534);
nor U11783 (N_11783,N_4539,N_2976);
xnor U11784 (N_11784,N_1865,N_2176);
and U11785 (N_11785,N_887,N_3700);
nor U11786 (N_11786,N_3285,N_4405);
nor U11787 (N_11787,N_3365,N_5123);
nor U11788 (N_11788,N_4566,N_1815);
nor U11789 (N_11789,N_6040,N_803);
nor U11790 (N_11790,N_5020,N_5164);
and U11791 (N_11791,N_5172,N_654);
and U11792 (N_11792,N_6119,N_2201);
xnor U11793 (N_11793,N_1326,N_1433);
xnor U11794 (N_11794,N_4513,N_4951);
and U11795 (N_11795,N_3795,N_708);
and U11796 (N_11796,N_4541,N_3060);
nand U11797 (N_11797,N_4316,N_3741);
nor U11798 (N_11798,N_5703,N_5941);
nor U11799 (N_11799,N_4621,N_2683);
nor U11800 (N_11800,N_2208,N_1210);
nor U11801 (N_11801,N_3138,N_1414);
nor U11802 (N_11802,N_1818,N_4335);
xor U11803 (N_11803,N_4143,N_2431);
or U11804 (N_11804,N_1019,N_816);
nor U11805 (N_11805,N_5868,N_3730);
nor U11806 (N_11806,N_5586,N_5942);
and U11807 (N_11807,N_191,N_4727);
xnor U11808 (N_11808,N_4173,N_648);
and U11809 (N_11809,N_6121,N_2876);
and U11810 (N_11810,N_1743,N_5973);
xor U11811 (N_11811,N_3285,N_5254);
xor U11812 (N_11812,N_1095,N_4199);
nor U11813 (N_11813,N_2736,N_5304);
and U11814 (N_11814,N_5004,N_4649);
nor U11815 (N_11815,N_5523,N_2589);
nor U11816 (N_11816,N_4200,N_3384);
nor U11817 (N_11817,N_5657,N_3517);
nand U11818 (N_11818,N_3265,N_5990);
and U11819 (N_11819,N_504,N_919);
nand U11820 (N_11820,N_789,N_2377);
xnor U11821 (N_11821,N_5354,N_1345);
nand U11822 (N_11822,N_3537,N_742);
nand U11823 (N_11823,N_1605,N_5801);
nor U11824 (N_11824,N_4593,N_5256);
nor U11825 (N_11825,N_1159,N_732);
or U11826 (N_11826,N_5703,N_2134);
nor U11827 (N_11827,N_31,N_2408);
and U11828 (N_11828,N_5444,N_3163);
or U11829 (N_11829,N_4659,N_242);
and U11830 (N_11830,N_3711,N_3222);
nor U11831 (N_11831,N_907,N_5528);
xnor U11832 (N_11832,N_2856,N_2797);
or U11833 (N_11833,N_4400,N_260);
or U11834 (N_11834,N_659,N_325);
xor U11835 (N_11835,N_3991,N_5058);
nand U11836 (N_11836,N_1940,N_5322);
nor U11837 (N_11837,N_5002,N_712);
nand U11838 (N_11838,N_4422,N_3048);
and U11839 (N_11839,N_3250,N_799);
nor U11840 (N_11840,N_2172,N_3370);
and U11841 (N_11841,N_5905,N_4065);
nor U11842 (N_11842,N_4272,N_1736);
nor U11843 (N_11843,N_6026,N_110);
nand U11844 (N_11844,N_3726,N_2246);
xor U11845 (N_11845,N_4326,N_174);
and U11846 (N_11846,N_534,N_5868);
nor U11847 (N_11847,N_3098,N_5371);
or U11848 (N_11848,N_2586,N_608);
or U11849 (N_11849,N_3528,N_2045);
xnor U11850 (N_11850,N_350,N_978);
and U11851 (N_11851,N_2940,N_2266);
and U11852 (N_11852,N_3254,N_3019);
and U11853 (N_11853,N_3226,N_954);
and U11854 (N_11854,N_4954,N_2811);
nand U11855 (N_11855,N_1976,N_2706);
nand U11856 (N_11856,N_5684,N_6012);
xor U11857 (N_11857,N_3184,N_418);
nand U11858 (N_11858,N_5082,N_1260);
nand U11859 (N_11859,N_5769,N_2806);
xnor U11860 (N_11860,N_4215,N_5696);
nor U11861 (N_11861,N_280,N_1223);
nand U11862 (N_11862,N_4044,N_5115);
xor U11863 (N_11863,N_6102,N_4342);
nor U11864 (N_11864,N_4933,N_4821);
nand U11865 (N_11865,N_3662,N_5607);
and U11866 (N_11866,N_5024,N_3260);
or U11867 (N_11867,N_1302,N_4823);
nor U11868 (N_11868,N_716,N_6220);
nand U11869 (N_11869,N_5573,N_1599);
nand U11870 (N_11870,N_3225,N_4946);
or U11871 (N_11871,N_5325,N_2909);
xnor U11872 (N_11872,N_2360,N_4544);
or U11873 (N_11873,N_4090,N_1776);
xnor U11874 (N_11874,N_3414,N_5401);
or U11875 (N_11875,N_2728,N_3442);
xnor U11876 (N_11876,N_5189,N_2159);
xor U11877 (N_11877,N_233,N_515);
xnor U11878 (N_11878,N_1304,N_6228);
xor U11879 (N_11879,N_1846,N_5535);
or U11880 (N_11880,N_2277,N_3119);
nand U11881 (N_11881,N_4040,N_5495);
nand U11882 (N_11882,N_1570,N_5043);
nor U11883 (N_11883,N_3165,N_2979);
xor U11884 (N_11884,N_6228,N_206);
xnor U11885 (N_11885,N_4160,N_3096);
xor U11886 (N_11886,N_1176,N_3835);
or U11887 (N_11887,N_249,N_1385);
nand U11888 (N_11888,N_5555,N_709);
xnor U11889 (N_11889,N_786,N_4291);
nor U11890 (N_11890,N_282,N_2288);
xor U11891 (N_11891,N_2487,N_3001);
nor U11892 (N_11892,N_1232,N_4589);
and U11893 (N_11893,N_1383,N_5765);
or U11894 (N_11894,N_4494,N_6228);
xnor U11895 (N_11895,N_4646,N_1065);
and U11896 (N_11896,N_5937,N_4576);
and U11897 (N_11897,N_5741,N_800);
xnor U11898 (N_11898,N_2171,N_5580);
nand U11899 (N_11899,N_1883,N_2409);
and U11900 (N_11900,N_2694,N_5011);
nand U11901 (N_11901,N_5934,N_3722);
nand U11902 (N_11902,N_1232,N_499);
xnor U11903 (N_11903,N_3194,N_4904);
and U11904 (N_11904,N_990,N_3929);
xnor U11905 (N_11905,N_5534,N_400);
nand U11906 (N_11906,N_4464,N_1616);
and U11907 (N_11907,N_6137,N_540);
and U11908 (N_11908,N_4683,N_4014);
and U11909 (N_11909,N_2908,N_1629);
or U11910 (N_11910,N_511,N_5445);
and U11911 (N_11911,N_2246,N_2596);
and U11912 (N_11912,N_865,N_2272);
or U11913 (N_11913,N_5272,N_3850);
xnor U11914 (N_11914,N_2569,N_2103);
and U11915 (N_11915,N_4846,N_6066);
nand U11916 (N_11916,N_1818,N_3866);
or U11917 (N_11917,N_458,N_3952);
nand U11918 (N_11918,N_3767,N_1507);
and U11919 (N_11919,N_3767,N_3726);
nand U11920 (N_11920,N_5269,N_5318);
nand U11921 (N_11921,N_4136,N_3525);
xnor U11922 (N_11922,N_2224,N_3173);
nand U11923 (N_11923,N_5559,N_2474);
or U11924 (N_11924,N_1013,N_3334);
and U11925 (N_11925,N_3417,N_1640);
and U11926 (N_11926,N_4541,N_3551);
or U11927 (N_11927,N_3962,N_2823);
or U11928 (N_11928,N_6063,N_5332);
and U11929 (N_11929,N_4345,N_5961);
nor U11930 (N_11930,N_4023,N_2038);
or U11931 (N_11931,N_5552,N_867);
or U11932 (N_11932,N_5915,N_6008);
nor U11933 (N_11933,N_5516,N_1453);
and U11934 (N_11934,N_4001,N_984);
and U11935 (N_11935,N_4158,N_5467);
nor U11936 (N_11936,N_2385,N_1450);
xor U11937 (N_11937,N_418,N_5914);
or U11938 (N_11938,N_5899,N_3772);
nor U11939 (N_11939,N_1200,N_5941);
or U11940 (N_11940,N_4143,N_1091);
nand U11941 (N_11941,N_5666,N_1665);
or U11942 (N_11942,N_1256,N_5718);
and U11943 (N_11943,N_3218,N_5584);
nor U11944 (N_11944,N_6065,N_3142);
xnor U11945 (N_11945,N_3840,N_3576);
nor U11946 (N_11946,N_407,N_2372);
or U11947 (N_11947,N_2302,N_1340);
and U11948 (N_11948,N_3975,N_3611);
nor U11949 (N_11949,N_914,N_4929);
nor U11950 (N_11950,N_59,N_3928);
xor U11951 (N_11951,N_632,N_1498);
or U11952 (N_11952,N_2237,N_2971);
nand U11953 (N_11953,N_6184,N_4294);
nand U11954 (N_11954,N_1745,N_4273);
and U11955 (N_11955,N_1022,N_1268);
and U11956 (N_11956,N_408,N_701);
nand U11957 (N_11957,N_1256,N_2660);
and U11958 (N_11958,N_4408,N_4366);
or U11959 (N_11959,N_5080,N_350);
xor U11960 (N_11960,N_3924,N_5920);
or U11961 (N_11961,N_4773,N_3716);
nand U11962 (N_11962,N_3850,N_5903);
and U11963 (N_11963,N_2357,N_799);
xnor U11964 (N_11964,N_2965,N_5896);
xor U11965 (N_11965,N_1445,N_5540);
nor U11966 (N_11966,N_1909,N_5551);
or U11967 (N_11967,N_4812,N_799);
nand U11968 (N_11968,N_2457,N_5310);
and U11969 (N_11969,N_6116,N_5826);
nor U11970 (N_11970,N_3368,N_4639);
or U11971 (N_11971,N_6016,N_2122);
and U11972 (N_11972,N_4559,N_1224);
and U11973 (N_11973,N_2565,N_721);
or U11974 (N_11974,N_2254,N_4572);
and U11975 (N_11975,N_3436,N_3417);
or U11976 (N_11976,N_3983,N_2712);
nand U11977 (N_11977,N_5027,N_1773);
or U11978 (N_11978,N_4770,N_4914);
xnor U11979 (N_11979,N_5668,N_943);
and U11980 (N_11980,N_1195,N_808);
and U11981 (N_11981,N_2468,N_6080);
nand U11982 (N_11982,N_2932,N_752);
nor U11983 (N_11983,N_144,N_1365);
nor U11984 (N_11984,N_5400,N_1314);
nor U11985 (N_11985,N_5183,N_1136);
nor U11986 (N_11986,N_82,N_5425);
and U11987 (N_11987,N_1334,N_2300);
xor U11988 (N_11988,N_992,N_1632);
xnor U11989 (N_11989,N_4759,N_709);
xnor U11990 (N_11990,N_284,N_3831);
or U11991 (N_11991,N_5537,N_891);
or U11992 (N_11992,N_551,N_4746);
nor U11993 (N_11993,N_3962,N_3139);
xnor U11994 (N_11994,N_2000,N_3616);
nor U11995 (N_11995,N_1021,N_1320);
xor U11996 (N_11996,N_2205,N_5848);
xnor U11997 (N_11997,N_2948,N_4703);
nand U11998 (N_11998,N_2997,N_5157);
or U11999 (N_11999,N_1015,N_6095);
and U12000 (N_12000,N_414,N_4318);
nor U12001 (N_12001,N_1721,N_884);
and U12002 (N_12002,N_6212,N_2941);
or U12003 (N_12003,N_4828,N_6102);
or U12004 (N_12004,N_1982,N_2084);
nand U12005 (N_12005,N_1858,N_3308);
nand U12006 (N_12006,N_5158,N_2927);
and U12007 (N_12007,N_750,N_1921);
nor U12008 (N_12008,N_1570,N_3164);
nor U12009 (N_12009,N_941,N_3749);
nand U12010 (N_12010,N_1383,N_5690);
and U12011 (N_12011,N_5664,N_5354);
or U12012 (N_12012,N_6040,N_2617);
and U12013 (N_12013,N_5790,N_2966);
nand U12014 (N_12014,N_646,N_717);
nor U12015 (N_12015,N_5539,N_1042);
nand U12016 (N_12016,N_5994,N_3689);
xnor U12017 (N_12017,N_4937,N_442);
nor U12018 (N_12018,N_1078,N_2576);
or U12019 (N_12019,N_22,N_1646);
nand U12020 (N_12020,N_441,N_4142);
nor U12021 (N_12021,N_3606,N_5185);
nand U12022 (N_12022,N_1373,N_5859);
and U12023 (N_12023,N_3040,N_2072);
and U12024 (N_12024,N_3145,N_1523);
nor U12025 (N_12025,N_371,N_3561);
nor U12026 (N_12026,N_2917,N_4502);
or U12027 (N_12027,N_3718,N_4171);
nor U12028 (N_12028,N_1607,N_689);
and U12029 (N_12029,N_1355,N_1715);
nor U12030 (N_12030,N_4889,N_1655);
nor U12031 (N_12031,N_2779,N_5747);
xor U12032 (N_12032,N_4392,N_1746);
xor U12033 (N_12033,N_321,N_2896);
nand U12034 (N_12034,N_3282,N_5057);
xnor U12035 (N_12035,N_3238,N_4566);
xor U12036 (N_12036,N_4797,N_6098);
xor U12037 (N_12037,N_6238,N_3865);
nand U12038 (N_12038,N_793,N_5449);
xor U12039 (N_12039,N_3082,N_4492);
and U12040 (N_12040,N_307,N_4882);
xnor U12041 (N_12041,N_76,N_3213);
and U12042 (N_12042,N_4734,N_5183);
or U12043 (N_12043,N_1352,N_1821);
nor U12044 (N_12044,N_4673,N_5300);
xnor U12045 (N_12045,N_2697,N_5278);
and U12046 (N_12046,N_1547,N_1781);
xor U12047 (N_12047,N_5223,N_5595);
nor U12048 (N_12048,N_1630,N_2237);
or U12049 (N_12049,N_817,N_1731);
xor U12050 (N_12050,N_2462,N_1069);
and U12051 (N_12051,N_1574,N_4688);
and U12052 (N_12052,N_2080,N_4930);
or U12053 (N_12053,N_2585,N_5970);
nand U12054 (N_12054,N_6195,N_5968);
or U12055 (N_12055,N_3255,N_5817);
xor U12056 (N_12056,N_2451,N_2533);
xnor U12057 (N_12057,N_19,N_1157);
nor U12058 (N_12058,N_6221,N_6186);
xnor U12059 (N_12059,N_3916,N_4146);
xor U12060 (N_12060,N_1818,N_3258);
nor U12061 (N_12061,N_278,N_628);
xor U12062 (N_12062,N_2486,N_561);
nor U12063 (N_12063,N_5930,N_3866);
and U12064 (N_12064,N_1754,N_3186);
nor U12065 (N_12065,N_4495,N_639);
nand U12066 (N_12066,N_3340,N_5964);
or U12067 (N_12067,N_1076,N_4429);
nor U12068 (N_12068,N_4094,N_268);
nand U12069 (N_12069,N_3248,N_1749);
nor U12070 (N_12070,N_2117,N_1176);
and U12071 (N_12071,N_62,N_4136);
xor U12072 (N_12072,N_41,N_4239);
or U12073 (N_12073,N_1463,N_4699);
nand U12074 (N_12074,N_2158,N_5209);
and U12075 (N_12075,N_467,N_6017);
and U12076 (N_12076,N_2455,N_1969);
or U12077 (N_12077,N_1518,N_522);
xor U12078 (N_12078,N_2423,N_1663);
or U12079 (N_12079,N_3235,N_5136);
nor U12080 (N_12080,N_1914,N_5149);
and U12081 (N_12081,N_4842,N_370);
and U12082 (N_12082,N_3663,N_459);
and U12083 (N_12083,N_3960,N_5230);
nand U12084 (N_12084,N_2996,N_5241);
nor U12085 (N_12085,N_203,N_136);
xor U12086 (N_12086,N_5085,N_4058);
or U12087 (N_12087,N_4727,N_2179);
nor U12088 (N_12088,N_237,N_5965);
xnor U12089 (N_12089,N_5155,N_4741);
nand U12090 (N_12090,N_3557,N_5796);
nand U12091 (N_12091,N_6211,N_219);
nand U12092 (N_12092,N_5105,N_4677);
nand U12093 (N_12093,N_4664,N_4351);
or U12094 (N_12094,N_719,N_780);
xnor U12095 (N_12095,N_5807,N_3595);
xor U12096 (N_12096,N_379,N_4938);
nor U12097 (N_12097,N_3903,N_2799);
nor U12098 (N_12098,N_5997,N_637);
or U12099 (N_12099,N_1173,N_6012);
xnor U12100 (N_12100,N_5481,N_2696);
nor U12101 (N_12101,N_3866,N_5266);
and U12102 (N_12102,N_830,N_112);
nor U12103 (N_12103,N_4705,N_2157);
xor U12104 (N_12104,N_5023,N_2551);
or U12105 (N_12105,N_4987,N_2669);
nand U12106 (N_12106,N_6007,N_6136);
nor U12107 (N_12107,N_2628,N_1649);
nand U12108 (N_12108,N_5590,N_3077);
or U12109 (N_12109,N_1489,N_1068);
nor U12110 (N_12110,N_3638,N_6033);
nand U12111 (N_12111,N_3342,N_3095);
and U12112 (N_12112,N_1518,N_4731);
or U12113 (N_12113,N_3299,N_4215);
xor U12114 (N_12114,N_2103,N_5574);
nand U12115 (N_12115,N_5441,N_4320);
nand U12116 (N_12116,N_5632,N_4917);
nand U12117 (N_12117,N_3804,N_1110);
or U12118 (N_12118,N_1066,N_3897);
xnor U12119 (N_12119,N_4595,N_1620);
nand U12120 (N_12120,N_4170,N_1320);
nand U12121 (N_12121,N_5090,N_2612);
nor U12122 (N_12122,N_4059,N_5924);
xor U12123 (N_12123,N_2690,N_2759);
and U12124 (N_12124,N_2895,N_4749);
and U12125 (N_12125,N_3260,N_901);
nor U12126 (N_12126,N_1065,N_791);
xor U12127 (N_12127,N_1378,N_3200);
or U12128 (N_12128,N_804,N_68);
and U12129 (N_12129,N_4170,N_4122);
nand U12130 (N_12130,N_2115,N_5703);
nor U12131 (N_12131,N_1436,N_5990);
nor U12132 (N_12132,N_4761,N_5991);
nand U12133 (N_12133,N_2371,N_2429);
or U12134 (N_12134,N_2080,N_314);
or U12135 (N_12135,N_5060,N_783);
or U12136 (N_12136,N_2727,N_889);
nor U12137 (N_12137,N_6179,N_2748);
xnor U12138 (N_12138,N_3806,N_3365);
and U12139 (N_12139,N_3385,N_6053);
xnor U12140 (N_12140,N_5882,N_4147);
nor U12141 (N_12141,N_4106,N_5620);
nor U12142 (N_12142,N_1202,N_2461);
or U12143 (N_12143,N_1130,N_5622);
and U12144 (N_12144,N_1935,N_5625);
and U12145 (N_12145,N_4153,N_1639);
nand U12146 (N_12146,N_2085,N_1663);
nor U12147 (N_12147,N_3780,N_5593);
nor U12148 (N_12148,N_4356,N_956);
nor U12149 (N_12149,N_3449,N_4274);
or U12150 (N_12150,N_5815,N_21);
nor U12151 (N_12151,N_4512,N_3354);
nand U12152 (N_12152,N_3078,N_6190);
or U12153 (N_12153,N_731,N_5117);
nor U12154 (N_12154,N_1225,N_257);
xnor U12155 (N_12155,N_2782,N_2351);
nand U12156 (N_12156,N_3921,N_3729);
or U12157 (N_12157,N_6173,N_1190);
nand U12158 (N_12158,N_2683,N_644);
nand U12159 (N_12159,N_4983,N_3358);
and U12160 (N_12160,N_2653,N_4464);
and U12161 (N_12161,N_6150,N_1264);
nor U12162 (N_12162,N_1337,N_3720);
nor U12163 (N_12163,N_1833,N_1707);
nor U12164 (N_12164,N_101,N_2557);
nor U12165 (N_12165,N_4832,N_5205);
nand U12166 (N_12166,N_2424,N_832);
or U12167 (N_12167,N_1788,N_1162);
xor U12168 (N_12168,N_1116,N_975);
nand U12169 (N_12169,N_5298,N_2297);
and U12170 (N_12170,N_3250,N_3295);
nand U12171 (N_12171,N_1194,N_3877);
nor U12172 (N_12172,N_758,N_4265);
nor U12173 (N_12173,N_5454,N_5476);
nand U12174 (N_12174,N_3080,N_5049);
and U12175 (N_12175,N_5523,N_3839);
and U12176 (N_12176,N_5532,N_3734);
xor U12177 (N_12177,N_1267,N_1705);
nor U12178 (N_12178,N_4007,N_2570);
nor U12179 (N_12179,N_2140,N_1513);
and U12180 (N_12180,N_3006,N_69);
nand U12181 (N_12181,N_245,N_4432);
and U12182 (N_12182,N_4217,N_1953);
nand U12183 (N_12183,N_2827,N_1793);
nand U12184 (N_12184,N_4671,N_3985);
or U12185 (N_12185,N_4003,N_103);
and U12186 (N_12186,N_4529,N_4157);
nand U12187 (N_12187,N_4118,N_6153);
and U12188 (N_12188,N_5665,N_1239);
and U12189 (N_12189,N_1989,N_3423);
or U12190 (N_12190,N_5580,N_881);
xnor U12191 (N_12191,N_1982,N_5949);
and U12192 (N_12192,N_3020,N_6039);
xor U12193 (N_12193,N_3678,N_1607);
nand U12194 (N_12194,N_5351,N_2743);
and U12195 (N_12195,N_1539,N_1837);
xor U12196 (N_12196,N_1945,N_4125);
and U12197 (N_12197,N_912,N_984);
xnor U12198 (N_12198,N_3499,N_3468);
nor U12199 (N_12199,N_1697,N_1104);
xnor U12200 (N_12200,N_5804,N_4864);
or U12201 (N_12201,N_1237,N_5446);
nand U12202 (N_12202,N_3185,N_1786);
and U12203 (N_12203,N_1845,N_2759);
nor U12204 (N_12204,N_5095,N_2246);
xnor U12205 (N_12205,N_5472,N_6241);
or U12206 (N_12206,N_5756,N_3521);
and U12207 (N_12207,N_6166,N_5552);
nor U12208 (N_12208,N_5823,N_976);
and U12209 (N_12209,N_2778,N_875);
nor U12210 (N_12210,N_5825,N_5230);
nor U12211 (N_12211,N_132,N_2099);
and U12212 (N_12212,N_2055,N_338);
xor U12213 (N_12213,N_1981,N_2201);
or U12214 (N_12214,N_3784,N_5126);
and U12215 (N_12215,N_897,N_760);
nand U12216 (N_12216,N_3283,N_3044);
nand U12217 (N_12217,N_4900,N_676);
or U12218 (N_12218,N_2973,N_4048);
and U12219 (N_12219,N_2666,N_5451);
nor U12220 (N_12220,N_5050,N_5778);
and U12221 (N_12221,N_3957,N_4544);
or U12222 (N_12222,N_3207,N_1462);
nand U12223 (N_12223,N_3790,N_5113);
and U12224 (N_12224,N_2602,N_2367);
or U12225 (N_12225,N_3106,N_4723);
xnor U12226 (N_12226,N_3538,N_1466);
nand U12227 (N_12227,N_3759,N_552);
xnor U12228 (N_12228,N_3133,N_2199);
or U12229 (N_12229,N_2232,N_2973);
xnor U12230 (N_12230,N_3505,N_3705);
and U12231 (N_12231,N_4300,N_4504);
xor U12232 (N_12232,N_5977,N_4148);
nor U12233 (N_12233,N_5505,N_3716);
nor U12234 (N_12234,N_2148,N_3865);
and U12235 (N_12235,N_3595,N_665);
and U12236 (N_12236,N_4423,N_6130);
and U12237 (N_12237,N_3580,N_4674);
nand U12238 (N_12238,N_851,N_2170);
and U12239 (N_12239,N_5735,N_1215);
and U12240 (N_12240,N_978,N_1440);
nand U12241 (N_12241,N_2215,N_2259);
nand U12242 (N_12242,N_2151,N_6095);
or U12243 (N_12243,N_923,N_5953);
nand U12244 (N_12244,N_3600,N_905);
or U12245 (N_12245,N_4184,N_4079);
and U12246 (N_12246,N_2551,N_6038);
and U12247 (N_12247,N_5008,N_722);
nor U12248 (N_12248,N_4933,N_1911);
and U12249 (N_12249,N_3165,N_4720);
nor U12250 (N_12250,N_2938,N_5076);
nand U12251 (N_12251,N_3385,N_6039);
or U12252 (N_12252,N_5353,N_4106);
nand U12253 (N_12253,N_103,N_1794);
and U12254 (N_12254,N_5638,N_3716);
or U12255 (N_12255,N_1904,N_4231);
and U12256 (N_12256,N_3320,N_137);
or U12257 (N_12257,N_6230,N_3987);
xor U12258 (N_12258,N_429,N_2174);
xnor U12259 (N_12259,N_6106,N_1551);
nand U12260 (N_12260,N_2359,N_4815);
nor U12261 (N_12261,N_2219,N_5519);
and U12262 (N_12262,N_1275,N_4627);
nand U12263 (N_12263,N_1226,N_5763);
nor U12264 (N_12264,N_3949,N_1350);
or U12265 (N_12265,N_5528,N_910);
nor U12266 (N_12266,N_5815,N_2905);
xnor U12267 (N_12267,N_1509,N_3682);
or U12268 (N_12268,N_5796,N_6022);
nor U12269 (N_12269,N_2232,N_4826);
or U12270 (N_12270,N_4407,N_3787);
nand U12271 (N_12271,N_2282,N_3943);
nand U12272 (N_12272,N_5779,N_415);
nand U12273 (N_12273,N_2902,N_436);
xnor U12274 (N_12274,N_156,N_2393);
nand U12275 (N_12275,N_936,N_3319);
or U12276 (N_12276,N_3404,N_4200);
or U12277 (N_12277,N_3433,N_2851);
xnor U12278 (N_12278,N_1918,N_5716);
nor U12279 (N_12279,N_1420,N_1921);
nand U12280 (N_12280,N_4415,N_4608);
nand U12281 (N_12281,N_3170,N_4871);
nor U12282 (N_12282,N_522,N_3814);
or U12283 (N_12283,N_2841,N_5154);
and U12284 (N_12284,N_1191,N_745);
xor U12285 (N_12285,N_4298,N_5906);
xor U12286 (N_12286,N_5660,N_3145);
or U12287 (N_12287,N_4582,N_1884);
or U12288 (N_12288,N_887,N_2848);
and U12289 (N_12289,N_4590,N_4624);
nor U12290 (N_12290,N_652,N_4675);
xor U12291 (N_12291,N_473,N_4365);
nand U12292 (N_12292,N_2300,N_4018);
or U12293 (N_12293,N_4571,N_3042);
or U12294 (N_12294,N_3288,N_1004);
xor U12295 (N_12295,N_939,N_3672);
nor U12296 (N_12296,N_1480,N_6023);
nand U12297 (N_12297,N_4911,N_3638);
nor U12298 (N_12298,N_1257,N_3889);
xnor U12299 (N_12299,N_2305,N_1504);
nand U12300 (N_12300,N_1930,N_2240);
xnor U12301 (N_12301,N_4629,N_4900);
xnor U12302 (N_12302,N_3964,N_4567);
nor U12303 (N_12303,N_1858,N_4750);
and U12304 (N_12304,N_4445,N_159);
xnor U12305 (N_12305,N_2724,N_1412);
nand U12306 (N_12306,N_5417,N_4038);
nand U12307 (N_12307,N_4207,N_1061);
xnor U12308 (N_12308,N_2555,N_3894);
or U12309 (N_12309,N_2975,N_3121);
and U12310 (N_12310,N_5282,N_5347);
nor U12311 (N_12311,N_4108,N_2884);
nor U12312 (N_12312,N_3888,N_752);
xor U12313 (N_12313,N_2625,N_4245);
nor U12314 (N_12314,N_3702,N_651);
xor U12315 (N_12315,N_5596,N_6067);
xor U12316 (N_12316,N_4329,N_1155);
xnor U12317 (N_12317,N_5207,N_5301);
and U12318 (N_12318,N_1960,N_1794);
nor U12319 (N_12319,N_5238,N_4160);
and U12320 (N_12320,N_5848,N_3430);
or U12321 (N_12321,N_6158,N_3065);
xor U12322 (N_12322,N_1109,N_1331);
nand U12323 (N_12323,N_2749,N_5759);
nor U12324 (N_12324,N_5324,N_3734);
nand U12325 (N_12325,N_1233,N_6024);
xor U12326 (N_12326,N_759,N_2695);
nand U12327 (N_12327,N_2723,N_640);
nor U12328 (N_12328,N_4426,N_2679);
nand U12329 (N_12329,N_6098,N_3498);
nor U12330 (N_12330,N_5897,N_5542);
nor U12331 (N_12331,N_5769,N_3990);
or U12332 (N_12332,N_5368,N_3489);
and U12333 (N_12333,N_3348,N_1635);
and U12334 (N_12334,N_1693,N_4413);
nor U12335 (N_12335,N_3289,N_5299);
nor U12336 (N_12336,N_1054,N_2977);
or U12337 (N_12337,N_1026,N_5160);
or U12338 (N_12338,N_3807,N_4748);
nor U12339 (N_12339,N_2632,N_6060);
xor U12340 (N_12340,N_4238,N_2083);
nand U12341 (N_12341,N_3436,N_220);
and U12342 (N_12342,N_4555,N_5438);
or U12343 (N_12343,N_1704,N_4780);
or U12344 (N_12344,N_2088,N_5712);
nand U12345 (N_12345,N_3226,N_832);
nand U12346 (N_12346,N_2644,N_5369);
or U12347 (N_12347,N_3136,N_5670);
nand U12348 (N_12348,N_3637,N_3930);
or U12349 (N_12349,N_3270,N_687);
nand U12350 (N_12350,N_149,N_4910);
xor U12351 (N_12351,N_558,N_5661);
nand U12352 (N_12352,N_3874,N_4181);
nor U12353 (N_12353,N_549,N_6033);
xnor U12354 (N_12354,N_1080,N_3140);
xnor U12355 (N_12355,N_3614,N_105);
nand U12356 (N_12356,N_2949,N_3284);
xor U12357 (N_12357,N_405,N_1024);
and U12358 (N_12358,N_1318,N_2982);
or U12359 (N_12359,N_4933,N_1858);
or U12360 (N_12360,N_1065,N_2018);
or U12361 (N_12361,N_3768,N_3446);
and U12362 (N_12362,N_2488,N_565);
xor U12363 (N_12363,N_44,N_3442);
nand U12364 (N_12364,N_3591,N_2318);
nand U12365 (N_12365,N_3578,N_2157);
or U12366 (N_12366,N_190,N_1293);
or U12367 (N_12367,N_2433,N_1685);
xor U12368 (N_12368,N_5772,N_861);
nand U12369 (N_12369,N_6099,N_2709);
and U12370 (N_12370,N_3573,N_1483);
nand U12371 (N_12371,N_5815,N_3339);
xnor U12372 (N_12372,N_2348,N_4039);
and U12373 (N_12373,N_1843,N_3972);
and U12374 (N_12374,N_2135,N_2530);
nor U12375 (N_12375,N_5060,N_4863);
nand U12376 (N_12376,N_5429,N_4383);
and U12377 (N_12377,N_855,N_1775);
xor U12378 (N_12378,N_3293,N_711);
or U12379 (N_12379,N_3042,N_5336);
xnor U12380 (N_12380,N_4878,N_2581);
nand U12381 (N_12381,N_5192,N_1040);
and U12382 (N_12382,N_4472,N_1498);
xnor U12383 (N_12383,N_1763,N_5661);
nor U12384 (N_12384,N_5940,N_3017);
xor U12385 (N_12385,N_3556,N_4004);
or U12386 (N_12386,N_4737,N_5392);
nand U12387 (N_12387,N_3135,N_3394);
or U12388 (N_12388,N_2409,N_5434);
and U12389 (N_12389,N_2326,N_1623);
nand U12390 (N_12390,N_1944,N_4399);
nor U12391 (N_12391,N_3289,N_356);
nor U12392 (N_12392,N_4806,N_430);
xnor U12393 (N_12393,N_4976,N_3527);
or U12394 (N_12394,N_997,N_2814);
and U12395 (N_12395,N_1429,N_4317);
or U12396 (N_12396,N_477,N_4649);
and U12397 (N_12397,N_4894,N_458);
nor U12398 (N_12398,N_310,N_471);
nor U12399 (N_12399,N_4888,N_1738);
nand U12400 (N_12400,N_6179,N_1637);
and U12401 (N_12401,N_1924,N_3336);
or U12402 (N_12402,N_1734,N_4927);
nand U12403 (N_12403,N_2572,N_4888);
xnor U12404 (N_12404,N_5327,N_5771);
or U12405 (N_12405,N_2574,N_365);
and U12406 (N_12406,N_3821,N_2938);
nor U12407 (N_12407,N_4490,N_6217);
and U12408 (N_12408,N_3333,N_6040);
xnor U12409 (N_12409,N_620,N_4643);
nor U12410 (N_12410,N_2510,N_5049);
or U12411 (N_12411,N_5959,N_5940);
and U12412 (N_12412,N_2222,N_3654);
and U12413 (N_12413,N_2009,N_323);
and U12414 (N_12414,N_4479,N_1086);
and U12415 (N_12415,N_5016,N_4644);
xnor U12416 (N_12416,N_2361,N_817);
and U12417 (N_12417,N_2057,N_4890);
nor U12418 (N_12418,N_1783,N_3366);
xor U12419 (N_12419,N_1415,N_2063);
or U12420 (N_12420,N_1225,N_3921);
nor U12421 (N_12421,N_4097,N_5772);
or U12422 (N_12422,N_425,N_969);
and U12423 (N_12423,N_4603,N_211);
or U12424 (N_12424,N_1453,N_4202);
and U12425 (N_12425,N_3191,N_3288);
and U12426 (N_12426,N_5067,N_5153);
and U12427 (N_12427,N_4419,N_223);
nand U12428 (N_12428,N_129,N_4212);
nand U12429 (N_12429,N_4173,N_2578);
or U12430 (N_12430,N_2574,N_2286);
and U12431 (N_12431,N_3354,N_5);
and U12432 (N_12432,N_6135,N_5757);
and U12433 (N_12433,N_2050,N_4765);
and U12434 (N_12434,N_1854,N_6148);
and U12435 (N_12435,N_4544,N_1813);
nand U12436 (N_12436,N_1924,N_1323);
nor U12437 (N_12437,N_3598,N_4652);
and U12438 (N_12438,N_3477,N_3539);
and U12439 (N_12439,N_5157,N_4260);
nor U12440 (N_12440,N_4959,N_5199);
and U12441 (N_12441,N_3923,N_5830);
nor U12442 (N_12442,N_2287,N_1233);
xnor U12443 (N_12443,N_4077,N_1738);
or U12444 (N_12444,N_699,N_133);
xnor U12445 (N_12445,N_4044,N_5073);
nand U12446 (N_12446,N_5315,N_3723);
or U12447 (N_12447,N_1017,N_412);
nor U12448 (N_12448,N_763,N_6024);
nor U12449 (N_12449,N_1005,N_2195);
or U12450 (N_12450,N_1079,N_795);
nor U12451 (N_12451,N_40,N_2047);
and U12452 (N_12452,N_2796,N_2461);
xor U12453 (N_12453,N_1210,N_3711);
nand U12454 (N_12454,N_1178,N_5670);
xor U12455 (N_12455,N_4096,N_4422);
and U12456 (N_12456,N_2875,N_338);
xnor U12457 (N_12457,N_225,N_5951);
nor U12458 (N_12458,N_4849,N_96);
nor U12459 (N_12459,N_2977,N_1615);
nand U12460 (N_12460,N_1645,N_5363);
or U12461 (N_12461,N_2435,N_1109);
and U12462 (N_12462,N_302,N_3915);
or U12463 (N_12463,N_26,N_2952);
and U12464 (N_12464,N_4528,N_3363);
and U12465 (N_12465,N_4890,N_5478);
nand U12466 (N_12466,N_3190,N_2807);
nor U12467 (N_12467,N_2419,N_2786);
xnor U12468 (N_12468,N_802,N_3563);
xnor U12469 (N_12469,N_3213,N_1891);
xnor U12470 (N_12470,N_4791,N_4596);
nor U12471 (N_12471,N_5148,N_5951);
and U12472 (N_12472,N_4324,N_1514);
nor U12473 (N_12473,N_2999,N_4497);
or U12474 (N_12474,N_2266,N_1681);
and U12475 (N_12475,N_503,N_1839);
nor U12476 (N_12476,N_2358,N_3554);
and U12477 (N_12477,N_3515,N_6062);
and U12478 (N_12478,N_6228,N_4905);
nand U12479 (N_12479,N_1568,N_2762);
and U12480 (N_12480,N_3825,N_795);
nand U12481 (N_12481,N_1563,N_508);
nor U12482 (N_12482,N_4675,N_3189);
nor U12483 (N_12483,N_799,N_1915);
or U12484 (N_12484,N_1191,N_4103);
and U12485 (N_12485,N_5179,N_5628);
nor U12486 (N_12486,N_2788,N_5161);
xnor U12487 (N_12487,N_3779,N_2330);
and U12488 (N_12488,N_4592,N_3025);
or U12489 (N_12489,N_108,N_6194);
and U12490 (N_12490,N_2501,N_6242);
or U12491 (N_12491,N_4951,N_85);
nand U12492 (N_12492,N_5174,N_3651);
nor U12493 (N_12493,N_3963,N_3207);
and U12494 (N_12494,N_5499,N_5862);
or U12495 (N_12495,N_4006,N_3144);
nor U12496 (N_12496,N_3837,N_4996);
nor U12497 (N_12497,N_1657,N_3928);
nand U12498 (N_12498,N_2483,N_1371);
nor U12499 (N_12499,N_5381,N_6219);
and U12500 (N_12500,N_10533,N_7323);
xnor U12501 (N_12501,N_11157,N_6696);
nor U12502 (N_12502,N_6965,N_8881);
or U12503 (N_12503,N_6959,N_7946);
nand U12504 (N_12504,N_9806,N_10670);
and U12505 (N_12505,N_8802,N_6885);
xnor U12506 (N_12506,N_8819,N_9769);
and U12507 (N_12507,N_11198,N_11541);
xnor U12508 (N_12508,N_10038,N_11059);
nor U12509 (N_12509,N_7704,N_7809);
and U12510 (N_12510,N_8124,N_6344);
and U12511 (N_12511,N_12275,N_12442);
nor U12512 (N_12512,N_11588,N_8277);
xor U12513 (N_12513,N_8414,N_8483);
xnor U12514 (N_12514,N_12139,N_6391);
nand U12515 (N_12515,N_11595,N_6454);
nor U12516 (N_12516,N_8168,N_9008);
nand U12517 (N_12517,N_8425,N_9719);
or U12518 (N_12518,N_12174,N_7249);
nand U12519 (N_12519,N_6772,N_9510);
xor U12520 (N_12520,N_10053,N_9032);
and U12521 (N_12521,N_8194,N_9748);
nor U12522 (N_12522,N_7676,N_9613);
nor U12523 (N_12523,N_6252,N_8803);
nor U12524 (N_12524,N_9069,N_11174);
nor U12525 (N_12525,N_9044,N_10994);
nand U12526 (N_12526,N_10530,N_9373);
and U12527 (N_12527,N_6783,N_11448);
xnor U12528 (N_12528,N_7525,N_11737);
nor U12529 (N_12529,N_8261,N_8291);
xor U12530 (N_12530,N_9565,N_9118);
nor U12531 (N_12531,N_7534,N_7682);
nand U12532 (N_12532,N_7816,N_11450);
xnor U12533 (N_12533,N_6397,N_11455);
xor U12534 (N_12534,N_6628,N_8929);
nor U12535 (N_12535,N_7983,N_10421);
nor U12536 (N_12536,N_8914,N_8569);
or U12537 (N_12537,N_11214,N_7545);
nand U12538 (N_12538,N_7931,N_10817);
nor U12539 (N_12539,N_7032,N_10506);
nand U12540 (N_12540,N_10606,N_8820);
and U12541 (N_12541,N_11547,N_7009);
nor U12542 (N_12542,N_9013,N_8413);
and U12543 (N_12543,N_9509,N_9796);
xnor U12544 (N_12544,N_8830,N_8645);
xor U12545 (N_12545,N_10652,N_9205);
xnor U12546 (N_12546,N_9910,N_10678);
nor U12547 (N_12547,N_10525,N_7184);
nor U12548 (N_12548,N_7125,N_10934);
xnor U12549 (N_12549,N_8763,N_8231);
and U12550 (N_12550,N_9786,N_6732);
nor U12551 (N_12551,N_8922,N_7936);
nor U12552 (N_12552,N_7537,N_11856);
nand U12553 (N_12553,N_7478,N_12039);
or U12554 (N_12554,N_9855,N_11335);
or U12555 (N_12555,N_9371,N_9107);
or U12556 (N_12556,N_11596,N_9632);
xnor U12557 (N_12557,N_10997,N_7105);
or U12558 (N_12558,N_9676,N_7022);
nor U12559 (N_12559,N_6301,N_10328);
xor U12560 (N_12560,N_7396,N_7647);
or U12561 (N_12561,N_10033,N_10389);
or U12562 (N_12562,N_9864,N_10473);
and U12563 (N_12563,N_7775,N_7577);
or U12564 (N_12564,N_11289,N_11216);
and U12565 (N_12565,N_6509,N_10518);
nand U12566 (N_12566,N_9805,N_9122);
xor U12567 (N_12567,N_10206,N_9985);
nand U12568 (N_12568,N_11070,N_10432);
and U12569 (N_12569,N_8462,N_12083);
and U12570 (N_12570,N_6986,N_11623);
or U12571 (N_12571,N_6283,N_12263);
or U12572 (N_12572,N_11614,N_8675);
xor U12573 (N_12573,N_11250,N_11167);
xor U12574 (N_12574,N_9182,N_6313);
nor U12575 (N_12575,N_6690,N_9502);
nand U12576 (N_12576,N_10594,N_11805);
or U12577 (N_12577,N_10509,N_11435);
or U12578 (N_12578,N_8834,N_11468);
and U12579 (N_12579,N_8682,N_12409);
xor U12580 (N_12580,N_9185,N_12448);
nand U12581 (N_12581,N_8740,N_6616);
and U12582 (N_12582,N_12484,N_12181);
xnor U12583 (N_12583,N_9701,N_11625);
and U12584 (N_12584,N_10927,N_12305);
xnor U12585 (N_12585,N_11437,N_7455);
nor U12586 (N_12586,N_7390,N_11754);
or U12587 (N_12587,N_11561,N_7239);
nand U12588 (N_12588,N_11039,N_11146);
and U12589 (N_12589,N_6861,N_8476);
and U12590 (N_12590,N_7302,N_12410);
nor U12591 (N_12591,N_8321,N_11814);
nor U12592 (N_12592,N_7089,N_12301);
and U12593 (N_12593,N_12488,N_11620);
nand U12594 (N_12594,N_11855,N_6493);
xor U12595 (N_12595,N_12408,N_11551);
nor U12596 (N_12596,N_9096,N_10369);
and U12597 (N_12597,N_9698,N_10885);
nand U12598 (N_12598,N_7793,N_9285);
and U12599 (N_12599,N_9359,N_8971);
nor U12600 (N_12600,N_7864,N_10460);
or U12601 (N_12601,N_8618,N_8005);
or U12602 (N_12602,N_11822,N_7643);
nor U12603 (N_12603,N_9619,N_8885);
or U12604 (N_12604,N_9920,N_10668);
nand U12605 (N_12605,N_12180,N_12001);
nand U12606 (N_12606,N_10596,N_10469);
nor U12607 (N_12607,N_6892,N_8771);
nand U12608 (N_12608,N_11131,N_8388);
nand U12609 (N_12609,N_10781,N_12045);
nand U12610 (N_12610,N_9184,N_11439);
or U12611 (N_12611,N_12162,N_11702);
nand U12612 (N_12612,N_10950,N_11274);
xor U12613 (N_12613,N_8353,N_6770);
nor U12614 (N_12614,N_7938,N_6864);
xor U12615 (N_12615,N_12102,N_7261);
nand U12616 (N_12616,N_10118,N_7941);
and U12617 (N_12617,N_7772,N_6284);
xor U12618 (N_12618,N_6365,N_8292);
nor U12619 (N_12619,N_7335,N_7144);
or U12620 (N_12620,N_12251,N_8192);
and U12621 (N_12621,N_7586,N_12179);
or U12622 (N_12622,N_6671,N_8322);
or U12623 (N_12623,N_7722,N_9942);
nand U12624 (N_12624,N_7994,N_12229);
nand U12625 (N_12625,N_12043,N_7221);
nand U12626 (N_12626,N_8006,N_12034);
or U12627 (N_12627,N_9423,N_11647);
nand U12628 (N_12628,N_9897,N_8375);
nor U12629 (N_12629,N_11441,N_8597);
xnor U12630 (N_12630,N_8259,N_10434);
nor U12631 (N_12631,N_7966,N_11655);
or U12632 (N_12632,N_11391,N_11612);
and U12633 (N_12633,N_7115,N_9955);
and U12634 (N_12634,N_10822,N_8826);
and U12635 (N_12635,N_9350,N_12441);
xnor U12636 (N_12636,N_7606,N_9007);
nand U12637 (N_12637,N_6253,N_9014);
nand U12638 (N_12638,N_6439,N_6479);
and U12639 (N_12639,N_9021,N_8519);
nor U12640 (N_12640,N_12461,N_8017);
nand U12641 (N_12641,N_7924,N_11063);
nor U12642 (N_12642,N_9574,N_10836);
and U12643 (N_12643,N_9583,N_10746);
nand U12644 (N_12644,N_8447,N_6495);
nand U12645 (N_12645,N_7686,N_8766);
nand U12646 (N_12646,N_7053,N_11918);
or U12647 (N_12647,N_8793,N_9011);
or U12648 (N_12648,N_9568,N_10635);
nand U12649 (N_12649,N_6514,N_10188);
xor U12650 (N_12650,N_9468,N_10039);
and U12651 (N_12651,N_10381,N_10189);
or U12652 (N_12652,N_6570,N_11905);
xnor U12653 (N_12653,N_6502,N_9586);
nand U12654 (N_12654,N_8683,N_8145);
nand U12655 (N_12655,N_12165,N_6682);
nand U12656 (N_12656,N_8021,N_11247);
or U12657 (N_12657,N_6600,N_6491);
and U12658 (N_12658,N_12021,N_7120);
or U12659 (N_12659,N_9344,N_10121);
or U12660 (N_12660,N_10797,N_8348);
xor U12661 (N_12661,N_9252,N_10623);
xnor U12662 (N_12662,N_7193,N_7055);
and U12663 (N_12663,N_6565,N_6273);
xor U12664 (N_12664,N_6335,N_6982);
nand U12665 (N_12665,N_6842,N_8454);
or U12666 (N_12666,N_7145,N_8711);
xnor U12667 (N_12667,N_10562,N_7490);
nand U12668 (N_12668,N_12027,N_10640);
xor U12669 (N_12669,N_10650,N_7067);
or U12670 (N_12670,N_9690,N_6715);
or U12671 (N_12671,N_11601,N_7202);
and U12672 (N_12672,N_10195,N_6809);
or U12673 (N_12673,N_9085,N_12363);
nand U12674 (N_12674,N_7524,N_6890);
or U12675 (N_12675,N_7395,N_9041);
xnor U12676 (N_12676,N_9139,N_11637);
or U12677 (N_12677,N_8373,N_8916);
xnor U12678 (N_12678,N_10583,N_11333);
nand U12679 (N_12679,N_6943,N_7020);
xnor U12680 (N_12680,N_6310,N_8727);
xnor U12681 (N_12681,N_8574,N_6623);
nor U12682 (N_12682,N_8724,N_8909);
nor U12683 (N_12683,N_6458,N_11538);
and U12684 (N_12684,N_10007,N_6779);
or U12685 (N_12685,N_10366,N_6680);
nor U12686 (N_12686,N_7191,N_9120);
and U12687 (N_12687,N_9869,N_9656);
or U12688 (N_12688,N_7319,N_8043);
or U12689 (N_12689,N_6385,N_9442);
and U12690 (N_12690,N_11325,N_6968);
xor U12691 (N_12691,N_10327,N_7712);
xnor U12692 (N_12692,N_9707,N_8113);
nand U12693 (N_12693,N_8081,N_12481);
nor U12694 (N_12694,N_6771,N_9800);
or U12695 (N_12695,N_12085,N_12469);
and U12696 (N_12696,N_8242,N_11715);
and U12697 (N_12697,N_9333,N_8190);
nand U12698 (N_12698,N_11338,N_10549);
or U12699 (N_12699,N_6728,N_10160);
nand U12700 (N_12700,N_9183,N_6289);
nand U12701 (N_12701,N_10021,N_11978);
nor U12702 (N_12702,N_8309,N_6387);
or U12703 (N_12703,N_10920,N_8792);
nor U12704 (N_12704,N_9461,N_6701);
or U12705 (N_12705,N_8632,N_9075);
or U12706 (N_12706,N_9347,N_9628);
nor U12707 (N_12707,N_6932,N_6359);
nand U12708 (N_12708,N_11374,N_9729);
or U12709 (N_12709,N_8137,N_10248);
or U12710 (N_12710,N_7497,N_11149);
nand U12711 (N_12711,N_9982,N_7522);
nand U12712 (N_12712,N_9038,N_7101);
nor U12713 (N_12713,N_11898,N_8274);
nor U12714 (N_12714,N_10896,N_9064);
xnor U12715 (N_12715,N_8888,N_9732);
or U12716 (N_12716,N_12244,N_6622);
or U12717 (N_12717,N_12345,N_6572);
and U12718 (N_12718,N_12022,N_6427);
nand U12719 (N_12719,N_9659,N_9703);
nand U12720 (N_12720,N_6720,N_9541);
xor U12721 (N_12721,N_6931,N_12192);
xor U12722 (N_12722,N_8823,N_9464);
or U12723 (N_12723,N_10575,N_7386);
and U12724 (N_12724,N_6567,N_11944);
or U12725 (N_12725,N_11550,N_7219);
nand U12726 (N_12726,N_8558,N_7849);
or U12727 (N_12727,N_8047,N_11979);
and U12728 (N_12728,N_7199,N_7257);
and U12729 (N_12729,N_9123,N_8620);
nand U12730 (N_12730,N_10490,N_8244);
xor U12731 (N_12731,N_8526,N_7458);
or U12732 (N_12732,N_10236,N_10353);
and U12733 (N_12733,N_10048,N_11150);
nor U12734 (N_12734,N_12234,N_11380);
and U12735 (N_12735,N_9970,N_11475);
nand U12736 (N_12736,N_6433,N_9481);
or U12737 (N_12737,N_12097,N_11718);
nand U12738 (N_12738,N_10253,N_9888);
and U12739 (N_12739,N_11183,N_10524);
or U12740 (N_12740,N_11611,N_8955);
xor U12741 (N_12741,N_9759,N_7289);
xor U12742 (N_12742,N_9266,N_7167);
and U12743 (N_12743,N_10799,N_6883);
nor U12744 (N_12744,N_8540,N_7540);
nor U12745 (N_12745,N_11656,N_7563);
nand U12746 (N_12746,N_11602,N_8845);
xnor U12747 (N_12747,N_6549,N_8427);
xnor U12748 (N_12748,N_6803,N_11329);
or U12749 (N_12749,N_9956,N_12321);
nand U12750 (N_12750,N_10698,N_11563);
nand U12751 (N_12751,N_10537,N_6738);
nor U12752 (N_12752,N_10361,N_6517);
nand U12753 (N_12753,N_6536,N_12205);
nor U12754 (N_12754,N_9989,N_9938);
nor U12755 (N_12755,N_12155,N_7488);
nor U12756 (N_12756,N_10061,N_8302);
or U12757 (N_12757,N_8416,N_10618);
or U12758 (N_12758,N_11094,N_8410);
nand U12759 (N_12759,N_10436,N_10829);
or U12760 (N_12760,N_9820,N_12443);
or U12761 (N_12761,N_11303,N_8831);
nor U12762 (N_12762,N_9638,N_7685);
and U12763 (N_12763,N_12052,N_9620);
xor U12764 (N_12764,N_7697,N_9900);
and U12765 (N_12765,N_8223,N_8110);
nand U12766 (N_12766,N_11082,N_10265);
nand U12767 (N_12767,N_8617,N_8814);
nand U12768 (N_12768,N_11050,N_6666);
or U12769 (N_12769,N_11580,N_8652);
xor U12770 (N_12770,N_9952,N_12067);
or U12771 (N_12771,N_8077,N_11461);
xor U12772 (N_12772,N_11415,N_7254);
and U12773 (N_12773,N_6322,N_8149);
and U12774 (N_12774,N_7515,N_11690);
xnor U12775 (N_12775,N_12452,N_10914);
nor U12776 (N_12776,N_9054,N_9336);
nor U12777 (N_12777,N_8878,N_9931);
nand U12778 (N_12778,N_7887,N_7436);
xnor U12779 (N_12779,N_10086,N_7517);
xor U12780 (N_12780,N_7131,N_11113);
nand U12781 (N_12781,N_9181,N_8835);
and U12782 (N_12782,N_9968,N_11949);
or U12783 (N_12783,N_10755,N_6657);
and U12784 (N_12784,N_6469,N_7664);
xnor U12785 (N_12785,N_10382,N_10619);
or U12786 (N_12786,N_7495,N_6956);
and U12787 (N_12787,N_11316,N_6800);
nor U12788 (N_12788,N_9368,N_8797);
xor U12789 (N_12789,N_7281,N_9207);
nand U12790 (N_12790,N_8440,N_11969);
or U12791 (N_12791,N_11554,N_11011);
nor U12792 (N_12792,N_7350,N_10256);
or U12793 (N_12793,N_7801,N_11252);
and U12794 (N_12794,N_6286,N_9080);
xnor U12795 (N_12795,N_11662,N_11869);
and U12796 (N_12796,N_6569,N_12421);
nor U12797 (N_12797,N_7449,N_7207);
nor U12798 (N_12798,N_6297,N_9849);
and U12799 (N_12799,N_10729,N_12336);
and U12800 (N_12800,N_8240,N_10901);
xor U12801 (N_12801,N_8537,N_9046);
or U12802 (N_12802,N_10002,N_6768);
or U12803 (N_12803,N_11189,N_7627);
and U12804 (N_12804,N_10093,N_10324);
nand U12805 (N_12805,N_6936,N_7619);
nor U12806 (N_12806,N_7729,N_10115);
nand U12807 (N_12807,N_11140,N_11743);
and U12808 (N_12808,N_8418,N_9886);
xnor U12809 (N_12809,N_8160,N_10461);
or U12810 (N_12810,N_8560,N_8721);
nor U12811 (N_12811,N_7036,N_10363);
or U12812 (N_12812,N_9517,N_6259);
xor U12813 (N_12813,N_11673,N_8225);
xor U12814 (N_12814,N_12230,N_8456);
nand U12815 (N_12815,N_10331,N_6703);
and U12816 (N_12816,N_9262,N_7910);
nand U12817 (N_12817,N_9558,N_7399);
or U12818 (N_12818,N_6533,N_8961);
xnor U12819 (N_12819,N_7960,N_12009);
and U12820 (N_12820,N_10742,N_9653);
nor U12821 (N_12821,N_10228,N_11211);
and U12822 (N_12822,N_10540,N_8434);
nand U12823 (N_12823,N_10319,N_10440);
and U12824 (N_12824,N_6326,N_11797);
nor U12825 (N_12825,N_11909,N_6908);
nand U12826 (N_12826,N_6523,N_11936);
xor U12827 (N_12827,N_9922,N_11607);
nor U12828 (N_12828,N_10539,N_8415);
and U12829 (N_12829,N_6945,N_10398);
nand U12830 (N_12830,N_6529,N_7259);
nor U12831 (N_12831,N_6323,N_7800);
xnor U12832 (N_12832,N_7286,N_6854);
xor U12833 (N_12833,N_8612,N_9348);
nand U12834 (N_12834,N_12289,N_7567);
nor U12835 (N_12835,N_6296,N_10957);
or U12836 (N_12836,N_8117,N_11863);
nand U12837 (N_12837,N_9249,N_9816);
xnor U12838 (N_12838,N_9728,N_8049);
or U12839 (N_12839,N_8957,N_11581);
nand U12840 (N_12840,N_9132,N_10548);
nor U12841 (N_12841,N_10791,N_9692);
and U12842 (N_12842,N_8324,N_10232);
xor U12843 (N_12843,N_7955,N_9608);
nand U12844 (N_12844,N_9335,N_7925);
nand U12845 (N_12845,N_6338,N_9440);
nand U12846 (N_12846,N_8948,N_8040);
or U12847 (N_12847,N_8263,N_7083);
xor U12848 (N_12848,N_10935,N_10333);
xnor U12849 (N_12849,N_7996,N_12435);
or U12850 (N_12850,N_10396,N_7283);
nand U12851 (N_12851,N_9253,N_12456);
xnor U12852 (N_12852,N_9229,N_7013);
xor U12853 (N_12853,N_8561,N_7473);
and U12854 (N_12854,N_9170,N_6884);
nor U12855 (N_12855,N_6309,N_9305);
or U12856 (N_12856,N_8382,N_11389);
xor U12857 (N_12857,N_7099,N_11932);
and U12858 (N_12858,N_11722,N_11407);
or U12859 (N_12859,N_6731,N_6827);
nor U12860 (N_12860,N_8482,N_11668);
nand U12861 (N_12861,N_11376,N_12103);
or U12862 (N_12862,N_8518,N_9553);
nor U12863 (N_12863,N_7632,N_11220);
or U12864 (N_12864,N_11457,N_10592);
nor U12865 (N_12865,N_9040,N_11721);
nand U12866 (N_12866,N_10146,N_6528);
or U12867 (N_12867,N_11309,N_11401);
or U12868 (N_12868,N_7003,N_6801);
nor U12869 (N_12869,N_11116,N_6461);
nor U12870 (N_12870,N_7084,N_8343);
xor U12871 (N_12871,N_11643,N_7300);
nand U12872 (N_12872,N_12256,N_11998);
and U12873 (N_12873,N_8852,N_9204);
nand U12874 (N_12874,N_10536,N_6994);
nor U12875 (N_12875,N_12249,N_9702);
and U12876 (N_12876,N_6710,N_9533);
or U12877 (N_12877,N_10963,N_10131);
nor U12878 (N_12878,N_6511,N_12259);
or U12879 (N_12879,N_11913,N_8810);
or U12880 (N_12880,N_9187,N_8094);
nor U12881 (N_12881,N_8829,N_11714);
xor U12882 (N_12882,N_11498,N_8705);
xnor U12883 (N_12883,N_8508,N_7654);
xor U12884 (N_12884,N_9921,N_10239);
nand U12885 (N_12885,N_9405,N_6524);
or U12886 (N_12886,N_10466,N_12166);
xnor U12887 (N_12887,N_9191,N_7166);
or U12888 (N_12888,N_7346,N_6954);
nand U12889 (N_12889,N_6813,N_9899);
xnor U12890 (N_12890,N_8898,N_7613);
and U12891 (N_12891,N_11850,N_8404);
nor U12892 (N_12892,N_11517,N_6635);
or U12893 (N_12893,N_8306,N_10811);
nand U12894 (N_12894,N_11412,N_12187);
and U12895 (N_12895,N_7097,N_6437);
or U12896 (N_12896,N_7523,N_7169);
xnor U12897 (N_12897,N_8520,N_7526);
nor U12898 (N_12898,N_10940,N_9918);
or U12899 (N_12899,N_6711,N_9898);
nor U12900 (N_12900,N_11486,N_9098);
and U12901 (N_12901,N_9251,N_6307);
nor U12902 (N_12902,N_7588,N_8604);
xor U12903 (N_12903,N_8411,N_10514);
xor U12904 (N_12904,N_7635,N_10102);
and U12905 (N_12905,N_10925,N_11594);
nand U12906 (N_12906,N_6918,N_12384);
xnor U12907 (N_12907,N_12489,N_8934);
nand U12908 (N_12908,N_8619,N_11197);
nor U12909 (N_12909,N_11337,N_10960);
and U12910 (N_12910,N_12079,N_8229);
nor U12911 (N_12911,N_7451,N_9647);
nor U12912 (N_12912,N_9554,N_11791);
and U12913 (N_12913,N_7905,N_11443);
and U12914 (N_12914,N_6345,N_11056);
nor U12915 (N_12915,N_6944,N_9436);
and U12916 (N_12916,N_6961,N_11422);
nand U12917 (N_12917,N_10100,N_12429);
and U12918 (N_12918,N_7038,N_8466);
xnor U12919 (N_12919,N_10664,N_7564);
nand U12920 (N_12920,N_8334,N_8853);
nand U12921 (N_12921,N_6367,N_11865);
or U12922 (N_12922,N_10835,N_10696);
nor U12923 (N_12923,N_8781,N_9273);
nor U12924 (N_12924,N_8202,N_11453);
nand U12925 (N_12925,N_10900,N_7496);
nand U12926 (N_12926,N_7837,N_8768);
nor U12927 (N_12927,N_11849,N_11915);
nor U12928 (N_12928,N_10939,N_10832);
nand U12929 (N_12929,N_12465,N_11416);
or U12930 (N_12930,N_8992,N_10283);
or U12931 (N_12931,N_10854,N_12040);
and U12932 (N_12932,N_7797,N_6428);
nor U12933 (N_12933,N_10437,N_6519);
xor U12934 (N_12934,N_11479,N_8813);
nand U12935 (N_12935,N_11474,N_12236);
and U12936 (N_12936,N_10011,N_9664);
nand U12937 (N_12937,N_7112,N_6423);
nor U12938 (N_12938,N_10495,N_10680);
and U12939 (N_12939,N_6880,N_11398);
nor U12940 (N_12940,N_6468,N_9760);
xor U12941 (N_12941,N_8087,N_6384);
nand U12942 (N_12942,N_6516,N_9893);
xor U12943 (N_12943,N_10789,N_7082);
xnor U12944 (N_12944,N_7598,N_7357);
or U12945 (N_12945,N_8770,N_12216);
nand U12946 (N_12946,N_10167,N_9953);
nor U12947 (N_12947,N_8686,N_11628);
nand U12948 (N_12948,N_10168,N_11795);
xnor U12949 (N_12949,N_6677,N_11777);
or U12950 (N_12950,N_12127,N_9057);
nand U12951 (N_12951,N_12226,N_8999);
and U12952 (N_12952,N_7419,N_9307);
or U12953 (N_12953,N_7116,N_6474);
and U12954 (N_12954,N_6399,N_12455);
nor U12955 (N_12955,N_10550,N_7535);
xnor U12956 (N_12956,N_12403,N_7918);
nor U12957 (N_12957,N_8036,N_8042);
nor U12958 (N_12958,N_10848,N_7786);
nor U12959 (N_12959,N_7050,N_10439);
or U12960 (N_12960,N_8027,N_9367);
nor U12961 (N_12961,N_12017,N_11449);
nand U12962 (N_12962,N_11811,N_8409);
nand U12963 (N_12963,N_6723,N_9003);
nor U12964 (N_12964,N_11745,N_11139);
nor U12965 (N_12965,N_8279,N_11980);
and U12966 (N_12966,N_7542,N_7782);
nor U12967 (N_12967,N_7649,N_7502);
or U12968 (N_12968,N_7409,N_10166);
and U12969 (N_12969,N_7514,N_6721);
and U12970 (N_12970,N_11187,N_11170);
nand U12971 (N_12971,N_7411,N_7761);
or U12972 (N_12972,N_9842,N_6416);
nand U12973 (N_12973,N_10467,N_6740);
nor U12974 (N_12974,N_7848,N_7511);
or U12975 (N_12975,N_9133,N_11971);
and U12976 (N_12976,N_7246,N_6531);
xor U12977 (N_12977,N_10679,N_7377);
or U12978 (N_12978,N_7406,N_11844);
nand U12979 (N_12979,N_7443,N_9562);
or U12980 (N_12980,N_11788,N_11049);
xor U12981 (N_12981,N_8278,N_6636);
and U12982 (N_12982,N_7764,N_12317);
and U12983 (N_12983,N_11560,N_10505);
nand U12984 (N_12984,N_7096,N_11096);
and U12985 (N_12985,N_6403,N_11032);
nor U12986 (N_12986,N_8850,N_6378);
nand U12987 (N_12987,N_12412,N_10633);
or U12988 (N_12988,N_10813,N_8968);
nor U12989 (N_12989,N_10591,N_11236);
or U12990 (N_12990,N_6821,N_9319);
or U12991 (N_12991,N_8088,N_11237);
and U12992 (N_12992,N_7306,N_11642);
and U12993 (N_12993,N_8442,N_9406);
or U12994 (N_12994,N_11185,N_10405);
or U12995 (N_12995,N_10977,N_7922);
xnor U12996 (N_12996,N_7776,N_11941);
and U12997 (N_12997,N_12416,N_10663);
and U12998 (N_12998,N_10272,N_7310);
and U12999 (N_12999,N_6634,N_8910);
and U13000 (N_13000,N_7315,N_8236);
or U13001 (N_13001,N_10037,N_7714);
nand U13002 (N_13002,N_7531,N_10788);
nor U13003 (N_13003,N_11728,N_9527);
xor U13004 (N_13004,N_10586,N_6704);
nand U13005 (N_13005,N_10733,N_8877);
and U13006 (N_13006,N_7652,N_11564);
and U13007 (N_13007,N_9018,N_7791);
and U13008 (N_13008,N_9490,N_11028);
nor U13009 (N_13009,N_10899,N_6805);
nor U13010 (N_13010,N_7446,N_10757);
nand U13011 (N_13011,N_10541,N_12440);
xor U13012 (N_13012,N_11425,N_10739);
nand U13013 (N_13013,N_7736,N_6318);
xnor U13014 (N_13014,N_10735,N_8001);
nand U13015 (N_13015,N_6866,N_11860);
xor U13016 (N_13016,N_10068,N_10703);
and U13017 (N_13017,N_11635,N_6718);
and U13018 (N_13018,N_10284,N_10806);
xnor U13019 (N_13019,N_9536,N_10648);
nand U13020 (N_13020,N_8698,N_8273);
nand U13021 (N_13021,N_9879,N_11841);
or U13022 (N_13022,N_7832,N_10750);
and U13023 (N_13023,N_6899,N_6625);
nor U13024 (N_13024,N_7416,N_9470);
and U13025 (N_13025,N_10207,N_9847);
nand U13026 (N_13026,N_11506,N_11024);
xnor U13027 (N_13027,N_9512,N_12073);
or U13028 (N_13028,N_10658,N_10446);
or U13029 (N_13029,N_9180,N_11205);
nor U13030 (N_13030,N_11332,N_9747);
or U13031 (N_13031,N_7351,N_10580);
and U13032 (N_13032,N_9724,N_7584);
or U13033 (N_13033,N_6436,N_8749);
nand U13034 (N_13034,N_9831,N_7519);
xor U13035 (N_13035,N_10169,N_11285);
xor U13036 (N_13036,N_8976,N_10494);
or U13037 (N_13037,N_10379,N_9658);
and U13038 (N_13038,N_7468,N_6925);
xnor U13039 (N_13039,N_8271,N_9084);
xor U13040 (N_13040,N_10094,N_8621);
xor U13041 (N_13041,N_11618,N_10270);
xnor U13042 (N_13042,N_9573,N_6924);
and U13043 (N_13043,N_8008,N_10574);
or U13044 (N_13044,N_6562,N_7194);
or U13045 (N_13045,N_8805,N_10222);
and U13046 (N_13046,N_9962,N_9372);
nand U13047 (N_13047,N_7285,N_6315);
or U13048 (N_13048,N_9648,N_6404);
or U13049 (N_13049,N_10254,N_12425);
xor U13050 (N_13050,N_9110,N_9854);
or U13051 (N_13051,N_9322,N_10981);
and U13052 (N_13052,N_11894,N_8173);
and U13053 (N_13053,N_7787,N_12374);
nand U13054 (N_13054,N_6586,N_10902);
xor U13055 (N_13055,N_6610,N_9885);
nor U13056 (N_13056,N_11883,N_6481);
or U13057 (N_13057,N_8403,N_12063);
nand U13058 (N_13058,N_6255,N_9173);
and U13059 (N_13059,N_12168,N_9168);
or U13060 (N_13060,N_11390,N_8233);
and U13061 (N_13061,N_10080,N_12120);
or U13062 (N_13062,N_6250,N_11911);
or U13063 (N_13063,N_9101,N_9267);
and U13064 (N_13064,N_12294,N_8818);
nand U13065 (N_13065,N_10295,N_6759);
and U13066 (N_13066,N_7817,N_10709);
nor U13067 (N_13067,N_6753,N_11923);
xnor U13068 (N_13068,N_6942,N_10572);
xnor U13069 (N_13069,N_10579,N_8114);
or U13070 (N_13070,N_6894,N_9666);
nand U13071 (N_13071,N_10252,N_8795);
and U13072 (N_13072,N_11484,N_10851);
and U13073 (N_13073,N_11687,N_9103);
or U13074 (N_13074,N_8352,N_8269);
and U13075 (N_13075,N_6321,N_11624);
nand U13076 (N_13076,N_12269,N_7336);
and U13077 (N_13077,N_10815,N_6689);
nor U13078 (N_13078,N_7726,N_6829);
and U13079 (N_13079,N_11436,N_6706);
nor U13080 (N_13080,N_7035,N_11350);
nand U13081 (N_13081,N_6447,N_11870);
and U13082 (N_13082,N_10138,N_10267);
nand U13083 (N_13083,N_9364,N_6614);
or U13084 (N_13084,N_11854,N_8502);
nand U13085 (N_13085,N_8120,N_9781);
and U13086 (N_13086,N_10223,N_7784);
nand U13087 (N_13087,N_8298,N_11137);
nand U13088 (N_13088,N_8772,N_7034);
xor U13089 (N_13089,N_11117,N_11046);
or U13090 (N_13090,N_8868,N_10560);
nand U13091 (N_13091,N_10212,N_6717);
and U13092 (N_13092,N_11991,N_8210);
nor U13093 (N_13093,N_8142,N_9772);
or U13094 (N_13094,N_8523,N_12360);
nor U13095 (N_13095,N_9292,N_8613);
nand U13096 (N_13096,N_12076,N_9286);
nand U13097 (N_13097,N_9740,N_9929);
or U13098 (N_13098,N_8270,N_7118);
nor U13099 (N_13099,N_10681,N_11562);
nand U13100 (N_13100,N_9113,N_12095);
xnor U13101 (N_13101,N_12104,N_9143);
nand U13102 (N_13102,N_7546,N_10529);
and U13103 (N_13103,N_8140,N_8363);
or U13104 (N_13104,N_6464,N_7264);
or U13105 (N_13105,N_8990,N_10111);
nor U13106 (N_13106,N_11202,N_7595);
or U13107 (N_13107,N_8494,N_8031);
and U13108 (N_13108,N_11308,N_7305);
or U13109 (N_13109,N_10783,N_10107);
xor U13110 (N_13110,N_11041,N_9127);
xor U13111 (N_13111,N_8433,N_6320);
xnor U13112 (N_13112,N_8908,N_6836);
and U13113 (N_13113,N_7002,N_9236);
nand U13114 (N_13114,N_9467,N_11759);
nand U13115 (N_13115,N_10173,N_7636);
or U13116 (N_13116,N_8241,N_8101);
xnor U13117 (N_13117,N_8395,N_9272);
and U13118 (N_13118,N_8362,N_8424);
nand U13119 (N_13119,N_11015,N_9835);
nand U13120 (N_13120,N_10804,N_6765);
and U13121 (N_13121,N_12044,N_9810);
and U13122 (N_13122,N_8285,N_11244);
nand U13123 (N_13123,N_9756,N_7225);
nand U13124 (N_13124,N_10535,N_12032);
nand U13125 (N_13125,N_10214,N_9901);
nand U13126 (N_13126,N_6268,N_10975);
and U13127 (N_13127,N_12003,N_10279);
xor U13128 (N_13128,N_9537,N_11408);
or U13129 (N_13129,N_7500,N_10348);
and U13130 (N_13130,N_7260,N_8350);
and U13131 (N_13131,N_11489,N_11592);
and U13132 (N_13132,N_8678,N_10046);
nor U13133 (N_13133,N_10299,N_6847);
or U13134 (N_13134,N_9317,N_10305);
nor U13135 (N_13135,N_10391,N_8673);
xor U13136 (N_13136,N_11394,N_6490);
nand U13137 (N_13137,N_8512,N_8441);
and U13138 (N_13138,N_10534,N_11199);
or U13139 (N_13139,N_10906,N_10042);
or U13140 (N_13140,N_8758,N_9341);
nor U13141 (N_13141,N_8970,N_6719);
or U13142 (N_13142,N_12483,N_12128);
and U13143 (N_13143,N_6432,N_11419);
nand U13144 (N_13144,N_11763,N_9160);
nor U13145 (N_13145,N_12303,N_9649);
nand U13146 (N_13146,N_7430,N_7298);
nor U13147 (N_13147,N_7041,N_8568);
nor U13148 (N_13148,N_8253,N_9679);
and U13149 (N_13149,N_8525,N_10844);
nor U13150 (N_13150,N_11817,N_7189);
xor U13151 (N_13151,N_10870,N_12077);
nor U13152 (N_13152,N_10288,N_9550);
nand U13153 (N_13153,N_6665,N_6487);
nand U13154 (N_13154,N_10304,N_9002);
and U13155 (N_13155,N_7504,N_9498);
and U13156 (N_13156,N_7394,N_11965);
or U13157 (N_13157,N_11597,N_8557);
nor U13158 (N_13158,N_12163,N_12285);
nand U13159 (N_13159,N_12049,N_9242);
nand U13160 (N_13160,N_10251,N_10413);
nor U13161 (N_13161,N_9940,N_10866);
or U13162 (N_13162,N_8355,N_9076);
and U13163 (N_13163,N_6691,N_11341);
nor U13164 (N_13164,N_12457,N_8012);
or U13165 (N_13165,N_9136,N_10113);
nor U13166 (N_13166,N_7266,N_7176);
nor U13167 (N_13167,N_6708,N_12293);
and U13168 (N_13168,N_9401,N_6807);
xnor U13169 (N_13169,N_10853,N_6643);
or U13170 (N_13170,N_9296,N_9736);
nand U13171 (N_13171,N_10082,N_8593);
nand U13172 (N_13172,N_10154,N_7232);
and U13173 (N_13173,N_7753,N_7968);
or U13174 (N_13174,N_12054,N_12453);
nor U13175 (N_13175,N_12471,N_7804);
xor U13176 (N_13176,N_9525,N_8435);
and U13177 (N_13177,N_10263,N_12101);
nand U13178 (N_13178,N_7591,N_6582);
nand U13179 (N_13179,N_11230,N_9145);
and U13180 (N_13180,N_12454,N_11099);
or U13181 (N_13181,N_10375,N_6264);
nand U13182 (N_13182,N_9635,N_7321);
and U13183 (N_13183,N_11842,N_12183);
or U13184 (N_13184,N_10847,N_6430);
nor U13185 (N_13185,N_6330,N_8326);
nand U13186 (N_13186,N_6272,N_12296);
nand U13187 (N_13187,N_9355,N_12389);
or U13188 (N_13188,N_7947,N_11903);
or U13189 (N_13189,N_8305,N_8663);
nor U13190 (N_13190,N_9245,N_7325);
xnor U13191 (N_13191,N_9395,N_8634);
or U13192 (N_13192,N_10816,N_11775);
or U13193 (N_13193,N_10163,N_11442);
nand U13194 (N_13194,N_6444,N_8422);
and U13195 (N_13195,N_7494,N_8799);
nand U13196 (N_13196,N_11279,N_12346);
nand U13197 (N_13197,N_8697,N_11179);
or U13198 (N_13198,N_12167,N_7562);
and U13199 (N_13199,N_8337,N_7465);
or U13200 (N_13200,N_11831,N_7731);
or U13201 (N_13201,N_6422,N_10078);
nand U13202 (N_13202,N_11300,N_10985);
or U13203 (N_13203,N_8755,N_9802);
nand U13204 (N_13204,N_11379,N_7061);
and U13205 (N_13205,N_12081,N_6955);
or U13206 (N_13206,N_12152,N_8247);
and U13207 (N_13207,N_7480,N_12014);
nand U13208 (N_13208,N_6845,N_7509);
xor U13209 (N_13209,N_10294,N_12460);
xnor U13210 (N_13210,N_7902,N_10216);
xnor U13211 (N_13211,N_12379,N_9435);
or U13212 (N_13212,N_7557,N_8776);
and U13213 (N_13213,N_7824,N_12090);
or U13214 (N_13214,N_6927,N_6853);
nand U13215 (N_13215,N_6887,N_8900);
and U13216 (N_13216,N_10544,N_8133);
xor U13217 (N_13217,N_8851,N_9661);
or U13218 (N_13218,N_6781,N_8547);
nand U13219 (N_13219,N_9758,N_11686);
nor U13220 (N_13220,N_7068,N_7295);
nand U13221 (N_13221,N_9172,N_10238);
or U13222 (N_13222,N_11879,N_11992);
and U13223 (N_13223,N_8671,N_8715);
xor U13224 (N_13224,N_9300,N_10649);
nor U13225 (N_13225,N_9569,N_11215);
and U13226 (N_13226,N_7078,N_9606);
and U13227 (N_13227,N_8630,N_10697);
and U13228 (N_13228,N_8832,N_9441);
xor U13229 (N_13229,N_11273,N_7213);
nor U13230 (N_13230,N_7743,N_6828);
and U13231 (N_13231,N_6831,N_6375);
nand U13232 (N_13232,N_9988,N_10448);
nand U13233 (N_13233,N_10843,N_8039);
xor U13234 (N_13234,N_8108,N_10988);
nand U13235 (N_13235,N_9836,N_8457);
nand U13236 (N_13236,N_10186,N_9294);
nor U13237 (N_13237,N_8336,N_9159);
nand U13238 (N_13238,N_8376,N_12208);
nand U13239 (N_13239,N_6515,N_6970);
and U13240 (N_13240,N_6425,N_7961);
or U13241 (N_13241,N_8346,N_7616);
nand U13242 (N_13242,N_6583,N_11080);
or U13243 (N_13243,N_12117,N_8387);
nand U13244 (N_13244,N_11483,N_7228);
or U13245 (N_13245,N_7997,N_11463);
or U13246 (N_13246,N_10502,N_8556);
or U13247 (N_13247,N_9599,N_8183);
nor U13248 (N_13248,N_11124,N_7882);
xnor U13249 (N_13249,N_11698,N_6638);
nor U13250 (N_13250,N_10062,N_9678);
xnor U13251 (N_13251,N_6911,N_7327);
nor U13252 (N_13252,N_6626,N_8566);
and U13253 (N_13253,N_6975,N_9351);
and U13254 (N_13254,N_9643,N_12123);
nand U13255 (N_13255,N_11472,N_8191);
or U13256 (N_13256,N_8288,N_9629);
nor U13257 (N_13257,N_10029,N_12059);
xnor U13258 (N_13258,N_11780,N_10488);
or U13259 (N_13259,N_11467,N_8886);
nor U13260 (N_13260,N_11530,N_8085);
nor U13261 (N_13261,N_10015,N_10229);
nor U13262 (N_13262,N_9179,N_10636);
xor U13263 (N_13263,N_11606,N_10577);
xor U13264 (N_13264,N_7212,N_8757);
or U13265 (N_13265,N_9112,N_10352);
nand U13266 (N_13266,N_12332,N_7610);
nor U13267 (N_13267,N_7951,N_11935);
nand U13268 (N_13268,N_10715,N_7284);
nor U13269 (N_13269,N_9496,N_12260);
and U13270 (N_13270,N_12434,N_9088);
xor U13271 (N_13271,N_11641,N_7989);
or U13272 (N_13272,N_6291,N_8171);
or U13273 (N_13273,N_8860,N_11106);
xor U13274 (N_13274,N_12381,N_10043);
nand U13275 (N_13275,N_11164,N_9754);
nand U13276 (N_13276,N_12404,N_11789);
nor U13277 (N_13277,N_8370,N_12341);
and U13278 (N_13278,N_10438,N_8014);
and U13279 (N_13279,N_8926,N_8380);
nand U13280 (N_13280,N_7328,N_11458);
nor U13281 (N_13281,N_8659,N_7571);
xor U13282 (N_13282,N_8491,N_10060);
xnor U13283 (N_13283,N_8158,N_9588);
xor U13284 (N_13284,N_8111,N_8399);
and U13285 (N_13285,N_6984,N_8756);
or U13286 (N_13286,N_9047,N_7907);
nor U13287 (N_13287,N_8449,N_8816);
xnor U13288 (N_13288,N_11328,N_9896);
and U13289 (N_13289,N_11853,N_7501);
and U13290 (N_13290,N_8402,N_8250);
nand U13291 (N_13291,N_8587,N_7437);
nand U13292 (N_13292,N_11302,N_6578);
or U13293 (N_13293,N_8116,N_11958);
and U13294 (N_13294,N_11083,N_11568);
nor U13295 (N_13295,N_11577,N_11331);
xnor U13296 (N_13296,N_10334,N_9020);
or U13297 (N_13297,N_8899,N_12156);
or U13298 (N_13298,N_8022,N_12413);
or U13299 (N_13299,N_9000,N_9090);
and U13300 (N_13300,N_9094,N_9135);
xnor U13301 (N_13301,N_6743,N_6263);
nand U13302 (N_13302,N_8513,N_11246);
nor U13303 (N_13303,N_8553,N_11283);
xor U13304 (N_13304,N_7128,N_12111);
xor U13305 (N_13305,N_10898,N_7637);
nor U13306 (N_13306,N_6566,N_9791);
nand U13307 (N_13307,N_9863,N_10954);
nor U13308 (N_13308,N_9950,N_11322);
nor U13309 (N_13309,N_9226,N_11723);
and U13310 (N_13310,N_11973,N_8975);
and U13311 (N_13311,N_6355,N_11809);
or U13312 (N_13312,N_7853,N_7371);
nor U13313 (N_13313,N_9811,N_9691);
nor U13314 (N_13314,N_11536,N_11585);
and U13315 (N_13315,N_8668,N_9592);
nand U13316 (N_13316,N_11533,N_10708);
xor U13317 (N_13317,N_10503,N_9834);
xor U13318 (N_13318,N_8463,N_11326);
or U13319 (N_13319,N_10026,N_7617);
or U13320 (N_13320,N_9564,N_6985);
and U13321 (N_13321,N_11510,N_10240);
xor U13322 (N_13322,N_7839,N_10419);
and U13323 (N_13323,N_9174,N_11946);
nand U13324 (N_13324,N_8717,N_6669);
or U13325 (N_13325,N_11630,N_9539);
nand U13326 (N_13326,N_9713,N_9268);
and U13327 (N_13327,N_7344,N_8930);
nor U13328 (N_13328,N_6921,N_7448);
or U13329 (N_13329,N_11707,N_12112);
nor U13330 (N_13330,N_7819,N_10172);
nand U13331 (N_13331,N_7831,N_7248);
xor U13332 (N_13332,N_11959,N_7464);
xnor U13333 (N_13333,N_10943,N_12492);
nand U13334 (N_13334,N_11892,N_8199);
nor U13335 (N_13335,N_8068,N_9042);
and U13336 (N_13336,N_6658,N_8707);
nor U13337 (N_13337,N_9710,N_9693);
nor U13338 (N_13338,N_8169,N_6798);
nand U13339 (N_13339,N_12451,N_8884);
xor U13340 (N_13340,N_12185,N_11679);
and U13341 (N_13341,N_11025,N_9803);
and U13342 (N_13342,N_8340,N_7746);
xor U13343 (N_13343,N_11864,N_6328);
nor U13344 (N_13344,N_9722,N_10508);
nand U13345 (N_13345,N_6640,N_9134);
nand U13346 (N_13346,N_6875,N_11207);
xor U13347 (N_13347,N_11636,N_10350);
xnor U13348 (N_13348,N_9244,N_6990);
or U13349 (N_13349,N_6878,N_12004);
nand U13350 (N_13350,N_9799,N_9396);
xor U13351 (N_13351,N_9447,N_10069);
nand U13352 (N_13352,N_12306,N_10462);
xor U13353 (N_13353,N_9444,N_10456);
or U13354 (N_13354,N_10587,N_6534);
nand U13355 (N_13355,N_9499,N_12390);
nand U13356 (N_13356,N_8728,N_11431);
and U13357 (N_13357,N_8912,N_8070);
or U13358 (N_13358,N_8915,N_6917);
and U13359 (N_13359,N_9451,N_8495);
and U13360 (N_13360,N_10982,N_8481);
and U13361 (N_13361,N_10442,N_6581);
and U13362 (N_13362,N_9585,N_9469);
or U13363 (N_13363,N_10004,N_9587);
nor U13364 (N_13364,N_10968,N_10769);
nand U13365 (N_13365,N_8703,N_9977);
and U13366 (N_13366,N_10394,N_9349);
nor U13367 (N_13367,N_6976,N_9686);
nor U13368 (N_13368,N_8486,N_11990);
nor U13369 (N_13369,N_7805,N_12333);
or U13370 (N_13370,N_7568,N_9163);
xor U13371 (N_13371,N_7127,N_10054);
and U13372 (N_13372,N_7222,N_11306);
nor U13373 (N_13373,N_9100,N_7163);
nor U13374 (N_13374,N_9387,N_10717);
xor U13375 (N_13375,N_11511,N_10915);
xor U13376 (N_13376,N_6431,N_8385);
or U13377 (N_13377,N_12309,N_8197);
or U13378 (N_13378,N_10280,N_7868);
or U13379 (N_13379,N_8331,N_6972);
nand U13380 (N_13380,N_8147,N_8809);
nor U13381 (N_13381,N_9033,N_8918);
and U13382 (N_13382,N_9460,N_7151);
xnor U13383 (N_13383,N_7603,N_9589);
nor U13384 (N_13384,N_9873,N_8662);
xor U13385 (N_13385,N_11985,N_9801);
nor U13386 (N_13386,N_7765,N_10753);
or U13387 (N_13387,N_11807,N_10860);
nor U13388 (N_13388,N_6683,N_8687);
nand U13389 (N_13389,N_6698,N_11321);
nor U13390 (N_13390,N_8965,N_11045);
nor U13391 (N_13391,N_10067,N_9544);
and U13392 (N_13392,N_9928,N_12053);
xnor U13393 (N_13393,N_10155,N_10455);
or U13394 (N_13394,N_10855,N_9969);
and U13395 (N_13395,N_11098,N_9755);
xnor U13396 (N_13396,N_10325,N_7425);
nor U13397 (N_13397,N_6526,N_12042);
or U13398 (N_13398,N_6438,N_7489);
nor U13399 (N_13399,N_9454,N_11760);
xor U13400 (N_13400,N_7934,N_10185);
nand U13401 (N_13401,N_12331,N_8396);
nand U13402 (N_13402,N_9514,N_11171);
or U13403 (N_13403,N_8938,N_11534);
nor U13404 (N_13404,N_8161,N_10776);
xnor U13405 (N_13405,N_11820,N_6811);
nand U13406 (N_13406,N_11779,N_7900);
and U13407 (N_13407,N_9495,N_6810);
or U13408 (N_13408,N_12444,N_7141);
nand U13409 (N_13409,N_12164,N_12322);
or U13410 (N_13410,N_9326,N_10425);
or U13411 (N_13411,N_10642,N_10598);
nand U13412 (N_13412,N_10097,N_10976);
and U13413 (N_13413,N_9767,N_11839);
or U13414 (N_13414,N_12347,N_6661);
and U13415 (N_13415,N_10754,N_9733);
nor U13416 (N_13416,N_6979,N_10865);
xnor U13417 (N_13417,N_7650,N_6537);
xor U13418 (N_13418,N_7757,N_8182);
nand U13419 (N_13419,N_12231,N_9449);
xor U13420 (N_13420,N_10364,N_9545);
xnor U13421 (N_13421,N_11180,N_12369);
nand U13422 (N_13422,N_9186,N_7706);
nand U13423 (N_13423,N_11238,N_9257);
or U13424 (N_13424,N_10368,N_7117);
or U13425 (N_13425,N_9843,N_8347);
or U13426 (N_13426,N_9994,N_8838);
and U13427 (N_13427,N_10886,N_9023);
nand U13428 (N_13428,N_11986,N_8559);
xor U13429 (N_13429,N_7707,N_9930);
nor U13430 (N_13430,N_8023,N_9878);
nand U13431 (N_13431,N_11370,N_7161);
nor U13432 (N_13432,N_11160,N_9626);
xnor U13433 (N_13433,N_10738,N_8200);
xor U13434 (N_13434,N_10259,N_12473);
or U13435 (N_13435,N_8460,N_9768);
xor U13436 (N_13436,N_7179,N_8939);
and U13437 (N_13437,N_10570,N_10718);
nor U13438 (N_13438,N_7609,N_6650);
or U13439 (N_13439,N_8599,N_8614);
and U13440 (N_13440,N_12356,N_12438);
nand U13441 (N_13441,N_8323,N_8203);
nor U13442 (N_13442,N_9433,N_10953);
xnor U13443 (N_13443,N_6484,N_9121);
xor U13444 (N_13444,N_11445,N_11294);
xor U13445 (N_13445,N_12047,N_11356);
or U13446 (N_13446,N_7499,N_12439);
nor U13447 (N_13447,N_11107,N_7404);
and U13448 (N_13448,N_11708,N_7885);
and U13449 (N_13449,N_7766,N_9815);
and U13450 (N_13450,N_11586,N_12218);
and U13451 (N_13451,N_8294,N_9082);
nand U13452 (N_13452,N_10492,N_6782);
or U13453 (N_13453,N_11426,N_10204);
and U13454 (N_13454,N_11794,N_9483);
or U13455 (N_13455,N_6408,N_8212);
xor U13456 (N_13456,N_8426,N_11799);
and U13457 (N_13457,N_7926,N_9178);
nor U13458 (N_13458,N_7029,N_11002);
nor U13459 (N_13459,N_12055,N_8714);
nand U13460 (N_13460,N_8532,N_11104);
and U13461 (N_13461,N_8623,N_9874);
or U13462 (N_13462,N_6560,N_7808);
or U13463 (N_13463,N_11427,N_11035);
xnor U13464 (N_13464,N_7196,N_9397);
nor U13465 (N_13465,N_10867,N_7388);
nor U13466 (N_13466,N_11512,N_11138);
xor U13467 (N_13467,N_8104,N_10158);
nor U13468 (N_13468,N_12154,N_9954);
nand U13469 (N_13469,N_9567,N_11344);
and U13470 (N_13470,N_6390,N_8048);
xnor U13471 (N_13471,N_8281,N_12376);
or U13472 (N_13472,N_10989,N_6857);
nand U13473 (N_13473,N_11268,N_11047);
nand U13474 (N_13474,N_7313,N_12329);
nand U13475 (N_13475,N_7268,N_12250);
or U13476 (N_13476,N_8498,N_9492);
xor U13477 (N_13477,N_9526,N_7387);
and U13478 (N_13478,N_12026,N_10351);
and U13479 (N_13479,N_10803,N_8172);
nor U13480 (N_13480,N_9083,N_11884);
or U13481 (N_13481,N_9363,N_7943);
or U13482 (N_13482,N_8238,N_9777);
and U13483 (N_13483,N_12291,N_7136);
nand U13484 (N_13484,N_11888,N_9386);
xnor U13485 (N_13485,N_7565,N_7979);
nor U13486 (N_13486,N_12036,N_8825);
nand U13487 (N_13487,N_7491,N_8846);
nor U13488 (N_13488,N_12274,N_12342);
xor U13489 (N_13489,N_9738,N_6544);
or U13490 (N_13490,N_6442,N_6879);
nor U13491 (N_13491,N_7211,N_7813);
nand U13492 (N_13492,N_11525,N_7091);
nand U13493 (N_13493,N_11816,N_9299);
nand U13494 (N_13494,N_7507,N_7576);
xor U13495 (N_13495,N_9717,N_11267);
xor U13496 (N_13496,N_8730,N_8458);
nand U13497 (N_13497,N_11756,N_8282);
or U13498 (N_13498,N_12248,N_11725);
and U13499 (N_13499,N_9824,N_10837);
nor U13500 (N_13500,N_11705,N_8296);
and U13501 (N_13501,N_10758,N_7276);
and U13502 (N_13502,N_10637,N_8764);
xnor U13503 (N_13503,N_10335,N_9936);
and U13504 (N_13504,N_10210,N_11386);
nand U13505 (N_13505,N_6652,N_11678);
and U13506 (N_13506,N_9337,N_7891);
or U13507 (N_13507,N_11967,N_7842);
nand U13508 (N_13508,N_10710,N_8822);
nor U13509 (N_13509,N_9818,N_10707);
nand U13510 (N_13510,N_7748,N_6760);
xnor U13511 (N_13511,N_11228,N_12270);
nand U13512 (N_13512,N_12493,N_8742);
or U13513 (N_13513,N_7671,N_12268);
or U13514 (N_13514,N_11726,N_9782);
xnor U13515 (N_13515,N_10523,N_7978);
and U13516 (N_13516,N_10445,N_10785);
nor U13517 (N_13517,N_11243,N_11837);
xnor U13518 (N_13518,N_7090,N_10825);
nand U13519 (N_13519,N_7153,N_6888);
nor U13520 (N_13520,N_11266,N_9522);
and U13521 (N_13521,N_6251,N_11460);
nor U13522 (N_13522,N_11502,N_6947);
and U13523 (N_13523,N_6999,N_11270);
nor U13524 (N_13524,N_11685,N_11454);
xnor U13525 (N_13525,N_10017,N_11209);
or U13526 (N_13526,N_6960,N_9670);
and U13527 (N_13527,N_8332,N_6992);
and U13528 (N_13528,N_10725,N_10607);
xor U13529 (N_13529,N_11774,N_9611);
nand U13530 (N_13530,N_7242,N_8501);
and U13531 (N_13531,N_10199,N_9012);
nor U13532 (N_13532,N_9745,N_9639);
and U13533 (N_13533,N_6774,N_7856);
or U13534 (N_13534,N_10385,N_10859);
nor U13535 (N_13535,N_8956,N_7263);
xnor U13536 (N_13536,N_11196,N_10627);
nor U13537 (N_13537,N_10959,N_10414);
nor U13538 (N_13538,N_11764,N_10845);
xor U13539 (N_13539,N_10878,N_9415);
nor U13540 (N_13540,N_8078,N_9688);
xor U13541 (N_13541,N_8299,N_10362);
or U13542 (N_13542,N_9871,N_10175);
nor U13543 (N_13543,N_8615,N_9164);
and U13544 (N_13544,N_9323,N_7293);
nor U13545 (N_13545,N_10430,N_6873);
or U13546 (N_13546,N_11166,N_6780);
or U13547 (N_13547,N_10103,N_7673);
nor U13548 (N_13548,N_7380,N_6906);
nand U13549 (N_13549,N_7383,N_10671);
xnor U13550 (N_13550,N_11487,N_7730);
and U13551 (N_13551,N_9894,N_12307);
and U13552 (N_13552,N_6588,N_7521);
nand U13553 (N_13553,N_11257,N_6406);
nor U13554 (N_13554,N_11933,N_10307);
or U13555 (N_13555,N_11916,N_11579);
nor U13556 (N_13556,N_11833,N_6869);
or U13557 (N_13557,N_7005,N_7329);
xnor U13558 (N_13558,N_6746,N_6656);
xnor U13559 (N_13559,N_10743,N_8807);
nor U13560 (N_13560,N_10264,N_7412);
nand U13561 (N_13561,N_12068,N_10630);
xor U13562 (N_13562,N_8865,N_8937);
or U13563 (N_13563,N_11900,N_10208);
xor U13564 (N_13564,N_8374,N_8545);
nand U13565 (N_13565,N_10684,N_10213);
xor U13566 (N_13566,N_12352,N_9718);
nand U13567 (N_13567,N_11832,N_11928);
or U13568 (N_13568,N_8034,N_11055);
nor U13569 (N_13569,N_9439,N_8903);
nor U13570 (N_13570,N_9814,N_12436);
nor U13571 (N_13571,N_8389,N_11671);
or U13572 (N_13572,N_6421,N_7362);
xnor U13573 (N_13573,N_10547,N_9053);
nand U13574 (N_13574,N_6364,N_7644);
and U13575 (N_13575,N_8641,N_12206);
or U13576 (N_13576,N_7758,N_9150);
and U13577 (N_13577,N_10625,N_6400);
nand U13578 (N_13578,N_8811,N_8661);
or U13579 (N_13579,N_11392,N_7527);
nor U13580 (N_13580,N_10507,N_7623);
nand U13581 (N_13581,N_8283,N_8090);
or U13582 (N_13582,N_9749,N_6987);
or U13583 (N_13583,N_9654,N_6377);
or U13584 (N_13584,N_9614,N_8390);
and U13585 (N_13585,N_8469,N_8365);
or U13586 (N_13586,N_8499,N_10120);
or U13587 (N_13587,N_9360,N_7967);
and U13588 (N_13588,N_11578,N_6555);
or U13589 (N_13589,N_12396,N_8864);
or U13590 (N_13590,N_7287,N_9247);
or U13591 (N_13591,N_6988,N_10933);
nand U13592 (N_13592,N_8125,N_11657);
nor U13593 (N_13593,N_6664,N_6592);
nand U13594 (N_13594,N_7838,N_10905);
or U13595 (N_13595,N_7622,N_8633);
nand U13596 (N_13596,N_9716,N_7532);
or U13597 (N_13597,N_10569,N_9434);
and U13598 (N_13598,N_7742,N_7093);
or U13599 (N_13599,N_6356,N_7320);
and U13600 (N_13600,N_10110,N_9610);
and U13601 (N_13601,N_9518,N_7689);
xor U13602 (N_13602,N_7944,N_12116);
nor U13603 (N_13603,N_9906,N_10181);
and U13604 (N_13604,N_8738,N_6546);
nor U13605 (N_13605,N_8300,N_7007);
xor U13606 (N_13606,N_11010,N_11646);
or U13607 (N_13607,N_6799,N_11014);
nor U13608 (N_13608,N_11315,N_11710);
nand U13609 (N_13609,N_9308,N_9581);
and U13610 (N_13610,N_12171,N_10310);
nor U13611 (N_13611,N_9775,N_6937);
nand U13612 (N_13612,N_9709,N_6337);
or U13613 (N_13613,N_11103,N_10309);
xor U13614 (N_13614,N_9230,N_7129);
nor U13615 (N_13615,N_8063,N_12035);
and U13616 (N_13616,N_12295,N_8262);
and U13617 (N_13617,N_9488,N_11917);
nor U13618 (N_13618,N_6678,N_11555);
nand U13619 (N_13619,N_10559,N_9524);
nor U13620 (N_13620,N_7754,N_11323);
or U13621 (N_13621,N_8762,N_7690);
xnor U13622 (N_13622,N_6293,N_11719);
or U13623 (N_13623,N_9215,N_7370);
or U13624 (N_13624,N_8468,N_10444);
nand U13625 (N_13625,N_10489,N_7431);
and U13626 (N_13626,N_10179,N_11348);
nor U13627 (N_13627,N_11478,N_9416);
or U13628 (N_13628,N_12235,N_12319);
nor U13629 (N_13629,N_8013,N_9288);
nor U13630 (N_13630,N_11276,N_10748);
nand U13631 (N_13631,N_7132,N_10292);
nand U13632 (N_13632,N_7043,N_12025);
and U13633 (N_13633,N_12046,N_9939);
nor U13634 (N_13634,N_12283,N_7172);
nor U13635 (N_13635,N_11684,N_10148);
nor U13636 (N_13636,N_11388,N_12367);
nand U13637 (N_13637,N_11119,N_6497);
nand U13638 (N_13638,N_12203,N_9325);
nor U13639 (N_13639,N_11670,N_7233);
and U13640 (N_13640,N_9092,N_10050);
nor U13641 (N_13641,N_6686,N_9231);
or U13642 (N_13642,N_9309,N_10719);
xor U13643 (N_13643,N_9523,N_12267);
xnor U13644 (N_13644,N_11031,N_8497);
xor U13645 (N_13645,N_11699,N_7159);
nand U13646 (N_13646,N_12276,N_9392);
and U13647 (N_13647,N_12124,N_12470);
nand U13648 (N_13648,N_6369,N_7760);
nor U13649 (N_13649,N_7389,N_9278);
nand U13650 (N_13650,N_8949,N_11029);
nor U13651 (N_13651,N_7674,N_7317);
nor U13652 (N_13652,N_8897,N_12143);
or U13653 (N_13653,N_6257,N_9511);
xnor U13654 (N_13654,N_8206,N_6910);
nor U13655 (N_13655,N_12495,N_10247);
nand U13656 (N_13656,N_8153,N_9125);
nand U13657 (N_13657,N_10429,N_7135);
and U13658 (N_13658,N_8339,N_11402);
nor U13659 (N_13659,N_10124,N_10682);
and U13660 (N_13660,N_10133,N_7023);
and U13661 (N_13661,N_7612,N_11920);
and U13662 (N_13662,N_11938,N_7288);
xnor U13663 (N_13663,N_7485,N_9477);
nor U13664 (N_13664,N_8102,N_8690);
nand U13665 (N_13665,N_8265,N_7720);
nor U13666 (N_13666,N_7162,N_12351);
and U13667 (N_13667,N_10293,N_9907);
and U13668 (N_13668,N_9161,N_10830);
or U13669 (N_13669,N_10098,N_8320);
nand U13670 (N_13670,N_10555,N_6417);
and U13671 (N_13671,N_11466,N_11134);
or U13672 (N_13672,N_11057,N_9486);
or U13673 (N_13673,N_9828,N_7744);
and U13674 (N_13674,N_12337,N_7170);
nor U13675 (N_13675,N_9987,N_9301);
nand U13676 (N_13676,N_8138,N_7379);
or U13677 (N_13677,N_7279,N_7641);
xor U13678 (N_13678,N_9452,N_9671);
and U13679 (N_13679,N_9823,N_8984);
or U13680 (N_13680,N_8920,N_8177);
nor U13681 (N_13681,N_9665,N_12499);
or U13682 (N_13682,N_7980,N_10584);
nor U13683 (N_13683,N_7678,N_8689);
nor U13684 (N_13684,N_9726,N_11133);
xor U13685 (N_13685,N_8582,N_11288);
or U13686 (N_13686,N_11038,N_6559);
nand U13687 (N_13687,N_9642,N_7481);
xnor U13688 (N_13688,N_11873,N_9382);
nor U13689 (N_13689,N_8349,N_10383);
xnor U13690 (N_13690,N_8530,N_11834);
xor U13691 (N_13691,N_10883,N_9482);
nand U13692 (N_13692,N_10647,N_7883);
and U13693 (N_13693,N_6603,N_8196);
and U13694 (N_13694,N_7349,N_9660);
nand U13695 (N_13695,N_7420,N_11514);
nor U13696 (N_13696,N_9050,N_11735);
nand U13697 (N_13697,N_11229,N_10415);
nor U13698 (N_13698,N_8033,N_9287);
xnor U13699 (N_13699,N_7415,N_10487);
nor U13700 (N_13700,N_10285,N_9903);
or U13701 (N_13701,N_8314,N_10913);
nand U13702 (N_13702,N_6287,N_11184);
and U13703 (N_13703,N_8546,N_11301);
and U13704 (N_13704,N_11169,N_10727);
xnor U13705 (N_13705,N_9563,N_11631);
nand U13706 (N_13706,N_10688,N_11893);
nor U13707 (N_13707,N_9022,N_6506);
and U13708 (N_13708,N_9773,N_9859);
or U13709 (N_13709,N_8889,N_12400);
nand U13710 (N_13710,N_6991,N_6958);
nor U13711 (N_13711,N_8748,N_8328);
nand U13712 (N_13712,N_11951,N_8222);
xor U13713 (N_13713,N_7407,N_10493);
or U13714 (N_13714,N_10170,N_11153);
or U13715 (N_13715,N_10140,N_6619);
xnor U13716 (N_13716,N_6773,N_12033);
xor U13717 (N_13717,N_11469,N_7439);
xor U13718 (N_13718,N_10770,N_8503);
and U13719 (N_13719,N_12417,N_8882);
nor U13720 (N_13720,N_7917,N_6312);
and U13721 (N_13721,N_7018,N_10109);
and U13722 (N_13722,N_11542,N_7543);
or U13723 (N_13723,N_11480,N_9313);
nor U13724 (N_13724,N_7825,N_9420);
nand U13725 (N_13725,N_10714,N_8905);
nor U13726 (N_13726,N_6727,N_11089);
and U13727 (N_13727,N_6483,N_10435);
and U13728 (N_13728,N_11007,N_10428);
nand U13729 (N_13729,N_8603,N_6964);
or U13730 (N_13730,N_11507,N_11446);
nand U13731 (N_13731,N_8564,N_6274);
xnor U13732 (N_13732,N_9822,N_12129);
xnor U13733 (N_13733,N_7708,N_12109);
and U13734 (N_13734,N_8232,N_11934);
and U13735 (N_13735,N_9986,N_6305);
xor U13736 (N_13736,N_8366,N_7301);
and U13737 (N_13737,N_6269,N_6935);
nor U13738 (N_13738,N_9379,N_9316);
nand U13739 (N_13739,N_9655,N_7087);
nor U13740 (N_13740,N_11523,N_10731);
nand U13741 (N_13741,N_7006,N_9275);
nor U13742 (N_13742,N_10187,N_10178);
and U13743 (N_13743,N_8921,N_9503);
or U13744 (N_13744,N_8239,N_10558);
nor U13745 (N_13745,N_7795,N_10274);
and U13746 (N_13746,N_6288,N_6648);
nand U13747 (N_13747,N_6357,N_11265);
nor U13748 (N_13748,N_6951,N_11914);
and U13749 (N_13749,N_9158,N_7679);
or U13750 (N_13750,N_10491,N_9073);
nor U13751 (N_13751,N_9697,N_11750);
xor U13752 (N_13752,N_9065,N_12237);
or U13753 (N_13753,N_6602,N_10686);
nor U13754 (N_13754,N_8325,N_7756);
nor U13755 (N_13755,N_9844,N_11071);
and U13756 (N_13756,N_11769,N_8052);
and U13757 (N_13757,N_7814,N_11218);
xor U13758 (N_13758,N_7653,N_10893);
or U13759 (N_13759,N_11194,N_7667);
or U13760 (N_13760,N_7292,N_8165);
xnor U13761 (N_13761,N_9389,N_10022);
xnor U13762 (N_13762,N_7347,N_12084);
or U13763 (N_13763,N_7695,N_10842);
xor U13764 (N_13764,N_8490,N_9192);
nand U13765 (N_13765,N_9432,N_9201);
or U13766 (N_13766,N_7530,N_10431);
nand U13767 (N_13767,N_11148,N_9861);
nand U13768 (N_13768,N_6554,N_10458);
xor U13769 (N_13769,N_9535,N_7137);
nand U13770 (N_13770,N_9165,N_11147);
or U13771 (N_13771,N_8293,N_8857);
and U13772 (N_13772,N_12006,N_8144);
nor U13773 (N_13773,N_6926,N_8091);
and U13774 (N_13774,N_10986,N_7134);
nor U13775 (N_13775,N_11086,N_10951);
or U13776 (N_13776,N_9681,N_8783);
xnor U13777 (N_13777,N_8644,N_10064);
xnor U13778 (N_13778,N_8150,N_7747);
xnor U13779 (N_13779,N_9577,N_7871);
and U13780 (N_13780,N_10593,N_7861);
nor U13781 (N_13781,N_8670,N_9398);
and U13782 (N_13782,N_9255,N_10367);
xor U13783 (N_13783,N_7956,N_10772);
and U13784 (N_13784,N_9304,N_11494);
and U13785 (N_13785,N_11451,N_11843);
or U13786 (N_13786,N_8500,N_7953);
xor U13787 (N_13787,N_7205,N_9478);
nor U13788 (N_13788,N_7594,N_10045);
and U13789 (N_13789,N_10084,N_7114);
nor U13790 (N_13790,N_11840,N_8493);
nor U13791 (N_13791,N_6260,N_9853);
xor U13792 (N_13792,N_6939,N_10200);
nor U13793 (N_13793,N_8978,N_11520);
nand U13794 (N_13794,N_12318,N_11634);
or U13795 (N_13795,N_12486,N_9283);
nand U13796 (N_13796,N_8051,N_7440);
or U13797 (N_13797,N_9714,N_8166);
xor U13798 (N_13798,N_9260,N_9250);
nand U13799 (N_13799,N_10744,N_9650);
nand U13800 (N_13800,N_11937,N_7363);
and U13801 (N_13801,N_7642,N_9875);
nor U13802 (N_13802,N_8736,N_12195);
xor U13803 (N_13803,N_11210,N_8188);
xor U13804 (N_13804,N_8496,N_7658);
or U13805 (N_13805,N_9254,N_10156);
nor U13806 (N_13806,N_9383,N_8551);
xnor U13807 (N_13807,N_8186,N_7631);
and U13808 (N_13808,N_6734,N_11259);
xnor U13809 (N_13809,N_7711,N_9981);
nor U13810 (N_13810,N_11241,N_8699);
xnor U13811 (N_13811,N_11093,N_8901);
and U13812 (N_13812,N_6791,N_8071);
or U13813 (N_13813,N_11186,N_7574);
xor U13814 (N_13814,N_7520,N_6456);
nand U13815 (N_13815,N_11195,N_8542);
nor U13816 (N_13816,N_12298,N_8511);
xor U13817 (N_13817,N_11111,N_10565);
and U13818 (N_13818,N_11748,N_6697);
or U13819 (N_13819,N_8983,N_9623);
and U13820 (N_13820,N_6271,N_7471);
xnor U13821 (N_13821,N_11734,N_9162);
and U13822 (N_13822,N_6613,N_7604);
nand U13823 (N_13823,N_8947,N_11861);
or U13824 (N_13824,N_8648,N_6608);
xnor U13825 (N_13825,N_12148,N_10946);
nor U13826 (N_13826,N_7962,N_12245);
nor U13827 (N_13827,N_6806,N_6621);
and U13828 (N_13828,N_12215,N_11067);
nand U13829 (N_13829,N_12136,N_10447);
nand U13830 (N_13830,N_11295,N_7269);
and U13831 (N_13831,N_10779,N_10090);
or U13832 (N_13832,N_9944,N_11501);
xor U13833 (N_13833,N_9246,N_12304);
xor U13834 (N_13834,N_9862,N_7126);
or U13835 (N_13835,N_8455,N_11852);
or U13836 (N_13836,N_8524,N_6604);
or U13837 (N_13837,N_10003,N_7074);
and U13838 (N_13838,N_8301,N_10824);
xor U13839 (N_13839,N_6512,N_10139);
or U13840 (N_13840,N_10653,N_11952);
or U13841 (N_13841,N_7959,N_7768);
or U13842 (N_13842,N_9543,N_11968);
or U13843 (N_13843,N_11792,N_7039);
nor U13844 (N_13844,N_10568,N_9068);
and U13845 (N_13845,N_9582,N_9636);
nand U13846 (N_13846,N_8935,N_10006);
nand U13847 (N_13847,N_11281,N_9071);
nor U13848 (N_13848,N_9789,N_6756);
and U13849 (N_13849,N_11053,N_9889);
nor U13850 (N_13850,N_8505,N_7391);
or U13851 (N_13851,N_11176,N_7734);
nor U13852 (N_13852,N_8688,N_8477);
and U13853 (N_13853,N_6896,N_12432);
xor U13854 (N_13854,N_11121,N_10326);
or U13855 (N_13855,N_10573,N_6872);
or U13856 (N_13856,N_9418,N_8407);
nor U13857 (N_13857,N_10557,N_9674);
and U13858 (N_13858,N_9225,N_9634);
nand U13859 (N_13859,N_6265,N_7620);
nand U13860 (N_13860,N_11666,N_6769);
nor U13861 (N_13861,N_7895,N_8863);
and U13862 (N_13862,N_7472,N_8079);
and U13863 (N_13863,N_10197,N_7826);
or U13864 (N_13864,N_7550,N_10798);
nand U13865 (N_13865,N_6966,N_10895);
or U13866 (N_13866,N_9067,N_9598);
and U13867 (N_13867,N_7037,N_6766);
and U13868 (N_13868,N_10416,N_12364);
nor U13869 (N_13869,N_7158,N_10602);
and U13870 (N_13870,N_9086,N_12078);
xnor U13871 (N_13871,N_9876,N_12201);
nand U13872 (N_13872,N_7672,N_9005);
xor U13873 (N_13873,N_10675,N_11122);
or U13874 (N_13874,N_12292,N_9422);
and U13875 (N_13875,N_7628,N_7080);
and U13876 (N_13876,N_7773,N_11882);
and U13877 (N_13877,N_7075,N_12094);
xor U13878 (N_13878,N_11340,N_10136);
nand U13879 (N_13879,N_11692,N_6660);
and U13880 (N_13880,N_11688,N_7811);
nand U13881 (N_13881,N_11078,N_9817);
nand U13882 (N_13882,N_11509,N_8789);
and U13883 (N_13883,N_11163,N_11717);
and U13884 (N_13884,N_10129,N_8765);
nand U13885 (N_13885,N_9675,N_10020);
nand U13886 (N_13886,N_10303,N_7930);
and U13887 (N_13887,N_6267,N_10058);
and U13888 (N_13888,N_9034,N_8421);
xnor U13889 (N_13889,N_8658,N_8024);
xnor U13890 (N_13890,N_8782,N_9557);
nand U13891 (N_13891,N_11826,N_7890);
and U13892 (N_13892,N_7589,N_7290);
nor U13893 (N_13893,N_8636,N_10117);
and U13894 (N_13894,N_9284,N_7592);
xnor U13895 (N_13895,N_10464,N_9734);
xnor U13896 (N_13896,N_6504,N_7382);
or U13897 (N_13897,N_10402,N_6856);
or U13898 (N_13898,N_6530,N_7771);
nor U13899 (N_13899,N_7197,N_11997);
xor U13900 (N_13900,N_9788,N_9621);
xor U13901 (N_13901,N_6709,N_9471);
nand U13902 (N_13902,N_8333,N_8107);
nor U13903 (N_13903,N_10841,N_10341);
and U13904 (N_13904,N_7236,N_9146);
nand U13905 (N_13905,N_6541,N_7846);
and U13906 (N_13906,N_11364,N_11232);
nand U13907 (N_13907,N_11473,N_9331);
and U13908 (N_13908,N_11296,N_10786);
xor U13909 (N_13909,N_7560,N_7599);
xor U13910 (N_13910,N_9407,N_12213);
or U13911 (N_13911,N_9048,N_11751);
or U13912 (N_13912,N_9332,N_8450);
or U13913 (N_13913,N_7901,N_8227);
nand U13914 (N_13914,N_9147,N_8429);
nor U13915 (N_13915,N_10055,N_11311);
or U13916 (N_13916,N_6587,N_7583);
xnor U13917 (N_13917,N_8216,N_10190);
nand U13918 (N_13918,N_11201,N_11627);
or U13919 (N_13919,N_7648,N_9829);
and U13920 (N_13920,N_6477,N_6929);
or U13921 (N_13921,N_10217,N_11385);
and U13922 (N_13922,N_6466,N_12300);
nor U13923 (N_13923,N_11847,N_8408);
nand U13924 (N_13924,N_11695,N_10371);
and U13925 (N_13925,N_7418,N_6564);
xnor U13926 (N_13926,N_11866,N_12015);
and U13927 (N_13927,N_10406,N_11192);
xor U13928 (N_13928,N_6694,N_9783);
nor U13929 (N_13929,N_11639,N_7539);
nor U13930 (N_13930,N_7086,N_9887);
or U13931 (N_13931,N_8824,N_7792);
nor U13932 (N_13932,N_7307,N_10685);
nor U13933 (N_13933,N_9884,N_7705);
nand U13934 (N_13934,N_12475,N_9063);
nor U13935 (N_13935,N_9725,N_6435);
nor U13936 (N_13936,N_8942,N_7798);
nor U13937 (N_13937,N_6612,N_7021);
nor U13938 (N_13938,N_6996,N_7265);
and U13939 (N_13939,N_6532,N_6632);
or U13940 (N_13940,N_6812,N_10554);
nor U13941 (N_13941,N_9591,N_8065);
nand U13942 (N_13942,N_9657,N_11193);
or U13943 (N_13943,N_8843,N_10921);
or U13944 (N_13944,N_10874,N_12071);
nor U13945 (N_13945,N_9547,N_9595);
xnor U13946 (N_13946,N_11716,N_10099);
or U13947 (N_13947,N_10152,N_11013);
nand U13948 (N_13948,N_11603,N_10882);
nand U13949 (N_13949,N_11411,N_10330);
or U13950 (N_13950,N_7174,N_9696);
xor U13951 (N_13951,N_7062,N_7789);
or U13952 (N_13952,N_6426,N_8430);
nor U13953 (N_13953,N_12247,N_6366);
and U13954 (N_13954,N_8681,N_10639);
nor U13955 (N_13955,N_6949,N_9340);
nand U13956 (N_13956,N_8516,N_6467);
and U13957 (N_13957,N_10864,N_6851);
or U13958 (N_13958,N_12261,N_11600);
nor U13959 (N_13959,N_9627,N_10995);
nand U13960 (N_13960,N_7291,N_7830);
or U13961 (N_13961,N_9455,N_8360);
nand U13962 (N_13962,N_6460,N_8002);
xnor U13963 (N_13963,N_10496,N_11648);
nor U13964 (N_13964,N_11375,N_10834);
and U13965 (N_13965,N_10654,N_7876);
xnor U13966 (N_13966,N_10884,N_11604);
or U13967 (N_13967,N_6510,N_8038);
xor U13968 (N_13968,N_11521,N_9631);
nand U13969 (N_13969,N_9616,N_6687);
or U13970 (N_13970,N_10794,N_11043);
xor U13971 (N_13971,N_7528,N_8585);
or U13972 (N_13972,N_9026,N_9819);
xnor U13973 (N_13973,N_8722,N_6647);
nand U13974 (N_13974,N_8401,N_6672);
and U13975 (N_13975,N_8952,N_10691);
or U13976 (N_13976,N_10828,N_7421);
and U13977 (N_13977,N_9840,N_9830);
nor U13978 (N_13978,N_8056,N_9281);
nor U13979 (N_13979,N_7218,N_8267);
nand U13980 (N_13980,N_10403,N_10342);
and U13981 (N_13981,N_11022,N_12175);
or U13982 (N_13982,N_10716,N_10393);
or U13983 (N_13983,N_10387,N_10945);
nand U13984 (N_13984,N_8701,N_8059);
nand U13985 (N_13985,N_8709,N_6485);
xor U13986 (N_13986,N_7921,N_11899);
and U13987 (N_13987,N_6699,N_10980);
nand U13988 (N_13988,N_12197,N_11481);
nand U13989 (N_13989,N_6508,N_6617);
or U13990 (N_13990,N_11558,N_8391);
nand U13991 (N_13991,N_6415,N_10269);
nor U13992 (N_13992,N_8625,N_6624);
or U13993 (N_13993,N_11280,N_6601);
xnor U13994 (N_13994,N_9519,N_10376);
xnor U13995 (N_13995,N_8295,N_6547);
xnor U13996 (N_13996,N_6642,N_10704);
or U13997 (N_13997,N_11158,N_9935);
nor U13998 (N_13998,N_10628,N_6596);
nand U13999 (N_13999,N_12028,N_10773);
nor U14000 (N_14000,N_10662,N_6556);
or U14001 (N_14001,N_10513,N_6507);
nand U14002 (N_14002,N_11654,N_8093);
xor U14003 (N_14003,N_10749,N_6398);
or U14004 (N_14004,N_11005,N_6676);
xor U14005 (N_14005,N_7942,N_8746);
nor U14006 (N_14006,N_12401,N_7054);
or U14007 (N_14007,N_6285,N_7778);
nor U14008 (N_14008,N_6615,N_9493);
or U14009 (N_14009,N_10849,N_6674);
xnor U14010 (N_14010,N_11088,N_8543);
nor U14011 (N_14011,N_10400,N_8844);
nor U14012 (N_14012,N_10116,N_12312);
xnor U14013 (N_14013,N_6449,N_7684);
xnor U14014 (N_14014,N_11314,N_10358);
xnor U14015 (N_14015,N_11403,N_8016);
xnor U14016 (N_14016,N_7634,N_11712);
and U14017 (N_14017,N_10302,N_6395);
and U14018 (N_14018,N_8341,N_8571);
nor U14019 (N_14019,N_8507,N_7326);
xor U14020 (N_14020,N_12479,N_7052);
nand U14021 (N_14021,N_7459,N_7173);
nor U14022 (N_14022,N_12096,N_7348);
and U14023 (N_14023,N_11954,N_9652);
xor U14024 (N_14024,N_8531,N_12467);
xor U14025 (N_14025,N_12463,N_11444);
xor U14026 (N_14026,N_9015,N_10918);
xnor U14027 (N_14027,N_11830,N_12189);
nor U14028 (N_14028,N_12207,N_8478);
or U14029 (N_14029,N_7110,N_7060);
and U14030 (N_14030,N_9534,N_9453);
and U14031 (N_14031,N_8894,N_9795);
or U14032 (N_14032,N_9149,N_8986);
xor U14033 (N_14033,N_8131,N_6420);
and U14034 (N_14034,N_7220,N_11042);
nor U14035 (N_14035,N_9601,N_10142);
nand U14036 (N_14036,N_10071,N_8141);
or U14037 (N_14037,N_10609,N_9114);
nor U14038 (N_14038,N_9197,N_11901);
and U14039 (N_14039,N_7727,N_7226);
or U14040 (N_14040,N_8228,N_9280);
xor U14041 (N_14041,N_9390,N_9466);
nand U14042 (N_14042,N_10929,N_8892);
nor U14043 (N_14043,N_10651,N_6797);
xnor U14044 (N_14044,N_10441,N_12122);
nand U14045 (N_14045,N_9381,N_10751);
xnor U14046 (N_14046,N_6488,N_10450);
or U14047 (N_14047,N_6778,N_8030);
or U14048 (N_14048,N_9343,N_6860);
or U14049 (N_14049,N_10392,N_12474);
nand U14050 (N_14050,N_7976,N_9792);
nor U14051 (N_14051,N_10008,N_9737);
and U14052 (N_14052,N_10705,N_9596);
xor U14053 (N_14053,N_7998,N_12228);
nand U14054 (N_14054,N_7888,N_9152);
xnor U14055 (N_14055,N_10766,N_11848);
or U14056 (N_14056,N_11897,N_7308);
nor U14057 (N_14057,N_9293,N_6350);
nand U14058 (N_14058,N_9852,N_10126);
nand U14059 (N_14059,N_8706,N_9559);
nand U14060 (N_14060,N_7243,N_8871);
nor U14061 (N_14061,N_7398,N_11785);
nand U14062 (N_14062,N_11548,N_10443);
nor U14063 (N_14063,N_8628,N_11343);
nor U14064 (N_14064,N_8072,N_9615);
xnor U14065 (N_14065,N_8643,N_8092);
or U14066 (N_14066,N_10095,N_10732);
nor U14067 (N_14067,N_12119,N_6755);
nand U14068 (N_14068,N_7051,N_7004);
and U14069 (N_14069,N_12423,N_12239);
nor U14070 (N_14070,N_8760,N_7898);
nor U14071 (N_14071,N_12191,N_6280);
xnor U14072 (N_14072,N_7554,N_9694);
nor U14073 (N_14073,N_12357,N_10347);
and U14074 (N_14074,N_8146,N_8189);
nand U14075 (N_14075,N_11672,N_8988);
xor U14076 (N_14076,N_8118,N_10215);
nand U14077 (N_14077,N_11527,N_9228);
nor U14078 (N_14078,N_11851,N_10132);
or U14079 (N_14079,N_7954,N_12160);
nor U14080 (N_14080,N_7755,N_11349);
nor U14081 (N_14081,N_7982,N_10763);
nor U14082 (N_14082,N_11553,N_9377);
nand U14083 (N_14083,N_12273,N_8692);
and U14084 (N_14084,N_6897,N_11810);
and U14085 (N_14085,N_11683,N_9872);
and U14086 (N_14086,N_8286,N_8162);
and U14087 (N_14087,N_8833,N_10796);
or U14088 (N_14088,N_9111,N_9833);
or U14089 (N_14089,N_12135,N_9561);
or U14090 (N_14090,N_9051,N_9365);
nand U14091 (N_14091,N_9102,N_10096);
xnor U14092 (N_14092,N_12480,N_12064);
or U14093 (N_14093,N_6381,N_10218);
nand U14094 (N_14094,N_6261,N_11761);
and U14095 (N_14095,N_6757,N_9804);
xor U14096 (N_14096,N_11526,N_8208);
xnor U14097 (N_14097,N_7698,N_7312);
nor U14098 (N_14098,N_11085,N_11544);
nor U14099 (N_14099,N_11569,N_10273);
or U14100 (N_14100,N_8126,N_8218);
or U14101 (N_14101,N_8127,N_12005);
and U14102 (N_14102,N_11665,N_8817);
nor U14103 (N_14103,N_11987,N_12324);
nor U14104 (N_14104,N_6824,N_10833);
xor U14105 (N_14105,N_6867,N_11405);
nand U14106 (N_14106,N_9752,N_11347);
xnor U14107 (N_14107,N_7862,N_11571);
and U14108 (N_14108,N_7318,N_9019);
xnor U14109 (N_14109,N_9282,N_6292);
nand U14110 (N_14110,N_9603,N_7630);
or U14111 (N_14111,N_8268,N_7614);
nor U14112 (N_14112,N_9391,N_11395);
or U14113 (N_14113,N_9327,N_7341);
or U14114 (N_14114,N_12406,N_12315);
and U14115 (N_14115,N_8492,N_10563);
nand U14116 (N_14116,N_11824,N_8963);
and U14117 (N_14117,N_12107,N_9265);
nand U14118 (N_14118,N_10123,N_10059);
and U14119 (N_14119,N_9644,N_8317);
nand U14120 (N_14120,N_7541,N_12170);
and U14121 (N_14121,N_9148,N_12258);
and U14122 (N_14122,N_11248,N_11307);
nor U14123 (N_14123,N_6909,N_11790);
or U14124 (N_14124,N_9105,N_8879);
xor U14125 (N_14125,N_11704,N_12146);
nand U14126 (N_14126,N_6998,N_10655);
or U14127 (N_14127,N_6574,N_6651);
or U14128 (N_14128,N_10194,N_7026);
nor U14129 (N_14129,N_9902,N_10470);
nor U14130 (N_14130,N_6590,N_11804);
and U14131 (N_14131,N_10220,N_7920);
and U14132 (N_14132,N_6605,N_7138);
xor U14133 (N_14133,N_7402,N_8887);
and U14134 (N_14134,N_12212,N_7354);
nor U14135 (N_14135,N_8876,N_11902);
xnor U14136 (N_14136,N_6368,N_10840);
and U14137 (N_14137,N_10971,N_7030);
nand U14138 (N_14138,N_8664,N_8319);
or U14139 (N_14139,N_12320,N_11638);
nor U14140 (N_14140,N_7204,N_8592);
or U14141 (N_14141,N_7227,N_10666);
nand U14142 (N_14142,N_7878,N_6463);
nand U14143 (N_14143,N_10373,N_11212);
nor U14144 (N_14144,N_6895,N_10891);
nor U14145 (N_14145,N_7807,N_9328);
or U14146 (N_14146,N_8602,N_7569);
nor U14147 (N_14147,N_11030,N_10315);
nand U14148 (N_14148,N_12011,N_6957);
or U14149 (N_14149,N_11649,N_7601);
nor U14150 (N_14150,N_7314,N_7855);
xor U14151 (N_14151,N_10721,N_12008);
and U14152 (N_14152,N_9868,N_6950);
or U14153 (N_14153,N_11136,N_7403);
and U14154 (N_14154,N_8954,N_7185);
nor U14155 (N_14155,N_9131,N_12427);
and U14156 (N_14156,N_9414,N_11557);
nor U14157 (N_14157,N_12280,N_11862);
nor U14158 (N_14158,N_9354,N_8164);
or U14159 (N_14159,N_10996,N_11264);
nand U14160 (N_14160,N_7638,N_10177);
or U14161 (N_14161,N_6353,N_10926);
and U14162 (N_14162,N_7717,N_8062);
and U14163 (N_14163,N_12091,N_12130);
nand U14164 (N_14164,N_12310,N_9941);
or U14165 (N_14165,N_9144,N_11773);
or U14166 (N_14166,N_12394,N_10922);
nor U14167 (N_14167,N_10983,N_8759);
or U14168 (N_14168,N_10941,N_12100);
nor U14169 (N_14169,N_12075,N_9998);
xor U14170 (N_14170,N_6973,N_9321);
nand U14171 (N_14171,N_9489,N_9009);
nor U14172 (N_14172,N_11940,N_8364);
nand U14173 (N_14173,N_6997,N_11747);
or U14174 (N_14174,N_8927,N_11680);
nand U14175 (N_14175,N_6303,N_11044);
xnor U14176 (N_14176,N_8423,N_7675);
xnor U14177 (N_14177,N_12089,N_6977);
nor U14178 (N_14178,N_10801,N_10740);
nand U14179 (N_14179,N_9062,N_7238);
nand U14180 (N_14180,N_9462,N_7977);
and U14181 (N_14181,N_9579,N_9947);
or U14182 (N_14182,N_9746,N_11733);
and U14183 (N_14183,N_11092,N_9990);
nand U14184 (N_14184,N_6548,N_10683);
nor U14185 (N_14185,N_6389,N_6914);
or U14186 (N_14186,N_9826,N_12131);
xor U14187 (N_14187,N_11669,N_11409);
xnor U14188 (N_14188,N_11605,N_12325);
xor U14189 (N_14189,N_8357,N_12265);
xor U14190 (N_14190,N_6324,N_9029);
and U14191 (N_14191,N_11621,N_9241);
or U14192 (N_14192,N_8195,N_7241);
or U14193 (N_14193,N_12018,N_7442);
nand U14194 (N_14194,N_10171,N_9578);
nor U14195 (N_14195,N_9914,N_12353);
and U14196 (N_14196,N_10657,N_7553);
nor U14197 (N_14197,N_11227,N_6256);
xor U14198 (N_14198,N_9790,N_7827);
xor U14199 (N_14199,N_12349,N_9880);
xnor U14200 (N_14200,N_10904,N_6761);
nor U14201 (N_14201,N_11572,N_10626);
xor U14202 (N_14202,N_9199,N_6361);
nand U14203 (N_14203,N_7474,N_6967);
and U14204 (N_14204,N_11988,N_9369);
nor U14205 (N_14205,N_11034,N_6332);
and U14206 (N_14206,N_7331,N_8902);
xnor U14207 (N_14207,N_11957,N_6304);
nand U14208 (N_14208,N_9881,N_10782);
xor U14209 (N_14209,N_9424,N_10521);
and U14210 (N_14210,N_8840,N_9324);
xor U14211 (N_14211,N_9515,N_12070);
and U14212 (N_14212,N_10499,N_7338);
nor U14213 (N_14213,N_10384,N_7358);
xor U14214 (N_14214,N_10700,N_10601);
xor U14215 (N_14215,N_11001,N_9866);
and U14216 (N_14216,N_11755,N_6862);
and U14217 (N_14217,N_10897,N_7851);
nor U14218 (N_14218,N_9411,N_10676);
nor U14219 (N_14219,N_8624,N_8471);
nand U14220 (N_14220,N_12477,N_10610);
nor U14221 (N_14221,N_9208,N_7581);
xnor U14222 (N_14222,N_10767,N_6539);
nor U14223 (N_14223,N_8487,N_8379);
or U14224 (N_14224,N_10880,N_12308);
nand U14225 (N_14225,N_8106,N_7322);
nor U14226 (N_14226,N_10611,N_6744);
and U14227 (N_14227,N_12430,N_7098);
and U14228 (N_14228,N_6451,N_9668);
or U14229 (N_14229,N_7108,N_9964);
and U14230 (N_14230,N_6667,N_9141);
xnor U14231 (N_14231,N_9689,N_7913);
nor U14232 (N_14232,N_7995,N_12138);
and U14233 (N_14233,N_8725,N_11224);
or U14234 (N_14234,N_12125,N_12223);
nor U14235 (N_14235,N_9630,N_8037);
nand U14236 (N_14236,N_7452,N_9618);
nand U14237 (N_14237,N_8796,N_9457);
nand U14238 (N_14238,N_8235,N_9776);
or U14239 (N_14239,N_11786,N_7914);
and U14240 (N_14240,N_6714,N_8679);
nor U14241 (N_14241,N_7001,N_8264);
and U14242 (N_14242,N_8448,N_6362);
xor U14243 (N_14243,N_7147,N_10863);
nand U14244 (N_14244,N_12072,N_9870);
and U14245 (N_14245,N_9637,N_10669);
nand U14246 (N_14246,N_11821,N_12240);
xnor U14247 (N_14247,N_10814,N_7081);
and U14248 (N_14248,N_11027,N_10378);
nand U14249 (N_14249,N_11381,N_6794);
or U14250 (N_14250,N_10999,N_11663);
and U14251 (N_14251,N_11829,N_9513);
xnor U14252 (N_14252,N_11342,N_11226);
xnor U14253 (N_14253,N_10643,N_8431);
nor U14254 (N_14254,N_10892,N_9375);
nor U14255 (N_14255,N_11757,N_10831);
nor U14256 (N_14256,N_11878,N_7602);
nand U14257 (N_14257,N_8307,N_12051);
or U14258 (N_14258,N_11927,N_8007);
and U14259 (N_14259,N_7889,N_6302);
xnor U14260 (N_14260,N_11845,N_8982);
nand U14261 (N_14261,N_6786,N_7369);
xor U14262 (N_14262,N_12050,N_6663);
nor U14263 (N_14263,N_7143,N_7342);
nand U14264 (N_14264,N_12392,N_7810);
and U14265 (N_14265,N_8020,N_10306);
nand U14266 (N_14266,N_11709,N_10701);
nor U14267 (N_14267,N_7533,N_9705);
or U14268 (N_14268,N_12159,N_7752);
xor U14269 (N_14269,N_8773,N_9984);
nand U14270 (N_14270,N_10282,N_7355);
or U14271 (N_14271,N_8769,N_7103);
xnor U14272 (N_14272,N_7011,N_11771);
or U14273 (N_14273,N_8539,N_9484);
or U14274 (N_14274,N_6571,N_8917);
and U14275 (N_14275,N_12433,N_8419);
or U14276 (N_14276,N_9116,N_8251);
nor U14277 (N_14277,N_11889,N_12424);
xor U14278 (N_14278,N_7065,N_7361);
and U14279 (N_14279,N_10340,N_6575);
nand U14280 (N_14280,N_9765,N_11152);
nor U14281 (N_14281,N_10546,N_6817);
nand U14282 (N_14282,N_7047,N_7909);
nand U14283 (N_14283,N_7016,N_9575);
nor U14284 (N_14284,N_10590,N_9978);
and U14285 (N_14285,N_7597,N_9302);
or U14286 (N_14286,N_10349,N_11235);
or U14287 (N_14287,N_11999,N_9222);
xor U14288 (N_14288,N_9093,N_10482);
nor U14289 (N_14289,N_10903,N_9504);
and U14290 (N_14290,N_7573,N_7094);
and U14291 (N_14291,N_9458,N_9506);
or U14292 (N_14292,N_6440,N_9270);
nor U14293 (N_14293,N_8784,N_6409);
nor U14294 (N_14294,N_10872,N_8204);
nor U14295 (N_14295,N_7229,N_11677);
xor U14296 (N_14296,N_6788,N_9546);
and U14297 (N_14297,N_9857,N_11433);
xor U14298 (N_14298,N_8694,N_11009);
and U14299 (N_14299,N_11378,N_6637);
nor U14300 (N_14300,N_8964,N_7575);
xor U14301 (N_14301,N_10690,N_10961);
or U14302 (N_14302,N_8381,N_8167);
and U14303 (N_14303,N_8647,N_11825);
and U14304 (N_14304,N_9310,N_10390);
xnor U14305 (N_14305,N_10164,N_12080);
nor U14306 (N_14306,N_10990,N_10354);
and U14307 (N_14307,N_8128,N_10510);
or U14308 (N_14308,N_10500,N_7896);
or U14309 (N_14309,N_9762,N_8974);
and U14310 (N_14310,N_11835,N_7470);
or U14311 (N_14311,N_11881,N_10504);
nand U14312 (N_14312,N_10070,N_6379);
xor U14313 (N_14313,N_12023,N_10949);
or U14314 (N_14314,N_6382,N_11528);
nand U14315 (N_14315,N_12210,N_8522);
and U14316 (N_14316,N_6962,N_7656);
nand U14317 (N_14317,N_10312,N_8836);
or U14318 (N_14318,N_10209,N_7165);
xor U14319 (N_14319,N_12485,N_7413);
or U14320 (N_14320,N_10044,N_6472);
or U14321 (N_14321,N_9500,N_7256);
nand U14322 (N_14322,N_7859,N_11823);
and U14323 (N_14323,N_8129,N_9832);
and U14324 (N_14324,N_10909,N_10150);
and U14325 (N_14325,N_8143,N_9570);
and U14326 (N_14326,N_6558,N_8997);
xor U14327 (N_14327,N_7552,N_7230);
xnor U14328 (N_14328,N_11061,N_9699);
nor U14329 (N_14329,N_11090,N_11644);
and U14330 (N_14330,N_8584,N_11652);
nor U14331 (N_14331,N_10974,N_10083);
xnor U14332 (N_14332,N_10784,N_11292);
nor U14333 (N_14333,N_9277,N_12278);
xor U14334 (N_14334,N_10329,N_10962);
and U14335 (N_14335,N_9973,N_9687);
and U14336 (N_14336,N_8737,N_10286);
or U14337 (N_14337,N_8504,N_12476);
xor U14338 (N_14338,N_6281,N_9778);
nand U14339 (N_14339,N_10372,N_6903);
xor U14340 (N_14340,N_9115,N_11661);
and U14341 (N_14341,N_11890,N_6407);
and U14342 (N_14342,N_6726,N_7587);
xnor U14343 (N_14343,N_6863,N_10085);
xor U14344 (N_14344,N_11567,N_6891);
or U14345 (N_14345,N_6724,N_8575);
xnor U14346 (N_14346,N_8577,N_10408);
xor U14347 (N_14347,N_11362,N_7028);
nand U14348 (N_14348,N_6550,N_10339);
nand U14349 (N_14349,N_8099,N_9501);
nand U14350 (N_14350,N_6333,N_7937);
or U14351 (N_14351,N_8872,N_6376);
and U14352 (N_14352,N_10242,N_8712);
xnor U14353 (N_14353,N_9376,N_7444);
or U14354 (N_14354,N_7984,N_7414);
or U14355 (N_14355,N_8358,N_10198);
nor U14356 (N_14356,N_7582,N_8310);
nor U14357 (N_14357,N_7780,N_11142);
and U14358 (N_14358,N_9016,N_9667);
xor U14359 (N_14359,N_8785,N_8946);
nand U14360 (N_14360,N_11102,N_6974);
and U14361 (N_14361,N_11079,N_8316);
nand U14362 (N_14362,N_11369,N_9933);
and U14363 (N_14363,N_7681,N_9198);
xor U14364 (N_14364,N_10603,N_8775);
and U14365 (N_14365,N_12359,N_11286);
and U14366 (N_14366,N_8245,N_8931);
and U14367 (N_14367,N_11989,N_12378);
nor U14368 (N_14368,N_11749,N_12365);
and U14369 (N_14369,N_10314,N_9821);
nand U14370 (N_14370,N_7845,N_7240);
xnor U14371 (N_14371,N_9055,N_9923);
xor U14372 (N_14372,N_11221,N_11262);
nor U14373 (N_14373,N_11766,N_7908);
nand U14374 (N_14374,N_7608,N_7385);
nor U14375 (N_14375,N_11535,N_9140);
nand U14376 (N_14376,N_7079,N_8629);
and U14377 (N_14377,N_11284,N_8252);
or U14378 (N_14378,N_10426,N_9594);
or U14379 (N_14379,N_7378,N_6855);
and U14380 (N_14380,N_8874,N_7952);
nand U14381 (N_14381,N_7450,N_9784);
or U14382 (N_14382,N_8734,N_7749);
and U14383 (N_14383,N_7365,N_8704);
xnor U14384 (N_14384,N_11076,N_11950);
nand U14385 (N_14385,N_12302,N_11162);
or U14386 (N_14386,N_8646,N_8953);
nand U14387 (N_14387,N_10388,N_8719);
or U14388 (N_14388,N_7311,N_7886);
and U14389 (N_14389,N_6540,N_9450);
and U14390 (N_14390,N_9721,N_9949);
xor U14391 (N_14391,N_7750,N_11172);
nand U14392 (N_14392,N_7130,N_6380);
nand U14393 (N_14393,N_11976,N_9193);
xnor U14394 (N_14394,N_7665,N_10567);
and U14395 (N_14395,N_11319,N_11428);
or U14396 (N_14396,N_11576,N_9882);
and U14397 (N_14397,N_10726,N_9221);
nor U14398 (N_14398,N_7933,N_7932);
or U14399 (N_14399,N_6882,N_11803);
or U14400 (N_14400,N_10978,N_11974);
xnor U14401 (N_14401,N_8720,N_10693);
nor U14402 (N_14402,N_7880,N_11961);
nand U14403 (N_14403,N_7033,N_8372);
nand U14404 (N_14404,N_6453,N_8651);
and U14405 (N_14405,N_11151,N_6742);
and U14406 (N_14406,N_7699,N_6764);
nor U14407 (N_14407,N_7186,N_8096);
and U14408 (N_14408,N_10774,N_11384);
nand U14409 (N_14409,N_10480,N_8180);
nor U14410 (N_14410,N_9770,N_9342);
and U14411 (N_14411,N_11175,N_11256);
and U14412 (N_14412,N_8936,N_6316);
nor U14413 (N_14413,N_11497,N_6589);
or U14414 (N_14414,N_8993,N_6787);
nor U14415 (N_14415,N_7683,N_8510);
nand U14416 (N_14416,N_8354,N_7973);
nand U14417 (N_14417,N_9750,N_9846);
and U14418 (N_14418,N_10000,N_10174);
nand U14419 (N_14419,N_7806,N_11297);
xnor U14420 (N_14420,N_9074,N_10644);
xor U14421 (N_14421,N_7456,N_6525);
xnor U14422 (N_14422,N_7963,N_11983);
nor U14423 (N_14423,N_6300,N_11062);
or U14424 (N_14424,N_8243,N_10241);
xnor U14425 (N_14425,N_11191,N_7462);
or U14426 (N_14426,N_11353,N_7303);
or U14427 (N_14427,N_11924,N_9508);
xnor U14428 (N_14428,N_10511,N_6745);
nor U14429 (N_14429,N_10631,N_8780);
xnor U14430 (N_14430,N_11420,N_8201);
or U14431 (N_14431,N_6343,N_9612);
xnor U14432 (N_14432,N_9735,N_11964);
nand U14433 (N_14433,N_6639,N_7677);
nor U14434 (N_14434,N_10907,N_7072);
and U14435 (N_14435,N_6874,N_7262);
and U14436 (N_14436,N_11701,N_8377);
or U14437 (N_14437,N_6314,N_7247);
nand U14438 (N_14438,N_9261,N_11217);
and U14439 (N_14439,N_9858,N_7992);
and U14440 (N_14440,N_10423,N_12282);
or U14441 (N_14441,N_11598,N_6796);
xnor U14442 (N_14442,N_10049,N_7208);
or U14443 (N_14443,N_11724,N_7529);
and U14444 (N_14444,N_8057,N_10255);
and U14445 (N_14445,N_7578,N_11020);
xnor U14446 (N_14446,N_7721,N_8919);
and U14447 (N_14447,N_9370,N_8439);
xor U14448 (N_14448,N_10692,N_7381);
or U14449 (N_14449,N_8175,N_11659);
or U14450 (N_14450,N_6971,N_9426);
and U14451 (N_14451,N_11583,N_10410);
or U14452 (N_14452,N_9673,N_10861);
or U14453 (N_14453,N_7477,N_8330);
nand U14454 (N_14454,N_10289,N_12264);
and U14455 (N_14455,N_6736,N_7187);
and U14456 (N_14456,N_8156,N_7475);
or U14457 (N_14457,N_9633,N_6501);
or U14458 (N_14458,N_8266,N_11689);
xor U14459 (N_14459,N_8950,N_7107);
or U14460 (N_14460,N_7874,N_11762);
nor U14461 (N_14461,N_11593,N_9339);
xnor U14462 (N_14462,N_8600,N_8702);
or U14463 (N_14463,N_7484,N_9825);
nor U14464 (N_14464,N_10620,N_11004);
nor U14465 (N_14465,N_6969,N_9976);
and U14466 (N_14466,N_11396,N_10501);
nand U14467 (N_14467,N_11051,N_8713);
nand U14468 (N_14468,N_10271,N_7680);
or U14469 (N_14469,N_7881,N_7024);
nand U14470 (N_14470,N_6401,N_10910);
or U14471 (N_14471,N_11768,N_10485);
xnor U14472 (N_14472,N_7272,N_7175);
and U14473 (N_14473,N_7299,N_8751);
xnor U14474 (N_14474,N_7716,N_7640);
nand U14475 (N_14475,N_12397,N_8891);
nor U14476 (N_14476,N_10621,N_9683);
or U14477 (N_14477,N_6983,N_8607);
and U14478 (N_14478,N_10025,N_12496);
nor U14479 (N_14479,N_8009,N_11503);
xor U14480 (N_14480,N_10919,N_11410);
or U14481 (N_14481,N_7401,N_9109);
and U14482 (N_14482,N_7077,N_9206);
and U14483 (N_14483,N_8933,N_10965);
xnor U14484 (N_14484,N_6870,N_10001);
nor U14485 (N_14485,N_11275,N_6542);
nand U14486 (N_14486,N_7639,N_9576);
xor U14487 (N_14487,N_11203,N_7618);
or U14488 (N_14488,N_11012,N_11559);
xnor U14489 (N_14489,N_8895,N_8514);
nand U14490 (N_14490,N_6278,N_11084);
nand U14491 (N_14491,N_11645,N_7343);
xnor U14492 (N_14492,N_11972,N_11922);
nand U14493 (N_14493,N_10246,N_7788);
nor U14494 (N_14494,N_12462,N_11574);
nor U14495 (N_14495,N_11159,N_12198);
xnor U14496 (N_14496,N_9358,N_10290);
or U14497 (N_14497,N_12219,N_6329);
or U14498 (N_14498,N_10595,N_8924);
xor U14499 (N_14499,N_11758,N_7662);
xnor U14500 (N_14500,N_9425,N_11161);
nand U14501 (N_14501,N_11582,N_9167);
nand U14502 (N_14502,N_9217,N_7857);
nand U14503 (N_14503,N_6876,N_9176);
or U14504 (N_14504,N_8848,N_9995);
and U14505 (N_14505,N_8069,N_12466);
nor U14506 (N_14506,N_7445,N_8589);
nor U14507 (N_14507,N_6631,N_8735);
nor U14508 (N_14508,N_11125,N_10889);
xor U14509 (N_14509,N_11493,N_8790);
nand U14510 (N_14510,N_11242,N_10756);
nand U14511 (N_14511,N_10395,N_12388);
nor U14512 (N_14512,N_9388,N_10079);
nor U14513 (N_14513,N_11513,N_7585);
and U14514 (N_14514,N_10257,N_11910);
nor U14515 (N_14515,N_6405,N_8654);
xor U14516 (N_14516,N_8284,N_9188);
xor U14517 (N_14517,N_8304,N_9763);
or U14518 (N_14518,N_8275,N_8249);
or U14519 (N_14519,N_8650,N_7879);
nor U14520 (N_14520,N_7739,N_9911);
xor U14521 (N_14521,N_7255,N_11651);
or U14522 (N_14522,N_11074,N_7668);
xor U14523 (N_14523,N_12082,N_8211);
xnor U14524 (N_14524,N_8870,N_9867);
or U14525 (N_14525,N_11060,N_10144);
nand U14526 (N_14526,N_9291,N_6702);
nand U14527 (N_14527,N_11994,N_12497);
or U14528 (N_14528,N_10451,N_10894);
nor U14529 (N_14529,N_8489,N_10761);
nor U14530 (N_14530,N_8393,N_8529);
and U14531 (N_14531,N_7770,N_10281);
nor U14532 (N_14532,N_6489,N_8944);
nor U14533 (N_14533,N_9813,N_11658);
nor U14534 (N_14534,N_6342,N_6563);
nand U14535 (N_14535,N_10192,N_9312);
or U14536 (N_14536,N_6334,N_9448);
nand U14537 (N_14537,N_11515,N_6741);
xor U14538 (N_14538,N_8550,N_8595);
nor U14539 (N_14539,N_7719,N_8989);
or U14540 (N_14540,N_8581,N_10992);
xnor U14541 (N_14541,N_6681,N_11626);
nand U14542 (N_14542,N_6737,N_9166);
and U14543 (N_14543,N_8880,N_10024);
or U14544 (N_14544,N_10313,N_6808);
or U14545 (N_14545,N_8962,N_9043);
xnor U14546 (N_14546,N_10645,N_9945);
nand U14547 (N_14547,N_11462,N_10998);
xnor U14548 (N_14548,N_11141,N_9087);
or U14549 (N_14549,N_9663,N_6846);
xor U14550 (N_14550,N_6308,N_6735);
nor U14551 (N_14551,N_6372,N_11674);
xor U14552 (N_14552,N_10984,N_8122);
nor U14553 (N_14553,N_10134,N_8977);
nand U14554 (N_14554,N_11299,N_11097);
xnor U14555 (N_14555,N_11324,N_10157);
xor U14556 (N_14556,N_6749,N_8710);
xnor U14557 (N_14557,N_8979,N_6841);
xor U14558 (N_14558,N_12498,N_7190);
nand U14559 (N_14559,N_9037,N_9289);
or U14560 (N_14560,N_6317,N_10741);
nand U14561 (N_14561,N_7799,N_9006);
xor U14562 (N_14562,N_12343,N_7410);
or U14563 (N_14563,N_10790,N_6802);
and U14564 (N_14564,N_6520,N_8464);
and U14565 (N_14565,N_8972,N_6633);
xnor U14566 (N_14566,N_12241,N_9540);
nor U14567 (N_14567,N_11278,N_6611);
nand U14568 (N_14568,N_9926,N_8718);
or U14569 (N_14569,N_9711,N_8221);
nand U14570 (N_14570,N_7375,N_9572);
and U14571 (N_14571,N_11556,N_8981);
xnor U14572 (N_14572,N_9948,N_9865);
and U14573 (N_14573,N_12287,N_6599);
nor U14574 (N_14574,N_7852,N_12145);
or U14575 (N_14575,N_10780,N_10809);
nand U14576 (N_14576,N_8083,N_9056);
nor U14577 (N_14577,N_9104,N_9218);
xor U14578 (N_14578,N_11129,N_8729);
and U14579 (N_14579,N_10777,N_10063);
xnor U14580 (N_14580,N_12238,N_11681);
nand U14581 (N_14581,N_12478,N_6904);
and U14582 (N_14582,N_10486,N_9264);
xor U14583 (N_14583,N_8417,N_11492);
or U14584 (N_14584,N_11930,N_8657);
nor U14585 (N_14585,N_7492,N_8923);
or U14586 (N_14586,N_8011,N_12361);
or U14587 (N_14587,N_10027,N_8338);
and U14588 (N_14588,N_10165,N_7155);
nand U14589 (N_14589,N_12150,N_12262);
xnor U14590 (N_14590,N_12002,N_7359);
nand U14591 (N_14591,N_12114,N_10723);
or U14592 (N_14592,N_10747,N_8313);
or U14593 (N_14593,N_10106,N_11943);
xor U14594 (N_14594,N_7424,N_10012);
or U14595 (N_14595,N_8753,N_8873);
or U14596 (N_14596,N_11711,N_6684);
xnor U14597 (N_14597,N_7356,N_7991);
or U14598 (N_14598,N_11566,N_8598);
nand U14599 (N_14599,N_12368,N_6424);
nor U14600 (N_14600,N_9428,N_9883);
nor U14601 (N_14601,N_8485,N_9427);
nand U14602 (N_14602,N_10125,N_8869);
nor U14603 (N_14603,N_9491,N_7893);
nand U14604 (N_14604,N_10411,N_8951);
or U14605 (N_14605,N_12199,N_9049);
nand U14606 (N_14606,N_6496,N_10016);
or U14607 (N_14607,N_7867,N_7548);
nor U14608 (N_14608,N_8745,N_6923);
nand U14609 (N_14609,N_7903,N_10258);
or U14610 (N_14610,N_6492,N_6327);
and U14611 (N_14611,N_6370,N_8573);
xnor U14612 (N_14612,N_7939,N_10966);
or U14613 (N_14613,N_6963,N_8135);
or U14614 (N_14614,N_10316,N_10730);
and U14615 (N_14615,N_8437,N_8105);
or U14616 (N_14616,N_6729,N_9946);
nand U14617 (N_14617,N_9070,N_11706);
nor U14618 (N_14618,N_11485,N_10958);
xor U14619 (N_14619,N_8806,N_10616);
xnor U14620 (N_14620,N_11874,N_7483);
xor U14621 (N_14621,N_7157,N_11108);
nand U14622 (N_14622,N_6584,N_11587);
xnor U14623 (N_14623,N_6418,N_10184);
and U14624 (N_14624,N_7935,N_8000);
and U14625 (N_14625,N_11190,N_8606);
nor U14626 (N_14626,N_11112,N_11225);
nor U14627 (N_14627,N_12227,N_7600);
or U14628 (N_14628,N_9089,N_10673);
or U14629 (N_14629,N_6905,N_9797);
and U14630 (N_14630,N_6819,N_12405);
xor U14631 (N_14631,N_10711,N_7869);
xnor U14632 (N_14632,N_11188,N_7066);
xor U14633 (N_14633,N_10112,N_10571);
and U14634 (N_14634,N_6915,N_6646);
xor U14635 (N_14635,N_11003,N_8528);
nand U14636 (N_14636,N_6419,N_9175);
and U14637 (N_14637,N_7070,N_11260);
xnor U14638 (N_14638,N_11887,N_12182);
or U14639 (N_14639,N_9210,N_11368);
xor U14640 (N_14640,N_10119,N_10072);
or U14641 (N_14641,N_10665,N_9904);
nand U14642 (N_14642,N_8966,N_7812);
nand U14643 (N_14643,N_10553,N_9290);
xnor U14644 (N_14644,N_9845,N_7198);
nand U14645 (N_14645,N_6859,N_8420);
nor U14646 (N_14646,N_12147,N_12450);
nand U14647 (N_14647,N_7149,N_12190);
or U14648 (N_14648,N_10498,N_11993);
nor U14649 (N_14649,N_10792,N_6363);
and U14650 (N_14650,N_9066,N_8003);
or U14651 (N_14651,N_6685,N_11868);
nor U14652 (N_14652,N_9992,N_12065);
and U14653 (N_14653,N_6775,N_9971);
or U14654 (N_14654,N_6371,N_7139);
or U14655 (N_14655,N_7790,N_7104);
nor U14656 (N_14656,N_10092,N_10928);
xor U14657 (N_14657,N_7435,N_6331);
xor U14658 (N_14658,N_6486,N_7723);
xor U14659 (N_14659,N_10127,N_11953);
or U14660 (N_14660,N_11054,N_10802);
xnor U14661 (N_14661,N_10013,N_8590);
xor U14662 (N_14662,N_10967,N_10291);
and U14663 (N_14663,N_9474,N_10404);
xor U14664 (N_14664,N_12126,N_7244);
xor U14665 (N_14665,N_9400,N_8798);
or U14666 (N_14666,N_10632,N_9720);
nor U14667 (N_14667,N_10613,N_6473);
nor U14668 (N_14668,N_6388,N_8596);
and U14669 (N_14669,N_11738,N_10300);
nand U14670 (N_14670,N_9274,N_10087);
and U14671 (N_14671,N_11018,N_9421);
and U14672 (N_14672,N_11269,N_11519);
or U14673 (N_14673,N_7148,N_6299);
nor U14674 (N_14674,N_12334,N_7870);
and U14675 (N_14675,N_7906,N_10528);
nand U14676 (N_14676,N_10871,N_6535);
or U14677 (N_14677,N_10128,N_9271);
nor U14678 (N_14678,N_7865,N_6543);
nor U14679 (N_14679,N_8616,N_7280);
nor U14680 (N_14680,N_11048,N_11880);
nor U14681 (N_14681,N_10917,N_9399);
nor U14682 (N_14682,N_9357,N_11895);
and U14683 (N_14683,N_11532,N_10775);
nor U14684 (N_14684,N_9212,N_10908);
xnor U14685 (N_14685,N_9958,N_8787);
xor U14686 (N_14686,N_6898,N_7715);
or U14687 (N_14687,N_6503,N_10604);
and U14688 (N_14688,N_11948,N_7364);
nor U14689 (N_14689,N_6476,N_7352);
or U14690 (N_14690,N_12254,N_12422);
and U14691 (N_14691,N_10641,N_9256);
nand U14692 (N_14692,N_9913,N_10608);
and U14693 (N_14693,N_8669,N_7071);
xor U14694 (N_14694,N_12279,N_10561);
nor U14695 (N_14695,N_9974,N_7781);
xnor U14696 (N_14696,N_6480,N_9972);
nor U14697 (N_14697,N_6594,N_7457);
nor U14698 (N_14698,N_10497,N_8327);
and U14699 (N_14699,N_11858,N_10868);
xnor U14700 (N_14700,N_8412,N_11590);
and U14701 (N_14701,N_6673,N_7076);
nor U14702 (N_14702,N_8890,N_11470);
and U14703 (N_14703,N_7493,N_7506);
nor U14704 (N_14704,N_8359,N_11414);
and U14705 (N_14705,N_11537,N_11127);
nand U14706 (N_14706,N_12271,N_11366);
nor U14707 (N_14707,N_10276,N_7102);
xnor U14708 (N_14708,N_7945,N_12354);
nand U14709 (N_14709,N_11204,N_11357);
nor U14710 (N_14710,N_10522,N_9909);
nand U14711 (N_14711,N_10465,N_11727);
or U14712 (N_14712,N_6386,N_8475);
xnor U14713 (N_14713,N_10629,N_6893);
xor U14714 (N_14714,N_12153,N_9479);
xnor U14715 (N_14715,N_12358,N_6577);
and U14716 (N_14716,N_9306,N_6946);
nand U14717 (N_14717,N_8723,N_7438);
nor U14718 (N_14718,N_9723,N_11393);
or U14719 (N_14719,N_10296,N_11846);
nand U14720 (N_14720,N_10308,N_10600);
nor U14721 (N_14721,N_10820,N_7970);
nand U14722 (N_14722,N_12242,N_7915);
nand U14723 (N_14723,N_11346,N_8054);
and U14724 (N_14724,N_10564,N_12257);
nand U14725 (N_14725,N_7505,N_10615);
xnor U14726 (N_14726,N_10475,N_8392);
or U14727 (N_14727,N_8176,N_11495);
xnor U14728 (N_14728,N_7168,N_7835);
and U14729 (N_14729,N_9685,N_12382);
or U14730 (N_14730,N_8209,N_11877);
nor U14731 (N_14731,N_8121,N_10931);
xnor U14732 (N_14732,N_11120,N_7854);
nor U14733 (N_14733,N_7957,N_9779);
and U14734 (N_14734,N_11145,N_8761);
nand U14735 (N_14735,N_6752,N_7693);
nand U14736 (N_14736,N_6258,N_10712);
nand U14737 (N_14737,N_6396,N_6830);
or U14738 (N_14738,N_6868,N_10526);
nand U14739 (N_14739,N_7408,N_11181);
nor U14740 (N_14740,N_6394,N_8985);
xor U14741 (N_14741,N_11075,N_11793);
xnor U14742 (N_14742,N_7203,N_9108);
nand U14743 (N_14743,N_12132,N_7498);
or U14744 (N_14744,N_11233,N_6790);
nand U14745 (N_14745,N_9142,N_11073);
or U14746 (N_14746,N_9169,N_10137);
and U14747 (N_14747,N_9130,N_9443);
nand U14748 (N_14748,N_12255,N_8178);
and U14749 (N_14749,N_10159,N_8053);
xnor U14750 (N_14750,N_11251,N_9329);
nand U14751 (N_14751,N_7759,N_10260);
nand U14752 (N_14752,N_10969,N_9625);
xnor U14753 (N_14753,N_11800,N_7709);
and U14754 (N_14754,N_11006,N_12186);
nor U14755 (N_14755,N_11132,N_6494);
or U14756 (N_14756,N_11490,N_8527);
nor U14757 (N_14757,N_10599,N_10433);
xnor U14758 (N_14758,N_6815,N_8398);
and U14759 (N_14759,N_12449,N_10018);
and U14760 (N_14760,N_10520,N_8075);
xor U14761 (N_14761,N_10581,N_6902);
or U14762 (N_14762,N_7828,N_6429);
and U14763 (N_14763,N_12391,N_7803);
xor U14764 (N_14764,N_7058,N_6413);
and U14765 (N_14765,N_12209,N_6659);
nor U14766 (N_14766,N_7850,N_7818);
or U14767 (N_14767,N_7872,N_6826);
nor U14768 (N_14768,N_8655,N_9593);
xnor U14769 (N_14769,N_7877,N_6989);
xnor U14770 (N_14770,N_7332,N_7156);
nand U14771 (N_14771,N_11720,N_8515);
or U14772 (N_14772,N_9404,N_7123);
xnor U14773 (N_14773,N_10052,N_11023);
nand U14774 (N_14774,N_8256,N_11608);
nor U14775 (N_14775,N_6580,N_11037);
xnor U14776 (N_14776,N_8847,N_6823);
nand U14777 (N_14777,N_7580,N_7316);
xor U14778 (N_14778,N_11397,N_10890);
nor U14779 (N_14779,N_11101,N_8637);
or U14780 (N_14780,N_10694,N_12118);
nor U14781 (N_14781,N_6552,N_10077);
nor U14782 (N_14782,N_12177,N_7008);
or U14783 (N_14783,N_6462,N_11875);
or U14784 (N_14784,N_12243,N_8215);
xor U14785 (N_14785,N_10852,N_7875);
nand U14786 (N_14786,N_10857,N_8287);
and U14787 (N_14787,N_9240,N_9248);
nor U14788 (N_14788,N_9194,N_11508);
and U14789 (N_14789,N_7012,N_6785);
or U14790 (N_14790,N_11667,N_8538);
or U14791 (N_14791,N_11339,N_8583);
or U14792 (N_14792,N_7294,N_10221);
nand U14793 (N_14793,N_10706,N_10202);
xnor U14794 (N_14794,N_11263,N_9651);
nand U14795 (N_14795,N_10869,N_6839);
and U14796 (N_14796,N_9743,N_6733);
xor U14797 (N_14797,N_7767,N_11482);
nor U14798 (N_14798,N_7049,N_12200);
nand U14799 (N_14799,N_7605,N_11334);
nor U14800 (N_14800,N_6266,N_11531);
nand U14801 (N_14801,N_6793,N_11676);
nand U14802 (N_14802,N_8640,N_11546);
nand U14803 (N_14803,N_9361,N_7278);
xor U14804 (N_14804,N_12380,N_6858);
xor U14805 (N_14805,N_8754,N_11330);
nand U14806 (N_14806,N_11424,N_7702);
xnor U14807 (N_14807,N_11016,N_10972);
or U14808 (N_14808,N_8733,N_11696);
nor U14809 (N_14809,N_8552,N_7393);
xnor U14810 (N_14810,N_12142,N_12058);
xor U14811 (N_14811,N_10409,N_8335);
nor U14812 (N_14812,N_9189,N_8405);
nor U14813 (N_14813,N_6254,N_7779);
nor U14814 (N_14814,N_9232,N_10268);
and U14815 (N_14815,N_7209,N_12038);
xor U14816 (N_14816,N_9276,N_9263);
xnor U14817 (N_14817,N_11178,N_9934);
or U14818 (N_14818,N_9580,N_11812);
or U14819 (N_14819,N_10075,N_12092);
or U14820 (N_14820,N_7551,N_9794);
or U14821 (N_14821,N_10104,N_6654);
or U14822 (N_14822,N_7339,N_6840);
nand U14823 (N_14823,N_7687,N_10374);
nor U14824 (N_14824,N_8297,N_6445);
and U14825 (N_14825,N_8801,N_7544);
nor U14826 (N_14826,N_7516,N_10991);
nor U14827 (N_14827,N_8622,N_9757);
and U14828 (N_14828,N_8777,N_7109);
nand U14829 (N_14829,N_10646,N_9560);
and U14830 (N_14830,N_11617,N_6618);
or U14831 (N_14831,N_6722,N_12069);
xor U14832 (N_14832,N_8911,N_12202);
and U14833 (N_14833,N_8680,N_10074);
nor U14834 (N_14834,N_7884,N_9708);
xor U14835 (N_14835,N_9960,N_7267);
or U14836 (N_14836,N_8134,N_10108);
nand U14837 (N_14837,N_9932,N_8170);
xor U14838 (N_14838,N_9521,N_6374);
nor U14839 (N_14839,N_11977,N_8812);
nor U14840 (N_14840,N_7696,N_6700);
nand U14841 (N_14841,N_7615,N_7296);
or U14842 (N_14842,N_12172,N_9684);
xor U14843 (N_14843,N_12087,N_8849);
and U14844 (N_14844,N_12445,N_11313);
or U14845 (N_14845,N_7250,N_8610);
or U14846 (N_14846,N_8044,N_11867);
nand U14847 (N_14847,N_6358,N_7251);
or U14848 (N_14848,N_6928,N_7815);
xnor U14849 (N_14849,N_8677,N_9124);
and U14850 (N_14850,N_7372,N_11017);
nand U14851 (N_14851,N_8676,N_10656);
nor U14852 (N_14852,N_9624,N_9314);
or U14853 (N_14853,N_6922,N_9730);
nor U14854 (N_14854,N_11234,N_8674);
or U14855 (N_14855,N_10808,N_6298);
xnor U14856 (N_14856,N_9605,N_11310);
or U14857 (N_14857,N_10459,N_10073);
and U14858 (N_14858,N_10838,N_7333);
or U14859 (N_14859,N_6948,N_7738);
and U14860 (N_14860,N_7048,N_10617);
or U14861 (N_14861,N_8484,N_7031);
or U14862 (N_14862,N_11540,N_7512);
or U14863 (N_14863,N_7732,N_6877);
xnor U14864 (N_14864,N_12012,N_11496);
nand U14865 (N_14865,N_6609,N_10964);
xor U14866 (N_14866,N_9915,N_11956);
or U14867 (N_14867,N_6716,N_9025);
and U14868 (N_14868,N_8626,N_6500);
or U14869 (N_14869,N_8741,N_10793);
nor U14870 (N_14870,N_9258,N_6705);
nor U14871 (N_14871,N_11984,N_10301);
nand U14872 (N_14872,N_10720,N_12327);
nor U14873 (N_14873,N_8517,N_9352);
xor U14874 (N_14874,N_9529,N_9991);
or U14875 (N_14875,N_10821,N_8535);
xnor U14876 (N_14876,N_12169,N_7570);
nor U14877 (N_14877,N_9027,N_10051);
nand U14878 (N_14878,N_8943,N_8862);
nand U14879 (N_14879,N_11505,N_9430);
nand U14880 (N_14880,N_11682,N_9095);
nor U14881 (N_14881,N_8866,N_7762);
or U14882 (N_14882,N_7345,N_9394);
xnor U14883 (N_14883,N_6993,N_10277);
nand U14884 (N_14884,N_8055,N_11258);
nand U14885 (N_14885,N_10262,N_9761);
xor U14886 (N_14886,N_8184,N_8119);
or U14887 (N_14887,N_10141,N_8452);
and U14888 (N_14888,N_10479,N_9937);
or U14889 (N_14889,N_12074,N_6522);
and U14890 (N_14890,N_7999,N_6649);
nor U14891 (N_14891,N_8058,N_11272);
or U14892 (N_14892,N_6751,N_6784);
nor U14893 (N_14893,N_8089,N_7958);
and U14894 (N_14894,N_7463,N_11500);
xnor U14895 (N_14895,N_12411,N_9157);
nor U14896 (N_14896,N_7820,N_10224);
nor U14897 (N_14897,N_6341,N_6348);
nor U14898 (N_14898,N_9741,N_11942);
and U14899 (N_14899,N_11240,N_11904);
nand U14900 (N_14900,N_12328,N_12459);
xnor U14901 (N_14901,N_10407,N_6934);
nand U14902 (N_14902,N_11081,N_6871);
and U14903 (N_14903,N_8858,N_7821);
or U14904 (N_14904,N_12037,N_8854);
nor U14905 (N_14905,N_8289,N_8973);
nor U14906 (N_14906,N_6995,N_11828);
and U14907 (N_14907,N_10846,N_11317);
nand U14908 (N_14908,N_6837,N_8554);
xnor U14909 (N_14909,N_8579,N_8368);
nand U14910 (N_14910,N_7940,N_6553);
and U14911 (N_14911,N_10227,N_7843);
nor U14912 (N_14912,N_6822,N_11765);
nor U14913 (N_14913,N_7433,N_10005);
xor U14914 (N_14914,N_8432,N_10942);
nand U14915 (N_14915,N_11156,N_12494);
and U14916 (N_14916,N_9532,N_9700);
nor U14917 (N_14917,N_8994,N_10543);
nand U14918 (N_14918,N_7235,N_7422);
or U14919 (N_14919,N_7700,N_7206);
nor U14920 (N_14920,N_8035,N_7911);
nand U14921 (N_14921,N_10143,N_9072);
nor U14922 (N_14922,N_7441,N_9052);
nand U14923 (N_14923,N_8667,N_10035);
nand U14924 (N_14924,N_11372,N_8842);
nor U14925 (N_14925,N_7596,N_12491);
nor U14926 (N_14926,N_8660,N_9213);
nor U14927 (N_14927,N_11619,N_11464);
or U14928 (N_14928,N_8378,N_8941);
or U14929 (N_14929,N_8344,N_7427);
nand U14930 (N_14930,N_8786,N_9409);
xnor U14931 (N_14931,N_11377,N_7579);
xnor U14932 (N_14932,N_8800,N_7660);
xor U14933 (N_14933,N_7916,N_7486);
xnor U14934 (N_14934,N_12348,N_12402);
and U14935 (N_14935,N_9566,N_8010);
xor U14936 (N_14936,N_7919,N_9151);
xnor U14937 (N_14937,N_10850,N_9556);
or U14938 (N_14938,N_8356,N_10589);
xor U14939 (N_14939,N_9672,N_11223);
and U14940 (N_14940,N_9706,N_9609);
nor U14941 (N_14941,N_11981,N_6545);
nand U14942 (N_14942,N_9542,N_7713);
nor U14943 (N_14943,N_7324,N_9235);
or U14944 (N_14944,N_7373,N_7146);
or U14945 (N_14945,N_11912,N_7428);
xor U14946 (N_14946,N_9731,N_9036);
and U14947 (N_14947,N_8074,N_6912);
nor U14948 (N_14948,N_7417,N_8386);
or U14949 (N_14949,N_7981,N_11629);
or U14950 (N_14950,N_7106,N_9156);
nand U14951 (N_14951,N_10161,N_9077);
and U14952 (N_14952,N_6679,N_7010);
nand U14953 (N_14953,N_7774,N_12057);
xnor U14954 (N_14954,N_12194,N_7844);
nor U14955 (N_14955,N_6579,N_9445);
nor U14956 (N_14956,N_9311,N_9856);
nor U14957 (N_14957,N_11746,N_7701);
or U14958 (N_14958,N_6653,N_10147);
xor U14959 (N_14959,N_9739,N_6763);
nor U14960 (N_14960,N_6527,N_6354);
xnor U14961 (N_14961,N_9640,N_7590);
nor U14962 (N_14962,N_12313,N_8436);
nand U14963 (N_14963,N_7892,N_9223);
nand U14964 (N_14964,N_7547,N_12204);
nor U14965 (N_14965,N_10912,N_7014);
or U14966 (N_14966,N_9004,N_7040);
or U14967 (N_14967,N_7223,N_11929);
nand U14968 (N_14968,N_11406,N_9402);
nor U14969 (N_14969,N_9138,N_12323);
and U14970 (N_14970,N_9602,N_7536);
and U14971 (N_14971,N_7073,N_8028);
nor U14972 (N_14972,N_10243,N_6938);
nor U14973 (N_14973,N_7741,N_12134);
or U14974 (N_14974,N_10614,N_10422);
and U14975 (N_14975,N_6916,N_8205);
nor U14976 (N_14976,N_6410,N_9078);
xor U14977 (N_14977,N_11130,N_10343);
nor U14978 (N_14978,N_10875,N_9196);
or U14979 (N_14979,N_7188,N_7044);
or U14980 (N_14980,N_9475,N_10201);
nand U14981 (N_14981,N_9417,N_8004);
nand U14982 (N_14982,N_9017,N_7447);
xor U14983 (N_14983,N_11784,N_11615);
nor U14984 (N_14984,N_8534,N_10032);
and U14985 (N_14985,N_7965,N_7894);
xnor U14986 (N_14986,N_7518,N_11452);
and U14987 (N_14987,N_6518,N_12010);
and U14988 (N_14988,N_8163,N_7912);
nor U14989 (N_14989,N_6981,N_10856);
and U14990 (N_14990,N_10818,N_7092);
and U14991 (N_14991,N_9330,N_10805);
and U14992 (N_14992,N_12281,N_8041);
nor U14993 (N_14993,N_9211,N_11095);
nand U14994 (N_14994,N_9234,N_10881);
or U14995 (N_14995,N_6452,N_10734);
and U14996 (N_14996,N_11477,N_9238);
or U14997 (N_14997,N_10076,N_7823);
nand U14998 (N_14998,N_9617,N_10225);
or U14999 (N_14999,N_10471,N_12196);
nor U15000 (N_15000,N_8248,N_11277);
nor U15001 (N_15001,N_7376,N_10737);
or U15002 (N_15002,N_7258,N_10752);
xor U15003 (N_15003,N_8691,N_9604);
xnor U15004 (N_15004,N_11144,N_8103);
or U15005 (N_15005,N_8318,N_9200);
xor U15006 (N_15006,N_7566,N_8896);
nand U15007 (N_15007,N_9463,N_8157);
xnor U15008 (N_15008,N_8649,N_9925);
nand U15009 (N_15009,N_8991,N_10056);
xor U15010 (N_15010,N_12335,N_9993);
nor U15011 (N_15011,N_7178,N_11664);
xor U15012 (N_15012,N_8181,N_12398);
or U15013 (N_15013,N_9860,N_11616);
nand U15014 (N_15014,N_9487,N_8794);
or U15015 (N_15015,N_6568,N_11287);
xnor U15016 (N_15016,N_9303,N_9571);
xnor U15017 (N_15017,N_6695,N_10810);
nor U15018 (N_15018,N_11891,N_9195);
nor U15019 (N_15019,N_7737,N_7216);
or U15020 (N_15020,N_11421,N_9905);
nand U15021 (N_15021,N_11077,N_6980);
xnor U15022 (N_15022,N_11154,N_6930);
nor U15023 (N_15023,N_10765,N_10768);
or U15024 (N_15024,N_10468,N_8342);
and U15025 (N_15025,N_11700,N_9465);
nand U15026 (N_15026,N_6482,N_8685);
nand U15027 (N_15027,N_8220,N_10538);
nand U15028 (N_15028,N_12468,N_10948);
xnor U15029 (N_15029,N_10800,N_8032);
and U15030 (N_15030,N_7836,N_11417);
or U15031 (N_15031,N_9438,N_7224);
nor U15032 (N_15032,N_7122,N_10453);
or U15033 (N_15033,N_8254,N_6538);
xnor U15034 (N_15034,N_7057,N_9641);
nand U15035 (N_15035,N_9366,N_10930);
and U15036 (N_15036,N_8998,N_10745);
and U15037 (N_15037,N_9552,N_7069);
and U15038 (N_15038,N_7214,N_9412);
and U15039 (N_15039,N_9431,N_9039);
or U15040 (N_15040,N_8893,N_9126);
and U15041 (N_15041,N_7045,N_12056);
or U15042 (N_15042,N_12290,N_8666);
and U15043 (N_15043,N_10089,N_12340);
xnor U15044 (N_15044,N_11491,N_7555);
and U15045 (N_15045,N_6730,N_8219);
xnor U15046 (N_15046,N_10477,N_6606);
nor U15047 (N_15047,N_8855,N_8193);
and U15048 (N_15048,N_7688,N_12428);
nand U15049 (N_15049,N_6475,N_11736);
or U15050 (N_15050,N_11447,N_7113);
or U15051 (N_15051,N_11373,N_10019);
nor U15052 (N_15052,N_11962,N_8638);
or U15053 (N_15053,N_10183,N_12173);
and U15054 (N_15054,N_12108,N_11168);
and U15055 (N_15055,N_10944,N_10674);
xnor U15056 (N_15056,N_12151,N_10287);
nand U15057 (N_15057,N_10938,N_9214);
xnor U15058 (N_15058,N_11110,N_7964);
nor U15059 (N_15059,N_10924,N_8827);
xor U15060 (N_15060,N_10481,N_10923);
xnor U15061 (N_15061,N_11660,N_10612);
and U15062 (N_15062,N_9001,N_10911);
or U15063 (N_15063,N_9877,N_10338);
and U15064 (N_15064,N_9408,N_7085);
or U15065 (N_15065,N_9662,N_10235);
xnor U15066 (N_15066,N_12386,N_8345);
or U15067 (N_15067,N_8631,N_9895);
or U15068 (N_15068,N_10023,N_10244);
and U15069 (N_15069,N_12350,N_11355);
nor U15070 (N_15070,N_11960,N_8555);
or U15071 (N_15071,N_10787,N_11732);
xor U15072 (N_15072,N_10040,N_6933);
nor U15073 (N_15073,N_6505,N_12472);
and U15074 (N_15074,N_12098,N_8098);
or U15075 (N_15075,N_8995,N_10512);
and U15076 (N_15076,N_7508,N_8061);
nor U15077 (N_15077,N_12061,N_8731);
and U15078 (N_15078,N_9106,N_10380);
and U15079 (N_15079,N_8136,N_9516);
nor U15080 (N_15080,N_11610,N_11312);
or U15081 (N_15081,N_10336,N_10877);
or U15082 (N_15082,N_7988,N_8445);
nand U15083 (N_15083,N_12113,N_9298);
or U15084 (N_15084,N_12311,N_11430);
or U15085 (N_15085,N_10687,N_6762);
or U15086 (N_15086,N_11827,N_10778);
xor U15087 (N_15087,N_9155,N_6655);
xnor U15088 (N_15088,N_11801,N_9851);
nor U15089 (N_15089,N_12326,N_9220);
xor U15090 (N_15090,N_6804,N_8029);
and U15091 (N_15091,N_9097,N_6276);
and U15092 (N_15092,N_11105,N_6978);
xor U15093 (N_15093,N_9190,N_10702);
nor U15094 (N_15094,N_8867,N_8045);
nor U15095 (N_15095,N_12214,N_6282);
and U15096 (N_15096,N_7948,N_11418);
xor U15097 (N_15097,N_7374,N_7661);
nand U15098 (N_15098,N_11818,N_7275);
nand U15099 (N_15099,N_9645,N_8925);
xnor U15100 (N_15100,N_11740,N_11352);
xnor U15101 (N_15101,N_8473,N_11290);
or U15102 (N_15102,N_6513,N_11399);
nor U15103 (N_15103,N_12184,N_11729);
nand U15104 (N_15104,N_8509,N_10463);
or U15105 (N_15105,N_12418,N_12464);
xnor U15106 (N_15106,N_9839,N_12110);
or U15107 (N_15107,N_11245,N_6295);
nand U15108 (N_15108,N_12316,N_8255);
or U15109 (N_15109,N_8018,N_7624);
or U15110 (N_15110,N_9742,N_11126);
nor U15111 (N_15111,N_7432,N_11886);
nand U15112 (N_15112,N_11925,N_11327);
xnor U15113 (N_15113,N_11072,N_6465);
and U15114 (N_15114,N_11213,N_10249);
or U15115 (N_15115,N_12099,N_7987);
nor U15116 (N_15116,N_10516,N_12024);
xnor U15117 (N_15117,N_7969,N_8521);
xnor U15118 (N_15118,N_6641,N_8565);
xnor U15119 (N_15119,N_11543,N_11565);
xnor U15120 (N_15120,N_11360,N_10359);
and U15121 (N_15121,N_8506,N_12217);
and U15122 (N_15122,N_8329,N_8290);
or U15123 (N_15123,N_11633,N_7829);
nor U15124 (N_15124,N_7833,N_10452);
nand U15125 (N_15125,N_7182,N_12288);
or U15126 (N_15126,N_6620,N_9485);
nor U15127 (N_15127,N_11591,N_12144);
nor U15128 (N_15128,N_12016,N_8945);
xnor U15129 (N_15129,N_11432,N_11008);
nand U15130 (N_15130,N_10153,N_8960);
xnor U15131 (N_15131,N_8472,N_8467);
or U15132 (N_15132,N_7200,N_7625);
nand U15133 (N_15133,N_7334,N_6373);
or U15134 (N_15134,N_8351,N_7949);
and U15135 (N_15135,N_8774,N_8601);
nand U15136 (N_15136,N_10344,N_7927);
xor U15137 (N_15137,N_11752,N_11128);
and U15138 (N_15138,N_6712,N_7860);
nor U15139 (N_15139,N_11806,N_7593);
xnor U15140 (N_15140,N_7384,N_11400);
nor U15141 (N_15141,N_11782,N_7434);
xnor U15142 (N_15142,N_9024,N_8548);
xnor U15143 (N_15143,N_9437,N_7253);
or U15144 (N_15144,N_10297,N_10484);
xor U15145 (N_15145,N_11970,N_11697);
nor U15146 (N_15146,N_12149,N_7904);
nand U15147 (N_15147,N_10386,N_7164);
nor U15148 (N_15148,N_8837,N_11255);
or U15149 (N_15149,N_10624,N_8856);
nand U15150 (N_15150,N_12431,N_9551);
xor U15151 (N_15151,N_7740,N_9807);
and U15152 (N_15152,N_8739,N_7271);
and U15153 (N_15153,N_11318,N_12158);
and U15154 (N_15154,N_10034,N_11293);
or U15155 (N_15155,N_8260,N_9429);
nand U15156 (N_15156,N_9793,N_11504);
and U15157 (N_15157,N_8461,N_11208);
nand U15158 (N_15158,N_8752,N_10130);
and U15159 (N_15159,N_6825,N_6352);
and U15160 (N_15160,N_9999,N_6346);
and U15161 (N_15161,N_11931,N_7142);
and U15162 (N_15162,N_9727,N_7027);
nor U15163 (N_15163,N_10101,N_7330);
nor U15164 (N_15164,N_11783,N_10827);
and U15165 (N_15165,N_12419,N_10234);
xnor U15166 (N_15166,N_6347,N_8148);
nor U15167 (N_15167,N_7466,N_11423);
or U15168 (N_15168,N_8732,N_11100);
and U15169 (N_15169,N_11440,N_8696);
xor U15170 (N_15170,N_7841,N_10041);
xnor U15171 (N_15171,N_9943,N_11798);
or U15172 (N_15172,N_10028,N_10760);
and U15173 (N_15173,N_10979,N_11069);
or U15174 (N_15174,N_7088,N_8025);
and U15175 (N_15175,N_11358,N_8907);
xor U15176 (N_15176,N_8470,N_11087);
nor U15177 (N_15177,N_9959,N_11438);
or U15178 (N_15178,N_7252,N_6591);
nand U15179 (N_15179,N_8174,N_7367);
and U15180 (N_15180,N_6852,N_8308);
and U15181 (N_15181,N_7231,N_10483);
xor U15182 (N_15182,N_8479,N_6630);
and U15183 (N_15183,N_7095,N_6627);
or U15184 (N_15184,N_9607,N_11640);
xnor U15185 (N_15185,N_9413,N_8578);
xor U15186 (N_15186,N_12041,N_8224);
or U15187 (N_15187,N_10823,N_10576);
xnor U15188 (N_15188,N_8544,N_10211);
xnor U15189 (N_15189,N_7847,N_9780);
xnor U15190 (N_15190,N_9848,N_11173);
or U15191 (N_15191,N_8549,N_6262);
nand U15192 (N_15192,N_9555,N_9530);
or U15193 (N_15193,N_8015,N_10205);
nand U15194 (N_15194,N_7000,N_12339);
nand U15195 (N_15195,N_11239,N_7368);
and U15196 (N_15196,N_9279,N_10231);
and U15197 (N_15197,N_9528,N_8821);
nor U15198 (N_15198,N_7733,N_8480);
nand U15199 (N_15199,N_6920,N_10519);
and U15200 (N_15200,N_9892,N_9548);
nand U15201 (N_15201,N_8397,N_7751);
nor U15202 (N_15202,N_7183,N_8904);
nor U15203 (N_15203,N_6325,N_8246);
or U15204 (N_15204,N_8019,N_10203);
or U15205 (N_15205,N_8541,N_8214);
nor U15206 (N_15206,N_11570,N_11808);
and U15207 (N_15207,N_10182,N_7559);
or U15208 (N_15208,N_8672,N_10762);
nand U15209 (N_15209,N_8369,N_8311);
nand U15210 (N_15210,N_7121,N_8591);
and U15211 (N_15211,N_7461,N_11065);
or U15212 (N_15212,N_12141,N_8488);
nor U15213 (N_15213,N_8716,N_10916);
xnor U15214 (N_15214,N_12277,N_9243);
and U15215 (N_15215,N_11143,N_8026);
nand U15216 (N_15216,N_6585,N_11336);
and U15217 (N_15217,N_7479,N_11552);
nand U15218 (N_15218,N_8151,N_11802);
or U15219 (N_15219,N_10332,N_8444);
nor U15220 (N_15220,N_9497,N_8050);
and U15221 (N_15221,N_10795,N_7274);
or U15222 (N_15222,N_6412,N_7353);
and U15223 (N_15223,N_7337,N_7237);
xor U15224 (N_15224,N_8642,N_12426);
nor U15225 (N_15225,N_9137,N_9259);
nand U15226 (N_15226,N_10196,N_12030);
and U15227 (N_15227,N_10418,N_7897);
or U15228 (N_15228,N_12362,N_11305);
or U15229 (N_15229,N_7923,N_6336);
nor U15230 (N_15230,N_7476,N_8361);
and U15231 (N_15231,N_8112,N_7234);
nor U15232 (N_15232,N_11982,N_11524);
and U15233 (N_15233,N_6688,N_10759);
nor U15234 (N_15234,N_9590,N_12093);
nand U15235 (N_15235,N_8750,N_7270);
xnor U15236 (N_15236,N_12284,N_11434);
nand U15237 (N_15237,N_6470,N_7866);
nor U15238 (N_15238,N_11222,N_8237);
xnor U15239 (N_15239,N_10887,N_6573);
xor U15240 (N_15240,N_7181,N_11365);
nor U15241 (N_15241,N_8073,N_10346);
nor U15242 (N_15242,N_10065,N_9669);
and U15243 (N_15243,N_12221,N_6662);
and U15244 (N_15244,N_11271,N_8095);
nor U15245 (N_15245,N_10622,N_8708);
and U15246 (N_15246,N_7971,N_10722);
nand U15247 (N_15247,N_10771,N_9028);
and U15248 (N_15248,N_12188,N_12193);
or U15249 (N_15249,N_9099,N_10551);
nor U15250 (N_15250,N_9403,N_11926);
nand U15251 (N_15251,N_8744,N_7645);
nand U15252 (N_15252,N_6340,N_7152);
xor U15253 (N_15253,N_9216,N_10449);
nand U15254 (N_15254,N_7423,N_9346);
and U15255 (N_15255,N_9597,N_6339);
nor U15256 (N_15256,N_11361,N_11135);
nor U15257 (N_15257,N_10237,N_7510);
and U15258 (N_15258,N_9695,N_12161);
nand U15259 (N_15259,N_7282,N_6795);
nor U15260 (N_15260,N_7460,N_10552);
or U15261 (N_15261,N_11693,N_7063);
xor U15262 (N_15262,N_9081,N_11838);
and U15263 (N_15263,N_10191,N_6319);
or U15264 (N_15264,N_11730,N_7273);
nand U15265 (N_15265,N_6471,N_9419);
xnor U15266 (N_15266,N_6907,N_10337);
and U15267 (N_15267,N_10876,N_9753);
xor U15268 (N_15268,N_11885,N_8996);
and U15269 (N_15269,N_11921,N_7140);
xor U15270 (N_15270,N_9227,N_10932);
and U15271 (N_15271,N_8207,N_7611);
and U15272 (N_15272,N_12106,N_6952);
xor U15273 (N_15273,N_9912,N_8406);
nor U15274 (N_15274,N_9584,N_11906);
nand U15275 (N_15275,N_11945,N_11857);
nor U15276 (N_15276,N_8967,N_9061);
and U15277 (N_15277,N_10105,N_9059);
xor U15278 (N_15278,N_12066,N_10699);
and U15279 (N_15279,N_6279,N_10457);
nand U15280 (N_15280,N_10066,N_9704);
and U15281 (N_15281,N_12482,N_8159);
xor U15282 (N_15282,N_9031,N_12088);
xnor U15283 (N_15283,N_9362,N_7015);
nand U15284 (N_15284,N_10858,N_11995);
xnor U15285 (N_15285,N_8875,N_10057);
nor U15286 (N_15286,N_12211,N_7633);
nand U15287 (N_15287,N_12020,N_11000);
nor U15288 (N_15288,N_6598,N_10515);
nor U15289 (N_15289,N_7692,N_9318);
xnor U15290 (N_15290,N_7626,N_6411);
xor U15291 (N_15291,N_11052,N_12366);
nor U15292 (N_15292,N_10311,N_6713);
xnor U15293 (N_15293,N_9353,N_10250);
and U15294 (N_15294,N_7745,N_7763);
nand U15295 (N_15295,N_11429,N_11584);
xor U15296 (N_15296,N_7691,N_8958);
xnor U15297 (N_15297,N_10081,N_12286);
and U15298 (N_15298,N_12338,N_12007);
or U15299 (N_15299,N_10298,N_9967);
nor U15300 (N_15300,N_7171,N_7621);
nor U15301 (N_15301,N_11713,N_7802);
nor U15302 (N_15302,N_9334,N_6789);
nand U15303 (N_15303,N_6707,N_11772);
and U15304 (N_15304,N_8747,N_9177);
xor U15305 (N_15305,N_10323,N_12297);
xor U15306 (N_15306,N_7834,N_7725);
or U15307 (N_15307,N_11609,N_6835);
nand U15308 (N_15308,N_8272,N_7482);
or U15309 (N_15309,N_7210,N_10317);
xor U15310 (N_15310,N_9827,N_6838);
or U15311 (N_15311,N_11599,N_12387);
nand U15312 (N_15312,N_10873,N_9808);
nand U15313 (N_15313,N_7666,N_6593);
or U15314 (N_15314,N_11575,N_10956);
and U15315 (N_15315,N_9035,N_11383);
nor U15316 (N_15316,N_11155,N_8594);
xnor U15317 (N_15317,N_12253,N_6919);
nor U15318 (N_15318,N_8187,N_11413);
nor U15319 (N_15319,N_10532,N_12222);
or U15320 (N_15320,N_12299,N_8576);
nand U15321 (N_15321,N_12458,N_11471);
nand U15322 (N_15322,N_9315,N_8656);
and U15323 (N_15323,N_11632,N_10036);
nor U15324 (N_15324,N_8217,N_7059);
and U15325 (N_15325,N_6693,N_9380);
or U15326 (N_15326,N_10427,N_11770);
xor U15327 (N_15327,N_6351,N_11219);
or U15328 (N_15328,N_11253,N_12029);
nor U15329 (N_15329,N_11996,N_8443);
and U15330 (N_15330,N_9505,N_6941);
nand U15331 (N_15331,N_11836,N_8700);
xor U15332 (N_15332,N_9153,N_11298);
or U15333 (N_15333,N_10695,N_8635);
or U15334 (N_15334,N_11516,N_8384);
and U15335 (N_15335,N_8064,N_11387);
nand U15336 (N_15336,N_11919,N_10370);
nand U15337 (N_15337,N_6668,N_6670);
or U15338 (N_15338,N_7659,N_10318);
xnor U15339 (N_15339,N_12407,N_6843);
and U15340 (N_15340,N_10266,N_6498);
xor U15341 (N_15341,N_9030,N_7607);
nand U15342 (N_15342,N_8315,N_10478);
or U15343 (N_15343,N_11456,N_7340);
xnor U15344 (N_15344,N_11359,N_9531);
and U15345 (N_15345,N_9224,N_6645);
xor U15346 (N_15346,N_7899,N_6383);
and U15347 (N_15347,N_7042,N_10355);
or U15348 (N_15348,N_9480,N_9919);
xnor U15349 (N_15349,N_8861,N_9295);
nand U15350 (N_15350,N_10412,N_11200);
or U15351 (N_15351,N_9356,N_8940);
and U15352 (N_15352,N_7056,N_8139);
xnor U15353 (N_15353,N_10322,N_9171);
nand U15354 (N_15354,N_7513,N_9476);
nor U15355 (N_15355,N_6747,N_10807);
xnor U15356 (N_15356,N_11545,N_8152);
xor U15357 (N_15357,N_7950,N_12019);
nand U15358 (N_15358,N_12377,N_9812);
xor U15359 (N_15359,N_10660,N_7728);
and U15360 (N_15360,N_10321,N_7710);
xnor U15361 (N_15361,N_6629,N_12224);
and U15362 (N_15362,N_10736,N_9520);
xnor U15363 (N_15363,N_8067,N_7972);
and U15364 (N_15364,N_10578,N_7655);
nand U15365 (N_15365,N_6820,N_11529);
or U15366 (N_15366,N_6478,N_8778);
nor U15367 (N_15367,N_8066,N_8258);
nor U15368 (N_15368,N_11019,N_9850);
or U15369 (N_15369,N_9209,N_7150);
nor U15370 (N_15370,N_6692,N_11345);
nor U15371 (N_15371,N_10993,N_9494);
nor U15372 (N_15372,N_7703,N_10345);
nor U15373 (N_15373,N_9766,N_6441);
or U15374 (N_15374,N_10088,N_6499);
and U15375 (N_15375,N_12487,N_10010);
xor U15376 (N_15376,N_8080,N_9129);
or U15377 (N_15377,N_8383,N_12446);
nor U15378 (N_15378,N_6597,N_8980);
xor U15379 (N_15379,N_7366,N_8828);
nand U15380 (N_15380,N_8155,N_11955);
or U15381 (N_15381,N_6901,N_8883);
nand U15382 (N_15382,N_9320,N_12115);
and U15383 (N_15383,N_7019,N_7873);
or U15384 (N_15384,N_10474,N_12373);
or U15385 (N_15385,N_7718,N_7735);
nor U15386 (N_15386,N_8115,N_7119);
nor U15387 (N_15387,N_6776,N_8609);
or U15388 (N_15388,N_7133,N_9966);
or U15389 (N_15389,N_6557,N_6832);
xor U15390 (N_15390,N_10180,N_6834);
xor U15391 (N_15391,N_9771,N_12395);
xnor U15392 (N_15392,N_9927,N_8665);
xor U15393 (N_15393,N_12060,N_8791);
or U15394 (N_15394,N_6576,N_12314);
xor U15395 (N_15395,N_7863,N_12232);
nand U15396 (N_15396,N_8639,N_9680);
and U15397 (N_15397,N_11767,N_11939);
nand U15398 (N_15398,N_7561,N_12415);
xor U15399 (N_15399,N_9841,N_7572);
and U15400 (N_15400,N_8185,N_6644);
and U15401 (N_15401,N_12252,N_6886);
nor U15402 (N_15402,N_9975,N_11026);
xnor U15403 (N_15403,N_12121,N_8367);
nand U15404 (N_15404,N_8084,N_11488);
and U15405 (N_15405,N_8312,N_9079);
nor U15406 (N_15406,N_10219,N_11404);
and U15407 (N_15407,N_9682,N_9751);
or U15408 (N_15408,N_10605,N_10819);
nand U15409 (N_15409,N_6767,N_6414);
or U15410 (N_15410,N_10176,N_10261);
and U15411 (N_15411,N_8788,N_10278);
nand U15412 (N_15412,N_7467,N_7453);
nor U15413 (N_15413,N_8400,N_8451);
xor U15414 (N_15414,N_10527,N_11304);
nor U15415 (N_15415,N_6277,N_9456);
xor U15416 (N_15416,N_11908,N_11499);
nor U15417 (N_15417,N_9010,N_8859);
nand U15418 (N_15418,N_10114,N_10713);
nand U15419 (N_15419,N_8605,N_7840);
and U15420 (N_15420,N_11123,N_9785);
nor U15421 (N_15421,N_7180,N_11907);
and U15422 (N_15422,N_11206,N_11966);
or U15423 (N_15423,N_10597,N_8465);
nor U15424 (N_15424,N_7556,N_12105);
or U15425 (N_15425,N_10659,N_8179);
or U15426 (N_15426,N_10091,N_11182);
and U15427 (N_15427,N_11781,N_8213);
nand U15428 (N_15428,N_8123,N_10320);
nor U15429 (N_15429,N_9965,N_11249);
xor U15430 (N_15430,N_8453,N_12086);
nor U15431 (N_15431,N_7487,N_6448);
nor U15432 (N_15432,N_8726,N_7651);
xor U15433 (N_15433,N_9119,N_9961);
or U15434 (N_15434,N_11354,N_9091);
xor U15435 (N_15435,N_10517,N_7929);
nor U15436 (N_15436,N_7046,N_6881);
nand U15437 (N_15437,N_6561,N_10193);
and U15438 (N_15438,N_6758,N_8743);
nor U15439 (N_15439,N_8198,N_12220);
xnor U15440 (N_15440,N_11382,N_11351);
nand U15441 (N_15441,N_11859,N_9385);
and U15442 (N_15442,N_9237,N_7297);
and U15443 (N_15443,N_6818,N_8653);
xnor U15444 (N_15444,N_11731,N_7177);
or U15445 (N_15445,N_11787,N_10970);
or U15446 (N_15446,N_8276,N_6275);
xnor U15447 (N_15447,N_11261,N_6848);
nand U15448 (N_15448,N_8536,N_7974);
and U15449 (N_15449,N_9393,N_8474);
and U15450 (N_15450,N_9117,N_11703);
nand U15451 (N_15451,N_10454,N_12371);
or U15452 (N_15452,N_11975,N_9917);
or U15453 (N_15453,N_9712,N_6816);
or U15454 (N_15454,N_11622,N_7694);
xor U15455 (N_15455,N_9239,N_10047);
and U15456 (N_15456,N_9963,N_6446);
or U15457 (N_15457,N_8132,N_6521);
or U15458 (N_15458,N_11091,N_12272);
nand U15459 (N_15459,N_8839,N_8459);
nor U15460 (N_15460,N_12225,N_11465);
and U15461 (N_15461,N_8257,N_11114);
or U15462 (N_15462,N_9219,N_12137);
or U15463 (N_15463,N_12414,N_10955);
nor U15464 (N_15464,N_10826,N_9715);
nand U15465 (N_15465,N_6595,N_9472);
or U15466 (N_15466,N_11675,N_12062);
nand U15467 (N_15467,N_9744,N_10839);
and U15468 (N_15468,N_10365,N_10151);
or U15469 (N_15469,N_8928,N_10230);
and U15470 (N_15470,N_10556,N_6844);
and U15471 (N_15471,N_6607,N_12437);
nor U15472 (N_15472,N_11815,N_10973);
nor U15473 (N_15473,N_8627,N_6443);
or U15474 (N_15474,N_9233,N_12000);
nand U15475 (N_15475,N_8394,N_8060);
nor U15476 (N_15476,N_8097,N_12330);
or U15477 (N_15477,N_9473,N_10724);
nor U15478 (N_15478,N_12370,N_7663);
nor U15479 (N_15479,N_12157,N_7858);
and U15480 (N_15480,N_8987,N_7629);
and U15481 (N_15481,N_6311,N_11518);
and U15482 (N_15482,N_12133,N_6739);
xnor U15483 (N_15483,N_9378,N_7392);
or U15484 (N_15484,N_9045,N_9980);
or U15485 (N_15485,N_9951,N_7429);
and U15486 (N_15486,N_8586,N_9997);
xnor U15487 (N_15487,N_9297,N_10226);
or U15488 (N_15488,N_7360,N_7304);
nand U15489 (N_15489,N_8280,N_7538);
and U15490 (N_15490,N_7558,N_11476);
nand U15491 (N_15491,N_7405,N_10420);
xor U15492 (N_15492,N_8234,N_11694);
nor U15493 (N_15493,N_11739,N_10531);
nor U15494 (N_15494,N_10689,N_7503);
nor U15495 (N_15495,N_6940,N_7769);
nand U15496 (N_15496,N_10472,N_11291);
or U15497 (N_15497,N_12266,N_9269);
or U15498 (N_15498,N_6294,N_7192);
nor U15499 (N_15499,N_8533,N_10030);
xor U15500 (N_15500,N_7309,N_11522);
and U15501 (N_15501,N_11573,N_10952);
and U15502 (N_15502,N_8130,N_9677);
nand U15503 (N_15503,N_11650,N_6290);
nor U15504 (N_15504,N_11033,N_9202);
or U15505 (N_15505,N_6889,N_7985);
xnor U15506 (N_15506,N_10542,N_11165);
and U15507 (N_15507,N_8230,N_12399);
nand U15508 (N_15508,N_10357,N_7245);
nand U15509 (N_15509,N_9774,N_6675);
xnor U15510 (N_15510,N_7201,N_10233);
nor U15511 (N_15511,N_8570,N_7975);
xnor U15512 (N_15512,N_9890,N_8303);
and U15513 (N_15513,N_9058,N_8046);
nand U15514 (N_15514,N_8913,N_12355);
nand U15515 (N_15515,N_10764,N_11744);
or U15516 (N_15516,N_10476,N_6953);
or U15517 (N_15517,N_12013,N_10862);
xnor U15518 (N_15518,N_7160,N_7195);
xnor U15519 (N_15519,N_7796,N_12344);
or U15520 (N_15520,N_6360,N_7794);
xnor U15521 (N_15521,N_9646,N_9924);
nor U15522 (N_15522,N_10566,N_8932);
nand U15523 (N_15523,N_11741,N_10677);
and U15524 (N_15524,N_9060,N_10936);
and U15525 (N_15525,N_11363,N_10588);
or U15526 (N_15526,N_9507,N_11115);
or U15527 (N_15527,N_10879,N_6748);
xor U15528 (N_15528,N_11371,N_11778);
xnor U15529 (N_15529,N_9538,N_6725);
or U15530 (N_15530,N_12176,N_7454);
nor U15531 (N_15531,N_8082,N_10399);
and U15532 (N_15532,N_6777,N_11742);
and U15533 (N_15533,N_6455,N_11177);
and U15534 (N_15534,N_7111,N_10162);
and U15535 (N_15535,N_9410,N_6393);
nand U15536 (N_15536,N_9446,N_7670);
and U15537 (N_15537,N_9957,N_10585);
nor U15538 (N_15538,N_11036,N_12420);
and U15539 (N_15539,N_8808,N_9764);
and U15540 (N_15540,N_10145,N_7669);
xor U15541 (N_15541,N_8767,N_11254);
or U15542 (N_15542,N_7785,N_10661);
nor U15543 (N_15543,N_8608,N_12393);
and U15544 (N_15544,N_10122,N_10728);
nor U15545 (N_15545,N_11819,N_11872);
and U15546 (N_15546,N_12490,N_9891);
nor U15547 (N_15547,N_12447,N_7124);
xnor U15548 (N_15548,N_7990,N_8100);
xor U15549 (N_15549,N_8428,N_7986);
and U15550 (N_15550,N_11549,N_12385);
or U15551 (N_15551,N_10987,N_6349);
xnor U15552 (N_15552,N_12233,N_6551);
or U15553 (N_15553,N_10360,N_9128);
or U15554 (N_15554,N_9996,N_11109);
nor U15555 (N_15555,N_7025,N_10377);
nand U15556 (N_15556,N_7724,N_6457);
or U15557 (N_15557,N_11876,N_6402);
or U15558 (N_15558,N_7397,N_6306);
nand U15559 (N_15559,N_8562,N_6865);
or U15560 (N_15560,N_9838,N_6900);
nand U15561 (N_15561,N_9203,N_12048);
and U15562 (N_15562,N_8076,N_8959);
and U15563 (N_15563,N_8563,N_7993);
and U15564 (N_15564,N_9983,N_9338);
or U15565 (N_15565,N_10397,N_11118);
nor U15566 (N_15566,N_8815,N_12178);
nand U15567 (N_15567,N_8611,N_12031);
nand U15568 (N_15568,N_10014,N_6434);
or U15569 (N_15569,N_12246,N_8906);
nand U15570 (N_15570,N_11896,N_7217);
and U15571 (N_15571,N_11459,N_12375);
or U15572 (N_15572,N_6833,N_10582);
nor U15573 (N_15573,N_11589,N_8684);
nor U15574 (N_15574,N_10638,N_10417);
nor U15575 (N_15575,N_10812,N_11231);
nand U15576 (N_15576,N_7657,N_7154);
nor U15577 (N_15577,N_11320,N_10424);
or U15578 (N_15578,N_10937,N_11776);
nor U15579 (N_15579,N_12140,N_9809);
nor U15580 (N_15580,N_6270,N_7215);
nand U15581 (N_15581,N_11064,N_11753);
nor U15582 (N_15582,N_7100,N_11066);
or U15583 (N_15583,N_9345,N_7549);
or U15584 (N_15584,N_11947,N_7822);
nor U15585 (N_15585,N_6850,N_11653);
nand U15586 (N_15586,N_8226,N_6754);
xnor U15587 (N_15587,N_11691,N_8567);
or U15588 (N_15588,N_7646,N_7064);
nand U15589 (N_15589,N_8446,N_6450);
nor U15590 (N_15590,N_8804,N_9837);
or U15591 (N_15591,N_10888,N_11367);
nand U15592 (N_15592,N_7400,N_8109);
xor U15593 (N_15593,N_6792,N_6849);
or U15594 (N_15594,N_11021,N_10009);
xor U15595 (N_15595,N_11613,N_8693);
or U15596 (N_15596,N_10672,N_9600);
nor U15597 (N_15597,N_9908,N_12372);
xnor U15598 (N_15598,N_11282,N_8969);
nor U15599 (N_15599,N_10245,N_7928);
xnor U15600 (N_15600,N_10275,N_6913);
nor U15601 (N_15601,N_8580,N_10149);
or U15602 (N_15602,N_8086,N_12383);
or U15603 (N_15603,N_11068,N_11963);
and U15604 (N_15604,N_9154,N_11796);
and U15605 (N_15605,N_10356,N_8588);
or U15606 (N_15606,N_11058,N_7469);
and U15607 (N_15607,N_7017,N_8841);
and U15608 (N_15608,N_10634,N_8695);
xor U15609 (N_15609,N_8371,N_7426);
or U15610 (N_15610,N_9622,N_10135);
xor U15611 (N_15611,N_9787,N_7777);
nor U15612 (N_15612,N_9916,N_8779);
or U15613 (N_15613,N_8154,N_10031);
nor U15614 (N_15614,N_11539,N_6750);
nor U15615 (N_15615,N_11040,N_7277);
nand U15616 (N_15616,N_7783,N_11813);
or U15617 (N_15617,N_6459,N_6814);
nand U15618 (N_15618,N_6392,N_9459);
xnor U15619 (N_15619,N_9549,N_10947);
xor U15620 (N_15620,N_11871,N_9979);
nand U15621 (N_15621,N_9374,N_9384);
or U15622 (N_15622,N_10401,N_10667);
nor U15623 (N_15623,N_8438,N_9798);
and U15624 (N_15624,N_10545,N_8572);
nor U15625 (N_15625,N_10861,N_7761);
xor U15626 (N_15626,N_9001,N_8000);
or U15627 (N_15627,N_7607,N_6883);
nor U15628 (N_15628,N_7390,N_7301);
and U15629 (N_15629,N_7514,N_10311);
nand U15630 (N_15630,N_12279,N_9205);
nor U15631 (N_15631,N_11693,N_11233);
nand U15632 (N_15632,N_9159,N_6570);
nor U15633 (N_15633,N_6548,N_10518);
xor U15634 (N_15634,N_7908,N_8334);
and U15635 (N_15635,N_7842,N_10659);
nand U15636 (N_15636,N_8273,N_6634);
xor U15637 (N_15637,N_9306,N_12117);
or U15638 (N_15638,N_11518,N_11549);
nor U15639 (N_15639,N_11250,N_8049);
or U15640 (N_15640,N_8622,N_10924);
xor U15641 (N_15641,N_8084,N_9500);
nor U15642 (N_15642,N_11984,N_7006);
or U15643 (N_15643,N_12421,N_11269);
and U15644 (N_15644,N_8663,N_6495);
and U15645 (N_15645,N_10727,N_9072);
xor U15646 (N_15646,N_10708,N_7011);
and U15647 (N_15647,N_10569,N_10737);
nor U15648 (N_15648,N_8540,N_6989);
xor U15649 (N_15649,N_8284,N_9421);
or U15650 (N_15650,N_10877,N_9733);
xnor U15651 (N_15651,N_8127,N_12186);
or U15652 (N_15652,N_7131,N_6860);
xnor U15653 (N_15653,N_7947,N_7710);
and U15654 (N_15654,N_7816,N_11287);
xnor U15655 (N_15655,N_12405,N_9623);
nand U15656 (N_15656,N_9329,N_8476);
or U15657 (N_15657,N_12352,N_8128);
nand U15658 (N_15658,N_8814,N_7998);
nand U15659 (N_15659,N_8156,N_9870);
nand U15660 (N_15660,N_10623,N_6619);
or U15661 (N_15661,N_12156,N_8731);
xnor U15662 (N_15662,N_10665,N_9884);
nand U15663 (N_15663,N_8120,N_9249);
and U15664 (N_15664,N_9978,N_9288);
or U15665 (N_15665,N_7260,N_6679);
or U15666 (N_15666,N_8956,N_11669);
nand U15667 (N_15667,N_11416,N_9088);
xnor U15668 (N_15668,N_11547,N_10290);
nor U15669 (N_15669,N_8387,N_11794);
and U15670 (N_15670,N_10962,N_6708);
or U15671 (N_15671,N_10112,N_11467);
and U15672 (N_15672,N_12495,N_12412);
or U15673 (N_15673,N_9347,N_11298);
and U15674 (N_15674,N_6323,N_9847);
nand U15675 (N_15675,N_9940,N_8518);
or U15676 (N_15676,N_9583,N_7577);
and U15677 (N_15677,N_12259,N_6731);
xor U15678 (N_15678,N_11864,N_12131);
nor U15679 (N_15679,N_8855,N_8531);
or U15680 (N_15680,N_7062,N_9040);
and U15681 (N_15681,N_6449,N_10803);
nor U15682 (N_15682,N_6259,N_7994);
nor U15683 (N_15683,N_7527,N_9534);
or U15684 (N_15684,N_8088,N_12459);
and U15685 (N_15685,N_10237,N_8519);
and U15686 (N_15686,N_9756,N_6326);
nor U15687 (N_15687,N_6755,N_7292);
nand U15688 (N_15688,N_11976,N_11032);
nor U15689 (N_15689,N_7891,N_7818);
xor U15690 (N_15690,N_12101,N_8855);
nor U15691 (N_15691,N_9303,N_12159);
or U15692 (N_15692,N_11941,N_8996);
or U15693 (N_15693,N_12415,N_11346);
xor U15694 (N_15694,N_6734,N_8436);
nand U15695 (N_15695,N_10434,N_10211);
and U15696 (N_15696,N_9973,N_11113);
nor U15697 (N_15697,N_9799,N_9330);
xnor U15698 (N_15698,N_10837,N_11542);
xnor U15699 (N_15699,N_11160,N_10901);
nand U15700 (N_15700,N_8507,N_6440);
or U15701 (N_15701,N_8292,N_11614);
or U15702 (N_15702,N_10022,N_8176);
xnor U15703 (N_15703,N_8618,N_9800);
or U15704 (N_15704,N_12081,N_11256);
and U15705 (N_15705,N_10308,N_8756);
nand U15706 (N_15706,N_8589,N_10483);
nor U15707 (N_15707,N_9733,N_11127);
xnor U15708 (N_15708,N_11408,N_9413);
and U15709 (N_15709,N_12344,N_9674);
nor U15710 (N_15710,N_6857,N_12331);
nor U15711 (N_15711,N_11199,N_9983);
nor U15712 (N_15712,N_9709,N_11596);
xnor U15713 (N_15713,N_8632,N_10433);
nand U15714 (N_15714,N_10609,N_6820);
or U15715 (N_15715,N_9029,N_11169);
nand U15716 (N_15716,N_11815,N_8663);
or U15717 (N_15717,N_6721,N_8721);
nand U15718 (N_15718,N_8151,N_9633);
nand U15719 (N_15719,N_7210,N_11246);
nand U15720 (N_15720,N_11149,N_8925);
nor U15721 (N_15721,N_12315,N_12206);
or U15722 (N_15722,N_9684,N_8834);
xor U15723 (N_15723,N_6622,N_10165);
nand U15724 (N_15724,N_10632,N_7198);
or U15725 (N_15725,N_9937,N_7889);
and U15726 (N_15726,N_8525,N_6577);
or U15727 (N_15727,N_6866,N_10466);
xor U15728 (N_15728,N_6304,N_11891);
and U15729 (N_15729,N_12189,N_10443);
and U15730 (N_15730,N_11066,N_10349);
nor U15731 (N_15731,N_11190,N_8533);
xnor U15732 (N_15732,N_8751,N_11801);
xor U15733 (N_15733,N_7804,N_6694);
and U15734 (N_15734,N_11877,N_8085);
nand U15735 (N_15735,N_7667,N_6600);
xor U15736 (N_15736,N_6454,N_10188);
or U15737 (N_15737,N_6514,N_7786);
or U15738 (N_15738,N_6970,N_12003);
xnor U15739 (N_15739,N_6496,N_7005);
or U15740 (N_15740,N_10724,N_8173);
nor U15741 (N_15741,N_10684,N_7784);
and U15742 (N_15742,N_11708,N_11464);
and U15743 (N_15743,N_6590,N_11633);
nand U15744 (N_15744,N_10328,N_9836);
and U15745 (N_15745,N_7006,N_6601);
nor U15746 (N_15746,N_7155,N_9292);
xor U15747 (N_15747,N_7410,N_6913);
nand U15748 (N_15748,N_7313,N_12012);
nand U15749 (N_15749,N_10670,N_10316);
nand U15750 (N_15750,N_8220,N_7389);
nor U15751 (N_15751,N_12266,N_12220);
xor U15752 (N_15752,N_12122,N_6501);
nand U15753 (N_15753,N_8908,N_11566);
or U15754 (N_15754,N_6703,N_8823);
or U15755 (N_15755,N_6961,N_7602);
nand U15756 (N_15756,N_11104,N_12484);
nor U15757 (N_15757,N_10284,N_6846);
nor U15758 (N_15758,N_9371,N_11081);
and U15759 (N_15759,N_7835,N_9763);
nor U15760 (N_15760,N_11095,N_9456);
nand U15761 (N_15761,N_8964,N_10145);
xnor U15762 (N_15762,N_9446,N_7144);
nor U15763 (N_15763,N_7785,N_9456);
or U15764 (N_15764,N_7371,N_9910);
and U15765 (N_15765,N_7113,N_7875);
or U15766 (N_15766,N_8923,N_9455);
xor U15767 (N_15767,N_9953,N_11596);
or U15768 (N_15768,N_6253,N_10620);
xnor U15769 (N_15769,N_9538,N_6943);
xnor U15770 (N_15770,N_9242,N_9865);
nor U15771 (N_15771,N_9581,N_6792);
or U15772 (N_15772,N_12273,N_6987);
and U15773 (N_15773,N_11379,N_9820);
xnor U15774 (N_15774,N_8390,N_10504);
nor U15775 (N_15775,N_8629,N_8324);
nand U15776 (N_15776,N_9108,N_10679);
or U15777 (N_15777,N_11265,N_10690);
xnor U15778 (N_15778,N_10355,N_10034);
and U15779 (N_15779,N_12283,N_12226);
nand U15780 (N_15780,N_9589,N_11039);
and U15781 (N_15781,N_8052,N_6634);
or U15782 (N_15782,N_6389,N_9959);
or U15783 (N_15783,N_11928,N_12155);
nand U15784 (N_15784,N_10969,N_6936);
nand U15785 (N_15785,N_7674,N_10890);
xnor U15786 (N_15786,N_11323,N_8381);
nor U15787 (N_15787,N_11622,N_8657);
xnor U15788 (N_15788,N_7097,N_9024);
or U15789 (N_15789,N_11688,N_12122);
or U15790 (N_15790,N_11024,N_8573);
xnor U15791 (N_15791,N_6734,N_10059);
or U15792 (N_15792,N_11581,N_11486);
xnor U15793 (N_15793,N_10536,N_8991);
xnor U15794 (N_15794,N_7678,N_9733);
or U15795 (N_15795,N_6438,N_11376);
nor U15796 (N_15796,N_9930,N_10010);
nor U15797 (N_15797,N_8856,N_6388);
nand U15798 (N_15798,N_9653,N_7911);
nor U15799 (N_15799,N_9088,N_7589);
xor U15800 (N_15800,N_9153,N_9719);
nor U15801 (N_15801,N_8847,N_9786);
xor U15802 (N_15802,N_6970,N_12091);
and U15803 (N_15803,N_8187,N_7438);
nor U15804 (N_15804,N_9668,N_8489);
xnor U15805 (N_15805,N_7901,N_9031);
nand U15806 (N_15806,N_8957,N_7308);
xnor U15807 (N_15807,N_9549,N_11838);
and U15808 (N_15808,N_8064,N_11330);
nand U15809 (N_15809,N_6558,N_11238);
xnor U15810 (N_15810,N_6392,N_12292);
and U15811 (N_15811,N_8236,N_6345);
nand U15812 (N_15812,N_6672,N_7619);
nor U15813 (N_15813,N_9035,N_7256);
nor U15814 (N_15814,N_6602,N_7134);
and U15815 (N_15815,N_12040,N_10015);
nor U15816 (N_15816,N_7889,N_9913);
or U15817 (N_15817,N_9275,N_10118);
and U15818 (N_15818,N_6400,N_6628);
xnor U15819 (N_15819,N_12361,N_7260);
and U15820 (N_15820,N_8140,N_6697);
or U15821 (N_15821,N_11407,N_11668);
or U15822 (N_15822,N_9323,N_6524);
and U15823 (N_15823,N_8427,N_12467);
nor U15824 (N_15824,N_8218,N_11443);
or U15825 (N_15825,N_12037,N_11013);
nor U15826 (N_15826,N_9653,N_6888);
and U15827 (N_15827,N_11929,N_10268);
nor U15828 (N_15828,N_6409,N_7665);
or U15829 (N_15829,N_8286,N_11793);
and U15830 (N_15830,N_8905,N_6990);
nor U15831 (N_15831,N_11601,N_9574);
and U15832 (N_15832,N_8177,N_11043);
xnor U15833 (N_15833,N_7129,N_10998);
and U15834 (N_15834,N_11189,N_10469);
xnor U15835 (N_15835,N_8369,N_12190);
nor U15836 (N_15836,N_12347,N_8648);
nand U15837 (N_15837,N_9158,N_10993);
or U15838 (N_15838,N_10370,N_9182);
xor U15839 (N_15839,N_7147,N_11887);
nor U15840 (N_15840,N_8477,N_6649);
and U15841 (N_15841,N_11729,N_9125);
nor U15842 (N_15842,N_9394,N_6877);
or U15843 (N_15843,N_8249,N_10767);
nor U15844 (N_15844,N_10062,N_10795);
nand U15845 (N_15845,N_8251,N_8363);
nor U15846 (N_15846,N_7079,N_8547);
xnor U15847 (N_15847,N_6378,N_9264);
nor U15848 (N_15848,N_11222,N_9150);
nor U15849 (N_15849,N_8212,N_6747);
xor U15850 (N_15850,N_11584,N_9671);
nand U15851 (N_15851,N_9217,N_7562);
or U15852 (N_15852,N_7637,N_10686);
or U15853 (N_15853,N_7783,N_11529);
and U15854 (N_15854,N_11620,N_6872);
nor U15855 (N_15855,N_10687,N_8112);
or U15856 (N_15856,N_9356,N_8677);
nor U15857 (N_15857,N_10310,N_11785);
or U15858 (N_15858,N_7711,N_7500);
nor U15859 (N_15859,N_8367,N_9514);
nand U15860 (N_15860,N_10672,N_8441);
nor U15861 (N_15861,N_11907,N_6705);
or U15862 (N_15862,N_7476,N_10902);
xor U15863 (N_15863,N_11173,N_7148);
nor U15864 (N_15864,N_9233,N_7741);
xnor U15865 (N_15865,N_10103,N_7063);
and U15866 (N_15866,N_11451,N_8101);
or U15867 (N_15867,N_11635,N_10531);
nand U15868 (N_15868,N_6504,N_10844);
or U15869 (N_15869,N_10011,N_9770);
and U15870 (N_15870,N_11677,N_10637);
nand U15871 (N_15871,N_7055,N_11821);
xnor U15872 (N_15872,N_10089,N_7920);
nand U15873 (N_15873,N_7937,N_9399);
nand U15874 (N_15874,N_10300,N_10639);
nor U15875 (N_15875,N_10019,N_6641);
and U15876 (N_15876,N_7912,N_8697);
nand U15877 (N_15877,N_9049,N_11259);
or U15878 (N_15878,N_10086,N_8383);
nor U15879 (N_15879,N_8854,N_10691);
nor U15880 (N_15880,N_10559,N_7043);
nor U15881 (N_15881,N_11467,N_6657);
nand U15882 (N_15882,N_7186,N_7420);
nand U15883 (N_15883,N_7270,N_10420);
nor U15884 (N_15884,N_9712,N_8370);
xor U15885 (N_15885,N_10961,N_8705);
and U15886 (N_15886,N_8532,N_7286);
nor U15887 (N_15887,N_7963,N_7565);
or U15888 (N_15888,N_7965,N_8249);
nand U15889 (N_15889,N_9345,N_9495);
nand U15890 (N_15890,N_11677,N_10704);
and U15891 (N_15891,N_7334,N_12402);
nand U15892 (N_15892,N_9845,N_10084);
nand U15893 (N_15893,N_10633,N_10310);
or U15894 (N_15894,N_10213,N_8138);
or U15895 (N_15895,N_8708,N_11169);
nand U15896 (N_15896,N_10334,N_9356);
nand U15897 (N_15897,N_12316,N_11855);
and U15898 (N_15898,N_8011,N_7847);
and U15899 (N_15899,N_10673,N_12059);
nand U15900 (N_15900,N_7457,N_7266);
nor U15901 (N_15901,N_7507,N_12171);
or U15902 (N_15902,N_9421,N_8761);
and U15903 (N_15903,N_11927,N_8449);
and U15904 (N_15904,N_7163,N_8171);
nand U15905 (N_15905,N_8867,N_10849);
nand U15906 (N_15906,N_11132,N_10455);
or U15907 (N_15907,N_6494,N_10537);
or U15908 (N_15908,N_7218,N_11235);
xnor U15909 (N_15909,N_7260,N_8434);
nand U15910 (N_15910,N_8909,N_12481);
xnor U15911 (N_15911,N_11763,N_10025);
nor U15912 (N_15912,N_10092,N_8960);
nor U15913 (N_15913,N_10272,N_7576);
nor U15914 (N_15914,N_9906,N_6306);
and U15915 (N_15915,N_10866,N_9108);
nor U15916 (N_15916,N_7146,N_10382);
or U15917 (N_15917,N_9399,N_7506);
nand U15918 (N_15918,N_11562,N_8767);
nor U15919 (N_15919,N_9977,N_6740);
nand U15920 (N_15920,N_7570,N_7475);
or U15921 (N_15921,N_6347,N_6700);
or U15922 (N_15922,N_11240,N_9092);
or U15923 (N_15923,N_7596,N_8816);
nor U15924 (N_15924,N_7208,N_7082);
nor U15925 (N_15925,N_8644,N_10389);
and U15926 (N_15926,N_10606,N_7205);
and U15927 (N_15927,N_6928,N_12047);
and U15928 (N_15928,N_7303,N_8723);
and U15929 (N_15929,N_10555,N_10848);
and U15930 (N_15930,N_11722,N_9198);
and U15931 (N_15931,N_7349,N_11796);
and U15932 (N_15932,N_9883,N_6604);
and U15933 (N_15933,N_9956,N_7083);
and U15934 (N_15934,N_6945,N_11378);
nand U15935 (N_15935,N_6813,N_8173);
nor U15936 (N_15936,N_10191,N_6976);
and U15937 (N_15937,N_12475,N_11317);
or U15938 (N_15938,N_10496,N_9987);
or U15939 (N_15939,N_11678,N_6821);
or U15940 (N_15940,N_11112,N_9747);
or U15941 (N_15941,N_7399,N_9266);
xnor U15942 (N_15942,N_10376,N_8125);
and U15943 (N_15943,N_10604,N_11566);
and U15944 (N_15944,N_9285,N_10944);
nand U15945 (N_15945,N_6893,N_10033);
xnor U15946 (N_15946,N_11503,N_10903);
or U15947 (N_15947,N_7824,N_12312);
xor U15948 (N_15948,N_8719,N_9992);
or U15949 (N_15949,N_7017,N_12455);
or U15950 (N_15950,N_10766,N_8051);
and U15951 (N_15951,N_8302,N_8500);
and U15952 (N_15952,N_9877,N_6267);
xnor U15953 (N_15953,N_11937,N_7980);
xnor U15954 (N_15954,N_10679,N_9336);
or U15955 (N_15955,N_12186,N_9173);
xor U15956 (N_15956,N_6641,N_6364);
xnor U15957 (N_15957,N_8243,N_8599);
nor U15958 (N_15958,N_6942,N_7984);
nor U15959 (N_15959,N_7637,N_11071);
nor U15960 (N_15960,N_9933,N_11011);
or U15961 (N_15961,N_10652,N_10774);
nor U15962 (N_15962,N_9478,N_12084);
and U15963 (N_15963,N_11297,N_10674);
or U15964 (N_15964,N_8884,N_6488);
and U15965 (N_15965,N_9435,N_9925);
and U15966 (N_15966,N_11101,N_9085);
nor U15967 (N_15967,N_11313,N_9035);
and U15968 (N_15968,N_9216,N_12497);
nand U15969 (N_15969,N_9157,N_11579);
or U15970 (N_15970,N_12098,N_6719);
nor U15971 (N_15971,N_8466,N_8410);
nand U15972 (N_15972,N_6408,N_9953);
or U15973 (N_15973,N_8621,N_7319);
nand U15974 (N_15974,N_9005,N_8369);
xor U15975 (N_15975,N_9589,N_8954);
nor U15976 (N_15976,N_8431,N_11532);
nand U15977 (N_15977,N_6473,N_8450);
nor U15978 (N_15978,N_11072,N_7247);
and U15979 (N_15979,N_7301,N_9089);
or U15980 (N_15980,N_9347,N_11783);
nand U15981 (N_15981,N_6882,N_11413);
xor U15982 (N_15982,N_6982,N_6294);
and U15983 (N_15983,N_7841,N_7296);
nand U15984 (N_15984,N_11318,N_11997);
xnor U15985 (N_15985,N_12227,N_7656);
xor U15986 (N_15986,N_10263,N_9181);
or U15987 (N_15987,N_6748,N_12216);
nand U15988 (N_15988,N_7777,N_11050);
nand U15989 (N_15989,N_11001,N_12035);
nand U15990 (N_15990,N_10491,N_10204);
xnor U15991 (N_15991,N_10930,N_6905);
and U15992 (N_15992,N_9828,N_6265);
and U15993 (N_15993,N_6780,N_6805);
nor U15994 (N_15994,N_11131,N_10759);
or U15995 (N_15995,N_9101,N_9075);
and U15996 (N_15996,N_8100,N_12113);
or U15997 (N_15997,N_11925,N_9567);
nand U15998 (N_15998,N_9311,N_11001);
and U15999 (N_15999,N_6750,N_9250);
and U16000 (N_16000,N_10315,N_10992);
or U16001 (N_16001,N_11235,N_10139);
and U16002 (N_16002,N_11597,N_10282);
and U16003 (N_16003,N_8121,N_6590);
nand U16004 (N_16004,N_8271,N_7280);
and U16005 (N_16005,N_10029,N_10430);
or U16006 (N_16006,N_11630,N_12166);
nand U16007 (N_16007,N_6274,N_7151);
or U16008 (N_16008,N_8643,N_7600);
or U16009 (N_16009,N_9291,N_7742);
and U16010 (N_16010,N_9466,N_10024);
xnor U16011 (N_16011,N_6898,N_12008);
or U16012 (N_16012,N_8952,N_9841);
nor U16013 (N_16013,N_9878,N_10016);
or U16014 (N_16014,N_10625,N_12257);
and U16015 (N_16015,N_9169,N_6861);
or U16016 (N_16016,N_12303,N_6902);
xnor U16017 (N_16017,N_8453,N_9337);
nand U16018 (N_16018,N_10828,N_7643);
or U16019 (N_16019,N_7233,N_9926);
nor U16020 (N_16020,N_8803,N_11017);
and U16021 (N_16021,N_9821,N_11410);
or U16022 (N_16022,N_7643,N_9853);
nand U16023 (N_16023,N_6627,N_6653);
xnor U16024 (N_16024,N_11831,N_10260);
and U16025 (N_16025,N_10124,N_7322);
xor U16026 (N_16026,N_10502,N_11967);
nand U16027 (N_16027,N_9973,N_10641);
nand U16028 (N_16028,N_6532,N_7914);
nand U16029 (N_16029,N_11919,N_11476);
or U16030 (N_16030,N_10474,N_7373);
nand U16031 (N_16031,N_8647,N_6450);
and U16032 (N_16032,N_11912,N_10677);
xnor U16033 (N_16033,N_12431,N_9662);
nor U16034 (N_16034,N_6337,N_9335);
nor U16035 (N_16035,N_7440,N_6302);
xnor U16036 (N_16036,N_7364,N_7129);
and U16037 (N_16037,N_7752,N_8549);
nor U16038 (N_16038,N_10935,N_7746);
xor U16039 (N_16039,N_11138,N_7739);
and U16040 (N_16040,N_7743,N_6954);
and U16041 (N_16041,N_9139,N_6834);
nor U16042 (N_16042,N_11021,N_8582);
nor U16043 (N_16043,N_11744,N_8416);
nand U16044 (N_16044,N_7496,N_8865);
or U16045 (N_16045,N_6492,N_8170);
nor U16046 (N_16046,N_7797,N_9985);
or U16047 (N_16047,N_12144,N_10854);
xor U16048 (N_16048,N_12378,N_6783);
or U16049 (N_16049,N_6791,N_12036);
xnor U16050 (N_16050,N_7228,N_8437);
or U16051 (N_16051,N_7101,N_11011);
or U16052 (N_16052,N_9282,N_8007);
nor U16053 (N_16053,N_9551,N_10473);
and U16054 (N_16054,N_10654,N_10208);
or U16055 (N_16055,N_9720,N_10790);
xor U16056 (N_16056,N_10875,N_11216);
xnor U16057 (N_16057,N_12468,N_10850);
or U16058 (N_16058,N_9569,N_10274);
nor U16059 (N_16059,N_9288,N_7030);
nand U16060 (N_16060,N_8217,N_12274);
nor U16061 (N_16061,N_10133,N_8864);
nor U16062 (N_16062,N_7029,N_11228);
and U16063 (N_16063,N_12385,N_6278);
nand U16064 (N_16064,N_6910,N_11247);
or U16065 (N_16065,N_10390,N_12473);
and U16066 (N_16066,N_8335,N_7289);
nand U16067 (N_16067,N_10397,N_12175);
or U16068 (N_16068,N_8093,N_10240);
nor U16069 (N_16069,N_9702,N_6349);
and U16070 (N_16070,N_10634,N_6856);
xnor U16071 (N_16071,N_7095,N_6512);
nand U16072 (N_16072,N_6883,N_8185);
and U16073 (N_16073,N_11294,N_11629);
xnor U16074 (N_16074,N_9271,N_10976);
nor U16075 (N_16075,N_10456,N_12086);
nand U16076 (N_16076,N_7341,N_10587);
nand U16077 (N_16077,N_11749,N_7559);
nand U16078 (N_16078,N_7008,N_9372);
or U16079 (N_16079,N_6942,N_12211);
nand U16080 (N_16080,N_9235,N_9429);
nor U16081 (N_16081,N_10053,N_12467);
nor U16082 (N_16082,N_10606,N_9484);
xor U16083 (N_16083,N_9376,N_6334);
and U16084 (N_16084,N_7198,N_9176);
or U16085 (N_16085,N_9629,N_11821);
and U16086 (N_16086,N_7101,N_10352);
and U16087 (N_16087,N_8614,N_8507);
nor U16088 (N_16088,N_10014,N_8996);
nand U16089 (N_16089,N_6553,N_7546);
or U16090 (N_16090,N_6689,N_12144);
xnor U16091 (N_16091,N_7710,N_9596);
and U16092 (N_16092,N_6318,N_7753);
nor U16093 (N_16093,N_8815,N_9829);
nor U16094 (N_16094,N_12077,N_10534);
nor U16095 (N_16095,N_8621,N_10335);
nand U16096 (N_16096,N_9033,N_7241);
xnor U16097 (N_16097,N_9186,N_8698);
nor U16098 (N_16098,N_11422,N_11513);
xnor U16099 (N_16099,N_8827,N_11658);
nand U16100 (N_16100,N_9382,N_8547);
nor U16101 (N_16101,N_7443,N_7292);
and U16102 (N_16102,N_11053,N_12263);
and U16103 (N_16103,N_8228,N_6909);
or U16104 (N_16104,N_11012,N_8481);
nor U16105 (N_16105,N_6967,N_10918);
nand U16106 (N_16106,N_7631,N_9151);
and U16107 (N_16107,N_10169,N_6832);
nor U16108 (N_16108,N_8577,N_6733);
or U16109 (N_16109,N_12305,N_9696);
nand U16110 (N_16110,N_9830,N_10335);
xor U16111 (N_16111,N_8595,N_7901);
or U16112 (N_16112,N_10760,N_10105);
and U16113 (N_16113,N_10210,N_7723);
nor U16114 (N_16114,N_11450,N_6308);
and U16115 (N_16115,N_6660,N_9760);
nor U16116 (N_16116,N_7963,N_9025);
and U16117 (N_16117,N_6877,N_8260);
or U16118 (N_16118,N_8929,N_9599);
xnor U16119 (N_16119,N_7936,N_8404);
and U16120 (N_16120,N_6512,N_10345);
nor U16121 (N_16121,N_8515,N_6833);
or U16122 (N_16122,N_8477,N_6508);
and U16123 (N_16123,N_8142,N_11375);
nand U16124 (N_16124,N_12442,N_6642);
xnor U16125 (N_16125,N_6615,N_10403);
and U16126 (N_16126,N_9012,N_9850);
xor U16127 (N_16127,N_9889,N_8990);
xnor U16128 (N_16128,N_9638,N_6815);
nor U16129 (N_16129,N_8003,N_8860);
or U16130 (N_16130,N_11484,N_12153);
xor U16131 (N_16131,N_6747,N_6285);
xnor U16132 (N_16132,N_6965,N_6303);
and U16133 (N_16133,N_12255,N_9751);
nand U16134 (N_16134,N_7584,N_8529);
xor U16135 (N_16135,N_8527,N_8790);
nand U16136 (N_16136,N_6629,N_8460);
xor U16137 (N_16137,N_10672,N_8127);
and U16138 (N_16138,N_11005,N_7182);
or U16139 (N_16139,N_6912,N_12203);
xnor U16140 (N_16140,N_10014,N_10113);
or U16141 (N_16141,N_8443,N_8748);
or U16142 (N_16142,N_10688,N_10778);
and U16143 (N_16143,N_10354,N_8654);
nor U16144 (N_16144,N_10131,N_10993);
or U16145 (N_16145,N_6977,N_9493);
or U16146 (N_16146,N_7641,N_10666);
xor U16147 (N_16147,N_11238,N_9061);
or U16148 (N_16148,N_10121,N_8817);
or U16149 (N_16149,N_9073,N_10227);
or U16150 (N_16150,N_7095,N_12244);
or U16151 (N_16151,N_8953,N_7452);
nor U16152 (N_16152,N_12384,N_9247);
and U16153 (N_16153,N_12334,N_11164);
nand U16154 (N_16154,N_10681,N_10123);
and U16155 (N_16155,N_9001,N_8040);
nor U16156 (N_16156,N_9233,N_12302);
xnor U16157 (N_16157,N_11301,N_9219);
or U16158 (N_16158,N_6399,N_8182);
and U16159 (N_16159,N_7611,N_7866);
and U16160 (N_16160,N_8600,N_9796);
nand U16161 (N_16161,N_6665,N_8399);
and U16162 (N_16162,N_10917,N_11092);
and U16163 (N_16163,N_10540,N_10165);
and U16164 (N_16164,N_8727,N_7731);
nor U16165 (N_16165,N_8331,N_9482);
nand U16166 (N_16166,N_7498,N_8680);
nand U16167 (N_16167,N_8012,N_7916);
xor U16168 (N_16168,N_8376,N_6263);
xor U16169 (N_16169,N_7600,N_6722);
or U16170 (N_16170,N_10890,N_8212);
and U16171 (N_16171,N_9072,N_7929);
and U16172 (N_16172,N_7239,N_11317);
or U16173 (N_16173,N_7298,N_9231);
xor U16174 (N_16174,N_7036,N_9281);
and U16175 (N_16175,N_12457,N_12091);
nor U16176 (N_16176,N_9664,N_7905);
or U16177 (N_16177,N_7565,N_10532);
nand U16178 (N_16178,N_6795,N_9694);
nand U16179 (N_16179,N_6893,N_8574);
or U16180 (N_16180,N_9665,N_11793);
nand U16181 (N_16181,N_9477,N_9671);
nand U16182 (N_16182,N_8870,N_6653);
xor U16183 (N_16183,N_11156,N_9989);
nand U16184 (N_16184,N_9122,N_11422);
or U16185 (N_16185,N_9446,N_8087);
nor U16186 (N_16186,N_11976,N_10136);
xnor U16187 (N_16187,N_6403,N_7036);
or U16188 (N_16188,N_8344,N_8041);
or U16189 (N_16189,N_11699,N_9660);
or U16190 (N_16190,N_7889,N_11411);
nand U16191 (N_16191,N_11658,N_10554);
and U16192 (N_16192,N_12186,N_7083);
nand U16193 (N_16193,N_11846,N_12096);
nor U16194 (N_16194,N_11833,N_12441);
nor U16195 (N_16195,N_10472,N_9935);
or U16196 (N_16196,N_11257,N_11168);
and U16197 (N_16197,N_9118,N_10776);
or U16198 (N_16198,N_7541,N_12363);
nand U16199 (N_16199,N_10162,N_6506);
nand U16200 (N_16200,N_12058,N_7841);
nor U16201 (N_16201,N_6872,N_9584);
and U16202 (N_16202,N_10493,N_8887);
nor U16203 (N_16203,N_9165,N_8849);
nand U16204 (N_16204,N_9900,N_9336);
and U16205 (N_16205,N_8976,N_8987);
xor U16206 (N_16206,N_9854,N_6506);
nor U16207 (N_16207,N_11161,N_7558);
or U16208 (N_16208,N_10447,N_10510);
or U16209 (N_16209,N_6960,N_7479);
and U16210 (N_16210,N_8234,N_8540);
xor U16211 (N_16211,N_11231,N_10339);
xor U16212 (N_16212,N_11623,N_12242);
nor U16213 (N_16213,N_9724,N_7165);
and U16214 (N_16214,N_10708,N_10977);
and U16215 (N_16215,N_10939,N_10120);
nor U16216 (N_16216,N_11093,N_7675);
and U16217 (N_16217,N_6337,N_7673);
xnor U16218 (N_16218,N_12339,N_8878);
nor U16219 (N_16219,N_11715,N_6945);
and U16220 (N_16220,N_7236,N_12012);
nor U16221 (N_16221,N_7287,N_9293);
nand U16222 (N_16222,N_6434,N_11608);
nor U16223 (N_16223,N_8078,N_6884);
xor U16224 (N_16224,N_7123,N_11725);
nand U16225 (N_16225,N_8343,N_7411);
xnor U16226 (N_16226,N_7010,N_8107);
nor U16227 (N_16227,N_8990,N_10647);
or U16228 (N_16228,N_6851,N_9540);
or U16229 (N_16229,N_8932,N_9387);
or U16230 (N_16230,N_9498,N_11102);
nor U16231 (N_16231,N_7306,N_11371);
or U16232 (N_16232,N_7959,N_7036);
nand U16233 (N_16233,N_11440,N_9935);
xor U16234 (N_16234,N_6741,N_11247);
and U16235 (N_16235,N_7597,N_8874);
nor U16236 (N_16236,N_11194,N_7181);
nor U16237 (N_16237,N_6888,N_9116);
xor U16238 (N_16238,N_7465,N_12109);
and U16239 (N_16239,N_9494,N_9238);
nand U16240 (N_16240,N_10553,N_8174);
xnor U16241 (N_16241,N_7283,N_7218);
xnor U16242 (N_16242,N_9880,N_7372);
xnor U16243 (N_16243,N_7590,N_11371);
nor U16244 (N_16244,N_10356,N_8742);
nand U16245 (N_16245,N_7662,N_6366);
xor U16246 (N_16246,N_8128,N_10394);
xnor U16247 (N_16247,N_7016,N_8666);
and U16248 (N_16248,N_9431,N_10420);
nand U16249 (N_16249,N_8293,N_8153);
and U16250 (N_16250,N_11941,N_8603);
and U16251 (N_16251,N_11849,N_6523);
or U16252 (N_16252,N_12231,N_8716);
xor U16253 (N_16253,N_8646,N_7800);
xor U16254 (N_16254,N_10150,N_8100);
xnor U16255 (N_16255,N_12297,N_11879);
and U16256 (N_16256,N_11180,N_11479);
xnor U16257 (N_16257,N_11913,N_8326);
nor U16258 (N_16258,N_10007,N_8332);
and U16259 (N_16259,N_10546,N_11479);
nor U16260 (N_16260,N_12162,N_10363);
or U16261 (N_16261,N_8164,N_10089);
nor U16262 (N_16262,N_6585,N_10836);
nand U16263 (N_16263,N_11296,N_8796);
or U16264 (N_16264,N_9968,N_10372);
nor U16265 (N_16265,N_9932,N_7596);
xor U16266 (N_16266,N_6926,N_10151);
and U16267 (N_16267,N_9606,N_10110);
or U16268 (N_16268,N_7374,N_8612);
or U16269 (N_16269,N_10308,N_8861);
and U16270 (N_16270,N_7643,N_11278);
nor U16271 (N_16271,N_10626,N_6837);
or U16272 (N_16272,N_10943,N_8641);
or U16273 (N_16273,N_8559,N_9936);
and U16274 (N_16274,N_7720,N_10076);
and U16275 (N_16275,N_12302,N_8261);
nor U16276 (N_16276,N_6298,N_12225);
xor U16277 (N_16277,N_9877,N_8792);
xor U16278 (N_16278,N_12236,N_6353);
nor U16279 (N_16279,N_10716,N_11949);
xor U16280 (N_16280,N_10670,N_12489);
and U16281 (N_16281,N_6562,N_10540);
nor U16282 (N_16282,N_8416,N_12043);
nor U16283 (N_16283,N_11573,N_8855);
or U16284 (N_16284,N_11740,N_6922);
or U16285 (N_16285,N_10586,N_11241);
nand U16286 (N_16286,N_12366,N_8983);
and U16287 (N_16287,N_10757,N_8333);
and U16288 (N_16288,N_7614,N_6325);
nand U16289 (N_16289,N_7312,N_7496);
nor U16290 (N_16290,N_8845,N_10227);
or U16291 (N_16291,N_9082,N_8597);
xor U16292 (N_16292,N_8414,N_7895);
xnor U16293 (N_16293,N_9928,N_10438);
or U16294 (N_16294,N_12127,N_8535);
and U16295 (N_16295,N_8908,N_6847);
or U16296 (N_16296,N_9129,N_10482);
xor U16297 (N_16297,N_7024,N_8160);
nor U16298 (N_16298,N_8173,N_10968);
nand U16299 (N_16299,N_9716,N_8087);
nor U16300 (N_16300,N_9702,N_11262);
nand U16301 (N_16301,N_10476,N_11461);
and U16302 (N_16302,N_9821,N_8560);
or U16303 (N_16303,N_9581,N_9452);
xor U16304 (N_16304,N_8027,N_8481);
xnor U16305 (N_16305,N_8901,N_12290);
or U16306 (N_16306,N_11247,N_10107);
nor U16307 (N_16307,N_9144,N_11253);
and U16308 (N_16308,N_6907,N_11363);
and U16309 (N_16309,N_7891,N_10152);
nor U16310 (N_16310,N_12074,N_7193);
nand U16311 (N_16311,N_12411,N_10788);
xor U16312 (N_16312,N_10243,N_7577);
or U16313 (N_16313,N_7442,N_10235);
or U16314 (N_16314,N_12360,N_8998);
nor U16315 (N_16315,N_7262,N_10121);
xnor U16316 (N_16316,N_6481,N_9836);
xnor U16317 (N_16317,N_11776,N_9467);
nor U16318 (N_16318,N_7574,N_6703);
and U16319 (N_16319,N_6815,N_9490);
or U16320 (N_16320,N_9936,N_7178);
xnor U16321 (N_16321,N_12408,N_6472);
and U16322 (N_16322,N_9629,N_7634);
xnor U16323 (N_16323,N_7480,N_7854);
nand U16324 (N_16324,N_8806,N_8845);
xor U16325 (N_16325,N_7329,N_12236);
nand U16326 (N_16326,N_11755,N_10456);
xnor U16327 (N_16327,N_6372,N_6536);
nand U16328 (N_16328,N_9701,N_9560);
nand U16329 (N_16329,N_7329,N_11119);
xor U16330 (N_16330,N_10145,N_11014);
xor U16331 (N_16331,N_11289,N_7797);
and U16332 (N_16332,N_7045,N_8469);
nand U16333 (N_16333,N_10895,N_10882);
nor U16334 (N_16334,N_7494,N_9344);
and U16335 (N_16335,N_11839,N_6989);
or U16336 (N_16336,N_11885,N_10189);
nand U16337 (N_16337,N_8067,N_9145);
xor U16338 (N_16338,N_8360,N_10480);
nor U16339 (N_16339,N_8310,N_11173);
xor U16340 (N_16340,N_10891,N_7605);
nor U16341 (N_16341,N_6346,N_11774);
or U16342 (N_16342,N_9247,N_10412);
nor U16343 (N_16343,N_9531,N_11348);
nand U16344 (N_16344,N_9404,N_7292);
nor U16345 (N_16345,N_10057,N_6677);
xnor U16346 (N_16346,N_6297,N_9530);
nand U16347 (N_16347,N_11910,N_6459);
or U16348 (N_16348,N_9698,N_10131);
and U16349 (N_16349,N_10949,N_10362);
xnor U16350 (N_16350,N_11790,N_11415);
xnor U16351 (N_16351,N_8321,N_10188);
nand U16352 (N_16352,N_8852,N_9207);
or U16353 (N_16353,N_7540,N_11214);
nand U16354 (N_16354,N_10786,N_9068);
xnor U16355 (N_16355,N_10630,N_7578);
nand U16356 (N_16356,N_8679,N_9331);
nor U16357 (N_16357,N_9756,N_10201);
nor U16358 (N_16358,N_11631,N_12492);
nand U16359 (N_16359,N_8517,N_10842);
and U16360 (N_16360,N_11455,N_9141);
and U16361 (N_16361,N_12256,N_7312);
xor U16362 (N_16362,N_9051,N_6424);
or U16363 (N_16363,N_11744,N_9412);
and U16364 (N_16364,N_12080,N_8136);
or U16365 (N_16365,N_9074,N_8615);
or U16366 (N_16366,N_7673,N_11072);
nor U16367 (N_16367,N_11269,N_12152);
nand U16368 (N_16368,N_11720,N_7342);
and U16369 (N_16369,N_11044,N_7200);
nand U16370 (N_16370,N_10893,N_7031);
or U16371 (N_16371,N_11783,N_7537);
or U16372 (N_16372,N_12308,N_12438);
and U16373 (N_16373,N_9975,N_9558);
xor U16374 (N_16374,N_9110,N_7003);
nor U16375 (N_16375,N_8127,N_7243);
or U16376 (N_16376,N_7675,N_11833);
xnor U16377 (N_16377,N_12440,N_9200);
nand U16378 (N_16378,N_8798,N_7308);
or U16379 (N_16379,N_11761,N_7435);
nand U16380 (N_16380,N_10393,N_9388);
or U16381 (N_16381,N_8134,N_8335);
xnor U16382 (N_16382,N_10411,N_10174);
and U16383 (N_16383,N_8753,N_12205);
nand U16384 (N_16384,N_11823,N_7327);
xor U16385 (N_16385,N_8658,N_6466);
nor U16386 (N_16386,N_11058,N_8963);
xnor U16387 (N_16387,N_10047,N_6743);
or U16388 (N_16388,N_7655,N_11557);
nor U16389 (N_16389,N_8816,N_9976);
nor U16390 (N_16390,N_9342,N_11745);
nand U16391 (N_16391,N_6436,N_6710);
and U16392 (N_16392,N_10715,N_7794);
and U16393 (N_16393,N_9665,N_9153);
or U16394 (N_16394,N_10075,N_8181);
nor U16395 (N_16395,N_11306,N_8451);
and U16396 (N_16396,N_7408,N_10920);
nand U16397 (N_16397,N_8966,N_9138);
nor U16398 (N_16398,N_7368,N_11329);
xor U16399 (N_16399,N_7784,N_11555);
nand U16400 (N_16400,N_10767,N_6504);
nor U16401 (N_16401,N_11438,N_10482);
and U16402 (N_16402,N_8667,N_8511);
xnor U16403 (N_16403,N_6314,N_10170);
or U16404 (N_16404,N_11772,N_6906);
and U16405 (N_16405,N_10221,N_7157);
or U16406 (N_16406,N_12181,N_9172);
nand U16407 (N_16407,N_8919,N_9864);
nor U16408 (N_16408,N_9952,N_6500);
xnor U16409 (N_16409,N_8375,N_11244);
xnor U16410 (N_16410,N_7436,N_8989);
or U16411 (N_16411,N_7573,N_10728);
nor U16412 (N_16412,N_12208,N_10323);
nor U16413 (N_16413,N_8419,N_9843);
nor U16414 (N_16414,N_10468,N_7587);
xnor U16415 (N_16415,N_9029,N_11066);
or U16416 (N_16416,N_8986,N_10009);
and U16417 (N_16417,N_6426,N_10486);
or U16418 (N_16418,N_6693,N_7515);
nor U16419 (N_16419,N_11980,N_6370);
nor U16420 (N_16420,N_9194,N_9972);
xor U16421 (N_16421,N_12389,N_12187);
nor U16422 (N_16422,N_10166,N_12324);
xor U16423 (N_16423,N_11277,N_6792);
nand U16424 (N_16424,N_10336,N_10758);
nor U16425 (N_16425,N_8704,N_7533);
and U16426 (N_16426,N_11235,N_11439);
and U16427 (N_16427,N_9911,N_10470);
and U16428 (N_16428,N_7245,N_10276);
and U16429 (N_16429,N_12365,N_10795);
nand U16430 (N_16430,N_9645,N_11560);
nand U16431 (N_16431,N_7063,N_10313);
xnor U16432 (N_16432,N_8277,N_6523);
xor U16433 (N_16433,N_11914,N_6968);
xnor U16434 (N_16434,N_9452,N_9134);
or U16435 (N_16435,N_9477,N_7000);
xor U16436 (N_16436,N_8222,N_7399);
nand U16437 (N_16437,N_9727,N_11677);
xnor U16438 (N_16438,N_8278,N_12017);
and U16439 (N_16439,N_12204,N_6354);
or U16440 (N_16440,N_11748,N_9878);
and U16441 (N_16441,N_7569,N_7822);
nor U16442 (N_16442,N_12017,N_10525);
nand U16443 (N_16443,N_7382,N_6302);
or U16444 (N_16444,N_9146,N_8915);
or U16445 (N_16445,N_8508,N_9252);
or U16446 (N_16446,N_9742,N_6737);
nor U16447 (N_16447,N_12246,N_10741);
and U16448 (N_16448,N_7282,N_9639);
xor U16449 (N_16449,N_10068,N_9945);
or U16450 (N_16450,N_7650,N_8364);
nor U16451 (N_16451,N_9864,N_8033);
and U16452 (N_16452,N_9846,N_9012);
nor U16453 (N_16453,N_7249,N_8520);
nand U16454 (N_16454,N_11021,N_6417);
nor U16455 (N_16455,N_9241,N_6504);
nand U16456 (N_16456,N_10044,N_6805);
nor U16457 (N_16457,N_8560,N_9713);
nand U16458 (N_16458,N_8635,N_8625);
nand U16459 (N_16459,N_10086,N_11509);
xor U16460 (N_16460,N_12135,N_8403);
nor U16461 (N_16461,N_9214,N_11686);
and U16462 (N_16462,N_6316,N_7002);
nor U16463 (N_16463,N_9135,N_9618);
xor U16464 (N_16464,N_10839,N_8688);
nor U16465 (N_16465,N_6444,N_7478);
or U16466 (N_16466,N_6995,N_8453);
and U16467 (N_16467,N_8720,N_11997);
xor U16468 (N_16468,N_11508,N_9306);
and U16469 (N_16469,N_12042,N_8899);
and U16470 (N_16470,N_11517,N_8617);
and U16471 (N_16471,N_8029,N_8958);
and U16472 (N_16472,N_11331,N_8257);
nor U16473 (N_16473,N_7981,N_11617);
xor U16474 (N_16474,N_10413,N_10404);
nor U16475 (N_16475,N_9399,N_7100);
and U16476 (N_16476,N_9616,N_6376);
or U16477 (N_16477,N_9605,N_11215);
xor U16478 (N_16478,N_6403,N_9357);
xor U16479 (N_16479,N_9669,N_7648);
nand U16480 (N_16480,N_9100,N_6976);
xnor U16481 (N_16481,N_9064,N_8482);
nor U16482 (N_16482,N_10953,N_12194);
or U16483 (N_16483,N_7212,N_6583);
nand U16484 (N_16484,N_11702,N_8399);
xnor U16485 (N_16485,N_7011,N_11528);
nand U16486 (N_16486,N_9244,N_10864);
or U16487 (N_16487,N_11818,N_6274);
and U16488 (N_16488,N_9353,N_6659);
xnor U16489 (N_16489,N_9086,N_9802);
xnor U16490 (N_16490,N_9829,N_6314);
xor U16491 (N_16491,N_8783,N_11581);
and U16492 (N_16492,N_11388,N_9747);
and U16493 (N_16493,N_9655,N_6446);
nor U16494 (N_16494,N_10500,N_10054);
nor U16495 (N_16495,N_11896,N_11264);
xor U16496 (N_16496,N_8664,N_8166);
or U16497 (N_16497,N_6341,N_9920);
nor U16498 (N_16498,N_9274,N_8740);
or U16499 (N_16499,N_6703,N_7091);
nor U16500 (N_16500,N_12327,N_8805);
and U16501 (N_16501,N_11246,N_8128);
nand U16502 (N_16502,N_10001,N_9274);
or U16503 (N_16503,N_11893,N_10536);
xor U16504 (N_16504,N_12299,N_11342);
nor U16505 (N_16505,N_7361,N_12476);
nand U16506 (N_16506,N_8880,N_11102);
nand U16507 (N_16507,N_6719,N_8990);
nand U16508 (N_16508,N_9120,N_6503);
xor U16509 (N_16509,N_12441,N_7815);
nand U16510 (N_16510,N_12090,N_6590);
nor U16511 (N_16511,N_10646,N_6987);
or U16512 (N_16512,N_7753,N_11375);
nand U16513 (N_16513,N_11049,N_12408);
and U16514 (N_16514,N_10312,N_6420);
or U16515 (N_16515,N_7629,N_11580);
xor U16516 (N_16516,N_12199,N_11019);
nand U16517 (N_16517,N_7477,N_6500);
or U16518 (N_16518,N_11185,N_8928);
and U16519 (N_16519,N_7376,N_7766);
and U16520 (N_16520,N_6345,N_7965);
or U16521 (N_16521,N_6679,N_8968);
nor U16522 (N_16522,N_12022,N_8890);
nor U16523 (N_16523,N_10608,N_10738);
nor U16524 (N_16524,N_12071,N_8185);
nor U16525 (N_16525,N_8950,N_7991);
or U16526 (N_16526,N_8023,N_8441);
or U16527 (N_16527,N_11470,N_11904);
nor U16528 (N_16528,N_12488,N_7042);
or U16529 (N_16529,N_7540,N_8292);
nand U16530 (N_16530,N_9551,N_12415);
xnor U16531 (N_16531,N_7005,N_7782);
nor U16532 (N_16532,N_9097,N_10026);
nor U16533 (N_16533,N_7835,N_9620);
nand U16534 (N_16534,N_9443,N_11955);
or U16535 (N_16535,N_7028,N_9099);
or U16536 (N_16536,N_9811,N_6978);
and U16537 (N_16537,N_7571,N_11297);
xnor U16538 (N_16538,N_10241,N_7721);
and U16539 (N_16539,N_7698,N_9609);
nand U16540 (N_16540,N_9616,N_6978);
xor U16541 (N_16541,N_6337,N_8213);
and U16542 (N_16542,N_6966,N_10782);
nor U16543 (N_16543,N_6258,N_7744);
or U16544 (N_16544,N_8108,N_6404);
and U16545 (N_16545,N_11362,N_8280);
and U16546 (N_16546,N_8831,N_12237);
or U16547 (N_16547,N_8743,N_7922);
nand U16548 (N_16548,N_6768,N_6321);
nand U16549 (N_16549,N_8608,N_12439);
nand U16550 (N_16550,N_7685,N_9882);
and U16551 (N_16551,N_9670,N_6539);
nor U16552 (N_16552,N_9052,N_7312);
and U16553 (N_16553,N_12067,N_6601);
nand U16554 (N_16554,N_8819,N_8061);
nor U16555 (N_16555,N_8871,N_11395);
xnor U16556 (N_16556,N_10966,N_8571);
or U16557 (N_16557,N_8183,N_12290);
xnor U16558 (N_16558,N_9600,N_8319);
and U16559 (N_16559,N_8417,N_8814);
nor U16560 (N_16560,N_7390,N_10353);
nor U16561 (N_16561,N_9597,N_6275);
nand U16562 (N_16562,N_10087,N_10608);
and U16563 (N_16563,N_6840,N_7604);
nor U16564 (N_16564,N_8343,N_10280);
or U16565 (N_16565,N_11728,N_10216);
and U16566 (N_16566,N_12189,N_7416);
and U16567 (N_16567,N_10626,N_11964);
or U16568 (N_16568,N_10521,N_7904);
nor U16569 (N_16569,N_9142,N_9814);
nor U16570 (N_16570,N_9205,N_12057);
or U16571 (N_16571,N_9343,N_9221);
and U16572 (N_16572,N_10514,N_7386);
or U16573 (N_16573,N_12216,N_9271);
xnor U16574 (N_16574,N_12288,N_10725);
or U16575 (N_16575,N_9106,N_6597);
or U16576 (N_16576,N_9880,N_9659);
and U16577 (N_16577,N_8130,N_11309);
xor U16578 (N_16578,N_8658,N_10351);
nor U16579 (N_16579,N_12249,N_7790);
xnor U16580 (N_16580,N_11897,N_10177);
or U16581 (N_16581,N_12296,N_8170);
and U16582 (N_16582,N_11331,N_7326);
nand U16583 (N_16583,N_8099,N_9842);
xnor U16584 (N_16584,N_9854,N_10392);
nor U16585 (N_16585,N_7144,N_6650);
nand U16586 (N_16586,N_12310,N_10907);
nand U16587 (N_16587,N_7197,N_7712);
nand U16588 (N_16588,N_9212,N_8454);
or U16589 (N_16589,N_12022,N_10267);
and U16590 (N_16590,N_9403,N_6599);
nor U16591 (N_16591,N_7453,N_11676);
xor U16592 (N_16592,N_10163,N_7330);
nor U16593 (N_16593,N_8694,N_8812);
nand U16594 (N_16594,N_12068,N_10859);
or U16595 (N_16595,N_7624,N_8890);
nand U16596 (N_16596,N_10671,N_11167);
xnor U16597 (N_16597,N_10096,N_7621);
nor U16598 (N_16598,N_8803,N_11658);
or U16599 (N_16599,N_10439,N_9021);
nor U16600 (N_16600,N_10665,N_12414);
or U16601 (N_16601,N_6828,N_12421);
and U16602 (N_16602,N_10837,N_7552);
nor U16603 (N_16603,N_11283,N_6574);
xor U16604 (N_16604,N_12471,N_10959);
nor U16605 (N_16605,N_8013,N_9298);
nor U16606 (N_16606,N_7994,N_9219);
and U16607 (N_16607,N_12187,N_11751);
and U16608 (N_16608,N_10760,N_6481);
or U16609 (N_16609,N_8217,N_9743);
nor U16610 (N_16610,N_10460,N_8026);
nand U16611 (N_16611,N_10698,N_9738);
nand U16612 (N_16612,N_8210,N_10460);
nor U16613 (N_16613,N_8723,N_8622);
or U16614 (N_16614,N_7579,N_9411);
xor U16615 (N_16615,N_8468,N_7230);
and U16616 (N_16616,N_8636,N_7949);
nor U16617 (N_16617,N_8006,N_9784);
and U16618 (N_16618,N_9489,N_11405);
nand U16619 (N_16619,N_10541,N_7411);
nand U16620 (N_16620,N_6796,N_9664);
or U16621 (N_16621,N_11234,N_8396);
or U16622 (N_16622,N_7339,N_6989);
and U16623 (N_16623,N_8353,N_8678);
xor U16624 (N_16624,N_8348,N_9358);
xor U16625 (N_16625,N_10795,N_9941);
or U16626 (N_16626,N_10868,N_9640);
or U16627 (N_16627,N_11353,N_9734);
xnor U16628 (N_16628,N_7600,N_7841);
and U16629 (N_16629,N_8168,N_6869);
nor U16630 (N_16630,N_11116,N_6373);
and U16631 (N_16631,N_9560,N_10080);
and U16632 (N_16632,N_8648,N_7738);
xnor U16633 (N_16633,N_8153,N_9510);
or U16634 (N_16634,N_9484,N_8864);
nand U16635 (N_16635,N_8172,N_8147);
nand U16636 (N_16636,N_11324,N_7533);
xnor U16637 (N_16637,N_12312,N_8778);
and U16638 (N_16638,N_7031,N_8985);
xor U16639 (N_16639,N_10529,N_9035);
xnor U16640 (N_16640,N_9374,N_10905);
or U16641 (N_16641,N_11273,N_8823);
nor U16642 (N_16642,N_8003,N_9695);
nand U16643 (N_16643,N_10031,N_9073);
xnor U16644 (N_16644,N_10861,N_6402);
xor U16645 (N_16645,N_11215,N_7082);
or U16646 (N_16646,N_9533,N_9895);
xor U16647 (N_16647,N_11177,N_11367);
nor U16648 (N_16648,N_7441,N_11627);
nor U16649 (N_16649,N_6959,N_6546);
nor U16650 (N_16650,N_11997,N_6375);
nand U16651 (N_16651,N_6817,N_7968);
or U16652 (N_16652,N_9882,N_6615);
nand U16653 (N_16653,N_10407,N_9933);
xor U16654 (N_16654,N_9992,N_11680);
or U16655 (N_16655,N_7260,N_8882);
and U16656 (N_16656,N_10438,N_7051);
nor U16657 (N_16657,N_7867,N_7329);
nand U16658 (N_16658,N_9994,N_6255);
or U16659 (N_16659,N_10020,N_6841);
or U16660 (N_16660,N_6996,N_10317);
or U16661 (N_16661,N_6586,N_11755);
nor U16662 (N_16662,N_11545,N_10370);
nor U16663 (N_16663,N_6453,N_10927);
nand U16664 (N_16664,N_7997,N_10530);
xnor U16665 (N_16665,N_12183,N_8788);
xor U16666 (N_16666,N_7405,N_7855);
xor U16667 (N_16667,N_6407,N_11925);
nor U16668 (N_16668,N_9380,N_11943);
and U16669 (N_16669,N_11650,N_12036);
and U16670 (N_16670,N_6657,N_9138);
nand U16671 (N_16671,N_8970,N_8109);
nor U16672 (N_16672,N_8973,N_12096);
nor U16673 (N_16673,N_10884,N_11473);
or U16674 (N_16674,N_12012,N_7562);
nor U16675 (N_16675,N_7329,N_8870);
nand U16676 (N_16676,N_9750,N_11048);
or U16677 (N_16677,N_12281,N_6765);
and U16678 (N_16678,N_7647,N_6628);
nand U16679 (N_16679,N_10696,N_6810);
xnor U16680 (N_16680,N_8845,N_6994);
and U16681 (N_16681,N_11175,N_6962);
and U16682 (N_16682,N_7451,N_10750);
nand U16683 (N_16683,N_11629,N_8411);
nor U16684 (N_16684,N_11539,N_7671);
nand U16685 (N_16685,N_9527,N_7022);
xor U16686 (N_16686,N_7510,N_11334);
and U16687 (N_16687,N_6378,N_8918);
nor U16688 (N_16688,N_7658,N_12128);
or U16689 (N_16689,N_7302,N_7953);
nand U16690 (N_16690,N_9840,N_11553);
or U16691 (N_16691,N_7697,N_7152);
xor U16692 (N_16692,N_10154,N_7438);
nor U16693 (N_16693,N_7280,N_12383);
or U16694 (N_16694,N_7646,N_12446);
or U16695 (N_16695,N_8150,N_12387);
xor U16696 (N_16696,N_8792,N_11562);
nand U16697 (N_16697,N_11447,N_10294);
xor U16698 (N_16698,N_11893,N_6355);
xor U16699 (N_16699,N_9506,N_8406);
xor U16700 (N_16700,N_8939,N_9326);
or U16701 (N_16701,N_11787,N_10059);
or U16702 (N_16702,N_6454,N_7231);
nand U16703 (N_16703,N_12131,N_12356);
or U16704 (N_16704,N_7711,N_8816);
nor U16705 (N_16705,N_12081,N_6818);
xnor U16706 (N_16706,N_7108,N_6962);
nor U16707 (N_16707,N_12410,N_7594);
or U16708 (N_16708,N_8171,N_9397);
or U16709 (N_16709,N_7846,N_9409);
nor U16710 (N_16710,N_7740,N_7159);
nand U16711 (N_16711,N_6474,N_10880);
nor U16712 (N_16712,N_6713,N_11118);
or U16713 (N_16713,N_8208,N_6566);
xnor U16714 (N_16714,N_7741,N_8805);
xor U16715 (N_16715,N_12092,N_12094);
xnor U16716 (N_16716,N_10355,N_12382);
and U16717 (N_16717,N_10903,N_9080);
or U16718 (N_16718,N_9726,N_9632);
nor U16719 (N_16719,N_10181,N_9841);
or U16720 (N_16720,N_11975,N_9635);
and U16721 (N_16721,N_6458,N_8132);
nand U16722 (N_16722,N_8576,N_6981);
nand U16723 (N_16723,N_7333,N_10785);
and U16724 (N_16724,N_10686,N_9178);
nand U16725 (N_16725,N_7927,N_8572);
xnor U16726 (N_16726,N_6924,N_8183);
or U16727 (N_16727,N_6783,N_10878);
or U16728 (N_16728,N_8915,N_9988);
xor U16729 (N_16729,N_6832,N_7134);
xor U16730 (N_16730,N_10200,N_7338);
or U16731 (N_16731,N_9909,N_6284);
xor U16732 (N_16732,N_12240,N_9543);
nor U16733 (N_16733,N_6279,N_6928);
nand U16734 (N_16734,N_8578,N_8856);
and U16735 (N_16735,N_7849,N_10198);
nand U16736 (N_16736,N_11639,N_12375);
or U16737 (N_16737,N_7662,N_7778);
nor U16738 (N_16738,N_10387,N_9496);
or U16739 (N_16739,N_11905,N_7971);
or U16740 (N_16740,N_7610,N_11317);
nor U16741 (N_16741,N_10141,N_12181);
and U16742 (N_16742,N_6616,N_8305);
and U16743 (N_16743,N_9792,N_10047);
nor U16744 (N_16744,N_6487,N_7159);
nand U16745 (N_16745,N_7493,N_10798);
nor U16746 (N_16746,N_12477,N_7326);
xor U16747 (N_16747,N_11048,N_9002);
nand U16748 (N_16748,N_10603,N_9787);
nor U16749 (N_16749,N_7520,N_7387);
and U16750 (N_16750,N_6320,N_11129);
nor U16751 (N_16751,N_9144,N_9788);
and U16752 (N_16752,N_9803,N_6481);
nor U16753 (N_16753,N_9526,N_11297);
nand U16754 (N_16754,N_6439,N_6840);
nor U16755 (N_16755,N_9286,N_9230);
and U16756 (N_16756,N_11566,N_10746);
nor U16757 (N_16757,N_10659,N_7693);
and U16758 (N_16758,N_8603,N_9829);
xor U16759 (N_16759,N_11868,N_11003);
xnor U16760 (N_16760,N_11670,N_9931);
nand U16761 (N_16761,N_6435,N_8971);
nand U16762 (N_16762,N_11354,N_6687);
and U16763 (N_16763,N_6822,N_11152);
and U16764 (N_16764,N_9014,N_10885);
xor U16765 (N_16765,N_6699,N_6681);
or U16766 (N_16766,N_9101,N_11241);
and U16767 (N_16767,N_8734,N_6744);
and U16768 (N_16768,N_7219,N_12436);
and U16769 (N_16769,N_10045,N_9474);
or U16770 (N_16770,N_7971,N_6662);
xnor U16771 (N_16771,N_10336,N_12335);
nor U16772 (N_16772,N_7165,N_6307);
xor U16773 (N_16773,N_6720,N_10924);
nor U16774 (N_16774,N_11037,N_6884);
nand U16775 (N_16775,N_11014,N_8107);
or U16776 (N_16776,N_10073,N_8734);
xnor U16777 (N_16777,N_10332,N_11506);
or U16778 (N_16778,N_9961,N_6930);
xor U16779 (N_16779,N_10168,N_10860);
nand U16780 (N_16780,N_8741,N_11904);
or U16781 (N_16781,N_11431,N_10244);
nand U16782 (N_16782,N_9982,N_11881);
nor U16783 (N_16783,N_10724,N_11203);
xor U16784 (N_16784,N_7926,N_7295);
or U16785 (N_16785,N_11274,N_8954);
nor U16786 (N_16786,N_9838,N_10260);
and U16787 (N_16787,N_12164,N_8318);
nand U16788 (N_16788,N_12107,N_9002);
nor U16789 (N_16789,N_6881,N_7347);
nand U16790 (N_16790,N_10317,N_7234);
and U16791 (N_16791,N_10003,N_9818);
nand U16792 (N_16792,N_7517,N_11083);
or U16793 (N_16793,N_11749,N_8615);
xor U16794 (N_16794,N_8265,N_7463);
xnor U16795 (N_16795,N_10668,N_7869);
xnor U16796 (N_16796,N_12271,N_7501);
nand U16797 (N_16797,N_12224,N_9643);
nor U16798 (N_16798,N_10720,N_10304);
and U16799 (N_16799,N_8825,N_11599);
nand U16800 (N_16800,N_10206,N_8472);
nor U16801 (N_16801,N_7913,N_12423);
and U16802 (N_16802,N_10066,N_6546);
nand U16803 (N_16803,N_10340,N_12105);
or U16804 (N_16804,N_6305,N_11551);
nor U16805 (N_16805,N_11733,N_7261);
and U16806 (N_16806,N_10717,N_12257);
or U16807 (N_16807,N_7111,N_7848);
nor U16808 (N_16808,N_12163,N_11174);
nor U16809 (N_16809,N_11133,N_8362);
xnor U16810 (N_16810,N_9286,N_10736);
and U16811 (N_16811,N_10426,N_7473);
nor U16812 (N_16812,N_9971,N_8941);
and U16813 (N_16813,N_10699,N_12175);
nor U16814 (N_16814,N_7498,N_9458);
xnor U16815 (N_16815,N_6671,N_7108);
and U16816 (N_16816,N_6539,N_6956);
or U16817 (N_16817,N_7175,N_12061);
nor U16818 (N_16818,N_7363,N_7744);
or U16819 (N_16819,N_11782,N_12233);
nor U16820 (N_16820,N_8812,N_6903);
nor U16821 (N_16821,N_12463,N_6597);
or U16822 (N_16822,N_11497,N_9810);
nor U16823 (N_16823,N_8292,N_12484);
or U16824 (N_16824,N_10666,N_9592);
nor U16825 (N_16825,N_11814,N_12047);
and U16826 (N_16826,N_9904,N_8664);
nor U16827 (N_16827,N_9765,N_9931);
xnor U16828 (N_16828,N_8726,N_7964);
or U16829 (N_16829,N_11327,N_9968);
and U16830 (N_16830,N_9777,N_6732);
nor U16831 (N_16831,N_11097,N_7655);
and U16832 (N_16832,N_11673,N_7879);
nand U16833 (N_16833,N_8095,N_8178);
nor U16834 (N_16834,N_6911,N_8095);
or U16835 (N_16835,N_11503,N_8113);
nor U16836 (N_16836,N_9766,N_7686);
nand U16837 (N_16837,N_7104,N_12165);
or U16838 (N_16838,N_9569,N_10458);
nor U16839 (N_16839,N_9531,N_7680);
xor U16840 (N_16840,N_9031,N_11625);
xor U16841 (N_16841,N_10921,N_6857);
and U16842 (N_16842,N_9434,N_6289);
or U16843 (N_16843,N_9761,N_8499);
nand U16844 (N_16844,N_9584,N_11096);
xor U16845 (N_16845,N_8237,N_10817);
nor U16846 (N_16846,N_8480,N_9035);
nor U16847 (N_16847,N_11393,N_11679);
nor U16848 (N_16848,N_9026,N_9111);
xor U16849 (N_16849,N_10074,N_8145);
or U16850 (N_16850,N_12437,N_8282);
or U16851 (N_16851,N_11040,N_12162);
nand U16852 (N_16852,N_12254,N_8900);
and U16853 (N_16853,N_11832,N_8986);
nand U16854 (N_16854,N_7375,N_9287);
and U16855 (N_16855,N_12401,N_10477);
or U16856 (N_16856,N_7078,N_10171);
or U16857 (N_16857,N_12385,N_12240);
nand U16858 (N_16858,N_12445,N_9924);
nand U16859 (N_16859,N_8751,N_8130);
nor U16860 (N_16860,N_8497,N_7404);
and U16861 (N_16861,N_10928,N_9963);
or U16862 (N_16862,N_10750,N_7812);
and U16863 (N_16863,N_6415,N_9804);
nor U16864 (N_16864,N_11478,N_9488);
and U16865 (N_16865,N_12169,N_8108);
nor U16866 (N_16866,N_10343,N_6614);
or U16867 (N_16867,N_9741,N_6282);
or U16868 (N_16868,N_12483,N_6610);
nand U16869 (N_16869,N_9338,N_11944);
and U16870 (N_16870,N_11594,N_11092);
xnor U16871 (N_16871,N_8643,N_12326);
and U16872 (N_16872,N_10527,N_9263);
xnor U16873 (N_16873,N_8523,N_9668);
nor U16874 (N_16874,N_6673,N_10782);
nand U16875 (N_16875,N_11723,N_7334);
and U16876 (N_16876,N_10280,N_10639);
and U16877 (N_16877,N_6399,N_7762);
xor U16878 (N_16878,N_8419,N_11504);
nand U16879 (N_16879,N_8808,N_11619);
nand U16880 (N_16880,N_8876,N_8718);
or U16881 (N_16881,N_6607,N_10073);
nand U16882 (N_16882,N_9500,N_11464);
nand U16883 (N_16883,N_9497,N_6870);
and U16884 (N_16884,N_11049,N_6672);
nand U16885 (N_16885,N_8258,N_9596);
or U16886 (N_16886,N_6615,N_9826);
or U16887 (N_16887,N_11992,N_12197);
and U16888 (N_16888,N_11309,N_12262);
and U16889 (N_16889,N_9903,N_10422);
nand U16890 (N_16890,N_11293,N_9623);
nor U16891 (N_16891,N_11283,N_9185);
or U16892 (N_16892,N_11259,N_10932);
nand U16893 (N_16893,N_6597,N_6950);
and U16894 (N_16894,N_12341,N_8269);
nor U16895 (N_16895,N_8429,N_6852);
nand U16896 (N_16896,N_9186,N_11676);
nand U16897 (N_16897,N_11133,N_8952);
nor U16898 (N_16898,N_10266,N_10279);
xor U16899 (N_16899,N_9362,N_8286);
nand U16900 (N_16900,N_7314,N_7536);
nand U16901 (N_16901,N_10916,N_12422);
xor U16902 (N_16902,N_10426,N_8575);
and U16903 (N_16903,N_11344,N_8196);
xnor U16904 (N_16904,N_8872,N_6888);
nor U16905 (N_16905,N_6688,N_6811);
nand U16906 (N_16906,N_11817,N_8507);
xor U16907 (N_16907,N_12254,N_7584);
nor U16908 (N_16908,N_6840,N_6316);
or U16909 (N_16909,N_6369,N_9580);
nand U16910 (N_16910,N_6315,N_8000);
xnor U16911 (N_16911,N_10914,N_9341);
or U16912 (N_16912,N_9200,N_9793);
nand U16913 (N_16913,N_12206,N_12391);
xor U16914 (N_16914,N_8357,N_8861);
nand U16915 (N_16915,N_8777,N_7161);
or U16916 (N_16916,N_11513,N_7074);
nand U16917 (N_16917,N_6988,N_10781);
xnor U16918 (N_16918,N_11740,N_10174);
xor U16919 (N_16919,N_12470,N_10527);
xnor U16920 (N_16920,N_7361,N_9882);
or U16921 (N_16921,N_9129,N_8335);
and U16922 (N_16922,N_11884,N_8190);
and U16923 (N_16923,N_9307,N_9944);
or U16924 (N_16924,N_7282,N_9153);
xor U16925 (N_16925,N_7190,N_6874);
and U16926 (N_16926,N_11223,N_8535);
and U16927 (N_16927,N_12077,N_6380);
nor U16928 (N_16928,N_9298,N_9984);
and U16929 (N_16929,N_9855,N_10968);
nand U16930 (N_16930,N_10616,N_9985);
xnor U16931 (N_16931,N_8409,N_9270);
and U16932 (N_16932,N_11135,N_6282);
nor U16933 (N_16933,N_12356,N_7340);
nand U16934 (N_16934,N_8648,N_10129);
nand U16935 (N_16935,N_9896,N_8714);
xnor U16936 (N_16936,N_10636,N_9243);
nor U16937 (N_16937,N_8455,N_7382);
or U16938 (N_16938,N_6728,N_8741);
or U16939 (N_16939,N_7980,N_7630);
or U16940 (N_16940,N_10823,N_9388);
xnor U16941 (N_16941,N_8511,N_6477);
nor U16942 (N_16942,N_12124,N_8437);
and U16943 (N_16943,N_6776,N_12425);
or U16944 (N_16944,N_7535,N_9215);
nand U16945 (N_16945,N_11294,N_12182);
and U16946 (N_16946,N_9942,N_8467);
nor U16947 (N_16947,N_7179,N_8925);
xnor U16948 (N_16948,N_12142,N_10042);
and U16949 (N_16949,N_9695,N_9162);
nand U16950 (N_16950,N_7829,N_11568);
nor U16951 (N_16951,N_11387,N_6948);
xor U16952 (N_16952,N_8377,N_7943);
and U16953 (N_16953,N_6404,N_7827);
and U16954 (N_16954,N_7622,N_11410);
nor U16955 (N_16955,N_12256,N_10031);
nand U16956 (N_16956,N_10739,N_8698);
nand U16957 (N_16957,N_6490,N_7002);
nor U16958 (N_16958,N_8904,N_10493);
or U16959 (N_16959,N_11091,N_9449);
and U16960 (N_16960,N_9089,N_11725);
nor U16961 (N_16961,N_10552,N_10789);
nand U16962 (N_16962,N_8302,N_12494);
nand U16963 (N_16963,N_7937,N_7074);
nand U16964 (N_16964,N_10471,N_12010);
nor U16965 (N_16965,N_7962,N_11468);
nor U16966 (N_16966,N_10090,N_10537);
nor U16967 (N_16967,N_11346,N_7669);
or U16968 (N_16968,N_11370,N_9015);
nor U16969 (N_16969,N_7129,N_6955);
nand U16970 (N_16970,N_11655,N_12202);
xnor U16971 (N_16971,N_8967,N_9871);
or U16972 (N_16972,N_8000,N_10041);
nand U16973 (N_16973,N_10236,N_11002);
nand U16974 (N_16974,N_7071,N_10372);
or U16975 (N_16975,N_8795,N_9582);
nand U16976 (N_16976,N_6599,N_10480);
or U16977 (N_16977,N_6277,N_6525);
nand U16978 (N_16978,N_11635,N_9114);
nand U16979 (N_16979,N_8510,N_7591);
nor U16980 (N_16980,N_8810,N_7211);
nor U16981 (N_16981,N_10387,N_10267);
and U16982 (N_16982,N_12050,N_10602);
nand U16983 (N_16983,N_12434,N_6466);
xnor U16984 (N_16984,N_10442,N_8173);
xnor U16985 (N_16985,N_8399,N_12144);
nand U16986 (N_16986,N_6876,N_9352);
or U16987 (N_16987,N_7932,N_6401);
nand U16988 (N_16988,N_10102,N_11368);
or U16989 (N_16989,N_9892,N_12464);
xor U16990 (N_16990,N_12477,N_7162);
xnor U16991 (N_16991,N_11484,N_11253);
nand U16992 (N_16992,N_8545,N_10698);
and U16993 (N_16993,N_7026,N_7758);
xor U16994 (N_16994,N_8135,N_8457);
nand U16995 (N_16995,N_11424,N_9130);
and U16996 (N_16996,N_8794,N_8446);
or U16997 (N_16997,N_8380,N_9532);
and U16998 (N_16998,N_8142,N_10076);
and U16999 (N_16999,N_11298,N_9933);
and U17000 (N_17000,N_9919,N_11880);
nand U17001 (N_17001,N_7331,N_10506);
nor U17002 (N_17002,N_11372,N_8330);
nand U17003 (N_17003,N_10608,N_11501);
nand U17004 (N_17004,N_11833,N_10549);
nor U17005 (N_17005,N_8268,N_7503);
or U17006 (N_17006,N_8606,N_8165);
xnor U17007 (N_17007,N_7235,N_8463);
nand U17008 (N_17008,N_6252,N_7911);
nand U17009 (N_17009,N_11045,N_12310);
and U17010 (N_17010,N_9571,N_11391);
xor U17011 (N_17011,N_7985,N_11385);
nand U17012 (N_17012,N_7149,N_11852);
and U17013 (N_17013,N_11874,N_6972);
nand U17014 (N_17014,N_7035,N_11846);
nand U17015 (N_17015,N_11114,N_7497);
and U17016 (N_17016,N_11958,N_10829);
nand U17017 (N_17017,N_10657,N_11671);
or U17018 (N_17018,N_9256,N_12192);
and U17019 (N_17019,N_12247,N_6474);
nor U17020 (N_17020,N_10273,N_8417);
or U17021 (N_17021,N_11636,N_12174);
nor U17022 (N_17022,N_8625,N_9590);
xor U17023 (N_17023,N_11983,N_11401);
and U17024 (N_17024,N_7541,N_9275);
nor U17025 (N_17025,N_8209,N_7713);
xnor U17026 (N_17026,N_8136,N_8522);
or U17027 (N_17027,N_7689,N_9353);
nor U17028 (N_17028,N_7779,N_7585);
xnor U17029 (N_17029,N_7898,N_10774);
and U17030 (N_17030,N_12407,N_11629);
nand U17031 (N_17031,N_11741,N_12267);
xnor U17032 (N_17032,N_6381,N_9834);
and U17033 (N_17033,N_7886,N_11503);
or U17034 (N_17034,N_8756,N_12194);
xnor U17035 (N_17035,N_8602,N_11858);
nor U17036 (N_17036,N_11576,N_12001);
nor U17037 (N_17037,N_6718,N_8795);
or U17038 (N_17038,N_9442,N_6409);
nand U17039 (N_17039,N_6888,N_11427);
xnor U17040 (N_17040,N_7040,N_11048);
and U17041 (N_17041,N_10015,N_8064);
xnor U17042 (N_17042,N_10852,N_11041);
nand U17043 (N_17043,N_11144,N_10866);
or U17044 (N_17044,N_8133,N_11697);
xnor U17045 (N_17045,N_8943,N_6565);
and U17046 (N_17046,N_11211,N_7319);
or U17047 (N_17047,N_10014,N_12132);
or U17048 (N_17048,N_6811,N_8134);
nand U17049 (N_17049,N_6350,N_12400);
or U17050 (N_17050,N_11813,N_8339);
nor U17051 (N_17051,N_11092,N_7725);
nor U17052 (N_17052,N_7377,N_7626);
and U17053 (N_17053,N_8572,N_10636);
or U17054 (N_17054,N_10678,N_11049);
nand U17055 (N_17055,N_9971,N_6567);
nor U17056 (N_17056,N_8621,N_10715);
or U17057 (N_17057,N_7269,N_8398);
nand U17058 (N_17058,N_11073,N_10090);
nor U17059 (N_17059,N_10931,N_6330);
nor U17060 (N_17060,N_6300,N_8233);
nor U17061 (N_17061,N_8763,N_8618);
and U17062 (N_17062,N_8610,N_9568);
xnor U17063 (N_17063,N_9266,N_11891);
xor U17064 (N_17064,N_10042,N_7606);
nand U17065 (N_17065,N_7336,N_12306);
or U17066 (N_17066,N_10339,N_7281);
or U17067 (N_17067,N_11656,N_7415);
and U17068 (N_17068,N_11400,N_9665);
or U17069 (N_17069,N_10626,N_6528);
nor U17070 (N_17070,N_8451,N_9410);
nor U17071 (N_17071,N_10057,N_9513);
nor U17072 (N_17072,N_10981,N_10826);
or U17073 (N_17073,N_6721,N_6464);
and U17074 (N_17074,N_8561,N_10745);
nor U17075 (N_17075,N_12352,N_6567);
nand U17076 (N_17076,N_10860,N_8287);
nand U17077 (N_17077,N_7338,N_11502);
or U17078 (N_17078,N_10353,N_8087);
nand U17079 (N_17079,N_9193,N_8850);
and U17080 (N_17080,N_11115,N_9558);
xor U17081 (N_17081,N_8847,N_8883);
nor U17082 (N_17082,N_6430,N_11978);
or U17083 (N_17083,N_9952,N_9538);
xnor U17084 (N_17084,N_8592,N_8133);
or U17085 (N_17085,N_8486,N_10689);
and U17086 (N_17086,N_12019,N_8791);
nand U17087 (N_17087,N_10036,N_8097);
xnor U17088 (N_17088,N_6870,N_6493);
nand U17089 (N_17089,N_8937,N_10117);
nor U17090 (N_17090,N_11025,N_8036);
and U17091 (N_17091,N_6545,N_9314);
nor U17092 (N_17092,N_11474,N_11206);
nand U17093 (N_17093,N_9133,N_11855);
xnor U17094 (N_17094,N_7172,N_8505);
nand U17095 (N_17095,N_7502,N_11326);
nor U17096 (N_17096,N_9601,N_11989);
and U17097 (N_17097,N_7998,N_10503);
xnor U17098 (N_17098,N_10420,N_9906);
xnor U17099 (N_17099,N_7963,N_12001);
nor U17100 (N_17100,N_8181,N_8812);
nand U17101 (N_17101,N_7132,N_7124);
and U17102 (N_17102,N_9514,N_11382);
xnor U17103 (N_17103,N_6409,N_10746);
xor U17104 (N_17104,N_8200,N_11415);
and U17105 (N_17105,N_7059,N_9551);
xor U17106 (N_17106,N_8946,N_6953);
or U17107 (N_17107,N_6994,N_7616);
nor U17108 (N_17108,N_9049,N_6519);
or U17109 (N_17109,N_7083,N_11452);
xnor U17110 (N_17110,N_8435,N_9125);
nand U17111 (N_17111,N_9772,N_7562);
nor U17112 (N_17112,N_10088,N_10740);
or U17113 (N_17113,N_10587,N_8424);
nand U17114 (N_17114,N_7639,N_11168);
and U17115 (N_17115,N_6867,N_7737);
nand U17116 (N_17116,N_6261,N_9026);
nand U17117 (N_17117,N_6877,N_11309);
or U17118 (N_17118,N_11057,N_11297);
xor U17119 (N_17119,N_10133,N_6789);
xor U17120 (N_17120,N_9888,N_7787);
or U17121 (N_17121,N_6811,N_9431);
nor U17122 (N_17122,N_6539,N_8463);
xnor U17123 (N_17123,N_6651,N_9852);
xnor U17124 (N_17124,N_6443,N_10438);
or U17125 (N_17125,N_6462,N_9870);
or U17126 (N_17126,N_7991,N_11862);
or U17127 (N_17127,N_11563,N_8670);
and U17128 (N_17128,N_8657,N_7261);
and U17129 (N_17129,N_8510,N_8172);
nor U17130 (N_17130,N_11968,N_11920);
nand U17131 (N_17131,N_11000,N_12458);
nand U17132 (N_17132,N_12080,N_8951);
nand U17133 (N_17133,N_10185,N_8565);
nor U17134 (N_17134,N_9069,N_10809);
nand U17135 (N_17135,N_10295,N_9383);
nor U17136 (N_17136,N_7169,N_10176);
xnor U17137 (N_17137,N_7300,N_8974);
nor U17138 (N_17138,N_8928,N_6293);
xor U17139 (N_17139,N_9841,N_8323);
nor U17140 (N_17140,N_6333,N_8231);
and U17141 (N_17141,N_7867,N_6410);
and U17142 (N_17142,N_7025,N_11444);
or U17143 (N_17143,N_7631,N_7338);
nand U17144 (N_17144,N_7895,N_6985);
or U17145 (N_17145,N_12335,N_11986);
or U17146 (N_17146,N_11964,N_6478);
or U17147 (N_17147,N_8179,N_11177);
or U17148 (N_17148,N_7028,N_10254);
or U17149 (N_17149,N_10609,N_12345);
and U17150 (N_17150,N_11776,N_8029);
xor U17151 (N_17151,N_6289,N_6344);
nor U17152 (N_17152,N_11847,N_8446);
nor U17153 (N_17153,N_6544,N_8840);
and U17154 (N_17154,N_7710,N_8741);
nor U17155 (N_17155,N_9208,N_9825);
nor U17156 (N_17156,N_7129,N_11783);
nor U17157 (N_17157,N_7783,N_7543);
nor U17158 (N_17158,N_9960,N_8700);
nand U17159 (N_17159,N_9934,N_8254);
or U17160 (N_17160,N_6499,N_8347);
and U17161 (N_17161,N_11615,N_8549);
nand U17162 (N_17162,N_10841,N_6531);
or U17163 (N_17163,N_7480,N_10157);
or U17164 (N_17164,N_7828,N_7032);
xor U17165 (N_17165,N_6873,N_8554);
nor U17166 (N_17166,N_7571,N_11602);
nand U17167 (N_17167,N_6371,N_11298);
nor U17168 (N_17168,N_12041,N_9681);
nor U17169 (N_17169,N_12232,N_9937);
xor U17170 (N_17170,N_7695,N_9409);
xnor U17171 (N_17171,N_11585,N_8942);
nor U17172 (N_17172,N_8283,N_6504);
xor U17173 (N_17173,N_6542,N_10249);
nand U17174 (N_17174,N_10528,N_12033);
nand U17175 (N_17175,N_9962,N_6896);
and U17176 (N_17176,N_12380,N_10690);
or U17177 (N_17177,N_11092,N_12166);
nand U17178 (N_17178,N_6326,N_6959);
and U17179 (N_17179,N_10930,N_11436);
or U17180 (N_17180,N_9325,N_9631);
or U17181 (N_17181,N_8134,N_9598);
nor U17182 (N_17182,N_8545,N_8517);
and U17183 (N_17183,N_7205,N_7344);
nor U17184 (N_17184,N_11093,N_7571);
nor U17185 (N_17185,N_8947,N_8320);
and U17186 (N_17186,N_7507,N_8338);
nand U17187 (N_17187,N_9972,N_9326);
nand U17188 (N_17188,N_8246,N_8243);
and U17189 (N_17189,N_10926,N_11167);
nor U17190 (N_17190,N_10526,N_10195);
nand U17191 (N_17191,N_9854,N_7896);
or U17192 (N_17192,N_8837,N_11003);
or U17193 (N_17193,N_11947,N_10915);
xor U17194 (N_17194,N_7783,N_11265);
nand U17195 (N_17195,N_6859,N_9427);
and U17196 (N_17196,N_6968,N_7864);
xor U17197 (N_17197,N_8234,N_11548);
or U17198 (N_17198,N_10059,N_8176);
and U17199 (N_17199,N_12080,N_8605);
and U17200 (N_17200,N_11246,N_7656);
nor U17201 (N_17201,N_10198,N_10716);
or U17202 (N_17202,N_11186,N_9803);
xor U17203 (N_17203,N_9301,N_7464);
xor U17204 (N_17204,N_9374,N_9857);
and U17205 (N_17205,N_8665,N_9185);
and U17206 (N_17206,N_10931,N_7582);
and U17207 (N_17207,N_8375,N_9284);
nor U17208 (N_17208,N_8614,N_9891);
nand U17209 (N_17209,N_7618,N_11060);
nand U17210 (N_17210,N_9828,N_10445);
nand U17211 (N_17211,N_8956,N_9103);
and U17212 (N_17212,N_7669,N_10737);
nor U17213 (N_17213,N_10548,N_11521);
and U17214 (N_17214,N_10363,N_8943);
or U17215 (N_17215,N_9101,N_6364);
or U17216 (N_17216,N_7792,N_10333);
and U17217 (N_17217,N_11581,N_10845);
and U17218 (N_17218,N_6740,N_12303);
xor U17219 (N_17219,N_9841,N_7443);
nor U17220 (N_17220,N_11605,N_8402);
or U17221 (N_17221,N_10600,N_9406);
nand U17222 (N_17222,N_7617,N_8933);
xnor U17223 (N_17223,N_8434,N_10441);
or U17224 (N_17224,N_11386,N_9841);
nor U17225 (N_17225,N_7063,N_7569);
or U17226 (N_17226,N_11328,N_11594);
or U17227 (N_17227,N_10403,N_11710);
nor U17228 (N_17228,N_10761,N_7451);
or U17229 (N_17229,N_9407,N_9851);
and U17230 (N_17230,N_12334,N_8930);
or U17231 (N_17231,N_8293,N_7371);
and U17232 (N_17232,N_8758,N_9919);
xor U17233 (N_17233,N_9438,N_11757);
or U17234 (N_17234,N_6926,N_7792);
nor U17235 (N_17235,N_8280,N_7466);
nor U17236 (N_17236,N_12250,N_9934);
nor U17237 (N_17237,N_6288,N_8827);
or U17238 (N_17238,N_7665,N_11119);
nor U17239 (N_17239,N_11341,N_10854);
nor U17240 (N_17240,N_9365,N_6289);
and U17241 (N_17241,N_7384,N_9452);
xnor U17242 (N_17242,N_7359,N_12489);
and U17243 (N_17243,N_8449,N_9752);
or U17244 (N_17244,N_7454,N_8485);
and U17245 (N_17245,N_9962,N_11576);
nor U17246 (N_17246,N_7870,N_11916);
nor U17247 (N_17247,N_8569,N_7569);
or U17248 (N_17248,N_9117,N_11158);
nor U17249 (N_17249,N_7101,N_9919);
nor U17250 (N_17250,N_9131,N_8795);
nor U17251 (N_17251,N_7451,N_6968);
nor U17252 (N_17252,N_6935,N_9235);
nand U17253 (N_17253,N_9657,N_10742);
nor U17254 (N_17254,N_10700,N_9166);
nor U17255 (N_17255,N_8767,N_6767);
and U17256 (N_17256,N_7013,N_12453);
nor U17257 (N_17257,N_11086,N_8997);
or U17258 (N_17258,N_9182,N_11486);
or U17259 (N_17259,N_8385,N_8885);
xnor U17260 (N_17260,N_8464,N_9574);
and U17261 (N_17261,N_11473,N_7289);
nor U17262 (N_17262,N_9409,N_11607);
xor U17263 (N_17263,N_10376,N_7349);
xor U17264 (N_17264,N_9951,N_6636);
xor U17265 (N_17265,N_10637,N_11245);
nor U17266 (N_17266,N_6763,N_11793);
nand U17267 (N_17267,N_7710,N_8533);
and U17268 (N_17268,N_6451,N_6355);
nor U17269 (N_17269,N_8785,N_6867);
and U17270 (N_17270,N_11279,N_8598);
nand U17271 (N_17271,N_10389,N_11893);
xor U17272 (N_17272,N_12454,N_11477);
nand U17273 (N_17273,N_10859,N_11968);
nand U17274 (N_17274,N_7201,N_10963);
xor U17275 (N_17275,N_12452,N_9195);
xnor U17276 (N_17276,N_10716,N_11441);
xor U17277 (N_17277,N_8052,N_10387);
or U17278 (N_17278,N_7675,N_9303);
and U17279 (N_17279,N_6436,N_10613);
nand U17280 (N_17280,N_11193,N_8519);
nand U17281 (N_17281,N_10782,N_8154);
xnor U17282 (N_17282,N_6654,N_8891);
nor U17283 (N_17283,N_11771,N_9094);
or U17284 (N_17284,N_9049,N_8988);
xnor U17285 (N_17285,N_9172,N_10837);
nor U17286 (N_17286,N_8366,N_8124);
xnor U17287 (N_17287,N_8478,N_8783);
nand U17288 (N_17288,N_10257,N_9886);
xor U17289 (N_17289,N_8718,N_7771);
nand U17290 (N_17290,N_8736,N_8633);
and U17291 (N_17291,N_11961,N_7463);
and U17292 (N_17292,N_11125,N_12355);
xnor U17293 (N_17293,N_7295,N_10016);
xor U17294 (N_17294,N_6797,N_6841);
and U17295 (N_17295,N_11538,N_12325);
nand U17296 (N_17296,N_6432,N_10842);
or U17297 (N_17297,N_7027,N_10656);
or U17298 (N_17298,N_7043,N_10409);
or U17299 (N_17299,N_10239,N_10338);
and U17300 (N_17300,N_7781,N_11418);
nor U17301 (N_17301,N_7662,N_8297);
and U17302 (N_17302,N_8279,N_8644);
nor U17303 (N_17303,N_12225,N_8257);
nor U17304 (N_17304,N_7615,N_11835);
or U17305 (N_17305,N_8366,N_11171);
nand U17306 (N_17306,N_10670,N_6479);
nor U17307 (N_17307,N_7500,N_6789);
and U17308 (N_17308,N_8248,N_6403);
or U17309 (N_17309,N_6387,N_11714);
and U17310 (N_17310,N_9181,N_9282);
and U17311 (N_17311,N_6371,N_12181);
nor U17312 (N_17312,N_9578,N_9023);
nand U17313 (N_17313,N_11290,N_10673);
nor U17314 (N_17314,N_6748,N_7884);
and U17315 (N_17315,N_12083,N_8288);
nor U17316 (N_17316,N_9014,N_9715);
xor U17317 (N_17317,N_11592,N_7152);
nand U17318 (N_17318,N_6388,N_11532);
and U17319 (N_17319,N_11707,N_11753);
nor U17320 (N_17320,N_9875,N_9953);
and U17321 (N_17321,N_8655,N_11067);
and U17322 (N_17322,N_8818,N_11542);
nor U17323 (N_17323,N_9931,N_8833);
nand U17324 (N_17324,N_7164,N_8127);
or U17325 (N_17325,N_7060,N_12235);
and U17326 (N_17326,N_8253,N_10139);
xnor U17327 (N_17327,N_12426,N_9840);
and U17328 (N_17328,N_7051,N_8070);
nand U17329 (N_17329,N_9361,N_6587);
or U17330 (N_17330,N_11483,N_6378);
and U17331 (N_17331,N_11309,N_7138);
nand U17332 (N_17332,N_10192,N_9872);
nand U17333 (N_17333,N_10431,N_11772);
or U17334 (N_17334,N_7669,N_9606);
or U17335 (N_17335,N_7414,N_7568);
and U17336 (N_17336,N_10203,N_12484);
xnor U17337 (N_17337,N_9366,N_12188);
nor U17338 (N_17338,N_9968,N_10200);
xnor U17339 (N_17339,N_11824,N_10975);
nor U17340 (N_17340,N_6647,N_9620);
xor U17341 (N_17341,N_7224,N_9373);
or U17342 (N_17342,N_11007,N_12356);
or U17343 (N_17343,N_11501,N_12301);
xnor U17344 (N_17344,N_9468,N_11473);
and U17345 (N_17345,N_7342,N_11273);
nand U17346 (N_17346,N_8361,N_10854);
and U17347 (N_17347,N_9495,N_9221);
nand U17348 (N_17348,N_11985,N_10494);
nand U17349 (N_17349,N_10771,N_11463);
nand U17350 (N_17350,N_12005,N_11575);
nand U17351 (N_17351,N_12001,N_11957);
and U17352 (N_17352,N_6471,N_9006);
or U17353 (N_17353,N_10005,N_9163);
xnor U17354 (N_17354,N_8170,N_9058);
nand U17355 (N_17355,N_8263,N_10724);
nor U17356 (N_17356,N_6699,N_11494);
xnor U17357 (N_17357,N_6342,N_8651);
nand U17358 (N_17358,N_7379,N_10185);
and U17359 (N_17359,N_10553,N_7848);
or U17360 (N_17360,N_6302,N_10183);
or U17361 (N_17361,N_9469,N_10542);
xnor U17362 (N_17362,N_6952,N_6708);
nor U17363 (N_17363,N_8238,N_8312);
xnor U17364 (N_17364,N_6960,N_11914);
and U17365 (N_17365,N_10838,N_9692);
nand U17366 (N_17366,N_9526,N_9306);
or U17367 (N_17367,N_10800,N_12103);
and U17368 (N_17368,N_10783,N_8131);
or U17369 (N_17369,N_8828,N_12152);
xor U17370 (N_17370,N_11693,N_6803);
and U17371 (N_17371,N_11838,N_10042);
nand U17372 (N_17372,N_7071,N_8313);
nand U17373 (N_17373,N_8003,N_7076);
and U17374 (N_17374,N_12357,N_9347);
xor U17375 (N_17375,N_12198,N_11638);
xor U17376 (N_17376,N_9217,N_8009);
and U17377 (N_17377,N_9701,N_7495);
nor U17378 (N_17378,N_7862,N_8198);
or U17379 (N_17379,N_8980,N_9337);
and U17380 (N_17380,N_8590,N_9204);
nor U17381 (N_17381,N_6292,N_7616);
nand U17382 (N_17382,N_8761,N_12076);
nor U17383 (N_17383,N_7226,N_7821);
or U17384 (N_17384,N_9772,N_8693);
xor U17385 (N_17385,N_10397,N_11950);
or U17386 (N_17386,N_10390,N_12276);
nand U17387 (N_17387,N_8553,N_8467);
and U17388 (N_17388,N_8975,N_6637);
nand U17389 (N_17389,N_6686,N_9744);
or U17390 (N_17390,N_11850,N_6474);
nand U17391 (N_17391,N_11716,N_7202);
or U17392 (N_17392,N_10465,N_10130);
xor U17393 (N_17393,N_6988,N_6471);
and U17394 (N_17394,N_11988,N_12297);
nor U17395 (N_17395,N_10242,N_9317);
or U17396 (N_17396,N_8532,N_11389);
or U17397 (N_17397,N_7860,N_10278);
and U17398 (N_17398,N_7209,N_6761);
xnor U17399 (N_17399,N_11046,N_8686);
nand U17400 (N_17400,N_6750,N_11398);
or U17401 (N_17401,N_9082,N_7056);
nor U17402 (N_17402,N_8382,N_8999);
nand U17403 (N_17403,N_6977,N_7257);
xor U17404 (N_17404,N_6589,N_9296);
nand U17405 (N_17405,N_10481,N_10488);
xnor U17406 (N_17406,N_12094,N_10505);
and U17407 (N_17407,N_12237,N_6742);
and U17408 (N_17408,N_9527,N_10132);
and U17409 (N_17409,N_8466,N_8655);
xor U17410 (N_17410,N_10534,N_9082);
and U17411 (N_17411,N_6586,N_9440);
or U17412 (N_17412,N_7848,N_8048);
nand U17413 (N_17413,N_8990,N_12020);
nor U17414 (N_17414,N_10272,N_12011);
or U17415 (N_17415,N_9809,N_12400);
nor U17416 (N_17416,N_9526,N_8939);
and U17417 (N_17417,N_10528,N_10232);
and U17418 (N_17418,N_11990,N_6305);
nor U17419 (N_17419,N_10204,N_7950);
nand U17420 (N_17420,N_12194,N_12293);
xor U17421 (N_17421,N_6380,N_11304);
nor U17422 (N_17422,N_10655,N_8725);
nand U17423 (N_17423,N_8685,N_6603);
and U17424 (N_17424,N_7881,N_11708);
nand U17425 (N_17425,N_8733,N_9708);
and U17426 (N_17426,N_8378,N_6659);
xnor U17427 (N_17427,N_11947,N_9651);
nor U17428 (N_17428,N_9786,N_7306);
or U17429 (N_17429,N_9376,N_11384);
xor U17430 (N_17430,N_7701,N_10927);
xor U17431 (N_17431,N_7054,N_10951);
or U17432 (N_17432,N_11548,N_6565);
xor U17433 (N_17433,N_9420,N_6518);
nor U17434 (N_17434,N_7991,N_10238);
and U17435 (N_17435,N_7976,N_8758);
nor U17436 (N_17436,N_8652,N_6538);
xor U17437 (N_17437,N_11416,N_8290);
nand U17438 (N_17438,N_11386,N_7589);
xnor U17439 (N_17439,N_11596,N_8541);
nand U17440 (N_17440,N_9824,N_6547);
xor U17441 (N_17441,N_8447,N_11045);
nor U17442 (N_17442,N_7974,N_8679);
or U17443 (N_17443,N_6979,N_12468);
xnor U17444 (N_17444,N_9948,N_8453);
and U17445 (N_17445,N_7835,N_8049);
xor U17446 (N_17446,N_7624,N_12431);
xor U17447 (N_17447,N_11111,N_9535);
or U17448 (N_17448,N_11498,N_12043);
nand U17449 (N_17449,N_9148,N_10059);
nand U17450 (N_17450,N_10439,N_9923);
or U17451 (N_17451,N_8255,N_7737);
and U17452 (N_17452,N_7953,N_6383);
and U17453 (N_17453,N_7112,N_11553);
and U17454 (N_17454,N_11122,N_9535);
xor U17455 (N_17455,N_11131,N_9265);
or U17456 (N_17456,N_10847,N_7850);
nor U17457 (N_17457,N_8481,N_10772);
nor U17458 (N_17458,N_11104,N_12405);
xor U17459 (N_17459,N_10798,N_10904);
xor U17460 (N_17460,N_10554,N_12166);
nor U17461 (N_17461,N_11664,N_11662);
xor U17462 (N_17462,N_11526,N_7262);
nand U17463 (N_17463,N_6947,N_6436);
and U17464 (N_17464,N_12060,N_7047);
nor U17465 (N_17465,N_10051,N_9761);
xor U17466 (N_17466,N_7504,N_10978);
xnor U17467 (N_17467,N_9968,N_9258);
and U17468 (N_17468,N_9105,N_9796);
nor U17469 (N_17469,N_7124,N_9321);
and U17470 (N_17470,N_10250,N_7275);
nand U17471 (N_17471,N_7643,N_12003);
or U17472 (N_17472,N_10004,N_8037);
and U17473 (N_17473,N_9377,N_9398);
nor U17474 (N_17474,N_10574,N_7674);
or U17475 (N_17475,N_9605,N_11364);
nor U17476 (N_17476,N_8623,N_9126);
nand U17477 (N_17477,N_11910,N_11468);
xnor U17478 (N_17478,N_11250,N_10636);
xor U17479 (N_17479,N_7939,N_12388);
and U17480 (N_17480,N_10313,N_11275);
nor U17481 (N_17481,N_6934,N_11646);
xor U17482 (N_17482,N_8293,N_7351);
and U17483 (N_17483,N_7608,N_7959);
nand U17484 (N_17484,N_10911,N_7937);
nor U17485 (N_17485,N_8805,N_8398);
and U17486 (N_17486,N_6643,N_6688);
nand U17487 (N_17487,N_11573,N_6805);
xor U17488 (N_17488,N_11201,N_8474);
and U17489 (N_17489,N_8711,N_9474);
nor U17490 (N_17490,N_12135,N_6455);
or U17491 (N_17491,N_8560,N_9559);
and U17492 (N_17492,N_6725,N_10714);
and U17493 (N_17493,N_12066,N_9055);
or U17494 (N_17494,N_6842,N_11962);
and U17495 (N_17495,N_7471,N_10012);
nand U17496 (N_17496,N_8837,N_9150);
and U17497 (N_17497,N_10367,N_8297);
and U17498 (N_17498,N_11736,N_6481);
nand U17499 (N_17499,N_7160,N_11992);
and U17500 (N_17500,N_11809,N_10225);
nand U17501 (N_17501,N_7528,N_10927);
nand U17502 (N_17502,N_7736,N_11216);
nor U17503 (N_17503,N_11452,N_8245);
and U17504 (N_17504,N_11640,N_9933);
nand U17505 (N_17505,N_10152,N_10857);
xnor U17506 (N_17506,N_6402,N_7174);
nor U17507 (N_17507,N_8031,N_12045);
xnor U17508 (N_17508,N_11185,N_10611);
nor U17509 (N_17509,N_9321,N_7890);
or U17510 (N_17510,N_9990,N_7490);
nand U17511 (N_17511,N_6942,N_10564);
xnor U17512 (N_17512,N_7996,N_7538);
nand U17513 (N_17513,N_11529,N_6967);
and U17514 (N_17514,N_8346,N_11185);
xnor U17515 (N_17515,N_6645,N_6363);
xor U17516 (N_17516,N_6554,N_6360);
xor U17517 (N_17517,N_10251,N_6726);
nor U17518 (N_17518,N_7923,N_11229);
and U17519 (N_17519,N_11400,N_7831);
nor U17520 (N_17520,N_10634,N_11335);
xnor U17521 (N_17521,N_12441,N_10444);
nor U17522 (N_17522,N_11220,N_7908);
and U17523 (N_17523,N_9217,N_10101);
nand U17524 (N_17524,N_6737,N_7086);
nor U17525 (N_17525,N_11716,N_6566);
nor U17526 (N_17526,N_8806,N_12010);
nand U17527 (N_17527,N_11747,N_10889);
xor U17528 (N_17528,N_12126,N_7093);
or U17529 (N_17529,N_8713,N_11655);
and U17530 (N_17530,N_10496,N_7875);
nand U17531 (N_17531,N_7174,N_10156);
xor U17532 (N_17532,N_9990,N_7096);
nand U17533 (N_17533,N_10838,N_7059);
xor U17534 (N_17534,N_7548,N_10117);
xor U17535 (N_17535,N_7588,N_6306);
and U17536 (N_17536,N_11961,N_8085);
or U17537 (N_17537,N_10992,N_7048);
and U17538 (N_17538,N_7981,N_12407);
and U17539 (N_17539,N_9853,N_11896);
and U17540 (N_17540,N_6831,N_9660);
nand U17541 (N_17541,N_7683,N_10938);
or U17542 (N_17542,N_7458,N_8748);
nand U17543 (N_17543,N_10835,N_8185);
nand U17544 (N_17544,N_11611,N_10391);
nand U17545 (N_17545,N_6279,N_7004);
or U17546 (N_17546,N_9445,N_7977);
or U17547 (N_17547,N_9092,N_8609);
xnor U17548 (N_17548,N_9000,N_10471);
nor U17549 (N_17549,N_11326,N_6610);
and U17550 (N_17550,N_8604,N_6427);
nand U17551 (N_17551,N_10835,N_11947);
xor U17552 (N_17552,N_9450,N_9405);
or U17553 (N_17553,N_6769,N_6522);
nor U17554 (N_17554,N_12113,N_12320);
or U17555 (N_17555,N_6791,N_11533);
xnor U17556 (N_17556,N_11547,N_10489);
nand U17557 (N_17557,N_12220,N_8838);
xor U17558 (N_17558,N_11906,N_10160);
xor U17559 (N_17559,N_7810,N_9301);
nor U17560 (N_17560,N_8616,N_6847);
nor U17561 (N_17561,N_6738,N_12228);
nand U17562 (N_17562,N_8740,N_11193);
and U17563 (N_17563,N_9719,N_11067);
nor U17564 (N_17564,N_9842,N_8371);
xor U17565 (N_17565,N_9054,N_10123);
nor U17566 (N_17566,N_8924,N_6442);
or U17567 (N_17567,N_7484,N_10153);
xor U17568 (N_17568,N_8210,N_10540);
xor U17569 (N_17569,N_11174,N_8939);
or U17570 (N_17570,N_12122,N_6350);
xnor U17571 (N_17571,N_10163,N_7782);
or U17572 (N_17572,N_9669,N_9038);
nand U17573 (N_17573,N_7302,N_8887);
nand U17574 (N_17574,N_11461,N_8803);
xor U17575 (N_17575,N_12197,N_7441);
and U17576 (N_17576,N_8122,N_7078);
or U17577 (N_17577,N_9806,N_9038);
nor U17578 (N_17578,N_10373,N_9726);
nand U17579 (N_17579,N_10146,N_10464);
or U17580 (N_17580,N_7742,N_12041);
nand U17581 (N_17581,N_9737,N_10164);
nand U17582 (N_17582,N_11019,N_7569);
xor U17583 (N_17583,N_7435,N_11015);
nand U17584 (N_17584,N_8067,N_6523);
nor U17585 (N_17585,N_7705,N_9820);
and U17586 (N_17586,N_8486,N_8098);
xnor U17587 (N_17587,N_8744,N_9587);
and U17588 (N_17588,N_11696,N_7361);
and U17589 (N_17589,N_7108,N_6284);
xor U17590 (N_17590,N_6627,N_6254);
nand U17591 (N_17591,N_6302,N_8060);
and U17592 (N_17592,N_11532,N_11014);
nor U17593 (N_17593,N_10715,N_9018);
nand U17594 (N_17594,N_9342,N_8174);
or U17595 (N_17595,N_10848,N_12226);
xnor U17596 (N_17596,N_12270,N_8905);
nor U17597 (N_17597,N_11582,N_7459);
nor U17598 (N_17598,N_8864,N_6620);
nand U17599 (N_17599,N_11830,N_6345);
xor U17600 (N_17600,N_10567,N_7138);
nand U17601 (N_17601,N_6404,N_10691);
nor U17602 (N_17602,N_9259,N_8464);
and U17603 (N_17603,N_10205,N_11642);
or U17604 (N_17604,N_11819,N_10868);
and U17605 (N_17605,N_10227,N_8404);
xnor U17606 (N_17606,N_8701,N_12397);
nand U17607 (N_17607,N_11842,N_12257);
xnor U17608 (N_17608,N_8945,N_12299);
nand U17609 (N_17609,N_8797,N_9351);
or U17610 (N_17610,N_11539,N_8827);
and U17611 (N_17611,N_8301,N_8289);
xnor U17612 (N_17612,N_7464,N_6904);
and U17613 (N_17613,N_6840,N_9441);
nand U17614 (N_17614,N_8489,N_7109);
or U17615 (N_17615,N_9858,N_11886);
and U17616 (N_17616,N_8777,N_9292);
nor U17617 (N_17617,N_8844,N_8568);
nand U17618 (N_17618,N_7462,N_7884);
nand U17619 (N_17619,N_10820,N_12333);
and U17620 (N_17620,N_11940,N_12444);
and U17621 (N_17621,N_9690,N_6433);
and U17622 (N_17622,N_12378,N_12202);
nor U17623 (N_17623,N_11011,N_11001);
nor U17624 (N_17624,N_8512,N_11714);
and U17625 (N_17625,N_10965,N_12331);
or U17626 (N_17626,N_7766,N_12039);
and U17627 (N_17627,N_7848,N_7706);
nand U17628 (N_17628,N_10035,N_10153);
or U17629 (N_17629,N_7430,N_12038);
and U17630 (N_17630,N_12463,N_9823);
nand U17631 (N_17631,N_10717,N_10460);
and U17632 (N_17632,N_8073,N_8686);
or U17633 (N_17633,N_8028,N_8965);
nor U17634 (N_17634,N_8267,N_10457);
nor U17635 (N_17635,N_6624,N_10167);
xor U17636 (N_17636,N_7837,N_9092);
or U17637 (N_17637,N_10055,N_6491);
nand U17638 (N_17638,N_10872,N_7856);
and U17639 (N_17639,N_10445,N_10898);
nand U17640 (N_17640,N_7325,N_7241);
or U17641 (N_17641,N_10271,N_11870);
nor U17642 (N_17642,N_11693,N_6936);
and U17643 (N_17643,N_10362,N_8297);
or U17644 (N_17644,N_7857,N_11695);
nand U17645 (N_17645,N_9248,N_8484);
and U17646 (N_17646,N_7574,N_9951);
nand U17647 (N_17647,N_11533,N_7643);
nor U17648 (N_17648,N_7365,N_11303);
xnor U17649 (N_17649,N_9137,N_10339);
xor U17650 (N_17650,N_10930,N_7774);
or U17651 (N_17651,N_9038,N_9999);
nand U17652 (N_17652,N_6981,N_6397);
and U17653 (N_17653,N_8244,N_7227);
and U17654 (N_17654,N_8376,N_11931);
nand U17655 (N_17655,N_9823,N_8389);
and U17656 (N_17656,N_7020,N_6270);
nor U17657 (N_17657,N_11376,N_8103);
nor U17658 (N_17658,N_6738,N_10689);
nand U17659 (N_17659,N_6763,N_11291);
or U17660 (N_17660,N_9883,N_9385);
nor U17661 (N_17661,N_10258,N_9838);
and U17662 (N_17662,N_7761,N_11728);
nor U17663 (N_17663,N_6660,N_11559);
nand U17664 (N_17664,N_9441,N_9578);
and U17665 (N_17665,N_6517,N_7606);
nand U17666 (N_17666,N_11443,N_10769);
xnor U17667 (N_17667,N_9292,N_11232);
and U17668 (N_17668,N_11818,N_11823);
xnor U17669 (N_17669,N_9482,N_7225);
or U17670 (N_17670,N_9540,N_7025);
xnor U17671 (N_17671,N_9659,N_10684);
nand U17672 (N_17672,N_10529,N_10567);
and U17673 (N_17673,N_9521,N_9921);
or U17674 (N_17674,N_7429,N_7246);
nand U17675 (N_17675,N_7696,N_8390);
xnor U17676 (N_17676,N_12061,N_10374);
and U17677 (N_17677,N_6302,N_11650);
nor U17678 (N_17678,N_7518,N_11364);
or U17679 (N_17679,N_7465,N_9701);
or U17680 (N_17680,N_7986,N_7349);
or U17681 (N_17681,N_8103,N_10503);
or U17682 (N_17682,N_8763,N_10176);
or U17683 (N_17683,N_9524,N_10299);
or U17684 (N_17684,N_11917,N_11656);
nor U17685 (N_17685,N_11608,N_6809);
xnor U17686 (N_17686,N_10515,N_9961);
xor U17687 (N_17687,N_7336,N_11820);
xor U17688 (N_17688,N_7519,N_11046);
and U17689 (N_17689,N_11854,N_8317);
or U17690 (N_17690,N_11274,N_8110);
nand U17691 (N_17691,N_8602,N_11176);
and U17692 (N_17692,N_9885,N_9573);
xor U17693 (N_17693,N_12048,N_8461);
nand U17694 (N_17694,N_10871,N_6455);
nand U17695 (N_17695,N_8863,N_12054);
nand U17696 (N_17696,N_11342,N_9631);
nor U17697 (N_17697,N_9546,N_6980);
nor U17698 (N_17698,N_8402,N_8919);
and U17699 (N_17699,N_9282,N_6913);
and U17700 (N_17700,N_7429,N_8304);
or U17701 (N_17701,N_11986,N_9330);
nand U17702 (N_17702,N_6304,N_10688);
or U17703 (N_17703,N_7782,N_10766);
or U17704 (N_17704,N_7201,N_9019);
and U17705 (N_17705,N_12252,N_8235);
and U17706 (N_17706,N_10080,N_7127);
xor U17707 (N_17707,N_11810,N_11240);
nor U17708 (N_17708,N_6647,N_10172);
or U17709 (N_17709,N_10731,N_7456);
xor U17710 (N_17710,N_6645,N_6304);
nor U17711 (N_17711,N_11418,N_10378);
nand U17712 (N_17712,N_10144,N_6288);
xor U17713 (N_17713,N_10101,N_7894);
nand U17714 (N_17714,N_9508,N_8444);
nand U17715 (N_17715,N_6925,N_10311);
nand U17716 (N_17716,N_11745,N_11788);
nand U17717 (N_17717,N_10977,N_8945);
nor U17718 (N_17718,N_6868,N_8588);
and U17719 (N_17719,N_7078,N_9771);
and U17720 (N_17720,N_6742,N_10081);
nor U17721 (N_17721,N_10787,N_10036);
and U17722 (N_17722,N_7478,N_6862);
or U17723 (N_17723,N_12329,N_10664);
nand U17724 (N_17724,N_8740,N_8996);
and U17725 (N_17725,N_8536,N_12036);
nand U17726 (N_17726,N_7059,N_9546);
and U17727 (N_17727,N_8219,N_6806);
nand U17728 (N_17728,N_6769,N_9287);
and U17729 (N_17729,N_8180,N_6482);
xor U17730 (N_17730,N_7803,N_9158);
or U17731 (N_17731,N_11931,N_7083);
nand U17732 (N_17732,N_7080,N_8743);
nand U17733 (N_17733,N_12270,N_7970);
nand U17734 (N_17734,N_11720,N_7462);
or U17735 (N_17735,N_9676,N_9720);
xor U17736 (N_17736,N_12033,N_11492);
nand U17737 (N_17737,N_12244,N_6384);
nand U17738 (N_17738,N_11650,N_11879);
nand U17739 (N_17739,N_8851,N_10897);
or U17740 (N_17740,N_12097,N_10311);
and U17741 (N_17741,N_9711,N_9809);
xor U17742 (N_17742,N_7193,N_10500);
nor U17743 (N_17743,N_8374,N_6874);
or U17744 (N_17744,N_8050,N_7487);
nand U17745 (N_17745,N_11283,N_10596);
xor U17746 (N_17746,N_11015,N_8565);
nand U17747 (N_17747,N_6282,N_10874);
xnor U17748 (N_17748,N_7347,N_9749);
or U17749 (N_17749,N_8630,N_10757);
xnor U17750 (N_17750,N_8533,N_8574);
nand U17751 (N_17751,N_10895,N_9648);
nand U17752 (N_17752,N_10657,N_11384);
nor U17753 (N_17753,N_7258,N_11682);
nor U17754 (N_17754,N_7074,N_10776);
or U17755 (N_17755,N_6640,N_8540);
nand U17756 (N_17756,N_9043,N_9009);
and U17757 (N_17757,N_11410,N_9955);
or U17758 (N_17758,N_9833,N_10601);
and U17759 (N_17759,N_9592,N_7504);
xor U17760 (N_17760,N_11356,N_9533);
xor U17761 (N_17761,N_8749,N_6362);
and U17762 (N_17762,N_9099,N_6714);
xor U17763 (N_17763,N_7033,N_7130);
and U17764 (N_17764,N_6644,N_11503);
nand U17765 (N_17765,N_10316,N_7944);
xnor U17766 (N_17766,N_9758,N_6334);
nand U17767 (N_17767,N_6575,N_7941);
nand U17768 (N_17768,N_8386,N_12160);
nand U17769 (N_17769,N_9675,N_11516);
and U17770 (N_17770,N_9839,N_9137);
nor U17771 (N_17771,N_12215,N_6285);
xor U17772 (N_17772,N_9466,N_6317);
and U17773 (N_17773,N_12151,N_10864);
and U17774 (N_17774,N_7950,N_10002);
nor U17775 (N_17775,N_7841,N_7280);
and U17776 (N_17776,N_8730,N_8655);
and U17777 (N_17777,N_10521,N_6960);
or U17778 (N_17778,N_7302,N_10587);
or U17779 (N_17779,N_6573,N_11063);
xnor U17780 (N_17780,N_6859,N_7460);
nand U17781 (N_17781,N_12249,N_7560);
nor U17782 (N_17782,N_8966,N_9933);
nand U17783 (N_17783,N_8943,N_8971);
xnor U17784 (N_17784,N_9992,N_12373);
nand U17785 (N_17785,N_6935,N_7359);
or U17786 (N_17786,N_7224,N_8816);
nand U17787 (N_17787,N_10836,N_10942);
and U17788 (N_17788,N_7275,N_11886);
and U17789 (N_17789,N_7599,N_12384);
and U17790 (N_17790,N_11840,N_11396);
or U17791 (N_17791,N_7786,N_8204);
nor U17792 (N_17792,N_8694,N_10378);
and U17793 (N_17793,N_11252,N_10266);
xnor U17794 (N_17794,N_9436,N_6509);
xnor U17795 (N_17795,N_9575,N_11916);
or U17796 (N_17796,N_9435,N_7114);
xor U17797 (N_17797,N_9698,N_9883);
or U17798 (N_17798,N_6255,N_8186);
nand U17799 (N_17799,N_9113,N_9750);
or U17800 (N_17800,N_8875,N_11762);
or U17801 (N_17801,N_7865,N_10538);
and U17802 (N_17802,N_8075,N_8318);
nand U17803 (N_17803,N_6463,N_11579);
or U17804 (N_17804,N_10413,N_10467);
and U17805 (N_17805,N_12367,N_7083);
nand U17806 (N_17806,N_11800,N_7400);
nor U17807 (N_17807,N_8928,N_9572);
or U17808 (N_17808,N_9737,N_12107);
nor U17809 (N_17809,N_7242,N_10660);
or U17810 (N_17810,N_10705,N_8244);
nor U17811 (N_17811,N_6720,N_9645);
nor U17812 (N_17812,N_11703,N_7763);
xnor U17813 (N_17813,N_11335,N_6374);
xnor U17814 (N_17814,N_6766,N_7347);
xor U17815 (N_17815,N_9038,N_10621);
xor U17816 (N_17816,N_6406,N_11642);
nand U17817 (N_17817,N_8095,N_7704);
nand U17818 (N_17818,N_10538,N_9298);
nand U17819 (N_17819,N_9736,N_9299);
or U17820 (N_17820,N_12469,N_6615);
nand U17821 (N_17821,N_10350,N_9667);
or U17822 (N_17822,N_7709,N_11227);
or U17823 (N_17823,N_7300,N_8918);
nor U17824 (N_17824,N_8931,N_8163);
nor U17825 (N_17825,N_10306,N_12363);
and U17826 (N_17826,N_10317,N_9855);
and U17827 (N_17827,N_9180,N_9508);
nor U17828 (N_17828,N_10601,N_12213);
nor U17829 (N_17829,N_8018,N_8832);
and U17830 (N_17830,N_9496,N_8887);
and U17831 (N_17831,N_10704,N_10177);
nor U17832 (N_17832,N_11189,N_6748);
nor U17833 (N_17833,N_8137,N_11162);
xor U17834 (N_17834,N_10997,N_6998);
xnor U17835 (N_17835,N_6490,N_10949);
xnor U17836 (N_17836,N_9437,N_9477);
xor U17837 (N_17837,N_9976,N_10597);
and U17838 (N_17838,N_12377,N_8731);
or U17839 (N_17839,N_9158,N_7430);
or U17840 (N_17840,N_8906,N_9402);
and U17841 (N_17841,N_9663,N_9380);
nor U17842 (N_17842,N_11831,N_6771);
and U17843 (N_17843,N_10595,N_12094);
nor U17844 (N_17844,N_9843,N_9708);
or U17845 (N_17845,N_12441,N_6313);
or U17846 (N_17846,N_12168,N_6993);
nor U17847 (N_17847,N_7832,N_8855);
and U17848 (N_17848,N_7914,N_6652);
xor U17849 (N_17849,N_9034,N_8760);
or U17850 (N_17850,N_9772,N_9184);
nand U17851 (N_17851,N_10590,N_11114);
or U17852 (N_17852,N_9090,N_7109);
or U17853 (N_17853,N_9458,N_10805);
xor U17854 (N_17854,N_6502,N_11242);
nand U17855 (N_17855,N_8803,N_7235);
nor U17856 (N_17856,N_11471,N_6487);
nand U17857 (N_17857,N_10403,N_6456);
nor U17858 (N_17858,N_6979,N_10065);
or U17859 (N_17859,N_9320,N_6480);
and U17860 (N_17860,N_6380,N_8391);
and U17861 (N_17861,N_7134,N_10383);
nand U17862 (N_17862,N_10051,N_7522);
and U17863 (N_17863,N_10247,N_8699);
or U17864 (N_17864,N_10872,N_7029);
nand U17865 (N_17865,N_8317,N_6254);
nand U17866 (N_17866,N_10102,N_7821);
or U17867 (N_17867,N_7722,N_11399);
nor U17868 (N_17868,N_8184,N_6528);
nor U17869 (N_17869,N_6319,N_10576);
and U17870 (N_17870,N_8051,N_12035);
nand U17871 (N_17871,N_8442,N_8432);
or U17872 (N_17872,N_7594,N_8687);
nor U17873 (N_17873,N_11701,N_12326);
or U17874 (N_17874,N_7461,N_10339);
xnor U17875 (N_17875,N_10068,N_8694);
or U17876 (N_17876,N_8734,N_9504);
nor U17877 (N_17877,N_9412,N_7536);
and U17878 (N_17878,N_6721,N_8798);
xnor U17879 (N_17879,N_7329,N_9568);
and U17880 (N_17880,N_10345,N_6936);
or U17881 (N_17881,N_7814,N_7476);
nand U17882 (N_17882,N_11972,N_10378);
nor U17883 (N_17883,N_11511,N_10327);
nor U17884 (N_17884,N_8811,N_6877);
xnor U17885 (N_17885,N_8473,N_10472);
xnor U17886 (N_17886,N_8066,N_11435);
nor U17887 (N_17887,N_10605,N_10906);
nor U17888 (N_17888,N_11848,N_9431);
nand U17889 (N_17889,N_7058,N_9785);
xor U17890 (N_17890,N_8240,N_8991);
nor U17891 (N_17891,N_9886,N_11399);
nand U17892 (N_17892,N_10807,N_7502);
or U17893 (N_17893,N_10077,N_8343);
nor U17894 (N_17894,N_9222,N_9021);
xor U17895 (N_17895,N_11017,N_7048);
or U17896 (N_17896,N_8445,N_11034);
xor U17897 (N_17897,N_8150,N_9402);
nor U17898 (N_17898,N_7906,N_8681);
and U17899 (N_17899,N_9681,N_11708);
and U17900 (N_17900,N_12423,N_11563);
xnor U17901 (N_17901,N_9967,N_10594);
nand U17902 (N_17902,N_12218,N_9104);
and U17903 (N_17903,N_11576,N_8949);
nor U17904 (N_17904,N_11168,N_9065);
nand U17905 (N_17905,N_11170,N_8030);
and U17906 (N_17906,N_9531,N_9578);
nand U17907 (N_17907,N_9410,N_8267);
or U17908 (N_17908,N_9430,N_11865);
nor U17909 (N_17909,N_9631,N_11087);
nand U17910 (N_17910,N_9334,N_12284);
nand U17911 (N_17911,N_10180,N_6299);
and U17912 (N_17912,N_11476,N_11346);
nor U17913 (N_17913,N_11222,N_11602);
nor U17914 (N_17914,N_10139,N_10849);
nor U17915 (N_17915,N_9410,N_6956);
and U17916 (N_17916,N_12193,N_8890);
or U17917 (N_17917,N_9256,N_10401);
and U17918 (N_17918,N_10933,N_12397);
nor U17919 (N_17919,N_8850,N_11786);
nor U17920 (N_17920,N_8812,N_9428);
and U17921 (N_17921,N_8164,N_12475);
nand U17922 (N_17922,N_11533,N_10698);
nor U17923 (N_17923,N_8931,N_8348);
and U17924 (N_17924,N_9757,N_10950);
nand U17925 (N_17925,N_11290,N_9717);
nor U17926 (N_17926,N_7673,N_7453);
xnor U17927 (N_17927,N_11432,N_9462);
nor U17928 (N_17928,N_11379,N_8950);
and U17929 (N_17929,N_6258,N_7159);
nor U17930 (N_17930,N_7737,N_10348);
nor U17931 (N_17931,N_9556,N_7541);
nand U17932 (N_17932,N_9334,N_10309);
nor U17933 (N_17933,N_8757,N_11707);
and U17934 (N_17934,N_8324,N_8687);
or U17935 (N_17935,N_7446,N_8339);
nor U17936 (N_17936,N_11927,N_11816);
and U17937 (N_17937,N_11995,N_7770);
or U17938 (N_17938,N_7105,N_7708);
nand U17939 (N_17939,N_10288,N_6995);
nor U17940 (N_17940,N_11906,N_6370);
xor U17941 (N_17941,N_8571,N_12398);
nand U17942 (N_17942,N_9766,N_12001);
nand U17943 (N_17943,N_8901,N_6319);
xnor U17944 (N_17944,N_8888,N_6629);
xor U17945 (N_17945,N_11518,N_9302);
nor U17946 (N_17946,N_7386,N_6438);
nor U17947 (N_17947,N_11120,N_7534);
and U17948 (N_17948,N_7390,N_9752);
xor U17949 (N_17949,N_8084,N_11392);
nor U17950 (N_17950,N_9835,N_9225);
xnor U17951 (N_17951,N_7228,N_7817);
nor U17952 (N_17952,N_9881,N_9926);
xnor U17953 (N_17953,N_7868,N_6686);
nand U17954 (N_17954,N_10508,N_10662);
or U17955 (N_17955,N_10158,N_10310);
or U17956 (N_17956,N_8024,N_7845);
and U17957 (N_17957,N_6334,N_6393);
nand U17958 (N_17958,N_7767,N_8962);
nand U17959 (N_17959,N_12128,N_10979);
and U17960 (N_17960,N_10569,N_7046);
and U17961 (N_17961,N_7900,N_6503);
nor U17962 (N_17962,N_7290,N_9526);
or U17963 (N_17963,N_10544,N_11051);
xor U17964 (N_17964,N_11410,N_7893);
and U17965 (N_17965,N_9398,N_11436);
nor U17966 (N_17966,N_9958,N_8240);
and U17967 (N_17967,N_8983,N_12208);
xor U17968 (N_17968,N_10221,N_9876);
nand U17969 (N_17969,N_8858,N_8130);
and U17970 (N_17970,N_10710,N_7124);
or U17971 (N_17971,N_6542,N_6254);
or U17972 (N_17972,N_7204,N_8361);
or U17973 (N_17973,N_10941,N_12162);
nand U17974 (N_17974,N_7637,N_12498);
nor U17975 (N_17975,N_6601,N_10515);
xnor U17976 (N_17976,N_7106,N_6441);
and U17977 (N_17977,N_6487,N_11747);
xor U17978 (N_17978,N_12237,N_9730);
and U17979 (N_17979,N_6274,N_11115);
nor U17980 (N_17980,N_9534,N_9865);
nand U17981 (N_17981,N_10264,N_7683);
nand U17982 (N_17982,N_9422,N_6980);
and U17983 (N_17983,N_8147,N_6518);
and U17984 (N_17984,N_6719,N_12342);
nor U17985 (N_17985,N_10525,N_10160);
nand U17986 (N_17986,N_10566,N_11722);
xor U17987 (N_17987,N_8390,N_10798);
xnor U17988 (N_17988,N_9038,N_11349);
and U17989 (N_17989,N_11000,N_11536);
or U17990 (N_17990,N_7450,N_9217);
or U17991 (N_17991,N_8163,N_7929);
xnor U17992 (N_17992,N_7271,N_12456);
nand U17993 (N_17993,N_8608,N_11440);
or U17994 (N_17994,N_9954,N_12218);
nor U17995 (N_17995,N_8147,N_8428);
or U17996 (N_17996,N_11103,N_8404);
xnor U17997 (N_17997,N_9741,N_9185);
nor U17998 (N_17998,N_7477,N_11439);
or U17999 (N_17999,N_10464,N_7569);
or U18000 (N_18000,N_12410,N_8656);
or U18001 (N_18001,N_10054,N_7110);
xnor U18002 (N_18002,N_11382,N_8828);
xnor U18003 (N_18003,N_6345,N_11755);
nor U18004 (N_18004,N_9289,N_12461);
and U18005 (N_18005,N_10022,N_8604);
xnor U18006 (N_18006,N_10005,N_6972);
nand U18007 (N_18007,N_11898,N_7443);
nor U18008 (N_18008,N_11559,N_6487);
nor U18009 (N_18009,N_11297,N_9435);
nor U18010 (N_18010,N_7588,N_6793);
nand U18011 (N_18011,N_9837,N_11384);
and U18012 (N_18012,N_11372,N_11606);
nand U18013 (N_18013,N_7985,N_7465);
or U18014 (N_18014,N_12202,N_11584);
and U18015 (N_18015,N_8162,N_8747);
xnor U18016 (N_18016,N_9816,N_10793);
xor U18017 (N_18017,N_7826,N_11202);
xnor U18018 (N_18018,N_11285,N_7612);
and U18019 (N_18019,N_6345,N_7301);
and U18020 (N_18020,N_6402,N_7024);
nor U18021 (N_18021,N_8633,N_7501);
xor U18022 (N_18022,N_9719,N_7531);
and U18023 (N_18023,N_10434,N_9137);
or U18024 (N_18024,N_10750,N_8990);
nor U18025 (N_18025,N_6802,N_11354);
and U18026 (N_18026,N_11023,N_11425);
and U18027 (N_18027,N_12033,N_9563);
xnor U18028 (N_18028,N_9227,N_6277);
nand U18029 (N_18029,N_10238,N_8181);
and U18030 (N_18030,N_7555,N_9485);
nand U18031 (N_18031,N_6644,N_10972);
xnor U18032 (N_18032,N_9326,N_8083);
nor U18033 (N_18033,N_10873,N_8789);
and U18034 (N_18034,N_6532,N_7224);
nand U18035 (N_18035,N_7171,N_8159);
and U18036 (N_18036,N_9916,N_9137);
nand U18037 (N_18037,N_8573,N_11555);
or U18038 (N_18038,N_8768,N_7403);
nand U18039 (N_18039,N_6417,N_10666);
xor U18040 (N_18040,N_12393,N_11725);
nor U18041 (N_18041,N_8660,N_11506);
xor U18042 (N_18042,N_12145,N_9555);
or U18043 (N_18043,N_12069,N_10235);
xor U18044 (N_18044,N_9252,N_7007);
nand U18045 (N_18045,N_12405,N_11215);
or U18046 (N_18046,N_8432,N_9450);
xor U18047 (N_18047,N_7164,N_6812);
xor U18048 (N_18048,N_10428,N_11707);
or U18049 (N_18049,N_7521,N_7820);
and U18050 (N_18050,N_10449,N_7403);
or U18051 (N_18051,N_12192,N_11273);
and U18052 (N_18052,N_10714,N_12456);
nand U18053 (N_18053,N_6310,N_9224);
or U18054 (N_18054,N_10897,N_8565);
and U18055 (N_18055,N_7307,N_9919);
and U18056 (N_18056,N_11661,N_6666);
nor U18057 (N_18057,N_7852,N_12343);
or U18058 (N_18058,N_7170,N_11138);
or U18059 (N_18059,N_10079,N_7937);
nand U18060 (N_18060,N_11128,N_11380);
nor U18061 (N_18061,N_8516,N_10962);
or U18062 (N_18062,N_8267,N_8500);
nand U18063 (N_18063,N_9174,N_12259);
xor U18064 (N_18064,N_10417,N_10865);
and U18065 (N_18065,N_9338,N_11562);
and U18066 (N_18066,N_10003,N_11260);
nor U18067 (N_18067,N_6334,N_8501);
xnor U18068 (N_18068,N_11724,N_11089);
xor U18069 (N_18069,N_9810,N_10595);
xor U18070 (N_18070,N_7393,N_11399);
xnor U18071 (N_18071,N_7911,N_7891);
xor U18072 (N_18072,N_10596,N_8155);
nor U18073 (N_18073,N_7392,N_6613);
or U18074 (N_18074,N_6941,N_9652);
nand U18075 (N_18075,N_7713,N_7963);
or U18076 (N_18076,N_7988,N_8722);
or U18077 (N_18077,N_9709,N_8803);
and U18078 (N_18078,N_12395,N_9232);
or U18079 (N_18079,N_10923,N_9510);
or U18080 (N_18080,N_12300,N_11868);
and U18081 (N_18081,N_6582,N_10675);
or U18082 (N_18082,N_11773,N_10089);
xnor U18083 (N_18083,N_7739,N_6977);
xor U18084 (N_18084,N_6572,N_8742);
nand U18085 (N_18085,N_8286,N_12034);
and U18086 (N_18086,N_8473,N_11051);
nor U18087 (N_18087,N_6435,N_12048);
nor U18088 (N_18088,N_6250,N_11395);
xnor U18089 (N_18089,N_7206,N_8878);
nand U18090 (N_18090,N_10488,N_9509);
or U18091 (N_18091,N_7218,N_9679);
xor U18092 (N_18092,N_11735,N_8625);
nor U18093 (N_18093,N_6429,N_12163);
or U18094 (N_18094,N_11579,N_10342);
and U18095 (N_18095,N_7328,N_12399);
nor U18096 (N_18096,N_11275,N_8861);
nand U18097 (N_18097,N_12058,N_11961);
and U18098 (N_18098,N_9216,N_6899);
and U18099 (N_18099,N_6451,N_9130);
nand U18100 (N_18100,N_11465,N_6705);
nand U18101 (N_18101,N_9775,N_11315);
or U18102 (N_18102,N_10171,N_6990);
nor U18103 (N_18103,N_8614,N_9420);
nor U18104 (N_18104,N_9101,N_10600);
nand U18105 (N_18105,N_11325,N_8846);
or U18106 (N_18106,N_6602,N_9502);
xnor U18107 (N_18107,N_8732,N_9811);
nor U18108 (N_18108,N_8329,N_7468);
and U18109 (N_18109,N_7895,N_7078);
or U18110 (N_18110,N_10396,N_11000);
nand U18111 (N_18111,N_6490,N_8357);
xnor U18112 (N_18112,N_10814,N_9141);
xnor U18113 (N_18113,N_11340,N_9826);
nand U18114 (N_18114,N_9380,N_6984);
or U18115 (N_18115,N_8570,N_11702);
nand U18116 (N_18116,N_9502,N_10656);
nand U18117 (N_18117,N_9047,N_6561);
or U18118 (N_18118,N_7595,N_10984);
nor U18119 (N_18119,N_8762,N_9784);
or U18120 (N_18120,N_9515,N_7271);
and U18121 (N_18121,N_7742,N_10418);
nand U18122 (N_18122,N_7005,N_9896);
nor U18123 (N_18123,N_7814,N_10328);
and U18124 (N_18124,N_6733,N_9074);
nand U18125 (N_18125,N_11644,N_10635);
and U18126 (N_18126,N_8224,N_10681);
and U18127 (N_18127,N_8239,N_7102);
and U18128 (N_18128,N_6672,N_9840);
xnor U18129 (N_18129,N_7528,N_6474);
or U18130 (N_18130,N_9369,N_11612);
nor U18131 (N_18131,N_10364,N_8949);
nand U18132 (N_18132,N_9153,N_10296);
nand U18133 (N_18133,N_7193,N_10672);
xor U18134 (N_18134,N_7199,N_11864);
xnor U18135 (N_18135,N_7512,N_9994);
or U18136 (N_18136,N_6700,N_8288);
xor U18137 (N_18137,N_8003,N_6338);
or U18138 (N_18138,N_10570,N_7497);
and U18139 (N_18139,N_11209,N_10976);
xor U18140 (N_18140,N_9264,N_12100);
nand U18141 (N_18141,N_6720,N_11020);
nand U18142 (N_18142,N_11811,N_6781);
xnor U18143 (N_18143,N_10807,N_7448);
nor U18144 (N_18144,N_10990,N_8996);
or U18145 (N_18145,N_7646,N_9770);
nand U18146 (N_18146,N_6866,N_8464);
nand U18147 (N_18147,N_9550,N_7588);
xnor U18148 (N_18148,N_11127,N_11292);
and U18149 (N_18149,N_8115,N_12197);
nor U18150 (N_18150,N_12135,N_7645);
or U18151 (N_18151,N_8023,N_11606);
xnor U18152 (N_18152,N_11814,N_9032);
xnor U18153 (N_18153,N_7217,N_8673);
nor U18154 (N_18154,N_9452,N_6809);
nor U18155 (N_18155,N_8918,N_11089);
or U18156 (N_18156,N_11699,N_12066);
and U18157 (N_18157,N_11275,N_7427);
or U18158 (N_18158,N_9402,N_7064);
and U18159 (N_18159,N_10959,N_11914);
xor U18160 (N_18160,N_9466,N_10463);
and U18161 (N_18161,N_8469,N_12094);
nand U18162 (N_18162,N_7215,N_10965);
nor U18163 (N_18163,N_11001,N_8877);
and U18164 (N_18164,N_9885,N_11211);
nand U18165 (N_18165,N_12337,N_9933);
xor U18166 (N_18166,N_11810,N_8310);
or U18167 (N_18167,N_7773,N_9687);
or U18168 (N_18168,N_6630,N_9486);
and U18169 (N_18169,N_11427,N_11188);
or U18170 (N_18170,N_10778,N_9432);
nor U18171 (N_18171,N_12499,N_11639);
and U18172 (N_18172,N_11564,N_11022);
nor U18173 (N_18173,N_9500,N_7740);
or U18174 (N_18174,N_7100,N_10153);
or U18175 (N_18175,N_8514,N_6774);
or U18176 (N_18176,N_7078,N_10815);
and U18177 (N_18177,N_8304,N_6692);
nand U18178 (N_18178,N_10120,N_8492);
nor U18179 (N_18179,N_6701,N_10157);
xor U18180 (N_18180,N_10688,N_9426);
nor U18181 (N_18181,N_6325,N_7277);
nand U18182 (N_18182,N_6459,N_9989);
nand U18183 (N_18183,N_6998,N_9892);
nand U18184 (N_18184,N_9106,N_8690);
nor U18185 (N_18185,N_8395,N_7004);
and U18186 (N_18186,N_6772,N_7206);
or U18187 (N_18187,N_11604,N_9887);
or U18188 (N_18188,N_11265,N_9602);
nand U18189 (N_18189,N_11147,N_11698);
nand U18190 (N_18190,N_6819,N_9893);
xnor U18191 (N_18191,N_9627,N_7782);
xor U18192 (N_18192,N_9369,N_9306);
nor U18193 (N_18193,N_11695,N_9109);
nor U18194 (N_18194,N_6852,N_12086);
nor U18195 (N_18195,N_10867,N_6508);
and U18196 (N_18196,N_7495,N_8878);
nand U18197 (N_18197,N_9396,N_8153);
and U18198 (N_18198,N_8444,N_10397);
or U18199 (N_18199,N_6584,N_7225);
xor U18200 (N_18200,N_10648,N_6367);
or U18201 (N_18201,N_7666,N_10777);
or U18202 (N_18202,N_11197,N_11399);
and U18203 (N_18203,N_8627,N_6464);
nand U18204 (N_18204,N_12147,N_12302);
and U18205 (N_18205,N_9940,N_11894);
nor U18206 (N_18206,N_8518,N_8405);
nand U18207 (N_18207,N_7044,N_6380);
nor U18208 (N_18208,N_7477,N_9353);
and U18209 (N_18209,N_11936,N_9867);
and U18210 (N_18210,N_12323,N_8451);
nor U18211 (N_18211,N_9310,N_12058);
and U18212 (N_18212,N_11187,N_9061);
or U18213 (N_18213,N_10033,N_9555);
or U18214 (N_18214,N_6512,N_8371);
and U18215 (N_18215,N_9893,N_9187);
and U18216 (N_18216,N_7658,N_9704);
xnor U18217 (N_18217,N_10634,N_8018);
or U18218 (N_18218,N_9056,N_7270);
xnor U18219 (N_18219,N_9031,N_8901);
nor U18220 (N_18220,N_7545,N_9388);
or U18221 (N_18221,N_11198,N_8100);
nor U18222 (N_18222,N_11918,N_10395);
or U18223 (N_18223,N_12096,N_8990);
or U18224 (N_18224,N_8912,N_6278);
xor U18225 (N_18225,N_10089,N_6609);
xor U18226 (N_18226,N_7068,N_8223);
nor U18227 (N_18227,N_6541,N_6668);
xnor U18228 (N_18228,N_9057,N_8565);
nor U18229 (N_18229,N_9711,N_12398);
nor U18230 (N_18230,N_7110,N_10793);
nor U18231 (N_18231,N_9675,N_7917);
nor U18232 (N_18232,N_9446,N_11121);
xnor U18233 (N_18233,N_9189,N_7325);
or U18234 (N_18234,N_9062,N_9572);
or U18235 (N_18235,N_10901,N_11983);
or U18236 (N_18236,N_6762,N_7022);
nor U18237 (N_18237,N_12403,N_8094);
nor U18238 (N_18238,N_10933,N_10644);
and U18239 (N_18239,N_9081,N_11635);
nor U18240 (N_18240,N_7574,N_10723);
nand U18241 (N_18241,N_9349,N_12015);
and U18242 (N_18242,N_8659,N_7210);
or U18243 (N_18243,N_7854,N_7524);
or U18244 (N_18244,N_10587,N_7689);
or U18245 (N_18245,N_11740,N_9436);
and U18246 (N_18246,N_7083,N_9336);
nor U18247 (N_18247,N_6741,N_6891);
nand U18248 (N_18248,N_10624,N_10303);
xnor U18249 (N_18249,N_11417,N_7030);
nand U18250 (N_18250,N_10892,N_6615);
nor U18251 (N_18251,N_6509,N_11820);
xor U18252 (N_18252,N_9961,N_8724);
and U18253 (N_18253,N_12116,N_11937);
nand U18254 (N_18254,N_11314,N_10395);
and U18255 (N_18255,N_12371,N_11791);
nand U18256 (N_18256,N_9715,N_7516);
nand U18257 (N_18257,N_9089,N_11133);
xor U18258 (N_18258,N_7059,N_7798);
nor U18259 (N_18259,N_8206,N_8114);
and U18260 (N_18260,N_6427,N_12400);
nor U18261 (N_18261,N_9081,N_7808);
nor U18262 (N_18262,N_6993,N_12429);
xnor U18263 (N_18263,N_6687,N_7888);
or U18264 (N_18264,N_10087,N_12291);
and U18265 (N_18265,N_10415,N_8967);
nor U18266 (N_18266,N_12059,N_12498);
nor U18267 (N_18267,N_12127,N_11233);
or U18268 (N_18268,N_10414,N_8641);
nand U18269 (N_18269,N_9059,N_12212);
nor U18270 (N_18270,N_8162,N_7618);
or U18271 (N_18271,N_12376,N_10547);
xnor U18272 (N_18272,N_7654,N_6469);
and U18273 (N_18273,N_9351,N_8237);
nor U18274 (N_18274,N_12119,N_6662);
or U18275 (N_18275,N_9687,N_6500);
nor U18276 (N_18276,N_9300,N_8772);
nor U18277 (N_18277,N_10583,N_7717);
nor U18278 (N_18278,N_9176,N_11846);
and U18279 (N_18279,N_11491,N_8253);
nor U18280 (N_18280,N_9799,N_8467);
nand U18281 (N_18281,N_7389,N_7961);
or U18282 (N_18282,N_7808,N_7971);
nor U18283 (N_18283,N_8416,N_8853);
and U18284 (N_18284,N_12117,N_10703);
and U18285 (N_18285,N_7762,N_9435);
nor U18286 (N_18286,N_10165,N_10246);
nor U18287 (N_18287,N_11238,N_9046);
nand U18288 (N_18288,N_10628,N_7506);
nand U18289 (N_18289,N_12478,N_11526);
or U18290 (N_18290,N_11048,N_8350);
xor U18291 (N_18291,N_10823,N_9998);
nand U18292 (N_18292,N_11165,N_10501);
xor U18293 (N_18293,N_9342,N_10169);
or U18294 (N_18294,N_9974,N_10566);
and U18295 (N_18295,N_7990,N_12423);
or U18296 (N_18296,N_7171,N_10731);
xnor U18297 (N_18297,N_10587,N_11691);
xor U18298 (N_18298,N_6272,N_11466);
nor U18299 (N_18299,N_8400,N_9318);
nand U18300 (N_18300,N_11206,N_11337);
xor U18301 (N_18301,N_11203,N_7158);
and U18302 (N_18302,N_8205,N_7031);
xnor U18303 (N_18303,N_6831,N_6463);
nand U18304 (N_18304,N_9793,N_12345);
nor U18305 (N_18305,N_6270,N_11724);
and U18306 (N_18306,N_7538,N_11502);
and U18307 (N_18307,N_7181,N_7546);
or U18308 (N_18308,N_11386,N_10973);
and U18309 (N_18309,N_6276,N_9206);
nor U18310 (N_18310,N_10713,N_6623);
nor U18311 (N_18311,N_11739,N_11275);
nor U18312 (N_18312,N_7477,N_11483);
xnor U18313 (N_18313,N_6899,N_8083);
nor U18314 (N_18314,N_7491,N_7084);
xnor U18315 (N_18315,N_9829,N_7572);
nand U18316 (N_18316,N_9619,N_9837);
xnor U18317 (N_18317,N_11451,N_9028);
nor U18318 (N_18318,N_12225,N_6374);
nor U18319 (N_18319,N_7481,N_8599);
nand U18320 (N_18320,N_7733,N_12410);
xnor U18321 (N_18321,N_8457,N_10864);
or U18322 (N_18322,N_6321,N_10923);
xnor U18323 (N_18323,N_6554,N_6992);
nor U18324 (N_18324,N_7552,N_9766);
nand U18325 (N_18325,N_6567,N_6886);
and U18326 (N_18326,N_7027,N_10024);
and U18327 (N_18327,N_7722,N_7810);
nor U18328 (N_18328,N_8909,N_9471);
or U18329 (N_18329,N_12366,N_9825);
nand U18330 (N_18330,N_9104,N_9483);
nand U18331 (N_18331,N_9929,N_10911);
or U18332 (N_18332,N_10782,N_10898);
or U18333 (N_18333,N_7395,N_8151);
nand U18334 (N_18334,N_10204,N_7396);
and U18335 (N_18335,N_10540,N_6406);
or U18336 (N_18336,N_9978,N_7780);
nand U18337 (N_18337,N_8451,N_8324);
or U18338 (N_18338,N_8802,N_8713);
or U18339 (N_18339,N_10572,N_11698);
or U18340 (N_18340,N_8096,N_11326);
and U18341 (N_18341,N_10914,N_9356);
nand U18342 (N_18342,N_7055,N_11430);
or U18343 (N_18343,N_6778,N_8666);
or U18344 (N_18344,N_7323,N_8992);
or U18345 (N_18345,N_9856,N_10160);
and U18346 (N_18346,N_9957,N_11583);
nand U18347 (N_18347,N_11289,N_6310);
nand U18348 (N_18348,N_9175,N_12258);
and U18349 (N_18349,N_11481,N_10654);
xnor U18350 (N_18350,N_12293,N_7753);
nand U18351 (N_18351,N_11648,N_11846);
nand U18352 (N_18352,N_9302,N_10530);
or U18353 (N_18353,N_8831,N_11047);
and U18354 (N_18354,N_10275,N_7584);
and U18355 (N_18355,N_9061,N_10426);
and U18356 (N_18356,N_6645,N_11773);
or U18357 (N_18357,N_9091,N_7696);
nand U18358 (N_18358,N_7802,N_10970);
nor U18359 (N_18359,N_6477,N_10585);
or U18360 (N_18360,N_10335,N_11773);
nor U18361 (N_18361,N_12251,N_10481);
nand U18362 (N_18362,N_7239,N_6510);
xnor U18363 (N_18363,N_9652,N_6806);
or U18364 (N_18364,N_12353,N_8496);
xor U18365 (N_18365,N_7033,N_11556);
and U18366 (N_18366,N_10986,N_10037);
nand U18367 (N_18367,N_6684,N_8661);
nand U18368 (N_18368,N_9170,N_12192);
nand U18369 (N_18369,N_6326,N_6580);
and U18370 (N_18370,N_6346,N_9791);
and U18371 (N_18371,N_10459,N_10747);
and U18372 (N_18372,N_6298,N_11084);
nor U18373 (N_18373,N_8342,N_12220);
and U18374 (N_18374,N_6437,N_7385);
nand U18375 (N_18375,N_10495,N_9967);
and U18376 (N_18376,N_7352,N_10533);
or U18377 (N_18377,N_10828,N_9686);
and U18378 (N_18378,N_11806,N_9820);
or U18379 (N_18379,N_7319,N_7789);
nor U18380 (N_18380,N_12115,N_7165);
or U18381 (N_18381,N_10961,N_6983);
and U18382 (N_18382,N_11637,N_11674);
nor U18383 (N_18383,N_12391,N_7536);
nand U18384 (N_18384,N_7414,N_10575);
xnor U18385 (N_18385,N_9319,N_8382);
nor U18386 (N_18386,N_8110,N_6593);
nor U18387 (N_18387,N_9949,N_8319);
or U18388 (N_18388,N_9179,N_10464);
or U18389 (N_18389,N_8596,N_6752);
nand U18390 (N_18390,N_10673,N_7590);
xor U18391 (N_18391,N_7791,N_12298);
or U18392 (N_18392,N_9524,N_6370);
or U18393 (N_18393,N_10863,N_10238);
nand U18394 (N_18394,N_7159,N_8787);
xnor U18395 (N_18395,N_6583,N_11540);
nor U18396 (N_18396,N_7176,N_10282);
or U18397 (N_18397,N_6597,N_11545);
or U18398 (N_18398,N_10319,N_8722);
xnor U18399 (N_18399,N_7296,N_9388);
or U18400 (N_18400,N_7800,N_9539);
xor U18401 (N_18401,N_12276,N_7815);
xnor U18402 (N_18402,N_11857,N_11310);
nor U18403 (N_18403,N_11246,N_6765);
or U18404 (N_18404,N_6989,N_7513);
and U18405 (N_18405,N_11432,N_10642);
nor U18406 (N_18406,N_9519,N_10166);
or U18407 (N_18407,N_10723,N_7870);
and U18408 (N_18408,N_10533,N_9622);
or U18409 (N_18409,N_11757,N_12467);
or U18410 (N_18410,N_11454,N_10703);
nand U18411 (N_18411,N_9331,N_12086);
and U18412 (N_18412,N_11645,N_12407);
nor U18413 (N_18413,N_7007,N_8892);
nor U18414 (N_18414,N_9464,N_6720);
nor U18415 (N_18415,N_9014,N_10239);
nand U18416 (N_18416,N_6697,N_11534);
and U18417 (N_18417,N_8023,N_7471);
and U18418 (N_18418,N_7149,N_11982);
and U18419 (N_18419,N_9620,N_6982);
nor U18420 (N_18420,N_6293,N_9879);
nor U18421 (N_18421,N_6692,N_7079);
nor U18422 (N_18422,N_7696,N_7439);
or U18423 (N_18423,N_10941,N_6560);
nor U18424 (N_18424,N_8688,N_8349);
xnor U18425 (N_18425,N_6660,N_9485);
nand U18426 (N_18426,N_8169,N_7339);
xnor U18427 (N_18427,N_12475,N_12012);
and U18428 (N_18428,N_8362,N_8289);
nand U18429 (N_18429,N_6475,N_7381);
or U18430 (N_18430,N_8694,N_6604);
nor U18431 (N_18431,N_11268,N_12057);
and U18432 (N_18432,N_8378,N_10673);
nor U18433 (N_18433,N_8798,N_7749);
or U18434 (N_18434,N_7962,N_11043);
nand U18435 (N_18435,N_10479,N_10529);
nor U18436 (N_18436,N_11971,N_9913);
and U18437 (N_18437,N_10432,N_6727);
and U18438 (N_18438,N_11757,N_9196);
or U18439 (N_18439,N_9893,N_7084);
nand U18440 (N_18440,N_10930,N_11798);
nand U18441 (N_18441,N_11009,N_10807);
or U18442 (N_18442,N_9689,N_7144);
nand U18443 (N_18443,N_6639,N_9757);
nor U18444 (N_18444,N_11288,N_8650);
nor U18445 (N_18445,N_6404,N_6403);
or U18446 (N_18446,N_12392,N_7084);
or U18447 (N_18447,N_11287,N_10218);
nor U18448 (N_18448,N_12109,N_11147);
xnor U18449 (N_18449,N_10122,N_8161);
xor U18450 (N_18450,N_12126,N_7393);
and U18451 (N_18451,N_9751,N_6486);
or U18452 (N_18452,N_11067,N_8084);
nor U18453 (N_18453,N_6377,N_10522);
xor U18454 (N_18454,N_8401,N_9646);
nor U18455 (N_18455,N_6310,N_11232);
and U18456 (N_18456,N_9356,N_11511);
or U18457 (N_18457,N_8456,N_10402);
xor U18458 (N_18458,N_12291,N_6626);
or U18459 (N_18459,N_6755,N_8557);
xor U18460 (N_18460,N_9606,N_9770);
nand U18461 (N_18461,N_10706,N_8962);
nor U18462 (N_18462,N_8583,N_11511);
xnor U18463 (N_18463,N_11515,N_6571);
nand U18464 (N_18464,N_8015,N_11167);
xor U18465 (N_18465,N_11407,N_11717);
or U18466 (N_18466,N_7181,N_8790);
nand U18467 (N_18467,N_6809,N_12006);
or U18468 (N_18468,N_11591,N_10012);
and U18469 (N_18469,N_7134,N_9026);
xnor U18470 (N_18470,N_8986,N_8250);
and U18471 (N_18471,N_9798,N_8264);
or U18472 (N_18472,N_6972,N_7965);
or U18473 (N_18473,N_9473,N_6596);
nor U18474 (N_18474,N_8554,N_11384);
nor U18475 (N_18475,N_9329,N_10864);
or U18476 (N_18476,N_10337,N_11040);
and U18477 (N_18477,N_6665,N_10839);
or U18478 (N_18478,N_12139,N_6357);
xor U18479 (N_18479,N_11596,N_10934);
nor U18480 (N_18480,N_12482,N_8870);
or U18481 (N_18481,N_6311,N_8604);
nor U18482 (N_18482,N_11838,N_10517);
xor U18483 (N_18483,N_6737,N_9762);
and U18484 (N_18484,N_10300,N_6414);
xnor U18485 (N_18485,N_9988,N_11055);
and U18486 (N_18486,N_6778,N_9205);
and U18487 (N_18487,N_12459,N_10941);
nand U18488 (N_18488,N_10837,N_10084);
nand U18489 (N_18489,N_8915,N_7624);
xor U18490 (N_18490,N_8738,N_10395);
nand U18491 (N_18491,N_9448,N_12250);
and U18492 (N_18492,N_7300,N_11179);
nand U18493 (N_18493,N_10724,N_9376);
nand U18494 (N_18494,N_10277,N_12248);
and U18495 (N_18495,N_6495,N_10565);
nand U18496 (N_18496,N_11518,N_6961);
nor U18497 (N_18497,N_10247,N_7875);
and U18498 (N_18498,N_11637,N_7313);
and U18499 (N_18499,N_11551,N_11762);
xor U18500 (N_18500,N_7437,N_10015);
xor U18501 (N_18501,N_9052,N_9431);
or U18502 (N_18502,N_10044,N_11901);
xnor U18503 (N_18503,N_8877,N_8918);
nand U18504 (N_18504,N_10761,N_6796);
and U18505 (N_18505,N_12284,N_9849);
and U18506 (N_18506,N_7891,N_12338);
nand U18507 (N_18507,N_8914,N_6454);
nand U18508 (N_18508,N_7457,N_6991);
nor U18509 (N_18509,N_6563,N_9069);
and U18510 (N_18510,N_10441,N_7601);
nand U18511 (N_18511,N_6338,N_10942);
nand U18512 (N_18512,N_7804,N_9717);
nor U18513 (N_18513,N_12151,N_8179);
and U18514 (N_18514,N_6852,N_10860);
nor U18515 (N_18515,N_9350,N_7828);
or U18516 (N_18516,N_7895,N_9598);
or U18517 (N_18517,N_11026,N_11139);
xor U18518 (N_18518,N_7162,N_11607);
or U18519 (N_18519,N_6787,N_12082);
nor U18520 (N_18520,N_9090,N_8809);
xnor U18521 (N_18521,N_7807,N_11188);
and U18522 (N_18522,N_8982,N_10830);
nor U18523 (N_18523,N_10875,N_8965);
nand U18524 (N_18524,N_12017,N_7870);
or U18525 (N_18525,N_7784,N_11735);
or U18526 (N_18526,N_6373,N_8630);
nor U18527 (N_18527,N_7885,N_9583);
or U18528 (N_18528,N_10276,N_10444);
xor U18529 (N_18529,N_7650,N_11807);
or U18530 (N_18530,N_10829,N_7862);
xnor U18531 (N_18531,N_12154,N_7148);
and U18532 (N_18532,N_11004,N_6762);
nor U18533 (N_18533,N_7096,N_9214);
and U18534 (N_18534,N_11621,N_9123);
nor U18535 (N_18535,N_9934,N_10609);
and U18536 (N_18536,N_7106,N_7474);
nand U18537 (N_18537,N_9692,N_10391);
nand U18538 (N_18538,N_9699,N_10466);
or U18539 (N_18539,N_6469,N_11183);
xor U18540 (N_18540,N_7428,N_7272);
and U18541 (N_18541,N_10510,N_6398);
nand U18542 (N_18542,N_10644,N_12075);
nand U18543 (N_18543,N_11374,N_10241);
nand U18544 (N_18544,N_7273,N_9535);
or U18545 (N_18545,N_6580,N_10090);
xnor U18546 (N_18546,N_9730,N_8745);
and U18547 (N_18547,N_11251,N_7199);
xor U18548 (N_18548,N_8325,N_8220);
xnor U18549 (N_18549,N_7230,N_11742);
nor U18550 (N_18550,N_11670,N_10268);
xnor U18551 (N_18551,N_10522,N_8034);
and U18552 (N_18552,N_11569,N_11600);
nand U18553 (N_18553,N_11358,N_11258);
and U18554 (N_18554,N_9044,N_8276);
and U18555 (N_18555,N_8340,N_9993);
nor U18556 (N_18556,N_7267,N_9665);
and U18557 (N_18557,N_11670,N_7245);
nor U18558 (N_18558,N_6855,N_8349);
nor U18559 (N_18559,N_10878,N_10551);
or U18560 (N_18560,N_7303,N_12202);
nor U18561 (N_18561,N_7213,N_8130);
or U18562 (N_18562,N_8975,N_11613);
xor U18563 (N_18563,N_7087,N_6919);
xnor U18564 (N_18564,N_8278,N_10724);
nand U18565 (N_18565,N_7598,N_11500);
nand U18566 (N_18566,N_8060,N_9630);
or U18567 (N_18567,N_9072,N_8408);
or U18568 (N_18568,N_11281,N_7060);
xor U18569 (N_18569,N_7477,N_9982);
or U18570 (N_18570,N_11120,N_9172);
nor U18571 (N_18571,N_6391,N_9413);
or U18572 (N_18572,N_12113,N_7587);
xor U18573 (N_18573,N_8797,N_7556);
nor U18574 (N_18574,N_10972,N_11780);
or U18575 (N_18575,N_7381,N_11798);
and U18576 (N_18576,N_8608,N_12448);
xnor U18577 (N_18577,N_7435,N_11828);
xnor U18578 (N_18578,N_12176,N_7007);
nand U18579 (N_18579,N_11173,N_6494);
nand U18580 (N_18580,N_8348,N_9547);
nand U18581 (N_18581,N_11156,N_9380);
nor U18582 (N_18582,N_12476,N_10515);
nand U18583 (N_18583,N_11081,N_11819);
xnor U18584 (N_18584,N_10002,N_11515);
nand U18585 (N_18585,N_7480,N_12182);
nor U18586 (N_18586,N_12295,N_11749);
or U18587 (N_18587,N_9130,N_10600);
nor U18588 (N_18588,N_9578,N_8093);
and U18589 (N_18589,N_12319,N_7422);
nand U18590 (N_18590,N_11081,N_9561);
nor U18591 (N_18591,N_12019,N_8564);
nand U18592 (N_18592,N_12171,N_8569);
or U18593 (N_18593,N_9881,N_10346);
nand U18594 (N_18594,N_7760,N_9815);
nor U18595 (N_18595,N_8746,N_9148);
xnor U18596 (N_18596,N_9312,N_7837);
nor U18597 (N_18597,N_7379,N_6585);
xnor U18598 (N_18598,N_11097,N_7394);
and U18599 (N_18599,N_9375,N_10883);
nor U18600 (N_18600,N_10140,N_12350);
nand U18601 (N_18601,N_11750,N_10235);
xor U18602 (N_18602,N_11606,N_10061);
nand U18603 (N_18603,N_7448,N_6947);
or U18604 (N_18604,N_6938,N_9557);
nor U18605 (N_18605,N_11012,N_7088);
nand U18606 (N_18606,N_12108,N_6981);
and U18607 (N_18607,N_11547,N_11601);
xor U18608 (N_18608,N_10300,N_10402);
nor U18609 (N_18609,N_10510,N_9521);
or U18610 (N_18610,N_12101,N_8714);
or U18611 (N_18611,N_7550,N_12148);
nand U18612 (N_18612,N_10528,N_11779);
nor U18613 (N_18613,N_7694,N_6256);
and U18614 (N_18614,N_11987,N_11623);
nor U18615 (N_18615,N_8251,N_6934);
nor U18616 (N_18616,N_9830,N_6902);
xor U18617 (N_18617,N_9439,N_7329);
nand U18618 (N_18618,N_7446,N_7894);
xor U18619 (N_18619,N_11504,N_12420);
nor U18620 (N_18620,N_9810,N_10380);
xnor U18621 (N_18621,N_7034,N_8433);
nand U18622 (N_18622,N_8266,N_11745);
and U18623 (N_18623,N_7463,N_10892);
or U18624 (N_18624,N_8156,N_9513);
nor U18625 (N_18625,N_7823,N_10754);
or U18626 (N_18626,N_9091,N_6438);
nand U18627 (N_18627,N_9550,N_12330);
nor U18628 (N_18628,N_7901,N_7232);
or U18629 (N_18629,N_7113,N_7312);
xor U18630 (N_18630,N_7917,N_8660);
nor U18631 (N_18631,N_6312,N_7348);
nor U18632 (N_18632,N_11589,N_6794);
nor U18633 (N_18633,N_7925,N_11339);
xnor U18634 (N_18634,N_12291,N_7687);
and U18635 (N_18635,N_11546,N_7940);
xor U18636 (N_18636,N_9773,N_7778);
nand U18637 (N_18637,N_7461,N_11679);
nor U18638 (N_18638,N_9285,N_12476);
nand U18639 (N_18639,N_12270,N_12082);
or U18640 (N_18640,N_10874,N_11410);
nor U18641 (N_18641,N_9080,N_9414);
xor U18642 (N_18642,N_7871,N_12140);
and U18643 (N_18643,N_8390,N_6652);
or U18644 (N_18644,N_8217,N_7536);
xor U18645 (N_18645,N_10310,N_12292);
nor U18646 (N_18646,N_9534,N_10320);
and U18647 (N_18647,N_9489,N_8726);
and U18648 (N_18648,N_6997,N_9503);
nor U18649 (N_18649,N_8586,N_10653);
and U18650 (N_18650,N_10289,N_9180);
nor U18651 (N_18651,N_7036,N_8478);
xor U18652 (N_18652,N_7366,N_8003);
nor U18653 (N_18653,N_9854,N_9275);
nor U18654 (N_18654,N_7837,N_10076);
or U18655 (N_18655,N_7602,N_6647);
and U18656 (N_18656,N_11867,N_9716);
xor U18657 (N_18657,N_10600,N_10573);
xor U18658 (N_18658,N_12440,N_9338);
nand U18659 (N_18659,N_7684,N_10861);
nor U18660 (N_18660,N_11476,N_10048);
or U18661 (N_18661,N_6820,N_9758);
xor U18662 (N_18662,N_10075,N_11772);
xor U18663 (N_18663,N_12180,N_10149);
nor U18664 (N_18664,N_8528,N_12116);
nor U18665 (N_18665,N_12434,N_9761);
xnor U18666 (N_18666,N_11223,N_8065);
and U18667 (N_18667,N_10771,N_11296);
xnor U18668 (N_18668,N_8022,N_10227);
or U18669 (N_18669,N_10298,N_7868);
nand U18670 (N_18670,N_8158,N_11145);
xor U18671 (N_18671,N_12032,N_7078);
xor U18672 (N_18672,N_11730,N_9864);
or U18673 (N_18673,N_6612,N_6954);
xnor U18674 (N_18674,N_12362,N_6792);
and U18675 (N_18675,N_11948,N_6989);
nor U18676 (N_18676,N_7356,N_7064);
and U18677 (N_18677,N_10806,N_6337);
or U18678 (N_18678,N_12081,N_9978);
nand U18679 (N_18679,N_6753,N_6781);
and U18680 (N_18680,N_7992,N_9259);
xnor U18681 (N_18681,N_11593,N_8700);
nor U18682 (N_18682,N_10406,N_6325);
nand U18683 (N_18683,N_7626,N_6517);
nor U18684 (N_18684,N_8063,N_12490);
or U18685 (N_18685,N_11023,N_9117);
or U18686 (N_18686,N_11542,N_7112);
or U18687 (N_18687,N_6672,N_7476);
and U18688 (N_18688,N_12153,N_6773);
nor U18689 (N_18689,N_12487,N_9556);
and U18690 (N_18690,N_8911,N_8282);
nand U18691 (N_18691,N_10901,N_7469);
or U18692 (N_18692,N_6424,N_7188);
xor U18693 (N_18693,N_10395,N_9842);
nor U18694 (N_18694,N_9405,N_8402);
xnor U18695 (N_18695,N_9987,N_9009);
and U18696 (N_18696,N_6395,N_11827);
nor U18697 (N_18697,N_9894,N_8803);
and U18698 (N_18698,N_11952,N_8732);
nand U18699 (N_18699,N_8668,N_10046);
nand U18700 (N_18700,N_11209,N_12252);
and U18701 (N_18701,N_7492,N_8530);
xnor U18702 (N_18702,N_8658,N_10846);
nand U18703 (N_18703,N_9554,N_7187);
xor U18704 (N_18704,N_11099,N_7746);
or U18705 (N_18705,N_9603,N_11576);
and U18706 (N_18706,N_6741,N_7391);
nor U18707 (N_18707,N_8949,N_8796);
or U18708 (N_18708,N_8097,N_6513);
or U18709 (N_18709,N_8966,N_11160);
xor U18710 (N_18710,N_11824,N_10756);
and U18711 (N_18711,N_6583,N_7833);
or U18712 (N_18712,N_8920,N_10813);
nor U18713 (N_18713,N_9068,N_8391);
nand U18714 (N_18714,N_10816,N_12393);
or U18715 (N_18715,N_10292,N_9601);
nor U18716 (N_18716,N_9677,N_9032);
or U18717 (N_18717,N_10434,N_9906);
xor U18718 (N_18718,N_9119,N_8193);
and U18719 (N_18719,N_8493,N_8014);
nor U18720 (N_18720,N_12410,N_12445);
or U18721 (N_18721,N_7249,N_11075);
nand U18722 (N_18722,N_9219,N_11572);
nor U18723 (N_18723,N_6385,N_11973);
or U18724 (N_18724,N_6605,N_11500);
nand U18725 (N_18725,N_7284,N_9492);
nor U18726 (N_18726,N_6749,N_7074);
nand U18727 (N_18727,N_8880,N_11926);
nor U18728 (N_18728,N_8074,N_10253);
nor U18729 (N_18729,N_6966,N_6910);
nand U18730 (N_18730,N_6455,N_10894);
nand U18731 (N_18731,N_11974,N_11611);
or U18732 (N_18732,N_9783,N_10126);
and U18733 (N_18733,N_11810,N_7674);
or U18734 (N_18734,N_8625,N_6628);
nand U18735 (N_18735,N_11890,N_6387);
or U18736 (N_18736,N_11169,N_12036);
nand U18737 (N_18737,N_10407,N_11328);
xor U18738 (N_18738,N_10674,N_9645);
xor U18739 (N_18739,N_9602,N_7336);
nand U18740 (N_18740,N_8336,N_10918);
nand U18741 (N_18741,N_6748,N_10068);
nand U18742 (N_18742,N_6647,N_7978);
nor U18743 (N_18743,N_9337,N_11848);
and U18744 (N_18744,N_8129,N_9426);
nor U18745 (N_18745,N_9755,N_10687);
and U18746 (N_18746,N_10624,N_8456);
and U18747 (N_18747,N_6908,N_11081);
or U18748 (N_18748,N_10716,N_6935);
and U18749 (N_18749,N_7708,N_10773);
nand U18750 (N_18750,N_12661,N_14744);
xnor U18751 (N_18751,N_16080,N_16225);
nor U18752 (N_18752,N_17505,N_17583);
nor U18753 (N_18753,N_13305,N_16731);
xor U18754 (N_18754,N_18134,N_16082);
nand U18755 (N_18755,N_15690,N_18691);
nor U18756 (N_18756,N_16973,N_16951);
or U18757 (N_18757,N_14764,N_15785);
nand U18758 (N_18758,N_16287,N_16255);
and U18759 (N_18759,N_14199,N_17330);
xor U18760 (N_18760,N_14702,N_15700);
and U18761 (N_18761,N_17300,N_12738);
and U18762 (N_18762,N_14988,N_17510);
and U18763 (N_18763,N_12806,N_16450);
and U18764 (N_18764,N_14382,N_18425);
nand U18765 (N_18765,N_16312,N_15272);
and U18766 (N_18766,N_13877,N_18522);
nand U18767 (N_18767,N_15220,N_14817);
nand U18768 (N_18768,N_18742,N_18566);
and U18769 (N_18769,N_16561,N_17060);
or U18770 (N_18770,N_17142,N_14556);
or U18771 (N_18771,N_18287,N_12531);
nand U18772 (N_18772,N_13430,N_14142);
xor U18773 (N_18773,N_18153,N_17246);
and U18774 (N_18774,N_13842,N_17382);
xor U18775 (N_18775,N_13288,N_15687);
nor U18776 (N_18776,N_15117,N_14624);
or U18777 (N_18777,N_17815,N_16228);
or U18778 (N_18778,N_16308,N_16949);
xor U18779 (N_18779,N_17813,N_14549);
and U18780 (N_18780,N_18587,N_12815);
and U18781 (N_18781,N_16587,N_17355);
nor U18782 (N_18782,N_15850,N_14467);
xnor U18783 (N_18783,N_18491,N_14376);
and U18784 (N_18784,N_13303,N_17974);
nand U18785 (N_18785,N_17597,N_16177);
nand U18786 (N_18786,N_14055,N_17801);
and U18787 (N_18787,N_17908,N_12640);
or U18788 (N_18788,N_15069,N_15842);
or U18789 (N_18789,N_12694,N_15134);
xor U18790 (N_18790,N_16376,N_14745);
nor U18791 (N_18791,N_18389,N_16291);
and U18792 (N_18792,N_15249,N_13289);
nand U18793 (N_18793,N_15759,N_13585);
nor U18794 (N_18794,N_16596,N_13043);
nand U18795 (N_18795,N_18246,N_16000);
nor U18796 (N_18796,N_16551,N_16491);
nor U18797 (N_18797,N_14909,N_13802);
and U18798 (N_18798,N_16845,N_17753);
and U18799 (N_18799,N_18125,N_14471);
and U18800 (N_18800,N_16186,N_12541);
xor U18801 (N_18801,N_16510,N_16410);
nor U18802 (N_18802,N_18527,N_12818);
and U18803 (N_18803,N_17742,N_14163);
or U18804 (N_18804,N_15814,N_16079);
or U18805 (N_18805,N_15379,N_16794);
nand U18806 (N_18806,N_13378,N_13488);
and U18807 (N_18807,N_14875,N_17206);
or U18808 (N_18808,N_16927,N_16547);
xor U18809 (N_18809,N_15870,N_14316);
xor U18810 (N_18810,N_16129,N_13906);
nor U18811 (N_18811,N_16728,N_15277);
xnor U18812 (N_18812,N_17290,N_14168);
or U18813 (N_18813,N_15823,N_16235);
and U18814 (N_18814,N_13092,N_12722);
or U18815 (N_18815,N_13533,N_14816);
or U18816 (N_18816,N_16691,N_15255);
nor U18817 (N_18817,N_17469,N_16555);
nand U18818 (N_18818,N_17244,N_17242);
and U18819 (N_18819,N_13326,N_16636);
nand U18820 (N_18820,N_16517,N_15103);
xnor U18821 (N_18821,N_13479,N_14231);
and U18822 (N_18822,N_15046,N_18734);
or U18823 (N_18823,N_16621,N_18362);
xor U18824 (N_18824,N_13546,N_18336);
or U18825 (N_18825,N_17618,N_16042);
or U18826 (N_18826,N_16207,N_17359);
xnor U18827 (N_18827,N_13205,N_17730);
and U18828 (N_18828,N_12718,N_16374);
nor U18829 (N_18829,N_16464,N_13821);
and U18830 (N_18830,N_17419,N_14511);
nand U18831 (N_18831,N_15080,N_15974);
or U18832 (N_18832,N_16895,N_13087);
xor U18833 (N_18833,N_12515,N_14703);
and U18834 (N_18834,N_15151,N_15705);
xor U18835 (N_18835,N_16124,N_18476);
xor U18836 (N_18836,N_13742,N_16036);
or U18837 (N_18837,N_18732,N_14783);
nor U18838 (N_18838,N_17691,N_13182);
nand U18839 (N_18839,N_14488,N_16777);
or U18840 (N_18840,N_14775,N_14041);
xnor U18841 (N_18841,N_13757,N_17724);
xor U18842 (N_18842,N_18297,N_14874);
and U18843 (N_18843,N_13295,N_18275);
nand U18844 (N_18844,N_14461,N_13299);
or U18845 (N_18845,N_13735,N_13807);
or U18846 (N_18846,N_13006,N_17828);
nor U18847 (N_18847,N_18117,N_18216);
or U18848 (N_18848,N_13148,N_15413);
nand U18849 (N_18849,N_14407,N_16418);
xnor U18850 (N_18850,N_13825,N_18489);
or U18851 (N_18851,N_18310,N_13457);
nand U18852 (N_18852,N_13294,N_13904);
nand U18853 (N_18853,N_15194,N_14265);
nand U18854 (N_18854,N_17091,N_12780);
or U18855 (N_18855,N_17861,N_13948);
nand U18856 (N_18856,N_12849,N_13634);
and U18857 (N_18857,N_13242,N_18159);
nor U18858 (N_18858,N_15939,N_15312);
nor U18859 (N_18859,N_17820,N_15386);
or U18860 (N_18860,N_13130,N_18724);
and U18861 (N_18861,N_18344,N_13373);
nor U18862 (N_18862,N_18409,N_18746);
nor U18863 (N_18863,N_16543,N_17571);
and U18864 (N_18864,N_16759,N_18473);
or U18865 (N_18865,N_17791,N_18552);
nand U18866 (N_18866,N_14321,N_14241);
nand U18867 (N_18867,N_16449,N_13764);
nor U18868 (N_18868,N_16979,N_14155);
and U18869 (N_18869,N_15412,N_13391);
nor U18870 (N_18870,N_15710,N_16836);
or U18871 (N_18871,N_13334,N_18047);
or U18872 (N_18872,N_13139,N_16842);
or U18873 (N_18873,N_13789,N_13893);
or U18874 (N_18874,N_16860,N_15660);
and U18875 (N_18875,N_17090,N_17208);
nand U18876 (N_18876,N_18225,N_18198);
or U18877 (N_18877,N_17825,N_13173);
nand U18878 (N_18878,N_18105,N_16882);
or U18879 (N_18879,N_13985,N_14340);
nand U18880 (N_18880,N_15865,N_16912);
xnor U18881 (N_18881,N_13292,N_14099);
or U18882 (N_18882,N_14635,N_15590);
nor U18883 (N_18883,N_16740,N_13360);
nand U18884 (N_18884,N_15755,N_16157);
nand U18885 (N_18885,N_15498,N_14262);
xor U18886 (N_18886,N_13744,N_12795);
xor U18887 (N_18887,N_13939,N_13409);
and U18888 (N_18888,N_14270,N_13267);
and U18889 (N_18889,N_17320,N_17291);
xor U18890 (N_18890,N_17700,N_13669);
and U18891 (N_18891,N_15706,N_16254);
nand U18892 (N_18892,N_16040,N_16196);
nand U18893 (N_18893,N_18418,N_15915);
and U18894 (N_18894,N_15029,N_17017);
and U18895 (N_18895,N_13860,N_13509);
nand U18896 (N_18896,N_18659,N_17192);
nor U18897 (N_18897,N_16689,N_18033);
xnor U18898 (N_18898,N_17258,N_13829);
xnor U18899 (N_18899,N_12704,N_14539);
or U18900 (N_18900,N_16280,N_15101);
nand U18901 (N_18901,N_15796,N_17444);
nand U18902 (N_18902,N_16874,N_15699);
xnor U18903 (N_18903,N_14620,N_15073);
or U18904 (N_18904,N_14259,N_13154);
xnor U18905 (N_18905,N_13787,N_13178);
xor U18906 (N_18906,N_16747,N_15247);
nand U18907 (N_18907,N_15956,N_18541);
and U18908 (N_18908,N_13121,N_14580);
and U18909 (N_18909,N_17488,N_16957);
nand U18910 (N_18910,N_18594,N_18030);
nand U18911 (N_18911,N_15256,N_14885);
xnor U18912 (N_18912,N_13819,N_18632);
xor U18913 (N_18913,N_15817,N_15780);
and U18914 (N_18914,N_17857,N_12526);
nor U18915 (N_18915,N_16578,N_17920);
or U18916 (N_18916,N_16574,N_14147);
xnor U18917 (N_18917,N_16294,N_12544);
or U18918 (N_18918,N_13311,N_16674);
nand U18919 (N_18919,N_14169,N_15455);
nor U18920 (N_18920,N_15716,N_14548);
nor U18921 (N_18921,N_18100,N_14111);
xor U18922 (N_18922,N_15535,N_15553);
xor U18923 (N_18923,N_15173,N_16875);
nand U18924 (N_18924,N_15869,N_17153);
and U18925 (N_18925,N_17454,N_13019);
nor U18926 (N_18926,N_13915,N_16852);
or U18927 (N_18927,N_13986,N_16813);
nand U18928 (N_18928,N_18689,N_13082);
nor U18929 (N_18929,N_15131,N_14158);
and U18930 (N_18930,N_14327,N_16765);
nand U18931 (N_18931,N_15383,N_13711);
nand U18932 (N_18932,N_14929,N_14748);
nand U18933 (N_18933,N_15343,N_16401);
nor U18934 (N_18934,N_16286,N_13371);
nand U18935 (N_18935,N_18382,N_17869);
and U18936 (N_18936,N_14081,N_15375);
xor U18937 (N_18937,N_17097,N_17521);
or U18938 (N_18938,N_18472,N_12508);
nor U18939 (N_18939,N_16370,N_13772);
and U18940 (N_18940,N_14489,N_14389);
nand U18941 (N_18941,N_16851,N_15799);
nor U18942 (N_18942,N_13515,N_17538);
xnor U18943 (N_18943,N_18373,N_12735);
and U18944 (N_18944,N_15691,N_16965);
xnor U18945 (N_18945,N_14989,N_12645);
nor U18946 (N_18946,N_15283,N_15506);
or U18947 (N_18947,N_13249,N_16353);
nor U18948 (N_18948,N_18682,N_14678);
xnor U18949 (N_18949,N_12622,N_14667);
or U18950 (N_18950,N_17081,N_13912);
and U18951 (N_18951,N_14789,N_16393);
nor U18952 (N_18952,N_16397,N_16382);
nand U18953 (N_18953,N_17342,N_17442);
xor U18954 (N_18954,N_17580,N_16609);
and U18955 (N_18955,N_14812,N_18678);
nor U18956 (N_18956,N_13049,N_15172);
or U18957 (N_18957,N_13762,N_18096);
or U18958 (N_18958,N_17564,N_15100);
or U18959 (N_18959,N_18116,N_15421);
nand U18960 (N_18960,N_16654,N_15952);
and U18961 (N_18961,N_12561,N_17685);
nor U18962 (N_18962,N_17032,N_16900);
nand U18963 (N_18963,N_15653,N_14979);
xor U18964 (N_18964,N_14519,N_16429);
or U18965 (N_18965,N_15463,N_12896);
nand U18966 (N_18966,N_13574,N_15568);
or U18967 (N_18967,N_14639,N_13489);
nand U18968 (N_18968,N_17709,N_15384);
and U18969 (N_18969,N_16829,N_18158);
and U18970 (N_18970,N_13959,N_15711);
nor U18971 (N_18971,N_17111,N_16901);
xor U18972 (N_18972,N_16527,N_15005);
or U18973 (N_18973,N_13203,N_14257);
xor U18974 (N_18974,N_12742,N_16877);
and U18975 (N_18975,N_16679,N_15563);
and U18976 (N_18976,N_13387,N_13962);
or U18977 (N_18977,N_18625,N_17862);
nand U18978 (N_18978,N_18679,N_13075);
nor U18979 (N_18979,N_13933,N_12554);
nand U18980 (N_18980,N_14757,N_18380);
or U18981 (N_18981,N_16172,N_13608);
nand U18982 (N_18982,N_18048,N_15536);
nand U18983 (N_18983,N_14857,N_15825);
or U18984 (N_18984,N_15887,N_15564);
nor U18985 (N_18985,N_18079,N_15457);
xnor U18986 (N_18986,N_13027,N_17399);
nand U18987 (N_18987,N_13238,N_13171);
xor U18988 (N_18988,N_14223,N_12506);
or U18989 (N_18989,N_13200,N_12709);
or U18990 (N_18990,N_17842,N_13197);
nor U18991 (N_18991,N_16320,N_15390);
and U18992 (N_18992,N_17392,N_13251);
xnor U18993 (N_18993,N_15736,N_13481);
xor U18994 (N_18994,N_16017,N_13752);
nand U18995 (N_18995,N_13706,N_18621);
nand U18996 (N_18996,N_14936,N_16760);
or U18997 (N_18997,N_16126,N_15133);
nand U18998 (N_18998,N_17752,N_13918);
xor U18999 (N_18999,N_17257,N_14114);
nor U19000 (N_19000,N_17340,N_15589);
or U19001 (N_19001,N_14436,N_13362);
or U19002 (N_19002,N_16701,N_12825);
or U19003 (N_19003,N_14798,N_18411);
xor U19004 (N_19004,N_12741,N_17123);
or U19005 (N_19005,N_17031,N_16662);
xor U19006 (N_19006,N_17174,N_14387);
and U19007 (N_19007,N_16425,N_15023);
nor U19008 (N_19008,N_16106,N_16583);
nor U19009 (N_19009,N_16642,N_17150);
or U19010 (N_19010,N_18169,N_13559);
nand U19011 (N_19011,N_16919,N_13452);
or U19012 (N_19012,N_13721,N_16170);
nand U19013 (N_19013,N_17947,N_15257);
nand U19014 (N_19014,N_16810,N_14189);
and U19015 (N_19015,N_13547,N_13313);
nor U19016 (N_19016,N_18662,N_13282);
xor U19017 (N_19017,N_17457,N_14933);
and U19018 (N_19018,N_18213,N_13624);
xnor U19019 (N_19019,N_13134,N_15862);
nand U19020 (N_19020,N_14584,N_15414);
and U19021 (N_19021,N_14156,N_15104);
nor U19022 (N_19022,N_14213,N_16730);
or U19023 (N_19023,N_18284,N_16092);
nand U19024 (N_19024,N_16439,N_16824);
nor U19025 (N_19025,N_13275,N_12611);
nor U19026 (N_19026,N_15372,N_14476);
xor U19027 (N_19027,N_17575,N_17059);
nor U19028 (N_19028,N_18049,N_13045);
or U19029 (N_19029,N_15357,N_14289);
nand U19030 (N_19030,N_12983,N_15578);
and U19031 (N_19031,N_17973,N_14131);
nor U19032 (N_19032,N_16763,N_15374);
or U19033 (N_19033,N_16745,N_16929);
nand U19034 (N_19034,N_14229,N_14473);
xnor U19035 (N_19035,N_12677,N_16270);
nor U19036 (N_19036,N_14709,N_14513);
nor U19037 (N_19037,N_16078,N_17196);
or U19038 (N_19038,N_13320,N_14557);
nand U19039 (N_19039,N_14239,N_12650);
or U19040 (N_19040,N_13977,N_16379);
nand U19041 (N_19041,N_15694,N_13616);
or U19042 (N_19042,N_15943,N_18528);
nand U19043 (N_19043,N_15062,N_12823);
and U19044 (N_19044,N_15895,N_15920);
nor U19045 (N_19045,N_12601,N_18328);
or U19046 (N_19046,N_13982,N_17911);
or U19047 (N_19047,N_15926,N_18077);
xnor U19048 (N_19048,N_13385,N_15561);
nand U19049 (N_19049,N_14258,N_13435);
xor U19050 (N_19050,N_16098,N_13351);
xnor U19051 (N_19051,N_16210,N_17903);
nor U19052 (N_19052,N_15505,N_13582);
or U19053 (N_19053,N_18186,N_12652);
nor U19054 (N_19054,N_13109,N_14809);
nand U19055 (N_19055,N_16061,N_13052);
nor U19056 (N_19056,N_18540,N_18633);
nor U19057 (N_19057,N_18504,N_14425);
nand U19058 (N_19058,N_17212,N_15471);
or U19059 (N_19059,N_18230,N_13403);
xnor U19060 (N_19060,N_12909,N_12789);
xnor U19061 (N_19061,N_17369,N_14947);
xnor U19062 (N_19062,N_15155,N_16970);
nand U19063 (N_19063,N_12770,N_15972);
xor U19064 (N_19064,N_17054,N_12636);
nor U19065 (N_19065,N_17231,N_17058);
nand U19066 (N_19066,N_13357,N_17967);
xor U19067 (N_19067,N_14713,N_16028);
xor U19068 (N_19068,N_18239,N_13639);
nand U19069 (N_19069,N_14255,N_13302);
nor U19070 (N_19070,N_13554,N_15917);
and U19071 (N_19071,N_12835,N_17020);
xor U19072 (N_19072,N_13895,N_12919);
and U19073 (N_19073,N_14707,N_13796);
or U19074 (N_19074,N_16703,N_15701);
or U19075 (N_19075,N_13503,N_13332);
xnor U19076 (N_19076,N_13529,N_14882);
and U19077 (N_19077,N_16651,N_17249);
and U19078 (N_19078,N_17494,N_16469);
xnor U19079 (N_19079,N_13964,N_13217);
or U19080 (N_19080,N_13056,N_12688);
and U19081 (N_19081,N_15108,N_16195);
xor U19082 (N_19082,N_17535,N_13650);
nor U19083 (N_19083,N_17837,N_16297);
or U19084 (N_19084,N_13186,N_15159);
nor U19085 (N_19085,N_14996,N_18251);
xnor U19086 (N_19086,N_12692,N_17190);
nand U19087 (N_19087,N_18684,N_18747);
xnor U19088 (N_19088,N_16476,N_15669);
nand U19089 (N_19089,N_15222,N_16190);
nor U19090 (N_19090,N_13972,N_13415);
xnor U19091 (N_19091,N_14522,N_12755);
and U19092 (N_19092,N_16735,N_16946);
and U19093 (N_19093,N_18267,N_16067);
and U19094 (N_19094,N_16342,N_18645);
xor U19095 (N_19095,N_17210,N_13505);
nor U19096 (N_19096,N_18130,N_15734);
nand U19097 (N_19097,N_17542,N_18417);
or U19098 (N_19098,N_13507,N_15233);
and U19099 (N_19099,N_15775,N_16584);
and U19100 (N_19100,N_14818,N_14881);
nand U19101 (N_19101,N_17871,N_16071);
nor U19102 (N_19102,N_15617,N_17586);
and U19103 (N_19103,N_17034,N_15309);
or U19104 (N_19104,N_16980,N_13621);
nand U19105 (N_19105,N_18238,N_18347);
xnor U19106 (N_19106,N_14483,N_14333);
nand U19107 (N_19107,N_18748,N_16140);
and U19108 (N_19108,N_16634,N_12679);
and U19109 (N_19109,N_16309,N_14330);
or U19110 (N_19110,N_13617,N_17805);
or U19111 (N_19111,N_15906,N_16127);
or U19112 (N_19112,N_16546,N_14866);
and U19113 (N_19113,N_17131,N_16554);
or U19114 (N_19114,N_12591,N_15400);
nand U19115 (N_19115,N_17958,N_14706);
nand U19116 (N_19116,N_17506,N_18143);
and U19117 (N_19117,N_15241,N_16683);
nor U19118 (N_19118,N_13455,N_15748);
and U19119 (N_19119,N_18636,N_18385);
nor U19120 (N_19120,N_14445,N_12890);
nor U19121 (N_19121,N_17572,N_14569);
or U19122 (N_19122,N_12588,N_15431);
xor U19123 (N_19123,N_15575,N_17205);
and U19124 (N_19124,N_15707,N_12997);
nor U19125 (N_19125,N_14191,N_13601);
nand U19126 (N_19126,N_14373,N_13036);
nand U19127 (N_19127,N_17600,N_18334);
and U19128 (N_19128,N_15962,N_16793);
and U19129 (N_19129,N_17439,N_13865);
xor U19130 (N_19130,N_18149,N_17026);
nand U19131 (N_19131,N_17325,N_18114);
xnor U19132 (N_19132,N_17721,N_13792);
xnor U19133 (N_19133,N_13717,N_13176);
or U19134 (N_19134,N_17484,N_14814);
xor U19135 (N_19135,N_16589,N_14284);
nand U19136 (N_19136,N_15427,N_17405);
or U19137 (N_19137,N_12627,N_12733);
nor U19138 (N_19138,N_13395,N_14849);
or U19139 (N_19139,N_15114,N_14883);
or U19140 (N_19140,N_13324,N_15064);
nor U19141 (N_19141,N_16620,N_17536);
nor U19142 (N_19142,N_14365,N_13284);
nor U19143 (N_19143,N_16688,N_12926);
nand U19144 (N_19144,N_18412,N_15976);
nor U19145 (N_19145,N_16166,N_16440);
nor U19146 (N_19146,N_12558,N_16118);
and U19147 (N_19147,N_17634,N_16566);
xnor U19148 (N_19148,N_15338,N_15628);
xnor U19149 (N_19149,N_14171,N_17066);
nor U19150 (N_19150,N_12880,N_15719);
nand U19151 (N_19151,N_15349,N_13279);
nand U19152 (N_19152,N_15299,N_13566);
and U19153 (N_19153,N_18383,N_16452);
and U19154 (N_19154,N_13485,N_12740);
xor U19155 (N_19155,N_13048,N_18535);
nor U19156 (N_19156,N_18580,N_16511);
nand U19157 (N_19157,N_14691,N_12595);
xor U19158 (N_19158,N_12839,N_12758);
nand U19159 (N_19159,N_13118,N_15878);
xnor U19160 (N_19160,N_18217,N_15264);
xor U19161 (N_19161,N_13607,N_12528);
xor U19162 (N_19162,N_14723,N_12571);
and U19163 (N_19163,N_15199,N_13994);
xor U19164 (N_19164,N_12563,N_18008);
nor U19165 (N_19165,N_17686,N_16378);
nand U19166 (N_19166,N_12821,N_12503);
nor U19167 (N_19167,N_16884,N_15336);
xnor U19168 (N_19168,N_13304,N_13946);
nor U19169 (N_19169,N_18578,N_12986);
xor U19170 (N_19170,N_15683,N_18027);
or U19171 (N_19171,N_18223,N_16076);
or U19172 (N_19172,N_17012,N_15541);
and U19173 (N_19173,N_13780,N_13552);
nand U19174 (N_19174,N_16560,N_17327);
and U19175 (N_19175,N_14220,N_18459);
nand U19176 (N_19176,N_13543,N_18591);
xnor U19177 (N_19177,N_15684,N_14045);
or U19178 (N_19178,N_18052,N_17492);
and U19179 (N_19179,N_18196,N_17978);
and U19180 (N_19180,N_13663,N_17447);
nor U19181 (N_19181,N_18352,N_14064);
or U19182 (N_19182,N_15833,N_15032);
nand U19183 (N_19183,N_13416,N_12930);
xor U19184 (N_19184,N_18556,N_15362);
xor U19185 (N_19185,N_13085,N_13308);
xor U19186 (N_19186,N_16796,N_17874);
nor U19187 (N_19187,N_17448,N_15467);
nor U19188 (N_19188,N_14182,N_16323);
or U19189 (N_19189,N_17671,N_13243);
or U19190 (N_19190,N_14767,N_15737);
xnor U19191 (N_19191,N_16215,N_17397);
nand U19192 (N_19192,N_16671,N_13545);
and U19193 (N_19193,N_13011,N_13595);
or U19194 (N_19194,N_16250,N_12917);
or U19195 (N_19195,N_18257,N_17799);
xor U19196 (N_19196,N_12946,N_16428);
nand U19197 (N_19197,N_16485,N_18062);
or U19198 (N_19198,N_13224,N_17158);
or U19199 (N_19199,N_15688,N_17140);
nand U19200 (N_19200,N_14640,N_18260);
xor U19201 (N_19201,N_14560,N_17648);
and U19202 (N_19202,N_12572,N_12727);
nor U19203 (N_19203,N_15677,N_15530);
and U19204 (N_19204,N_13928,N_13594);
and U19205 (N_19205,N_17170,N_18087);
nor U19206 (N_19206,N_16271,N_17228);
xnor U19207 (N_19207,N_17687,N_16015);
or U19208 (N_19208,N_12646,N_17339);
or U19209 (N_19209,N_14253,N_16849);
or U19210 (N_19210,N_13323,N_16976);
and U19211 (N_19211,N_14423,N_18075);
nor U19212 (N_19212,N_17764,N_13705);
and U19213 (N_19213,N_12974,N_12728);
nand U19214 (N_19214,N_15847,N_13494);
nand U19215 (N_19215,N_15116,N_16360);
or U19216 (N_19216,N_13809,N_16776);
nand U19217 (N_19217,N_16841,N_15063);
xor U19218 (N_19218,N_13530,N_17818);
or U19219 (N_19219,N_17311,N_13888);
nand U19220 (N_19220,N_15528,N_18650);
nand U19221 (N_19221,N_18692,N_17627);
nor U19222 (N_19222,N_15866,N_17723);
nor U19223 (N_19223,N_14617,N_16152);
or U19224 (N_19224,N_14546,N_14503);
and U19225 (N_19225,N_13033,N_13953);
and U19226 (N_19226,N_18563,N_16497);
nor U19227 (N_19227,N_17582,N_14932);
nor U19228 (N_19228,N_15950,N_18168);
nor U19229 (N_19229,N_18111,N_17269);
nand U19230 (N_19230,N_17446,N_13723);
or U19231 (N_19231,N_17476,N_18124);
or U19232 (N_19232,N_14224,N_16415);
xnor U19233 (N_19233,N_16736,N_18640);
and U19234 (N_19234,N_17649,N_15610);
and U19235 (N_19235,N_18513,N_16542);
nor U19236 (N_19236,N_13141,N_14235);
nor U19237 (N_19237,N_16212,N_14611);
nor U19238 (N_19238,N_13472,N_12540);
xor U19239 (N_19239,N_12786,N_17534);
nor U19240 (N_19240,N_16381,N_14899);
and U19241 (N_19241,N_17643,N_14102);
xor U19242 (N_19242,N_14338,N_12502);
nor U19243 (N_19243,N_15472,N_15794);
or U19244 (N_19244,N_16831,N_15411);
and U19245 (N_19245,N_18082,N_17255);
nand U19246 (N_19246,N_18144,N_13907);
and U19247 (N_19247,N_13336,N_15788);
and U19248 (N_19248,N_13655,N_14810);
and U19249 (N_19249,N_18210,N_14065);
and U19250 (N_19250,N_14090,N_18097);
nor U19251 (N_19251,N_17201,N_17356);
nand U19252 (N_19252,N_14559,N_16661);
nor U19253 (N_19253,N_14700,N_15355);
nand U19254 (N_19254,N_15315,N_17126);
and U19255 (N_19255,N_16515,N_15028);
nand U19256 (N_19256,N_18067,N_14370);
xor U19257 (N_19257,N_16508,N_17647);
or U19258 (N_19258,N_14161,N_14558);
and U19259 (N_19259,N_17578,N_12803);
nor U19260 (N_19260,N_14962,N_14344);
xnor U19261 (N_19261,N_17599,N_14037);
or U19262 (N_19262,N_13880,N_15370);
or U19263 (N_19263,N_12523,N_15981);
nand U19264 (N_19264,N_16887,N_16607);
nor U19265 (N_19265,N_16380,N_15227);
nand U19266 (N_19266,N_18333,N_16402);
and U19267 (N_19267,N_13136,N_13031);
nor U19268 (N_19268,N_14832,N_15809);
and U19269 (N_19269,N_17470,N_15876);
xor U19270 (N_19270,N_14547,N_14508);
or U19271 (N_19271,N_15948,N_17921);
nand U19272 (N_19272,N_17577,N_16663);
or U19273 (N_19273,N_14015,N_17675);
nor U19274 (N_19274,N_14804,N_17239);
nor U19275 (N_19275,N_12576,N_17553);
nor U19276 (N_19276,N_14915,N_18278);
nor U19277 (N_19277,N_14658,N_15109);
and U19278 (N_19278,N_17778,N_13874);
nor U19279 (N_19279,N_18113,N_13152);
and U19280 (N_19280,N_13795,N_15686);
nor U19281 (N_19281,N_17986,N_12536);
or U19282 (N_19282,N_15006,N_16245);
nor U19283 (N_19283,N_18646,N_15096);
nand U19284 (N_19284,N_17133,N_12855);
xor U19285 (N_19285,N_12841,N_15793);
xnor U19286 (N_19286,N_12509,N_18235);
nand U19287 (N_19287,N_13908,N_12979);
xnor U19288 (N_19288,N_13042,N_12912);
nor U19289 (N_19289,N_13719,N_15250);
and U19290 (N_19290,N_17800,N_15650);
nor U19291 (N_19291,N_13555,N_14564);
nand U19292 (N_19292,N_14762,N_16790);
nand U19293 (N_19293,N_16311,N_17194);
or U19294 (N_19294,N_12959,N_13233);
nor U19295 (N_19295,N_13088,N_13382);
nand U19296 (N_19296,N_14146,N_13438);
or U19297 (N_19297,N_16459,N_13140);
or U19298 (N_19298,N_14346,N_16339);
and U19299 (N_19299,N_17107,N_15461);
nand U19300 (N_19300,N_13414,N_18330);
xor U19301 (N_19301,N_14778,N_17016);
nor U19302 (N_19302,N_18693,N_16183);
nand U19303 (N_19303,N_16302,N_14132);
xor U19304 (N_19304,N_13040,N_12982);
and U19305 (N_19305,N_16009,N_15864);
or U19306 (N_19306,N_17219,N_12724);
nand U19307 (N_19307,N_14429,N_14368);
and U19308 (N_19308,N_16644,N_16426);
nor U19309 (N_19309,N_16012,N_16417);
nor U19310 (N_19310,N_13408,N_16395);
or U19311 (N_19311,N_12649,N_14834);
or U19312 (N_19312,N_16928,N_13029);
or U19313 (N_19313,N_17424,N_15758);
xor U19314 (N_19314,N_12899,N_17297);
xor U19315 (N_19315,N_18601,N_17179);
nor U19316 (N_19316,N_14317,N_14103);
xnor U19317 (N_19317,N_13638,N_18437);
xnor U19318 (N_19318,N_18604,N_14714);
nor U19319 (N_19319,N_13722,N_14543);
nor U19320 (N_19320,N_18256,N_18658);
xnor U19321 (N_19321,N_16633,N_14502);
xnor U19322 (N_19322,N_15821,N_16984);
or U19323 (N_19323,N_16966,N_16138);
and U19324 (N_19324,N_16160,N_17462);
xor U19325 (N_19325,N_17819,N_15652);
or U19326 (N_19326,N_13673,N_16692);
and U19327 (N_19327,N_13469,N_15989);
nand U19328 (N_19328,N_16502,N_13064);
or U19329 (N_19329,N_17357,N_18064);
or U19330 (N_19330,N_13593,N_15416);
xnor U19331 (N_19331,N_13331,N_13235);
xor U19332 (N_19332,N_15061,N_14821);
xnor U19333 (N_19333,N_14492,N_13526);
or U19334 (N_19334,N_13256,N_12666);
or U19335 (N_19335,N_15351,N_15176);
nor U19336 (N_19336,N_14731,N_18183);
or U19337 (N_19337,N_13114,N_14104);
nand U19338 (N_19338,N_16289,N_14016);
or U19339 (N_19339,N_18146,N_13445);
or U19340 (N_19340,N_16338,N_14997);
and U19341 (N_19341,N_17240,N_15945);
or U19342 (N_19342,N_17427,N_18317);
nor U19343 (N_19343,N_17692,N_18652);
nand U19344 (N_19344,N_12964,N_15102);
nor U19345 (N_19345,N_16182,N_13597);
or U19346 (N_19346,N_12977,N_16941);
and U19347 (N_19347,N_14763,N_12701);
nand U19348 (N_19348,N_13606,N_14615);
nand U19349 (N_19349,N_16390,N_16767);
xnor U19350 (N_19350,N_15018,N_16333);
xor U19351 (N_19351,N_18674,N_18629);
or U19352 (N_19352,N_13710,N_14772);
and U19353 (N_19353,N_14602,N_16635);
nor U19354 (N_19354,N_12861,N_17585);
and U19355 (N_19355,N_15486,N_12639);
or U19356 (N_19356,N_17930,N_18712);
nor U19357 (N_19357,N_15562,N_15086);
or U19358 (N_19358,N_18253,N_18228);
nand U19359 (N_19359,N_18005,N_13724);
and U19360 (N_19360,N_13851,N_15066);
nor U19361 (N_19361,N_18057,N_14324);
nor U19362 (N_19362,N_14073,N_14251);
xnor U19363 (N_19363,N_13812,N_14180);
xnor U19364 (N_19364,N_16606,N_15293);
and U19365 (N_19365,N_13262,N_17475);
nand U19366 (N_19366,N_15129,N_18307);
nand U19367 (N_19367,N_12597,N_14341);
and U19368 (N_19368,N_14009,N_17898);
nand U19369 (N_19369,N_14674,N_16154);
nand U19370 (N_19370,N_14059,N_14035);
nor U19371 (N_19371,N_13831,N_15881);
nor U19372 (N_19372,N_18593,N_15958);
and U19373 (N_19373,N_16773,N_18557);
or U19374 (N_19374,N_16306,N_15285);
and U19375 (N_19375,N_17659,N_14946);
xnor U19376 (N_19376,N_17347,N_15678);
or U19377 (N_19377,N_17948,N_15534);
nor U19378 (N_19378,N_18400,N_18306);
or U19379 (N_19379,N_14271,N_18714);
and U19380 (N_19380,N_13935,N_14401);
and U19381 (N_19381,N_14299,N_17332);
and U19382 (N_19382,N_18635,N_18526);
and U19383 (N_19383,N_14733,N_13799);
or U19384 (N_19384,N_13798,N_15037);
nand U19385 (N_19385,N_15767,N_13189);
and U19386 (N_19386,N_12586,N_18607);
or U19387 (N_19387,N_13390,N_12857);
and U19388 (N_19388,N_12555,N_13017);
or U19389 (N_19389,N_18368,N_14150);
nand U19390 (N_19390,N_14970,N_13063);
nor U19391 (N_19391,N_18584,N_14138);
or U19392 (N_19392,N_12577,N_15326);
or U19393 (N_19393,N_17633,N_14441);
or U19394 (N_19394,N_15296,N_16359);
nor U19395 (N_19395,N_18280,N_12587);
xnor U19396 (N_19396,N_17189,N_13979);
nand U19397 (N_19397,N_14388,N_16617);
and U19398 (N_19398,N_17005,N_13818);
and U19399 (N_19399,N_16048,N_15404);
xnor U19400 (N_19400,N_15648,N_17626);
nor U19401 (N_19401,N_15844,N_18208);
xor U19402 (N_19402,N_18500,N_15871);
and U19403 (N_19403,N_12657,N_16670);
xnor U19404 (N_19404,N_17729,N_12734);
nor U19405 (N_19405,N_16463,N_16164);
nand U19406 (N_19406,N_13832,N_15499);
xnor U19407 (N_19407,N_13811,N_12749);
nand U19408 (N_19408,N_18061,N_14957);
nor U19409 (N_19409,N_15666,N_14805);
xor U19410 (N_19410,N_18749,N_14018);
nand U19411 (N_19411,N_15604,N_13884);
xnor U19412 (N_19412,N_18314,N_17949);
or U19413 (N_19413,N_16724,N_17363);
xnor U19414 (N_19414,N_13751,N_12767);
xor U19415 (N_19415,N_13718,N_17410);
xor U19416 (N_19416,N_16897,N_13855);
xor U19417 (N_19417,N_17983,N_17784);
nor U19418 (N_19418,N_17048,N_12744);
xor U19419 (N_19419,N_12864,N_13779);
xor U19420 (N_19420,N_14968,N_17316);
nor U19421 (N_19421,N_13450,N_15317);
and U19422 (N_19422,N_17855,N_13328);
nor U19423 (N_19423,N_14083,N_13454);
or U19424 (N_19424,N_15637,N_15373);
nand U19425 (N_19425,N_13836,N_16603);
and U19426 (N_19426,N_18441,N_18147);
nor U19427 (N_19427,N_17102,N_12972);
or U19428 (N_19428,N_16865,N_14826);
and U19429 (N_19429,N_14001,N_13000);
or U19430 (N_19430,N_15508,N_14485);
xnor U19431 (N_19431,N_14204,N_16577);
or U19432 (N_19432,N_12761,N_16404);
nor U19433 (N_19433,N_16480,N_15601);
and U19434 (N_19434,N_14893,N_13519);
nor U19435 (N_19435,N_13456,N_14948);
xnor U19436 (N_19436,N_16820,N_12893);
nand U19437 (N_19437,N_13212,N_14390);
or U19438 (N_19438,N_16142,N_18525);
nor U19439 (N_19439,N_18243,N_14486);
or U19440 (N_19440,N_12578,N_16041);
nand U19441 (N_19441,N_15803,N_18657);
xnor U19442 (N_19442,N_17843,N_18354);
nor U19443 (N_19443,N_13406,N_12916);
or U19444 (N_19444,N_18053,N_16815);
and U19445 (N_19445,N_14005,N_13398);
nand U19446 (N_19446,N_12796,N_16677);
nor U19447 (N_19447,N_18366,N_14943);
nor U19448 (N_19448,N_14236,N_15090);
and U19449 (N_19449,N_13388,N_14019);
or U19450 (N_19450,N_17824,N_15165);
or U19451 (N_19451,N_15420,N_17501);
nor U19452 (N_19452,N_15656,N_15524);
xnor U19453 (N_19453,N_15550,N_17846);
xnor U19454 (N_19454,N_13206,N_16066);
xor U19455 (N_19455,N_17341,N_12765);
nor U19456 (N_19456,N_17420,N_18126);
and U19457 (N_19457,N_16614,N_12989);
and U19458 (N_19458,N_15837,N_18568);
xor U19459 (N_19459,N_18236,N_17039);
nand U19460 (N_19460,N_16343,N_15447);
nand U19461 (N_19461,N_14124,N_13968);
nor U19462 (N_19462,N_18731,N_12984);
nand U19463 (N_19463,N_15070,N_16423);
nand U19464 (N_19464,N_15845,N_13321);
xor U19465 (N_19465,N_18145,N_16335);
and U19466 (N_19466,N_15475,N_14985);
nor U19467 (N_19467,N_15921,N_13346);
and U19468 (N_19468,N_18537,N_16605);
or U19469 (N_19469,N_14438,N_12676);
or U19470 (N_19470,N_14550,N_13591);
nand U19471 (N_19471,N_14054,N_14243);
and U19472 (N_19472,N_15964,N_17881);
nor U19473 (N_19473,N_16026,N_16403);
and U19474 (N_19474,N_15797,N_17227);
or U19475 (N_19475,N_18439,N_13670);
xnor U19476 (N_19476,N_17902,N_14369);
xnor U19477 (N_19477,N_14004,N_14266);
xor U19478 (N_19478,N_15135,N_13892);
nor U19479 (N_19479,N_13493,N_17605);
nand U19480 (N_19480,N_18739,N_18327);
nor U19481 (N_19481,N_16285,N_13263);
nor U19482 (N_19482,N_17071,N_13848);
and U19483 (N_19483,N_13666,N_13990);
xnor U19484 (N_19484,N_15880,N_12863);
nor U19485 (N_19485,N_12871,N_15197);
or U19486 (N_19486,N_17472,N_16111);
xnor U19487 (N_19487,N_14588,N_16902);
nand U19488 (N_19488,N_15497,N_14515);
or U19489 (N_19489,N_14276,N_13782);
xor U19490 (N_19490,N_14926,N_17830);
nand U19491 (N_19491,N_17714,N_16969);
nand U19492 (N_19492,N_16065,N_12543);
or U19493 (N_19493,N_15019,N_14607);
xnor U19494 (N_19494,N_18505,N_15609);
nand U19495 (N_19495,N_15662,N_16771);
xnor U19496 (N_19496,N_15787,N_16103);
nor U19497 (N_19497,N_14753,N_17217);
xnor U19498 (N_19498,N_15462,N_16322);
xnor U19499 (N_19499,N_18606,N_13147);
xor U19500 (N_19500,N_16037,N_12801);
nor U19501 (N_19501,N_16305,N_14087);
or U19502 (N_19502,N_14653,N_16668);
nor U19503 (N_19503,N_15640,N_15522);
xnor U19504 (N_19504,N_18219,N_13604);
xnor U19505 (N_19505,N_18074,N_15305);
xnor U19506 (N_19506,N_12775,N_15994);
nor U19507 (N_19507,N_13866,N_17285);
and U19508 (N_19508,N_16173,N_13372);
nand U19509 (N_19509,N_18583,N_16447);
xnor U19510 (N_19510,N_14465,N_17337);
xor U19511 (N_19511,N_13883,N_15205);
nor U19512 (N_19512,N_14527,N_16385);
nor U19513 (N_19513,N_17028,N_16650);
nor U19514 (N_19514,N_13658,N_13930);
and U19515 (N_19515,N_13815,N_13891);
or U19516 (N_19516,N_14208,N_17321);
nor U19517 (N_19517,N_18542,N_13844);
xnor U19518 (N_19518,N_18157,N_15052);
and U19519 (N_19519,N_12532,N_18506);
xor U19520 (N_19520,N_12908,N_13736);
and U19521 (N_19521,N_14201,N_15314);
or U19522 (N_19522,N_16224,N_16952);
and U19523 (N_19523,N_12620,N_13333);
xnor U19524 (N_19524,N_16413,N_17877);
nor U19525 (N_19525,N_18653,N_18022);
xnor U19526 (N_19526,N_18665,N_16131);
nor U19527 (N_19527,N_14612,N_14434);
nand U19528 (N_19528,N_17080,N_18534);
nand U19529 (N_19529,N_17412,N_13433);
xor U19530 (N_19530,N_14518,N_14118);
nand U19531 (N_19531,N_15094,N_15860);
and U19532 (N_19532,N_14914,N_17411);
nor U19533 (N_19533,N_12799,N_15565);
nor U19534 (N_19534,N_16907,N_18449);
xnor U19535 (N_19535,N_13854,N_12606);
and U19536 (N_19536,N_16181,N_13486);
nor U19537 (N_19537,N_12746,N_17765);
xnor U19538 (N_19538,N_17707,N_14795);
xor U19539 (N_19539,N_15012,N_18545);
xnor U19540 (N_19540,N_17587,N_17072);
xnor U19541 (N_19541,N_13689,N_16732);
nand U19542 (N_19542,N_17408,N_12790);
and U19543 (N_19543,N_17566,N_14935);
nand U19544 (N_19544,N_15681,N_18670);
nand U19545 (N_19545,N_13680,N_12872);
nor U19546 (N_19546,N_13426,N_18735);
nand U19547 (N_19547,N_13225,N_15083);
or U19548 (N_19548,N_13869,N_14911);
or U19549 (N_19549,N_15181,N_12826);
nor U19550 (N_19550,N_13648,N_13247);
or U19551 (N_19551,N_13688,N_13380);
xor U19552 (N_19552,N_18581,N_17343);
or U19553 (N_19553,N_16623,N_16582);
xnor U19554 (N_19554,N_12697,N_14586);
or U19555 (N_19555,N_17460,N_17416);
and U19556 (N_19556,N_15896,N_14673);
nor U19557 (N_19557,N_16005,N_13028);
or U19558 (N_19558,N_18432,N_14153);
and U19559 (N_19559,N_12547,N_13358);
xor U19560 (N_19560,N_17909,N_16593);
or U19561 (N_19561,N_15680,N_18374);
nand U19562 (N_19562,N_14600,N_17944);
and U19563 (N_19563,N_18184,N_15358);
nand U19564 (N_19564,N_12764,N_13227);
nand U19565 (N_19565,N_13644,N_13327);
or U19566 (N_19566,N_14836,N_17745);
xnor U19567 (N_19567,N_17811,N_13053);
nor U19568 (N_19568,N_18560,N_14773);
or U19569 (N_19569,N_16315,N_13571);
and U19570 (N_19570,N_18544,N_12949);
and U19571 (N_19571,N_13352,N_15231);
or U19572 (N_19572,N_12980,N_14443);
xnor U19573 (N_19573,N_17502,N_13786);
nor U19574 (N_19574,N_13693,N_15477);
nand U19575 (N_19575,N_16242,N_14475);
or U19576 (N_19576,N_16389,N_15933);
or U19577 (N_19577,N_16367,N_18553);
and U19578 (N_19578,N_14941,N_15572);
xor U19579 (N_19579,N_16371,N_13468);
nor U19580 (N_19580,N_16693,N_16500);
nand U19581 (N_19581,N_12811,N_16214);
nand U19582 (N_19582,N_17867,N_12665);
xnor U19583 (N_19583,N_13287,N_16325);
or U19584 (N_19584,N_15042,N_14540);
nor U19585 (N_19585,N_14982,N_14043);
xnor U19586 (N_19586,N_17118,N_14190);
nor U19587 (N_19587,N_15465,N_17364);
and U19588 (N_19588,N_16538,N_14123);
nand U19589 (N_19589,N_14280,N_15345);
and U19590 (N_19590,N_15132,N_13077);
xor U19591 (N_19591,N_13459,N_16598);
xor U19592 (N_19592,N_15928,N_17785);
or U19593 (N_19593,N_16317,N_13341);
or U19594 (N_19594,N_16788,N_16288);
or U19595 (N_19595,N_18201,N_18660);
and U19596 (N_19596,N_15000,N_13576);
xnor U19597 (N_19597,N_17136,N_16355);
nand U19598 (N_19598,N_17668,N_18511);
nor U19599 (N_19599,N_13484,N_16122);
and U19600 (N_19600,N_17798,N_13540);
nand U19601 (N_19601,N_18574,N_14575);
and U19602 (N_19602,N_13337,N_17435);
nor U19603 (N_19603,N_16601,N_15446);
nand U19604 (N_19604,N_13575,N_16721);
or U19605 (N_19605,N_13009,N_16521);
nand U19606 (N_19606,N_13682,N_14652);
or U19607 (N_19607,N_12927,N_18661);
or U19608 (N_19608,N_14395,N_12853);
and U19609 (N_19609,N_17814,N_14524);
and U19610 (N_19610,N_13770,N_17936);
xnor U19611 (N_19611,N_17367,N_14592);
nor U19612 (N_19612,N_16296,N_16616);
and U19613 (N_19613,N_15323,N_18687);
nand U19614 (N_19614,N_18531,N_16750);
xnor U19615 (N_19615,N_16978,N_17083);
and U19616 (N_19616,N_16498,N_18414);
xnor U19617 (N_19617,N_17971,N_16749);
nand U19618 (N_19618,N_15999,N_16918);
xnor U19619 (N_19619,N_17278,N_12580);
xnor U19620 (N_19620,N_17354,N_16427);
xnor U19621 (N_19621,N_18138,N_17895);
or U19622 (N_19622,N_13640,N_15883);
and U19623 (N_19623,N_18638,N_13269);
and U19624 (N_19624,N_17518,N_17245);
xor U19625 (N_19625,N_13926,N_18501);
and U19626 (N_19626,N_13924,N_14323);
or U19627 (N_19627,N_16579,N_17471);
nand U19628 (N_19628,N_15418,N_14755);
nor U19629 (N_19629,N_14050,N_14487);
nor U19630 (N_19630,N_17304,N_14568);
nor U19631 (N_19631,N_13058,N_13602);
nor U19632 (N_19632,N_17899,N_16130);
nand U19633 (N_19633,N_13330,N_16913);
and U19634 (N_19634,N_13692,N_15608);
and U19635 (N_19635,N_12748,N_18012);
xor U19636 (N_19636,N_18006,N_13005);
or U19637 (N_19637,N_13843,N_13899);
or U19638 (N_19638,N_14777,N_14993);
nor U19639 (N_19639,N_17713,N_14855);
and U19640 (N_19640,N_17197,N_13542);
and U19641 (N_19641,N_15739,N_14398);
xor U19642 (N_19642,N_15890,N_17038);
nor U19643 (N_19643,N_16774,N_15060);
xnor U19644 (N_19644,N_17496,N_18156);
or U19645 (N_19645,N_17165,N_17844);
or U19646 (N_19646,N_18381,N_17719);
and U19647 (N_19647,N_14453,N_16295);
nand U19648 (N_19648,N_17500,N_12630);
and U19649 (N_19649,N_16995,N_18532);
and U19650 (N_19650,N_14181,N_15646);
nor U19651 (N_19651,N_14339,N_17084);
nor U19652 (N_19652,N_13447,N_17749);
nor U19653 (N_19653,N_18175,N_17461);
xor U19654 (N_19654,N_17298,N_13974);
nor U19655 (N_19655,N_15452,N_12953);
xor U19656 (N_19656,N_15428,N_17113);
and U19657 (N_19657,N_15366,N_15750);
nand U19658 (N_19658,N_17863,N_14374);
or U19659 (N_19659,N_16512,N_15033);
nor U19660 (N_19660,N_16156,N_17615);
and U19661 (N_19661,N_17995,N_12960);
and U19662 (N_19662,N_13830,N_18405);
or U19663 (N_19663,N_14221,N_14319);
xor U19664 (N_19664,N_17073,N_17540);
or U19665 (N_19665,N_13401,N_15657);
xnor U19666 (N_19666,N_13465,N_18426);
or U19667 (N_19667,N_14177,N_13732);
nand U19668 (N_19668,N_17622,N_17892);
and U19669 (N_19669,N_13541,N_13202);
xnor U19670 (N_19670,N_18129,N_13900);
nand U19671 (N_19671,N_18249,N_16544);
xor U19672 (N_19672,N_12889,N_14392);
nor U19673 (N_19673,N_13805,N_16352);
xor U19674 (N_19674,N_16377,N_17848);
xnor U19675 (N_19675,N_16441,N_14718);
or U19676 (N_19676,N_17409,N_15118);
nor U19677 (N_19677,N_17570,N_13344);
nand U19678 (N_19678,N_14149,N_15882);
xor U19679 (N_19679,N_12719,N_16020);
or U19680 (N_19680,N_12683,N_17323);
xor U19681 (N_19681,N_14112,N_18248);
xnor U19682 (N_19682,N_17087,N_14622);
nand U19683 (N_19683,N_15615,N_15605);
or U19684 (N_19684,N_15478,N_15329);
xor U19685 (N_19685,N_15458,N_17628);
xor U19686 (N_19686,N_13592,N_18469);
xor U19687 (N_19687,N_16102,N_13065);
nor U19688 (N_19688,N_13325,N_12660);
nand U19689 (N_19689,N_13677,N_13179);
nor U19690 (N_19690,N_13209,N_15969);
nand U19691 (N_19691,N_16751,N_14071);
nand U19692 (N_19692,N_15957,N_16526);
nor U19693 (N_19693,N_18637,N_17757);
nor U19694 (N_19694,N_13436,N_17346);
or U19695 (N_19695,N_12714,N_16516);
xor U19696 (N_19696,N_16891,N_14137);
or U19697 (N_19697,N_14228,N_15437);
and U19698 (N_19698,N_14076,N_13174);
or U19699 (N_19699,N_13917,N_15904);
or U19700 (N_19700,N_18404,N_18038);
xnor U19701 (N_19701,N_14992,N_16161);
and U19702 (N_19702,N_18071,N_14165);
and U19703 (N_19703,N_17726,N_17135);
nor U19704 (N_19704,N_16278,N_18298);
nor U19705 (N_19705,N_17044,N_16084);
xnor U19706 (N_19706,N_18741,N_14100);
nor U19707 (N_19707,N_17455,N_17508);
nor U19708 (N_19708,N_12794,N_15318);
nor U19709 (N_19709,N_16602,N_12537);
nor U19710 (N_19710,N_15740,N_14534);
nand U19711 (N_19711,N_17985,N_17994);
or U19712 (N_19712,N_14940,N_15754);
and U19713 (N_19713,N_16997,N_12702);
nand U19714 (N_19714,N_16424,N_18273);
xnor U19715 (N_19715,N_13421,N_16434);
or U19716 (N_19716,N_14922,N_12573);
nor U19717 (N_19717,N_16261,N_15692);
and U19718 (N_19718,N_13902,N_18312);
nor U19719 (N_19719,N_14710,N_13950);
and U19720 (N_19720,N_14405,N_16723);
nor U19721 (N_19721,N_16920,N_14196);
or U19722 (N_19722,N_18648,N_14942);
nand U19723 (N_19723,N_17235,N_14837);
or U19724 (N_19724,N_13995,N_15998);
nor U19725 (N_19725,N_12995,N_14646);
nor U19726 (N_19726,N_14116,N_13464);
or U19727 (N_19727,N_17295,N_14572);
xnor U19728 (N_19728,N_14372,N_16908);
nor U19729 (N_19729,N_18465,N_18019);
or U19730 (N_19730,N_15555,N_13335);
nor U19731 (N_19731,N_18479,N_15959);
and U19732 (N_19732,N_18173,N_18705);
xor U19733 (N_19733,N_17378,N_18034);
xnor U19734 (N_19734,N_14632,N_16321);
nor U19735 (N_19735,N_17635,N_13778);
nor U19736 (N_19736,N_15922,N_15433);
and U19737 (N_19737,N_12664,N_12604);
nor U19738 (N_19738,N_18028,N_17803);
or U19739 (N_19739,N_14545,N_16468);
and U19740 (N_19740,N_13151,N_18010);
nor U19741 (N_19741,N_17216,N_13016);
nand U19742 (N_19742,N_14164,N_12938);
xnor U19743 (N_19743,N_18189,N_16797);
nor U19744 (N_19744,N_15831,N_13765);
nor U19745 (N_19745,N_15055,N_17823);
xnor U19746 (N_19746,N_12970,N_15269);
nand U19747 (N_19747,N_17563,N_16817);
and U19748 (N_19748,N_16540,N_16258);
xnor U19749 (N_19749,N_16657,N_17121);
and U19750 (N_19750,N_17906,N_18458);
xor U19751 (N_19751,N_15776,N_13577);
or U19752 (N_19752,N_17666,N_14737);
and U19753 (N_19753,N_16932,N_17393);
xnor U19754 (N_19754,N_16075,N_16905);
nor U19755 (N_19755,N_16990,N_15341);
nand U19756 (N_19756,N_15262,N_14910);
nor U19757 (N_19757,N_16146,N_13794);
nor U19758 (N_19758,N_18490,N_16806);
or U19759 (N_19759,N_17456,N_15460);
or U19760 (N_19760,N_18586,N_17381);
nor U19761 (N_19761,N_16807,N_13153);
nor U19762 (N_19762,N_12730,N_16840);
and U19763 (N_19763,N_13030,N_12944);
nand U19764 (N_19764,N_12534,N_15072);
or U19765 (N_19765,N_13820,N_16785);
or U19766 (N_19766,N_14945,N_15822);
and U19767 (N_19767,N_16963,N_17253);
or U19768 (N_19768,N_16804,N_14375);
xor U19769 (N_19769,N_18565,N_18000);
and U19770 (N_19770,N_15909,N_18627);
xor U19771 (N_19771,N_17388,N_17676);
nand U19772 (N_19772,N_14491,N_14450);
nand U19773 (N_19773,N_17996,N_13384);
or U19774 (N_19774,N_17969,N_14699);
and U19775 (N_19775,N_15321,N_13568);
nor U19776 (N_19776,N_12598,N_14170);
nand U19777 (N_19777,N_17710,N_18597);
and U19778 (N_19778,N_14408,N_14807);
and U19779 (N_19779,N_18647,N_17706);
nor U19780 (N_19780,N_17527,N_12610);
nor U19781 (N_19781,N_17195,N_15085);
xor U19782 (N_19782,N_13690,N_13047);
nor U19783 (N_19783,N_12763,N_15558);
or U19784 (N_19784,N_17306,N_14790);
and U19785 (N_19785,N_12832,N_12725);
and U19786 (N_19786,N_14120,N_17151);
xor U19787 (N_19787,N_16708,N_12519);
nand U19788 (N_19788,N_18358,N_16921);
or U19789 (N_19789,N_16938,N_18686);
and U19790 (N_19790,N_15746,N_13366);
nor U19791 (N_19791,N_16930,N_16094);
nor U19792 (N_19792,N_14871,N_14919);
and U19793 (N_19793,N_14462,N_16873);
nor U19794 (N_19794,N_18575,N_17695);
or U19795 (N_19795,N_17840,N_15485);
and U19796 (N_19796,N_15170,N_12612);
nor U19797 (N_19797,N_17318,N_15749);
or U19798 (N_19798,N_16187,N_15897);
or U19799 (N_19799,N_16519,N_14066);
nor U19800 (N_19800,N_14536,N_14442);
nor U19801 (N_19801,N_15675,N_17105);
xor U19802 (N_19802,N_12754,N_17303);
nor U19803 (N_19803,N_12766,N_15539);
nor U19804 (N_19804,N_18442,N_12726);
nor U19805 (N_19805,N_13054,N_13383);
nand U19806 (N_19806,N_16898,N_13103);
nor U19807 (N_19807,N_15632,N_14062);
nand U19808 (N_19808,N_14458,N_13458);
nand U19809 (N_19809,N_13659,N_17225);
nand U19810 (N_19810,N_17989,N_16059);
xor U19811 (N_19811,N_12817,N_13375);
nand U19812 (N_19812,N_13422,N_16314);
nand U19813 (N_19813,N_16368,N_17959);
xnor U19814 (N_19814,N_17774,N_14905);
or U19815 (N_19815,N_14136,N_14582);
xnor U19816 (N_19816,N_15025,N_17096);
xnor U19817 (N_19817,N_16208,N_16917);
nand U19818 (N_19818,N_15908,N_14198);
or U19819 (N_19819,N_16625,N_18202);
and U19820 (N_19820,N_14916,N_15004);
and U19821 (N_19821,N_16494,N_14591);
xor U19822 (N_19822,N_18649,N_12850);
nand U19823 (N_19823,N_17976,N_14918);
nor U19824 (N_19824,N_15188,N_16823);
or U19825 (N_19825,N_14096,N_17832);
and U19826 (N_19826,N_15816,N_13562);
nand U19827 (N_19827,N_12904,N_18392);
or U19828 (N_19828,N_16178,N_15941);
nor U19829 (N_19829,N_16741,N_18332);
and U19830 (N_19830,N_15527,N_14468);
and U19831 (N_19831,N_17276,N_12706);
and U19832 (N_19832,N_17184,N_15337);
nand U19833 (N_19833,N_14085,N_12991);
or U19834 (N_19834,N_17716,N_14292);
and U19835 (N_19835,N_12671,N_18345);
and U19836 (N_19836,N_13266,N_18205);
nand U19837 (N_19837,N_16977,N_13730);
xor U19838 (N_19838,N_14013,N_12596);
xnor U19839 (N_19839,N_15284,N_12951);
xor U19840 (N_19840,N_17529,N_13858);
or U19841 (N_19841,N_18242,N_17531);
nor U19842 (N_19842,N_13177,N_13898);
xnor U19843 (N_19843,N_13766,N_13001);
nand U19844 (N_19844,N_13556,N_13589);
nor U19845 (N_19845,N_13317,N_16192);
nor U19846 (N_19846,N_18119,N_14420);
or U19847 (N_19847,N_17115,N_13499);
and U19848 (N_19848,N_16149,N_17551);
and U19849 (N_19849,N_17261,N_17762);
xnor U19850 (N_19850,N_17612,N_12760);
and U19851 (N_19851,N_12525,N_16221);
nor U19852 (N_19852,N_17452,N_14449);
and U19853 (N_19853,N_15961,N_13578);
or U19854 (N_19854,N_17657,N_15929);
nand U19855 (N_19855,N_18065,N_12647);
xor U19856 (N_19856,N_14192,N_16155);
nand U19857 (N_19857,N_17061,N_18524);
and U19858 (N_19858,N_18598,N_17573);
nor U19859 (N_19859,N_16386,N_13374);
or U19860 (N_19860,N_18599,N_18152);
and U19861 (N_19861,N_12772,N_16307);
nand U19862 (N_19862,N_12840,N_17793);
xor U19863 (N_19863,N_14335,N_17561);
nor U19864 (N_19864,N_14860,N_14743);
nor U19865 (N_19865,N_14819,N_14361);
nor U19866 (N_19866,N_17391,N_13978);
xor U19867 (N_19867,N_17001,N_18212);
and U19868 (N_19868,N_18446,N_15971);
nand U19869 (N_19869,N_16687,N_13258);
nor U19870 (N_19870,N_17503,N_14981);
nor U19871 (N_19871,N_14629,N_13516);
nor U19872 (N_19872,N_15111,N_14525);
or U19873 (N_19873,N_16351,N_15017);
or U19874 (N_19874,N_17826,N_17414);
nor U19875 (N_19875,N_17007,N_14887);
nor U19876 (N_19876,N_14995,N_14815);
or U19877 (N_19877,N_18579,N_12847);
nand U19878 (N_19878,N_17746,N_17351);
or U19879 (N_19879,N_14261,N_17767);
xor U19880 (N_19880,N_16229,N_12797);
nor U19881 (N_19881,N_16588,N_13756);
nor U19882 (N_19882,N_18559,N_15048);
or U19883 (N_19883,N_13098,N_12903);
xnor U19884 (N_19884,N_17809,N_12836);
nor U19885 (N_19885,N_13873,N_14058);
nor U19886 (N_19886,N_17795,N_12721);
nor U19887 (N_19887,N_18514,N_13635);
or U19888 (N_19888,N_17596,N_16240);
or U19889 (N_19889,N_15840,N_14966);
nand U19890 (N_19890,N_18390,N_18339);
nand U19891 (N_19891,N_13149,N_15398);
nand U19892 (N_19892,N_16801,N_15599);
or U19893 (N_19893,N_18669,N_16273);
or U19894 (N_19894,N_14227,N_17932);
nor U19895 (N_19895,N_16742,N_13760);
xor U19896 (N_19896,N_18369,N_16529);
nor U19897 (N_19897,N_16272,N_13506);
nand U19898 (N_19898,N_16981,N_16373);
nand U19899 (N_19899,N_16128,N_16752);
and U19900 (N_19900,N_18419,N_17498);
or U19901 (N_19901,N_18577,N_12662);
nor U19902 (N_19902,N_14601,N_16504);
nor U19903 (N_19903,N_17467,N_14606);
nor U19904 (N_19904,N_16328,N_13755);
xor U19905 (N_19905,N_15808,N_14846);
nand U19906 (N_19906,N_16926,N_18220);
nor U19907 (N_19907,N_17368,N_12574);
xnor U19908 (N_19908,N_15275,N_13712);
xnor U19909 (N_19909,N_18656,N_13894);
nor U19910 (N_19910,N_14061,N_17423);
and U19911 (N_19911,N_17036,N_18515);
nor U19912 (N_19912,N_18286,N_14175);
and U19913 (N_19913,N_13890,N_12691);
xnor U19914 (N_19914,N_15381,N_15757);
or U19915 (N_19915,N_15886,N_12762);
and U19916 (N_19916,N_18042,N_16779);
or U19917 (N_19917,N_17543,N_13002);
and U19918 (N_19918,N_15034,N_15811);
or U19919 (N_19919,N_17526,N_15624);
nor U19920 (N_19920,N_14938,N_12773);
or U19921 (N_19921,N_12584,N_16243);
xor U19922 (N_19922,N_14694,N_14758);
nand U19923 (N_19923,N_16139,N_18452);
xnor U19924 (N_19924,N_15644,N_15798);
or U19925 (N_19925,N_15879,N_13096);
xnor U19926 (N_19926,N_14516,N_17374);
and U19927 (N_19927,N_14040,N_17271);
nor U19928 (N_19928,N_16830,N_13444);
or U19929 (N_19929,N_17178,N_16761);
xnor U19930 (N_19930,N_14554,N_15294);
nor U19931 (N_19931,N_18713,N_14172);
nor U19932 (N_19932,N_15540,N_15300);
and U19933 (N_19933,N_14254,N_18264);
nand U19934 (N_19934,N_14288,N_13612);
or U19935 (N_19935,N_14482,N_16611);
and U19936 (N_19936,N_18372,N_17214);
xor U19937 (N_19937,N_15146,N_13090);
xnor U19938 (N_19938,N_12599,N_14219);
nand U19939 (N_19939,N_17624,N_13633);
and U19940 (N_19940,N_13381,N_14020);
or U19941 (N_19941,N_17065,N_18341);
nand U19942 (N_19942,N_14167,N_15219);
nand U19943 (N_19943,N_16675,N_16446);
nor U19944 (N_19944,N_12814,N_18304);
or U19945 (N_19945,N_18743,N_18063);
or U19946 (N_19946,N_17267,N_13885);
and U19947 (N_19947,N_16705,N_13239);
or U19948 (N_19948,N_16141,N_13810);
nand U19949 (N_19949,N_13731,N_18001);
and U19950 (N_19950,N_12870,N_18717);
or U19951 (N_19951,N_13340,N_13394);
nor U19952 (N_19952,N_12512,N_15685);
or U19953 (N_19953,N_16478,N_16839);
nand U19954 (N_19954,N_14484,N_16828);
nand U19955 (N_19955,N_13747,N_15051);
nor U19956 (N_19956,N_18456,N_12653);
nand U19957 (N_19957,N_18296,N_13253);
nor U19958 (N_19958,N_15942,N_17955);
nor U19959 (N_19959,N_13500,N_17835);
or U19960 (N_19960,N_12511,N_14859);
nor U19961 (N_19961,N_13230,N_16791);
nor U19962 (N_19962,N_14619,N_15946);
nor U19963 (N_19963,N_14424,N_15859);
xor U19964 (N_19964,N_15733,N_17787);
nand U19965 (N_19965,N_13580,N_18517);
or U19966 (N_19966,N_17385,N_16935);
nand U19967 (N_19967,N_15801,N_14820);
nor U19968 (N_19968,N_16029,N_18311);
nand U19969 (N_19969,N_18546,N_17120);
nand U19970 (N_19970,N_16720,N_16466);
and U19971 (N_19971,N_13941,N_18391);
xor U19972 (N_19972,N_12808,N_14603);
nand U19973 (N_19973,N_13069,N_14354);
xnor U19974 (N_19974,N_16496,N_13237);
xor U19975 (N_19975,N_16419,N_13567);
and U19976 (N_19976,N_18396,N_18244);
nand U19977 (N_19977,N_16805,N_14098);
nand U19978 (N_19978,N_14677,N_14282);
nand U19979 (N_19979,N_14792,N_15308);
and U19980 (N_19980,N_15380,N_14121);
nand U19981 (N_19981,N_16557,N_16523);
nor U19982 (N_19982,N_16881,N_14174);
nand U19983 (N_19983,N_12804,N_13834);
and U19984 (N_19984,N_18274,N_16669);
xnor U19985 (N_19985,N_15150,N_18103);
and U19986 (N_19986,N_16108,N_13301);
nor U19987 (N_19987,N_14750,N_15036);
or U19988 (N_19988,N_12942,N_17609);
nor U19989 (N_19989,N_14215,N_18316);
nor U19990 (N_19990,N_14980,N_17546);
nand U19991 (N_19991,N_13322,N_12800);
and U19992 (N_19992,N_16431,N_16121);
and U19993 (N_19993,N_16545,N_18706);
and U19994 (N_19994,N_17931,N_15243);
and U19995 (N_19995,N_13954,N_17528);
and U19996 (N_19996,N_14675,N_18044);
or U19997 (N_19997,N_13700,N_17132);
xnor U19998 (N_19998,N_14332,N_17565);
xor U19999 (N_19999,N_15913,N_16392);
and U20000 (N_20000,N_13674,N_15664);
and U20001 (N_20001,N_13482,N_16153);
or U20002 (N_20002,N_12784,N_15178);
or U20003 (N_20003,N_14057,N_13777);
and U20004 (N_20004,N_18011,N_14433);
nand U20005 (N_20005,N_16608,N_18321);
nor U20006 (N_20006,N_15763,N_15289);
nor U20007 (N_20007,N_16509,N_16477);
nor U20008 (N_20008,N_17477,N_18172);
or U20009 (N_20009,N_17642,N_17243);
nor U20010 (N_20010,N_16789,N_17681);
xnor U20011 (N_20011,N_14977,N_13497);
and U20012 (N_20012,N_17697,N_18337);
and U20013 (N_20013,N_18569,N_15319);
and U20014 (N_20014,N_18688,N_18408);
xnor U20015 (N_20015,N_12648,N_18070);
or U20016 (N_20016,N_15196,N_14139);
or U20017 (N_20017,N_17705,N_15614);
or U20018 (N_20018,N_16524,N_18313);
nand U20019 (N_20019,N_14833,N_18174);
xor U20020 (N_20020,N_15161,N_13172);
nor U20021 (N_20021,N_18090,N_15849);
xnor U20022 (N_20022,N_12569,N_13991);
nand U20023 (N_20023,N_14969,N_16685);
xnor U20024 (N_20024,N_12570,N_15537);
nand U20025 (N_20025,N_16968,N_15805);
and U20026 (N_20026,N_13348,N_17302);
nand U20027 (N_20027,N_18346,N_18101);
xor U20028 (N_20028,N_13708,N_13823);
or U20029 (N_20029,N_15888,N_14012);
xor U20030 (N_20030,N_16275,N_16032);
and U20031 (N_20031,N_18013,N_16894);
and U20032 (N_20032,N_13010,N_15057);
xnor U20033 (N_20033,N_18262,N_18093);
nor U20034 (N_20034,N_15207,N_18178);
xor U20035 (N_20035,N_13268,N_17299);
xor U20036 (N_20036,N_16070,N_14079);
and U20037 (N_20037,N_15713,N_17040);
nand U20038 (N_20038,N_13449,N_16231);
and U20039 (N_20039,N_18634,N_17937);
nand U20040 (N_20040,N_16565,N_17853);
and U20041 (N_20041,N_17614,N_17292);
nand U20042 (N_20042,N_15885,N_12894);
xnor U20043 (N_20043,N_13013,N_15986);
or U20044 (N_20044,N_18644,N_13439);
or U20045 (N_20045,N_15238,N_13826);
xnor U20046 (N_20046,N_15812,N_15068);
nor U20047 (N_20047,N_12700,N_15518);
nor U20048 (N_20048,N_14566,N_14419);
and U20049 (N_20049,N_16757,N_18187);
xor U20050 (N_20050,N_16034,N_13738);
or U20051 (N_20051,N_17396,N_15391);
or U20052 (N_20052,N_17099,N_13845);
xor U20053 (N_20053,N_13318,N_16619);
nand U20054 (N_20054,N_14811,N_13695);
or U20055 (N_20055,N_14256,N_18530);
nor U20056 (N_20056,N_14695,N_14410);
or U20057 (N_20057,N_16802,N_17775);
nand U20058 (N_20058,N_18643,N_12914);
xor U20059 (N_20059,N_17672,N_17797);
and U20060 (N_20060,N_15980,N_18171);
and U20061 (N_20061,N_17592,N_18348);
xor U20062 (N_20062,N_15977,N_16011);
nor U20063 (N_20063,N_14642,N_12670);
or U20064 (N_20064,N_18571,N_12829);
xor U20065 (N_20065,N_15975,N_18137);
nor U20066 (N_20066,N_17569,N_14384);
xnor U20067 (N_20067,N_15526,N_16711);
and U20068 (N_20068,N_13259,N_12750);
or U20069 (N_20069,N_13231,N_14377);
nand U20070 (N_20070,N_15827,N_18685);
and U20071 (N_20071,N_18122,N_18440);
nor U20072 (N_20072,N_13356,N_13849);
or U20073 (N_20073,N_18360,N_17317);
and U20074 (N_20074,N_13437,N_15122);
and U20075 (N_20075,N_14952,N_14593);
nand U20076 (N_20076,N_18361,N_13379);
or U20077 (N_20077,N_14297,N_18199);
and U20078 (N_20078,N_15279,N_12538);
nand U20079 (N_20079,N_15596,N_15092);
xnor U20080 (N_20080,N_14234,N_16667);
and U20081 (N_20081,N_15352,N_16702);
xor U20082 (N_20082,N_18014,N_14596);
nor U20083 (N_20083,N_17545,N_13338);
nor U20084 (N_20084,N_15873,N_14721);
or U20085 (N_20085,N_15967,N_17788);
nor U20086 (N_20086,N_15704,N_12935);
and U20087 (N_20087,N_16630,N_13857);
or U20088 (N_20088,N_12834,N_17193);
and U20089 (N_20089,N_12868,N_12962);
nor U20090 (N_20090,N_16340,N_15752);
xor U20091 (N_20091,N_12862,N_14006);
nand U20092 (N_20092,N_17831,N_15542);
and U20093 (N_20093,N_15244,N_15211);
nand U20094 (N_20094,N_15180,N_18421);
xnor U20095 (N_20095,N_12513,N_16843);
or U20096 (N_20096,N_15693,N_14844);
nand U20097 (N_20097,N_14576,N_17914);
nor U20098 (N_20098,N_16247,N_12918);
nand U20099 (N_20099,N_14978,N_15786);
nor U20100 (N_20100,N_13143,N_16962);
nand U20101 (N_20101,N_16961,N_12752);
nand U20102 (N_20102,N_14735,N_15445);
or U20103 (N_20103,N_13790,N_18471);
or U20104 (N_20104,N_15489,N_12602);
nand U20105 (N_20105,N_16915,N_16682);
and U20106 (N_20106,N_16482,N_16475);
nor U20107 (N_20107,N_13155,N_14027);
xnor U20108 (N_20108,N_15620,N_14459);
and U20109 (N_20109,N_15001,N_15186);
xnor U20110 (N_20110,N_18695,N_16716);
or U20111 (N_20111,N_12833,N_15698);
xor U20112 (N_20112,N_15679,N_14894);
nor U20113 (N_20113,N_13630,N_15819);
nor U20114 (N_20114,N_18707,N_14872);
xor U20115 (N_20115,N_13195,N_12717);
nand U20116 (N_20116,N_16471,N_15440);
nand U20117 (N_20117,N_14448,N_13672);
nand U20118 (N_20118,N_15841,N_18351);
nand U20119 (N_20119,N_15200,N_12716);
nor U20120 (N_20120,N_15450,N_17884);
nor U20121 (N_20121,N_15830,N_16659);
or U20122 (N_20122,N_17783,N_18250);
nand U20123 (N_20123,N_15468,N_12842);
nor U20124 (N_20124,N_17755,N_14604);
nor U20125 (N_20125,N_16202,N_14162);
nor U20126 (N_20126,N_17519,N_17379);
nand U20127 (N_20127,N_14145,N_16193);
nand U20128 (N_20128,N_15715,N_14383);
and U20129 (N_20129,N_15802,N_18016);
and U20130 (N_20130,N_17418,N_16706);
nor U20131 (N_20131,N_12968,N_17013);
nor U20132 (N_20132,N_18447,N_16088);
nand U20133 (N_20133,N_15966,N_12973);
or U20134 (N_20134,N_15839,N_16649);
xnor U20135 (N_20135,N_13667,N_13976);
or U20136 (N_20136,N_18407,N_14529);
xnor U20137 (N_20137,N_13745,N_17900);
and U20138 (N_20138,N_16484,N_13701);
or U20139 (N_20139,N_18608,N_14203);
nor U20140 (N_20140,N_13534,N_16045);
and U20141 (N_20141,N_13702,N_17443);
nor U20142 (N_20142,N_13473,N_14217);
nand U20143 (N_20143,N_16203,N_14379);
xnor U20144 (N_20144,N_13590,N_13349);
or U20145 (N_20145,N_17876,N_18558);
xnor U20146 (N_20146,N_17022,N_15931);
nor U20147 (N_20147,N_14847,N_15955);
nor U20148 (N_20148,N_16337,N_16768);
xnor U20149 (N_20149,N_12971,N_12966);
xor U20150 (N_20150,N_12860,N_17966);
nor U20151 (N_20151,N_13508,N_15654);
and U20152 (N_20152,N_12658,N_12851);
nor U20153 (N_20153,N_14637,N_15600);
nor U20154 (N_20154,N_14494,N_18204);
or U20155 (N_20155,N_13716,N_15996);
xor U20156 (N_20156,N_14210,N_17638);
nand U20157 (N_20157,N_17613,N_15729);
nor U20158 (N_20158,N_14084,N_17064);
and U20159 (N_20159,N_16488,N_18673);
or U20160 (N_20160,N_13038,N_18494);
nor U20161 (N_20161,N_17160,N_18107);
or U20162 (N_20162,N_16627,N_15894);
and U20163 (N_20163,N_17489,N_16031);
nor U20164 (N_20164,N_18444,N_14520);
nand U20165 (N_20165,N_14595,N_15560);
and U20166 (N_20166,N_15718,N_14312);
nand U20167 (N_20167,N_14294,N_14421);
and U20168 (N_20168,N_17893,N_17845);
nand U20169 (N_20169,N_12798,N_17314);
nor U20170 (N_20170,N_12813,N_14920);
nor U20171 (N_20171,N_13277,N_13425);
and U20172 (N_20172,N_16489,N_15417);
nor U20173 (N_20173,N_17739,N_14886);
nor U20174 (N_20174,N_17279,N_14802);
or U20175 (N_20175,N_16265,N_16062);
nor U20176 (N_20176,N_13861,N_18589);
nor U20177 (N_20177,N_15239,N_18508);
nor U20178 (N_20178,N_18164,N_18701);
or U20179 (N_20179,N_18431,N_17458);
nand U20180 (N_20180,N_14951,N_13410);
xnor U20181 (N_20181,N_15784,N_17006);
nor U20182 (N_20182,N_14285,N_15905);
nand U20183 (N_20183,N_16050,N_14521);
and U20184 (N_20184,N_16541,N_13018);
or U20185 (N_20185,N_15762,N_17234);
nand U20186 (N_20186,N_16890,N_18496);
and U20187 (N_20187,N_14785,N_14417);
nor U20188 (N_20188,N_12678,N_15949);
xor U20189 (N_20189,N_17555,N_16772);
xnor U20190 (N_20190,N_16700,N_12939);
or U20191 (N_20191,N_17683,N_18365);
and U20192 (N_20192,N_14683,N_17619);
and U20193 (N_20193,N_12827,N_15204);
and U20194 (N_20194,N_16880,N_15074);
or U20195 (N_20195,N_17712,N_15727);
and U20196 (N_20196,N_13656,N_14853);
nor U20197 (N_20197,N_15448,N_15053);
or U20198 (N_20198,N_12897,N_14680);
and U20199 (N_20199,N_13240,N_13159);
nand U20200 (N_20200,N_14638,N_17629);
or U20201 (N_20201,N_15835,N_13254);
nand U20202 (N_20202,N_15521,N_17049);
xnor U20203 (N_20203,N_17322,N_18240);
and U20204 (N_20204,N_16144,N_17394);
nand U20205 (N_20205,N_14200,N_15611);
nand U20206 (N_20206,N_15228,N_15332);
and U20207 (N_20207,N_15240,N_15303);
and U20208 (N_20208,N_16366,N_18003);
nor U20209 (N_20209,N_13123,N_13691);
and U20210 (N_20210,N_13281,N_17980);
and U20211 (N_20211,N_17282,N_13476);
nor U20212 (N_20212,N_15265,N_18203);
nor U20213 (N_20213,N_17894,N_16293);
nand U20214 (N_20214,N_15979,N_16350);
and U20215 (N_20215,N_14360,N_12618);
or U20216 (N_20216,N_13035,N_16878);
nor U20217 (N_20217,N_15378,N_12774);
nand U20218 (N_20218,N_13709,N_17281);
and U20219 (N_20219,N_12878,N_15189);
and U20220 (N_20220,N_16047,N_13081);
nor U20221 (N_20221,N_17866,N_15235);
nor U20222 (N_20222,N_13089,N_14225);
and U20223 (N_20223,N_14697,N_14868);
and U20224 (N_20224,N_13838,N_17779);
or U20225 (N_20225,N_12607,N_17041);
nor U20226 (N_20226,N_13653,N_15320);
and U20227 (N_20227,N_17849,N_15984);
xnor U20228 (N_20228,N_14466,N_15121);
nor U20229 (N_20229,N_12824,N_15731);
nor U20230 (N_20230,N_17737,N_18617);
and U20231 (N_20231,N_14501,N_18595);
and U20232 (N_20232,N_13771,N_12844);
and U20233 (N_20233,N_17806,N_13998);
or U20234 (N_20234,N_13106,N_16060);
and U20235 (N_20235,N_18402,N_13248);
and U20236 (N_20236,N_15934,N_14663);
xnor U20237 (N_20237,N_15807,N_15732);
nand U20238 (N_20238,N_16643,N_12810);
nand U20239 (N_20239,N_15221,N_16004);
and U20240 (N_20240,N_14002,N_12567);
nor U20241 (N_20241,N_16868,N_18529);
nor U20242 (N_20242,N_16013,N_16786);
and U20243 (N_20243,N_16406,N_15990);
and U20244 (N_20244,N_17011,N_17089);
nor U20245 (N_20245,N_14927,N_17660);
xnor U20246 (N_20246,N_17371,N_14140);
nor U20247 (N_20247,N_13668,N_14760);
and U20248 (N_20248,N_15570,N_12644);
nand U20249 (N_20249,N_14671,N_15992);
or U20250 (N_20250,N_18302,N_15525);
nand U20251 (N_20251,N_17101,N_18376);
or U20252 (N_20252,N_13470,N_16876);
nor U20253 (N_20253,N_14406,N_14456);
or U20254 (N_20254,N_16781,N_16465);
and U20255 (N_20255,N_17769,N_12667);
nor U20256 (N_20256,N_13399,N_15923);
nor U20257 (N_20257,N_16552,N_18484);
and U20258 (N_20258,N_15924,N_14931);
xnor U20259 (N_20259,N_14803,N_15493);
and U20260 (N_20260,N_16445,N_17052);
xor U20261 (N_20261,N_13080,N_14711);
nor U20262 (N_20262,N_15368,N_17747);
nor U20263 (N_20263,N_12831,N_15987);
nand U20264 (N_20264,N_13988,N_12629);
nor U20265 (N_20265,N_18277,N_17232);
and U20266 (N_20266,N_17215,N_13822);
and U20267 (N_20267,N_14283,N_15753);
or U20268 (N_20268,N_14347,N_12505);
and U20269 (N_20269,N_13285,N_15813);
or U20270 (N_20270,N_13560,N_17468);
nor U20271 (N_20271,N_14014,N_18470);
or U20272 (N_20272,N_15723,N_17241);
or U20273 (N_20273,N_16442,N_16435);
or U20274 (N_20274,N_17689,N_12830);
nand U20275 (N_20275,N_13355,N_15106);
or U20276 (N_20276,N_12549,N_16169);
nand U20277 (N_20277,N_15586,N_14431);
and U20278 (N_20278,N_17544,N_17677);
or U20279 (N_20279,N_13032,N_17890);
xor U20280 (N_20280,N_14628,N_14302);
nand U20281 (N_20281,N_14924,N_16888);
xnor U20282 (N_20282,N_16943,N_15935);
xnor U20283 (N_20283,N_14728,N_18200);
xnor U20284 (N_20284,N_13875,N_15789);
xnor U20285 (N_20285,N_18475,N_13491);
xnor U20286 (N_20286,N_18177,N_16916);
nor U20287 (N_20287,N_15960,N_18319);
or U20288 (N_20288,N_18102,N_12516);
xnor U20289 (N_20289,N_18521,N_14010);
and U20290 (N_20290,N_17905,N_13839);
and U20291 (N_20291,N_13271,N_14928);
nor U20292 (N_20292,N_13389,N_17694);
nand U20293 (N_20293,N_18104,N_15166);
or U20294 (N_20294,N_13647,N_14371);
and U20295 (N_20295,N_17425,N_15580);
and U20296 (N_20296,N_17568,N_16622);
or U20297 (N_20297,N_18499,N_15449);
nor U20298 (N_20298,N_16087,N_15503);
or U20299 (N_20299,N_18176,N_16834);
xor U20300 (N_20300,N_18745,N_17485);
nor U20301 (N_20301,N_13413,N_17077);
nand U20302 (N_20302,N_17512,N_17211);
nand U20303 (N_20303,N_17002,N_13319);
nand U20304 (N_20304,N_16832,N_15639);
and U20305 (N_20305,N_17925,N_15722);
xor U20306 (N_20306,N_12689,N_18066);
nand U20307 (N_20307,N_16100,N_13720);
or U20308 (N_20308,N_14541,N_17426);
and U20309 (N_20309,N_14903,N_14839);
or U20310 (N_20310,N_12812,N_16838);
nand U20311 (N_20311,N_13116,N_13646);
or U20312 (N_20312,N_16007,N_18474);
nor U20313 (N_20313,N_15182,N_18520);
xor U20314 (N_20314,N_12617,N_15324);
nand U20315 (N_20315,N_16848,N_16704);
nand U20316 (N_20316,N_13008,N_14643);
xnor U20317 (N_20317,N_16816,N_16341);
nor U20318 (N_20318,N_16924,N_17260);
nand U20319 (N_20319,N_17104,N_18237);
and U20320 (N_20320,N_13626,N_17313);
nor U20321 (N_20321,N_13965,N_18331);
or U20322 (N_20322,N_16680,N_17702);
or U20323 (N_20323,N_18572,N_13175);
xor U20324 (N_20324,N_16416,N_17387);
nand U20325 (N_20325,N_16975,N_14630);
nand U20326 (N_20326,N_15003,N_16664);
nor U20327 (N_20327,N_13427,N_17449);
and U20328 (N_20328,N_17109,N_14496);
xor U20329 (N_20329,N_12641,N_17218);
or U20330 (N_20330,N_13214,N_18265);
or U20331 (N_20331,N_17230,N_18356);
or U20332 (N_20332,N_13652,N_18247);
nand U20333 (N_20333,N_13938,N_15479);
nor U20334 (N_20334,N_14325,N_17069);
nor U20335 (N_20335,N_14863,N_17085);
xnor U20336 (N_20336,N_16592,N_18018);
nand U20337 (N_20337,N_16495,N_13512);
and U20338 (N_20338,N_16145,N_16744);
or U20339 (N_20339,N_14901,N_15910);
and U20340 (N_20340,N_15021,N_12695);
or U20341 (N_20341,N_14890,N_15307);
or U20342 (N_20342,N_17124,N_17878);
nand U20343 (N_20343,N_17975,N_14446);
nor U20344 (N_20344,N_12967,N_17463);
or U20345 (N_20345,N_14898,N_13161);
or U20346 (N_20346,N_12710,N_18133);
and U20347 (N_20347,N_18293,N_13922);
and U20348 (N_20348,N_12751,N_13272);
and U20349 (N_20349,N_16073,N_18068);
xor U20350 (N_20350,N_15772,N_16585);
nand U20351 (N_20351,N_15829,N_12759);
and U20352 (N_20352,N_16863,N_15832);
nand U20353 (N_20353,N_14509,N_18180);
or U20354 (N_20354,N_16284,N_17407);
nor U20355 (N_20355,N_13581,N_13714);
xnor U20356 (N_20356,N_14232,N_16738);
nor U20357 (N_20357,N_15078,N_18612);
or U20358 (N_20358,N_13598,N_15002);
xor U20359 (N_20359,N_18740,N_13675);
xor U20360 (N_20360,N_14651,N_12564);
nor U20361 (N_20361,N_14598,N_18007);
and U20362 (N_20362,N_16853,N_12673);
and U20363 (N_20363,N_18151,N_14965);
nor U20364 (N_20364,N_15673,N_18676);
or U20365 (N_20365,N_15041,N_14659);
xor U20366 (N_20366,N_16443,N_17743);
xor U20367 (N_20367,N_16091,N_13913);
or U20368 (N_20368,N_16472,N_14030);
and U20369 (N_20369,N_13190,N_17617);
nand U20370 (N_20370,N_13934,N_15551);
nor U20371 (N_20371,N_14300,N_17067);
or U20372 (N_20372,N_16399,N_12884);
xnor U20373 (N_20373,N_13392,N_13734);
xnor U20374 (N_20374,N_15217,N_15520);
nor U20375 (N_20375,N_13971,N_14435);
nor U20376 (N_20376,N_15510,N_16632);
and U20377 (N_20377,N_17114,N_13713);
or U20378 (N_20378,N_14538,N_16955);
or U20379 (N_20379,N_15348,N_15770);
nor U20380 (N_20380,N_16281,N_16227);
and U20381 (N_20381,N_14585,N_13188);
or U20382 (N_20382,N_16799,N_16266);
nand U20383 (N_20383,N_14328,N_15419);
nor U20384 (N_20384,N_15901,N_17652);
nor U20385 (N_20385,N_12858,N_17025);
nor U20386 (N_20386,N_15191,N_17897);
xor U20387 (N_20387,N_16327,N_12659);
nand U20388 (N_20388,N_13783,N_13863);
nand U20389 (N_20389,N_17515,N_13520);
nand U20390 (N_20390,N_15311,N_14666);
nand U20391 (N_20391,N_13023,N_17259);
and U20392 (N_20392,N_13661,N_14402);
xnor U20393 (N_20393,N_14314,N_12931);
xnor U20394 (N_20394,N_16077,N_13743);
xnor U20395 (N_20395,N_17924,N_12869);
nor U20396 (N_20396,N_14152,N_15044);
nand U20397 (N_20397,N_16234,N_13649);
or U20398 (N_20398,N_15792,N_18507);
xor U20399 (N_20399,N_13847,N_15203);
or U20400 (N_20400,N_12816,N_13553);
or U20401 (N_20401,N_14544,N_17263);
and U20402 (N_20402,N_16448,N_16717);
xnor U20403 (N_20403,N_17928,N_18241);
nand U20404 (N_20404,N_13122,N_18291);
or U20405 (N_20405,N_16081,N_15242);
and U20406 (N_20406,N_18227,N_18017);
and U20407 (N_20407,N_18554,N_15208);
xor U20408 (N_20408,N_17495,N_17451);
and U20409 (N_20409,N_14696,N_14953);
xor U20410 (N_20410,N_17509,N_18699);
and U20411 (N_20411,N_14759,N_17865);
nand U20412 (N_20412,N_12514,N_17068);
xor U20413 (N_20413,N_16163,N_15721);
or U20414 (N_20414,N_17478,N_12792);
xnor U20415 (N_20415,N_12731,N_16487);
and U20416 (N_20416,N_17766,N_17106);
nor U20417 (N_20417,N_14305,N_15344);
nand U20418 (N_20418,N_15306,N_15488);
nand U20419 (N_20419,N_16686,N_13999);
xnor U20420 (N_20420,N_15647,N_16490);
and U20421 (N_20421,N_14129,N_14672);
and U20422 (N_20422,N_17758,N_18020);
xor U20423 (N_20423,N_16737,N_17965);
nand U20424 (N_20424,N_15140,N_15804);
nand U20425 (N_20425,N_15330,N_12901);
nand U20426 (N_20426,N_14732,N_14650);
nand U20427 (N_20427,N_14393,N_15773);
xnor U20428 (N_20428,N_14080,N_16513);
and U20429 (N_20429,N_17082,N_17157);
nand U20430 (N_20430,N_17164,N_12600);
nand U20431 (N_20431,N_15875,N_14742);
nor U20432 (N_20432,N_16893,N_16553);
and U20433 (N_20433,N_16528,N_16994);
xnor U20434 (N_20434,N_17344,N_16755);
xnor U20435 (N_20435,N_13216,N_14571);
and U20436 (N_20436,N_17247,N_13925);
or U20437 (N_20437,N_14895,N_18040);
and U20438 (N_20438,N_17887,N_18095);
xnor U20439 (N_20439,N_12553,N_18276);
nand U20440 (N_20440,N_15735,N_15245);
nor U20441 (N_20441,N_15951,N_16909);
xor U20442 (N_20442,N_18231,N_13314);
xor U20443 (N_20443,N_12546,N_16318);
xnor U20444 (N_20444,N_15514,N_13852);
xor U20445 (N_20445,N_15274,N_13487);
nor U20446 (N_20446,N_13510,N_18478);
xnor U20447 (N_20447,N_14038,N_14222);
nor U20448 (N_20448,N_15997,N_14752);
nand U20449 (N_20449,N_15703,N_14359);
and U20450 (N_20450,N_17574,N_12693);
and U20451 (N_20451,N_17119,N_16972);
xnor U20452 (N_20452,N_17620,N_18497);
xor U20453 (N_20453,N_12941,N_12745);
nor U20454 (N_20454,N_17935,N_14216);
nor U20455 (N_20455,N_16734,N_17266);
nand U20456 (N_20456,N_16857,N_17350);
nand U20457 (N_20457,N_18190,N_15126);
or U20458 (N_20458,N_16822,N_14668);
nor U20459 (N_20459,N_14523,N_12822);
nand U20460 (N_20460,N_16748,N_18106);
and U20461 (N_20461,N_16244,N_12626);
xnor U20462 (N_20462,N_18427,N_17156);
nand U20463 (N_20463,N_14211,N_15153);
and U20464 (N_20464,N_17552,N_15098);
nand U20465 (N_20465,N_16055,N_18150);
xnor U20466 (N_20466,N_16694,N_15224);
nor U20467 (N_20467,N_17108,N_15039);
or U20468 (N_20468,N_13236,N_18165);
nand U20469 (N_20469,N_17138,N_12687);
nand U20470 (N_20470,N_13419,N_14399);
nand U20471 (N_20471,N_13835,N_12895);
nor U20472 (N_20472,N_14279,N_17864);
or U20473 (N_20473,N_13910,N_14218);
nand U20474 (N_20474,N_15893,N_17092);
nor U20475 (N_20475,N_14594,N_17491);
and U20476 (N_20476,N_14851,N_15764);
nand U20477 (N_20477,N_13264,N_18091);
and U20478 (N_20478,N_15434,N_17238);
xor U20479 (N_20479,N_13804,N_18320);
nand U20480 (N_20480,N_17168,N_17493);
or U20481 (N_20481,N_14867,N_15663);
or U20482 (N_20482,N_15430,N_17722);
nor U20483 (N_20483,N_13987,N_17942);
or U20484 (N_20484,N_17646,N_16191);
nand U20485 (N_20485,N_17621,N_18523);
xnor U20486 (N_20486,N_14440,N_13316);
nand U20487 (N_20487,N_12781,N_12624);
xnor U20488 (N_20488,N_14738,N_16230);
nor U20489 (N_20489,N_12779,N_14975);
and U20490 (N_20490,N_17589,N_15128);
and U20491 (N_20491,N_17662,N_13273);
xor U20492 (N_20492,N_16109,N_15280);
xnor U20493 (N_20493,N_14031,N_18424);
nand U20494 (N_20494,N_15367,N_16989);
xnor U20495 (N_20495,N_18616,N_14244);
nor U20496 (N_20496,N_18281,N_13194);
or U20497 (N_20497,N_15607,N_13397);
nor U20498 (N_20498,N_16069,N_15918);
xor U20499 (N_20499,N_17365,N_17093);
and U20500 (N_20500,N_12987,N_14412);
nor U20501 (N_20501,N_16241,N_16180);
xor U20502 (N_20502,N_15790,N_18086);
or U20503 (N_20503,N_15815,N_14669);
or U20504 (N_20504,N_12906,N_15603);
nand U20505 (N_20505,N_14493,N_13564);
nor U20506 (N_20506,N_14896,N_14961);
or U20507 (N_20507,N_13280,N_12669);
and U20508 (N_20508,N_13969,N_14452);
or U20509 (N_20509,N_18485,N_15071);
nor U20510 (N_20510,N_18308,N_17383);
nor U20511 (N_20511,N_16967,N_14091);
and U20512 (N_20512,N_12539,N_18036);
nor U20513 (N_20513,N_14378,N_12921);
xnor U20514 (N_20514,N_17858,N_18072);
and U20515 (N_20515,N_18663,N_14355);
xor U20516 (N_20516,N_14178,N_12582);
and U20517 (N_20517,N_13068,N_16462);
xnor U20518 (N_20518,N_14574,N_18655);
or U20519 (N_20519,N_16758,N_14955);
or U20520 (N_20520,N_18738,N_16248);
nand U20521 (N_20521,N_12924,N_15973);
nand U20522 (N_20522,N_13046,N_13220);
nand U20523 (N_20523,N_17051,N_15696);
nor U20524 (N_20524,N_14825,N_14007);
xnor U20525 (N_20525,N_15504,N_13623);
and U20526 (N_20526,N_18510,N_15263);
nand U20527 (N_20527,N_18487,N_18234);
and U20528 (N_20528,N_15643,N_15676);
and U20529 (N_20529,N_16300,N_13086);
xnor U20530 (N_20530,N_14342,N_16194);
and U20531 (N_20531,N_16982,N_12581);
xor U20532 (N_20532,N_15342,N_17421);
nand U20533 (N_20533,N_18547,N_16914);
and U20534 (N_20534,N_18618,N_17334);
xnor U20535 (N_20535,N_16467,N_17400);
nor U20536 (N_20536,N_15077,N_18233);
or U20537 (N_20537,N_14287,N_12805);
xor U20538 (N_20538,N_16571,N_16147);
or U20539 (N_20539,N_13347,N_13662);
xnor U20540 (N_20540,N_12900,N_15587);
or U20541 (N_20541,N_13193,N_16695);
and U20542 (N_20542,N_17432,N_12565);
nand U20543 (N_20543,N_13707,N_18386);
nand U20544 (N_20544,N_17796,N_16025);
or U20545 (N_20545,N_18696,N_18626);
nand U20546 (N_20546,N_14154,N_18624);
and U20547 (N_20547,N_14963,N_18378);
xor U20548 (N_20548,N_14046,N_12787);
or U20549 (N_20549,N_14533,N_15954);
nor U20550 (N_20550,N_15515,N_14827);
and U20551 (N_20551,N_17137,N_18737);
or U20552 (N_20552,N_12699,N_12883);
nor U20553 (N_20553,N_12837,N_16304);
xnor U20554 (N_20554,N_14052,N_13511);
nand U20555 (N_20555,N_12625,N_16259);
or U20556 (N_20556,N_13309,N_12707);
nor U20557 (N_20557,N_14976,N_14581);
nor U20558 (N_20558,N_16064,N_18073);
nand U20559 (N_20559,N_17632,N_17326);
xnor U20560 (N_20560,N_16211,N_14661);
and U20561 (N_20561,N_15253,N_14971);
nor U20562 (N_20562,N_15725,N_17172);
or U20563 (N_20563,N_15435,N_16536);
xnor U20564 (N_20564,N_18094,N_14776);
or U20565 (N_20565,N_13126,N_13060);
or U20566 (N_20566,N_18683,N_17019);
and U20567 (N_20567,N_15415,N_15008);
xor U20568 (N_20568,N_13402,N_15212);
nor U20569 (N_20569,N_12668,N_15501);
nor U20570 (N_20570,N_18379,N_14490);
or U20571 (N_20571,N_15353,N_18285);
or U20572 (N_20572,N_12768,N_13004);
or U20573 (N_20573,N_13157,N_13228);
nand U20574 (N_20574,N_15089,N_14246);
and U20575 (N_20575,N_15027,N_16518);
xor U20576 (N_20576,N_14274,N_15720);
xor U20577 (N_20577,N_15407,N_14843);
xnor U20578 (N_20578,N_14173,N_16864);
and U20579 (N_20579,N_16421,N_15399);
and U20580 (N_20580,N_18131,N_18435);
or U20581 (N_20581,N_16176,N_15993);
and U20582 (N_20582,N_12510,N_17441);
nand U20583 (N_20583,N_14813,N_13184);
xnor U20584 (N_20584,N_15634,N_17053);
or U20585 (N_20585,N_16150,N_17827);
and U20586 (N_20586,N_13014,N_12848);
and U20587 (N_20587,N_13059,N_17296);
nor U20588 (N_20588,N_15552,N_18305);
and U20589 (N_20589,N_15868,N_14747);
nor U20590 (N_20590,N_18355,N_18309);
nor U20591 (N_20591,N_13551,N_13198);
or U20592 (N_20592,N_15267,N_16729);
nor U20593 (N_20593,N_13784,N_14226);
or U20594 (N_20594,N_17727,N_17268);
and U20595 (N_20595,N_16698,N_17035);
nand U20596 (N_20596,N_12782,N_15919);
and U20597 (N_20597,N_14082,N_16539);
or U20598 (N_20598,N_13613,N_13104);
and U20599 (N_20599,N_15045,N_15474);
or U20600 (N_20600,N_15988,N_18463);
nand U20601 (N_20601,N_16590,N_12713);
or U20602 (N_20602,N_15995,N_18118);
and U20603 (N_20603,N_14105,N_13241);
and U20604 (N_20604,N_14298,N_14263);
nor U20605 (N_20605,N_17018,N_13522);
or U20606 (N_20606,N_16637,N_17516);
and U20607 (N_20607,N_17199,N_12550);
nor U20608 (N_20608,N_15225,N_16697);
or U20609 (N_20609,N_14693,N_18726);
nor U20610 (N_20610,N_14097,N_18269);
and U20611 (N_20611,N_15927,N_18292);
nand U20612 (N_20612,N_17539,N_16220);
and U20613 (N_20613,N_15863,N_16334);
or U20614 (N_20614,N_16993,N_18564);
nor U20615 (N_20615,N_14310,N_13423);
nor U20616 (N_20616,N_16206,N_16407);
and U20617 (N_20617,N_16699,N_13474);
and U20618 (N_20618,N_13296,N_12948);
and U20619 (N_20619,N_16422,N_12642);
xnor U20620 (N_20620,N_15661,N_17110);
xor U20621 (N_20621,N_15481,N_16357);
xnor U20622 (N_20622,N_14352,N_12729);
nand U20623 (N_20623,N_15356,N_15857);
xor U20624 (N_20624,N_14655,N_15466);
nor U20625 (N_20625,N_14609,N_15495);
xnor U20626 (N_20626,N_17913,N_15183);
and U20627 (N_20627,N_14329,N_16175);
xor U20628 (N_20628,N_17532,N_14353);
or U20629 (N_20629,N_14641,N_18069);
and U20630 (N_20630,N_16626,N_15548);
or U20631 (N_20631,N_18725,N_13183);
and U20632 (N_20632,N_18718,N_16344);
xnor U20633 (N_20633,N_16937,N_16213);
or U20634 (N_20634,N_17946,N_16709);
or U20635 (N_20635,N_18155,N_13806);
or U20636 (N_20636,N_14357,N_16093);
and U20637 (N_20637,N_14437,N_18338);
xor U20638 (N_20638,N_12785,N_16136);
nand U20639 (N_20639,N_16559,N_15009);
or U20640 (N_20640,N_13523,N_15867);
nand U20641 (N_20641,N_16715,N_17086);
xnor U20642 (N_20642,N_14278,N_14029);
xor U20643 (N_20643,N_14573,N_18092);
xor U20644 (N_20644,N_16956,N_17637);
nor U20645 (N_20645,N_13927,N_12788);
nand U20646 (N_20646,N_13611,N_12954);
nand U20647 (N_20647,N_13739,N_16054);
nand U20648 (N_20648,N_13726,N_17916);
nand U20649 (N_20649,N_12530,N_13400);
nand U20650 (N_20650,N_13480,N_12592);
nor U20651 (N_20651,N_17953,N_12619);
and U20652 (N_20652,N_17786,N_14797);
and U20653 (N_20653,N_13698,N_14708);
and U20654 (N_20654,N_17698,N_14400);
nand U20655 (N_20655,N_17328,N_16872);
nor U20656 (N_20656,N_13307,N_18664);
xor U20657 (N_20657,N_15851,N_15288);
xor U20658 (N_20658,N_16290,N_15838);
or U20659 (N_20659,N_17910,N_18140);
and U20660 (N_20660,N_13636,N_17701);
or U20661 (N_20661,N_13451,N_14047);
nand U20662 (N_20662,N_16861,N_13226);
nand U20663 (N_20663,N_14086,N_13637);
or U20664 (N_20664,N_16531,N_18179);
nor U20665 (N_20665,N_14404,N_15500);
xor U20666 (N_20666,N_15828,N_14530);
nand U20667 (N_20667,N_16629,N_14892);
nand U20668 (N_20668,N_16870,N_18539);
and U20669 (N_20669,N_16886,N_14769);
xnor U20670 (N_20670,N_14782,N_18139);
nor U20671 (N_20671,N_15331,N_14973);
nand U20672 (N_20672,N_13687,N_14318);
and U20673 (N_20673,N_15771,N_17984);
nand U20674 (N_20674,N_18263,N_17152);
or U20675 (N_20675,N_15724,N_13213);
nand U20676 (N_20676,N_15145,N_17345);
or U20677 (N_20677,N_12684,N_13343);
and U20678 (N_20678,N_18588,N_17272);
and U20679 (N_20679,N_12628,N_15582);
nor U20680 (N_20680,N_15254,N_17708);
xor U20681 (N_20681,N_17665,N_17504);
nand U20682 (N_20682,N_17403,N_12548);
nand U20683 (N_20683,N_12965,N_17880);
and U20684 (N_20684,N_12867,N_17352);
nor U20685 (N_20685,N_18467,N_16096);
xor U20686 (N_20686,N_18163,N_18466);
and U20687 (N_20687,N_16712,N_16400);
and U20688 (N_20688,N_13133,N_13565);
nor U20689 (N_20689,N_17445,N_17923);
or U20690 (N_20690,N_18288,N_14682);
and U20691 (N_20691,N_18384,N_16958);
or U20692 (N_20692,N_17200,N_18232);
and U20693 (N_20693,N_18651,N_18367);
xor U20694 (N_20694,N_15237,N_17286);
or U20695 (N_20695,N_14715,N_15179);
xnor U20696 (N_20696,N_17957,N_13021);
and U20697 (N_20697,N_16201,N_14512);
xnor U20698 (N_20698,N_13498,N_13131);
or U20699 (N_20699,N_14093,N_17821);
xnor U20700 (N_20700,N_17740,N_18498);
and U20701 (N_20701,N_16501,N_13776);
xor U20702 (N_20702,N_14032,N_15059);
nor U20703 (N_20703,N_14176,N_17333);
xor U20704 (N_20704,N_12737,N_14645);
nand U20705 (N_20705,N_18495,N_13619);
xor U20706 (N_20706,N_12743,N_14722);
or U20707 (N_20707,N_13132,N_14796);
nand U20708 (N_20708,N_17079,N_13572);
xnor U20709 (N_20709,N_15287,N_16753);
nor U20710 (N_20710,N_14286,N_17717);
nand U20711 (N_20711,N_17198,N_17856);
xnor U20712 (N_20712,N_14039,N_18434);
xnor U20713 (N_20713,N_18406,N_17074);
and U20714 (N_20714,N_16570,N_12996);
nand U20715 (N_20715,N_15160,N_15543);
nand U20716 (N_20716,N_18209,N_15093);
nand U20717 (N_20717,N_16114,N_14159);
nor U20718 (N_20718,N_16408,N_17885);
nand U20719 (N_20719,N_17159,N_18192);
nand U20720 (N_20720,N_13012,N_13896);
or U20721 (N_20721,N_14907,N_13412);
xnor U20722 (N_20722,N_12791,N_15198);
and U20723 (N_20723,N_14470,N_15760);
nor U20724 (N_20724,N_15709,N_13749);
xnor U20725 (N_20725,N_14727,N_13310);
xor U20726 (N_20726,N_18206,N_15573);
xnor U20727 (N_20727,N_15035,N_14309);
nand U20728 (N_20728,N_13093,N_17353);
xnor U20729 (N_20729,N_18730,N_13170);
nand U20730 (N_20730,N_15105,N_12937);
nand U20731 (N_20731,N_14730,N_17929);
nand U20732 (N_20732,N_17372,N_14852);
xor U20733 (N_20733,N_16277,N_14555);
xnor U20734 (N_20734,N_15482,N_16624);
nand U20735 (N_20735,N_14949,N_14049);
nor U20736 (N_20736,N_16018,N_17187);
xnor U20737 (N_20737,N_14664,N_14526);
xnor U20738 (N_20738,N_18613,N_13610);
and U20739 (N_20739,N_16458,N_16133);
nor U20740 (N_20740,N_17130,N_14311);
and U20741 (N_20741,N_12828,N_17988);
nor U20742 (N_20742,N_17711,N_18721);
nor U20743 (N_20743,N_12945,N_15141);
and U20744 (N_20744,N_14051,N_14036);
and U20745 (N_20745,N_14252,N_17175);
nand U20746 (N_20746,N_14422,N_17951);
and U20747 (N_20747,N_16569,N_16558);
or U20748 (N_20748,N_18551,N_12616);
nor U20749 (N_20749,N_17181,N_13368);
nand U20750 (N_20750,N_14106,N_16896);
nand U20751 (N_20751,N_12845,N_16354);
or U20752 (N_20752,N_13981,N_15689);
nor U20753 (N_20753,N_15742,N_13144);
xor U20754 (N_20754,N_17037,N_12875);
xor U20755 (N_20755,N_18221,N_17735);
and U20756 (N_20756,N_17009,N_15156);
or U20757 (N_20757,N_13785,N_18516);
or U20758 (N_20758,N_17654,N_15282);
nor U20759 (N_20759,N_14472,N_14720);
or U20760 (N_20760,N_14464,N_18641);
nand U20761 (N_20761,N_16035,N_16276);
nand U20762 (N_20762,N_13278,N_16811);
and U20763 (N_20763,N_15441,N_17718);
nor U20764 (N_20764,N_14240,N_15556);
xor U20765 (N_20765,N_16369,N_15523);
nand U20766 (N_20766,N_17057,N_16818);
or U20767 (N_20767,N_13532,N_16101);
nand U20768 (N_20768,N_14613,N_18397);
nand U20769 (N_20769,N_17264,N_16003);
nor U20770 (N_20770,N_15631,N_13127);
nor U20771 (N_20771,N_15766,N_13587);
xnor U20772 (N_20772,N_17595,N_14127);
or U20773 (N_20773,N_17307,N_15765);
and U20774 (N_20774,N_15982,N_16964);
and U20775 (N_20775,N_17376,N_17358);
nor U20776 (N_20776,N_14956,N_17917);
nand U20777 (N_20777,N_18193,N_17270);
or U20778 (N_20778,N_18197,N_18422);
xor U20779 (N_20779,N_13681,N_13686);
and U20780 (N_20780,N_15297,N_13957);
xnor U20781 (N_20781,N_13872,N_16039);
nor U20782 (N_20782,N_15717,N_15712);
or U20783 (N_20783,N_17517,N_17229);
nor U20784 (N_20784,N_14771,N_17616);
and U20785 (N_20785,N_13916,N_18614);
nor U20786 (N_20786,N_16727,N_14186);
xor U20787 (N_20787,N_13942,N_13168);
nor U20788 (N_20788,N_17301,N_16639);
xor U20789 (N_20789,N_16470,N_15175);
and U20790 (N_20790,N_13490,N_13539);
nor U20791 (N_20791,N_17560,N_18315);
and U20792 (N_20792,N_15409,N_12545);
nand U20793 (N_20793,N_13740,N_16336);
nor U20794 (N_20794,N_16432,N_17640);
or U20795 (N_20795,N_13868,N_17252);
or U20796 (N_20796,N_14532,N_14937);
nand U20797 (N_20797,N_16454,N_13025);
xor U20798 (N_20798,N_18519,N_16493);
or U20799 (N_20799,N_12501,N_17934);
xor U20800 (N_20800,N_17438,N_18488);
and U20801 (N_20801,N_17738,N_15579);
nor U20802 (N_20802,N_17139,N_13632);
or U20803 (N_20803,N_16137,N_17680);
xor U20804 (N_20804,N_17593,N_14088);
nand U20805 (N_20805,N_15290,N_17015);
nor U20806 (N_20806,N_13992,N_14578);
xor U20807 (N_20807,N_15911,N_16903);
nand U20808 (N_20808,N_16960,N_17465);
or U20809 (N_20809,N_13495,N_14331);
or U20810 (N_20810,N_17380,N_13246);
or U20811 (N_20811,N_15091,N_14230);
or U20812 (N_20812,N_14385,N_14644);
and U20813 (N_20813,N_16505,N_13222);
xor U20814 (N_20814,N_13274,N_13527);
and U20815 (N_20815,N_14044,N_18710);
and U20816 (N_20816,N_13460,N_15438);
xnor U20817 (N_20817,N_14260,N_12757);
or U20818 (N_20818,N_18211,N_17684);
nor U20819 (N_20819,N_15286,N_18451);
xnor U20820 (N_20820,N_15364,N_16262);
nand U20821 (N_20821,N_15496,N_18214);
and U20822 (N_20822,N_12632,N_13833);
xnor U20823 (N_20823,N_12557,N_13671);
and U20824 (N_20824,N_17520,N_14306);
or U20825 (N_20825,N_14610,N_14729);
or U20826 (N_20826,N_16361,N_14958);
nand U20827 (N_20827,N_16548,N_17794);
nor U20828 (N_20828,N_18371,N_13903);
and U20829 (N_20829,N_15301,N_14135);
and U20830 (N_20830,N_17567,N_15248);
or U20831 (N_20831,N_14416,N_17386);
or U20832 (N_20832,N_16090,N_14621);
and U20833 (N_20833,N_15099,N_12907);
or U20834 (N_20834,N_13022,N_15137);
xnor U20835 (N_20835,N_13404,N_17254);
nand U20836 (N_20836,N_17176,N_13919);
and U20837 (N_20837,N_14478,N_16530);
or U20838 (N_20838,N_17319,N_15834);
xnor U20839 (N_20839,N_15371,N_12999);
nand U20840 (N_20840,N_12859,N_16844);
xnor U20841 (N_20841,N_17981,N_13250);
xor U20842 (N_20842,N_16433,N_13932);
or U20843 (N_20843,N_14864,N_16942);
nand U20844 (N_20844,N_16762,N_17674);
xnor U20845 (N_20845,N_18415,N_12793);
and U20846 (N_20846,N_15142,N_16479);
nand U20847 (N_20847,N_13097,N_15013);
or U20848 (N_20848,N_15423,N_13781);
nand U20849 (N_20849,N_13628,N_12686);
xnor U20850 (N_20850,N_16534,N_14024);
and U20851 (N_20851,N_17655,N_15726);
nand U20852 (N_20852,N_13067,N_18349);
nor U20853 (N_20853,N_18628,N_16827);
nor U20854 (N_20854,N_12928,N_14247);
and U20855 (N_20855,N_17804,N_14537);
and U20856 (N_20856,N_15056,N_15854);
or U20857 (N_20857,N_16346,N_18460);
and U20858 (N_20858,N_17889,N_16573);
or U20859 (N_20859,N_17576,N_15223);
and U20860 (N_20860,N_15322,N_12955);
or U20861 (N_20861,N_17483,N_12560);
xnor U20862 (N_20862,N_16506,N_12552);
nand U20863 (N_20863,N_15810,N_17972);
or U20864 (N_20864,N_17579,N_15618);
nand U20865 (N_20865,N_14447,N_13105);
or U20866 (N_20866,N_13538,N_18004);
xor U20867 (N_20867,N_17474,N_13945);
and U20868 (N_20868,N_14614,N_17029);
xor U20869 (N_20869,N_14724,N_17436);
nand U20870 (N_20870,N_16396,N_15571);
nand U20871 (N_20871,N_12854,N_14128);
xnor U20872 (N_20872,N_17324,N_17030);
xor U20873 (N_20873,N_15115,N_12708);
and U20874 (N_20874,N_15333,N_13569);
xor U20875 (N_20875,N_16209,N_13163);
or U20876 (N_20876,N_14631,N_14779);
nand U20877 (N_20877,N_18736,N_17915);
or U20878 (N_20878,N_16074,N_13312);
xor U20879 (N_20879,N_17003,N_18301);
xor U20880 (N_20880,N_12593,N_17415);
and U20881 (N_20881,N_13618,N_14293);
xor U20882 (N_20882,N_17497,N_13600);
or U20883 (N_20883,N_12969,N_17982);
and U20884 (N_20884,N_13704,N_18462);
nor U20885 (N_20885,N_13078,N_18120);
and U20886 (N_20886,N_16326,N_13958);
or U20887 (N_20887,N_14498,N_15401);
and U20888 (N_20888,N_14391,N_13660);
and U20889 (N_20889,N_18394,N_12603);
and U20890 (N_20890,N_15007,N_18401);
nor U20891 (N_20891,N_15594,N_16798);
xnor U20892 (N_20892,N_13418,N_14774);
xor U20893 (N_20893,N_16866,N_13079);
or U20894 (N_20894,N_18037,N_15852);
nand U20895 (N_20895,N_12998,N_16409);
nand U20896 (N_20896,N_15432,N_17122);
nor U20897 (N_20897,N_17663,N_15902);
xnor U20898 (N_20898,N_15425,N_17221);
nand U20899 (N_20899,N_16645,N_13290);
nor U20900 (N_20900,N_17095,N_17185);
and U20901 (N_20901,N_13956,N_18055);
or U20902 (N_20902,N_16405,N_17406);
or U20903 (N_20903,N_18226,N_17777);
nand U20904 (N_20904,N_13657,N_18493);
xnor U20905 (N_20905,N_13664,N_15625);
or U20906 (N_20906,N_16274,N_15209);
nor U20907 (N_20907,N_12769,N_15791);
xor U20908 (N_20908,N_15406,N_15855);
and U20909 (N_20909,N_12886,N_14845);
nand U20910 (N_20910,N_17728,N_13066);
and U20911 (N_20911,N_13850,N_16263);
and U20912 (N_20912,N_16189,N_16549);
nand U20913 (N_20913,N_17293,N_15050);
nand U20914 (N_20914,N_17789,N_15246);
xor U20915 (N_20915,N_16456,N_17550);
nand U20916 (N_20916,N_13631,N_14739);
xnor U20917 (N_20917,N_13234,N_15965);
xnor U20918 (N_20918,N_14689,N_14781);
xor U20919 (N_20919,N_17094,N_14684);
xor U20920 (N_20920,N_13101,N_15768);
and U20921 (N_20921,N_17100,N_14649);
xor U20922 (N_20922,N_16999,N_17941);
nor U20923 (N_20923,N_18215,N_13407);
or U20924 (N_20924,N_17305,N_13940);
or U20925 (N_20925,N_17558,N_14605);
or U20926 (N_20926,N_16120,N_15874);
nand U20927 (N_20927,N_14426,N_17851);
or U20928 (N_20928,N_15925,N_17429);
xor U20929 (N_20929,N_17603,N_15783);
and U20930 (N_20930,N_14334,N_16733);
or U20931 (N_20931,N_17223,N_14095);
nand U20932 (N_20932,N_16922,N_14122);
nand U20933 (N_20933,N_15258,N_14108);
or U20934 (N_20934,N_14770,N_16303);
nand U20935 (N_20935,N_16331,N_13477);
nand U20936 (N_20936,N_17952,N_17653);
or U20937 (N_20937,N_17673,N_15195);
nor U20938 (N_20938,N_15774,N_18694);
or U20939 (N_20939,N_15316,N_13596);
xnor U20940 (N_20940,N_15387,N_15668);
and U20941 (N_20941,N_12712,N_13753);
and U20942 (N_20942,N_17171,N_15507);
nor U20943 (N_20943,N_17977,N_14835);
and U20944 (N_20944,N_12739,N_14552);
and U20945 (N_20945,N_18229,N_12961);
or U20946 (N_20946,N_15861,N_14967);
or U20947 (N_20947,N_17277,N_14070);
xor U20948 (N_20948,N_18690,N_17522);
and U20949 (N_20949,N_16648,N_13905);
or U20950 (N_20950,N_14808,N_17720);
nand U20951 (N_20951,N_12877,N_13255);
nor U20952 (N_20952,N_15082,N_15067);
nand U20953 (N_20953,N_13286,N_15234);
nor U20954 (N_20954,N_18031,N_17530);
and U20955 (N_20955,N_16437,N_17872);
nand U20956 (N_20956,N_12947,N_16330);
nor U20957 (N_20957,N_15110,N_18711);
or U20958 (N_20958,N_18503,N_14562);
nand U20959 (N_20959,N_12936,N_13393);
and U20960 (N_20960,N_17027,N_17507);
nand U20961 (N_20961,N_13192,N_14380);
and U20962 (N_20962,N_17690,N_15335);
xnor U20963 (N_20963,N_16112,N_14077);
nor U20964 (N_20964,N_17315,N_15641);
and U20965 (N_20965,N_16001,N_14656);
nand U20966 (N_20966,N_17125,N_18548);
xor U20967 (N_20967,N_13625,N_14322);
nor U20968 (N_20968,N_12891,N_17336);
nand U20969 (N_20969,N_16681,N_17486);
nor U20970 (N_20970,N_17310,N_13367);
or U20971 (N_20971,N_18224,N_16988);
or U20972 (N_20972,N_15394,N_16038);
nor U20973 (N_20973,N_14308,N_13219);
and U20974 (N_20974,N_16684,N_15229);
xor U20975 (N_20975,N_13440,N_16097);
or U20976 (N_20976,N_13003,N_18675);
or U20977 (N_20977,N_15800,N_14060);
xor U20978 (N_20978,N_14403,N_15439);
or U20979 (N_20979,N_17998,N_16086);
and U20980 (N_20980,N_14301,N_18303);
and U20981 (N_20981,N_13879,N_13361);
nand U20982 (N_20982,N_14148,N_16363);
nand U20983 (N_20983,N_16430,N_15513);
nor U20984 (N_20984,N_14647,N_14479);
xnor U20985 (N_20985,N_13814,N_12637);
or U20986 (N_20986,N_14841,N_12500);
or U20987 (N_20987,N_12819,N_15898);
nor U20988 (N_20988,N_17598,N_15125);
or U20989 (N_20989,N_15991,N_17348);
nand U20990 (N_20990,N_17256,N_12685);
nor U20991 (N_20991,N_17395,N_17251);
nor U20992 (N_20992,N_18561,N_13573);
nor U20993 (N_20993,N_13293,N_12507);
or U20994 (N_20994,N_16923,N_18261);
and U20995 (N_20995,N_13196,N_15026);
and U20996 (N_20996,N_17541,N_13201);
nand U20997 (N_20997,N_15622,N_16944);
xnor U20998 (N_20998,N_12633,N_18294);
or U20999 (N_20999,N_17859,N_15152);
and U21000 (N_21000,N_13496,N_15581);
xnor U21001 (N_21001,N_13859,N_12802);
and U21002 (N_21002,N_18481,N_13897);
xor U21003 (N_21003,N_17836,N_15123);
nand U21004 (N_21004,N_13142,N_18195);
nor U21005 (N_21005,N_14891,N_12956);
and U21006 (N_21006,N_13699,N_17312);
or U21007 (N_21007,N_17127,N_14687);
nor U21008 (N_21008,N_16883,N_17287);
or U21009 (N_21009,N_16520,N_16461);
and U21010 (N_21010,N_16394,N_14023);
nand U21011 (N_21011,N_17511,N_16171);
nor U21012 (N_21012,N_15670,N_15031);
nor U21013 (N_21013,N_15193,N_16239);
xnor U21014 (N_21014,N_14917,N_17112);
nor U21015 (N_21015,N_15584,N_13727);
nand U21016 (N_21016,N_12905,N_15426);
nand U21017 (N_21017,N_15456,N_18509);
or U21018 (N_21018,N_15592,N_16713);
nor U21019 (N_21019,N_16672,N_14053);
xor U21020 (N_21020,N_16612,N_16362);
or U21021 (N_21021,N_17116,N_14823);
nor U21022 (N_21022,N_18654,N_14734);
and U21023 (N_21023,N_17792,N_18700);
nand U21024 (N_21024,N_18719,N_16162);
nand U21025 (N_21025,N_17117,N_12551);
and U21026 (N_21026,N_18076,N_16089);
nand U21027 (N_21027,N_13557,N_13099);
xnor U21028 (N_21028,N_18132,N_13741);
and U21029 (N_21029,N_16722,N_16591);
nand U21030 (N_21030,N_14264,N_15214);
nor U21031 (N_21031,N_17839,N_18342);
nand U21032 (N_21032,N_18085,N_16535);
nand U21033 (N_21033,N_14577,N_13057);
xnor U21034 (N_21034,N_13871,N_13386);
and U21035 (N_21035,N_16068,N_16948);
xnor U21036 (N_21036,N_18191,N_13146);
nor U21037 (N_21037,N_16072,N_14784);
or U21038 (N_21038,N_16052,N_13828);
nand U21039 (N_21039,N_16710,N_14912);
nor U21040 (N_21040,N_12623,N_17602);
nand U21041 (N_21041,N_14801,N_15616);
nand U21042 (N_21042,N_17610,N_17207);
nor U21043 (N_21043,N_13034,N_13697);
or U21044 (N_21044,N_15252,N_15429);
nand U21045 (N_21045,N_18609,N_16444);
xnor U21046 (N_21046,N_16754,N_12615);
xor U21047 (N_21047,N_15751,N_17968);
xnor U21048 (N_21048,N_13429,N_16537);
or U21049 (N_21049,N_15778,N_15930);
and U21050 (N_21050,N_14856,N_14705);
nand U21051 (N_21051,N_16507,N_17623);
or U21052 (N_21052,N_17896,N_17265);
and U21053 (N_21053,N_13471,N_12614);
or U21054 (N_21054,N_17918,N_13678);
or U21055 (N_21055,N_15230,N_15347);
nor U21056 (N_21056,N_15185,N_14008);
xor U21057 (N_21057,N_15511,N_14022);
or U21058 (N_21058,N_14381,N_16572);
xor U21059 (N_21059,N_14861,N_15745);
and U21060 (N_21060,N_18698,N_13936);
or U21061 (N_21061,N_13210,N_18194);
or U21062 (N_21062,N_17919,N_17891);
nand U21063 (N_21063,N_12978,N_14141);
nor U21064 (N_21064,N_12654,N_16766);
nor U21065 (N_21065,N_15015,N_15365);
xnor U21066 (N_21066,N_13769,N_18395);
or U21067 (N_21067,N_14822,N_17154);
nand U21068 (N_21068,N_18185,N_17533);
and U21069 (N_21069,N_18218,N_14480);
and U21070 (N_21070,N_18702,N_17514);
nor U21071 (N_21071,N_17760,N_15291);
nor U21072 (N_21072,N_17224,N_13725);
nor U21073 (N_21073,N_14889,N_17772);
nor U21074 (N_21074,N_15728,N_17641);
xor U21075 (N_21075,N_15162,N_18188);
nand U21076 (N_21076,N_14657,N_13537);
nor U21077 (N_21077,N_13609,N_13074);
nand U21078 (N_21078,N_14067,N_14648);
xnor U21079 (N_21079,N_14345,N_15148);
nor U21080 (N_21080,N_13377,N_18112);
and U21081 (N_21081,N_12517,N_16778);
nor U21082 (N_21082,N_13549,N_14583);
xor U21083 (N_21083,N_17776,N_15232);
xnor U21084 (N_21084,N_15623,N_15983);
xor U21085 (N_21085,N_14313,N_13129);
and U21086 (N_21086,N_13614,N_16653);
and U21087 (N_21087,N_13694,N_14415);
xnor U21088 (N_21088,N_17162,N_17431);
nor U21089 (N_21089,N_14418,N_14944);
xnor U21090 (N_21090,N_16936,N_14056);
xnor U21091 (N_21091,N_18098,N_14134);
nand U21092 (N_21092,N_13475,N_17960);
nand U21093 (N_21093,N_14984,N_15187);
nor U21094 (N_21094,N_14193,N_13091);
nor U21095 (N_21095,N_14273,N_16016);
xnor U21096 (N_21096,N_16391,N_17024);
nand U21097 (N_21097,N_14160,N_18032);
nand U21098 (N_21098,N_15944,N_14791);
nor U21099 (N_21099,N_14179,N_12852);
or U21100 (N_21100,N_14717,N_18671);
or U21101 (N_21101,N_17756,N_16940);
nand U21102 (N_21102,N_18026,N_18448);
and U21103 (N_21103,N_15633,N_18343);
nor U21104 (N_21104,N_16825,N_13218);
and U21105 (N_21105,N_12672,N_17361);
and U21106 (N_21106,N_14507,N_16985);
and U21107 (N_21107,N_15359,N_13824);
nor U21108 (N_21108,N_17146,N_16532);
or U21109 (N_21109,N_16024,N_14788);
and U21110 (N_21110,N_18550,N_13128);
and U21111 (N_21111,N_15354,N_15010);
nand U21112 (N_21112,N_13768,N_14411);
and U21113 (N_21113,N_14741,N_14042);
or U21114 (N_21114,N_14904,N_18002);
nand U21115 (N_21115,N_15517,N_15226);
or U21116 (N_21116,N_18300,N_17070);
nand U21117 (N_21117,N_16132,N_17487);
xor U21118 (N_21118,N_12876,N_14570);
or U21119 (N_21119,N_13261,N_14625);
nor U21120 (N_21120,N_16251,N_13921);
or U21121 (N_21121,N_17023,N_15671);
xnor U21122 (N_21122,N_14455,N_14195);
nor U21123 (N_21123,N_14908,N_18715);
and U21124 (N_21124,N_18398,N_16819);
or U21125 (N_21125,N_17608,N_13949);
and U21126 (N_21126,N_15963,N_17389);
xor U21127 (N_21127,N_13039,N_13773);
nor U21128 (N_21128,N_13643,N_13544);
xnor U21129 (N_21129,N_17703,N_18438);
nor U21130 (N_21130,N_17733,N_13502);
xnor U21131 (N_21131,N_13342,N_13622);
xnor U21132 (N_21132,N_17790,N_18272);
or U21133 (N_21133,N_14126,N_16260);
nand U21134 (N_21134,N_15163,N_14842);
nand U21135 (N_21135,N_14991,N_18370);
xnor U21136 (N_21136,N_14428,N_14430);
xnor U21137 (N_21137,N_17822,N_14364);
nand U21138 (N_21138,N_12696,N_13579);
nand U21139 (N_21139,N_13889,N_14900);
nand U21140 (N_21140,N_17191,N_17166);
xnor U21141 (N_21141,N_12990,N_13996);
and U21142 (N_21142,N_15756,N_18024);
nand U21143 (N_21143,N_15968,N_14212);
nor U21144 (N_21144,N_18703,N_13514);
xnor U21145 (N_21145,N_13943,N_14660);
or U21146 (N_21146,N_13629,N_16223);
nand U21147 (N_21147,N_13466,N_16933);
nor U21148 (N_21148,N_15583,N_13696);
xor U21149 (N_21149,N_17145,N_14686);
nor U21150 (N_21150,N_13570,N_16232);
nor U21151 (N_21151,N_12656,N_16987);
or U21152 (N_21152,N_13405,N_17331);
or U21153 (N_21153,N_13911,N_13169);
and U21154 (N_21154,N_13808,N_14281);
and U21155 (N_21155,N_16219,N_14994);
and U21156 (N_21156,N_13816,N_13685);
and U21157 (N_21157,N_15442,N_18318);
or U21158 (N_21158,N_17250,N_13548);
nand U21159 (N_21159,N_18015,N_14205);
and U21160 (N_21160,N_15884,N_15494);
and U21161 (N_21161,N_17810,N_15334);
or U21162 (N_21162,N_17607,N_17838);
or U21163 (N_21163,N_13967,N_14451);
or U21164 (N_21164,N_14531,N_13973);
xor U21165 (N_21165,N_16384,N_18335);
xor U21166 (N_21166,N_18570,N_18727);
nor U21167 (N_21167,N_13265,N_16595);
xor U21168 (N_21168,N_12992,N_16499);
xnor U21169 (N_21169,N_16971,N_15119);
xnor U21170 (N_21170,N_18266,N_13997);
or U21171 (N_21171,N_18576,N_18639);
nand U21172 (N_21172,N_16436,N_14337);
xnor U21173 (N_21173,N_15651,N_14025);
nand U21174 (N_21174,N_15602,N_17759);
xor U21175 (N_21175,N_13862,N_15598);
and U21176 (N_21176,N_17682,N_13993);
xor U21177 (N_21177,N_17964,N_14291);
and U21178 (N_21178,N_13050,N_16364);
or U21179 (N_21179,N_12943,N_16814);
nand U21180 (N_21180,N_14983,N_12776);
and U21181 (N_21181,N_14858,N_16301);
or U21182 (N_21182,N_15154,N_15636);
or U21183 (N_21183,N_14879,N_17398);
or U21184 (N_21184,N_16714,N_18127);
or U21185 (N_21185,N_16200,N_15388);
and U21186 (N_21186,N_17237,N_13931);
nor U21187 (N_21187,N_12609,N_17479);
xnor U21188 (N_21188,N_13117,N_14972);
nor U21189 (N_21189,N_16719,N_16238);
xnor U21190 (N_21190,N_13462,N_12527);
nand U21191 (N_21191,N_15127,N_15595);
nor U21192 (N_21192,N_18115,N_14793);
or U21193 (N_21193,N_16647,N_16597);
nor U21194 (N_21194,N_14034,N_13162);
and U21195 (N_21195,N_17062,N_17954);
nand U21196 (N_21196,N_15304,N_17604);
or U21197 (N_21197,N_18630,N_13180);
nand U21198 (N_21198,N_16119,N_17679);
nand U21199 (N_21199,N_15075,N_12723);
nor U21200 (N_21200,N_12711,N_14766);
nor U21201 (N_21201,N_16253,N_18602);
nor U21202 (N_21202,N_16604,N_15626);
or U21203 (N_21203,N_13164,N_15741);
nand U21204 (N_21204,N_17606,N_17284);
nor U21205 (N_21205,N_13684,N_13434);
xor U21206 (N_21206,N_16299,N_18258);
xor U21207 (N_21207,N_18486,N_13024);
and U21208 (N_21208,N_14850,N_15655);
nand U21209 (N_21209,N_13232,N_13966);
xnor U21210 (N_21210,N_13791,N_15395);
and U21211 (N_21211,N_18148,N_15627);
or U21212 (N_21212,N_16809,N_12929);
xnor U21213 (N_21213,N_14237,N_15453);
xnor U21214 (N_21214,N_18538,N_12925);
and U21215 (N_21215,N_14829,N_17912);
nand U21216 (N_21216,N_18387,N_16486);
xor U21217 (N_21217,N_13853,N_16780);
or U21218 (N_21218,N_16533,N_14636);
nand U21219 (N_21219,N_15824,N_13803);
or U21220 (N_21220,N_13737,N_12922);
or U21221 (N_21221,N_15079,N_13944);
nand U21222 (N_21222,N_18454,N_18416);
nand U21223 (N_21223,N_17226,N_17834);
nand U21224 (N_21224,N_13257,N_17741);
nor U21225 (N_21225,N_17280,N_12621);
nand U21226 (N_21226,N_16237,N_12866);
xnor U21227 (N_21227,N_17004,N_17464);
and U21228 (N_21228,N_14197,N_17644);
and U21229 (N_21229,N_15389,N_17033);
xor U21230 (N_21230,N_16113,N_16002);
nor U21231 (N_21231,N_13886,N_14295);
nor U21232 (N_21232,N_13984,N_17513);
and U21233 (N_21233,N_12566,N_16051);
xor U21234 (N_21234,N_18364,N_16269);
or U21235 (N_21235,N_15843,N_17274);
or U21236 (N_21236,N_14726,N_14427);
xor U21237 (N_21237,N_16056,N_16085);
nor U21238 (N_21238,N_12892,N_14986);
nand U21239 (N_21239,N_13051,N_17780);
or U21240 (N_21240,N_16282,N_16867);
and U21241 (N_21241,N_17562,N_13870);
or U21242 (N_21242,N_17050,N_17782);
nand U21243 (N_21243,N_17763,N_16046);
nand U21244 (N_21244,N_14725,N_15402);
xnor U21245 (N_21245,N_18622,N_18667);
and U21246 (N_21246,N_13586,N_16782);
xor U21247 (N_21247,N_13583,N_17148);
or U21248 (N_21248,N_16457,N_18035);
nor U21249 (N_21249,N_15369,N_14184);
and U21250 (N_21250,N_14765,N_18135);
nor U21251 (N_21251,N_18403,N_13453);
or U21252 (N_21252,N_13645,N_15273);
or U21253 (N_21253,N_16010,N_13923);
nor U21254 (N_21254,N_16105,N_13961);
or U21255 (N_21255,N_15516,N_14394);
and U21256 (N_21256,N_13428,N_16006);
xnor U21257 (N_21257,N_14267,N_12663);
xor U21258 (N_21258,N_14740,N_15424);
nand U21259 (N_21259,N_17943,N_13055);
nand U21260 (N_21260,N_16455,N_17868);
xor U21261 (N_21261,N_14143,N_16575);
nor U21262 (N_21262,N_15491,N_16856);
or U21263 (N_21263,N_13124,N_13531);
nand U21264 (N_21264,N_15184,N_14396);
and U21265 (N_21265,N_17236,N_16199);
and U21266 (N_21266,N_16821,N_12575);
and U21267 (N_21267,N_14627,N_15695);
nand U21268 (N_21268,N_15576,N_13229);
and U21269 (N_21269,N_16725,N_17088);
xor U21270 (N_21270,N_16185,N_15138);
nand U21271 (N_21271,N_13563,N_15361);
and U21272 (N_21272,N_13759,N_14756);
or U21273 (N_21273,N_16690,N_15470);
and U21274 (N_21274,N_16610,N_18502);
nand U21275 (N_21275,N_14623,N_18723);
xor U21276 (N_21276,N_13627,N_15120);
or U21277 (N_21277,N_13483,N_18039);
nand U21278 (N_21278,N_18283,N_18681);
nand U21279 (N_21279,N_16996,N_15124);
or U21280 (N_21280,N_13364,N_13420);
nand U21281 (N_21281,N_15206,N_12865);
xnor U21282 (N_21282,N_15292,N_17422);
nand U21283 (N_21283,N_15858,N_12736);
and U21284 (N_21284,N_17883,N_15761);
and U21285 (N_21285,N_16492,N_13951);
nor U21286 (N_21286,N_14144,N_17650);
nor U21287 (N_21287,N_17401,N_17812);
nand U21288 (N_21288,N_13339,N_16678);
and U21289 (N_21289,N_17888,N_18271);
nand U21290 (N_21290,N_15310,N_17047);
xor U21291 (N_21291,N_13167,N_16906);
or U21292 (N_21292,N_13642,N_18605);
nor U21293 (N_21293,N_13007,N_13150);
nor U21294 (N_21294,N_15097,N_15266);
and U21295 (N_21295,N_16764,N_18029);
xnor U21296 (N_21296,N_13703,N_18680);
nand U21297 (N_21297,N_13156,N_14457);
nor U21298 (N_21298,N_17870,N_16159);
nor U21299 (N_21299,N_15509,N_14716);
and U21300 (N_21300,N_18512,N_13223);
and U21301 (N_21301,N_18359,N_12887);
and U21302 (N_21302,N_18562,N_16707);
nand U21303 (N_21303,N_18099,N_17390);
or U21304 (N_21304,N_16783,N_14238);
and U21305 (N_21305,N_16319,N_15585);
and U21306 (N_21306,N_18363,N_16959);
or U21307 (N_21307,N_17808,N_18123);
nand U21308 (N_21308,N_18492,N_17045);
xnor U21309 (N_21309,N_18436,N_16483);
or U21310 (N_21310,N_13442,N_17063);
and U21311 (N_21311,N_16613,N_17275);
or U21312 (N_21312,N_12881,N_17664);
nand U21313 (N_21313,N_15738,N_16983);
or U21314 (N_21314,N_15538,N_17450);
and U21315 (N_21315,N_16420,N_14187);
and U21316 (N_21316,N_16125,N_15260);
or U21317 (N_21317,N_17021,N_16383);
xnor U21318 (N_21318,N_14990,N_17480);
nor U21319 (N_21319,N_17417,N_12535);
nand U21320 (N_21320,N_14854,N_17273);
nor U21321 (N_21321,N_13754,N_15544);
xor U21322 (N_21322,N_17669,N_13191);
nand U21323 (N_21323,N_12874,N_14026);
and U21324 (N_21324,N_18573,N_12608);
nor U21325 (N_21325,N_16835,N_17781);
and U21326 (N_21326,N_14072,N_16236);
and U21327 (N_21327,N_17490,N_16655);
xnor U21328 (N_21328,N_14497,N_16316);
nor U21329 (N_21329,N_16217,N_15377);
xor U21330 (N_21330,N_14528,N_13463);
nand U21331 (N_21331,N_18170,N_18060);
nand U21332 (N_21332,N_14320,N_14551);
or U21333 (N_21333,N_16586,N_18668);
and U21334 (N_21334,N_14074,N_15363);
nand U21335 (N_21335,N_14565,N_13775);
nor U21336 (N_21336,N_15281,N_15038);
xnor U21337 (N_21337,N_14597,N_16743);
nand U21338 (N_21338,N_14495,N_17055);
or U21339 (N_21339,N_14690,N_16998);
or U21340 (N_21340,N_17362,N_18433);
and U21341 (N_21341,N_18056,N_17338);
nor U21342 (N_21342,N_15177,N_12562);
xor U21343 (N_21343,N_12963,N_15872);
nor U21344 (N_21344,N_12583,N_16167);
nor U21345 (N_21345,N_16021,N_18611);
xor U21346 (N_21346,N_17699,N_14151);
and U21347 (N_21347,N_13467,N_12993);
xor U21348 (N_21348,N_13788,N_18582);
nand U21349 (N_21349,N_16812,N_15613);
xnor U21350 (N_21350,N_13599,N_16599);
xor U21351 (N_21351,N_17992,N_15218);
or U21352 (N_21352,N_14504,N_16954);
and U21353 (N_21353,N_17149,N_16833);
nor U21354 (N_21354,N_17222,N_13947);
nand U21355 (N_21355,N_12613,N_14397);
nand U21356 (N_21356,N_15985,N_13108);
or U21357 (N_21357,N_13975,N_15144);
nor U21358 (N_21358,N_17377,N_18615);
nor U21359 (N_21359,N_16950,N_15672);
and U21360 (N_21360,N_15149,N_18326);
nor U21361 (N_21361,N_14787,N_13728);
and U21362 (N_21362,N_18413,N_14616);
and U21363 (N_21363,N_14587,N_14469);
nand U21364 (N_21364,N_14921,N_13102);
nor U21365 (N_21365,N_14934,N_13448);
nand U21366 (N_21366,N_18252,N_13733);
or U21367 (N_21367,N_16188,N_16184);
and U21368 (N_21368,N_13041,N_14654);
and U21369 (N_21369,N_13185,N_14761);
and U21370 (N_21370,N_18051,N_15397);
nand U21371 (N_21371,N_15588,N_17203);
and U21372 (N_21372,N_16945,N_16356);
and U21373 (N_21373,N_17688,N_15846);
nand U21374 (N_21374,N_15385,N_14626);
and U21375 (N_21375,N_12655,N_12940);
xnor U21376 (N_21376,N_16205,N_15820);
and U21377 (N_21377,N_13558,N_12898);
or U21378 (N_21378,N_13095,N_15806);
nor U21379 (N_21379,N_16871,N_17204);
xnor U21380 (N_21380,N_15697,N_12674);
and U21381 (N_21381,N_15403,N_16556);
or U21382 (N_21382,N_14089,N_18023);
nor U21383 (N_21383,N_15473,N_15095);
and U21384 (N_21384,N_15877,N_13504);
and U21385 (N_21385,N_18666,N_17186);
nor U21386 (N_21386,N_14272,N_16899);
nor U21387 (N_21387,N_13676,N_12651);
nand U21388 (N_21388,N_13270,N_18322);
xnor U21389 (N_21389,N_16095,N_13651);
nor U21390 (N_21390,N_17043,N_14048);
xnor U21391 (N_21391,N_16854,N_12975);
or U21392 (N_21392,N_14510,N_18350);
or U21393 (N_21393,N_18423,N_17997);
nand U21394 (N_21394,N_15612,N_14249);
xor U21395 (N_21395,N_15065,N_12783);
or U21396 (N_21396,N_16134,N_15638);
and U21397 (N_21397,N_17926,N_18720);
and U21398 (N_21398,N_18722,N_13878);
xnor U21399 (N_21399,N_12976,N_16974);
or U21400 (N_21400,N_17384,N_15682);
and U21401 (N_21401,N_17134,N_16451);
and U21402 (N_21402,N_18081,N_15658);
xnor U21403 (N_21403,N_17904,N_14794);
xnor U21404 (N_21404,N_15916,N_14590);
xor U21405 (N_21405,N_15454,N_13165);
or U21406 (N_21406,N_13221,N_16746);
nand U21407 (N_21407,N_13076,N_16049);
nor U21408 (N_21408,N_16673,N_13135);
and U21409 (N_21409,N_14685,N_17678);
xnor U21410 (N_21410,N_17549,N_16083);
or U21411 (N_21411,N_12950,N_16053);
or U21412 (N_21412,N_16151,N_16388);
xnor U21413 (N_21413,N_14888,N_16660);
and U21414 (N_21414,N_16014,N_14561);
xnor U21415 (N_21415,N_16787,N_18043);
or U21416 (N_21416,N_14206,N_14786);
nand U21417 (N_21417,N_14183,N_18323);
nor U21418 (N_21418,N_14028,N_12879);
nor U21419 (N_21419,N_16739,N_13525);
and U21420 (N_21420,N_18357,N_16104);
or U21421 (N_21421,N_15856,N_15903);
nor U21422 (N_21422,N_14463,N_13980);
and U21423 (N_21423,N_16218,N_18428);
xnor U21424 (N_21424,N_15547,N_15702);
nor U21425 (N_21425,N_16563,N_14092);
xnor U21426 (N_21426,N_17927,N_13207);
nand U21427 (N_21427,N_16628,N_14107);
nor U21428 (N_21428,N_16252,N_16019);
or U21429 (N_21429,N_14800,N_14848);
nor U21430 (N_21430,N_16310,N_17141);
and U21431 (N_21431,N_13920,N_15392);
nor U21432 (N_21432,N_18549,N_17907);
or U21433 (N_21433,N_17525,N_16676);
or U21434 (N_21434,N_18161,N_15559);
nor U21435 (N_21435,N_13641,N_12579);
and U21436 (N_21436,N_14688,N_12873);
or U21437 (N_21437,N_12981,N_18443);
or U21438 (N_21438,N_15936,N_16934);
xnor U21439 (N_21439,N_13113,N_18399);
xnor U21440 (N_21440,N_12682,N_17816);
xnor U21441 (N_21441,N_14925,N_13354);
or U21442 (N_21442,N_18059,N_16879);
nand U21443 (N_21443,N_16576,N_15302);
nand U21444 (N_21444,N_13767,N_16168);
nand U21445 (N_21445,N_13561,N_16116);
and U21446 (N_21446,N_14884,N_15024);
or U21447 (N_21447,N_14535,N_18464);
or U21448 (N_21448,N_12910,N_15853);
nand U21449 (N_21449,N_17990,N_18672);
or U21450 (N_21450,N_14409,N_18110);
and U21451 (N_21451,N_18245,N_17428);
and U21452 (N_21452,N_12756,N_18041);
or U21453 (N_21453,N_18592,N_17103);
and U21454 (N_21454,N_16226,N_17349);
or U21455 (N_21455,N_17940,N_13797);
nor U21456 (N_21456,N_14877,N_16666);
and U21457 (N_21457,N_17014,N_16784);
or U21458 (N_21458,N_17854,N_14326);
xor U21459 (N_21459,N_16058,N_14618);
nand U21460 (N_21460,N_17144,N_15665);
nor U21461 (N_21461,N_18078,N_16550);
nor U21462 (N_21462,N_14780,N_13411);
and U21463 (N_21463,N_16869,N_18468);
or U21464 (N_21464,N_13083,N_17547);
or U21465 (N_21465,N_17611,N_15531);
nor U21466 (N_21466,N_17588,N_14906);
nor U21467 (N_21467,N_14950,N_13881);
nand U21468 (N_21468,N_13603,N_16398);
or U21469 (N_21469,N_14115,N_17581);
nor U21470 (N_21470,N_12680,N_15088);
and U21471 (N_21471,N_14166,N_17213);
nor U21472 (N_21472,N_16414,N_15339);
nand U21473 (N_21473,N_13683,N_17482);
xor U21474 (N_21474,N_18619,N_13715);
or U21475 (N_21475,N_16107,N_13517);
or U21476 (N_21476,N_16652,N_17294);
or U21477 (N_21477,N_16204,N_15169);
or U21478 (N_21478,N_18025,N_15030);
nor U21479 (N_21479,N_15769,N_17636);
and U21480 (N_21480,N_14351,N_17143);
nor U21481 (N_21481,N_13120,N_14665);
nor U21482 (N_21482,N_14662,N_12594);
nor U21483 (N_21483,N_18457,N_18109);
xnor U21484 (N_21484,N_17556,N_12681);
and U21485 (N_21485,N_16770,N_15278);
nand U21486 (N_21486,N_15107,N_13211);
nor U21487 (N_21487,N_15325,N_17129);
or U21488 (N_21488,N_17147,N_16222);
xor U21489 (N_21489,N_15215,N_16460);
and U21490 (N_21490,N_15360,N_17289);
nand U21491 (N_21491,N_14069,N_15016);
and U21492 (N_21492,N_18136,N_18697);
or U21493 (N_21493,N_18388,N_15781);
or U21494 (N_21494,N_13443,N_17594);
xor U21495 (N_21495,N_12932,N_16641);
nor U21496 (N_21496,N_17829,N_13110);
or U21497 (N_21497,N_12915,N_17309);
and U21498 (N_21498,N_18270,N_17329);
nand U21499 (N_21499,N_14514,N_15081);
nor U21500 (N_21500,N_16696,N_17524);
or U21501 (N_21501,N_14268,N_13417);
xnor U21502 (N_21502,N_17879,N_18631);
xor U21503 (N_21503,N_17744,N_13746);
and U21504 (N_21504,N_13160,N_16855);
and U21505 (N_21505,N_17770,N_15529);
and U21506 (N_21506,N_14698,N_18518);
or U21507 (N_21507,N_15444,N_17771);
nor U21508 (N_21508,N_14481,N_14011);
xnor U21509 (N_21509,N_17736,N_18050);
xor U21510 (N_21510,N_13396,N_18181);
nand U21511 (N_21511,N_14831,N_17402);
nor U21512 (N_21512,N_13837,N_17288);
nor U21513 (N_21513,N_14634,N_14608);
nand U21514 (N_21514,N_15606,N_18450);
xnor U21515 (N_21515,N_13431,N_16264);
xor U21516 (N_21516,N_16387,N_15047);
or U21517 (N_21517,N_14157,N_13929);
nand U21518 (N_21518,N_17076,N_13501);
and U21519 (N_21519,N_16197,N_16803);
xor U21520 (N_21520,N_16892,N_16904);
xnor U21521 (N_21521,N_17557,N_13615);
or U21522 (N_21522,N_17370,N_12518);
or U21523 (N_21523,N_18585,N_18596);
nor U21524 (N_21524,N_18167,N_15464);
nand U21525 (N_21525,N_16600,N_18483);
xor U21526 (N_21526,N_15192,N_17473);
xnor U21527 (N_21527,N_16640,N_17631);
or U21528 (N_21528,N_16911,N_15597);
and U21529 (N_21529,N_13252,N_18430);
or U21530 (N_21530,N_15171,N_16800);
nor U21531 (N_21531,N_17335,N_13817);
nor U21532 (N_21532,N_15659,N_13204);
nand U21533 (N_21533,N_14902,N_16358);
nand U21534 (N_21534,N_17882,N_17731);
nand U21535 (N_21535,N_12720,N_13963);
and U21536 (N_21536,N_14960,N_14068);
xor U21537 (N_21537,N_13350,N_15577);
or U21538 (N_21538,N_13306,N_13882);
nor U21539 (N_21539,N_15889,N_15782);
and U21540 (N_21540,N_18377,N_14838);
and U21541 (N_21541,N_14356,N_12638);
xnor U21542 (N_21542,N_14499,N_18567);
xnor U21543 (N_21543,N_17725,N_17183);
or U21544 (N_21544,N_14125,N_12920);
nand U21545 (N_21545,N_12902,N_15451);
nor U21546 (N_21546,N_16022,N_15276);
or U21547 (N_21547,N_17308,N_17715);
nor U21548 (N_21548,N_17453,N_18555);
nor U21549 (N_21549,N_17559,N_15167);
and U21550 (N_21550,N_16991,N_17639);
nand U21551 (N_21551,N_17042,N_15405);
or U21552 (N_21552,N_14075,N_15469);
xor U21553 (N_21553,N_13260,N_14505);
nor U21554 (N_21554,N_15393,N_13276);
nor U21555 (N_21555,N_14679,N_17761);
or U21556 (N_21556,N_13665,N_15667);
or U21557 (N_21557,N_18477,N_16474);
xor U21558 (N_21558,N_14930,N_18543);
nand U21559 (N_21559,N_16233,N_15040);
nand U21560 (N_21560,N_16158,N_17262);
or U21561 (N_21561,N_15743,N_14432);
or U21562 (N_21562,N_17704,N_14194);
nor U21563 (N_21563,N_17645,N_17875);
and U21564 (N_21564,N_14999,N_16174);
nand U21565 (N_21565,N_13867,N_16568);
nand U21566 (N_21566,N_17010,N_17220);
xor U21567 (N_21567,N_12911,N_17169);
nor U21568 (N_21568,N_14207,N_15566);
and U21569 (N_21569,N_16718,N_13245);
nor U21570 (N_21570,N_13446,N_16313);
nand U21571 (N_21571,N_16594,N_15593);
or U21572 (N_21572,N_18733,N_16564);
or U21573 (N_21573,N_15410,N_14063);
and U21574 (N_21574,N_15270,N_14296);
xnor U21575 (N_21575,N_12675,N_14830);
or U21576 (N_21576,N_18590,N_15043);
or U21577 (N_21577,N_15143,N_17046);
nor U21578 (N_21578,N_16033,N_15190);
or U21579 (N_21579,N_14799,N_14553);
and U21580 (N_21580,N_15259,N_18623);
or U21581 (N_21581,N_15642,N_13989);
xor U21582 (N_21582,N_17661,N_13353);
xnor U21583 (N_21583,N_16438,N_14133);
xor U21584 (N_21584,N_14998,N_16885);
or U21585 (N_21585,N_17656,N_16216);
or U21586 (N_21586,N_13072,N_17963);
nor U21587 (N_21587,N_17008,N_17933);
nand U21588 (N_21588,N_15630,N_15022);
and U21589 (N_21589,N_16348,N_17434);
and U21590 (N_21590,N_18058,N_15619);
nand U21591 (N_21591,N_18128,N_17078);
nor U21592 (N_21592,N_17817,N_17950);
or U21593 (N_21593,N_15932,N_16615);
and U21594 (N_21594,N_12590,N_18325);
and U21595 (N_21595,N_15635,N_13158);
or U21596 (N_21596,N_16859,N_18620);
nor U21597 (N_21597,N_13605,N_15076);
xor U21598 (N_21598,N_18141,N_13528);
nand U21599 (N_21599,N_17537,N_12957);
nor U21600 (N_21600,N_17956,N_12585);
nor U21601 (N_21601,N_14751,N_17768);
and U21602 (N_21602,N_17696,N_18704);
or U21603 (N_21603,N_15569,N_13584);
and U21604 (N_21604,N_13952,N_14358);
nor U21605 (N_21605,N_15502,N_17182);
nand U21606 (N_21606,N_18677,N_16332);
nand U21607 (N_21607,N_13840,N_14676);
nand U21608 (N_21608,N_18222,N_17987);
or U21609 (N_21609,N_14454,N_18045);
nand U21610 (N_21610,N_13937,N_18708);
xnor U21611 (N_21611,N_15953,N_14712);
xor U21612 (N_21612,N_16283,N_15574);
or U21613 (N_21613,N_14870,N_15268);
nor U21614 (N_21614,N_14110,N_17161);
nand U21615 (N_21615,N_13283,N_18716);
and U21616 (N_21616,N_12988,N_12690);
nor U21617 (N_21617,N_16198,N_17437);
and U21618 (N_21618,N_13800,N_17999);
or U21619 (N_21619,N_18420,N_15327);
nor U21620 (N_21620,N_16372,N_13887);
and U21621 (N_21621,N_14349,N_15382);
nor U21622 (N_21622,N_16658,N_17188);
nor U21623 (N_21623,N_15533,N_14880);
nor U21624 (N_21624,N_12703,N_15139);
nor U21625 (N_21625,N_13376,N_18533);
and U21626 (N_21626,N_15900,N_16514);
xnor U21627 (N_21627,N_17732,N_12589);
or U21628 (N_21628,N_15708,N_14304);
or U21629 (N_21629,N_18329,N_15396);
xor U21630 (N_21630,N_12958,N_16453);
nor U21631 (N_21631,N_12994,N_17773);
or U21632 (N_21632,N_17233,N_15459);
xnor U21633 (N_21633,N_17860,N_16324);
xnor U21634 (N_21634,N_14897,N_17000);
nand U21635 (N_21635,N_18080,N_16808);
xor U21636 (N_21636,N_17979,N_17440);
and U21637 (N_21637,N_13107,N_16846);
and U21638 (N_21638,N_15350,N_18709);
and U21639 (N_21639,N_17886,N_15210);
or U21640 (N_21640,N_14363,N_14840);
xnor U21641 (N_21641,N_18455,N_14704);
xnor U21642 (N_21642,N_14033,N_16769);
and U21643 (N_21643,N_13763,N_15483);
or U21644 (N_21644,N_15645,N_18340);
nor U21645 (N_21645,N_13588,N_14873);
and U21646 (N_21646,N_15937,N_16365);
and U21647 (N_21647,N_13801,N_17670);
or U21648 (N_21648,N_15777,N_16581);
and U21649 (N_21649,N_13315,N_13112);
nand U21650 (N_21650,N_12843,N_14386);
and U21651 (N_21651,N_14101,N_13208);
xnor U21652 (N_21652,N_13359,N_17833);
nor U21653 (N_21653,N_15443,N_16826);
nand U21654 (N_21654,N_14563,N_13015);
or U21655 (N_21655,N_14824,N_16567);
xor U21656 (N_21656,N_14248,N_14754);
and U21657 (N_21657,N_13061,N_15629);
xnor U21658 (N_21658,N_17693,N_16792);
xor U21659 (N_21659,N_18729,N_17754);
xor U21660 (N_21660,N_12888,N_18160);
nor U21661 (N_21661,N_15907,N_13550);
nor U21662 (N_21662,N_17180,N_13441);
nand U21663 (N_21663,N_17404,N_14290);
or U21664 (N_21664,N_14277,N_14413);
xnor U21665 (N_21665,N_12520,N_13365);
and U21666 (N_21666,N_15147,N_15747);
nor U21667 (N_21667,N_18480,N_17938);
and U21668 (N_21668,N_13115,N_16115);
and U21669 (N_21669,N_16279,N_14878);
or U21670 (N_21670,N_16246,N_12838);
or U21671 (N_21671,N_15168,N_14275);
nand U21672 (N_21672,N_15795,N_15554);
or U21673 (N_21673,N_18162,N_15213);
nand U21674 (N_21674,N_14130,N_18375);
xor U21675 (N_21675,N_16249,N_14567);
nand U21676 (N_21676,N_14477,N_14589);
nor U21677 (N_21677,N_12952,N_12635);
xnor U21678 (N_21678,N_16522,N_13300);
or U21679 (N_21679,N_15912,N_15848);
nand U21680 (N_21680,N_13914,N_13345);
nor U21681 (N_21681,N_12923,N_17939);
and U21682 (N_21682,N_14987,N_17601);
xnor U21683 (N_21683,N_18461,N_14862);
or U21684 (N_21684,N_17459,N_18744);
nand U21685 (N_21685,N_14119,N_14460);
or U21686 (N_21686,N_17098,N_17466);
xnor U21687 (N_21687,N_18154,N_14736);
and U21688 (N_21688,N_16638,N_16117);
xnor U21689 (N_21689,N_15346,N_15978);
nand U21690 (N_21690,N_15591,N_15940);
and U21691 (N_21691,N_12529,N_14245);
xnor U21692 (N_21692,N_15532,N_14959);
or U21693 (N_21693,N_15020,N_17847);
nand U21694 (N_21694,N_16656,N_15947);
nor U21695 (N_21695,N_15519,N_17173);
xor U21696 (N_21696,N_12698,N_17807);
and U21697 (N_21697,N_18453,N_18410);
or U21698 (N_21698,N_14869,N_15340);
nand U21699 (N_21699,N_15892,N_13478);
and U21700 (N_21700,N_13370,N_13654);
and U21701 (N_21701,N_14506,N_15216);
or U21702 (N_21702,N_18482,N_17413);
or U21703 (N_21703,N_12715,N_14078);
xnor U21704 (N_21704,N_16646,N_17750);
xor U21705 (N_21705,N_16726,N_18046);
nand U21706 (N_21706,N_17075,N_14343);
or U21707 (N_21707,N_16631,N_17873);
nor U21708 (N_21708,N_18600,N_14017);
and U21709 (N_21709,N_18054,N_14954);
xnor U21710 (N_21710,N_12631,N_18009);
nor U21711 (N_21711,N_13044,N_12809);
or U21712 (N_21712,N_18083,N_15970);
xor U21713 (N_21713,N_15049,N_12542);
nor U21714 (N_21714,N_13518,N_13813);
or U21715 (N_21715,N_13297,N_17630);
and U21716 (N_21716,N_13729,N_16947);
and U21717 (N_21717,N_16256,N_15779);
or U21718 (N_21718,N_15201,N_15174);
or U21719 (N_21719,N_15084,N_18108);
nor U21720 (N_21720,N_17841,N_16030);
xor U21721 (N_21721,N_16412,N_17658);
nand U21722 (N_21722,N_12634,N_17248);
nand U21723 (N_21723,N_14303,N_16910);
xor U21724 (N_21724,N_17523,N_15730);
and U21725 (N_21725,N_16847,N_16837);
or U21726 (N_21726,N_13244,N_17360);
xor U21727 (N_21727,N_12732,N_14117);
or U21728 (N_21728,N_14242,N_17499);
nand U21729 (N_21729,N_16931,N_13841);
and U21730 (N_21730,N_16148,N_13750);
or U21731 (N_21731,N_13363,N_15298);
or U21732 (N_21732,N_18255,N_12524);
nor U21733 (N_21733,N_12643,N_16889);
and U21734 (N_21734,N_12521,N_18279);
nor U21735 (N_21735,N_14923,N_14913);
xnor U21736 (N_21736,N_14185,N_13037);
nor U21737 (N_21737,N_16347,N_13955);
nor U21738 (N_21738,N_14113,N_18642);
or U21739 (N_21739,N_17375,N_16503);
xor U21740 (N_21740,N_13062,N_16858);
and U21741 (N_21741,N_14974,N_13679);
xor U21742 (N_21742,N_14439,N_13111);
and U21743 (N_21743,N_15011,N_17202);
nand U21744 (N_21744,N_16008,N_15295);
nor U21745 (N_21745,N_14701,N_17366);
xor U21746 (N_21746,N_13793,N_12753);
nor U21747 (N_21747,N_12605,N_16043);
nor U21748 (N_21748,N_15476,N_16986);
or U21749 (N_21749,N_17481,N_18610);
xor U21750 (N_21750,N_17554,N_15376);
or U21751 (N_21751,N_17734,N_13026);
and U21752 (N_21752,N_15714,N_14500);
and U21753 (N_21753,N_15087,N_13199);
xor U21754 (N_21754,N_15826,N_14579);
or U21755 (N_21755,N_14517,N_14865);
xnor U21756 (N_21756,N_14768,N_12559);
nand U21757 (N_21757,N_13960,N_13876);
or U21758 (N_21758,N_14209,N_12747);
nor U21759 (N_21759,N_15236,N_17591);
nand U21760 (N_21760,N_17922,N_12913);
nand U21761 (N_21761,N_18295,N_15492);
xor U21762 (N_21762,N_16562,N_15164);
nand U21763 (N_21763,N_12533,N_15251);
nand U21764 (N_21764,N_18324,N_13461);
nor U21765 (N_21765,N_14021,N_13432);
or U21766 (N_21766,N_15408,N_17901);
nor U21767 (N_21767,N_13084,N_14633);
or U21768 (N_21768,N_17209,N_13513);
and U21769 (N_21769,N_15674,N_13369);
nor U21770 (N_21770,N_14806,N_13329);
and U21771 (N_21771,N_15818,N_14362);
xor U21772 (N_21772,N_15202,N_15914);
xor U21773 (N_21773,N_13138,N_14202);
and U21774 (N_21774,N_18254,N_13983);
and U21775 (N_21775,N_14670,N_17991);
or U21776 (N_21776,N_12778,N_14366);
or U21777 (N_21777,N_16027,N_16179);
nand U21778 (N_21778,N_17852,N_13125);
nor U21779 (N_21779,N_13181,N_12504);
or U21780 (N_21780,N_14719,N_15157);
and U21781 (N_21781,N_15014,N_18121);
xnor U21782 (N_21782,N_17961,N_18166);
or U21783 (N_21783,N_13748,N_14307);
nor U21784 (N_21784,N_18259,N_13524);
and U21785 (N_21785,N_14000,N_13073);
nor U21786 (N_21786,N_16481,N_13020);
nor U21787 (N_21787,N_12985,N_15891);
or U21788 (N_21788,N_13070,N_16057);
xnor U21789 (N_21789,N_14214,N_15158);
and U21790 (N_21790,N_16123,N_14350);
nand U21791 (N_21791,N_17430,N_17584);
or U21792 (N_21792,N_15938,N_17751);
nor U21793 (N_21793,N_14269,N_14939);
xor U21794 (N_21794,N_14542,N_18142);
nand U21795 (N_21795,N_13137,N_14749);
nand U21796 (N_21796,N_15621,N_13166);
nor U21797 (N_21797,N_17962,N_15136);
nand U21798 (N_21798,N_16268,N_17970);
xnor U21799 (N_21799,N_15313,N_14188);
or U21800 (N_21800,N_16992,N_18536);
or U21801 (N_21801,N_16298,N_13291);
nand U21802 (N_21802,N_16580,N_16143);
or U21803 (N_21803,N_12705,N_16925);
nand U21804 (N_21804,N_15484,N_18393);
xor U21805 (N_21805,N_17590,N_13536);
nand U21806 (N_21806,N_16099,N_13970);
nand U21807 (N_21807,N_16165,N_15490);
nand U21808 (N_21808,N_13774,N_16473);
nor U21809 (N_21809,N_15512,N_16775);
and U21810 (N_21810,N_15567,N_17625);
and U21811 (N_21811,N_18021,N_14367);
and U21812 (N_21812,N_15836,N_16618);
and U21813 (N_21813,N_14336,N_13424);
or U21814 (N_21814,N_14109,N_16257);
xor U21815 (N_21815,N_15557,N_13864);
or U21816 (N_21816,N_12934,N_16411);
or U21817 (N_21817,N_13620,N_14315);
or U21818 (N_21818,N_14681,N_17128);
or U21819 (N_21819,N_12522,N_13215);
xor U21820 (N_21820,N_12820,N_12807);
xnor U21821 (N_21821,N_16349,N_18353);
nor U21822 (N_21822,N_12556,N_18603);
nand U21823 (N_21823,N_17167,N_17945);
and U21824 (N_21824,N_16023,N_16862);
xor U21825 (N_21825,N_15480,N_13535);
nand U21826 (N_21826,N_13145,N_16525);
nand U21827 (N_21827,N_14599,N_16292);
nor U21828 (N_21828,N_17850,N_18290);
xor U21829 (N_21829,N_13521,N_13094);
or U21830 (N_21830,N_17373,N_14444);
and U21831 (N_21831,N_13761,N_16665);
xor U21832 (N_21832,N_14876,N_17177);
and U21833 (N_21833,N_14692,N_12777);
nand U21834 (N_21834,N_14828,N_18728);
or U21835 (N_21835,N_12771,N_15112);
xnor U21836 (N_21836,N_15549,N_13758);
and U21837 (N_21837,N_15130,N_13846);
nor U21838 (N_21838,N_17802,N_14250);
xor U21839 (N_21839,N_18299,N_16329);
or U21840 (N_21840,N_16267,N_14964);
nor U21841 (N_21841,N_15058,N_17651);
and U21842 (N_21842,N_17667,N_13187);
nor U21843 (N_21843,N_15261,N_14746);
nor U21844 (N_21844,N_13071,N_14003);
or U21845 (N_21845,N_18207,N_12568);
nor U21846 (N_21846,N_12885,N_15649);
xor U21847 (N_21847,N_18089,N_15744);
nor U21848 (N_21848,N_17163,N_12933);
xor U21849 (N_21849,N_17748,N_16135);
xor U21850 (N_21850,N_16375,N_16795);
and U21851 (N_21851,N_18445,N_18268);
nand U21852 (N_21852,N_16044,N_13298);
or U21853 (N_21853,N_13100,N_13119);
nor U21854 (N_21854,N_16110,N_13492);
nand U21855 (N_21855,N_13909,N_18088);
nor U21856 (N_21856,N_16850,N_15271);
nand U21857 (N_21857,N_14233,N_18282);
nand U21858 (N_21858,N_12846,N_15487);
and U21859 (N_21859,N_17155,N_15546);
and U21860 (N_21860,N_16953,N_17548);
and U21861 (N_21861,N_12882,N_15436);
nor U21862 (N_21862,N_17433,N_16063);
nor U21863 (N_21863,N_14474,N_16756);
nor U21864 (N_21864,N_13827,N_17993);
nand U21865 (N_21865,N_17056,N_13856);
xnor U21866 (N_21866,N_17283,N_16345);
or U21867 (N_21867,N_15054,N_14348);
nor U21868 (N_21868,N_16939,N_18429);
nand U21869 (N_21869,N_15328,N_13901);
and U21870 (N_21870,N_18289,N_15422);
nor U21871 (N_21871,N_15899,N_12856);
or U21872 (N_21872,N_18084,N_14094);
nand U21873 (N_21873,N_18182,N_15113);
nor U21874 (N_21874,N_14414,N_15545);
or U21875 (N_21875,N_17934,N_15989);
and U21876 (N_21876,N_14581,N_17541);
or U21877 (N_21877,N_13817,N_18033);
or U21878 (N_21878,N_17353,N_13199);
nor U21879 (N_21879,N_12706,N_15864);
xor U21880 (N_21880,N_14990,N_17930);
nand U21881 (N_21881,N_15945,N_17794);
or U21882 (N_21882,N_15822,N_16059);
xnor U21883 (N_21883,N_14917,N_14723);
nor U21884 (N_21884,N_14479,N_14209);
and U21885 (N_21885,N_15957,N_15730);
nand U21886 (N_21886,N_14695,N_17260);
xor U21887 (N_21887,N_17108,N_15290);
nor U21888 (N_21888,N_13909,N_13164);
xnor U21889 (N_21889,N_17981,N_13324);
xnor U21890 (N_21890,N_17255,N_17268);
nand U21891 (N_21891,N_14929,N_16177);
nor U21892 (N_21892,N_15944,N_12915);
or U21893 (N_21893,N_15642,N_16362);
and U21894 (N_21894,N_14039,N_14096);
nor U21895 (N_21895,N_17587,N_13247);
xnor U21896 (N_21896,N_12565,N_18124);
xor U21897 (N_21897,N_12621,N_12948);
or U21898 (N_21898,N_12764,N_15870);
or U21899 (N_21899,N_15760,N_12893);
and U21900 (N_21900,N_12954,N_16815);
nor U21901 (N_21901,N_13405,N_18516);
or U21902 (N_21902,N_16064,N_18460);
xnor U21903 (N_21903,N_14150,N_13979);
xnor U21904 (N_21904,N_18021,N_13207);
and U21905 (N_21905,N_13226,N_16195);
xor U21906 (N_21906,N_14683,N_14343);
or U21907 (N_21907,N_13167,N_14626);
xor U21908 (N_21908,N_14348,N_16688);
xor U21909 (N_21909,N_18375,N_13053);
or U21910 (N_21910,N_17437,N_13080);
and U21911 (N_21911,N_16367,N_12654);
and U21912 (N_21912,N_13082,N_17955);
or U21913 (N_21913,N_15934,N_15744);
and U21914 (N_21914,N_17858,N_16817);
xnor U21915 (N_21915,N_12997,N_16994);
nor U21916 (N_21916,N_13453,N_12532);
and U21917 (N_21917,N_15891,N_13589);
or U21918 (N_21918,N_13658,N_16801);
or U21919 (N_21919,N_17476,N_13377);
and U21920 (N_21920,N_14867,N_16355);
and U21921 (N_21921,N_17058,N_18494);
xor U21922 (N_21922,N_13664,N_12886);
nor U21923 (N_21923,N_16479,N_18431);
xnor U21924 (N_21924,N_13854,N_18267);
nand U21925 (N_21925,N_16469,N_15300);
nand U21926 (N_21926,N_15632,N_15057);
xor U21927 (N_21927,N_16820,N_13859);
and U21928 (N_21928,N_13655,N_15801);
nor U21929 (N_21929,N_14893,N_18645);
and U21930 (N_21930,N_13115,N_15695);
xnor U21931 (N_21931,N_14152,N_18670);
nor U21932 (N_21932,N_15161,N_17423);
and U21933 (N_21933,N_17618,N_18080);
and U21934 (N_21934,N_18228,N_17148);
or U21935 (N_21935,N_18026,N_12502);
and U21936 (N_21936,N_15039,N_12718);
xnor U21937 (N_21937,N_16694,N_16621);
or U21938 (N_21938,N_15944,N_14079);
or U21939 (N_21939,N_14188,N_16164);
or U21940 (N_21940,N_12613,N_13547);
or U21941 (N_21941,N_16396,N_14116);
and U21942 (N_21942,N_18649,N_13746);
and U21943 (N_21943,N_16368,N_13892);
nand U21944 (N_21944,N_17521,N_15909);
and U21945 (N_21945,N_15366,N_15857);
nor U21946 (N_21946,N_18404,N_16629);
nor U21947 (N_21947,N_18540,N_15975);
and U21948 (N_21948,N_12508,N_13587);
or U21949 (N_21949,N_14471,N_16676);
nand U21950 (N_21950,N_15900,N_13045);
nand U21951 (N_21951,N_16448,N_12880);
xor U21952 (N_21952,N_18062,N_16204);
nor U21953 (N_21953,N_14909,N_16607);
xnor U21954 (N_21954,N_15574,N_12583);
xor U21955 (N_21955,N_18688,N_15730);
nand U21956 (N_21956,N_14223,N_18313);
or U21957 (N_21957,N_13798,N_16692);
or U21958 (N_21958,N_17679,N_18657);
xnor U21959 (N_21959,N_14175,N_16819);
xnor U21960 (N_21960,N_12564,N_13221);
and U21961 (N_21961,N_14613,N_14608);
or U21962 (N_21962,N_14189,N_16054);
and U21963 (N_21963,N_13665,N_17329);
and U21964 (N_21964,N_14652,N_12759);
nand U21965 (N_21965,N_18708,N_16277);
or U21966 (N_21966,N_16353,N_17045);
or U21967 (N_21967,N_17632,N_16831);
nor U21968 (N_21968,N_13450,N_14528);
and U21969 (N_21969,N_15589,N_14104);
nor U21970 (N_21970,N_12841,N_15368);
xor U21971 (N_21971,N_17363,N_13110);
xnor U21972 (N_21972,N_16534,N_12634);
xor U21973 (N_21973,N_13460,N_13905);
or U21974 (N_21974,N_18003,N_18043);
or U21975 (N_21975,N_18573,N_12880);
xnor U21976 (N_21976,N_14908,N_15027);
nand U21977 (N_21977,N_15532,N_18015);
and U21978 (N_21978,N_15118,N_17329);
nand U21979 (N_21979,N_18038,N_12956);
nor U21980 (N_21980,N_12638,N_13851);
nand U21981 (N_21981,N_14143,N_16476);
xor U21982 (N_21982,N_13295,N_14232);
or U21983 (N_21983,N_15436,N_14351);
and U21984 (N_21984,N_17801,N_12983);
or U21985 (N_21985,N_18269,N_15995);
nand U21986 (N_21986,N_18686,N_12792);
or U21987 (N_21987,N_17810,N_16499);
xnor U21988 (N_21988,N_13865,N_16616);
nand U21989 (N_21989,N_13959,N_15410);
nand U21990 (N_21990,N_14538,N_14894);
nand U21991 (N_21991,N_15071,N_14250);
xnor U21992 (N_21992,N_17667,N_13777);
nand U21993 (N_21993,N_18665,N_13657);
or U21994 (N_21994,N_16622,N_14729);
nand U21995 (N_21995,N_13105,N_14934);
nor U21996 (N_21996,N_17612,N_13962);
or U21997 (N_21997,N_16987,N_13044);
or U21998 (N_21998,N_17417,N_12549);
nand U21999 (N_21999,N_12755,N_17981);
and U22000 (N_22000,N_16967,N_12901);
xnor U22001 (N_22001,N_17169,N_14346);
or U22002 (N_22002,N_14072,N_13136);
nand U22003 (N_22003,N_15085,N_18310);
and U22004 (N_22004,N_15239,N_15667);
nand U22005 (N_22005,N_13597,N_18352);
nor U22006 (N_22006,N_16468,N_13832);
and U22007 (N_22007,N_18284,N_18330);
or U22008 (N_22008,N_15064,N_16600);
or U22009 (N_22009,N_15156,N_12525);
or U22010 (N_22010,N_13391,N_14508);
or U22011 (N_22011,N_13719,N_16444);
and U22012 (N_22012,N_18344,N_15418);
nor U22013 (N_22013,N_14940,N_13423);
and U22014 (N_22014,N_15260,N_14703);
or U22015 (N_22015,N_14242,N_15003);
nor U22016 (N_22016,N_14583,N_14007);
and U22017 (N_22017,N_15469,N_18055);
and U22018 (N_22018,N_12720,N_13994);
or U22019 (N_22019,N_12769,N_14262);
nand U22020 (N_22020,N_13156,N_15372);
and U22021 (N_22021,N_18260,N_16150);
or U22022 (N_22022,N_13677,N_18316);
and U22023 (N_22023,N_12832,N_14717);
xor U22024 (N_22024,N_15807,N_14397);
xnor U22025 (N_22025,N_12508,N_17338);
and U22026 (N_22026,N_16474,N_17569);
and U22027 (N_22027,N_13255,N_18128);
xnor U22028 (N_22028,N_14603,N_18011);
xnor U22029 (N_22029,N_16051,N_16999);
nand U22030 (N_22030,N_14339,N_15109);
or U22031 (N_22031,N_14125,N_17257);
nand U22032 (N_22032,N_18705,N_17874);
xnor U22033 (N_22033,N_17660,N_14624);
and U22034 (N_22034,N_14391,N_16732);
and U22035 (N_22035,N_14473,N_16284);
nor U22036 (N_22036,N_15528,N_17002);
nand U22037 (N_22037,N_15964,N_13026);
xor U22038 (N_22038,N_14508,N_12602);
and U22039 (N_22039,N_17239,N_14850);
nand U22040 (N_22040,N_12576,N_18002);
and U22041 (N_22041,N_14717,N_12794);
nand U22042 (N_22042,N_13261,N_13445);
xnor U22043 (N_22043,N_15489,N_17033);
nor U22044 (N_22044,N_17401,N_14063);
and U22045 (N_22045,N_13320,N_12686);
nand U22046 (N_22046,N_17393,N_16974);
and U22047 (N_22047,N_16123,N_15391);
nor U22048 (N_22048,N_14661,N_15801);
xor U22049 (N_22049,N_14589,N_13687);
and U22050 (N_22050,N_13263,N_16854);
nor U22051 (N_22051,N_14465,N_18497);
xnor U22052 (N_22052,N_13379,N_14964);
or U22053 (N_22053,N_18671,N_15051);
xnor U22054 (N_22054,N_14921,N_18021);
nand U22055 (N_22055,N_18398,N_13390);
nor U22056 (N_22056,N_18264,N_16266);
and U22057 (N_22057,N_14377,N_14072);
nor U22058 (N_22058,N_12979,N_18128);
nor U22059 (N_22059,N_12769,N_13329);
xnor U22060 (N_22060,N_14194,N_18199);
and U22061 (N_22061,N_15137,N_15343);
and U22062 (N_22062,N_15676,N_14602);
xor U22063 (N_22063,N_18214,N_16836);
nor U22064 (N_22064,N_12533,N_15815);
nand U22065 (N_22065,N_12993,N_13573);
xor U22066 (N_22066,N_14974,N_13847);
or U22067 (N_22067,N_15993,N_14359);
nand U22068 (N_22068,N_16218,N_14334);
nor U22069 (N_22069,N_13853,N_13694);
nor U22070 (N_22070,N_16081,N_18566);
nor U22071 (N_22071,N_17064,N_15978);
nor U22072 (N_22072,N_17795,N_12568);
nand U22073 (N_22073,N_17816,N_15969);
or U22074 (N_22074,N_18314,N_14675);
xor U22075 (N_22075,N_16869,N_12654);
or U22076 (N_22076,N_14290,N_17377);
nor U22077 (N_22077,N_13293,N_12531);
or U22078 (N_22078,N_17627,N_16047);
or U22079 (N_22079,N_14121,N_14768);
or U22080 (N_22080,N_18425,N_16701);
nand U22081 (N_22081,N_14801,N_16661);
nand U22082 (N_22082,N_17764,N_13625);
or U22083 (N_22083,N_14477,N_13632);
nand U22084 (N_22084,N_13851,N_15875);
or U22085 (N_22085,N_16980,N_13699);
nand U22086 (N_22086,N_12932,N_15530);
and U22087 (N_22087,N_15299,N_17519);
or U22088 (N_22088,N_17270,N_18352);
nand U22089 (N_22089,N_13325,N_15808);
xnor U22090 (N_22090,N_13886,N_17234);
or U22091 (N_22091,N_18050,N_12509);
nand U22092 (N_22092,N_12731,N_14320);
nand U22093 (N_22093,N_18240,N_16323);
nand U22094 (N_22094,N_16689,N_14014);
and U22095 (N_22095,N_16245,N_12626);
nor U22096 (N_22096,N_14164,N_12863);
xor U22097 (N_22097,N_12844,N_15106);
or U22098 (N_22098,N_17435,N_14973);
and U22099 (N_22099,N_16110,N_14410);
or U22100 (N_22100,N_16174,N_16389);
and U22101 (N_22101,N_18624,N_15923);
nor U22102 (N_22102,N_17077,N_18272);
nor U22103 (N_22103,N_14719,N_17625);
and U22104 (N_22104,N_13988,N_16513);
and U22105 (N_22105,N_16851,N_15406);
or U22106 (N_22106,N_12655,N_14746);
nor U22107 (N_22107,N_12885,N_15662);
nand U22108 (N_22108,N_17352,N_15132);
and U22109 (N_22109,N_15006,N_13085);
and U22110 (N_22110,N_14899,N_15750);
nor U22111 (N_22111,N_18241,N_14854);
nand U22112 (N_22112,N_14829,N_14414);
nand U22113 (N_22113,N_17302,N_14921);
or U22114 (N_22114,N_12809,N_16659);
and U22115 (N_22115,N_13974,N_17802);
or U22116 (N_22116,N_17080,N_14148);
nor U22117 (N_22117,N_18063,N_15984);
or U22118 (N_22118,N_12623,N_12954);
xor U22119 (N_22119,N_13484,N_18359);
nand U22120 (N_22120,N_14317,N_15417);
nor U22121 (N_22121,N_17302,N_12778);
nor U22122 (N_22122,N_18018,N_17028);
or U22123 (N_22123,N_15362,N_13808);
or U22124 (N_22124,N_13405,N_14098);
nor U22125 (N_22125,N_14543,N_17094);
nand U22126 (N_22126,N_12763,N_16560);
nor U22127 (N_22127,N_16983,N_16324);
xor U22128 (N_22128,N_18745,N_16737);
or U22129 (N_22129,N_16022,N_15974);
nor U22130 (N_22130,N_15957,N_17016);
or U22131 (N_22131,N_12884,N_15291);
nand U22132 (N_22132,N_14242,N_13559);
xnor U22133 (N_22133,N_13544,N_15846);
nand U22134 (N_22134,N_16202,N_16554);
xor U22135 (N_22135,N_17779,N_13090);
xnor U22136 (N_22136,N_15979,N_13768);
xor U22137 (N_22137,N_17736,N_17924);
nand U22138 (N_22138,N_13173,N_12910);
and U22139 (N_22139,N_12778,N_13677);
and U22140 (N_22140,N_13406,N_16957);
and U22141 (N_22141,N_16931,N_13322);
xnor U22142 (N_22142,N_14105,N_17956);
and U22143 (N_22143,N_15544,N_12783);
and U22144 (N_22144,N_14600,N_17816);
xnor U22145 (N_22145,N_14553,N_12813);
xor U22146 (N_22146,N_16018,N_14874);
nand U22147 (N_22147,N_18468,N_16392);
or U22148 (N_22148,N_15966,N_15841);
nor U22149 (N_22149,N_14952,N_17463);
xnor U22150 (N_22150,N_16324,N_16878);
xnor U22151 (N_22151,N_13924,N_15530);
and U22152 (N_22152,N_18442,N_14378);
or U22153 (N_22153,N_16748,N_17245);
and U22154 (N_22154,N_15191,N_16431);
and U22155 (N_22155,N_18612,N_15114);
nand U22156 (N_22156,N_12827,N_14348);
xnor U22157 (N_22157,N_13837,N_17415);
nor U22158 (N_22158,N_13378,N_17428);
and U22159 (N_22159,N_16055,N_13216);
and U22160 (N_22160,N_15948,N_17265);
nand U22161 (N_22161,N_16226,N_17979);
and U22162 (N_22162,N_17603,N_12597);
and U22163 (N_22163,N_15083,N_13116);
xnor U22164 (N_22164,N_17650,N_14873);
nand U22165 (N_22165,N_12646,N_14471);
xnor U22166 (N_22166,N_15978,N_16765);
or U22167 (N_22167,N_14354,N_12686);
and U22168 (N_22168,N_12650,N_16737);
xnor U22169 (N_22169,N_17196,N_13233);
and U22170 (N_22170,N_17152,N_13272);
nor U22171 (N_22171,N_17273,N_17825);
xnor U22172 (N_22172,N_14289,N_16840);
nor U22173 (N_22173,N_17051,N_16242);
and U22174 (N_22174,N_13676,N_17605);
xor U22175 (N_22175,N_15000,N_12880);
and U22176 (N_22176,N_16010,N_18142);
nor U22177 (N_22177,N_14319,N_13712);
nor U22178 (N_22178,N_17540,N_18434);
or U22179 (N_22179,N_14502,N_14308);
xnor U22180 (N_22180,N_13336,N_13505);
xor U22181 (N_22181,N_13081,N_12956);
and U22182 (N_22182,N_16116,N_14466);
and U22183 (N_22183,N_12839,N_15070);
nand U22184 (N_22184,N_12739,N_14824);
and U22185 (N_22185,N_17756,N_12778);
or U22186 (N_22186,N_13618,N_18223);
or U22187 (N_22187,N_17947,N_16245);
or U22188 (N_22188,N_15502,N_18589);
or U22189 (N_22189,N_17122,N_15523);
xor U22190 (N_22190,N_16554,N_16056);
nor U22191 (N_22191,N_17022,N_13725);
or U22192 (N_22192,N_12913,N_18654);
or U22193 (N_22193,N_13202,N_16866);
nand U22194 (N_22194,N_13364,N_13610);
and U22195 (N_22195,N_15376,N_14533);
or U22196 (N_22196,N_18306,N_17202);
nor U22197 (N_22197,N_16496,N_13946);
nand U22198 (N_22198,N_17102,N_12892);
xnor U22199 (N_22199,N_13033,N_15425);
nor U22200 (N_22200,N_16660,N_14262);
xor U22201 (N_22201,N_12854,N_13763);
and U22202 (N_22202,N_13921,N_18286);
nor U22203 (N_22203,N_16631,N_15263);
nor U22204 (N_22204,N_17756,N_16233);
nand U22205 (N_22205,N_13159,N_15349);
nand U22206 (N_22206,N_15622,N_15215);
and U22207 (N_22207,N_15213,N_18749);
and U22208 (N_22208,N_13688,N_16633);
and U22209 (N_22209,N_14409,N_16150);
or U22210 (N_22210,N_13178,N_14818);
or U22211 (N_22211,N_12944,N_13593);
and U22212 (N_22212,N_16188,N_16067);
nor U22213 (N_22213,N_16593,N_17162);
xor U22214 (N_22214,N_15535,N_17077);
or U22215 (N_22215,N_15255,N_18701);
and U22216 (N_22216,N_16560,N_18440);
nand U22217 (N_22217,N_13611,N_14084);
xnor U22218 (N_22218,N_14259,N_16423);
and U22219 (N_22219,N_15778,N_15622);
xor U22220 (N_22220,N_15843,N_14778);
nor U22221 (N_22221,N_14278,N_17181);
and U22222 (N_22222,N_16993,N_16499);
and U22223 (N_22223,N_13314,N_14287);
and U22224 (N_22224,N_13455,N_17923);
or U22225 (N_22225,N_16477,N_16162);
nand U22226 (N_22226,N_16940,N_16382);
and U22227 (N_22227,N_14924,N_17285);
nor U22228 (N_22228,N_13258,N_18296);
nor U22229 (N_22229,N_15189,N_16025);
xor U22230 (N_22230,N_15485,N_13530);
nand U22231 (N_22231,N_16388,N_14541);
xor U22232 (N_22232,N_14141,N_14417);
nand U22233 (N_22233,N_15312,N_16940);
xor U22234 (N_22234,N_13722,N_13730);
nand U22235 (N_22235,N_17655,N_16111);
and U22236 (N_22236,N_13311,N_13667);
and U22237 (N_22237,N_15615,N_15767);
or U22238 (N_22238,N_14036,N_13416);
xor U22239 (N_22239,N_17814,N_16052);
and U22240 (N_22240,N_13605,N_18604);
xor U22241 (N_22241,N_16713,N_16339);
or U22242 (N_22242,N_14963,N_12859);
and U22243 (N_22243,N_14943,N_13152);
and U22244 (N_22244,N_15425,N_14243);
or U22245 (N_22245,N_14527,N_13197);
nor U22246 (N_22246,N_18584,N_14578);
or U22247 (N_22247,N_13357,N_14784);
or U22248 (N_22248,N_16906,N_13055);
or U22249 (N_22249,N_16314,N_13645);
xor U22250 (N_22250,N_13995,N_14916);
or U22251 (N_22251,N_17045,N_14924);
nand U22252 (N_22252,N_18189,N_15361);
nand U22253 (N_22253,N_13308,N_17094);
or U22254 (N_22254,N_17999,N_16065);
or U22255 (N_22255,N_16234,N_14125);
or U22256 (N_22256,N_15282,N_13240);
nor U22257 (N_22257,N_15745,N_14547);
xnor U22258 (N_22258,N_14748,N_18697);
xor U22259 (N_22259,N_18727,N_12654);
nand U22260 (N_22260,N_15718,N_14962);
nand U22261 (N_22261,N_17431,N_14021);
xor U22262 (N_22262,N_15244,N_12921);
or U22263 (N_22263,N_16782,N_18190);
and U22264 (N_22264,N_14958,N_15482);
or U22265 (N_22265,N_16514,N_16851);
and U22266 (N_22266,N_17839,N_12816);
xnor U22267 (N_22267,N_14922,N_17721);
or U22268 (N_22268,N_18348,N_13095);
xor U22269 (N_22269,N_15324,N_15368);
xor U22270 (N_22270,N_13556,N_15772);
xnor U22271 (N_22271,N_14765,N_13005);
xnor U22272 (N_22272,N_17931,N_16990);
nand U22273 (N_22273,N_15572,N_13591);
nor U22274 (N_22274,N_14741,N_14967);
or U22275 (N_22275,N_13612,N_15408);
xnor U22276 (N_22276,N_16753,N_12806);
and U22277 (N_22277,N_13973,N_15906);
and U22278 (N_22278,N_12970,N_16966);
or U22279 (N_22279,N_14805,N_17066);
nand U22280 (N_22280,N_13146,N_15906);
and U22281 (N_22281,N_17410,N_18513);
nor U22282 (N_22282,N_16983,N_14697);
nor U22283 (N_22283,N_16524,N_14585);
xnor U22284 (N_22284,N_17964,N_12529);
nor U22285 (N_22285,N_15280,N_16465);
nand U22286 (N_22286,N_12797,N_17328);
nand U22287 (N_22287,N_13617,N_18223);
nor U22288 (N_22288,N_13739,N_15336);
nor U22289 (N_22289,N_16357,N_16846);
xor U22290 (N_22290,N_12616,N_18298);
xnor U22291 (N_22291,N_18073,N_16874);
nor U22292 (N_22292,N_12622,N_14794);
xor U22293 (N_22293,N_15298,N_17898);
nand U22294 (N_22294,N_16106,N_17265);
nand U22295 (N_22295,N_15396,N_13299);
and U22296 (N_22296,N_16465,N_14400);
or U22297 (N_22297,N_17635,N_18245);
or U22298 (N_22298,N_17212,N_17609);
xor U22299 (N_22299,N_17879,N_18190);
and U22300 (N_22300,N_13658,N_14395);
or U22301 (N_22301,N_15618,N_16861);
xnor U22302 (N_22302,N_13993,N_15763);
nor U22303 (N_22303,N_13936,N_13167);
nor U22304 (N_22304,N_15649,N_15324);
and U22305 (N_22305,N_16922,N_18392);
or U22306 (N_22306,N_17940,N_15349);
nor U22307 (N_22307,N_12874,N_18366);
xor U22308 (N_22308,N_18264,N_13346);
nor U22309 (N_22309,N_15457,N_17794);
nor U22310 (N_22310,N_14374,N_16991);
xnor U22311 (N_22311,N_17191,N_15378);
xnor U22312 (N_22312,N_12836,N_15081);
and U22313 (N_22313,N_17245,N_18007);
and U22314 (N_22314,N_16079,N_17377);
or U22315 (N_22315,N_13735,N_16724);
nor U22316 (N_22316,N_17963,N_13070);
xor U22317 (N_22317,N_13862,N_17610);
nand U22318 (N_22318,N_13124,N_16619);
nand U22319 (N_22319,N_17277,N_18409);
xnor U22320 (N_22320,N_14101,N_14333);
xnor U22321 (N_22321,N_18334,N_14556);
xnor U22322 (N_22322,N_12745,N_14661);
nor U22323 (N_22323,N_12899,N_16656);
and U22324 (N_22324,N_18062,N_18161);
nor U22325 (N_22325,N_12640,N_18369);
nand U22326 (N_22326,N_16912,N_15251);
xnor U22327 (N_22327,N_12951,N_12549);
xnor U22328 (N_22328,N_17226,N_13600);
and U22329 (N_22329,N_12992,N_13340);
or U22330 (N_22330,N_12997,N_13101);
nor U22331 (N_22331,N_15008,N_13072);
and U22332 (N_22332,N_14842,N_13332);
or U22333 (N_22333,N_14537,N_13859);
and U22334 (N_22334,N_14189,N_14981);
and U22335 (N_22335,N_15280,N_15367);
or U22336 (N_22336,N_15880,N_17801);
and U22337 (N_22337,N_17906,N_16063);
and U22338 (N_22338,N_15610,N_13709);
xor U22339 (N_22339,N_13109,N_16744);
or U22340 (N_22340,N_12646,N_13771);
or U22341 (N_22341,N_18428,N_16897);
nand U22342 (N_22342,N_14074,N_13350);
xnor U22343 (N_22343,N_18524,N_13453);
nor U22344 (N_22344,N_14603,N_17196);
xnor U22345 (N_22345,N_15670,N_17786);
xor U22346 (N_22346,N_14911,N_16733);
or U22347 (N_22347,N_13626,N_12719);
and U22348 (N_22348,N_16779,N_16590);
nor U22349 (N_22349,N_18295,N_14584);
or U22350 (N_22350,N_18014,N_18076);
nand U22351 (N_22351,N_16516,N_14424);
nor U22352 (N_22352,N_14522,N_13451);
nand U22353 (N_22353,N_16250,N_16660);
nand U22354 (N_22354,N_14392,N_15766);
xor U22355 (N_22355,N_18112,N_17412);
nand U22356 (N_22356,N_15606,N_16412);
nor U22357 (N_22357,N_14502,N_17250);
xnor U22358 (N_22358,N_15083,N_15234);
nor U22359 (N_22359,N_13877,N_17206);
or U22360 (N_22360,N_17178,N_16624);
or U22361 (N_22361,N_17833,N_15460);
nor U22362 (N_22362,N_14133,N_12636);
nor U22363 (N_22363,N_14772,N_18173);
nor U22364 (N_22364,N_18590,N_17707);
nor U22365 (N_22365,N_13805,N_17827);
nand U22366 (N_22366,N_15702,N_17430);
xnor U22367 (N_22367,N_16643,N_13114);
nand U22368 (N_22368,N_14075,N_18334);
and U22369 (N_22369,N_16036,N_16802);
nand U22370 (N_22370,N_18592,N_16519);
xnor U22371 (N_22371,N_16621,N_16181);
xnor U22372 (N_22372,N_13870,N_13256);
xor U22373 (N_22373,N_14240,N_12587);
nor U22374 (N_22374,N_14550,N_17802);
and U22375 (N_22375,N_17620,N_17952);
and U22376 (N_22376,N_13908,N_15927);
xor U22377 (N_22377,N_13723,N_13668);
nand U22378 (N_22378,N_13875,N_15962);
or U22379 (N_22379,N_15207,N_12623);
nand U22380 (N_22380,N_13782,N_15412);
nor U22381 (N_22381,N_17999,N_18077);
nor U22382 (N_22382,N_14052,N_16147);
xor U22383 (N_22383,N_16254,N_15460);
nor U22384 (N_22384,N_14883,N_17863);
and U22385 (N_22385,N_17432,N_15573);
and U22386 (N_22386,N_15883,N_18087);
or U22387 (N_22387,N_14687,N_16368);
xnor U22388 (N_22388,N_18681,N_14296);
nand U22389 (N_22389,N_13004,N_16876);
nand U22390 (N_22390,N_15340,N_18700);
and U22391 (N_22391,N_18422,N_12514);
xor U22392 (N_22392,N_16405,N_15113);
nand U22393 (N_22393,N_14711,N_16080);
or U22394 (N_22394,N_16249,N_14919);
or U22395 (N_22395,N_16048,N_18338);
and U22396 (N_22396,N_13658,N_13194);
nor U22397 (N_22397,N_16337,N_14504);
and U22398 (N_22398,N_16984,N_17039);
nor U22399 (N_22399,N_17337,N_16782);
and U22400 (N_22400,N_17908,N_14588);
nand U22401 (N_22401,N_18255,N_17092);
xor U22402 (N_22402,N_13633,N_17842);
nor U22403 (N_22403,N_18675,N_16495);
or U22404 (N_22404,N_14415,N_13156);
xor U22405 (N_22405,N_17033,N_13897);
or U22406 (N_22406,N_13563,N_16572);
and U22407 (N_22407,N_13956,N_13735);
nor U22408 (N_22408,N_16609,N_18609);
or U22409 (N_22409,N_12836,N_18012);
or U22410 (N_22410,N_16708,N_17463);
nor U22411 (N_22411,N_18545,N_15338);
xnor U22412 (N_22412,N_16824,N_17619);
nor U22413 (N_22413,N_14468,N_17320);
or U22414 (N_22414,N_13878,N_18580);
and U22415 (N_22415,N_12887,N_18614);
and U22416 (N_22416,N_18434,N_15567);
xnor U22417 (N_22417,N_15592,N_14796);
nand U22418 (N_22418,N_12854,N_14606);
or U22419 (N_22419,N_12879,N_14096);
and U22420 (N_22420,N_17050,N_15083);
or U22421 (N_22421,N_13243,N_13828);
nor U22422 (N_22422,N_12513,N_14664);
or U22423 (N_22423,N_13360,N_18520);
xor U22424 (N_22424,N_16373,N_15656);
nor U22425 (N_22425,N_15613,N_12719);
or U22426 (N_22426,N_17834,N_15432);
or U22427 (N_22427,N_12593,N_13065);
xor U22428 (N_22428,N_17108,N_14905);
and U22429 (N_22429,N_13326,N_14079);
and U22430 (N_22430,N_15245,N_12972);
nor U22431 (N_22431,N_13146,N_14724);
or U22432 (N_22432,N_12974,N_14880);
and U22433 (N_22433,N_15209,N_13044);
or U22434 (N_22434,N_17376,N_16003);
and U22435 (N_22435,N_13084,N_17928);
xor U22436 (N_22436,N_18638,N_13117);
nand U22437 (N_22437,N_12658,N_16198);
xnor U22438 (N_22438,N_15040,N_15325);
xor U22439 (N_22439,N_12638,N_13712);
or U22440 (N_22440,N_17369,N_18071);
nand U22441 (N_22441,N_13296,N_14515);
nor U22442 (N_22442,N_15460,N_13056);
nor U22443 (N_22443,N_16034,N_17104);
or U22444 (N_22444,N_17419,N_18716);
and U22445 (N_22445,N_15135,N_17168);
nand U22446 (N_22446,N_13748,N_13457);
xor U22447 (N_22447,N_17610,N_15225);
or U22448 (N_22448,N_16024,N_17052);
and U22449 (N_22449,N_14262,N_17058);
nor U22450 (N_22450,N_17139,N_14554);
nor U22451 (N_22451,N_14078,N_18133);
nand U22452 (N_22452,N_14620,N_17780);
and U22453 (N_22453,N_17938,N_17565);
nand U22454 (N_22454,N_15281,N_12954);
nor U22455 (N_22455,N_12639,N_14087);
nand U22456 (N_22456,N_18237,N_13474);
or U22457 (N_22457,N_13670,N_15634);
and U22458 (N_22458,N_14619,N_12945);
and U22459 (N_22459,N_18098,N_12780);
xnor U22460 (N_22460,N_16775,N_12539);
nor U22461 (N_22461,N_12737,N_18130);
and U22462 (N_22462,N_15632,N_15769);
or U22463 (N_22463,N_17045,N_18166);
nand U22464 (N_22464,N_17719,N_18498);
or U22465 (N_22465,N_17710,N_12509);
and U22466 (N_22466,N_13213,N_16448);
or U22467 (N_22467,N_17313,N_14043);
and U22468 (N_22468,N_18201,N_15002);
xor U22469 (N_22469,N_13652,N_14746);
xor U22470 (N_22470,N_14161,N_16365);
or U22471 (N_22471,N_14925,N_15395);
nor U22472 (N_22472,N_17240,N_16960);
nand U22473 (N_22473,N_13079,N_13685);
xnor U22474 (N_22474,N_13491,N_15794);
or U22475 (N_22475,N_15082,N_16587);
nand U22476 (N_22476,N_13990,N_17064);
xnor U22477 (N_22477,N_16065,N_17606);
xnor U22478 (N_22478,N_13639,N_17020);
and U22479 (N_22479,N_17925,N_15191);
nor U22480 (N_22480,N_13389,N_17621);
and U22481 (N_22481,N_15998,N_15961);
nand U22482 (N_22482,N_18633,N_17656);
and U22483 (N_22483,N_17689,N_16276);
nor U22484 (N_22484,N_17572,N_14344);
xnor U22485 (N_22485,N_13574,N_14665);
nand U22486 (N_22486,N_16724,N_14362);
or U22487 (N_22487,N_14841,N_18653);
nor U22488 (N_22488,N_17285,N_18142);
nor U22489 (N_22489,N_17788,N_18609);
or U22490 (N_22490,N_14847,N_16626);
xnor U22491 (N_22491,N_14215,N_18720);
or U22492 (N_22492,N_13686,N_16636);
xnor U22493 (N_22493,N_15981,N_17698);
or U22494 (N_22494,N_12634,N_13138);
and U22495 (N_22495,N_17946,N_14533);
nand U22496 (N_22496,N_16883,N_16334);
and U22497 (N_22497,N_12615,N_14572);
and U22498 (N_22498,N_13818,N_17726);
xnor U22499 (N_22499,N_14546,N_13371);
xor U22500 (N_22500,N_12548,N_13335);
xor U22501 (N_22501,N_15834,N_15355);
or U22502 (N_22502,N_18635,N_12763);
nand U22503 (N_22503,N_13125,N_18200);
or U22504 (N_22504,N_13926,N_13525);
nand U22505 (N_22505,N_17297,N_12529);
and U22506 (N_22506,N_16132,N_16331);
nor U22507 (N_22507,N_13539,N_15242);
nor U22508 (N_22508,N_12848,N_17907);
and U22509 (N_22509,N_15572,N_17903);
xnor U22510 (N_22510,N_14675,N_17148);
nor U22511 (N_22511,N_15649,N_18256);
xor U22512 (N_22512,N_14694,N_15093);
nand U22513 (N_22513,N_16301,N_16431);
nor U22514 (N_22514,N_16945,N_13340);
or U22515 (N_22515,N_16534,N_18479);
xnor U22516 (N_22516,N_18275,N_17186);
or U22517 (N_22517,N_15356,N_13120);
nor U22518 (N_22518,N_15050,N_15306);
nor U22519 (N_22519,N_18479,N_15560);
or U22520 (N_22520,N_16677,N_16805);
nand U22521 (N_22521,N_16481,N_14627);
xnor U22522 (N_22522,N_17918,N_17942);
and U22523 (N_22523,N_17663,N_14164);
nand U22524 (N_22524,N_15433,N_17351);
nor U22525 (N_22525,N_15058,N_16924);
and U22526 (N_22526,N_17734,N_13163);
and U22527 (N_22527,N_16383,N_13747);
nor U22528 (N_22528,N_16373,N_12645);
nor U22529 (N_22529,N_18560,N_16865);
or U22530 (N_22530,N_16962,N_16112);
or U22531 (N_22531,N_12503,N_14721);
nand U22532 (N_22532,N_13815,N_18744);
nand U22533 (N_22533,N_17741,N_16112);
or U22534 (N_22534,N_13646,N_18677);
or U22535 (N_22535,N_17187,N_15994);
nand U22536 (N_22536,N_18071,N_13914);
or U22537 (N_22537,N_13069,N_12868);
or U22538 (N_22538,N_16665,N_15047);
and U22539 (N_22539,N_15642,N_18160);
nand U22540 (N_22540,N_13250,N_17776);
nand U22541 (N_22541,N_16952,N_16558);
and U22542 (N_22542,N_15764,N_15291);
xnor U22543 (N_22543,N_14639,N_18652);
nand U22544 (N_22544,N_18365,N_12523);
and U22545 (N_22545,N_17898,N_15865);
xor U22546 (N_22546,N_17195,N_14542);
nor U22547 (N_22547,N_14769,N_14905);
or U22548 (N_22548,N_17660,N_16290);
or U22549 (N_22549,N_18697,N_16789);
nand U22550 (N_22550,N_13478,N_16173);
xnor U22551 (N_22551,N_16265,N_16858);
nand U22552 (N_22552,N_12894,N_13635);
nor U22553 (N_22553,N_18740,N_14459);
xnor U22554 (N_22554,N_13199,N_15343);
nand U22555 (N_22555,N_18609,N_15982);
or U22556 (N_22556,N_14407,N_12838);
and U22557 (N_22557,N_12746,N_18327);
nand U22558 (N_22558,N_14295,N_15630);
and U22559 (N_22559,N_17474,N_13999);
nor U22560 (N_22560,N_16275,N_12565);
and U22561 (N_22561,N_15015,N_14408);
nor U22562 (N_22562,N_17935,N_17271);
nor U22563 (N_22563,N_17562,N_13930);
nand U22564 (N_22564,N_14458,N_14517);
or U22565 (N_22565,N_16536,N_15191);
nor U22566 (N_22566,N_13725,N_14463);
nand U22567 (N_22567,N_16502,N_16568);
or U22568 (N_22568,N_14612,N_12809);
xnor U22569 (N_22569,N_14978,N_15619);
or U22570 (N_22570,N_14925,N_17499);
or U22571 (N_22571,N_16906,N_15409);
nor U22572 (N_22572,N_12642,N_15472);
nor U22573 (N_22573,N_12885,N_15449);
nor U22574 (N_22574,N_13524,N_13196);
or U22575 (N_22575,N_16441,N_17406);
and U22576 (N_22576,N_18564,N_16617);
nand U22577 (N_22577,N_14517,N_18602);
nand U22578 (N_22578,N_17942,N_18386);
or U22579 (N_22579,N_14539,N_17211);
nor U22580 (N_22580,N_14344,N_15109);
or U22581 (N_22581,N_13876,N_14072);
or U22582 (N_22582,N_14983,N_15081);
xnor U22583 (N_22583,N_16340,N_13785);
nor U22584 (N_22584,N_13360,N_15427);
nor U22585 (N_22585,N_14975,N_18503);
nand U22586 (N_22586,N_12640,N_15617);
nor U22587 (N_22587,N_14979,N_15716);
nor U22588 (N_22588,N_13368,N_14984);
nand U22589 (N_22589,N_18654,N_14511);
and U22590 (N_22590,N_16663,N_15665);
xor U22591 (N_22591,N_15976,N_15669);
or U22592 (N_22592,N_18314,N_17515);
or U22593 (N_22593,N_17855,N_17691);
xnor U22594 (N_22594,N_12856,N_18319);
or U22595 (N_22595,N_13983,N_13337);
and U22596 (N_22596,N_14876,N_12909);
xnor U22597 (N_22597,N_17996,N_17493);
and U22598 (N_22598,N_14906,N_17721);
xnor U22599 (N_22599,N_13710,N_15077);
xor U22600 (N_22600,N_16925,N_14535);
nand U22601 (N_22601,N_14466,N_16673);
nor U22602 (N_22602,N_17187,N_16719);
or U22603 (N_22603,N_18717,N_18218);
and U22604 (N_22604,N_13556,N_13165);
xor U22605 (N_22605,N_12679,N_18049);
or U22606 (N_22606,N_14625,N_13959);
or U22607 (N_22607,N_18523,N_13354);
xor U22608 (N_22608,N_17007,N_18700);
and U22609 (N_22609,N_14358,N_15172);
xor U22610 (N_22610,N_16781,N_17056);
or U22611 (N_22611,N_14248,N_13784);
nand U22612 (N_22612,N_18377,N_15421);
xor U22613 (N_22613,N_13858,N_15995);
nor U22614 (N_22614,N_16514,N_14885);
or U22615 (N_22615,N_13036,N_16369);
and U22616 (N_22616,N_16434,N_16984);
and U22617 (N_22617,N_15705,N_14836);
or U22618 (N_22618,N_18275,N_17608);
and U22619 (N_22619,N_17443,N_14365);
or U22620 (N_22620,N_12816,N_18335);
or U22621 (N_22621,N_15042,N_18613);
nand U22622 (N_22622,N_13301,N_16366);
xnor U22623 (N_22623,N_16497,N_15187);
and U22624 (N_22624,N_13016,N_17585);
and U22625 (N_22625,N_17788,N_18201);
and U22626 (N_22626,N_12731,N_14950);
nor U22627 (N_22627,N_16081,N_18053);
and U22628 (N_22628,N_16218,N_14817);
xnor U22629 (N_22629,N_18170,N_14194);
or U22630 (N_22630,N_16835,N_17871);
xnor U22631 (N_22631,N_14527,N_12909);
nor U22632 (N_22632,N_14123,N_14577);
or U22633 (N_22633,N_18106,N_14930);
and U22634 (N_22634,N_12787,N_15627);
and U22635 (N_22635,N_13720,N_12760);
xnor U22636 (N_22636,N_13861,N_13962);
xor U22637 (N_22637,N_12859,N_17980);
and U22638 (N_22638,N_14309,N_13983);
nand U22639 (N_22639,N_18716,N_14106);
nand U22640 (N_22640,N_13945,N_16171);
nor U22641 (N_22641,N_18645,N_18692);
nor U22642 (N_22642,N_16951,N_17569);
nor U22643 (N_22643,N_14149,N_15544);
xnor U22644 (N_22644,N_18739,N_15765);
nand U22645 (N_22645,N_16502,N_14445);
and U22646 (N_22646,N_12737,N_17391);
nand U22647 (N_22647,N_12638,N_17988);
or U22648 (N_22648,N_18677,N_13945);
xnor U22649 (N_22649,N_12611,N_13293);
or U22650 (N_22650,N_18225,N_15672);
or U22651 (N_22651,N_17102,N_16050);
nand U22652 (N_22652,N_18053,N_16359);
and U22653 (N_22653,N_12613,N_15981);
or U22654 (N_22654,N_17820,N_16592);
or U22655 (N_22655,N_15980,N_15282);
or U22656 (N_22656,N_15161,N_17053);
and U22657 (N_22657,N_18558,N_14584);
nand U22658 (N_22658,N_16295,N_13395);
or U22659 (N_22659,N_13718,N_17609);
and U22660 (N_22660,N_18735,N_14816);
and U22661 (N_22661,N_13305,N_15476);
xor U22662 (N_22662,N_14594,N_13805);
nand U22663 (N_22663,N_18691,N_15638);
nor U22664 (N_22664,N_16387,N_13630);
nand U22665 (N_22665,N_13253,N_14091);
nor U22666 (N_22666,N_15922,N_13931);
nand U22667 (N_22667,N_17793,N_12831);
nand U22668 (N_22668,N_13534,N_12826);
and U22669 (N_22669,N_13957,N_14860);
nor U22670 (N_22670,N_15721,N_14746);
nor U22671 (N_22671,N_14214,N_15681);
nor U22672 (N_22672,N_17086,N_16622);
or U22673 (N_22673,N_13164,N_18682);
xor U22674 (N_22674,N_13528,N_15744);
and U22675 (N_22675,N_18170,N_16372);
nor U22676 (N_22676,N_16253,N_18072);
xnor U22677 (N_22677,N_14850,N_14213);
or U22678 (N_22678,N_12553,N_12640);
and U22679 (N_22679,N_15302,N_16788);
xnor U22680 (N_22680,N_14252,N_18436);
nor U22681 (N_22681,N_14541,N_18020);
nand U22682 (N_22682,N_18196,N_16376);
nor U22683 (N_22683,N_13867,N_16344);
nand U22684 (N_22684,N_15149,N_15883);
and U22685 (N_22685,N_16325,N_17011);
or U22686 (N_22686,N_14294,N_16805);
and U22687 (N_22687,N_17940,N_16188);
or U22688 (N_22688,N_13913,N_18511);
nand U22689 (N_22689,N_12887,N_17621);
xor U22690 (N_22690,N_13178,N_16169);
xor U22691 (N_22691,N_17698,N_12841);
nand U22692 (N_22692,N_12703,N_16999);
xnor U22693 (N_22693,N_17755,N_15908);
or U22694 (N_22694,N_14162,N_14053);
or U22695 (N_22695,N_13550,N_13734);
and U22696 (N_22696,N_13164,N_15429);
xnor U22697 (N_22697,N_15906,N_15933);
xnor U22698 (N_22698,N_15816,N_12613);
and U22699 (N_22699,N_17375,N_14414);
nor U22700 (N_22700,N_13225,N_16020);
nor U22701 (N_22701,N_14106,N_18301);
xnor U22702 (N_22702,N_13172,N_12875);
nor U22703 (N_22703,N_18663,N_17429);
and U22704 (N_22704,N_15207,N_17613);
and U22705 (N_22705,N_14943,N_14994);
nand U22706 (N_22706,N_14732,N_12562);
or U22707 (N_22707,N_14852,N_16988);
and U22708 (N_22708,N_14953,N_15515);
xnor U22709 (N_22709,N_16922,N_17731);
and U22710 (N_22710,N_15700,N_13715);
or U22711 (N_22711,N_13083,N_17564);
nor U22712 (N_22712,N_17586,N_16025);
and U22713 (N_22713,N_13399,N_12763);
nand U22714 (N_22714,N_12884,N_13766);
nand U22715 (N_22715,N_15158,N_13985);
and U22716 (N_22716,N_13604,N_18031);
xor U22717 (N_22717,N_13238,N_16325);
and U22718 (N_22718,N_17825,N_14772);
xnor U22719 (N_22719,N_13127,N_15974);
xnor U22720 (N_22720,N_14143,N_18637);
xnor U22721 (N_22721,N_17240,N_18054);
nor U22722 (N_22722,N_18218,N_13327);
nand U22723 (N_22723,N_13929,N_17710);
xor U22724 (N_22724,N_14377,N_15696);
nand U22725 (N_22725,N_12584,N_13537);
nand U22726 (N_22726,N_15839,N_14255);
or U22727 (N_22727,N_15177,N_17555);
and U22728 (N_22728,N_12706,N_14591);
nand U22729 (N_22729,N_12949,N_16422);
nor U22730 (N_22730,N_13856,N_12823);
xor U22731 (N_22731,N_12893,N_13522);
nor U22732 (N_22732,N_17983,N_16238);
nor U22733 (N_22733,N_18612,N_14883);
nor U22734 (N_22734,N_14250,N_12574);
xor U22735 (N_22735,N_13022,N_16423);
xor U22736 (N_22736,N_12644,N_14019);
nand U22737 (N_22737,N_17128,N_12946);
or U22738 (N_22738,N_16630,N_17839);
or U22739 (N_22739,N_14368,N_16872);
or U22740 (N_22740,N_18231,N_17622);
or U22741 (N_22741,N_15734,N_12984);
and U22742 (N_22742,N_18647,N_15813);
and U22743 (N_22743,N_13037,N_14956);
nand U22744 (N_22744,N_16689,N_13765);
xor U22745 (N_22745,N_18036,N_15785);
and U22746 (N_22746,N_17238,N_18110);
nand U22747 (N_22747,N_14004,N_13824);
nor U22748 (N_22748,N_15016,N_14288);
nand U22749 (N_22749,N_16145,N_13587);
or U22750 (N_22750,N_14090,N_14275);
and U22751 (N_22751,N_16282,N_15935);
and U22752 (N_22752,N_14283,N_13213);
nor U22753 (N_22753,N_14176,N_13224);
nand U22754 (N_22754,N_17820,N_17356);
and U22755 (N_22755,N_17621,N_16051);
nand U22756 (N_22756,N_14135,N_14695);
and U22757 (N_22757,N_12560,N_15407);
nor U22758 (N_22758,N_17648,N_15775);
nor U22759 (N_22759,N_12535,N_15874);
or U22760 (N_22760,N_14982,N_17544);
nor U22761 (N_22761,N_12664,N_14672);
nor U22762 (N_22762,N_12700,N_18649);
nor U22763 (N_22763,N_14381,N_15017);
nor U22764 (N_22764,N_13874,N_14909);
and U22765 (N_22765,N_17385,N_14753);
or U22766 (N_22766,N_13281,N_17925);
nand U22767 (N_22767,N_13858,N_14948);
nor U22768 (N_22768,N_12937,N_17933);
nor U22769 (N_22769,N_18499,N_16730);
and U22770 (N_22770,N_15613,N_15336);
or U22771 (N_22771,N_15074,N_16954);
or U22772 (N_22772,N_18614,N_18659);
xnor U22773 (N_22773,N_18170,N_14838);
or U22774 (N_22774,N_12563,N_16282);
nand U22775 (N_22775,N_16797,N_15057);
and U22776 (N_22776,N_15412,N_13967);
xor U22777 (N_22777,N_12570,N_14142);
nand U22778 (N_22778,N_14889,N_17382);
xnor U22779 (N_22779,N_12545,N_13755);
xor U22780 (N_22780,N_15584,N_15352);
nor U22781 (N_22781,N_12665,N_16641);
xor U22782 (N_22782,N_13746,N_17020);
nand U22783 (N_22783,N_18346,N_15678);
and U22784 (N_22784,N_17655,N_16388);
and U22785 (N_22785,N_12682,N_14610);
and U22786 (N_22786,N_16135,N_13857);
xor U22787 (N_22787,N_13262,N_13982);
nor U22788 (N_22788,N_14565,N_13860);
xor U22789 (N_22789,N_13667,N_15876);
nand U22790 (N_22790,N_17977,N_12776);
or U22791 (N_22791,N_16759,N_14027);
nand U22792 (N_22792,N_17860,N_13462);
nor U22793 (N_22793,N_12519,N_15049);
nand U22794 (N_22794,N_16154,N_14771);
and U22795 (N_22795,N_15149,N_13204);
xnor U22796 (N_22796,N_15330,N_16610);
xor U22797 (N_22797,N_17012,N_17873);
and U22798 (N_22798,N_16516,N_15090);
xnor U22799 (N_22799,N_12706,N_14374);
nand U22800 (N_22800,N_14912,N_13482);
nand U22801 (N_22801,N_14351,N_17243);
nand U22802 (N_22802,N_18522,N_14613);
nor U22803 (N_22803,N_17747,N_16831);
xnor U22804 (N_22804,N_14870,N_16940);
or U22805 (N_22805,N_16228,N_15538);
xnor U22806 (N_22806,N_15026,N_17805);
or U22807 (N_22807,N_13890,N_13933);
nor U22808 (N_22808,N_15129,N_16093);
nand U22809 (N_22809,N_18409,N_17407);
xor U22810 (N_22810,N_15309,N_18583);
nand U22811 (N_22811,N_14582,N_17453);
and U22812 (N_22812,N_16957,N_13455);
or U22813 (N_22813,N_12564,N_14254);
or U22814 (N_22814,N_14995,N_18082);
nand U22815 (N_22815,N_17920,N_13351);
and U22816 (N_22816,N_15181,N_15299);
and U22817 (N_22817,N_14982,N_18594);
nand U22818 (N_22818,N_12875,N_15896);
and U22819 (N_22819,N_16285,N_17175);
xor U22820 (N_22820,N_15931,N_12725);
xnor U22821 (N_22821,N_14753,N_14711);
nor U22822 (N_22822,N_15829,N_14515);
and U22823 (N_22823,N_15506,N_15258);
nand U22824 (N_22824,N_17977,N_15913);
and U22825 (N_22825,N_16892,N_15823);
nand U22826 (N_22826,N_15592,N_16368);
nor U22827 (N_22827,N_15544,N_12786);
and U22828 (N_22828,N_13249,N_14730);
nor U22829 (N_22829,N_15233,N_15528);
and U22830 (N_22830,N_16392,N_15920);
nand U22831 (N_22831,N_15089,N_15873);
or U22832 (N_22832,N_16623,N_16108);
nor U22833 (N_22833,N_17228,N_13806);
nand U22834 (N_22834,N_13495,N_13673);
or U22835 (N_22835,N_18246,N_12843);
xnor U22836 (N_22836,N_18556,N_15055);
nor U22837 (N_22837,N_18707,N_15073);
and U22838 (N_22838,N_18303,N_16109);
xnor U22839 (N_22839,N_15667,N_14949);
or U22840 (N_22840,N_18709,N_16629);
and U22841 (N_22841,N_17074,N_14900);
and U22842 (N_22842,N_15050,N_13644);
nand U22843 (N_22843,N_17506,N_17468);
and U22844 (N_22844,N_16543,N_12910);
or U22845 (N_22845,N_17241,N_17765);
nor U22846 (N_22846,N_17759,N_15878);
or U22847 (N_22847,N_12632,N_17144);
xor U22848 (N_22848,N_14765,N_13597);
nand U22849 (N_22849,N_18553,N_18462);
nand U22850 (N_22850,N_15658,N_16944);
nor U22851 (N_22851,N_17357,N_14303);
xnor U22852 (N_22852,N_14675,N_13708);
nor U22853 (N_22853,N_12561,N_15593);
nor U22854 (N_22854,N_17539,N_16702);
nor U22855 (N_22855,N_15417,N_17193);
nor U22856 (N_22856,N_12517,N_16544);
or U22857 (N_22857,N_12511,N_18193);
nor U22858 (N_22858,N_12678,N_14717);
xor U22859 (N_22859,N_14262,N_18738);
or U22860 (N_22860,N_17755,N_13689);
nor U22861 (N_22861,N_16473,N_13730);
nand U22862 (N_22862,N_12753,N_14959);
nor U22863 (N_22863,N_16218,N_13688);
nand U22864 (N_22864,N_15758,N_14718);
nor U22865 (N_22865,N_15656,N_15348);
nand U22866 (N_22866,N_17777,N_12823);
nand U22867 (N_22867,N_18677,N_15154);
nor U22868 (N_22868,N_14527,N_16085);
xnor U22869 (N_22869,N_17107,N_15290);
and U22870 (N_22870,N_16042,N_15083);
nor U22871 (N_22871,N_16943,N_12621);
or U22872 (N_22872,N_18252,N_15865);
or U22873 (N_22873,N_13515,N_16617);
xnor U22874 (N_22874,N_13309,N_15773);
nand U22875 (N_22875,N_14004,N_16904);
nor U22876 (N_22876,N_12799,N_15417);
nand U22877 (N_22877,N_15647,N_15262);
or U22878 (N_22878,N_16137,N_17260);
nor U22879 (N_22879,N_13632,N_15062);
or U22880 (N_22880,N_15547,N_17914);
nor U22881 (N_22881,N_13993,N_16009);
xnor U22882 (N_22882,N_16715,N_17270);
nor U22883 (N_22883,N_18648,N_13940);
xor U22884 (N_22884,N_18708,N_18155);
xor U22885 (N_22885,N_17799,N_16814);
and U22886 (N_22886,N_14678,N_14834);
nand U22887 (N_22887,N_14743,N_17676);
nand U22888 (N_22888,N_17955,N_13533);
nor U22889 (N_22889,N_17678,N_12889);
or U22890 (N_22890,N_17182,N_16674);
nor U22891 (N_22891,N_15652,N_15538);
xor U22892 (N_22892,N_17671,N_14496);
and U22893 (N_22893,N_18161,N_14220);
or U22894 (N_22894,N_15841,N_15347);
and U22895 (N_22895,N_16555,N_16670);
or U22896 (N_22896,N_13649,N_15359);
xor U22897 (N_22897,N_15424,N_18399);
xnor U22898 (N_22898,N_18627,N_16999);
nand U22899 (N_22899,N_12545,N_17290);
xor U22900 (N_22900,N_12530,N_14677);
or U22901 (N_22901,N_15799,N_15781);
or U22902 (N_22902,N_18109,N_15609);
nor U22903 (N_22903,N_16715,N_15638);
xnor U22904 (N_22904,N_13685,N_13864);
and U22905 (N_22905,N_16175,N_13055);
or U22906 (N_22906,N_14147,N_16874);
nand U22907 (N_22907,N_16953,N_12885);
and U22908 (N_22908,N_13487,N_18534);
or U22909 (N_22909,N_18155,N_16680);
or U22910 (N_22910,N_13646,N_14786);
nand U22911 (N_22911,N_16545,N_12842);
and U22912 (N_22912,N_13518,N_13849);
xnor U22913 (N_22913,N_14344,N_14913);
and U22914 (N_22914,N_17893,N_14328);
nor U22915 (N_22915,N_17813,N_16748);
nand U22916 (N_22916,N_17557,N_17764);
or U22917 (N_22917,N_18471,N_14120);
nor U22918 (N_22918,N_13456,N_15331);
nand U22919 (N_22919,N_14707,N_18139);
or U22920 (N_22920,N_18637,N_15053);
nand U22921 (N_22921,N_16151,N_13794);
nand U22922 (N_22922,N_16547,N_14689);
nand U22923 (N_22923,N_18725,N_17279);
nand U22924 (N_22924,N_13317,N_16694);
or U22925 (N_22925,N_14777,N_12765);
and U22926 (N_22926,N_16182,N_18528);
or U22927 (N_22927,N_15476,N_18379);
nand U22928 (N_22928,N_17367,N_15951);
xor U22929 (N_22929,N_15399,N_14074);
xnor U22930 (N_22930,N_17854,N_18108);
or U22931 (N_22931,N_14224,N_14441);
nor U22932 (N_22932,N_15039,N_14486);
or U22933 (N_22933,N_18215,N_14072);
xor U22934 (N_22934,N_14121,N_15348);
nor U22935 (N_22935,N_17889,N_15596);
xnor U22936 (N_22936,N_17227,N_12717);
and U22937 (N_22937,N_13234,N_17393);
xnor U22938 (N_22938,N_16929,N_15987);
and U22939 (N_22939,N_12986,N_16020);
nor U22940 (N_22940,N_18405,N_17315);
nor U22941 (N_22941,N_13797,N_15186);
nand U22942 (N_22942,N_13717,N_13035);
nand U22943 (N_22943,N_15422,N_14695);
xnor U22944 (N_22944,N_12506,N_17698);
nor U22945 (N_22945,N_16440,N_15495);
nand U22946 (N_22946,N_14193,N_13326);
or U22947 (N_22947,N_16904,N_14466);
and U22948 (N_22948,N_16306,N_16258);
and U22949 (N_22949,N_15167,N_13850);
nor U22950 (N_22950,N_16194,N_15496);
or U22951 (N_22951,N_14032,N_15478);
and U22952 (N_22952,N_15393,N_16231);
nor U22953 (N_22953,N_15072,N_12763);
and U22954 (N_22954,N_17542,N_14184);
nand U22955 (N_22955,N_14955,N_15038);
nor U22956 (N_22956,N_15662,N_15291);
or U22957 (N_22957,N_15188,N_18619);
or U22958 (N_22958,N_16988,N_18180);
and U22959 (N_22959,N_13950,N_18472);
nand U22960 (N_22960,N_15911,N_13464);
nand U22961 (N_22961,N_12845,N_17384);
or U22962 (N_22962,N_12606,N_13346);
or U22963 (N_22963,N_14128,N_17540);
or U22964 (N_22964,N_14639,N_14798);
and U22965 (N_22965,N_12750,N_18187);
nand U22966 (N_22966,N_15278,N_14578);
xor U22967 (N_22967,N_13141,N_15675);
xor U22968 (N_22968,N_16021,N_18116);
and U22969 (N_22969,N_12909,N_17138);
nand U22970 (N_22970,N_14005,N_15257);
nand U22971 (N_22971,N_13852,N_14049);
nand U22972 (N_22972,N_17350,N_14767);
or U22973 (N_22973,N_13282,N_13715);
xor U22974 (N_22974,N_14342,N_17421);
xor U22975 (N_22975,N_15628,N_14679);
xnor U22976 (N_22976,N_15902,N_16624);
nor U22977 (N_22977,N_17600,N_14638);
xor U22978 (N_22978,N_17845,N_15272);
and U22979 (N_22979,N_14751,N_17227);
nor U22980 (N_22980,N_13129,N_14059);
nor U22981 (N_22981,N_16278,N_17443);
nand U22982 (N_22982,N_14727,N_16292);
nor U22983 (N_22983,N_14378,N_14318);
or U22984 (N_22984,N_14582,N_14480);
and U22985 (N_22985,N_17188,N_14903);
nand U22986 (N_22986,N_15590,N_14645);
or U22987 (N_22987,N_13078,N_18405);
nor U22988 (N_22988,N_15040,N_12822);
nand U22989 (N_22989,N_18427,N_13763);
xnor U22990 (N_22990,N_17976,N_15182);
nand U22991 (N_22991,N_14584,N_15255);
nand U22992 (N_22992,N_13694,N_14943);
nor U22993 (N_22993,N_13226,N_18385);
and U22994 (N_22994,N_17807,N_16047);
xnor U22995 (N_22995,N_12987,N_15135);
and U22996 (N_22996,N_14514,N_16014);
or U22997 (N_22997,N_17791,N_13723);
nand U22998 (N_22998,N_14826,N_18330);
nand U22999 (N_22999,N_18573,N_13723);
nor U23000 (N_23000,N_18604,N_16946);
or U23001 (N_23001,N_14836,N_14981);
and U23002 (N_23002,N_13836,N_15991);
or U23003 (N_23003,N_16922,N_14430);
or U23004 (N_23004,N_13577,N_18015);
nor U23005 (N_23005,N_13459,N_17058);
nand U23006 (N_23006,N_15821,N_13454);
or U23007 (N_23007,N_14240,N_12958);
nor U23008 (N_23008,N_15267,N_13120);
nor U23009 (N_23009,N_18727,N_14942);
or U23010 (N_23010,N_15226,N_14488);
nor U23011 (N_23011,N_12734,N_18451);
and U23012 (N_23012,N_16746,N_18376);
nor U23013 (N_23013,N_17070,N_17040);
or U23014 (N_23014,N_12733,N_17097);
nand U23015 (N_23015,N_14176,N_14472);
or U23016 (N_23016,N_13377,N_14277);
and U23017 (N_23017,N_15512,N_13124);
xnor U23018 (N_23018,N_13161,N_14695);
nand U23019 (N_23019,N_13508,N_12632);
and U23020 (N_23020,N_18501,N_15448);
nor U23021 (N_23021,N_17242,N_14510);
and U23022 (N_23022,N_18471,N_12737);
nand U23023 (N_23023,N_14197,N_17540);
or U23024 (N_23024,N_13448,N_17928);
and U23025 (N_23025,N_17332,N_14339);
nor U23026 (N_23026,N_14679,N_13460);
and U23027 (N_23027,N_15829,N_13006);
nor U23028 (N_23028,N_14927,N_15229);
and U23029 (N_23029,N_16136,N_14226);
and U23030 (N_23030,N_16781,N_13108);
nor U23031 (N_23031,N_13420,N_17237);
xnor U23032 (N_23032,N_14433,N_16291);
nand U23033 (N_23033,N_17966,N_15332);
xnor U23034 (N_23034,N_16594,N_14284);
or U23035 (N_23035,N_18312,N_14348);
or U23036 (N_23036,N_18725,N_16995);
or U23037 (N_23037,N_16360,N_15984);
nor U23038 (N_23038,N_12849,N_18402);
xor U23039 (N_23039,N_12507,N_14549);
nand U23040 (N_23040,N_18147,N_15964);
nand U23041 (N_23041,N_13774,N_14653);
xnor U23042 (N_23042,N_18529,N_13291);
nand U23043 (N_23043,N_17737,N_13950);
and U23044 (N_23044,N_18383,N_13409);
nand U23045 (N_23045,N_13479,N_15017);
nor U23046 (N_23046,N_14613,N_17934);
and U23047 (N_23047,N_14068,N_13982);
and U23048 (N_23048,N_15092,N_13306);
nor U23049 (N_23049,N_14505,N_12785);
nand U23050 (N_23050,N_15730,N_17562);
and U23051 (N_23051,N_17067,N_16160);
and U23052 (N_23052,N_12689,N_17367);
or U23053 (N_23053,N_15561,N_12593);
nor U23054 (N_23054,N_18458,N_17827);
and U23055 (N_23055,N_12877,N_15210);
or U23056 (N_23056,N_16444,N_14790);
or U23057 (N_23057,N_16345,N_15010);
xnor U23058 (N_23058,N_16963,N_13793);
nand U23059 (N_23059,N_16316,N_17279);
or U23060 (N_23060,N_18461,N_16299);
nand U23061 (N_23061,N_13162,N_14162);
xnor U23062 (N_23062,N_13893,N_13896);
and U23063 (N_23063,N_18087,N_15020);
xnor U23064 (N_23064,N_18403,N_12854);
nor U23065 (N_23065,N_14205,N_15768);
xor U23066 (N_23066,N_17390,N_15030);
xnor U23067 (N_23067,N_18732,N_16966);
xnor U23068 (N_23068,N_15174,N_17455);
and U23069 (N_23069,N_12552,N_16218);
nor U23070 (N_23070,N_18535,N_18203);
nand U23071 (N_23071,N_18223,N_15889);
nor U23072 (N_23072,N_17802,N_13368);
and U23073 (N_23073,N_14847,N_17958);
and U23074 (N_23074,N_18603,N_13411);
or U23075 (N_23075,N_15186,N_14044);
nand U23076 (N_23076,N_13961,N_17647);
xor U23077 (N_23077,N_15424,N_18496);
xnor U23078 (N_23078,N_16254,N_13268);
nor U23079 (N_23079,N_18652,N_16223);
nand U23080 (N_23080,N_13687,N_16550);
nand U23081 (N_23081,N_13799,N_15807);
nor U23082 (N_23082,N_15084,N_16206);
or U23083 (N_23083,N_15971,N_17901);
and U23084 (N_23084,N_12953,N_16697);
nor U23085 (N_23085,N_13600,N_15993);
and U23086 (N_23086,N_14519,N_14408);
nand U23087 (N_23087,N_13326,N_17475);
nand U23088 (N_23088,N_17838,N_16076);
or U23089 (N_23089,N_18561,N_14184);
or U23090 (N_23090,N_13023,N_15905);
or U23091 (N_23091,N_17719,N_16888);
or U23092 (N_23092,N_14101,N_17791);
xor U23093 (N_23093,N_18398,N_13161);
xnor U23094 (N_23094,N_16923,N_13077);
nand U23095 (N_23095,N_12977,N_12756);
xnor U23096 (N_23096,N_14772,N_13294);
and U23097 (N_23097,N_18495,N_17239);
and U23098 (N_23098,N_14172,N_15089);
nor U23099 (N_23099,N_16803,N_12644);
or U23100 (N_23100,N_16307,N_13071);
nor U23101 (N_23101,N_16519,N_15073);
nor U23102 (N_23102,N_16861,N_12581);
xor U23103 (N_23103,N_14809,N_12982);
nand U23104 (N_23104,N_18315,N_14580);
nor U23105 (N_23105,N_17412,N_17418);
and U23106 (N_23106,N_12892,N_15108);
nand U23107 (N_23107,N_18705,N_16902);
nor U23108 (N_23108,N_15158,N_16514);
nand U23109 (N_23109,N_17437,N_18580);
xor U23110 (N_23110,N_17678,N_14935);
nand U23111 (N_23111,N_13940,N_17559);
nor U23112 (N_23112,N_18220,N_13396);
xor U23113 (N_23113,N_16194,N_18587);
nor U23114 (N_23114,N_12910,N_18122);
and U23115 (N_23115,N_13142,N_13275);
or U23116 (N_23116,N_16126,N_18572);
or U23117 (N_23117,N_16574,N_15378);
nor U23118 (N_23118,N_16120,N_14971);
and U23119 (N_23119,N_17317,N_17524);
nor U23120 (N_23120,N_18327,N_12735);
xnor U23121 (N_23121,N_13527,N_16125);
nand U23122 (N_23122,N_15072,N_15138);
and U23123 (N_23123,N_17676,N_16452);
and U23124 (N_23124,N_14331,N_12863);
nand U23125 (N_23125,N_18221,N_17580);
nand U23126 (N_23126,N_17918,N_12634);
xor U23127 (N_23127,N_12676,N_17579);
xor U23128 (N_23128,N_15957,N_14655);
nand U23129 (N_23129,N_15445,N_17969);
nor U23130 (N_23130,N_16517,N_16876);
xnor U23131 (N_23131,N_13319,N_15096);
nor U23132 (N_23132,N_15745,N_14541);
and U23133 (N_23133,N_14147,N_17786);
xor U23134 (N_23134,N_13405,N_13915);
nor U23135 (N_23135,N_12770,N_16434);
nor U23136 (N_23136,N_13185,N_12747);
nand U23137 (N_23137,N_17328,N_17863);
nor U23138 (N_23138,N_12555,N_13080);
nor U23139 (N_23139,N_16646,N_12904);
and U23140 (N_23140,N_17619,N_14068);
xnor U23141 (N_23141,N_12735,N_13106);
or U23142 (N_23142,N_13067,N_16079);
and U23143 (N_23143,N_14570,N_18627);
nand U23144 (N_23144,N_14144,N_17548);
nor U23145 (N_23145,N_14834,N_12741);
and U23146 (N_23146,N_12992,N_15797);
or U23147 (N_23147,N_17903,N_18252);
and U23148 (N_23148,N_13683,N_17751);
nor U23149 (N_23149,N_15362,N_17332);
nor U23150 (N_23150,N_17833,N_14039);
and U23151 (N_23151,N_17305,N_17079);
nor U23152 (N_23152,N_18744,N_15804);
xnor U23153 (N_23153,N_15609,N_17383);
nand U23154 (N_23154,N_17864,N_17986);
nor U23155 (N_23155,N_12835,N_18591);
or U23156 (N_23156,N_12671,N_16846);
nand U23157 (N_23157,N_15949,N_14956);
nor U23158 (N_23158,N_16482,N_15459);
or U23159 (N_23159,N_15124,N_14516);
xnor U23160 (N_23160,N_15937,N_13431);
xor U23161 (N_23161,N_12508,N_13605);
and U23162 (N_23162,N_16737,N_12565);
or U23163 (N_23163,N_16644,N_13608);
nand U23164 (N_23164,N_13323,N_13961);
nand U23165 (N_23165,N_12510,N_18737);
and U23166 (N_23166,N_15652,N_17824);
and U23167 (N_23167,N_17253,N_12751);
nand U23168 (N_23168,N_15252,N_13262);
or U23169 (N_23169,N_12536,N_15642);
xnor U23170 (N_23170,N_18486,N_14026);
and U23171 (N_23171,N_13206,N_16262);
xor U23172 (N_23172,N_14021,N_13986);
and U23173 (N_23173,N_13383,N_15109);
or U23174 (N_23174,N_14174,N_18508);
or U23175 (N_23175,N_16088,N_12742);
and U23176 (N_23176,N_12970,N_16002);
xnor U23177 (N_23177,N_16590,N_15603);
and U23178 (N_23178,N_18404,N_17544);
and U23179 (N_23179,N_14391,N_14484);
and U23180 (N_23180,N_12521,N_13906);
xor U23181 (N_23181,N_16595,N_16811);
nand U23182 (N_23182,N_14368,N_17262);
xor U23183 (N_23183,N_18449,N_15496);
nand U23184 (N_23184,N_12882,N_17781);
and U23185 (N_23185,N_14771,N_17507);
nor U23186 (N_23186,N_17250,N_13439);
or U23187 (N_23187,N_16288,N_18747);
nor U23188 (N_23188,N_15882,N_13748);
or U23189 (N_23189,N_18226,N_15002);
nand U23190 (N_23190,N_15174,N_15306);
and U23191 (N_23191,N_15791,N_14606);
or U23192 (N_23192,N_12555,N_18679);
or U23193 (N_23193,N_18031,N_13411);
xnor U23194 (N_23194,N_14158,N_12813);
and U23195 (N_23195,N_14618,N_18267);
or U23196 (N_23196,N_13068,N_14683);
or U23197 (N_23197,N_16127,N_17700);
and U23198 (N_23198,N_15854,N_14233);
xor U23199 (N_23199,N_16446,N_15558);
nand U23200 (N_23200,N_15384,N_16013);
nor U23201 (N_23201,N_15170,N_13180);
nand U23202 (N_23202,N_16848,N_16453);
or U23203 (N_23203,N_15993,N_14102);
nor U23204 (N_23204,N_13358,N_14322);
nand U23205 (N_23205,N_18730,N_13701);
and U23206 (N_23206,N_18466,N_18273);
or U23207 (N_23207,N_18677,N_18202);
xnor U23208 (N_23208,N_18003,N_17224);
and U23209 (N_23209,N_18450,N_14029);
nand U23210 (N_23210,N_14816,N_15566);
nand U23211 (N_23211,N_14812,N_16614);
xnor U23212 (N_23212,N_15278,N_16913);
nor U23213 (N_23213,N_14018,N_16036);
nand U23214 (N_23214,N_16133,N_18102);
xor U23215 (N_23215,N_12581,N_13599);
and U23216 (N_23216,N_14097,N_17433);
nand U23217 (N_23217,N_16744,N_13382);
nand U23218 (N_23218,N_12515,N_14035);
or U23219 (N_23219,N_13946,N_13997);
and U23220 (N_23220,N_16266,N_18113);
or U23221 (N_23221,N_18634,N_15517);
nor U23222 (N_23222,N_14935,N_14343);
nor U23223 (N_23223,N_12585,N_15197);
or U23224 (N_23224,N_14956,N_18467);
xor U23225 (N_23225,N_15626,N_17846);
and U23226 (N_23226,N_16552,N_18344);
and U23227 (N_23227,N_13366,N_15736);
xor U23228 (N_23228,N_14124,N_13513);
nor U23229 (N_23229,N_18696,N_14183);
or U23230 (N_23230,N_18356,N_14560);
nor U23231 (N_23231,N_14365,N_17547);
nand U23232 (N_23232,N_14348,N_17896);
nand U23233 (N_23233,N_14641,N_18584);
or U23234 (N_23234,N_16250,N_15879);
or U23235 (N_23235,N_14837,N_12710);
or U23236 (N_23236,N_12723,N_12525);
xor U23237 (N_23237,N_17458,N_16563);
or U23238 (N_23238,N_16462,N_17579);
or U23239 (N_23239,N_12607,N_12791);
xor U23240 (N_23240,N_16516,N_15931);
xnor U23241 (N_23241,N_12958,N_13237);
nand U23242 (N_23242,N_17464,N_15422);
nor U23243 (N_23243,N_13958,N_17695);
xnor U23244 (N_23244,N_14503,N_16922);
nor U23245 (N_23245,N_18391,N_14147);
and U23246 (N_23246,N_14624,N_13201);
nor U23247 (N_23247,N_17901,N_14270);
and U23248 (N_23248,N_14711,N_14997);
and U23249 (N_23249,N_15493,N_18689);
or U23250 (N_23250,N_12553,N_18279);
xnor U23251 (N_23251,N_18258,N_14295);
nor U23252 (N_23252,N_18710,N_17702);
or U23253 (N_23253,N_15138,N_17231);
nand U23254 (N_23254,N_14149,N_13713);
and U23255 (N_23255,N_16759,N_18568);
or U23256 (N_23256,N_16203,N_12955);
xnor U23257 (N_23257,N_13774,N_18038);
and U23258 (N_23258,N_14502,N_15131);
xnor U23259 (N_23259,N_12857,N_15904);
or U23260 (N_23260,N_15154,N_14870);
nand U23261 (N_23261,N_13818,N_14873);
xor U23262 (N_23262,N_14631,N_14573);
and U23263 (N_23263,N_15262,N_13645);
or U23264 (N_23264,N_13802,N_14247);
and U23265 (N_23265,N_14549,N_16600);
and U23266 (N_23266,N_18226,N_16963);
and U23267 (N_23267,N_14472,N_13161);
nor U23268 (N_23268,N_18546,N_15582);
or U23269 (N_23269,N_16814,N_13142);
nor U23270 (N_23270,N_13835,N_15698);
or U23271 (N_23271,N_13842,N_12516);
nand U23272 (N_23272,N_18532,N_14612);
xor U23273 (N_23273,N_15561,N_14095);
xor U23274 (N_23274,N_13867,N_13375);
xnor U23275 (N_23275,N_18563,N_14743);
or U23276 (N_23276,N_14102,N_13992);
xor U23277 (N_23277,N_14944,N_12671);
nand U23278 (N_23278,N_13127,N_16442);
nor U23279 (N_23279,N_16886,N_15587);
xnor U23280 (N_23280,N_15610,N_14384);
xnor U23281 (N_23281,N_13055,N_15831);
nand U23282 (N_23282,N_17066,N_12969);
xor U23283 (N_23283,N_18505,N_17300);
nand U23284 (N_23284,N_15906,N_17756);
or U23285 (N_23285,N_14699,N_18694);
xnor U23286 (N_23286,N_13175,N_12747);
or U23287 (N_23287,N_13943,N_18576);
xor U23288 (N_23288,N_15725,N_15649);
nor U23289 (N_23289,N_15596,N_15071);
and U23290 (N_23290,N_12928,N_18694);
xnor U23291 (N_23291,N_15366,N_15436);
nand U23292 (N_23292,N_16439,N_15529);
nor U23293 (N_23293,N_17303,N_16868);
xor U23294 (N_23294,N_15487,N_13231);
and U23295 (N_23295,N_17214,N_16827);
nand U23296 (N_23296,N_14744,N_12835);
nor U23297 (N_23297,N_14294,N_14243);
nor U23298 (N_23298,N_18121,N_13393);
and U23299 (N_23299,N_15930,N_15310);
or U23300 (N_23300,N_14698,N_18724);
and U23301 (N_23301,N_16240,N_15352);
nand U23302 (N_23302,N_17479,N_18208);
and U23303 (N_23303,N_16422,N_16014);
or U23304 (N_23304,N_17784,N_18131);
nor U23305 (N_23305,N_14729,N_17975);
nand U23306 (N_23306,N_13882,N_18341);
or U23307 (N_23307,N_17618,N_15577);
and U23308 (N_23308,N_13437,N_15375);
nand U23309 (N_23309,N_17463,N_18696);
nand U23310 (N_23310,N_17917,N_18181);
xor U23311 (N_23311,N_18528,N_14545);
or U23312 (N_23312,N_16351,N_17788);
or U23313 (N_23313,N_14358,N_18613);
or U23314 (N_23314,N_17726,N_18612);
and U23315 (N_23315,N_14403,N_13722);
xnor U23316 (N_23316,N_13428,N_15358);
nor U23317 (N_23317,N_16533,N_17857);
or U23318 (N_23318,N_15308,N_14527);
and U23319 (N_23319,N_15645,N_13932);
or U23320 (N_23320,N_17706,N_17255);
or U23321 (N_23321,N_16998,N_12804);
nor U23322 (N_23322,N_15404,N_17660);
nand U23323 (N_23323,N_18648,N_17740);
nor U23324 (N_23324,N_14286,N_17608);
or U23325 (N_23325,N_17377,N_14022);
and U23326 (N_23326,N_15183,N_15797);
or U23327 (N_23327,N_16211,N_14141);
and U23328 (N_23328,N_14974,N_14453);
nor U23329 (N_23329,N_15525,N_18012);
xnor U23330 (N_23330,N_16695,N_16621);
xnor U23331 (N_23331,N_12997,N_12984);
or U23332 (N_23332,N_15735,N_16787);
and U23333 (N_23333,N_14607,N_12936);
and U23334 (N_23334,N_17416,N_13436);
or U23335 (N_23335,N_16365,N_15503);
nor U23336 (N_23336,N_17944,N_16687);
nor U23337 (N_23337,N_16913,N_13574);
or U23338 (N_23338,N_14290,N_13175);
or U23339 (N_23339,N_16191,N_16077);
and U23340 (N_23340,N_13843,N_17336);
or U23341 (N_23341,N_18403,N_14864);
xor U23342 (N_23342,N_15557,N_13305);
or U23343 (N_23343,N_16113,N_17373);
xor U23344 (N_23344,N_14659,N_17957);
and U23345 (N_23345,N_14197,N_15051);
nand U23346 (N_23346,N_18674,N_13482);
nor U23347 (N_23347,N_12595,N_17925);
or U23348 (N_23348,N_14866,N_14200);
nor U23349 (N_23349,N_17405,N_15848);
nor U23350 (N_23350,N_15088,N_14775);
and U23351 (N_23351,N_13638,N_12828);
and U23352 (N_23352,N_15860,N_12685);
nand U23353 (N_23353,N_14615,N_16388);
or U23354 (N_23354,N_14816,N_16828);
xnor U23355 (N_23355,N_16456,N_16967);
and U23356 (N_23356,N_16452,N_15007);
xor U23357 (N_23357,N_15660,N_13420);
nor U23358 (N_23358,N_14499,N_14384);
or U23359 (N_23359,N_14393,N_16911);
or U23360 (N_23360,N_17789,N_16443);
or U23361 (N_23361,N_17184,N_15027);
xor U23362 (N_23362,N_13815,N_13845);
nand U23363 (N_23363,N_14358,N_13833);
and U23364 (N_23364,N_12767,N_13529);
or U23365 (N_23365,N_15777,N_17211);
and U23366 (N_23366,N_12929,N_13091);
or U23367 (N_23367,N_14565,N_15674);
xor U23368 (N_23368,N_13022,N_15792);
nor U23369 (N_23369,N_16468,N_18231);
nor U23370 (N_23370,N_16660,N_14968);
or U23371 (N_23371,N_13510,N_16300);
or U23372 (N_23372,N_13599,N_17617);
nand U23373 (N_23373,N_13091,N_17115);
xor U23374 (N_23374,N_12818,N_18575);
or U23375 (N_23375,N_14981,N_14528);
nand U23376 (N_23376,N_17076,N_18209);
and U23377 (N_23377,N_13880,N_12851);
nor U23378 (N_23378,N_16674,N_14447);
and U23379 (N_23379,N_16643,N_14487);
and U23380 (N_23380,N_15667,N_16111);
nand U23381 (N_23381,N_14087,N_17493);
nand U23382 (N_23382,N_17131,N_15030);
nor U23383 (N_23383,N_17547,N_14038);
and U23384 (N_23384,N_12814,N_16935);
and U23385 (N_23385,N_15879,N_17537);
or U23386 (N_23386,N_16124,N_16652);
or U23387 (N_23387,N_14194,N_15859);
or U23388 (N_23388,N_17093,N_14230);
and U23389 (N_23389,N_17919,N_16304);
nor U23390 (N_23390,N_13139,N_13177);
or U23391 (N_23391,N_13871,N_15077);
nand U23392 (N_23392,N_14253,N_17480);
or U23393 (N_23393,N_16452,N_14176);
xor U23394 (N_23394,N_15064,N_15708);
xnor U23395 (N_23395,N_16049,N_16558);
nor U23396 (N_23396,N_12599,N_15943);
and U23397 (N_23397,N_15692,N_14038);
nand U23398 (N_23398,N_13001,N_18247);
and U23399 (N_23399,N_15956,N_16626);
nor U23400 (N_23400,N_17711,N_13182);
and U23401 (N_23401,N_14270,N_17016);
xnor U23402 (N_23402,N_17183,N_17756);
and U23403 (N_23403,N_18407,N_14313);
xnor U23404 (N_23404,N_16883,N_16938);
nor U23405 (N_23405,N_16340,N_16268);
nand U23406 (N_23406,N_12761,N_14902);
nor U23407 (N_23407,N_15012,N_15493);
or U23408 (N_23408,N_14126,N_18293);
nand U23409 (N_23409,N_14784,N_15528);
or U23410 (N_23410,N_18565,N_15344);
nand U23411 (N_23411,N_14315,N_18379);
nand U23412 (N_23412,N_15906,N_15711);
xnor U23413 (N_23413,N_18250,N_17059);
nand U23414 (N_23414,N_17482,N_16237);
nand U23415 (N_23415,N_16978,N_18523);
xnor U23416 (N_23416,N_13246,N_12865);
nand U23417 (N_23417,N_15578,N_15499);
nand U23418 (N_23418,N_17766,N_18091);
xnor U23419 (N_23419,N_14996,N_12606);
xnor U23420 (N_23420,N_17540,N_13001);
or U23421 (N_23421,N_13556,N_14178);
nand U23422 (N_23422,N_14564,N_15645);
nand U23423 (N_23423,N_13746,N_12912);
or U23424 (N_23424,N_16408,N_14243);
or U23425 (N_23425,N_18484,N_13925);
nand U23426 (N_23426,N_13290,N_15611);
nor U23427 (N_23427,N_12864,N_16430);
and U23428 (N_23428,N_13046,N_18209);
or U23429 (N_23429,N_18573,N_17753);
nor U23430 (N_23430,N_14091,N_18631);
and U23431 (N_23431,N_17337,N_12660);
nand U23432 (N_23432,N_15071,N_15718);
nand U23433 (N_23433,N_13812,N_18320);
nand U23434 (N_23434,N_17641,N_13680);
nor U23435 (N_23435,N_16078,N_17739);
nand U23436 (N_23436,N_12981,N_17905);
and U23437 (N_23437,N_18608,N_16893);
and U23438 (N_23438,N_18120,N_16056);
nor U23439 (N_23439,N_18484,N_18535);
and U23440 (N_23440,N_13921,N_18530);
nor U23441 (N_23441,N_15893,N_14499);
nand U23442 (N_23442,N_17090,N_16888);
or U23443 (N_23443,N_16487,N_12868);
or U23444 (N_23444,N_18151,N_12970);
xor U23445 (N_23445,N_14076,N_17349);
and U23446 (N_23446,N_14931,N_14612);
or U23447 (N_23447,N_13003,N_15781);
xor U23448 (N_23448,N_17199,N_17984);
nor U23449 (N_23449,N_14571,N_17790);
or U23450 (N_23450,N_16594,N_16214);
nand U23451 (N_23451,N_16795,N_17676);
or U23452 (N_23452,N_17620,N_16339);
xor U23453 (N_23453,N_12952,N_13506);
xor U23454 (N_23454,N_15591,N_14181);
xnor U23455 (N_23455,N_16544,N_12841);
nand U23456 (N_23456,N_14923,N_18354);
xnor U23457 (N_23457,N_15434,N_15163);
nor U23458 (N_23458,N_14094,N_18455);
and U23459 (N_23459,N_15916,N_14124);
xor U23460 (N_23460,N_13984,N_16611);
nand U23461 (N_23461,N_18054,N_14143);
xor U23462 (N_23462,N_16239,N_12579);
nor U23463 (N_23463,N_18270,N_16178);
nand U23464 (N_23464,N_16430,N_15253);
nand U23465 (N_23465,N_16750,N_12830);
xor U23466 (N_23466,N_17376,N_13899);
or U23467 (N_23467,N_14630,N_18240);
and U23468 (N_23468,N_17244,N_12629);
xor U23469 (N_23469,N_17984,N_12839);
nand U23470 (N_23470,N_16840,N_16048);
xor U23471 (N_23471,N_14276,N_14179);
and U23472 (N_23472,N_17584,N_13703);
nor U23473 (N_23473,N_16950,N_16894);
nor U23474 (N_23474,N_14096,N_15609);
nand U23475 (N_23475,N_16872,N_12805);
nor U23476 (N_23476,N_14324,N_17929);
xor U23477 (N_23477,N_13856,N_16710);
or U23478 (N_23478,N_16760,N_15026);
nand U23479 (N_23479,N_15213,N_18500);
or U23480 (N_23480,N_15301,N_17160);
or U23481 (N_23481,N_13210,N_14097);
nor U23482 (N_23482,N_18317,N_12734);
xor U23483 (N_23483,N_12885,N_13900);
and U23484 (N_23484,N_14387,N_18227);
nor U23485 (N_23485,N_13456,N_18335);
nand U23486 (N_23486,N_15731,N_15332);
or U23487 (N_23487,N_14632,N_13496);
or U23488 (N_23488,N_18685,N_18484);
or U23489 (N_23489,N_18091,N_18708);
and U23490 (N_23490,N_14124,N_15891);
and U23491 (N_23491,N_13928,N_13707);
and U23492 (N_23492,N_13004,N_18213);
xnor U23493 (N_23493,N_14819,N_16303);
xor U23494 (N_23494,N_15791,N_17515);
or U23495 (N_23495,N_18092,N_13767);
and U23496 (N_23496,N_18488,N_14992);
nor U23497 (N_23497,N_14846,N_17841);
and U23498 (N_23498,N_14305,N_16849);
and U23499 (N_23499,N_16595,N_16681);
and U23500 (N_23500,N_14009,N_14217);
nor U23501 (N_23501,N_14236,N_13262);
nor U23502 (N_23502,N_16188,N_13807);
xnor U23503 (N_23503,N_17153,N_16100);
nand U23504 (N_23504,N_13929,N_16330);
nor U23505 (N_23505,N_14363,N_17732);
or U23506 (N_23506,N_13272,N_17184);
nand U23507 (N_23507,N_13826,N_16451);
or U23508 (N_23508,N_14031,N_14845);
or U23509 (N_23509,N_15307,N_13963);
xnor U23510 (N_23510,N_17545,N_14464);
nor U23511 (N_23511,N_14575,N_16030);
nand U23512 (N_23512,N_14734,N_17182);
nor U23513 (N_23513,N_15891,N_17752);
and U23514 (N_23514,N_15645,N_14054);
xnor U23515 (N_23515,N_15277,N_16908);
or U23516 (N_23516,N_17651,N_13618);
nor U23517 (N_23517,N_15208,N_12766);
nand U23518 (N_23518,N_18294,N_13235);
nor U23519 (N_23519,N_16724,N_18326);
xor U23520 (N_23520,N_18705,N_12913);
nand U23521 (N_23521,N_16361,N_15879);
xor U23522 (N_23522,N_15571,N_18677);
xnor U23523 (N_23523,N_17522,N_17891);
or U23524 (N_23524,N_18311,N_12511);
nor U23525 (N_23525,N_13386,N_15205);
and U23526 (N_23526,N_16497,N_18004);
nor U23527 (N_23527,N_16009,N_17436);
and U23528 (N_23528,N_13271,N_15548);
nor U23529 (N_23529,N_17000,N_15415);
nand U23530 (N_23530,N_15370,N_15466);
nor U23531 (N_23531,N_14633,N_16785);
and U23532 (N_23532,N_15367,N_14973);
or U23533 (N_23533,N_14541,N_14631);
nor U23534 (N_23534,N_13649,N_18376);
xnor U23535 (N_23535,N_18357,N_16598);
and U23536 (N_23536,N_14902,N_12677);
xor U23537 (N_23537,N_15009,N_16464);
nor U23538 (N_23538,N_15597,N_14827);
xnor U23539 (N_23539,N_13011,N_13341);
or U23540 (N_23540,N_14002,N_13404);
xnor U23541 (N_23541,N_12800,N_15260);
nand U23542 (N_23542,N_17555,N_13151);
nor U23543 (N_23543,N_16854,N_18542);
nor U23544 (N_23544,N_18260,N_16568);
xnor U23545 (N_23545,N_17024,N_14212);
or U23546 (N_23546,N_16208,N_12844);
xor U23547 (N_23547,N_12526,N_17005);
or U23548 (N_23548,N_14435,N_15165);
or U23549 (N_23549,N_17869,N_18125);
and U23550 (N_23550,N_14553,N_13112);
xnor U23551 (N_23551,N_16739,N_17022);
nand U23552 (N_23552,N_13573,N_12940);
or U23553 (N_23553,N_13498,N_13053);
nand U23554 (N_23554,N_12920,N_14578);
nand U23555 (N_23555,N_14938,N_16944);
nand U23556 (N_23556,N_12569,N_16852);
xnor U23557 (N_23557,N_13908,N_17602);
or U23558 (N_23558,N_14708,N_16860);
nand U23559 (N_23559,N_13598,N_17217);
nand U23560 (N_23560,N_17855,N_13515);
or U23561 (N_23561,N_16198,N_17767);
or U23562 (N_23562,N_15525,N_13672);
xnor U23563 (N_23563,N_17145,N_14515);
nand U23564 (N_23564,N_17032,N_12924);
xnor U23565 (N_23565,N_15695,N_17989);
and U23566 (N_23566,N_17467,N_17839);
xnor U23567 (N_23567,N_14128,N_14245);
nor U23568 (N_23568,N_18573,N_15097);
and U23569 (N_23569,N_16663,N_16913);
nand U23570 (N_23570,N_15002,N_13836);
or U23571 (N_23571,N_18382,N_13634);
or U23572 (N_23572,N_14247,N_16561);
or U23573 (N_23573,N_15684,N_14046);
xnor U23574 (N_23574,N_17656,N_17311);
and U23575 (N_23575,N_16663,N_13899);
nand U23576 (N_23576,N_16463,N_17830);
nand U23577 (N_23577,N_16433,N_14738);
xor U23578 (N_23578,N_13217,N_17467);
or U23579 (N_23579,N_15258,N_16078);
and U23580 (N_23580,N_15232,N_12999);
and U23581 (N_23581,N_12569,N_14982);
xor U23582 (N_23582,N_13901,N_17625);
and U23583 (N_23583,N_14070,N_15407);
xnor U23584 (N_23584,N_14310,N_18712);
or U23585 (N_23585,N_14637,N_18340);
nor U23586 (N_23586,N_13845,N_15039);
and U23587 (N_23587,N_13056,N_15585);
and U23588 (N_23588,N_15512,N_15883);
or U23589 (N_23589,N_15922,N_18000);
xor U23590 (N_23590,N_16349,N_15588);
nor U23591 (N_23591,N_18283,N_17370);
or U23592 (N_23592,N_15616,N_17090);
xor U23593 (N_23593,N_17428,N_15358);
nand U23594 (N_23594,N_15758,N_18335);
xor U23595 (N_23595,N_18511,N_12944);
and U23596 (N_23596,N_13812,N_17407);
xor U23597 (N_23597,N_12509,N_15914);
nand U23598 (N_23598,N_16058,N_18438);
and U23599 (N_23599,N_14166,N_12985);
and U23600 (N_23600,N_16407,N_12890);
nand U23601 (N_23601,N_14952,N_15806);
or U23602 (N_23602,N_13754,N_15756);
and U23603 (N_23603,N_13306,N_17735);
nor U23604 (N_23604,N_18718,N_15192);
nand U23605 (N_23605,N_17253,N_17567);
nor U23606 (N_23606,N_14648,N_13656);
nor U23607 (N_23607,N_15693,N_13939);
and U23608 (N_23608,N_17786,N_15919);
xor U23609 (N_23609,N_14230,N_15484);
and U23610 (N_23610,N_17365,N_14977);
nand U23611 (N_23611,N_18418,N_18700);
nand U23612 (N_23612,N_15210,N_16838);
nor U23613 (N_23613,N_14822,N_15501);
or U23614 (N_23614,N_14900,N_18737);
and U23615 (N_23615,N_18112,N_17758);
or U23616 (N_23616,N_13469,N_13785);
xor U23617 (N_23617,N_12625,N_13363);
nand U23618 (N_23618,N_17909,N_16380);
or U23619 (N_23619,N_18600,N_17594);
or U23620 (N_23620,N_12614,N_12721);
nor U23621 (N_23621,N_15465,N_15178);
nand U23622 (N_23622,N_17717,N_13825);
nor U23623 (N_23623,N_13478,N_15103);
or U23624 (N_23624,N_17114,N_18091);
nand U23625 (N_23625,N_14167,N_18165);
nand U23626 (N_23626,N_12734,N_14301);
or U23627 (N_23627,N_17751,N_16486);
xnor U23628 (N_23628,N_14382,N_14676);
and U23629 (N_23629,N_15402,N_17739);
xnor U23630 (N_23630,N_13195,N_13733);
xor U23631 (N_23631,N_16593,N_18313);
or U23632 (N_23632,N_13373,N_16138);
and U23633 (N_23633,N_12730,N_14913);
xnor U23634 (N_23634,N_14023,N_18238);
nand U23635 (N_23635,N_13747,N_17841);
xor U23636 (N_23636,N_17148,N_15809);
nand U23637 (N_23637,N_15814,N_16557);
nand U23638 (N_23638,N_14159,N_15566);
or U23639 (N_23639,N_18734,N_17271);
nor U23640 (N_23640,N_15325,N_13594);
nor U23641 (N_23641,N_17017,N_13804);
nor U23642 (N_23642,N_12959,N_16116);
xnor U23643 (N_23643,N_17110,N_17060);
nand U23644 (N_23644,N_16356,N_15716);
nand U23645 (N_23645,N_13833,N_15416);
nand U23646 (N_23646,N_12536,N_17107);
and U23647 (N_23647,N_17352,N_16402);
nor U23648 (N_23648,N_18081,N_16838);
nor U23649 (N_23649,N_17538,N_18248);
nor U23650 (N_23650,N_18306,N_14221);
nor U23651 (N_23651,N_18387,N_16404);
xnor U23652 (N_23652,N_18411,N_15253);
nor U23653 (N_23653,N_14930,N_18166);
or U23654 (N_23654,N_13151,N_12557);
or U23655 (N_23655,N_16368,N_16588);
or U23656 (N_23656,N_17714,N_14532);
or U23657 (N_23657,N_18379,N_14735);
nor U23658 (N_23658,N_13984,N_17050);
nand U23659 (N_23659,N_16593,N_14944);
or U23660 (N_23660,N_15953,N_15128);
and U23661 (N_23661,N_12624,N_18030);
nor U23662 (N_23662,N_16112,N_18741);
nor U23663 (N_23663,N_14334,N_17133);
nand U23664 (N_23664,N_14850,N_13993);
xor U23665 (N_23665,N_17359,N_15975);
and U23666 (N_23666,N_17308,N_15111);
or U23667 (N_23667,N_14535,N_16056);
and U23668 (N_23668,N_16121,N_13537);
and U23669 (N_23669,N_15320,N_14329);
xor U23670 (N_23670,N_15414,N_17703);
nand U23671 (N_23671,N_16813,N_14124);
and U23672 (N_23672,N_18557,N_15499);
and U23673 (N_23673,N_15803,N_15397);
and U23674 (N_23674,N_17860,N_15368);
xor U23675 (N_23675,N_17221,N_13030);
xor U23676 (N_23676,N_17115,N_17792);
and U23677 (N_23677,N_17058,N_16573);
and U23678 (N_23678,N_16212,N_18273);
nor U23679 (N_23679,N_14500,N_12576);
xnor U23680 (N_23680,N_18519,N_13787);
and U23681 (N_23681,N_13828,N_15206);
nand U23682 (N_23682,N_17931,N_12751);
and U23683 (N_23683,N_13536,N_14504);
and U23684 (N_23684,N_14423,N_14843);
xnor U23685 (N_23685,N_16939,N_17281);
nand U23686 (N_23686,N_17652,N_16728);
or U23687 (N_23687,N_14872,N_14776);
and U23688 (N_23688,N_13496,N_14911);
and U23689 (N_23689,N_13499,N_14826);
nor U23690 (N_23690,N_16810,N_15893);
nor U23691 (N_23691,N_13316,N_13543);
and U23692 (N_23692,N_12886,N_14144);
and U23693 (N_23693,N_16142,N_15557);
or U23694 (N_23694,N_15053,N_18573);
nand U23695 (N_23695,N_14774,N_12978);
nand U23696 (N_23696,N_14769,N_12708);
and U23697 (N_23697,N_14401,N_12790);
and U23698 (N_23698,N_17492,N_17403);
and U23699 (N_23699,N_17834,N_15264);
nand U23700 (N_23700,N_13092,N_18417);
nand U23701 (N_23701,N_14917,N_18277);
or U23702 (N_23702,N_13164,N_13240);
and U23703 (N_23703,N_17235,N_18521);
and U23704 (N_23704,N_13041,N_17894);
xor U23705 (N_23705,N_16101,N_17895);
or U23706 (N_23706,N_15933,N_16122);
or U23707 (N_23707,N_13309,N_18565);
and U23708 (N_23708,N_17269,N_17075);
and U23709 (N_23709,N_12912,N_16749);
and U23710 (N_23710,N_13315,N_15539);
or U23711 (N_23711,N_16321,N_18291);
xnor U23712 (N_23712,N_15228,N_17482);
nand U23713 (N_23713,N_17259,N_14976);
xor U23714 (N_23714,N_14603,N_16141);
and U23715 (N_23715,N_12650,N_12953);
or U23716 (N_23716,N_13827,N_18066);
or U23717 (N_23717,N_18032,N_16710);
or U23718 (N_23718,N_16270,N_15398);
nor U23719 (N_23719,N_17449,N_13759);
xnor U23720 (N_23720,N_14585,N_16706);
xor U23721 (N_23721,N_14447,N_14475);
or U23722 (N_23722,N_12567,N_14424);
nand U23723 (N_23723,N_14506,N_17064);
and U23724 (N_23724,N_13695,N_16180);
or U23725 (N_23725,N_13405,N_15300);
or U23726 (N_23726,N_14301,N_13380);
or U23727 (N_23727,N_17673,N_13649);
and U23728 (N_23728,N_15065,N_12920);
xnor U23729 (N_23729,N_15889,N_17378);
or U23730 (N_23730,N_16576,N_14762);
or U23731 (N_23731,N_17389,N_14831);
nand U23732 (N_23732,N_14378,N_16543);
and U23733 (N_23733,N_14249,N_13242);
and U23734 (N_23734,N_15367,N_17321);
xor U23735 (N_23735,N_15354,N_14816);
or U23736 (N_23736,N_18003,N_16740);
or U23737 (N_23737,N_17562,N_16218);
nand U23738 (N_23738,N_16802,N_14896);
nor U23739 (N_23739,N_16725,N_14569);
and U23740 (N_23740,N_14651,N_17137);
and U23741 (N_23741,N_14336,N_15087);
and U23742 (N_23742,N_16222,N_16214);
or U23743 (N_23743,N_17521,N_12597);
and U23744 (N_23744,N_12992,N_17326);
and U23745 (N_23745,N_14491,N_15262);
nor U23746 (N_23746,N_18535,N_13699);
or U23747 (N_23747,N_18594,N_14553);
and U23748 (N_23748,N_15769,N_17737);
xnor U23749 (N_23749,N_16895,N_18725);
nand U23750 (N_23750,N_13465,N_12973);
nor U23751 (N_23751,N_18683,N_18531);
and U23752 (N_23752,N_13479,N_18533);
nand U23753 (N_23753,N_14003,N_13080);
nand U23754 (N_23754,N_18110,N_18058);
or U23755 (N_23755,N_13877,N_14465);
and U23756 (N_23756,N_13503,N_15831);
and U23757 (N_23757,N_14583,N_12928);
or U23758 (N_23758,N_18062,N_12775);
or U23759 (N_23759,N_16106,N_18462);
xor U23760 (N_23760,N_14241,N_12547);
nand U23761 (N_23761,N_12853,N_17130);
and U23762 (N_23762,N_17411,N_17615);
nor U23763 (N_23763,N_16123,N_13807);
nand U23764 (N_23764,N_16883,N_15609);
nand U23765 (N_23765,N_13486,N_13353);
xnor U23766 (N_23766,N_16653,N_18320);
nand U23767 (N_23767,N_18390,N_17152);
nand U23768 (N_23768,N_12713,N_13438);
nand U23769 (N_23769,N_14222,N_17696);
and U23770 (N_23770,N_14756,N_13707);
xnor U23771 (N_23771,N_16610,N_16222);
nor U23772 (N_23772,N_15383,N_15032);
xor U23773 (N_23773,N_16745,N_15505);
nand U23774 (N_23774,N_12928,N_13244);
or U23775 (N_23775,N_18694,N_17669);
nor U23776 (N_23776,N_14763,N_17224);
and U23777 (N_23777,N_13027,N_17639);
nand U23778 (N_23778,N_14849,N_16544);
nand U23779 (N_23779,N_16612,N_16784);
nand U23780 (N_23780,N_14016,N_17368);
xnor U23781 (N_23781,N_13711,N_14103);
or U23782 (N_23782,N_16108,N_14136);
xor U23783 (N_23783,N_16482,N_13524);
xor U23784 (N_23784,N_18483,N_13414);
xor U23785 (N_23785,N_14555,N_18289);
nor U23786 (N_23786,N_16336,N_17287);
or U23787 (N_23787,N_15520,N_13838);
nor U23788 (N_23788,N_12645,N_13572);
nor U23789 (N_23789,N_14856,N_13881);
and U23790 (N_23790,N_16092,N_17443);
xor U23791 (N_23791,N_12628,N_17416);
and U23792 (N_23792,N_14465,N_15642);
xnor U23793 (N_23793,N_13849,N_12513);
or U23794 (N_23794,N_12692,N_15244);
and U23795 (N_23795,N_18631,N_13028);
nor U23796 (N_23796,N_14077,N_16330);
nor U23797 (N_23797,N_16120,N_13990);
or U23798 (N_23798,N_13148,N_17859);
xnor U23799 (N_23799,N_18698,N_16010);
and U23800 (N_23800,N_14879,N_14598);
and U23801 (N_23801,N_18649,N_13942);
or U23802 (N_23802,N_14875,N_14238);
or U23803 (N_23803,N_14608,N_18103);
nor U23804 (N_23804,N_12775,N_13159);
nand U23805 (N_23805,N_14798,N_12700);
xnor U23806 (N_23806,N_15079,N_16431);
and U23807 (N_23807,N_17708,N_17901);
nor U23808 (N_23808,N_14326,N_15689);
nand U23809 (N_23809,N_16654,N_14259);
nand U23810 (N_23810,N_16175,N_17376);
xor U23811 (N_23811,N_18082,N_17434);
xor U23812 (N_23812,N_15046,N_12829);
or U23813 (N_23813,N_17961,N_15524);
nand U23814 (N_23814,N_16726,N_15309);
nand U23815 (N_23815,N_18228,N_16632);
nand U23816 (N_23816,N_14252,N_17072);
nand U23817 (N_23817,N_15862,N_14946);
nand U23818 (N_23818,N_17262,N_15023);
or U23819 (N_23819,N_16109,N_12798);
and U23820 (N_23820,N_16236,N_12539);
nor U23821 (N_23821,N_17522,N_16007);
xnor U23822 (N_23822,N_13182,N_16586);
nor U23823 (N_23823,N_18211,N_17421);
or U23824 (N_23824,N_12815,N_15700);
or U23825 (N_23825,N_15899,N_12941);
nor U23826 (N_23826,N_17545,N_16307);
and U23827 (N_23827,N_15959,N_15068);
nor U23828 (N_23828,N_17971,N_17545);
nor U23829 (N_23829,N_16195,N_15113);
or U23830 (N_23830,N_14291,N_14697);
nor U23831 (N_23831,N_14759,N_13267);
or U23832 (N_23832,N_15463,N_18748);
nor U23833 (N_23833,N_14526,N_12956);
xor U23834 (N_23834,N_15574,N_16724);
or U23835 (N_23835,N_13945,N_13579);
and U23836 (N_23836,N_16835,N_14298);
or U23837 (N_23837,N_17477,N_14548);
nand U23838 (N_23838,N_17630,N_14092);
nor U23839 (N_23839,N_17284,N_16773);
nor U23840 (N_23840,N_14530,N_18250);
nor U23841 (N_23841,N_18314,N_15032);
or U23842 (N_23842,N_18296,N_12771);
xor U23843 (N_23843,N_14868,N_17619);
nor U23844 (N_23844,N_17969,N_15654);
xnor U23845 (N_23845,N_15129,N_14723);
xnor U23846 (N_23846,N_14611,N_18258);
or U23847 (N_23847,N_12789,N_14839);
nand U23848 (N_23848,N_14858,N_13710);
xnor U23849 (N_23849,N_17924,N_13008);
xor U23850 (N_23850,N_13987,N_16344);
nand U23851 (N_23851,N_13436,N_14225);
xnor U23852 (N_23852,N_14929,N_17698);
and U23853 (N_23853,N_13368,N_14045);
or U23854 (N_23854,N_15127,N_12796);
nand U23855 (N_23855,N_15542,N_16739);
nor U23856 (N_23856,N_15298,N_13171);
xor U23857 (N_23857,N_17438,N_14252);
or U23858 (N_23858,N_15810,N_16669);
nor U23859 (N_23859,N_12669,N_16091);
or U23860 (N_23860,N_14588,N_14268);
nor U23861 (N_23861,N_14827,N_17972);
or U23862 (N_23862,N_17824,N_16269);
nor U23863 (N_23863,N_15252,N_17431);
nand U23864 (N_23864,N_14224,N_14573);
nor U23865 (N_23865,N_14886,N_15325);
or U23866 (N_23866,N_15824,N_17942);
nor U23867 (N_23867,N_14064,N_15100);
and U23868 (N_23868,N_13578,N_14600);
nand U23869 (N_23869,N_13240,N_16690);
nand U23870 (N_23870,N_14343,N_14902);
and U23871 (N_23871,N_13620,N_17294);
nor U23872 (N_23872,N_16989,N_15022);
nand U23873 (N_23873,N_18456,N_13455);
xor U23874 (N_23874,N_15394,N_13523);
and U23875 (N_23875,N_13024,N_17801);
nor U23876 (N_23876,N_17694,N_15980);
xnor U23877 (N_23877,N_14956,N_18649);
nor U23878 (N_23878,N_17255,N_12750);
and U23879 (N_23879,N_13023,N_17868);
nor U23880 (N_23880,N_15278,N_18510);
nand U23881 (N_23881,N_15876,N_18277);
or U23882 (N_23882,N_12622,N_17327);
nor U23883 (N_23883,N_16896,N_14086);
nor U23884 (N_23884,N_18455,N_17452);
nor U23885 (N_23885,N_17503,N_13602);
nand U23886 (N_23886,N_18493,N_17028);
nand U23887 (N_23887,N_17756,N_13518);
or U23888 (N_23888,N_12792,N_13916);
nand U23889 (N_23889,N_18239,N_14927);
and U23890 (N_23890,N_13820,N_14081);
xnor U23891 (N_23891,N_12924,N_13354);
nand U23892 (N_23892,N_16627,N_15949);
nand U23893 (N_23893,N_17100,N_12978);
nor U23894 (N_23894,N_17135,N_17593);
and U23895 (N_23895,N_16841,N_14346);
nor U23896 (N_23896,N_14027,N_16972);
nand U23897 (N_23897,N_17327,N_15880);
nor U23898 (N_23898,N_18415,N_17742);
nand U23899 (N_23899,N_15494,N_18626);
nand U23900 (N_23900,N_12637,N_16262);
nand U23901 (N_23901,N_14182,N_15592);
and U23902 (N_23902,N_16368,N_16223);
and U23903 (N_23903,N_13515,N_17026);
nor U23904 (N_23904,N_16003,N_17418);
or U23905 (N_23905,N_18127,N_16718);
xor U23906 (N_23906,N_15033,N_14065);
or U23907 (N_23907,N_13661,N_18037);
nor U23908 (N_23908,N_17215,N_15970);
nor U23909 (N_23909,N_14517,N_16939);
or U23910 (N_23910,N_15369,N_17113);
xor U23911 (N_23911,N_14045,N_13198);
nand U23912 (N_23912,N_18747,N_14592);
nor U23913 (N_23913,N_18132,N_15511);
nor U23914 (N_23914,N_16850,N_13449);
nor U23915 (N_23915,N_12643,N_16552);
xnor U23916 (N_23916,N_13412,N_16210);
nor U23917 (N_23917,N_18734,N_12950);
and U23918 (N_23918,N_13939,N_12821);
and U23919 (N_23919,N_13575,N_15512);
nor U23920 (N_23920,N_13649,N_13876);
nand U23921 (N_23921,N_13693,N_12783);
nand U23922 (N_23922,N_15564,N_13031);
nor U23923 (N_23923,N_15449,N_13568);
nand U23924 (N_23924,N_17451,N_15080);
and U23925 (N_23925,N_17948,N_14635);
xnor U23926 (N_23926,N_13644,N_13680);
and U23927 (N_23927,N_15964,N_15196);
nor U23928 (N_23928,N_17455,N_13932);
or U23929 (N_23929,N_15312,N_16458);
nor U23930 (N_23930,N_18556,N_16189);
nor U23931 (N_23931,N_17351,N_17090);
nor U23932 (N_23932,N_17992,N_12616);
nor U23933 (N_23933,N_17226,N_18555);
nor U23934 (N_23934,N_16789,N_16551);
nand U23935 (N_23935,N_12687,N_17730);
xnor U23936 (N_23936,N_13254,N_14631);
nand U23937 (N_23937,N_14026,N_13915);
xor U23938 (N_23938,N_17747,N_16559);
nor U23939 (N_23939,N_18325,N_13780);
or U23940 (N_23940,N_14582,N_15343);
or U23941 (N_23941,N_17877,N_17665);
or U23942 (N_23942,N_12718,N_18039);
nor U23943 (N_23943,N_17605,N_13793);
nor U23944 (N_23944,N_14462,N_17644);
nand U23945 (N_23945,N_17728,N_15003);
or U23946 (N_23946,N_13892,N_17094);
and U23947 (N_23947,N_13853,N_13121);
and U23948 (N_23948,N_15642,N_18405);
or U23949 (N_23949,N_14020,N_13994);
xnor U23950 (N_23950,N_15187,N_16566);
and U23951 (N_23951,N_14787,N_16845);
and U23952 (N_23952,N_18169,N_13479);
nor U23953 (N_23953,N_15701,N_18085);
or U23954 (N_23954,N_15356,N_13062);
nor U23955 (N_23955,N_14820,N_15462);
xor U23956 (N_23956,N_16209,N_15654);
nor U23957 (N_23957,N_14525,N_14096);
nand U23958 (N_23958,N_16219,N_15817);
xnor U23959 (N_23959,N_12714,N_16772);
xnor U23960 (N_23960,N_17895,N_15237);
and U23961 (N_23961,N_12993,N_13006);
and U23962 (N_23962,N_16456,N_14314);
xor U23963 (N_23963,N_16326,N_15317);
and U23964 (N_23964,N_15048,N_14920);
nor U23965 (N_23965,N_13368,N_13669);
and U23966 (N_23966,N_13665,N_18504);
or U23967 (N_23967,N_16051,N_17371);
nor U23968 (N_23968,N_16115,N_14840);
nor U23969 (N_23969,N_16230,N_12852);
and U23970 (N_23970,N_14438,N_14442);
or U23971 (N_23971,N_14359,N_15034);
or U23972 (N_23972,N_18315,N_16398);
and U23973 (N_23973,N_18245,N_15905);
xnor U23974 (N_23974,N_12819,N_13930);
and U23975 (N_23975,N_12919,N_13511);
nor U23976 (N_23976,N_12936,N_16120);
xor U23977 (N_23977,N_18517,N_13912);
and U23978 (N_23978,N_15890,N_18636);
xor U23979 (N_23979,N_14328,N_16785);
or U23980 (N_23980,N_18066,N_14675);
nor U23981 (N_23981,N_13212,N_14948);
nand U23982 (N_23982,N_12512,N_14731);
nand U23983 (N_23983,N_16132,N_15480);
nand U23984 (N_23984,N_12559,N_17917);
and U23985 (N_23985,N_13142,N_17067);
nand U23986 (N_23986,N_17412,N_12913);
xnor U23987 (N_23987,N_12546,N_17936);
xnor U23988 (N_23988,N_13174,N_15378);
nand U23989 (N_23989,N_15387,N_15593);
xor U23990 (N_23990,N_16714,N_16013);
nand U23991 (N_23991,N_15435,N_16887);
and U23992 (N_23992,N_18463,N_18070);
or U23993 (N_23993,N_13776,N_18049);
and U23994 (N_23994,N_12681,N_17427);
and U23995 (N_23995,N_13113,N_13186);
nand U23996 (N_23996,N_13263,N_12861);
nor U23997 (N_23997,N_18435,N_18091);
nor U23998 (N_23998,N_15968,N_18303);
nor U23999 (N_23999,N_17453,N_18069);
nor U24000 (N_24000,N_13460,N_12570);
nand U24001 (N_24001,N_16581,N_17345);
and U24002 (N_24002,N_16051,N_13477);
xor U24003 (N_24003,N_18135,N_13879);
nor U24004 (N_24004,N_15815,N_15096);
or U24005 (N_24005,N_15095,N_14530);
xnor U24006 (N_24006,N_18190,N_14445);
or U24007 (N_24007,N_16605,N_13770);
and U24008 (N_24008,N_14428,N_14632);
nand U24009 (N_24009,N_13630,N_16515);
and U24010 (N_24010,N_13635,N_16731);
xor U24011 (N_24011,N_16133,N_13882);
xor U24012 (N_24012,N_14373,N_12931);
and U24013 (N_24013,N_17216,N_15186);
or U24014 (N_24014,N_14788,N_12687);
nand U24015 (N_24015,N_17732,N_18226);
nor U24016 (N_24016,N_17495,N_16287);
and U24017 (N_24017,N_14529,N_14281);
and U24018 (N_24018,N_16193,N_16007);
nor U24019 (N_24019,N_18440,N_13585);
xor U24020 (N_24020,N_15811,N_13154);
nand U24021 (N_24021,N_17285,N_18211);
or U24022 (N_24022,N_16390,N_13537);
nor U24023 (N_24023,N_14379,N_17583);
nand U24024 (N_24024,N_17877,N_17438);
and U24025 (N_24025,N_14128,N_17585);
xor U24026 (N_24026,N_18145,N_17366);
and U24027 (N_24027,N_14227,N_17873);
and U24028 (N_24028,N_17991,N_17181);
nand U24029 (N_24029,N_12931,N_14920);
and U24030 (N_24030,N_12555,N_16494);
or U24031 (N_24031,N_17437,N_17135);
nor U24032 (N_24032,N_18651,N_13381);
and U24033 (N_24033,N_16941,N_14346);
nor U24034 (N_24034,N_12925,N_15502);
nor U24035 (N_24035,N_18271,N_14799);
and U24036 (N_24036,N_14579,N_17857);
or U24037 (N_24037,N_15702,N_18680);
nor U24038 (N_24038,N_15945,N_13880);
nor U24039 (N_24039,N_13309,N_16283);
and U24040 (N_24040,N_17511,N_15248);
and U24041 (N_24041,N_16922,N_14032);
nand U24042 (N_24042,N_14822,N_12674);
and U24043 (N_24043,N_17633,N_13525);
and U24044 (N_24044,N_13761,N_15960);
nor U24045 (N_24045,N_16460,N_14597);
nand U24046 (N_24046,N_14366,N_17455);
xnor U24047 (N_24047,N_13270,N_15261);
and U24048 (N_24048,N_12629,N_14839);
nor U24049 (N_24049,N_14154,N_16280);
and U24050 (N_24050,N_16669,N_17870);
nor U24051 (N_24051,N_16595,N_17216);
xnor U24052 (N_24052,N_13648,N_13244);
xor U24053 (N_24053,N_16323,N_15096);
or U24054 (N_24054,N_15842,N_13352);
and U24055 (N_24055,N_15236,N_14198);
or U24056 (N_24056,N_15773,N_16544);
nor U24057 (N_24057,N_15015,N_14820);
xor U24058 (N_24058,N_16706,N_18138);
xor U24059 (N_24059,N_14770,N_18410);
or U24060 (N_24060,N_16750,N_16541);
or U24061 (N_24061,N_16230,N_13366);
or U24062 (N_24062,N_16716,N_18598);
and U24063 (N_24063,N_12687,N_16376);
or U24064 (N_24064,N_15014,N_16706);
and U24065 (N_24065,N_17766,N_18189);
and U24066 (N_24066,N_14701,N_13633);
nor U24067 (N_24067,N_18291,N_16996);
xor U24068 (N_24068,N_16399,N_16680);
and U24069 (N_24069,N_13758,N_13060);
and U24070 (N_24070,N_12563,N_14694);
xnor U24071 (N_24071,N_12511,N_15127);
xnor U24072 (N_24072,N_13058,N_14335);
or U24073 (N_24073,N_13793,N_16943);
nand U24074 (N_24074,N_16640,N_15548);
nand U24075 (N_24075,N_14661,N_15483);
nand U24076 (N_24076,N_15182,N_17485);
nor U24077 (N_24077,N_17369,N_12716);
and U24078 (N_24078,N_15789,N_17037);
and U24079 (N_24079,N_16668,N_17371);
nand U24080 (N_24080,N_17952,N_13150);
and U24081 (N_24081,N_14588,N_13356);
or U24082 (N_24082,N_13323,N_14400);
and U24083 (N_24083,N_12624,N_16409);
or U24084 (N_24084,N_16367,N_15591);
nand U24085 (N_24085,N_12918,N_14718);
or U24086 (N_24086,N_18323,N_15955);
or U24087 (N_24087,N_18339,N_14281);
nand U24088 (N_24088,N_18240,N_17386);
xnor U24089 (N_24089,N_14961,N_12685);
nor U24090 (N_24090,N_12840,N_18172);
nor U24091 (N_24091,N_18139,N_13410);
or U24092 (N_24092,N_18699,N_15565);
or U24093 (N_24093,N_16051,N_16795);
nor U24094 (N_24094,N_12631,N_13604);
nand U24095 (N_24095,N_16912,N_12829);
and U24096 (N_24096,N_15784,N_17414);
nand U24097 (N_24097,N_15473,N_14438);
or U24098 (N_24098,N_16605,N_16051);
or U24099 (N_24099,N_17349,N_15266);
or U24100 (N_24100,N_12719,N_15469);
xnor U24101 (N_24101,N_16321,N_14023);
xor U24102 (N_24102,N_14889,N_15605);
nand U24103 (N_24103,N_15075,N_13286);
nor U24104 (N_24104,N_13132,N_16751);
and U24105 (N_24105,N_17085,N_18652);
and U24106 (N_24106,N_13477,N_18638);
nor U24107 (N_24107,N_13274,N_14599);
nand U24108 (N_24108,N_18376,N_17379);
nor U24109 (N_24109,N_13442,N_14220);
or U24110 (N_24110,N_12741,N_18158);
nand U24111 (N_24111,N_18688,N_13306);
nand U24112 (N_24112,N_14936,N_13171);
nand U24113 (N_24113,N_17401,N_15996);
nand U24114 (N_24114,N_12918,N_13136);
and U24115 (N_24115,N_12822,N_15116);
xor U24116 (N_24116,N_18625,N_15482);
and U24117 (N_24117,N_17650,N_12924);
xnor U24118 (N_24118,N_15070,N_15590);
and U24119 (N_24119,N_17047,N_15427);
nand U24120 (N_24120,N_13812,N_17074);
or U24121 (N_24121,N_17112,N_13530);
and U24122 (N_24122,N_17859,N_14261);
xnor U24123 (N_24123,N_17321,N_16452);
xnor U24124 (N_24124,N_16189,N_13514);
and U24125 (N_24125,N_16004,N_15537);
nand U24126 (N_24126,N_15797,N_14148);
xnor U24127 (N_24127,N_13104,N_13884);
and U24128 (N_24128,N_15269,N_14581);
nor U24129 (N_24129,N_15058,N_14208);
or U24130 (N_24130,N_15595,N_13073);
or U24131 (N_24131,N_17507,N_16713);
nor U24132 (N_24132,N_12997,N_14796);
or U24133 (N_24133,N_13303,N_16047);
or U24134 (N_24134,N_14909,N_16566);
or U24135 (N_24135,N_17647,N_12540);
xnor U24136 (N_24136,N_18027,N_15847);
xnor U24137 (N_24137,N_12569,N_13921);
nor U24138 (N_24138,N_14728,N_15542);
nor U24139 (N_24139,N_17147,N_13355);
nand U24140 (N_24140,N_15186,N_13773);
nand U24141 (N_24141,N_13922,N_16195);
or U24142 (N_24142,N_14082,N_17688);
xnor U24143 (N_24143,N_16722,N_16321);
nand U24144 (N_24144,N_14205,N_14963);
xnor U24145 (N_24145,N_17452,N_16772);
nand U24146 (N_24146,N_13755,N_14724);
xnor U24147 (N_24147,N_13143,N_16365);
nor U24148 (N_24148,N_16371,N_15364);
nand U24149 (N_24149,N_18167,N_17007);
nor U24150 (N_24150,N_17666,N_17034);
nor U24151 (N_24151,N_15829,N_15873);
and U24152 (N_24152,N_16449,N_16078);
nand U24153 (N_24153,N_16805,N_14536);
and U24154 (N_24154,N_15023,N_13750);
nor U24155 (N_24155,N_15371,N_14233);
xnor U24156 (N_24156,N_13006,N_16229);
or U24157 (N_24157,N_15294,N_13531);
nor U24158 (N_24158,N_14687,N_15345);
nand U24159 (N_24159,N_14675,N_18311);
nor U24160 (N_24160,N_15057,N_14906);
or U24161 (N_24161,N_17016,N_16908);
and U24162 (N_24162,N_14030,N_13153);
and U24163 (N_24163,N_18672,N_13142);
nor U24164 (N_24164,N_15332,N_18489);
or U24165 (N_24165,N_13119,N_12625);
nor U24166 (N_24166,N_17824,N_18505);
nand U24167 (N_24167,N_14740,N_15539);
or U24168 (N_24168,N_18012,N_14727);
xnor U24169 (N_24169,N_15048,N_13813);
nor U24170 (N_24170,N_16626,N_13864);
and U24171 (N_24171,N_16251,N_18067);
or U24172 (N_24172,N_14141,N_13112);
nor U24173 (N_24173,N_17129,N_16640);
and U24174 (N_24174,N_18049,N_13813);
xnor U24175 (N_24175,N_18615,N_16258);
nand U24176 (N_24176,N_13837,N_13468);
and U24177 (N_24177,N_15578,N_16706);
nand U24178 (N_24178,N_17947,N_16481);
nand U24179 (N_24179,N_18482,N_14821);
or U24180 (N_24180,N_14907,N_17645);
or U24181 (N_24181,N_12723,N_17532);
nand U24182 (N_24182,N_15355,N_16358);
nand U24183 (N_24183,N_14416,N_18497);
xor U24184 (N_24184,N_16929,N_16575);
or U24185 (N_24185,N_16094,N_16145);
nor U24186 (N_24186,N_16380,N_13844);
or U24187 (N_24187,N_16052,N_12668);
nor U24188 (N_24188,N_15482,N_17054);
nand U24189 (N_24189,N_18123,N_12556);
or U24190 (N_24190,N_15637,N_13817);
and U24191 (N_24191,N_12997,N_15553);
nor U24192 (N_24192,N_13571,N_14797);
xor U24193 (N_24193,N_12791,N_13527);
nor U24194 (N_24194,N_17087,N_17489);
nor U24195 (N_24195,N_14126,N_16599);
xor U24196 (N_24196,N_17821,N_13571);
nor U24197 (N_24197,N_14749,N_15194);
xnor U24198 (N_24198,N_15672,N_18237);
xor U24199 (N_24199,N_16426,N_15159);
and U24200 (N_24200,N_14844,N_14682);
nand U24201 (N_24201,N_16466,N_17262);
nand U24202 (N_24202,N_17145,N_16061);
nand U24203 (N_24203,N_14782,N_16896);
and U24204 (N_24204,N_14514,N_16277);
nor U24205 (N_24205,N_15363,N_16128);
xor U24206 (N_24206,N_18418,N_18709);
and U24207 (N_24207,N_13688,N_14500);
xor U24208 (N_24208,N_18437,N_15188);
nand U24209 (N_24209,N_15216,N_17792);
and U24210 (N_24210,N_13271,N_15301);
nand U24211 (N_24211,N_14280,N_12878);
or U24212 (N_24212,N_17426,N_15276);
nand U24213 (N_24213,N_12984,N_16305);
nor U24214 (N_24214,N_13163,N_14890);
or U24215 (N_24215,N_13053,N_17196);
or U24216 (N_24216,N_13291,N_13464);
xor U24217 (N_24217,N_16877,N_13578);
and U24218 (N_24218,N_16761,N_14730);
nand U24219 (N_24219,N_12557,N_18688);
xnor U24220 (N_24220,N_17050,N_14172);
and U24221 (N_24221,N_17937,N_13514);
or U24222 (N_24222,N_18048,N_16444);
or U24223 (N_24223,N_13353,N_12677);
xnor U24224 (N_24224,N_16002,N_13529);
nor U24225 (N_24225,N_15786,N_13374);
xnor U24226 (N_24226,N_17355,N_16442);
xor U24227 (N_24227,N_17908,N_15422);
nand U24228 (N_24228,N_12570,N_13128);
nor U24229 (N_24229,N_12754,N_16101);
xnor U24230 (N_24230,N_16308,N_16861);
nor U24231 (N_24231,N_13659,N_15532);
and U24232 (N_24232,N_16661,N_12616);
nor U24233 (N_24233,N_13285,N_14614);
and U24234 (N_24234,N_13758,N_15448);
nor U24235 (N_24235,N_13799,N_17948);
nor U24236 (N_24236,N_17162,N_17659);
nand U24237 (N_24237,N_13276,N_15596);
xor U24238 (N_24238,N_15550,N_17646);
or U24239 (N_24239,N_12582,N_15964);
nor U24240 (N_24240,N_13923,N_12667);
or U24241 (N_24241,N_18626,N_17876);
or U24242 (N_24242,N_16402,N_13236);
nor U24243 (N_24243,N_12632,N_14551);
or U24244 (N_24244,N_15283,N_17495);
nor U24245 (N_24245,N_18124,N_12868);
nand U24246 (N_24246,N_17060,N_15999);
xnor U24247 (N_24247,N_17377,N_18583);
nor U24248 (N_24248,N_17039,N_13664);
xor U24249 (N_24249,N_13870,N_14187);
and U24250 (N_24250,N_13386,N_17033);
nand U24251 (N_24251,N_18247,N_15043);
xnor U24252 (N_24252,N_13887,N_13634);
xor U24253 (N_24253,N_15935,N_17179);
or U24254 (N_24254,N_14716,N_18434);
or U24255 (N_24255,N_18023,N_15924);
xor U24256 (N_24256,N_13628,N_17839);
nand U24257 (N_24257,N_14418,N_16024);
and U24258 (N_24258,N_16530,N_16851);
nor U24259 (N_24259,N_14629,N_14341);
nand U24260 (N_24260,N_18171,N_12976);
nor U24261 (N_24261,N_16930,N_17768);
nor U24262 (N_24262,N_16689,N_13465);
or U24263 (N_24263,N_15392,N_16820);
nor U24264 (N_24264,N_15500,N_13733);
xnor U24265 (N_24265,N_12677,N_17700);
or U24266 (N_24266,N_14401,N_17330);
nor U24267 (N_24267,N_15448,N_16370);
nor U24268 (N_24268,N_12705,N_15697);
nand U24269 (N_24269,N_15772,N_12813);
and U24270 (N_24270,N_14189,N_12606);
nor U24271 (N_24271,N_14743,N_15378);
and U24272 (N_24272,N_14405,N_13711);
and U24273 (N_24273,N_16496,N_16633);
and U24274 (N_24274,N_13402,N_13744);
or U24275 (N_24275,N_15154,N_18520);
nor U24276 (N_24276,N_17531,N_16785);
nand U24277 (N_24277,N_18498,N_12565);
nand U24278 (N_24278,N_17012,N_16717);
or U24279 (N_24279,N_12617,N_13243);
and U24280 (N_24280,N_15704,N_15343);
and U24281 (N_24281,N_17509,N_16590);
nor U24282 (N_24282,N_18382,N_14901);
and U24283 (N_24283,N_14876,N_15975);
nand U24284 (N_24284,N_14443,N_12779);
xor U24285 (N_24285,N_15507,N_12947);
nor U24286 (N_24286,N_15276,N_14958);
nor U24287 (N_24287,N_14029,N_15605);
xor U24288 (N_24288,N_14594,N_17974);
and U24289 (N_24289,N_13857,N_16722);
nor U24290 (N_24290,N_17918,N_15763);
xnor U24291 (N_24291,N_13578,N_18346);
xor U24292 (N_24292,N_13486,N_12565);
nand U24293 (N_24293,N_13038,N_18674);
nand U24294 (N_24294,N_16089,N_15585);
and U24295 (N_24295,N_16333,N_17810);
xor U24296 (N_24296,N_16848,N_14380);
xnor U24297 (N_24297,N_17299,N_12662);
or U24298 (N_24298,N_16419,N_14553);
or U24299 (N_24299,N_13272,N_13256);
xnor U24300 (N_24300,N_15606,N_17792);
nand U24301 (N_24301,N_15037,N_12712);
nor U24302 (N_24302,N_12697,N_14428);
or U24303 (N_24303,N_13724,N_18389);
nand U24304 (N_24304,N_15615,N_13549);
or U24305 (N_24305,N_17087,N_13777);
or U24306 (N_24306,N_12831,N_14771);
and U24307 (N_24307,N_16628,N_18202);
and U24308 (N_24308,N_16748,N_16186);
xor U24309 (N_24309,N_12808,N_15971);
nand U24310 (N_24310,N_14751,N_18207);
or U24311 (N_24311,N_16215,N_15747);
or U24312 (N_24312,N_18657,N_15383);
xnor U24313 (N_24313,N_18057,N_16637);
nand U24314 (N_24314,N_16480,N_13470);
nor U24315 (N_24315,N_17861,N_15451);
or U24316 (N_24316,N_13684,N_18108);
xor U24317 (N_24317,N_13780,N_18541);
nand U24318 (N_24318,N_15466,N_13251);
or U24319 (N_24319,N_14249,N_14027);
and U24320 (N_24320,N_13279,N_15336);
xor U24321 (N_24321,N_16708,N_13167);
xor U24322 (N_24322,N_17455,N_18623);
nor U24323 (N_24323,N_15369,N_14182);
nand U24324 (N_24324,N_15489,N_16056);
or U24325 (N_24325,N_13619,N_15743);
nor U24326 (N_24326,N_16558,N_17244);
or U24327 (N_24327,N_15660,N_17308);
nor U24328 (N_24328,N_16431,N_15632);
or U24329 (N_24329,N_13676,N_14578);
nand U24330 (N_24330,N_15673,N_14586);
xnor U24331 (N_24331,N_15479,N_14805);
or U24332 (N_24332,N_18627,N_18007);
xnor U24333 (N_24333,N_15571,N_18188);
and U24334 (N_24334,N_13774,N_16771);
and U24335 (N_24335,N_15737,N_13739);
nand U24336 (N_24336,N_17246,N_18087);
or U24337 (N_24337,N_16492,N_16057);
and U24338 (N_24338,N_17641,N_13717);
nand U24339 (N_24339,N_17202,N_13385);
or U24340 (N_24340,N_14693,N_17887);
xnor U24341 (N_24341,N_13964,N_17759);
and U24342 (N_24342,N_17380,N_17438);
nand U24343 (N_24343,N_13489,N_16553);
or U24344 (N_24344,N_17926,N_17508);
xnor U24345 (N_24345,N_17421,N_12950);
nor U24346 (N_24346,N_17210,N_15373);
and U24347 (N_24347,N_16527,N_13243);
xnor U24348 (N_24348,N_15198,N_13738);
and U24349 (N_24349,N_13982,N_14151);
nor U24350 (N_24350,N_17424,N_15098);
xnor U24351 (N_24351,N_18337,N_16864);
nor U24352 (N_24352,N_14143,N_18144);
or U24353 (N_24353,N_14149,N_12954);
nand U24354 (N_24354,N_13202,N_14056);
xnor U24355 (N_24355,N_15488,N_15031);
xnor U24356 (N_24356,N_13451,N_15264);
or U24357 (N_24357,N_14302,N_13275);
and U24358 (N_24358,N_15170,N_15718);
nor U24359 (N_24359,N_14961,N_16142);
or U24360 (N_24360,N_13668,N_15728);
nand U24361 (N_24361,N_15107,N_13044);
nand U24362 (N_24362,N_17376,N_15148);
and U24363 (N_24363,N_17246,N_15359);
nand U24364 (N_24364,N_14394,N_12584);
or U24365 (N_24365,N_16606,N_18073);
nand U24366 (N_24366,N_15339,N_17614);
nor U24367 (N_24367,N_13889,N_17780);
xor U24368 (N_24368,N_14533,N_17355);
xor U24369 (N_24369,N_18726,N_16207);
xnor U24370 (N_24370,N_16490,N_17446);
nor U24371 (N_24371,N_13574,N_14418);
xnor U24372 (N_24372,N_13930,N_14423);
nand U24373 (N_24373,N_15900,N_16126);
xnor U24374 (N_24374,N_13463,N_16038);
nand U24375 (N_24375,N_13889,N_15371);
or U24376 (N_24376,N_13910,N_15398);
or U24377 (N_24377,N_13270,N_17607);
nor U24378 (N_24378,N_18708,N_17029);
nand U24379 (N_24379,N_13106,N_17413);
nor U24380 (N_24380,N_14794,N_15796);
or U24381 (N_24381,N_16709,N_17152);
and U24382 (N_24382,N_18311,N_17119);
xnor U24383 (N_24383,N_14846,N_14233);
nor U24384 (N_24384,N_13085,N_16455);
nor U24385 (N_24385,N_14079,N_15770);
or U24386 (N_24386,N_18194,N_13292);
nand U24387 (N_24387,N_13629,N_17310);
nand U24388 (N_24388,N_14171,N_18633);
nand U24389 (N_24389,N_16267,N_15695);
nand U24390 (N_24390,N_17561,N_18224);
and U24391 (N_24391,N_12505,N_13721);
nand U24392 (N_24392,N_17451,N_16900);
and U24393 (N_24393,N_13048,N_15646);
and U24394 (N_24394,N_14076,N_13194);
nor U24395 (N_24395,N_15509,N_17686);
nor U24396 (N_24396,N_17220,N_13448);
or U24397 (N_24397,N_16386,N_13829);
nor U24398 (N_24398,N_17073,N_17605);
xnor U24399 (N_24399,N_13517,N_17240);
and U24400 (N_24400,N_17119,N_14021);
or U24401 (N_24401,N_17436,N_15674);
xnor U24402 (N_24402,N_14886,N_13918);
xnor U24403 (N_24403,N_13559,N_18023);
xor U24404 (N_24404,N_14483,N_13828);
xor U24405 (N_24405,N_15091,N_16672);
nand U24406 (N_24406,N_12664,N_14540);
nor U24407 (N_24407,N_14229,N_15527);
nand U24408 (N_24408,N_14291,N_13712);
or U24409 (N_24409,N_16331,N_15437);
nand U24410 (N_24410,N_17433,N_12936);
nor U24411 (N_24411,N_13682,N_12567);
nor U24412 (N_24412,N_13152,N_16527);
and U24413 (N_24413,N_16063,N_18610);
nand U24414 (N_24414,N_16282,N_17112);
and U24415 (N_24415,N_17999,N_14594);
or U24416 (N_24416,N_14199,N_14119);
xnor U24417 (N_24417,N_16163,N_16020);
or U24418 (N_24418,N_16350,N_15052);
or U24419 (N_24419,N_17084,N_13702);
or U24420 (N_24420,N_14341,N_17832);
xnor U24421 (N_24421,N_16778,N_15485);
and U24422 (N_24422,N_14144,N_13991);
or U24423 (N_24423,N_18535,N_16306);
and U24424 (N_24424,N_17924,N_18019);
or U24425 (N_24425,N_16347,N_13262);
nand U24426 (N_24426,N_13109,N_16445);
and U24427 (N_24427,N_13749,N_18154);
xor U24428 (N_24428,N_17004,N_15456);
nand U24429 (N_24429,N_12831,N_17703);
and U24430 (N_24430,N_14140,N_14950);
nand U24431 (N_24431,N_14239,N_12501);
and U24432 (N_24432,N_16343,N_17939);
and U24433 (N_24433,N_15158,N_17928);
xnor U24434 (N_24434,N_17616,N_13740);
or U24435 (N_24435,N_16960,N_14126);
nor U24436 (N_24436,N_16692,N_14637);
and U24437 (N_24437,N_14734,N_13203);
nor U24438 (N_24438,N_13672,N_12795);
xnor U24439 (N_24439,N_16276,N_13096);
nor U24440 (N_24440,N_13511,N_12900);
or U24441 (N_24441,N_13968,N_13993);
and U24442 (N_24442,N_14077,N_14201);
nand U24443 (N_24443,N_13965,N_15982);
or U24444 (N_24444,N_13236,N_17494);
and U24445 (N_24445,N_17299,N_18232);
or U24446 (N_24446,N_14206,N_17585);
or U24447 (N_24447,N_13008,N_16114);
or U24448 (N_24448,N_13988,N_13084);
xor U24449 (N_24449,N_12676,N_13633);
xor U24450 (N_24450,N_13159,N_13214);
xnor U24451 (N_24451,N_16910,N_16710);
nor U24452 (N_24452,N_12683,N_15138);
nand U24453 (N_24453,N_12970,N_17600);
and U24454 (N_24454,N_16024,N_16614);
or U24455 (N_24455,N_17819,N_13724);
and U24456 (N_24456,N_14687,N_18189);
or U24457 (N_24457,N_18570,N_18626);
xnor U24458 (N_24458,N_16569,N_13061);
xor U24459 (N_24459,N_17379,N_16472);
nand U24460 (N_24460,N_14621,N_14206);
nand U24461 (N_24461,N_14353,N_17560);
nor U24462 (N_24462,N_18712,N_15117);
nor U24463 (N_24463,N_13780,N_13215);
xor U24464 (N_24464,N_12821,N_18096);
and U24465 (N_24465,N_17055,N_14926);
nor U24466 (N_24466,N_16837,N_17545);
or U24467 (N_24467,N_17294,N_15491);
or U24468 (N_24468,N_14782,N_12958);
and U24469 (N_24469,N_15629,N_15074);
xnor U24470 (N_24470,N_13561,N_16562);
nand U24471 (N_24471,N_15674,N_18321);
xor U24472 (N_24472,N_17513,N_15557);
xnor U24473 (N_24473,N_17347,N_12820);
and U24474 (N_24474,N_16619,N_13274);
nor U24475 (N_24475,N_18712,N_15226);
xor U24476 (N_24476,N_14683,N_15763);
nand U24477 (N_24477,N_18288,N_15218);
nand U24478 (N_24478,N_16596,N_15120);
or U24479 (N_24479,N_15470,N_13231);
nand U24480 (N_24480,N_15648,N_17252);
xor U24481 (N_24481,N_17494,N_15875);
or U24482 (N_24482,N_17410,N_13532);
nand U24483 (N_24483,N_16640,N_16170);
or U24484 (N_24484,N_15793,N_15261);
and U24485 (N_24485,N_15494,N_17902);
or U24486 (N_24486,N_17227,N_16040);
nand U24487 (N_24487,N_14075,N_16192);
xnor U24488 (N_24488,N_17568,N_12719);
nor U24489 (N_24489,N_17955,N_14313);
nor U24490 (N_24490,N_14489,N_16600);
xnor U24491 (N_24491,N_14855,N_14305);
or U24492 (N_24492,N_15422,N_16990);
or U24493 (N_24493,N_17521,N_18465);
nor U24494 (N_24494,N_13373,N_18216);
and U24495 (N_24495,N_17886,N_15747);
nand U24496 (N_24496,N_15982,N_17242);
and U24497 (N_24497,N_15864,N_15515);
nand U24498 (N_24498,N_15113,N_12669);
or U24499 (N_24499,N_16920,N_12788);
nand U24500 (N_24500,N_13192,N_13613);
nand U24501 (N_24501,N_15474,N_12899);
or U24502 (N_24502,N_16204,N_15607);
nand U24503 (N_24503,N_18353,N_14590);
nor U24504 (N_24504,N_14563,N_12999);
nor U24505 (N_24505,N_13199,N_16051);
nand U24506 (N_24506,N_13180,N_17533);
xnor U24507 (N_24507,N_15216,N_17251);
or U24508 (N_24508,N_16466,N_17170);
nand U24509 (N_24509,N_14105,N_13251);
nand U24510 (N_24510,N_15620,N_15266);
nor U24511 (N_24511,N_12721,N_18338);
nor U24512 (N_24512,N_17041,N_18433);
and U24513 (N_24513,N_18399,N_13429);
nand U24514 (N_24514,N_18125,N_13761);
nor U24515 (N_24515,N_14162,N_18485);
nor U24516 (N_24516,N_17715,N_15980);
and U24517 (N_24517,N_16401,N_17712);
nor U24518 (N_24518,N_17182,N_13093);
or U24519 (N_24519,N_17029,N_12693);
nand U24520 (N_24520,N_15029,N_18378);
and U24521 (N_24521,N_14237,N_17929);
xnor U24522 (N_24522,N_14395,N_12609);
and U24523 (N_24523,N_18184,N_13789);
or U24524 (N_24524,N_16086,N_14477);
or U24525 (N_24525,N_13782,N_13354);
nor U24526 (N_24526,N_18406,N_18403);
nand U24527 (N_24527,N_14042,N_18296);
xnor U24528 (N_24528,N_18658,N_16938);
and U24529 (N_24529,N_18153,N_14072);
or U24530 (N_24530,N_14648,N_13972);
or U24531 (N_24531,N_16086,N_16691);
and U24532 (N_24532,N_14998,N_12836);
and U24533 (N_24533,N_17464,N_12928);
or U24534 (N_24534,N_13290,N_13844);
and U24535 (N_24535,N_13990,N_18529);
nor U24536 (N_24536,N_18592,N_16269);
and U24537 (N_24537,N_15910,N_18180);
nand U24538 (N_24538,N_17691,N_14578);
nor U24539 (N_24539,N_13826,N_15708);
nor U24540 (N_24540,N_16183,N_17687);
nand U24541 (N_24541,N_13129,N_18044);
nor U24542 (N_24542,N_18529,N_16904);
xor U24543 (N_24543,N_16283,N_13895);
or U24544 (N_24544,N_13488,N_13424);
nor U24545 (N_24545,N_14362,N_13430);
nor U24546 (N_24546,N_16015,N_18045);
xnor U24547 (N_24547,N_13164,N_14505);
xnor U24548 (N_24548,N_16088,N_16734);
or U24549 (N_24549,N_17002,N_17402);
nand U24550 (N_24550,N_12834,N_15058);
nor U24551 (N_24551,N_15911,N_13063);
and U24552 (N_24552,N_13958,N_13860);
nor U24553 (N_24553,N_13155,N_17977);
and U24554 (N_24554,N_15272,N_12763);
nand U24555 (N_24555,N_16933,N_16714);
nand U24556 (N_24556,N_15250,N_14280);
and U24557 (N_24557,N_12817,N_13464);
nand U24558 (N_24558,N_13881,N_16539);
or U24559 (N_24559,N_13862,N_14071);
xor U24560 (N_24560,N_18296,N_18469);
nor U24561 (N_24561,N_16261,N_12661);
and U24562 (N_24562,N_17319,N_13312);
and U24563 (N_24563,N_17644,N_15998);
nand U24564 (N_24564,N_16559,N_16166);
and U24565 (N_24565,N_12563,N_13364);
nand U24566 (N_24566,N_18440,N_17581);
and U24567 (N_24567,N_15329,N_15806);
or U24568 (N_24568,N_14634,N_13300);
nand U24569 (N_24569,N_12776,N_14663);
nor U24570 (N_24570,N_16801,N_15961);
xnor U24571 (N_24571,N_16086,N_15390);
nor U24572 (N_24572,N_14840,N_15173);
nand U24573 (N_24573,N_18410,N_13495);
nand U24574 (N_24574,N_17896,N_15231);
xor U24575 (N_24575,N_17337,N_16273);
or U24576 (N_24576,N_14712,N_17439);
xnor U24577 (N_24577,N_18723,N_14411);
nor U24578 (N_24578,N_14011,N_13569);
nor U24579 (N_24579,N_17407,N_16288);
and U24580 (N_24580,N_18428,N_16647);
nor U24581 (N_24581,N_16143,N_12636);
nor U24582 (N_24582,N_15594,N_15348);
nand U24583 (N_24583,N_17518,N_16843);
nor U24584 (N_24584,N_17216,N_16808);
or U24585 (N_24585,N_17101,N_18696);
nand U24586 (N_24586,N_16194,N_15651);
xor U24587 (N_24587,N_13397,N_16950);
or U24588 (N_24588,N_16851,N_13096);
xor U24589 (N_24589,N_14208,N_17643);
nand U24590 (N_24590,N_13992,N_16024);
nor U24591 (N_24591,N_13127,N_15674);
or U24592 (N_24592,N_15629,N_13594);
nor U24593 (N_24593,N_13357,N_13594);
and U24594 (N_24594,N_13705,N_18060);
nand U24595 (N_24595,N_18453,N_14003);
nor U24596 (N_24596,N_15170,N_14331);
or U24597 (N_24597,N_18051,N_16742);
nor U24598 (N_24598,N_16516,N_17295);
or U24599 (N_24599,N_13936,N_14136);
nand U24600 (N_24600,N_13587,N_18542);
xor U24601 (N_24601,N_16998,N_18182);
and U24602 (N_24602,N_13213,N_18477);
and U24603 (N_24603,N_18149,N_14895);
or U24604 (N_24604,N_16269,N_16948);
nand U24605 (N_24605,N_15174,N_13568);
nor U24606 (N_24606,N_18520,N_15518);
and U24607 (N_24607,N_13537,N_13553);
or U24608 (N_24608,N_16309,N_15299);
nor U24609 (N_24609,N_16102,N_13093);
or U24610 (N_24610,N_17069,N_17278);
xor U24611 (N_24611,N_14337,N_13884);
nand U24612 (N_24612,N_18683,N_15620);
xor U24613 (N_24613,N_16935,N_13478);
nand U24614 (N_24614,N_16538,N_17868);
nor U24615 (N_24615,N_17159,N_14422);
or U24616 (N_24616,N_15929,N_14345);
and U24617 (N_24617,N_17660,N_17600);
xnor U24618 (N_24618,N_16799,N_18472);
or U24619 (N_24619,N_15468,N_13270);
nor U24620 (N_24620,N_16139,N_15804);
or U24621 (N_24621,N_14429,N_15038);
xnor U24622 (N_24622,N_15376,N_13046);
or U24623 (N_24623,N_14793,N_15213);
nand U24624 (N_24624,N_14818,N_12739);
nand U24625 (N_24625,N_14406,N_15853);
and U24626 (N_24626,N_17372,N_15990);
or U24627 (N_24627,N_15225,N_15641);
and U24628 (N_24628,N_12608,N_17123);
nor U24629 (N_24629,N_14792,N_18699);
or U24630 (N_24630,N_18033,N_16449);
xnor U24631 (N_24631,N_14567,N_17598);
nand U24632 (N_24632,N_18726,N_14221);
nand U24633 (N_24633,N_14982,N_13605);
nand U24634 (N_24634,N_12541,N_17163);
or U24635 (N_24635,N_14786,N_15702);
and U24636 (N_24636,N_17001,N_15092);
nor U24637 (N_24637,N_14371,N_14785);
or U24638 (N_24638,N_16776,N_17574);
or U24639 (N_24639,N_16822,N_14331);
nand U24640 (N_24640,N_17741,N_13064);
nor U24641 (N_24641,N_14544,N_14622);
and U24642 (N_24642,N_13915,N_15736);
xor U24643 (N_24643,N_18166,N_16683);
and U24644 (N_24644,N_17918,N_16788);
nor U24645 (N_24645,N_16526,N_15487);
nand U24646 (N_24646,N_15133,N_13490);
and U24647 (N_24647,N_17629,N_14081);
xor U24648 (N_24648,N_17318,N_13028);
and U24649 (N_24649,N_12738,N_13510);
or U24650 (N_24650,N_12979,N_18109);
nand U24651 (N_24651,N_14862,N_12988);
or U24652 (N_24652,N_17743,N_12884);
and U24653 (N_24653,N_18012,N_15270);
or U24654 (N_24654,N_16995,N_16571);
nand U24655 (N_24655,N_14109,N_17604);
nor U24656 (N_24656,N_18182,N_15227);
nor U24657 (N_24657,N_13104,N_13840);
nand U24658 (N_24658,N_13635,N_16971);
nand U24659 (N_24659,N_17871,N_16417);
and U24660 (N_24660,N_13725,N_16978);
or U24661 (N_24661,N_16011,N_16190);
and U24662 (N_24662,N_15861,N_16953);
xnor U24663 (N_24663,N_14196,N_16320);
or U24664 (N_24664,N_15265,N_18113);
or U24665 (N_24665,N_14819,N_13720);
or U24666 (N_24666,N_15075,N_13445);
or U24667 (N_24667,N_18322,N_18335);
or U24668 (N_24668,N_15139,N_18051);
nor U24669 (N_24669,N_14503,N_14258);
nand U24670 (N_24670,N_15012,N_14834);
and U24671 (N_24671,N_13758,N_13853);
nor U24672 (N_24672,N_17090,N_12962);
xor U24673 (N_24673,N_18217,N_14247);
xor U24674 (N_24674,N_18643,N_15766);
nor U24675 (N_24675,N_16677,N_13902);
xnor U24676 (N_24676,N_18412,N_17451);
nand U24677 (N_24677,N_16316,N_14537);
nor U24678 (N_24678,N_14269,N_14739);
and U24679 (N_24679,N_15698,N_18404);
and U24680 (N_24680,N_16217,N_16651);
or U24681 (N_24681,N_14751,N_17958);
or U24682 (N_24682,N_15686,N_15876);
xnor U24683 (N_24683,N_14660,N_13033);
nor U24684 (N_24684,N_13601,N_17537);
nor U24685 (N_24685,N_13363,N_15869);
and U24686 (N_24686,N_13810,N_15129);
and U24687 (N_24687,N_14517,N_17837);
nor U24688 (N_24688,N_18256,N_18524);
or U24689 (N_24689,N_18364,N_14742);
nand U24690 (N_24690,N_14955,N_15374);
or U24691 (N_24691,N_12654,N_16155);
xnor U24692 (N_24692,N_12533,N_16796);
xor U24693 (N_24693,N_15731,N_15268);
nor U24694 (N_24694,N_14547,N_13691);
or U24695 (N_24695,N_12702,N_17337);
and U24696 (N_24696,N_13683,N_17778);
xor U24697 (N_24697,N_18221,N_17212);
or U24698 (N_24698,N_13050,N_14137);
or U24699 (N_24699,N_14947,N_13874);
xnor U24700 (N_24700,N_18749,N_14078);
and U24701 (N_24701,N_12573,N_17868);
or U24702 (N_24702,N_15465,N_13351);
nand U24703 (N_24703,N_16644,N_17339);
nor U24704 (N_24704,N_18293,N_18672);
nor U24705 (N_24705,N_16716,N_18025);
nand U24706 (N_24706,N_13226,N_12810);
nand U24707 (N_24707,N_16899,N_13989);
nand U24708 (N_24708,N_14164,N_15067);
nor U24709 (N_24709,N_14235,N_17092);
nand U24710 (N_24710,N_14665,N_16692);
nor U24711 (N_24711,N_14623,N_15199);
xnor U24712 (N_24712,N_12929,N_16637);
xor U24713 (N_24713,N_14936,N_17440);
xnor U24714 (N_24714,N_18560,N_17243);
and U24715 (N_24715,N_17917,N_15684);
nand U24716 (N_24716,N_17482,N_13270);
xnor U24717 (N_24717,N_18018,N_14146);
nand U24718 (N_24718,N_17097,N_16973);
nor U24719 (N_24719,N_13155,N_12884);
nor U24720 (N_24720,N_18315,N_17717);
xor U24721 (N_24721,N_17765,N_14317);
nand U24722 (N_24722,N_16658,N_16555);
or U24723 (N_24723,N_15864,N_13761);
xnor U24724 (N_24724,N_16443,N_13045);
nor U24725 (N_24725,N_12959,N_13290);
and U24726 (N_24726,N_12614,N_12611);
nor U24727 (N_24727,N_17876,N_15741);
or U24728 (N_24728,N_12729,N_15011);
or U24729 (N_24729,N_17203,N_13824);
and U24730 (N_24730,N_18341,N_16687);
nor U24731 (N_24731,N_13178,N_14589);
or U24732 (N_24732,N_15208,N_18625);
nor U24733 (N_24733,N_18276,N_13286);
nand U24734 (N_24734,N_14155,N_14379);
nand U24735 (N_24735,N_13248,N_14436);
nand U24736 (N_24736,N_16669,N_14461);
xnor U24737 (N_24737,N_18216,N_13658);
xor U24738 (N_24738,N_12519,N_15812);
nor U24739 (N_24739,N_16139,N_18200);
nand U24740 (N_24740,N_17582,N_15508);
nand U24741 (N_24741,N_17835,N_18401);
or U24742 (N_24742,N_14086,N_16542);
and U24743 (N_24743,N_13415,N_14418);
xnor U24744 (N_24744,N_17782,N_14439);
xor U24745 (N_24745,N_13335,N_15064);
nand U24746 (N_24746,N_16838,N_18084);
nor U24747 (N_24747,N_16598,N_13615);
and U24748 (N_24748,N_13184,N_12691);
nor U24749 (N_24749,N_16910,N_16734);
nand U24750 (N_24750,N_14344,N_18062);
xor U24751 (N_24751,N_14065,N_17092);
nand U24752 (N_24752,N_12792,N_14522);
nor U24753 (N_24753,N_17799,N_14584);
nor U24754 (N_24754,N_14317,N_15908);
nor U24755 (N_24755,N_16881,N_15472);
or U24756 (N_24756,N_14994,N_16661);
nand U24757 (N_24757,N_12929,N_16948);
or U24758 (N_24758,N_17878,N_16308);
and U24759 (N_24759,N_17191,N_13317);
or U24760 (N_24760,N_16156,N_13120);
nor U24761 (N_24761,N_14610,N_17665);
nand U24762 (N_24762,N_16695,N_13649);
nor U24763 (N_24763,N_17225,N_18012);
and U24764 (N_24764,N_15583,N_17916);
or U24765 (N_24765,N_17431,N_14776);
nand U24766 (N_24766,N_15897,N_15511);
and U24767 (N_24767,N_13217,N_16484);
or U24768 (N_24768,N_17312,N_17041);
xnor U24769 (N_24769,N_17594,N_13239);
xor U24770 (N_24770,N_13961,N_12913);
xor U24771 (N_24771,N_15506,N_17495);
nand U24772 (N_24772,N_18666,N_15359);
nor U24773 (N_24773,N_13774,N_15108);
nor U24774 (N_24774,N_13038,N_15161);
or U24775 (N_24775,N_13911,N_14431);
nor U24776 (N_24776,N_14792,N_14501);
xnor U24777 (N_24777,N_16653,N_13956);
nor U24778 (N_24778,N_12555,N_15924);
xor U24779 (N_24779,N_17663,N_17418);
nor U24780 (N_24780,N_17481,N_13349);
nand U24781 (N_24781,N_12847,N_18519);
and U24782 (N_24782,N_14207,N_14247);
xnor U24783 (N_24783,N_14951,N_18078);
and U24784 (N_24784,N_15567,N_17694);
and U24785 (N_24785,N_13335,N_18676);
nor U24786 (N_24786,N_13307,N_16673);
and U24787 (N_24787,N_14451,N_12763);
or U24788 (N_24788,N_15483,N_12606);
nor U24789 (N_24789,N_14686,N_16533);
xnor U24790 (N_24790,N_15084,N_13867);
nor U24791 (N_24791,N_13323,N_12986);
or U24792 (N_24792,N_18085,N_14309);
or U24793 (N_24793,N_13602,N_17702);
xnor U24794 (N_24794,N_15399,N_13917);
xnor U24795 (N_24795,N_13061,N_12868);
and U24796 (N_24796,N_17532,N_15514);
nor U24797 (N_24797,N_13719,N_17450);
and U24798 (N_24798,N_14895,N_13161);
and U24799 (N_24799,N_14400,N_16615);
and U24800 (N_24800,N_13358,N_15128);
nand U24801 (N_24801,N_12950,N_18406);
or U24802 (N_24802,N_18700,N_18045);
nand U24803 (N_24803,N_15535,N_16927);
nor U24804 (N_24804,N_14918,N_13917);
xnor U24805 (N_24805,N_13655,N_15038);
or U24806 (N_24806,N_14262,N_17501);
nor U24807 (N_24807,N_18327,N_16328);
or U24808 (N_24808,N_12969,N_13852);
nor U24809 (N_24809,N_17950,N_17845);
nor U24810 (N_24810,N_13994,N_12890);
and U24811 (N_24811,N_13530,N_13508);
xor U24812 (N_24812,N_18508,N_16193);
xnor U24813 (N_24813,N_15623,N_17242);
nand U24814 (N_24814,N_14383,N_18587);
and U24815 (N_24815,N_18400,N_14958);
xnor U24816 (N_24816,N_17982,N_18253);
and U24817 (N_24817,N_16484,N_13943);
xnor U24818 (N_24818,N_17059,N_14252);
nand U24819 (N_24819,N_16524,N_13493);
nor U24820 (N_24820,N_18226,N_14107);
nor U24821 (N_24821,N_13801,N_12817);
or U24822 (N_24822,N_16851,N_13800);
or U24823 (N_24823,N_13420,N_14915);
xor U24824 (N_24824,N_16291,N_15926);
nand U24825 (N_24825,N_17678,N_13920);
and U24826 (N_24826,N_18333,N_13164);
xnor U24827 (N_24827,N_13797,N_13332);
and U24828 (N_24828,N_15163,N_12603);
or U24829 (N_24829,N_16167,N_14967);
nor U24830 (N_24830,N_13181,N_14236);
xor U24831 (N_24831,N_16638,N_17799);
nand U24832 (N_24832,N_18019,N_14520);
or U24833 (N_24833,N_18440,N_15388);
and U24834 (N_24834,N_18094,N_18211);
nor U24835 (N_24835,N_14492,N_17654);
nand U24836 (N_24836,N_14778,N_13284);
and U24837 (N_24837,N_17615,N_16477);
or U24838 (N_24838,N_15696,N_18716);
and U24839 (N_24839,N_15072,N_16322);
nor U24840 (N_24840,N_15162,N_16414);
xnor U24841 (N_24841,N_13738,N_12653);
or U24842 (N_24842,N_12908,N_15253);
nand U24843 (N_24843,N_13371,N_12849);
xnor U24844 (N_24844,N_14474,N_13862);
xnor U24845 (N_24845,N_14075,N_16152);
xor U24846 (N_24846,N_18533,N_18432);
nand U24847 (N_24847,N_12596,N_12954);
nor U24848 (N_24848,N_13211,N_16585);
nor U24849 (N_24849,N_13245,N_18457);
nor U24850 (N_24850,N_15176,N_18484);
xor U24851 (N_24851,N_15183,N_13069);
nor U24852 (N_24852,N_15845,N_15681);
xor U24853 (N_24853,N_15777,N_18726);
nand U24854 (N_24854,N_13401,N_18575);
xnor U24855 (N_24855,N_14545,N_16970);
or U24856 (N_24856,N_16912,N_14082);
or U24857 (N_24857,N_13762,N_12600);
and U24858 (N_24858,N_15312,N_15585);
and U24859 (N_24859,N_18313,N_15840);
and U24860 (N_24860,N_17007,N_13150);
xor U24861 (N_24861,N_17597,N_14400);
nand U24862 (N_24862,N_12832,N_13491);
xnor U24863 (N_24863,N_17495,N_14952);
xor U24864 (N_24864,N_14105,N_12705);
nor U24865 (N_24865,N_13180,N_18117);
nor U24866 (N_24866,N_18623,N_17832);
or U24867 (N_24867,N_13715,N_15627);
or U24868 (N_24868,N_17637,N_12797);
and U24869 (N_24869,N_17035,N_15865);
xor U24870 (N_24870,N_13009,N_16547);
nand U24871 (N_24871,N_14746,N_14494);
nor U24872 (N_24872,N_16602,N_14503);
nor U24873 (N_24873,N_14809,N_14355);
nor U24874 (N_24874,N_13151,N_13818);
nor U24875 (N_24875,N_14868,N_16858);
or U24876 (N_24876,N_17601,N_12893);
and U24877 (N_24877,N_13207,N_15010);
or U24878 (N_24878,N_15235,N_14386);
xor U24879 (N_24879,N_13227,N_16431);
nand U24880 (N_24880,N_16188,N_13440);
or U24881 (N_24881,N_17813,N_16560);
nand U24882 (N_24882,N_16522,N_17003);
xor U24883 (N_24883,N_13100,N_12549);
xnor U24884 (N_24884,N_15361,N_15072);
or U24885 (N_24885,N_16465,N_17182);
nand U24886 (N_24886,N_14662,N_17701);
and U24887 (N_24887,N_13756,N_15113);
and U24888 (N_24888,N_17541,N_17830);
nor U24889 (N_24889,N_14911,N_14241);
xnor U24890 (N_24890,N_17665,N_14952);
and U24891 (N_24891,N_16744,N_17881);
nor U24892 (N_24892,N_14938,N_14225);
nand U24893 (N_24893,N_15859,N_18076);
nor U24894 (N_24894,N_15206,N_13069);
or U24895 (N_24895,N_18652,N_13880);
nor U24896 (N_24896,N_15523,N_17134);
nor U24897 (N_24897,N_18607,N_16368);
xnor U24898 (N_24898,N_17737,N_15187);
and U24899 (N_24899,N_14689,N_17259);
nand U24900 (N_24900,N_12666,N_15543);
nand U24901 (N_24901,N_15143,N_13484);
nand U24902 (N_24902,N_18519,N_18507);
nor U24903 (N_24903,N_17441,N_15352);
or U24904 (N_24904,N_17057,N_14124);
or U24905 (N_24905,N_16111,N_13177);
xor U24906 (N_24906,N_16060,N_17517);
nor U24907 (N_24907,N_16866,N_16527);
or U24908 (N_24908,N_13726,N_18660);
or U24909 (N_24909,N_18035,N_14651);
and U24910 (N_24910,N_14979,N_15526);
nand U24911 (N_24911,N_16370,N_18382);
nand U24912 (N_24912,N_17650,N_18329);
nor U24913 (N_24913,N_12890,N_13387);
nor U24914 (N_24914,N_14811,N_14201);
and U24915 (N_24915,N_16245,N_13217);
nor U24916 (N_24916,N_12650,N_13826);
nor U24917 (N_24917,N_16103,N_14271);
and U24918 (N_24918,N_13733,N_14764);
nand U24919 (N_24919,N_14751,N_12747);
nand U24920 (N_24920,N_16382,N_15038);
or U24921 (N_24921,N_15228,N_17069);
or U24922 (N_24922,N_15048,N_15525);
or U24923 (N_24923,N_12742,N_13998);
and U24924 (N_24924,N_13007,N_16537);
and U24925 (N_24925,N_14514,N_18616);
xnor U24926 (N_24926,N_13914,N_18511);
or U24927 (N_24927,N_15306,N_12874);
nand U24928 (N_24928,N_16891,N_14899);
and U24929 (N_24929,N_14571,N_15690);
xnor U24930 (N_24930,N_16059,N_12971);
or U24931 (N_24931,N_16057,N_17655);
or U24932 (N_24932,N_13155,N_12702);
nand U24933 (N_24933,N_12724,N_17799);
or U24934 (N_24934,N_16418,N_13396);
or U24935 (N_24935,N_15939,N_15488);
nand U24936 (N_24936,N_14914,N_13022);
nand U24937 (N_24937,N_13579,N_15100);
or U24938 (N_24938,N_13566,N_13784);
nand U24939 (N_24939,N_17831,N_14129);
or U24940 (N_24940,N_16133,N_14979);
xor U24941 (N_24941,N_13829,N_16613);
nor U24942 (N_24942,N_14544,N_14703);
nand U24943 (N_24943,N_13108,N_15523);
or U24944 (N_24944,N_16376,N_13931);
nand U24945 (N_24945,N_16222,N_15446);
and U24946 (N_24946,N_15169,N_18288);
xor U24947 (N_24947,N_18063,N_18534);
or U24948 (N_24948,N_18283,N_16394);
or U24949 (N_24949,N_18561,N_16031);
xor U24950 (N_24950,N_18060,N_17558);
or U24951 (N_24951,N_14906,N_14335);
xor U24952 (N_24952,N_17123,N_15236);
nor U24953 (N_24953,N_16416,N_15882);
nand U24954 (N_24954,N_16618,N_14892);
or U24955 (N_24955,N_12787,N_14600);
and U24956 (N_24956,N_12890,N_16376);
or U24957 (N_24957,N_13559,N_13091);
nor U24958 (N_24958,N_17010,N_16894);
xor U24959 (N_24959,N_17590,N_18039);
nand U24960 (N_24960,N_13785,N_17055);
or U24961 (N_24961,N_15131,N_12698);
nor U24962 (N_24962,N_17585,N_13775);
nand U24963 (N_24963,N_13574,N_14791);
nor U24964 (N_24964,N_15235,N_16377);
or U24965 (N_24965,N_15818,N_14287);
xnor U24966 (N_24966,N_15751,N_12718);
nand U24967 (N_24967,N_13910,N_17311);
or U24968 (N_24968,N_17475,N_17573);
nor U24969 (N_24969,N_18376,N_16407);
xnor U24970 (N_24970,N_15391,N_14683);
nand U24971 (N_24971,N_16118,N_17092);
nor U24972 (N_24972,N_17444,N_12927);
xor U24973 (N_24973,N_14338,N_15716);
nand U24974 (N_24974,N_17126,N_17794);
nor U24975 (N_24975,N_12751,N_13584);
nor U24976 (N_24976,N_18196,N_12773);
or U24977 (N_24977,N_14442,N_14862);
nor U24978 (N_24978,N_13210,N_14216);
or U24979 (N_24979,N_14410,N_17954);
nand U24980 (N_24980,N_12863,N_15511);
nor U24981 (N_24981,N_12819,N_13789);
or U24982 (N_24982,N_13727,N_13247);
and U24983 (N_24983,N_18402,N_16320);
or U24984 (N_24984,N_14669,N_16273);
nand U24985 (N_24985,N_12854,N_18367);
nand U24986 (N_24986,N_17847,N_12627);
or U24987 (N_24987,N_15800,N_13540);
or U24988 (N_24988,N_13234,N_17048);
xnor U24989 (N_24989,N_13218,N_17722);
xor U24990 (N_24990,N_17118,N_15367);
and U24991 (N_24991,N_17542,N_16709);
nand U24992 (N_24992,N_17025,N_14257);
nand U24993 (N_24993,N_18252,N_17095);
xnor U24994 (N_24994,N_17301,N_16808);
nor U24995 (N_24995,N_15925,N_17139);
nand U24996 (N_24996,N_15592,N_16638);
and U24997 (N_24997,N_18156,N_13657);
and U24998 (N_24998,N_13567,N_17895);
nor U24999 (N_24999,N_15096,N_15456);
or UO_0 (O_0,N_19328,N_24782);
nand UO_1 (O_1,N_19029,N_23013);
and UO_2 (O_2,N_23706,N_22502);
or UO_3 (O_3,N_22556,N_24762);
and UO_4 (O_4,N_24417,N_20248);
nand UO_5 (O_5,N_24586,N_20759);
and UO_6 (O_6,N_22444,N_19018);
and UO_7 (O_7,N_20305,N_24617);
nor UO_8 (O_8,N_20447,N_24907);
and UO_9 (O_9,N_22697,N_21661);
nor UO_10 (O_10,N_22861,N_20843);
xor UO_11 (O_11,N_20198,N_21639);
and UO_12 (O_12,N_20584,N_21276);
xor UO_13 (O_13,N_24802,N_24518);
xnor UO_14 (O_14,N_21966,N_23730);
or UO_15 (O_15,N_19418,N_21588);
and UO_16 (O_16,N_20822,N_19823);
xor UO_17 (O_17,N_24777,N_24727);
and UO_18 (O_18,N_23046,N_18941);
nand UO_19 (O_19,N_24489,N_19549);
nand UO_20 (O_20,N_19233,N_23161);
or UO_21 (O_21,N_23908,N_23763);
or UO_22 (O_22,N_20910,N_20098);
and UO_23 (O_23,N_21616,N_20211);
and UO_24 (O_24,N_22156,N_19753);
nor UO_25 (O_25,N_22165,N_20336);
xnor UO_26 (O_26,N_21222,N_22467);
or UO_27 (O_27,N_24277,N_21043);
or UO_28 (O_28,N_24382,N_19963);
xor UO_29 (O_29,N_23236,N_24060);
or UO_30 (O_30,N_24042,N_20527);
xor UO_31 (O_31,N_22016,N_19196);
or UO_32 (O_32,N_21817,N_24288);
nand UO_33 (O_33,N_22990,N_24707);
or UO_34 (O_34,N_22186,N_19281);
nand UO_35 (O_35,N_23915,N_19271);
nor UO_36 (O_36,N_24068,N_22857);
and UO_37 (O_37,N_19745,N_22942);
nand UO_38 (O_38,N_22080,N_23426);
nor UO_39 (O_39,N_21064,N_21181);
or UO_40 (O_40,N_21049,N_19080);
and UO_41 (O_41,N_19353,N_24211);
nand UO_42 (O_42,N_20048,N_22635);
nor UO_43 (O_43,N_24520,N_21145);
and UO_44 (O_44,N_21589,N_18849);
or UO_45 (O_45,N_19439,N_21005);
nand UO_46 (O_46,N_22718,N_23647);
nand UO_47 (O_47,N_19369,N_23901);
and UO_48 (O_48,N_22298,N_23356);
xnor UO_49 (O_49,N_19969,N_24569);
or UO_50 (O_50,N_21576,N_20990);
nand UO_51 (O_51,N_19816,N_23207);
or UO_52 (O_52,N_22243,N_20650);
nand UO_53 (O_53,N_24840,N_19175);
or UO_54 (O_54,N_23009,N_18765);
and UO_55 (O_55,N_20823,N_22076);
nand UO_56 (O_56,N_24602,N_20763);
xor UO_57 (O_57,N_19895,N_23537);
or UO_58 (O_58,N_18993,N_23972);
nand UO_59 (O_59,N_22272,N_20637);
nor UO_60 (O_60,N_19038,N_19257);
nor UO_61 (O_61,N_21165,N_22501);
nor UO_62 (O_62,N_19164,N_22085);
and UO_63 (O_63,N_23484,N_19903);
nand UO_64 (O_64,N_21266,N_20927);
and UO_65 (O_65,N_23867,N_21082);
nor UO_66 (O_66,N_21006,N_23401);
xnor UO_67 (O_67,N_23181,N_18850);
nand UO_68 (O_68,N_23290,N_19800);
nor UO_69 (O_69,N_21887,N_19635);
or UO_70 (O_70,N_24089,N_23542);
or UO_71 (O_71,N_21171,N_23215);
nand UO_72 (O_72,N_21342,N_18790);
or UO_73 (O_73,N_20804,N_21925);
or UO_74 (O_74,N_22258,N_19775);
nand UO_75 (O_75,N_21126,N_23228);
and UO_76 (O_76,N_23053,N_24126);
xnor UO_77 (O_77,N_19146,N_22565);
nand UO_78 (O_78,N_23322,N_19151);
and UO_79 (O_79,N_21139,N_21875);
nand UO_80 (O_80,N_18878,N_21620);
xnor UO_81 (O_81,N_23131,N_18986);
nor UO_82 (O_82,N_19651,N_21728);
xnor UO_83 (O_83,N_24379,N_21448);
nor UO_84 (O_84,N_23240,N_23648);
or UO_85 (O_85,N_23944,N_20112);
or UO_86 (O_86,N_23381,N_20391);
nand UO_87 (O_87,N_21852,N_24553);
nor UO_88 (O_88,N_19299,N_24452);
xor UO_89 (O_89,N_22630,N_19639);
nor UO_90 (O_90,N_19646,N_18983);
or UO_91 (O_91,N_22349,N_23510);
or UO_92 (O_92,N_23835,N_22644);
nand UO_93 (O_93,N_18817,N_20782);
nand UO_94 (O_94,N_20644,N_22285);
or UO_95 (O_95,N_19998,N_23591);
or UO_96 (O_96,N_23079,N_21940);
xnor UO_97 (O_97,N_24665,N_19493);
and UO_98 (O_98,N_19324,N_22372);
and UO_99 (O_99,N_20912,N_20406);
or UO_100 (O_100,N_23932,N_22503);
or UO_101 (O_101,N_18798,N_20877);
nand UO_102 (O_102,N_22054,N_21409);
or UO_103 (O_103,N_21060,N_19055);
nand UO_104 (O_104,N_23808,N_21054);
and UO_105 (O_105,N_22541,N_23012);
nor UO_106 (O_106,N_23738,N_20466);
nand UO_107 (O_107,N_20742,N_21882);
or UO_108 (O_108,N_19276,N_23249);
nor UO_109 (O_109,N_22177,N_21317);
or UO_110 (O_110,N_19723,N_21377);
nand UO_111 (O_111,N_19932,N_23097);
nand UO_112 (O_112,N_22577,N_24831);
nor UO_113 (O_113,N_23801,N_21028);
nand UO_114 (O_114,N_21854,N_24138);
and UO_115 (O_115,N_22267,N_24273);
nor UO_116 (O_116,N_20239,N_21952);
nand UO_117 (O_117,N_22595,N_22129);
or UO_118 (O_118,N_20163,N_23747);
nand UO_119 (O_119,N_24749,N_19312);
and UO_120 (O_120,N_24685,N_20178);
nor UO_121 (O_121,N_20328,N_21295);
and UO_122 (O_122,N_21233,N_23736);
xnor UO_123 (O_123,N_24580,N_18877);
or UO_124 (O_124,N_23552,N_18928);
nor UO_125 (O_125,N_22708,N_19384);
nand UO_126 (O_126,N_23470,N_23128);
xnor UO_127 (O_127,N_22189,N_20977);
nand UO_128 (O_128,N_24920,N_24186);
and UO_129 (O_129,N_24212,N_24978);
or UO_130 (O_130,N_19781,N_21236);
nand UO_131 (O_131,N_19189,N_22506);
nand UO_132 (O_132,N_20709,N_18873);
nand UO_133 (O_133,N_19171,N_23869);
xor UO_134 (O_134,N_22803,N_23540);
nor UO_135 (O_135,N_23694,N_23597);
or UO_136 (O_136,N_23672,N_19769);
nor UO_137 (O_137,N_22031,N_19143);
and UO_138 (O_138,N_23882,N_24041);
and UO_139 (O_139,N_24483,N_24949);
nand UO_140 (O_140,N_23222,N_20740);
nand UO_141 (O_141,N_22905,N_19943);
nor UO_142 (O_142,N_23538,N_19843);
nor UO_143 (O_143,N_18914,N_20933);
xnor UO_144 (O_144,N_22801,N_19047);
or UO_145 (O_145,N_24613,N_24704);
or UO_146 (O_146,N_24551,N_18962);
and UO_147 (O_147,N_22854,N_19313);
nor UO_148 (O_148,N_24645,N_24303);
nand UO_149 (O_149,N_18769,N_21474);
and UO_150 (O_150,N_23146,N_24000);
nor UO_151 (O_151,N_23898,N_23057);
and UO_152 (O_152,N_19004,N_22877);
nor UO_153 (O_153,N_20777,N_24440);
nor UO_154 (O_154,N_21623,N_19126);
nand UO_155 (O_155,N_23091,N_23567);
and UO_156 (O_156,N_20187,N_22005);
or UO_157 (O_157,N_23216,N_19341);
nand UO_158 (O_158,N_20593,N_21085);
nor UO_159 (O_159,N_23679,N_22217);
and UO_160 (O_160,N_23986,N_23230);
xor UO_161 (O_161,N_21155,N_21142);
nor UO_162 (O_162,N_19455,N_21821);
nand UO_163 (O_163,N_20561,N_19444);
or UO_164 (O_164,N_20497,N_22432);
xor UO_165 (O_165,N_21938,N_24479);
xnor UO_166 (O_166,N_22423,N_20284);
and UO_167 (O_167,N_24540,N_20087);
nor UO_168 (O_168,N_20318,N_20224);
or UO_169 (O_169,N_24607,N_24110);
xnor UO_170 (O_170,N_23757,N_20199);
xnor UO_171 (O_171,N_22131,N_19459);
nand UO_172 (O_172,N_19861,N_24106);
or UO_173 (O_173,N_19794,N_23967);
nand UO_174 (O_174,N_20312,N_20660);
or UO_175 (O_175,N_24221,N_21964);
and UO_176 (O_176,N_19486,N_19584);
nand UO_177 (O_177,N_20510,N_24087);
or UO_178 (O_178,N_22188,N_24485);
nand UO_179 (O_179,N_21238,N_20322);
or UO_180 (O_180,N_24388,N_22769);
or UO_181 (O_181,N_23776,N_20960);
nand UO_182 (O_182,N_21723,N_22438);
or UO_183 (O_183,N_20619,N_24400);
nand UO_184 (O_184,N_22086,N_19757);
or UO_185 (O_185,N_21449,N_23366);
or UO_186 (O_186,N_21184,N_22344);
nand UO_187 (O_187,N_22914,N_23008);
nand UO_188 (O_188,N_18751,N_24732);
nor UO_189 (O_189,N_23572,N_24583);
nand UO_190 (O_190,N_22487,N_22961);
nand UO_191 (O_191,N_22239,N_20119);
nand UO_192 (O_192,N_23785,N_19037);
xnor UO_193 (O_193,N_20071,N_23697);
xnor UO_194 (O_194,N_22985,N_24958);
xnor UO_195 (O_195,N_20184,N_21844);
nor UO_196 (O_196,N_18978,N_20417);
and UO_197 (O_197,N_21009,N_24990);
nand UO_198 (O_198,N_19468,N_19566);
nand UO_199 (O_199,N_21129,N_21038);
nand UO_200 (O_200,N_19934,N_21579);
nand UO_201 (O_201,N_24472,N_20679);
nor UO_202 (O_202,N_23621,N_24204);
and UO_203 (O_203,N_22172,N_19526);
and UO_204 (O_204,N_19501,N_18801);
nand UO_205 (O_205,N_21700,N_19929);
and UO_206 (O_206,N_22709,N_22325);
xor UO_207 (O_207,N_20330,N_20281);
xnor UO_208 (O_208,N_22232,N_19691);
or UO_209 (O_209,N_24250,N_23098);
or UO_210 (O_210,N_21625,N_22822);
and UO_211 (O_211,N_24092,N_23622);
or UO_212 (O_212,N_22616,N_21857);
or UO_213 (O_213,N_23943,N_19093);
and UO_214 (O_214,N_23545,N_24023);
nand UO_215 (O_215,N_21841,N_21785);
nand UO_216 (O_216,N_24073,N_19531);
nand UO_217 (O_217,N_23047,N_21806);
xnor UO_218 (O_218,N_21895,N_23305);
or UO_219 (O_219,N_19590,N_21663);
nor UO_220 (O_220,N_22557,N_20247);
or UO_221 (O_221,N_24812,N_20196);
and UO_222 (O_222,N_21051,N_20753);
xnor UO_223 (O_223,N_22802,N_20344);
xnor UO_224 (O_224,N_23522,N_21983);
and UO_225 (O_225,N_22870,N_21715);
xor UO_226 (O_226,N_22437,N_19064);
nand UO_227 (O_227,N_20925,N_18960);
or UO_228 (O_228,N_20842,N_20065);
or UO_229 (O_229,N_20646,N_19655);
or UO_230 (O_230,N_23549,N_22166);
xor UO_231 (O_231,N_21019,N_23947);
or UO_232 (O_232,N_22868,N_19389);
nor UO_233 (O_233,N_20105,N_23383);
xnor UO_234 (O_234,N_19116,N_24450);
nand UO_235 (O_235,N_23384,N_24562);
nand UO_236 (O_236,N_22138,N_20875);
nor UO_237 (O_237,N_22287,N_22661);
nor UO_238 (O_238,N_21725,N_20208);
and UO_239 (O_239,N_20427,N_20773);
nand UO_240 (O_240,N_23171,N_21626);
and UO_241 (O_241,N_19227,N_19669);
nor UO_242 (O_242,N_20939,N_22458);
nand UO_243 (O_243,N_19846,N_20082);
xnor UO_244 (O_244,N_24584,N_20160);
xor UO_245 (O_245,N_23719,N_24251);
xnor UO_246 (O_246,N_22899,N_21702);
xor UO_247 (O_247,N_21297,N_18967);
nor UO_248 (O_248,N_19518,N_21619);
xor UO_249 (O_249,N_21513,N_23420);
or UO_250 (O_250,N_23821,N_24494);
xnor UO_251 (O_251,N_19693,N_23543);
xnor UO_252 (O_252,N_19755,N_21225);
xor UO_253 (O_253,N_18782,N_24497);
nand UO_254 (O_254,N_21826,N_19565);
xnor UO_255 (O_255,N_21269,N_18806);
nand UO_256 (O_256,N_24879,N_21779);
and UO_257 (O_257,N_23805,N_24002);
nor UO_258 (O_258,N_22509,N_19911);
and UO_259 (O_259,N_22969,N_19332);
nor UO_260 (O_260,N_22452,N_21713);
xnor UO_261 (O_261,N_24844,N_20546);
nand UO_262 (O_262,N_19585,N_19904);
and UO_263 (O_263,N_19979,N_24940);
nor UO_264 (O_264,N_19256,N_18864);
and UO_265 (O_265,N_21534,N_19202);
nand UO_266 (O_266,N_23289,N_22976);
nand UO_267 (O_267,N_21587,N_22093);
and UO_268 (O_268,N_22346,N_21402);
xnor UO_269 (O_269,N_21662,N_21041);
and UO_270 (O_270,N_21760,N_20407);
or UO_271 (O_271,N_21419,N_22362);
nor UO_272 (O_272,N_20422,N_20780);
and UO_273 (O_273,N_19153,N_22701);
or UO_274 (O_274,N_24968,N_22040);
and UO_275 (O_275,N_22064,N_22626);
nand UO_276 (O_276,N_21629,N_24107);
or UO_277 (O_277,N_19326,N_20651);
and UO_278 (O_278,N_21967,N_24716);
nor UO_279 (O_279,N_22855,N_19070);
nand UO_280 (O_280,N_21924,N_20325);
and UO_281 (O_281,N_22489,N_23993);
xnor UO_282 (O_282,N_20226,N_18952);
or UO_283 (O_283,N_18870,N_22240);
nand UO_284 (O_284,N_21694,N_19410);
xor UO_285 (O_285,N_20360,N_21791);
nand UO_286 (O_286,N_20693,N_20061);
nor UO_287 (O_287,N_22500,N_21563);
and UO_288 (O_288,N_24960,N_18780);
nor UO_289 (O_289,N_19322,N_22686);
and UO_290 (O_290,N_22132,N_21767);
and UO_291 (O_291,N_22401,N_23663);
xor UO_292 (O_292,N_21511,N_24402);
xnor UO_293 (O_293,N_22035,N_21018);
or UO_294 (O_294,N_18977,N_22561);
or UO_295 (O_295,N_19329,N_23204);
nand UO_296 (O_296,N_22968,N_19849);
and UO_297 (O_297,N_19716,N_23594);
and UO_298 (O_298,N_22691,N_22116);
xnor UO_299 (O_299,N_22864,N_20476);
and UO_300 (O_300,N_18825,N_21193);
nand UO_301 (O_301,N_23134,N_21721);
nand UO_302 (O_302,N_18963,N_22315);
nand UO_303 (O_303,N_21649,N_20726);
and UO_304 (O_304,N_22218,N_24750);
or UO_305 (O_305,N_21315,N_21761);
and UO_306 (O_306,N_21605,N_19790);
nand UO_307 (O_307,N_19947,N_19228);
nand UO_308 (O_308,N_24375,N_22765);
nor UO_309 (O_309,N_21530,N_19300);
xor UO_310 (O_310,N_24367,N_22988);
or UO_311 (O_311,N_22789,N_18866);
nor UO_312 (O_312,N_20575,N_20755);
nor UO_313 (O_313,N_20648,N_19944);
and UO_314 (O_314,N_19851,N_21246);
and UO_315 (O_315,N_23130,N_22780);
or UO_316 (O_316,N_19690,N_21950);
xnor UO_317 (O_317,N_21187,N_19964);
nor UO_318 (O_318,N_24284,N_20157);
or UO_319 (O_319,N_19482,N_24541);
or UO_320 (O_320,N_20775,N_22846);
nand UO_321 (O_321,N_20081,N_23795);
nand UO_322 (O_322,N_23819,N_22453);
nor UO_323 (O_323,N_22830,N_22021);
nand UO_324 (O_324,N_20761,N_20181);
or UO_325 (O_325,N_23950,N_24117);
and UO_326 (O_326,N_22030,N_23499);
or UO_327 (O_327,N_23377,N_22125);
xor UO_328 (O_328,N_19351,N_24604);
and UO_329 (O_329,N_24672,N_20806);
nand UO_330 (O_330,N_24528,N_21306);
and UO_331 (O_331,N_20365,N_20671);
nand UO_332 (O_332,N_20701,N_22073);
xnor UO_333 (O_333,N_19152,N_24931);
and UO_334 (O_334,N_24587,N_21197);
nand UO_335 (O_335,N_21332,N_20586);
xor UO_336 (O_336,N_23772,N_21052);
nand UO_337 (O_337,N_21674,N_23189);
xnor UO_338 (O_338,N_24357,N_23880);
xnor UO_339 (O_339,N_20741,N_20978);
nand UO_340 (O_340,N_21128,N_22429);
and UO_341 (O_341,N_21598,N_23606);
or UO_342 (O_342,N_22746,N_23996);
xor UO_343 (O_343,N_23961,N_20382);
xor UO_344 (O_344,N_19619,N_23214);
or UO_345 (O_345,N_22527,N_23406);
xnor UO_346 (O_346,N_20049,N_24778);
nand UO_347 (O_347,N_24736,N_19742);
xor UO_348 (O_348,N_24136,N_20276);
nand UO_349 (O_349,N_23177,N_18786);
or UO_350 (O_350,N_24619,N_19304);
xor UO_351 (O_351,N_24745,N_20362);
nor UO_352 (O_352,N_20841,N_19124);
nand UO_353 (O_353,N_23589,N_24537);
nor UO_354 (O_354,N_24453,N_21683);
nand UO_355 (O_355,N_19535,N_20275);
nand UO_356 (O_356,N_24090,N_20244);
and UO_357 (O_357,N_18797,N_23242);
and UO_358 (O_358,N_20778,N_19182);
xnor UO_359 (O_359,N_24546,N_20713);
nand UO_360 (O_360,N_23065,N_19251);
or UO_361 (O_361,N_20310,N_23044);
nand UO_362 (O_362,N_24011,N_21370);
and UO_363 (O_363,N_21979,N_24150);
nor UO_364 (O_364,N_18821,N_21135);
or UO_365 (O_365,N_19764,N_21989);
xor UO_366 (O_366,N_21740,N_21098);
or UO_367 (O_367,N_20717,N_19466);
or UO_368 (O_368,N_21220,N_22774);
xnor UO_369 (O_369,N_24398,N_21538);
nand UO_370 (O_370,N_22374,N_19395);
xor UO_371 (O_371,N_21635,N_22796);
or UO_372 (O_372,N_22679,N_19048);
and UO_373 (O_373,N_22548,N_21546);
nor UO_374 (O_374,N_22029,N_20499);
nor UO_375 (O_375,N_24547,N_22482);
nand UO_376 (O_376,N_22282,N_22687);
or UO_377 (O_377,N_22529,N_23565);
xor UO_378 (O_378,N_24156,N_19561);
or UO_379 (O_379,N_20959,N_22462);
nor UO_380 (O_380,N_20571,N_24237);
nand UO_381 (O_381,N_19088,N_24294);
xor UO_382 (O_382,N_21672,N_19978);
nand UO_383 (O_383,N_19442,N_20390);
and UO_384 (O_384,N_19789,N_23331);
and UO_385 (O_385,N_20824,N_19971);
nand UO_386 (O_386,N_23528,N_20902);
and UO_387 (O_387,N_23077,N_21480);
and UO_388 (O_388,N_23203,N_20869);
or UO_389 (O_389,N_24721,N_19259);
nor UO_390 (O_390,N_21633,N_23132);
nand UO_391 (O_391,N_23300,N_24374);
or UO_392 (O_392,N_19719,N_20946);
and UO_393 (O_393,N_20558,N_24696);
or UO_394 (O_394,N_22853,N_18945);
nor UO_395 (O_395,N_22212,N_22614);
and UO_396 (O_396,N_24337,N_24993);
and UO_397 (O_397,N_24193,N_20015);
nand UO_398 (O_398,N_23725,N_24733);
or UO_399 (O_399,N_23011,N_24194);
xor UO_400 (O_400,N_20642,N_18857);
nand UO_401 (O_401,N_22301,N_21828);
and UO_402 (O_402,N_21050,N_20676);
xnor UO_403 (O_403,N_23197,N_23575);
nand UO_404 (O_404,N_24614,N_21078);
nor UO_405 (O_405,N_24019,N_23710);
and UO_406 (O_406,N_21999,N_18950);
xnor UO_407 (O_407,N_20901,N_19279);
or UO_408 (O_408,N_18753,N_21400);
and UO_409 (O_409,N_21354,N_24301);
nand UO_410 (O_410,N_19623,N_23749);
xor UO_411 (O_411,N_24141,N_22963);
xnor UO_412 (O_412,N_23078,N_21754);
nand UO_413 (O_413,N_19484,N_24281);
nand UO_414 (O_414,N_20723,N_24225);
or UO_415 (O_415,N_22304,N_22752);
xnor UO_416 (O_416,N_19137,N_19681);
and UO_417 (O_417,N_23125,N_21170);
nand UO_418 (O_418,N_21809,N_23348);
nor UO_419 (O_419,N_21219,N_19672);
xnor UO_420 (O_420,N_22645,N_22168);
or UO_421 (O_421,N_20080,N_19598);
nand UO_422 (O_422,N_24434,N_23443);
and UO_423 (O_423,N_22024,N_22335);
nand UO_424 (O_424,N_22631,N_21506);
xor UO_425 (O_425,N_22371,N_20398);
xnor UO_426 (O_426,N_24809,N_22551);
and UO_427 (O_427,N_20996,N_20550);
and UO_428 (O_428,N_22533,N_24325);
or UO_429 (O_429,N_23583,N_20278);
nand UO_430 (O_430,N_24845,N_21045);
or UO_431 (O_431,N_24228,N_24677);
and UO_432 (O_432,N_19458,N_23396);
and UO_433 (O_433,N_20212,N_23870);
nand UO_434 (O_434,N_23140,N_23632);
xor UO_435 (O_435,N_20616,N_21404);
or UO_436 (O_436,N_19051,N_19330);
nand UO_437 (O_437,N_20522,N_23464);
and UO_438 (O_438,N_24737,N_19758);
nand UO_439 (O_439,N_19784,N_21729);
xor UO_440 (O_440,N_19144,N_19292);
nand UO_441 (O_441,N_20250,N_24380);
xor UO_442 (O_442,N_19207,N_22422);
nand UO_443 (O_443,N_19890,N_24408);
and UO_444 (O_444,N_21473,N_19751);
nand UO_445 (O_445,N_22747,N_23992);
nand UO_446 (O_446,N_21363,N_22713);
nand UO_447 (O_447,N_19169,N_19948);
nor UO_448 (O_448,N_22339,N_19006);
nand UO_449 (O_449,N_18889,N_24188);
nand UO_450 (O_450,N_19650,N_24903);
or UO_451 (O_451,N_23779,N_24869);
nor UO_452 (O_452,N_23367,N_23989);
or UO_453 (O_453,N_19665,N_22979);
xnor UO_454 (O_454,N_18858,N_23612);
and UO_455 (O_455,N_19335,N_21947);
nor UO_456 (O_456,N_21917,N_23745);
and UO_457 (O_457,N_20712,N_19926);
nor UO_458 (O_458,N_23902,N_24058);
xor UO_459 (O_459,N_22715,N_20203);
or UO_460 (O_460,N_19521,N_23103);
nand UO_461 (O_461,N_20699,N_24558);
or UO_462 (O_462,N_23728,N_21612);
and UO_463 (O_463,N_24895,N_21003);
nor UO_464 (O_464,N_18922,N_19238);
nand UO_465 (O_465,N_23003,N_24446);
nand UO_466 (O_466,N_23831,N_20023);
nand UO_467 (O_467,N_21503,N_19625);
nor UO_468 (O_468,N_23891,N_23655);
and UO_469 (O_469,N_21395,N_22729);
nand UO_470 (O_470,N_20935,N_24873);
or UO_471 (O_471,N_23111,N_21011);
and UO_472 (O_472,N_20132,N_21037);
and UO_473 (O_473,N_24952,N_19604);
or UO_474 (O_474,N_20460,N_23699);
xnor UO_475 (O_475,N_24512,N_19917);
and UO_476 (O_476,N_23068,N_18819);
xor UO_477 (O_477,N_21951,N_21608);
or UO_478 (O_478,N_24169,N_22992);
nor UO_479 (O_479,N_24063,N_22411);
nand UO_480 (O_480,N_20079,N_24729);
xnor UO_481 (O_481,N_23681,N_20641);
xnor UO_482 (O_482,N_24649,N_23350);
nand UO_483 (O_483,N_19877,N_24226);
xnor UO_484 (O_484,N_22824,N_24815);
and UO_485 (O_485,N_20057,N_21023);
or UO_486 (O_486,N_24003,N_22705);
xnor UO_487 (O_487,N_21680,N_22292);
nand UO_488 (O_488,N_19432,N_18981);
or UO_489 (O_489,N_24643,N_19698);
xnor UO_490 (O_490,N_19722,N_23850);
nor UO_491 (O_491,N_19872,N_18848);
nor UO_492 (O_492,N_21256,N_23615);
and UO_493 (O_493,N_21497,N_22930);
xnor UO_494 (O_494,N_23255,N_24673);
and UO_495 (O_495,N_21932,N_22268);
nor UO_496 (O_496,N_23015,N_21777);
or UO_497 (O_497,N_21300,N_20176);
or UO_498 (O_498,N_24373,N_20492);
nand UO_499 (O_499,N_20147,N_24102);
nor UO_500 (O_500,N_24246,N_24425);
nor UO_501 (O_501,N_21012,N_21901);
xor UO_502 (O_502,N_19931,N_20991);
and UO_503 (O_503,N_21816,N_23048);
nand UO_504 (O_504,N_19264,N_23781);
and UO_505 (O_505,N_24217,N_21237);
nor UO_506 (O_506,N_21535,N_24244);
and UO_507 (O_507,N_19562,N_24333);
or UO_508 (O_508,N_21988,N_23372);
xor UO_509 (O_509,N_20025,N_20519);
xnor UO_510 (O_510,N_24418,N_22844);
or UO_511 (O_511,N_19889,N_23887);
xor UO_512 (O_512,N_20215,N_22481);
xnor UO_513 (O_513,N_24948,N_23347);
and UO_514 (O_514,N_21542,N_20458);
nand UO_515 (O_515,N_23539,N_21040);
nor UO_516 (O_516,N_23937,N_24804);
or UO_517 (O_517,N_21211,N_21601);
nor UO_518 (O_518,N_24764,N_24459);
xnor UO_519 (O_519,N_18988,N_21850);
and UO_520 (O_520,N_24793,N_20658);
and UO_521 (O_521,N_23459,N_21460);
or UO_522 (O_522,N_21234,N_20677);
and UO_523 (O_523,N_20152,N_24030);
xor UO_524 (O_524,N_19888,N_21697);
and UO_525 (O_525,N_23453,N_21438);
xor UO_526 (O_526,N_22751,N_23778);
xnor UO_527 (O_527,N_19022,N_23629);
nor UO_528 (O_528,N_21447,N_18859);
xnor UO_529 (O_529,N_22216,N_22749);
xnor UO_530 (O_530,N_21446,N_19415);
and UO_531 (O_531,N_22934,N_19833);
nand UO_532 (O_532,N_24932,N_23531);
or UO_533 (O_533,N_19013,N_21937);
and UO_534 (O_534,N_22307,N_22296);
xnor UO_535 (O_535,N_24921,N_19505);
nor UO_536 (O_536,N_21196,N_20604);
xnor UO_537 (O_537,N_24177,N_23185);
nand UO_538 (O_538,N_23601,N_22209);
xnor UO_539 (O_539,N_24897,N_21732);
nor UO_540 (O_540,N_19508,N_19239);
or UO_541 (O_541,N_19778,N_20088);
nor UO_542 (O_542,N_19197,N_22526);
nand UO_543 (O_543,N_22654,N_23273);
nand UO_544 (O_544,N_21773,N_24045);
and UO_545 (O_545,N_21643,N_24312);
xnor UO_546 (O_546,N_18917,N_21496);
nand UO_547 (O_547,N_22978,N_23382);
xor UO_548 (O_548,N_21328,N_20298);
xnor UO_549 (O_549,N_22478,N_23462);
nand UO_550 (O_550,N_24647,N_23392);
xor UO_551 (O_551,N_22757,N_23557);
nand UO_552 (O_552,N_22998,N_23447);
xnor UO_553 (O_553,N_19558,N_22612);
xor UO_554 (O_554,N_18874,N_19166);
nand UO_555 (O_555,N_19488,N_23371);
xnor UO_556 (O_556,N_21415,N_22202);
and UO_557 (O_557,N_20748,N_23741);
or UO_558 (O_558,N_20092,N_19813);
xnor UO_559 (O_559,N_24519,N_23688);
and UO_560 (O_560,N_20915,N_19956);
nand UO_561 (O_561,N_23686,N_20192);
nor UO_562 (O_562,N_18779,N_21066);
xnor UO_563 (O_563,N_21575,N_24972);
nand UO_564 (O_564,N_23452,N_20636);
nand UO_565 (O_565,N_23337,N_22062);
xor UO_566 (O_566,N_21552,N_20785);
nand UO_567 (O_567,N_19249,N_20289);
and UO_568 (O_568,N_23276,N_23118);
or UO_569 (O_569,N_23262,N_22337);
xnor UO_570 (O_570,N_23683,N_20124);
nand UO_571 (O_571,N_22767,N_18997);
or UO_572 (O_572,N_24914,N_22257);
nand UO_573 (O_573,N_23798,N_22314);
nand UO_574 (O_574,N_21871,N_21144);
and UO_575 (O_575,N_22688,N_20142);
or UO_576 (O_576,N_21281,N_24353);
and UO_577 (O_577,N_19617,N_20821);
nor UO_578 (O_578,N_19959,N_20467);
or UO_579 (O_579,N_22305,N_24208);
xor UO_580 (O_580,N_22164,N_23456);
and UO_581 (O_581,N_19504,N_20078);
xnor UO_582 (O_582,N_19241,N_20858);
or UO_583 (O_583,N_22194,N_23917);
nor UO_584 (O_584,N_20828,N_19933);
nor UO_585 (O_585,N_20591,N_20565);
xnor UO_586 (O_586,N_20523,N_24361);
nand UO_587 (O_587,N_19624,N_21077);
nor UO_588 (O_588,N_18867,N_20610);
nand UO_589 (O_589,N_24910,N_24658);
or UO_590 (O_590,N_23949,N_22417);
xnor UO_591 (O_591,N_21454,N_24571);
and UO_592 (O_592,N_23116,N_19481);
xor UO_593 (O_593,N_21762,N_23005);
xnor UO_594 (O_594,N_21159,N_24984);
xnor UO_595 (O_595,N_20691,N_19627);
xnor UO_596 (O_596,N_19277,N_23623);
or UO_597 (O_597,N_24490,N_21425);
nor UO_598 (O_598,N_21630,N_20323);
nor UO_599 (O_599,N_23573,N_23147);
nor UO_600 (O_600,N_19897,N_24172);
nand UO_601 (O_601,N_21437,N_20412);
nor UO_602 (O_602,N_19016,N_24043);
xnor UO_603 (O_603,N_19920,N_24842);
and UO_604 (O_604,N_19295,N_23909);
nor UO_605 (O_605,N_22028,N_23024);
nand UO_606 (O_606,N_19863,N_23436);
xnor UO_607 (O_607,N_23875,N_23114);
xor UO_608 (O_608,N_20622,N_19125);
nor UO_609 (O_609,N_22171,N_22773);
or UO_610 (O_610,N_21618,N_20953);
nor UO_611 (O_611,N_21031,N_18895);
nor UO_612 (O_612,N_19052,N_21292);
xnor UO_613 (O_613,N_23174,N_23198);
nand UO_614 (O_614,N_23159,N_21693);
nor UO_615 (O_615,N_24539,N_23722);
nor UO_616 (O_616,N_22133,N_21688);
xnor UO_617 (O_617,N_21559,N_24461);
and UO_618 (O_618,N_23871,N_20682);
nor UO_619 (O_619,N_22714,N_23713);
and UO_620 (O_620,N_20032,N_19513);
xor UO_621 (O_621,N_22706,N_24936);
xor UO_622 (O_622,N_22926,N_19763);
xnor UO_623 (O_623,N_24533,N_24059);
nand UO_624 (O_624,N_21800,N_19866);
or UO_625 (O_625,N_20008,N_21529);
or UO_626 (O_626,N_22279,N_24139);
or UO_627 (O_627,N_19883,N_19223);
and UO_628 (O_628,N_20577,N_22837);
and UO_629 (O_629,N_18772,N_19747);
xor UO_630 (O_630,N_23286,N_20002);
nand UO_631 (O_631,N_22648,N_19483);
and UO_632 (O_632,N_20464,N_22762);
and UO_633 (O_633,N_22542,N_21682);
and UO_634 (O_634,N_22681,N_21709);
xnor UO_635 (O_635,N_19771,N_24598);
nand UO_636 (O_636,N_23899,N_24444);
nor UO_637 (O_637,N_22295,N_20881);
xnor UO_638 (O_638,N_24475,N_19390);
xor UO_639 (O_639,N_22136,N_18776);
and UO_640 (O_640,N_22804,N_21868);
nor UO_641 (O_641,N_24293,N_21788);
or UO_642 (O_642,N_20300,N_21792);
or UO_643 (O_643,N_19377,N_23284);
and UO_644 (O_644,N_24791,N_24124);
nand UO_645 (O_645,N_18915,N_20273);
and UO_646 (O_646,N_24708,N_19403);
and UO_647 (O_647,N_21084,N_24753);
xor UO_648 (O_648,N_20317,N_23884);
or UO_649 (O_649,N_19575,N_24074);
nand UO_650 (O_650,N_20058,N_22492);
or UO_651 (O_651,N_21822,N_21519);
or UO_652 (O_652,N_18762,N_23698);
or UO_653 (O_653,N_21162,N_21897);
xor UO_654 (O_654,N_19480,N_23380);
and UO_655 (O_655,N_24698,N_21692);
or UO_656 (O_656,N_24018,N_22892);
or UO_657 (O_657,N_22309,N_21190);
or UO_658 (O_658,N_22673,N_20425);
nand UO_659 (O_659,N_19066,N_20678);
nor UO_660 (O_660,N_19776,N_21798);
or UO_661 (O_661,N_19557,N_19127);
xnor UO_662 (O_662,N_21248,N_19419);
nand UO_663 (O_663,N_22269,N_20907);
xnor UO_664 (O_664,N_20768,N_24849);
nor UO_665 (O_665,N_19629,N_19297);
nand UO_666 (O_666,N_21094,N_24431);
xor UO_667 (O_667,N_22621,N_20805);
xnor UO_668 (O_668,N_21730,N_23178);
and UO_669 (O_669,N_23913,N_19511);
and UO_670 (O_670,N_22039,N_22377);
and UO_671 (O_671,N_21515,N_21093);
or UO_672 (O_672,N_23004,N_21805);
nor UO_673 (O_673,N_21894,N_19555);
or UO_674 (O_674,N_24690,N_22387);
xnor UO_675 (O_675,N_21622,N_24828);
nand UO_676 (O_676,N_20486,N_19008);
nor UO_677 (O_677,N_22038,N_22395);
or UO_678 (O_678,N_24399,N_20718);
xnor UO_679 (O_679,N_19291,N_24635);
nand UO_680 (O_680,N_23138,N_21442);
xnor UO_681 (O_681,N_20480,N_22816);
nor UO_682 (O_682,N_19858,N_19431);
and UO_683 (O_683,N_23939,N_23938);
xor UO_684 (O_684,N_20054,N_20667);
xor UO_685 (O_685,N_21710,N_23006);
nand UO_686 (O_686,N_21765,N_20093);
and UO_687 (O_687,N_23029,N_23554);
and UO_688 (O_688,N_23751,N_24702);
xor UO_689 (O_689,N_20436,N_22419);
nor UO_690 (O_690,N_21888,N_21180);
nor UO_691 (O_691,N_22716,N_20614);
nand UO_692 (O_692,N_19765,N_18777);
or UO_693 (O_693,N_23405,N_20745);
or UO_694 (O_694,N_19670,N_22465);
xor UO_695 (O_695,N_24320,N_21804);
or UO_696 (O_696,N_22360,N_23001);
and UO_697 (O_697,N_20271,N_20257);
and UO_698 (O_698,N_23746,N_20972);
xnor UO_699 (O_699,N_21468,N_20156);
or UO_700 (O_700,N_22664,N_24548);
nor UO_701 (O_701,N_22882,N_19172);
xnor UO_702 (O_702,N_24022,N_24101);
xnor UO_703 (O_703,N_24545,N_21731);
and UO_704 (O_704,N_22871,N_19710);
and UO_705 (O_705,N_19059,N_19730);
and UO_706 (O_706,N_22903,N_24637);
xnor UO_707 (O_707,N_24061,N_23912);
and UO_708 (O_708,N_20468,N_21067);
xnor UO_709 (O_709,N_20973,N_19095);
and UO_710 (O_710,N_24767,N_20272);
or UO_711 (O_711,N_23677,N_23075);
nand UO_712 (O_712,N_21632,N_24760);
and UO_713 (O_713,N_24370,N_23854);
nand UO_714 (O_714,N_24616,N_23379);
nand UO_715 (O_715,N_20779,N_24240);
nor UO_716 (O_716,N_18893,N_24310);
or UO_717 (O_717,N_18781,N_24624);
nand UO_718 (O_718,N_24977,N_22604);
nor UO_719 (O_719,N_21724,N_19777);
xor UO_720 (O_720,N_22966,N_22091);
nor UO_721 (O_721,N_19613,N_21200);
or UO_722 (O_722,N_22678,N_19460);
or UO_723 (O_723,N_20728,N_20094);
nand UO_724 (O_724,N_24340,N_19308);
xnor UO_725 (O_725,N_21357,N_24864);
nand UO_726 (O_726,N_24395,N_21013);
nor UO_727 (O_727,N_23229,N_24148);
or UO_728 (O_728,N_24119,N_21975);
xor UO_729 (O_729,N_22727,N_24476);
nand UO_730 (O_730,N_19782,N_21061);
xnor UO_731 (O_731,N_24860,N_19406);
or UO_732 (O_732,N_22955,N_22745);
nand UO_733 (O_733,N_20452,N_20331);
and UO_734 (O_734,N_24153,N_20041);
and UO_735 (O_735,N_21026,N_20911);
nand UO_736 (O_736,N_23769,N_20433);
and UO_737 (O_737,N_19552,N_21982);
xnor UO_738 (O_738,N_21735,N_21312);
and UO_739 (O_739,N_24180,N_23104);
xnor UO_740 (O_740,N_23876,N_19750);
xor UO_741 (O_741,N_18865,N_19731);
nor UO_742 (O_742,N_23434,N_22986);
or UO_743 (O_743,N_22246,N_24454);
nor UO_744 (O_744,N_22723,N_21056);
nand UO_745 (O_745,N_22370,N_23175);
nor UO_746 (O_746,N_19168,N_20632);
xor UO_747 (O_747,N_21908,N_20228);
xnor UO_748 (O_748,N_23856,N_19834);
or UO_749 (O_749,N_22015,N_20954);
and UO_750 (O_750,N_19438,N_24823);
or UO_751 (O_751,N_19367,N_22543);
nand UO_752 (O_752,N_21379,N_24667);
and UO_753 (O_753,N_24255,N_19305);
or UO_754 (O_754,N_23498,N_20418);
xnor UO_755 (O_755,N_22019,N_18946);
and UO_756 (O_756,N_19302,N_21252);
nand UO_757 (O_757,N_24053,N_20031);
nand UO_758 (O_758,N_23723,N_20020);
nand UO_759 (O_759,N_22071,N_24684);
or UO_760 (O_760,N_18756,N_20700);
xnor UO_761 (O_761,N_23469,N_24332);
xnor UO_762 (O_762,N_20385,N_19011);
and UO_763 (O_763,N_24419,N_21750);
or UO_764 (O_764,N_20168,N_20932);
nor UO_765 (O_765,N_20813,N_19735);
nor UO_766 (O_766,N_23792,N_20304);
nand UO_767 (O_767,N_24116,N_21691);
and UO_768 (O_768,N_23759,N_20258);
xnor UO_769 (O_769,N_20624,N_21824);
and UO_770 (O_770,N_23761,N_21943);
and UO_771 (O_771,N_24013,N_19547);
xnor UO_772 (O_772,N_24681,N_20148);
nor UO_773 (O_773,N_23900,N_23933);
and UO_774 (O_774,N_19475,N_23731);
xor UO_775 (O_775,N_24471,N_22271);
and UO_776 (O_776,N_20440,N_21873);
and UO_777 (O_777,N_22790,N_21703);
or UO_778 (O_778,N_23151,N_23235);
and UO_779 (O_779,N_22777,N_20264);
or UO_780 (O_780,N_20689,N_24631);
xnor UO_781 (O_781,N_24300,N_22977);
xor UO_782 (O_782,N_19633,N_24722);
nand UO_783 (O_783,N_20729,N_20043);
or UO_784 (O_784,N_21778,N_23223);
nor UO_785 (O_785,N_22540,N_24848);
nor UO_786 (O_786,N_21820,N_23524);
nor UO_787 (O_787,N_19366,N_21324);
or UO_788 (O_788,N_18814,N_21573);
or UO_789 (O_789,N_19798,N_22858);
and UO_790 (O_790,N_22149,N_21478);
nand UO_791 (O_791,N_23444,N_24508);
nand UO_792 (O_792,N_21008,N_23948);
nor UO_793 (O_793,N_19900,N_23476);
and UO_794 (O_794,N_24634,N_19808);
and UO_795 (O_795,N_20788,N_21569);
nand UO_796 (O_796,N_22121,N_20930);
or UO_797 (O_797,N_23251,N_23709);
xnor UO_798 (O_798,N_19539,N_21574);
nand UO_799 (O_799,N_24096,N_22638);
and UO_800 (O_800,N_18911,N_19337);
xnor UO_801 (O_801,N_20885,N_20976);
nand UO_802 (O_802,N_22013,N_22699);
xor UO_803 (O_803,N_22569,N_20000);
and UO_804 (O_804,N_19560,N_22842);
nor UO_805 (O_805,N_19357,N_21000);
xnor UO_806 (O_806,N_19157,N_19853);
and UO_807 (O_807,N_24238,N_18860);
nand UO_808 (O_808,N_22032,N_24052);
nor UO_809 (O_809,N_23355,N_24794);
xor UO_810 (O_810,N_19430,N_20692);
and UO_811 (O_811,N_21673,N_22178);
nor UO_812 (O_812,N_22210,N_23605);
xnor UO_813 (O_813,N_20807,N_22011);
and UO_814 (O_814,N_21585,N_18835);
nand UO_815 (O_815,N_22238,N_20267);
nor UO_816 (O_816,N_19601,N_22169);
nand UO_817 (O_817,N_19579,N_21776);
nor UO_818 (O_818,N_20149,N_18879);
nor UO_819 (O_819,N_20450,N_20814);
nand UO_820 (O_820,N_20340,N_20765);
nand UO_821 (O_821,N_22581,N_21501);
or UO_822 (O_822,N_20026,N_21341);
or UO_823 (O_823,N_24286,N_19054);
or UO_824 (O_824,N_22819,N_19138);
xnor UO_825 (O_825,N_23239,N_20299);
nor UO_826 (O_826,N_19413,N_24426);
xnor UO_827 (O_827,N_24334,N_22208);
or UO_828 (O_828,N_22841,N_24044);
nor UO_829 (O_829,N_22646,N_21469);
or UO_830 (O_830,N_24964,N_24710);
nor UO_831 (O_831,N_24348,N_20207);
nand UO_832 (O_832,N_20500,N_21151);
or UO_833 (O_833,N_22682,N_19595);
xor UO_834 (O_834,N_20102,N_21638);
nand UO_835 (O_835,N_21939,N_22034);
xnor UO_836 (O_836,N_21208,N_23495);
or UO_837 (O_837,N_22836,N_22356);
or UO_838 (O_838,N_20889,N_19129);
nand UO_839 (O_839,N_24975,N_22656);
nand UO_840 (O_840,N_24344,N_24953);
and UO_841 (O_841,N_24377,N_23020);
nand UO_842 (O_842,N_23962,N_22469);
nand UO_843 (O_843,N_20846,N_22464);
nor UO_844 (O_844,N_19993,N_22704);
xnor UO_845 (O_845,N_24071,N_22758);
or UO_846 (O_846,N_20415,N_20921);
or UO_847 (O_847,N_23979,N_23056);
nor UO_848 (O_848,N_22354,N_24996);
or UO_849 (O_849,N_19568,N_18810);
nand UO_850 (O_850,N_19147,N_22220);
or UO_851 (O_851,N_22376,N_20702);
nor UO_852 (O_852,N_22303,N_21823);
nor UO_853 (O_853,N_22405,N_19411);
and UO_854 (O_854,N_22135,N_20793);
and UO_855 (O_855,N_22812,N_23339);
and UO_856 (O_856,N_19709,N_22698);
and UO_857 (O_857,N_20227,N_23811);
nor UO_858 (O_858,N_21436,N_20206);
nor UO_859 (O_859,N_19178,N_23315);
or UO_860 (O_860,N_18965,N_19773);
and UO_861 (O_861,N_20014,N_23270);
and UO_862 (O_862,N_20876,N_19695);
xor UO_863 (O_863,N_22984,N_23458);
xnor UO_864 (O_864,N_22154,N_23368);
nand UO_865 (O_865,N_21178,N_19072);
nand UO_866 (O_866,N_20585,N_19510);
or UO_867 (O_867,N_21617,N_21912);
nand UO_868 (O_868,N_24424,N_19974);
and UO_869 (O_869,N_24534,N_24219);
xnor UO_870 (O_870,N_20837,N_23463);
nor UO_871 (O_871,N_20361,N_24363);
xnor UO_872 (O_872,N_20923,N_19951);
or UO_873 (O_873,N_22607,N_22112);
or UO_874 (O_874,N_20789,N_20085);
nor UO_875 (O_875,N_19350,N_20568);
nand UO_876 (O_876,N_19401,N_21784);
and UO_877 (O_877,N_21183,N_23985);
and UO_878 (O_878,N_22211,N_20291);
or UO_879 (O_879,N_24816,N_24771);
and UO_880 (O_880,N_24739,N_22883);
nand UO_881 (O_881,N_19033,N_19461);
or UO_882 (O_882,N_22863,N_21091);
and UO_883 (O_883,N_23312,N_20413);
xor UO_884 (O_884,N_24438,N_23834);
nor UO_885 (O_885,N_24442,N_23303);
xnor UO_886 (O_886,N_18803,N_22920);
or UO_887 (O_887,N_22317,N_22587);
and UO_888 (O_888,N_20983,N_21095);
and UO_889 (O_889,N_19656,N_18898);
or UO_890 (O_890,N_21972,N_20351);
nor UO_891 (O_891,N_19424,N_19131);
or UO_892 (O_892,N_23064,N_23043);
nand UO_893 (O_893,N_19972,N_19186);
nand UO_894 (O_894,N_24055,N_22468);
or UO_895 (O_895,N_20410,N_22907);
nor UO_896 (O_896,N_20261,N_22277);
nand UO_897 (O_897,N_20818,N_22941);
or UO_898 (O_898,N_21073,N_24819);
nor UO_899 (O_899,N_22847,N_22262);
nand UO_900 (O_900,N_20277,N_22668);
xor UO_901 (O_901,N_22316,N_19570);
and UO_902 (O_902,N_24383,N_22550);
nand UO_903 (O_903,N_24198,N_22794);
and UO_904 (O_904,N_18891,N_23244);
nor UO_905 (O_905,N_20509,N_24761);
xor UO_906 (O_906,N_18802,N_22663);
nand UO_907 (O_907,N_22229,N_24467);
or UO_908 (O_908,N_23771,N_21475);
xor UO_909 (O_909,N_23923,N_23465);
nor UO_910 (O_910,N_20150,N_22620);
or UO_911 (O_911,N_22050,N_24299);
and UO_912 (O_912,N_21512,N_18990);
or UO_913 (O_913,N_21247,N_21640);
xor UO_914 (O_914,N_23314,N_22450);
nand UO_915 (O_915,N_20485,N_19728);
and UO_916 (O_916,N_20487,N_22311);
xor UO_917 (O_917,N_23395,N_21571);
nor UO_918 (O_918,N_20653,N_19523);
nor UO_919 (O_919,N_21381,N_22471);
nor UO_920 (O_920,N_22510,N_20399);
nand UO_921 (O_921,N_19532,N_24233);
nand UO_922 (O_922,N_20165,N_22615);
xor UO_923 (O_923,N_23861,N_23378);
xnor UO_924 (O_924,N_24805,N_21592);
nand UO_925 (O_925,N_19519,N_22632);
nor UO_926 (O_926,N_20601,N_22960);
nor UO_927 (O_927,N_23828,N_21564);
nor UO_928 (O_928,N_20620,N_21763);
and UO_929 (O_929,N_19325,N_23477);
and UO_930 (O_930,N_18882,N_22049);
or UO_931 (O_931,N_24773,N_20243);
nand UO_932 (O_932,N_20539,N_22677);
and UO_933 (O_933,N_24473,N_23080);
xor UO_934 (O_934,N_20952,N_22460);
xnor UO_935 (O_935,N_21406,N_20513);
nor UO_936 (O_936,N_23299,N_23165);
or UO_937 (O_937,N_20838,N_23364);
nor UO_938 (O_938,N_23599,N_20984);
nand UO_939 (O_939,N_23560,N_24712);
or UO_940 (O_940,N_23288,N_21965);
nor UO_941 (O_941,N_18855,N_21285);
and UO_942 (O_942,N_21267,N_23129);
and UO_943 (O_943,N_22181,N_20067);
nand UO_944 (O_944,N_22971,N_20801);
xor UO_945 (O_945,N_24621,N_24271);
and UO_946 (O_946,N_23145,N_20180);
nand UO_947 (O_947,N_24252,N_23021);
nor UO_948 (O_948,N_21755,N_23506);
and UO_949 (O_949,N_22957,N_20588);
or UO_950 (O_950,N_22042,N_23267);
xor UO_951 (O_951,N_23791,N_22726);
nand UO_952 (O_952,N_20999,N_22402);
xnor UO_953 (O_953,N_20341,N_22791);
and UO_954 (O_954,N_22110,N_21556);
nand UO_955 (O_955,N_22114,N_19630);
and UO_956 (O_956,N_19333,N_22743);
and UO_957 (O_957,N_18804,N_24366);
and UO_958 (O_958,N_21329,N_24915);
xor UO_959 (O_959,N_22308,N_20400);
and UO_960 (O_960,N_23432,N_23758);
and UO_961 (O_961,N_24752,N_21991);
and UO_962 (O_962,N_21224,N_21081);
nor UO_963 (O_963,N_24898,N_22869);
nor UO_964 (O_964,N_23714,N_23890);
nor UO_965 (O_965,N_22755,N_20209);
or UO_966 (O_966,N_23855,N_20223);
nor UO_967 (O_967,N_21304,N_24115);
or UO_968 (O_968,N_19949,N_23610);
nor UO_969 (O_969,N_19417,N_24428);
xor UO_970 (O_970,N_22495,N_23360);
and UO_971 (O_971,N_24850,N_24725);
and UO_972 (O_972,N_24207,N_24474);
or UO_973 (O_973,N_19024,N_21790);
nand UO_974 (O_974,N_22650,N_23019);
and UO_975 (O_975,N_21491,N_19495);
xor UO_976 (O_976,N_23588,N_21793);
xor UO_977 (O_977,N_20242,N_22591);
nor UO_978 (O_978,N_21388,N_18949);
nand UO_979 (O_979,N_21685,N_23136);
xnor UO_980 (O_980,N_21919,N_18761);
xnor UO_981 (O_981,N_20762,N_21314);
or UO_982 (O_982,N_23297,N_24095);
or UO_983 (O_983,N_21768,N_21811);
nand UO_984 (O_984,N_20238,N_22902);
nor UO_985 (O_985,N_20489,N_24086);
nor UO_986 (O_986,N_23283,N_24679);
or UO_987 (O_987,N_24799,N_21827);
nor UO_988 (O_988,N_23478,N_19573);
nor UO_989 (O_989,N_23903,N_20557);
nor UO_990 (O_990,N_24057,N_23293);
and UO_991 (O_991,N_19477,N_23519);
nor UO_992 (O_992,N_23953,N_19820);
nor UO_993 (O_993,N_23975,N_24132);
nand UO_994 (O_994,N_21087,N_20955);
nand UO_995 (O_995,N_20733,N_22430);
nand UO_996 (O_996,N_22283,N_18842);
nand UO_997 (O_997,N_20766,N_22414);
nand UO_998 (O_998,N_21386,N_24943);
xor UO_999 (O_999,N_23752,N_21435);
nor UO_1000 (O_1000,N_23182,N_24397);
or UO_1001 (O_1001,N_23994,N_22608);
and UO_1002 (O_1002,N_19803,N_23577);
or UO_1003 (O_1003,N_22025,N_24088);
or UO_1004 (O_1004,N_22579,N_21380);
or UO_1005 (O_1005,N_20146,N_23582);
or UO_1006 (O_1006,N_23788,N_22900);
or UO_1007 (O_1007,N_19856,N_24610);
or UO_1008 (O_1008,N_24021,N_22451);
xnor UO_1009 (O_1009,N_23375,N_21780);
xnor UO_1010 (O_1010,N_23211,N_20847);
or UO_1011 (O_1011,N_22554,N_19839);
nand UO_1012 (O_1012,N_22585,N_24109);
or UO_1013 (O_1013,N_22660,N_23700);
xor UO_1014 (O_1014,N_20083,N_24623);
nor UO_1015 (O_1015,N_24403,N_22951);
xor UO_1016 (O_1016,N_21408,N_24856);
or UO_1017 (O_1017,N_20076,N_20516);
nand UO_1018 (O_1018,N_22962,N_19541);
or UO_1019 (O_1019,N_22623,N_23265);
or UO_1020 (O_1020,N_24262,N_22056);
or UO_1021 (O_1021,N_24846,N_22103);
and UO_1022 (O_1022,N_24149,N_19636);
and UO_1023 (O_1023,N_24544,N_19824);
nand UO_1024 (O_1024,N_18794,N_19176);
or UO_1025 (O_1025,N_22162,N_18791);
nor UO_1026 (O_1026,N_23413,N_22627);
or UO_1027 (O_1027,N_23581,N_21839);
xor UO_1028 (O_1028,N_23563,N_22908);
or UO_1029 (O_1029,N_19840,N_20366);
or UO_1030 (O_1030,N_24430,N_19844);
xnor UO_1031 (O_1031,N_19076,N_21560);
or UO_1032 (O_1032,N_23219,N_19334);
and UO_1033 (O_1033,N_24048,N_20784);
xor UO_1034 (O_1034,N_23206,N_23200);
or UO_1035 (O_1035,N_22795,N_23866);
nand UO_1036 (O_1036,N_20303,N_19310);
and UO_1037 (O_1037,N_19039,N_21743);
xor UO_1038 (O_1038,N_19828,N_21899);
or UO_1039 (O_1039,N_22927,N_19859);
nor UO_1040 (O_1040,N_19689,N_24296);
and UO_1041 (O_1041,N_21390,N_21719);
or UO_1042 (O_1042,N_20758,N_20060);
and UO_1043 (O_1043,N_19572,N_21973);
xor UO_1044 (O_1044,N_18999,N_19167);
or UO_1045 (O_1045,N_18989,N_20734);
xnor UO_1046 (O_1046,N_21372,N_23243);
nor UO_1047 (O_1047,N_23839,N_20288);
or UO_1048 (O_1048,N_20047,N_23234);
nor UO_1049 (O_1049,N_21044,N_19492);
nand UO_1050 (O_1050,N_23535,N_22290);
nor UO_1051 (O_1051,N_23152,N_20849);
nand UO_1052 (O_1052,N_21909,N_20764);
nor UO_1053 (O_1053,N_20495,N_24309);
xnor UO_1054 (O_1054,N_23209,N_24409);
or UO_1055 (O_1055,N_21244,N_20293);
nor UO_1056 (O_1056,N_23541,N_23645);
nand UO_1057 (O_1057,N_23737,N_24145);
nor UO_1058 (O_1058,N_19718,N_22255);
nor UO_1059 (O_1059,N_24420,N_22815);
xnor UO_1060 (O_1060,N_23323,N_20517);
or UO_1061 (O_1061,N_20347,N_21364);
or UO_1062 (O_1062,N_24254,N_19814);
xnor UO_1063 (O_1063,N_22490,N_22852);
and UO_1064 (O_1064,N_22721,N_20890);
or UO_1065 (O_1065,N_23259,N_20618);
or UO_1066 (O_1066,N_23067,N_24772);
nand UO_1067 (O_1067,N_21903,N_21457);
nor UO_1068 (O_1068,N_24706,N_22066);
xor UO_1069 (O_1069,N_22179,N_24785);
and UO_1070 (O_1070,N_24875,N_24429);
nor UO_1071 (O_1071,N_24973,N_24386);
nor UO_1072 (O_1072,N_23361,N_21359);
nand UO_1073 (O_1073,N_23934,N_23782);
nor UO_1074 (O_1074,N_19362,N_18998);
or UO_1075 (O_1075,N_22893,N_23652);
nor UO_1076 (O_1076,N_20280,N_19314);
xor UO_1077 (O_1077,N_21245,N_20052);
and UO_1078 (O_1078,N_23682,N_24360);
xor UO_1079 (O_1079,N_24611,N_22694);
xor UO_1080 (O_1080,N_19832,N_24191);
and UO_1081 (O_1081,N_20301,N_23852);
nand UO_1082 (O_1082,N_23983,N_22888);
nand UO_1083 (O_1083,N_21333,N_20521);
nand UO_1084 (O_1084,N_21383,N_18763);
nor UO_1085 (O_1085,N_24882,N_20559);
nor UO_1086 (O_1086,N_22000,N_18768);
nand UO_1087 (O_1087,N_20265,N_23394);
xor UO_1088 (O_1088,N_20388,N_24503);
or UO_1089 (O_1089,N_18900,N_24445);
nand UO_1090 (O_1090,N_19809,N_20320);
nor UO_1091 (O_1091,N_19502,N_23889);
or UO_1092 (O_1092,N_24034,N_24097);
or UO_1093 (O_1093,N_21326,N_23311);
nand UO_1094 (O_1094,N_20193,N_24001);
nor UO_1095 (O_1095,N_24573,N_23892);
xnor UO_1096 (O_1096,N_20980,N_21034);
nor UO_1097 (O_1097,N_21484,N_22911);
and UO_1098 (O_1098,N_24687,N_19108);
nand UO_1099 (O_1099,N_22431,N_24853);
nand UO_1100 (O_1100,N_21161,N_23489);
and UO_1101 (O_1101,N_20459,N_22399);
or UO_1102 (O_1102,N_18912,N_20378);
and UO_1103 (O_1103,N_23387,N_23715);
xnor UO_1104 (O_1104,N_24572,N_21007);
nor UO_1105 (O_1105,N_20908,N_18880);
nor UO_1106 (O_1106,N_23318,N_20830);
xnor UO_1107 (O_1107,N_23691,N_24401);
nand UO_1108 (O_1108,N_24974,N_21394);
xnor UO_1109 (O_1109,N_21192,N_23153);
or UO_1110 (O_1110,N_20369,N_24196);
or UO_1111 (O_1111,N_22873,N_24356);
xor UO_1112 (O_1112,N_21157,N_19620);
and UO_1113 (O_1113,N_24713,N_22596);
and UO_1114 (O_1114,N_21834,N_22286);
xnor UO_1115 (O_1115,N_22123,N_19044);
or UO_1116 (O_1116,N_24830,N_23957);
and UO_1117 (O_1117,N_23864,N_24161);
nor UO_1118 (O_1118,N_24448,N_21278);
and UO_1119 (O_1119,N_21257,N_20965);
or UO_1120 (O_1120,N_20608,N_21881);
nand UO_1121 (O_1121,N_24274,N_22890);
and UO_1122 (O_1122,N_19580,N_22134);
nand UO_1123 (O_1123,N_24336,N_20356);
or UO_1124 (O_1124,N_19586,N_24959);
nand UO_1125 (O_1125,N_19023,N_23674);
nand UO_1126 (O_1126,N_20992,N_23121);
xor UO_1127 (O_1127,N_24266,N_22288);
nand UO_1128 (O_1128,N_20089,N_22672);
nor UO_1129 (O_1129,N_20866,N_24157);
and UO_1130 (O_1130,N_20714,N_19868);
and UO_1131 (O_1131,N_19996,N_20719);
nor UO_1132 (O_1132,N_21651,N_24560);
nand UO_1133 (O_1133,N_24084,N_23580);
xnor UO_1134 (O_1134,N_20829,N_18961);
and UO_1135 (O_1135,N_20016,N_23281);
nand UO_1136 (O_1136,N_24652,N_23885);
nand UO_1137 (O_1137,N_24112,N_24067);
or UO_1138 (O_1138,N_24748,N_22094);
xor UO_1139 (O_1139,N_20698,N_23163);
xor UO_1140 (O_1140,N_24938,N_23441);
or UO_1141 (O_1141,N_21321,N_24335);
nor UO_1142 (O_1142,N_18788,N_21149);
xnor UO_1143 (O_1143,N_20672,N_20661);
nor UO_1144 (O_1144,N_21707,N_19425);
or UO_1145 (O_1145,N_20036,N_24980);
or UO_1146 (O_1146,N_19923,N_21347);
nand UO_1147 (O_1147,N_19485,N_18992);
xor UO_1148 (O_1148,N_21686,N_20868);
xnor UO_1149 (O_1149,N_23956,N_24662);
and UO_1150 (O_1150,N_23416,N_23261);
or UO_1151 (O_1151,N_23633,N_20349);
nand UO_1152 (O_1152,N_23224,N_19306);
nor UO_1153 (O_1153,N_22545,N_21520);
xnor UO_1154 (O_1154,N_24522,N_21554);
or UO_1155 (O_1155,N_21074,N_20944);
nor UO_1156 (O_1156,N_23062,N_19217);
nand UO_1157 (O_1157,N_19423,N_22574);
nand UO_1158 (O_1158,N_18951,N_20791);
nand UO_1159 (O_1159,N_23352,N_23974);
nand UO_1160 (O_1160,N_18919,N_21275);
xor UO_1161 (O_1161,N_19826,N_19640);
nor UO_1162 (O_1162,N_22918,N_21350);
and UO_1163 (O_1163,N_21122,N_21258);
and UO_1164 (O_1164,N_19290,N_20776);
xor UO_1165 (O_1165,N_20233,N_21179);
xor UO_1166 (O_1166,N_24241,N_22270);
xor UO_1167 (O_1167,N_24887,N_20030);
nand UO_1168 (O_1168,N_22874,N_21970);
and UO_1169 (O_1169,N_19211,N_22617);
or UO_1170 (O_1170,N_21416,N_18771);
and UO_1171 (O_1171,N_19220,N_20259);
nand UO_1172 (O_1172,N_22214,N_21230);
xor UO_1173 (O_1173,N_22108,N_21614);
xor UO_1174 (O_1174,N_21106,N_19838);
xnor UO_1175 (O_1175,N_20154,N_22634);
nor UO_1176 (O_1176,N_18811,N_24263);
nor UO_1177 (O_1177,N_23278,N_18905);
and UO_1178 (O_1178,N_19109,N_24594);
or UO_1179 (O_1179,N_20851,N_20697);
or UO_1180 (O_1180,N_21855,N_24464);
or UO_1181 (O_1181,N_23193,N_21108);
and UO_1182 (O_1182,N_21136,N_23292);
or UO_1183 (O_1183,N_22711,N_22332);
nor UO_1184 (O_1184,N_24549,N_24641);
xor UO_1185 (O_1185,N_19714,N_19928);
xnor UO_1186 (O_1186,N_20475,N_21815);
or UO_1187 (O_1187,N_20705,N_21101);
nand UO_1188 (O_1188,N_22428,N_23940);
and UO_1189 (O_1189,N_20969,N_19244);
and UO_1190 (O_1190,N_21900,N_23858);
or UO_1191 (O_1191,N_23810,N_22738);
nor UO_1192 (O_1192,N_24056,N_24597);
xor UO_1193 (O_1193,N_23673,N_24037);
nand UO_1194 (O_1194,N_22754,N_21426);
nand UO_1195 (O_1195,N_23271,N_21311);
nand UO_1196 (O_1196,N_23649,N_22763);
or UO_1197 (O_1197,N_21260,N_20799);
xor UO_1198 (O_1198,N_19336,N_19180);
xor UO_1199 (O_1199,N_22823,N_23925);
or UO_1200 (O_1200,N_23799,N_24538);
or UO_1201 (O_1201,N_19342,N_20326);
nor UO_1202 (O_1202,N_19795,N_23822);
nand UO_1203 (O_1203,N_21103,N_22840);
and UO_1204 (O_1204,N_22817,N_23755);
nor UO_1205 (O_1205,N_22273,N_22593);
and UO_1206 (O_1206,N_22326,N_18899);
nand UO_1207 (O_1207,N_22037,N_23141);
nor UO_1208 (O_1208,N_24756,N_19376);
xor UO_1209 (O_1209,N_22602,N_24892);
and UO_1210 (O_1210,N_22659,N_23507);
nor UO_1211 (O_1211,N_21545,N_24603);
or UO_1212 (O_1212,N_24878,N_23676);
xor UO_1213 (O_1213,N_23753,N_21621);
nor UO_1214 (O_1214,N_23167,N_24646);
and UO_1215 (O_1215,N_19788,N_24369);
xnor UO_1216 (O_1216,N_24691,N_24248);
nor UO_1217 (O_1217,N_21288,N_20066);
nor UO_1218 (O_1218,N_24197,N_19721);
nor UO_1219 (O_1219,N_22400,N_20321);
and UO_1220 (O_1220,N_22580,N_19380);
xor UO_1221 (O_1221,N_18921,N_20772);
and UO_1222 (O_1222,N_22880,N_22046);
nor UO_1223 (O_1223,N_19273,N_18958);
nor UO_1224 (O_1224,N_19680,N_20860);
or UO_1225 (O_1225,N_24801,N_22667);
xor UO_1226 (O_1226,N_19534,N_22161);
xnor UO_1227 (O_1227,N_19878,N_20820);
nand UO_1228 (O_1228,N_19912,N_23739);
nand UO_1229 (O_1229,N_22516,N_19232);
and UO_1230 (O_1230,N_21287,N_23905);
nand UO_1231 (O_1231,N_19319,N_22843);
or UO_1232 (O_1232,N_19117,N_21452);
and UO_1233 (O_1233,N_21189,N_23279);
and UO_1234 (O_1234,N_22055,N_23973);
nor UO_1235 (O_1235,N_19114,N_23054);
nor UO_1236 (O_1236,N_24477,N_19882);
and UO_1237 (O_1237,N_18787,N_24970);
nor UO_1238 (O_1238,N_23142,N_19699);
nand UO_1239 (O_1239,N_23037,N_20339);
or UO_1240 (O_1240,N_19441,N_19287);
nor UO_1241 (O_1241,N_24550,N_19242);
and UO_1242 (O_1242,N_20189,N_23072);
nand UO_1243 (O_1243,N_20465,N_23664);
and UO_1244 (O_1244,N_19248,N_21387);
xor UO_1245 (O_1245,N_23143,N_22938);
or UO_1246 (O_1246,N_21993,N_19822);
and UO_1247 (O_1247,N_18964,N_23237);
nor UO_1248 (O_1248,N_23965,N_22159);
xor UO_1249 (O_1249,N_21676,N_20507);
and UO_1250 (O_1250,N_19847,N_19454);
nand UO_1251 (O_1251,N_24966,N_24381);
nand UO_1252 (O_1252,N_18904,N_23837);
and UO_1253 (O_1253,N_20942,N_21981);
or UO_1254 (O_1254,N_22618,N_22106);
nor UO_1255 (O_1255,N_20895,N_24181);
nand UO_1256 (O_1256,N_21665,N_23995);
and UO_1257 (O_1257,N_24912,N_23051);
and UO_1258 (O_1258,N_21148,N_21866);
nand UO_1259 (O_1259,N_23210,N_22200);
or UO_1260 (O_1260,N_19436,N_20262);
nand UO_1261 (O_1261,N_21907,N_19724);
xor UO_1262 (O_1262,N_21343,N_23783);
or UO_1263 (O_1263,N_19612,N_20496);
nand UO_1264 (O_1264,N_19183,N_22633);
nand UO_1265 (O_1265,N_19663,N_23941);
or UO_1266 (O_1266,N_20656,N_24224);
xor UO_1267 (O_1267,N_24715,N_21606);
and UO_1268 (O_1268,N_22396,N_19077);
or UO_1269 (O_1269,N_19902,N_21796);
nand UO_1270 (O_1270,N_19240,N_24028);
nand UO_1271 (O_1271,N_22191,N_24870);
and UO_1272 (O_1272,N_19582,N_24510);
xor UO_1273 (O_1273,N_24513,N_22924);
or UO_1274 (O_1274,N_23928,N_18757);
nand UO_1275 (O_1275,N_18764,N_19345);
or UO_1276 (O_1276,N_22299,N_22065);
nor UO_1277 (O_1277,N_20518,N_21558);
nand UO_1278 (O_1278,N_18959,N_21218);
and UO_1279 (O_1279,N_24625,N_20638);
or UO_1280 (O_1280,N_24317,N_20770);
and UO_1281 (O_1281,N_19266,N_20013);
and UO_1282 (O_1282,N_21677,N_24582);
and UO_1283 (O_1283,N_23076,N_22798);
nor UO_1284 (O_1284,N_24433,N_22140);
and UO_1285 (O_1285,N_19961,N_18901);
or UO_1286 (O_1286,N_21891,N_23551);
nor UO_1287 (O_1287,N_24118,N_24552);
or UO_1288 (O_1288,N_24585,N_24695);
and UO_1289 (O_1289,N_22230,N_22408);
xnor UO_1290 (O_1290,N_23556,N_21636);
nand UO_1291 (O_1291,N_18830,N_21642);
and UO_1292 (O_1292,N_22473,N_23423);
xnor UO_1293 (O_1293,N_21726,N_19499);
and UO_1294 (O_1294,N_23106,N_23906);
or UO_1295 (O_1295,N_22583,N_23630);
xnor UO_1296 (O_1296,N_23365,N_20839);
xnor UO_1297 (O_1297,N_21956,N_24327);
nor UO_1298 (O_1298,N_19286,N_19162);
nand UO_1299 (O_1299,N_18942,N_22045);
nor UO_1300 (O_1300,N_22100,N_21872);
nor UO_1301 (O_1301,N_21679,N_24443);
xnor UO_1302 (O_1302,N_24836,N_23483);
xor UO_1303 (O_1303,N_24655,N_20582);
nand UO_1304 (O_1304,N_22418,N_24901);
xor UO_1305 (O_1305,N_19696,N_23643);
and UO_1306 (O_1306,N_23332,N_23809);
and UO_1307 (O_1307,N_24342,N_23653);
xor UO_1308 (O_1308,N_19017,N_21859);
nor UO_1309 (O_1309,N_19315,N_20333);
or UO_1310 (O_1310,N_20707,N_20844);
nor UO_1311 (O_1311,N_19739,N_23183);
or UO_1312 (O_1312,N_24111,N_19567);
and UO_1313 (O_1313,N_23921,N_19272);
xnor UO_1314 (O_1314,N_23620,N_20501);
or UO_1315 (O_1315,N_21213,N_19416);
and UO_1316 (O_1316,N_24660,N_22061);
or UO_1317 (O_1317,N_19644,N_21022);
or UO_1318 (O_1318,N_19284,N_20583);
or UO_1319 (O_1319,N_19712,N_21132);
xnor UO_1320 (O_1320,N_21843,N_21812);
xor UO_1321 (O_1321,N_24983,N_19226);
xor UO_1322 (O_1322,N_24858,N_20282);
xor UO_1323 (O_1323,N_19071,N_22068);
and UO_1324 (O_1324,N_19688,N_23086);
or UO_1325 (O_1325,N_18930,N_24575);
xor UO_1326 (O_1326,N_23930,N_22250);
nor UO_1327 (O_1327,N_22345,N_20205);
and UO_1328 (O_1328,N_24209,N_20929);
or UO_1329 (O_1329,N_21134,N_19647);
xnor UO_1330 (O_1330,N_20357,N_19587);
and UO_1331 (O_1331,N_23806,N_18923);
nand UO_1332 (O_1332,N_19134,N_18800);
xor UO_1333 (O_1333,N_19098,N_22917);
or UO_1334 (O_1334,N_19019,N_21120);
nand UO_1335 (O_1335,N_24565,N_23485);
or UO_1336 (O_1336,N_24339,N_20744);
nand UO_1337 (O_1337,N_18897,N_22023);
and UO_1338 (O_1338,N_20928,N_24278);
xnor UO_1339 (O_1339,N_21756,N_23695);
or UO_1340 (O_1340,N_20576,N_22811);
and UO_1341 (O_1341,N_20162,N_23654);
nand UO_1342 (O_1342,N_23275,N_22879);
nor UO_1343 (O_1343,N_20039,N_24880);
or UO_1344 (O_1344,N_22898,N_23041);
nor UO_1345 (O_1345,N_21191,N_24009);
nand UO_1346 (O_1346,N_23873,N_22434);
or UO_1347 (O_1347,N_23448,N_24222);
nand UO_1348 (O_1348,N_22358,N_23087);
nor UO_1349 (O_1349,N_23853,N_22532);
and UO_1350 (O_1350,N_20567,N_21794);
xor UO_1351 (O_1351,N_19837,N_21570);
xor UO_1352 (O_1352,N_24505,N_19218);
or UO_1353 (O_1353,N_19783,N_19005);
nor UO_1354 (O_1354,N_23848,N_22499);
nor UO_1355 (O_1355,N_20241,N_24321);
and UO_1356 (O_1356,N_24020,N_24159);
xor UO_1357 (O_1357,N_21653,N_21168);
nor UO_1358 (O_1358,N_20225,N_22069);
nor UO_1359 (O_1359,N_18851,N_24839);
xnor UO_1360 (O_1360,N_24412,N_23574);
nand UO_1361 (O_1361,N_24123,N_22474);
and UO_1362 (O_1362,N_20430,N_23807);
or UO_1363 (O_1363,N_22592,N_19762);
and UO_1364 (O_1364,N_22359,N_22261);
nand UO_1365 (O_1365,N_24803,N_24364);
xnor UO_1366 (O_1366,N_23665,N_21337);
xor UO_1367 (O_1367,N_22525,N_20649);
xnor UO_1368 (O_1368,N_23487,N_21650);
nor UO_1369 (O_1369,N_24916,N_21069);
xnor UO_1370 (O_1370,N_22022,N_23248);
xor UO_1371 (O_1371,N_24162,N_23675);
nor UO_1372 (O_1372,N_18752,N_23626);
and UO_1373 (O_1373,N_24098,N_24659);
nand UO_1374 (O_1374,N_23414,N_21392);
and UO_1375 (O_1375,N_20848,N_23424);
nor UO_1376 (O_1376,N_19453,N_21174);
and UO_1377 (O_1377,N_19825,N_22578);
nor UO_1378 (O_1378,N_21580,N_22702);
and UO_1379 (O_1379,N_22740,N_21163);
or UO_1380 (O_1380,N_24265,N_24267);
nor UO_1381 (O_1381,N_24027,N_19648);
or UO_1382 (O_1382,N_20471,N_22343);
nand UO_1383 (O_1383,N_18844,N_18862);
and UO_1384 (O_1384,N_23390,N_19970);
and UO_1385 (O_1385,N_20615,N_20100);
xnor UO_1386 (O_1386,N_20117,N_21215);
or UO_1387 (O_1387,N_22563,N_22331);
nand UO_1388 (O_1388,N_18909,N_20574);
xor UO_1389 (O_1389,N_22008,N_20872);
nand UO_1390 (O_1390,N_22327,N_20139);
or UO_1391 (O_1391,N_20544,N_24352);
nor UO_1392 (O_1392,N_20626,N_24470);
nor UO_1393 (O_1393,N_22476,N_24345);
nor UO_1394 (O_1394,N_21105,N_22084);
xnor UO_1395 (O_1395,N_21293,N_24855);
or UO_1396 (O_1396,N_24786,N_22931);
nor UO_1397 (O_1397,N_21316,N_19845);
or UO_1398 (O_1398,N_24173,N_23052);
or UO_1399 (O_1399,N_21323,N_23227);
xnor UO_1400 (O_1400,N_24908,N_24291);
nor UO_1401 (O_1401,N_18853,N_21305);
and UO_1402 (O_1402,N_23160,N_23217);
xor UO_1403 (O_1403,N_21483,N_23602);
nor UO_1404 (O_1404,N_20514,N_19609);
nor UO_1405 (O_1405,N_21062,N_24663);
or UO_1406 (O_1406,N_21927,N_19083);
nor UO_1407 (O_1407,N_22912,N_19715);
xor UO_1408 (O_1408,N_19546,N_23796);
nand UO_1409 (O_1409,N_20335,N_22887);
and UO_1410 (O_1410,N_20781,N_18750);
nand UO_1411 (O_1411,N_23298,N_19155);
xnor UO_1412 (O_1412,N_22300,N_18935);
nor UO_1413 (O_1413,N_23123,N_22845);
nand UO_1414 (O_1414,N_24929,N_22180);
nor UO_1415 (O_1415,N_19741,N_22044);
xnor UO_1416 (O_1416,N_24814,N_20864);
nand UO_1417 (O_1417,N_20274,N_20861);
nor UO_1418 (O_1418,N_22130,N_19678);
and UO_1419 (O_1419,N_20254,N_22098);
or UO_1420 (O_1420,N_24039,N_24405);
nand UO_1421 (O_1421,N_23088,N_19941);
nand UO_1422 (O_1422,N_18976,N_22146);
xor UO_1423 (O_1423,N_20256,N_22350);
nor UO_1424 (O_1424,N_19359,N_18916);
xor UO_1425 (O_1425,N_20253,N_20370);
or UO_1426 (O_1426,N_18831,N_23058);
and UO_1427 (O_1427,N_24081,N_22223);
xor UO_1428 (O_1428,N_20255,N_21864);
nor UO_1429 (O_1429,N_20034,N_24866);
or UO_1430 (O_1430,N_20355,N_24046);
xnor UO_1431 (O_1431,N_24313,N_22074);
nor UO_1432 (O_1432,N_22625,N_19026);
and UO_1433 (O_1433,N_19865,N_21789);
nand UO_1434 (O_1434,N_23980,N_21079);
xnor UO_1435 (O_1435,N_23523,N_24220);
and UO_1436 (O_1436,N_20769,N_19942);
and UO_1437 (O_1437,N_21227,N_22433);
nand UO_1438 (O_1438,N_22278,N_19641);
xnor UO_1439 (O_1439,N_20316,N_20096);
xnor UO_1440 (O_1440,N_20989,N_19743);
nand UO_1441 (O_1441,N_21711,N_22051);
and UO_1442 (O_1442,N_24877,N_21423);
nor UO_1443 (O_1443,N_19229,N_22226);
nand UO_1444 (O_1444,N_24979,N_22571);
and UO_1445 (O_1445,N_21934,N_20155);
and UO_1446 (O_1446,N_22190,N_20603);
or UO_1447 (O_1447,N_21562,N_20945);
nor UO_1448 (O_1448,N_21111,N_22365);
or UO_1449 (O_1449,N_24670,N_20796);
or UO_1450 (O_1450,N_20962,N_23571);
nand UO_1451 (O_1451,N_22351,N_18829);
xor UO_1452 (O_1452,N_21923,N_24349);
nand UO_1453 (O_1453,N_24195,N_22312);
nand UO_1454 (O_1454,N_24140,N_19122);
and UO_1455 (O_1455,N_24202,N_24627);
or UO_1456 (O_1456,N_18834,N_20453);
nor UO_1457 (O_1457,N_24924,N_18852);
or UO_1458 (O_1458,N_19069,N_19940);
xnor UO_1459 (O_1459,N_21433,N_20134);
nor UO_1460 (O_1460,N_23340,N_23619);
and UO_1461 (O_1461,N_20645,N_21714);
nand UO_1462 (O_1462,N_21770,N_19245);
and UO_1463 (O_1463,N_23018,N_23346);
nor UO_1464 (O_1464,N_24811,N_23439);
and UO_1465 (O_1465,N_24468,N_23302);
xor UO_1466 (O_1466,N_21481,N_21695);
xnor UO_1467 (O_1467,N_22310,N_22753);
nor UO_1468 (O_1468,N_20454,N_19706);
xor UO_1469 (O_1469,N_18969,N_21962);
xor UO_1470 (O_1470,N_22324,N_24175);
nor UO_1471 (O_1471,N_22818,N_20787);
nor UO_1472 (O_1472,N_20437,N_22964);
xor UO_1473 (O_1473,N_21455,N_19096);
nand UO_1474 (O_1474,N_23050,N_20408);
and UO_1475 (O_1475,N_24302,N_20859);
xnor UO_1476 (O_1476,N_20431,N_20401);
or UO_1477 (O_1477,N_18770,N_24775);
and UO_1478 (O_1478,N_24680,N_21968);
xor UO_1479 (O_1479,N_19733,N_19870);
nor UO_1480 (O_1480,N_20669,N_19049);
nand UO_1481 (O_1481,N_21166,N_20873);
xnor UO_1482 (O_1482,N_21831,N_20800);
or UO_1483 (O_1483,N_21119,N_24947);
xor UO_1484 (O_1484,N_22568,N_23617);
nor UO_1485 (O_1485,N_20414,N_23598);
and UO_1486 (O_1486,N_19082,N_24253);
and UO_1487 (O_1487,N_21202,N_21206);
or UO_1488 (O_1488,N_24638,N_22141);
nand UO_1489 (O_1489,N_22518,N_21996);
xnor UO_1490 (O_1490,N_22523,N_21581);
or UO_1491 (O_1491,N_24618,N_22994);
nand UO_1492 (O_1492,N_22967,N_21867);
nor UO_1493 (O_1493,N_22003,N_20551);
and UO_1494 (O_1494,N_24066,N_20504);
xnor UO_1495 (O_1495,N_21753,N_21097);
nand UO_1496 (O_1496,N_18980,N_22600);
and UO_1497 (O_1497,N_22096,N_22886);
or UO_1498 (O_1498,N_18823,N_19554);
nor UO_1499 (O_1499,N_23263,N_19412);
or UO_1500 (O_1500,N_22060,N_22204);
nand UO_1501 (O_1501,N_23651,N_21599);
xnor UO_1502 (O_1502,N_22072,N_19381);
and UO_1503 (O_1503,N_20542,N_20898);
nor UO_1504 (O_1504,N_21953,N_23952);
nand UO_1505 (O_1505,N_22834,N_24178);
nor UO_1506 (O_1506,N_20695,N_23460);
nor UO_1507 (O_1507,N_21664,N_23687);
nor UO_1508 (O_1508,N_24524,N_24888);
or UO_1509 (O_1509,N_24697,N_22599);
nand UO_1510 (O_1510,N_24788,N_19491);
and UO_1511 (O_1511,N_22567,N_22416);
xor UO_1512 (O_1512,N_20099,N_22786);
xor UO_1513 (O_1513,N_20783,N_18995);
and UO_1514 (O_1514,N_23034,N_24862);
or UO_1515 (O_1515,N_21164,N_22732);
nor UO_1516 (O_1516,N_22851,N_22470);
or UO_1517 (O_1517,N_21479,N_21035);
nor UO_1518 (O_1518,N_22603,N_21922);
and UO_1519 (O_1519,N_21531,N_21977);
nand UO_1520 (O_1520,N_19603,N_24891);
or UO_1521 (O_1521,N_23954,N_20009);
nand UO_1522 (O_1522,N_20725,N_22415);
and UO_1523 (O_1523,N_23110,N_24135);
and UO_1524 (O_1524,N_24499,N_21528);
nor UO_1525 (O_1525,N_20950,N_19779);
or UO_1526 (O_1526,N_24029,N_18807);
or UO_1527 (O_1527,N_22784,N_22734);
or UO_1528 (O_1528,N_19785,N_22566);
or UO_1529 (O_1529,N_21393,N_21470);
or UO_1530 (O_1530,N_19626,N_22090);
nor UO_1531 (O_1531,N_21376,N_19702);
and UO_1532 (O_1532,N_21137,N_21930);
nand UO_1533 (O_1533,N_23748,N_23468);
nor UO_1534 (O_1534,N_22466,N_23353);
and UO_1535 (O_1535,N_20073,N_19694);
xnor UO_1536 (O_1536,N_21296,N_20438);
and UO_1537 (O_1537,N_24396,N_19209);
nand UO_1538 (O_1538,N_24904,N_24516);
and UO_1539 (O_1539,N_19818,N_23157);
xnor UO_1540 (O_1540,N_22389,N_24032);
or UO_1541 (O_1541,N_19192,N_22392);
or UO_1542 (O_1542,N_23176,N_24744);
and UO_1543 (O_1543,N_24894,N_23843);
xor UO_1544 (O_1544,N_19805,N_19854);
nor UO_1545 (O_1545,N_21905,N_22089);
or UO_1546 (O_1546,N_24599,N_20183);
xor UO_1547 (O_1547,N_18838,N_21880);
nand UO_1548 (O_1548,N_20743,N_22519);
and UO_1549 (O_1549,N_24014,N_20472);
nor UO_1550 (O_1550,N_20230,N_21385);
xor UO_1551 (O_1551,N_22352,N_22496);
and UO_1552 (O_1552,N_20217,N_22426);
nor UO_1553 (O_1553,N_24678,N_24355);
or UO_1554 (O_1554,N_18847,N_23449);
xor UO_1555 (O_1555,N_23391,N_19185);
nor UO_1556 (O_1556,N_20662,N_18937);
and UO_1557 (O_1557,N_19343,N_22461);
nor UO_1558 (O_1558,N_23735,N_22082);
and UO_1559 (O_1559,N_21522,N_23168);
nor UO_1560 (O_1560,N_23927,N_22318);
xor UO_1561 (O_1561,N_21893,N_24012);
nand UO_1562 (O_1562,N_19035,N_21915);
xor UO_1563 (O_1563,N_19074,N_23306);
or UO_1564 (O_1564,N_24163,N_23473);
or UO_1565 (O_1565,N_24006,N_18881);
xor UO_1566 (O_1566,N_23527,N_24235);
or UO_1567 (O_1567,N_23074,N_20751);
nor UO_1568 (O_1568,N_23984,N_23849);
nor UO_1569 (O_1569,N_22680,N_19449);
or UO_1570 (O_1570,N_21109,N_20308);
xor UO_1571 (O_1571,N_23190,N_19860);
and UO_1572 (O_1572,N_23218,N_18886);
nor UO_1573 (O_1573,N_22564,N_20809);
or UO_1574 (O_1574,N_19427,N_23525);
xnor UO_1575 (O_1575,N_21353,N_19780);
and UO_1576 (O_1576,N_19405,N_20831);
and UO_1577 (O_1577,N_24456,N_22302);
and UO_1578 (O_1578,N_19927,N_24466);
nor UO_1579 (O_1579,N_24488,N_20021);
nand UO_1580 (O_1580,N_23614,N_24790);
or UO_1581 (O_1581,N_21641,N_22391);
nand UO_1582 (O_1582,N_23148,N_24911);
nand UO_1583 (O_1583,N_23309,N_24626);
and UO_1584 (O_1584,N_19130,N_22605);
xor UO_1585 (O_1585,N_21352,N_23877);
or UO_1586 (O_1586,N_18973,N_23258);
and UO_1587 (O_1587,N_24925,N_19007);
nand UO_1588 (O_1588,N_19894,N_24343);
and UO_1589 (O_1589,N_22207,N_19520);
or UO_1590 (O_1590,N_20245,N_20880);
xor UO_1591 (O_1591,N_24358,N_20903);
or UO_1592 (O_1592,N_21322,N_21648);
xor UO_1593 (O_1593,N_24167,N_21889);
and UO_1594 (O_1594,N_19981,N_22797);
xnor UO_1595 (O_1595,N_21949,N_22807);
xor UO_1596 (O_1596,N_20145,N_19542);
nor UO_1597 (O_1597,N_24529,N_22512);
xor UO_1598 (O_1598,N_24605,N_24563);
nor UO_1599 (O_1599,N_21366,N_20605);
and UO_1600 (O_1600,N_20109,N_24082);
xor UO_1601 (O_1601,N_24287,N_24385);
nor UO_1602 (O_1602,N_18766,N_20195);
nor UO_1603 (O_1603,N_23445,N_19852);
nor UO_1604 (O_1604,N_19204,N_21186);
nor UO_1605 (O_1605,N_23740,N_21282);
nand UO_1606 (O_1606,N_20792,N_22637);
nor UO_1607 (O_1607,N_19149,N_21420);
xnor UO_1608 (O_1608,N_20668,N_21667);
xor UO_1609 (O_1609,N_21771,N_20592);
or UO_1610 (O_1610,N_20315,N_24437);
or UO_1611 (O_1611,N_23512,N_22594);
and UO_1612 (O_1612,N_20524,N_20266);
and UO_1613 (O_1613,N_20541,N_19014);
and UO_1614 (O_1614,N_22275,N_24561);
or UO_1615 (O_1615,N_20072,N_19301);
nor UO_1616 (O_1616,N_20957,N_20892);
xnor UO_1617 (O_1617,N_21150,N_23662);
or UO_1618 (O_1618,N_20232,N_24955);
or UO_1619 (O_1619,N_21865,N_20063);
and UO_1620 (O_1620,N_22531,N_24954);
or UO_1621 (O_1621,N_21758,N_23982);
xnor UO_1622 (O_1622,N_19364,N_23154);
nand UO_1623 (O_1623,N_20529,N_21207);
nor UO_1624 (O_1624,N_20987,N_19980);
nor UO_1625 (O_1625,N_19361,N_22367);
nand UO_1626 (O_1626,N_21113,N_24189);
nand UO_1627 (O_1627,N_21814,N_20564);
xor UO_1628 (O_1628,N_22010,N_21369);
or UO_1629 (O_1629,N_24094,N_21870);
nand UO_1630 (O_1630,N_21781,N_19512);
and UO_1631 (O_1631,N_20958,N_20204);
xor UO_1632 (O_1632,N_23842,N_22201);
and UO_1633 (O_1633,N_23231,N_22104);
or UO_1634 (O_1634,N_24632,N_20130);
and UO_1635 (O_1635,N_20001,N_19729);
or UO_1636 (O_1636,N_23959,N_24079);
or UO_1637 (O_1637,N_19864,N_24797);
xor UO_1638 (O_1638,N_22264,N_22333);
and UO_1639 (O_1639,N_21976,N_20675);
and UO_1640 (O_1640,N_23033,N_19914);
and UO_1641 (O_1641,N_20432,N_20917);
nand UO_1642 (O_1642,N_20970,N_20019);
nand UO_1643 (O_1643,N_23186,N_19010);
nor UO_1644 (O_1644,N_19659,N_19473);
xor UO_1645 (O_1645,N_21429,N_21185);
nand UO_1646 (O_1646,N_24308,N_20835);
xor UO_1647 (O_1647,N_24854,N_22759);
nand UO_1648 (O_1648,N_22989,N_19041);
or UO_1649 (O_1649,N_20064,N_20123);
nor UO_1650 (O_1650,N_21624,N_23308);
and UO_1651 (O_1651,N_19767,N_22597);
nor UO_1652 (O_1652,N_21361,N_23513);
and UO_1653 (O_1653,N_19462,N_19210);
and UO_1654 (O_1654,N_21963,N_18925);
and UO_1655 (O_1655,N_20884,N_24941);
or UO_1656 (O_1656,N_24885,N_23285);
xnor UO_1657 (O_1657,N_24168,N_21869);
or UO_1658 (O_1658,N_24731,N_19170);
xor UO_1659 (O_1659,N_20441,N_19255);
and UO_1660 (O_1660,N_21055,N_24720);
xnor UO_1661 (O_1661,N_20137,N_19602);
or UO_1662 (O_1662,N_24666,N_20240);
xnor UO_1663 (O_1663,N_21848,N_21582);
xor UO_1664 (O_1664,N_24832,N_18836);
and UO_1665 (O_1665,N_20680,N_20380);
or UO_1666 (O_1666,N_21941,N_23500);
xor UO_1667 (O_1667,N_23039,N_20359);
xnor UO_1668 (O_1668,N_24121,N_19685);
nor UO_1669 (O_1669,N_21896,N_22157);
nor UO_1670 (O_1670,N_20511,N_21039);
and UO_1671 (O_1671,N_19812,N_22079);
and UO_1672 (O_1672,N_24763,N_21681);
xnor UO_1673 (O_1673,N_24504,N_21440);
or UO_1674 (O_1674,N_19103,N_23199);
or UO_1675 (O_1675,N_23886,N_22472);
and UO_1676 (O_1676,N_24229,N_19819);
and UO_1677 (O_1677,N_19469,N_23108);
and UO_1678 (O_1678,N_19953,N_23085);
or UO_1679 (O_1679,N_18841,N_19443);
xor UO_1680 (O_1680,N_20625,N_21405);
and UO_1681 (O_1681,N_24155,N_23349);
or UO_1682 (O_1682,N_20294,N_20153);
and UO_1683 (O_1683,N_24393,N_19215);
nor UO_1684 (O_1684,N_22829,N_21351);
and UO_1685 (O_1685,N_23987,N_21846);
nor UO_1686 (O_1686,N_21118,N_22624);
and UO_1687 (O_1687,N_20126,N_21271);
or UO_1688 (O_1688,N_19605,N_24808);
and UO_1689 (O_1689,N_24787,N_19994);
xor UO_1690 (O_1690,N_24570,N_21335);
nand UO_1691 (O_1691,N_18939,N_21928);
xnor UO_1692 (O_1692,N_19031,N_22077);
or UO_1693 (O_1693,N_22348,N_21243);
nand UO_1694 (O_1694,N_22781,N_18822);
nor UO_1695 (O_1695,N_22524,N_21308);
nand UO_1696 (O_1696,N_21836,N_19801);
nor UO_1697 (O_1697,N_24506,N_24085);
xor UO_1698 (O_1698,N_19298,N_19296);
and UO_1699 (O_1699,N_24183,N_22144);
and UO_1700 (O_1700,N_23173,N_19545);
nor UO_1701 (O_1701,N_23127,N_22256);
or UO_1702 (O_1702,N_20046,N_22195);
or UO_1703 (O_1703,N_22741,N_23637);
nor UO_1704 (O_1704,N_19992,N_23031);
and UO_1705 (O_1705,N_22953,N_19746);
nand UO_1706 (O_1706,N_22552,N_20897);
or UO_1707 (O_1707,N_24591,N_18979);
or UO_1708 (O_1708,N_23122,N_22328);
nor UO_1709 (O_1709,N_18795,N_23238);
or UO_1710 (O_1710,N_19262,N_19983);
nand UO_1711 (O_1711,N_19599,N_21858);
or UO_1712 (O_1712,N_22265,N_24218);
or UO_1713 (O_1713,N_24104,N_20270);
nand UO_1714 (O_1714,N_23398,N_23536);
xor UO_1715 (O_1715,N_24813,N_20135);
nor UO_1716 (O_1716,N_24492,N_23762);
nand UO_1717 (O_1717,N_22613,N_20633);
xor UO_1718 (O_1718,N_21742,N_20213);
nor UO_1719 (O_1719,N_24069,N_22027);
or UO_1720 (O_1720,N_21401,N_21421);
nand UO_1721 (O_1721,N_21090,N_22147);
xor UO_1722 (O_1722,N_19768,N_19236);
nand UO_1723 (O_1723,N_20343,N_22925);
nand UO_1724 (O_1724,N_19774,N_22404);
and UO_1725 (O_1725,N_19677,N_20377);
or UO_1726 (O_1726,N_23404,N_19032);
nor UO_1727 (O_1727,N_23369,N_19950);
or UO_1728 (O_1728,N_19682,N_23787);
xor UO_1729 (O_1729,N_20424,N_23812);
and UO_1730 (O_1730,N_21769,N_24606);
or UO_1731 (O_1731,N_20334,N_23427);
and UO_1732 (O_1732,N_21239,N_21525);
nand UO_1733 (O_1733,N_24517,N_23014);
or UO_1734 (O_1734,N_24934,N_21644);
nor UO_1735 (O_1735,N_19571,N_19628);
and UO_1736 (O_1736,N_19945,N_21367);
nand UO_1737 (O_1737,N_21313,N_21153);
xnor UO_1738 (O_1738,N_22390,N_21874);
xnor UO_1739 (O_1739,N_20397,N_19939);
nand UO_1740 (O_1740,N_21647,N_22148);
nand UO_1741 (O_1741,N_19527,N_22364);
nor UO_1742 (O_1742,N_22584,N_22736);
nand UO_1743 (O_1743,N_24969,N_23501);
nor UO_1744 (O_1744,N_23497,N_20666);
and UO_1745 (O_1745,N_24963,N_21523);
nand UO_1746 (O_1746,N_21349,N_20358);
nand UO_1747 (O_1747,N_19317,N_18854);
and UO_1748 (O_1748,N_24127,N_22231);
and UO_1749 (O_1749,N_19804,N_20704);
or UO_1750 (O_1750,N_23282,N_24798);
nand UO_1751 (O_1751,N_22213,N_19615);
and UO_1752 (O_1752,N_22813,N_18755);
or UO_1753 (O_1753,N_23301,N_19464);
nor UO_1754 (O_1754,N_21001,N_24719);
and UO_1755 (O_1755,N_23897,N_24555);
and UO_1756 (O_1756,N_19577,N_21969);
and UO_1757 (O_1757,N_20363,N_23945);
nor UO_1758 (O_1758,N_19394,N_23330);
or UO_1759 (O_1759,N_21024,N_22833);
or UO_1760 (O_1760,N_24780,N_19267);
xnor UO_1761 (O_1761,N_20028,N_19559);
xnor UO_1762 (O_1762,N_19396,N_24259);
xnor UO_1763 (O_1763,N_24323,N_19589);
nor UO_1764 (O_1764,N_21766,N_19976);
or UO_1765 (O_1765,N_22850,N_20201);
nand UO_1766 (O_1766,N_22933,N_23099);
nand UO_1767 (O_1767,N_24566,N_22070);
nand UO_1768 (O_1768,N_22378,N_21532);
xnor UO_1769 (O_1769,N_23385,N_22111);
nand UO_1770 (O_1770,N_22342,N_20936);
nor UO_1771 (O_1771,N_22088,N_21799);
and UO_1772 (O_1772,N_24285,N_18953);
nand UO_1773 (O_1773,N_24579,N_24436);
or UO_1774 (O_1774,N_19265,N_19340);
xnor UO_1775 (O_1775,N_18924,N_22505);
nand UO_1776 (O_1776,N_23455,N_24414);
and UO_1777 (O_1777,N_24496,N_24779);
or UO_1778 (O_1778,N_22170,N_19548);
xor UO_1779 (O_1779,N_22776,N_24295);
and UO_1780 (O_1780,N_19653,N_21736);
nand UO_1781 (O_1781,N_23981,N_20797);
nor UO_1782 (O_1782,N_22412,N_21509);
and UO_1783 (O_1783,N_22175,N_18890);
or UO_1784 (O_1784,N_24035,N_23025);
nand UO_1785 (O_1785,N_19036,N_20904);
xor UO_1786 (O_1786,N_20834,N_22684);
or UO_1787 (O_1787,N_20587,N_19181);
or UO_1788 (O_1788,N_21916,N_24125);
nor UO_1789 (O_1789,N_19622,N_23250);
nand UO_1790 (O_1790,N_21593,N_21358);
and UO_1791 (O_1791,N_22782,N_23094);
nand UO_1792 (O_1792,N_20617,N_21764);
and UO_1793 (O_1793,N_19748,N_24935);
or UO_1794 (O_1794,N_20647,N_21089);
nand UO_1795 (O_1795,N_18775,N_24164);
nor UO_1796 (O_1796,N_24574,N_23307);
nand UO_1797 (O_1797,N_22244,N_24368);
and UO_1798 (O_1798,N_19085,N_20174);
nand UO_1799 (O_1799,N_19919,N_21998);
nor UO_1800 (O_1800,N_21320,N_19807);
nand UO_1801 (O_1801,N_23107,N_20703);
xnor UO_1802 (O_1802,N_20570,N_20606);
nand UO_1803 (O_1803,N_21590,N_19429);
and UO_1804 (O_1804,N_20673,N_23430);
or UO_1805 (O_1805,N_24410,N_20750);
and UO_1806 (O_1806,N_23205,N_19388);
xnor UO_1807 (O_1807,N_24615,N_21946);
xor UO_1808 (O_1808,N_24674,N_23187);
xnor UO_1809 (O_1809,N_22355,N_21173);
xor UO_1810 (O_1810,N_24694,N_21104);
xor UO_1811 (O_1811,N_22341,N_19408);
nor UO_1812 (O_1812,N_21251,N_20027);
or UO_1813 (O_1813,N_22897,N_23446);
or UO_1814 (O_1814,N_24648,N_21143);
or UO_1815 (O_1815,N_23827,N_21906);
nor UO_1816 (O_1816,N_18948,N_23137);
nor UO_1817 (O_1817,N_24609,N_18827);
nor UO_1818 (O_1818,N_20611,N_19203);
nand UO_1819 (O_1819,N_22693,N_23333);
nor UO_1820 (O_1820,N_19756,N_20754);
xnor UO_1821 (O_1821,N_23659,N_23313);
nor UO_1822 (O_1822,N_20997,N_20479);
nor UO_1823 (O_1823,N_24523,N_22859);
and UO_1824 (O_1824,N_20110,N_19899);
and UO_1825 (O_1825,N_22805,N_19578);
and UO_1826 (O_1826,N_19957,N_19487);
or UO_1827 (O_1827,N_19514,N_23440);
xnor UO_1828 (O_1828,N_19045,N_20599);
nand UO_1829 (O_1829,N_23532,N_20421);
or UO_1830 (O_1830,N_24292,N_21203);
or UO_1831 (O_1831,N_20882,N_19216);
nor UO_1832 (O_1832,N_19285,N_21058);
and UO_1833 (O_1833,N_21160,N_20802);
and UO_1834 (O_1834,N_19206,N_23727);
nor UO_1835 (O_1835,N_24203,N_20865);
xor UO_1836 (O_1836,N_21010,N_21507);
nand UO_1837 (O_1837,N_19015,N_20986);
and UO_1838 (O_1838,N_20429,N_21526);
or UO_1839 (O_1839,N_20234,N_20737);
nand UO_1840 (O_1840,N_22766,N_21325);
xor UO_1841 (O_1841,N_24351,N_24578);
or UO_1842 (O_1842,N_24675,N_19606);
and UO_1843 (O_1843,N_21944,N_23935);
nand UO_1844 (O_1844,N_24007,N_23851);
or UO_1845 (O_1845,N_24692,N_23964);
and UO_1846 (O_1846,N_19128,N_23461);
nor UO_1847 (O_1847,N_19283,N_22915);
nand UO_1848 (O_1848,N_23773,N_24817);
xnor UO_1849 (O_1849,N_22221,N_24200);
and UO_1850 (O_1850,N_20979,N_19988);
nor UO_1851 (O_1851,N_19638,N_24701);
xnor UO_1852 (O_1852,N_24957,N_24620);
nor UO_1853 (O_1853,N_24187,N_24770);
or UO_1854 (O_1854,N_23991,N_20735);
nand UO_1855 (O_1855,N_19365,N_22291);
nand UO_1856 (O_1856,N_22547,N_22122);
and UO_1857 (O_1857,N_21825,N_19373);
or UO_1858 (O_1858,N_21355,N_21708);
or UO_1859 (O_1859,N_21430,N_21751);
or UO_1860 (O_1860,N_20368,N_23479);
nand UO_1861 (O_1861,N_21205,N_23608);
nand UO_1862 (O_1862,N_20448,N_23971);
nor UO_1863 (O_1863,N_18883,N_19550);
and UO_1864 (O_1864,N_24754,N_20493);
or UO_1865 (O_1865,N_22017,N_19121);
nand UO_1866 (O_1866,N_24992,N_21063);
and UO_1867 (O_1867,N_22719,N_22590);
nand UO_1868 (O_1868,N_22263,N_21340);
or UO_1869 (O_1869,N_22598,N_23070);
or UO_1870 (O_1870,N_23049,N_21268);
nand UO_1871 (O_1871,N_21658,N_22394);
or UO_1872 (O_1872,N_21744,N_23685);
nand UO_1873 (O_1873,N_19793,N_23790);
nor UO_1874 (O_1874,N_23593,N_21070);
nor UO_1875 (O_1875,N_21498,N_22940);
nor UO_1876 (O_1876,N_19399,N_20190);
nor UO_1877 (O_1877,N_23359,N_24527);
nor UO_1878 (O_1878,N_21114,N_21961);
or UO_1879 (O_1879,N_19472,N_23520);
nand UO_1880 (O_1880,N_21931,N_21704);
and UO_1881 (O_1881,N_19830,N_20290);
xor UO_1882 (O_1882,N_21441,N_24276);
nand UO_1883 (O_1883,N_24987,N_20202);
or UO_1884 (O_1884,N_24532,N_20811);
xor UO_1885 (O_1885,N_23707,N_20263);
or UO_1886 (O_1886,N_22760,N_22454);
nor UO_1887 (O_1887,N_19607,N_19995);
nor UO_1888 (O_1888,N_22779,N_20512);
nand UO_1889 (O_1889,N_22606,N_20353);
nand UO_1890 (O_1890,N_24718,N_20188);
nand UO_1891 (O_1891,N_24439,N_21130);
or UO_1892 (O_1892,N_22983,N_24884);
and UO_1893 (O_1893,N_19224,N_20191);
and UO_1894 (O_1894,N_24622,N_20103);
or UO_1895 (O_1895,N_22546,N_23600);
or UO_1896 (O_1896,N_18892,N_19243);
nor UO_1897 (O_1897,N_20007,N_18996);
nand UO_1898 (O_1898,N_22313,N_22067);
nand UO_1899 (O_1899,N_22622,N_23280);
nor UO_1900 (O_1900,N_19086,N_24190);
and UO_1901 (O_1901,N_19621,N_20115);
or UO_1902 (O_1902,N_20995,N_20613);
and UO_1903 (O_1903,N_22628,N_20338);
or UO_1904 (O_1904,N_24387,N_24991);
xnor UO_1905 (O_1905,N_23865,N_21169);
xnor UO_1906 (O_1906,N_22913,N_19020);
and UO_1907 (O_1907,N_19841,N_19989);
or UO_1908 (O_1908,N_20231,N_23780);
xnor UO_1909 (O_1909,N_22832,N_24593);
nor UO_1910 (O_1910,N_24122,N_21494);
xor UO_1911 (O_1911,N_22425,N_22916);
xnor UO_1912 (O_1912,N_22936,N_22196);
nor UO_1913 (O_1913,N_20982,N_22826);
nor UO_1914 (O_1914,N_23970,N_21543);
nor UO_1915 (O_1915,N_21339,N_24305);
xnor UO_1916 (O_1916,N_19161,N_22639);
or UO_1917 (O_1917,N_21117,N_20985);
xor UO_1918 (O_1918,N_23883,N_22182);
nor UO_1919 (O_1919,N_24160,N_22860);
nor UO_1920 (O_1920,N_22521,N_18934);
or UO_1921 (O_1921,N_22363,N_19909);
or UO_1922 (O_1922,N_24676,N_23155);
or UO_1923 (O_1923,N_20449,N_19193);
nand UO_1924 (O_1924,N_22353,N_19614);
and UO_1925 (O_1925,N_18974,N_19905);
nand UO_1926 (O_1926,N_19349,N_19494);
or UO_1927 (O_1927,N_20035,N_21154);
nor UO_1928 (O_1928,N_19811,N_20128);
xor UO_1929 (O_1929,N_21738,N_21652);
nor UO_1930 (O_1930,N_20484,N_21913);
xor UO_1931 (O_1931,N_23997,N_20319);
xnor UO_1932 (O_1932,N_22053,N_23701);
xnor UO_1933 (O_1933,N_19848,N_19440);
nor UO_1934 (O_1934,N_19525,N_22320);
or UO_1935 (O_1935,N_18832,N_20070);
nand UO_1936 (O_1936,N_19451,N_20883);
or UO_1937 (O_1937,N_20720,N_23358);
xor UO_1938 (O_1938,N_22183,N_22756);
nor UO_1939 (O_1939,N_24824,N_19701);
nor UO_1940 (O_1940,N_22203,N_21489);
and UO_1941 (O_1941,N_23083,N_20279);
nor UO_1942 (O_1942,N_20690,N_23627);
nand UO_1943 (O_1943,N_22895,N_22009);
xnor UO_1944 (O_1944,N_20494,N_22193);
and UO_1945 (O_1945,N_19752,N_22517);
or UO_1946 (O_1946,N_20114,N_21125);
and UO_1947 (O_1947,N_22457,N_21502);
xnor UO_1948 (O_1948,N_21782,N_18783);
nand UO_1949 (O_1949,N_22236,N_20566);
nor UO_1950 (O_1950,N_21568,N_22508);
and UO_1951 (O_1951,N_24982,N_24070);
xnor UO_1952 (O_1952,N_21829,N_22252);
nand UO_1953 (O_1953,N_22479,N_19428);
or UO_1954 (O_1954,N_24834,N_23661);
or UO_1955 (O_1955,N_23640,N_23830);
nor UO_1956 (O_1956,N_19563,N_18826);
nor UO_1957 (O_1957,N_21995,N_19470);
and UO_1958 (O_1958,N_19634,N_20386);
nand UO_1959 (O_1959,N_20136,N_23611);
and UO_1960 (O_1960,N_24511,N_20543);
nand UO_1961 (O_1961,N_20602,N_19112);
or UO_1962 (O_1962,N_19321,N_23711);
nand UO_1963 (O_1963,N_20121,N_20684);
and UO_1964 (O_1964,N_23998,N_22440);
xor UO_1965 (O_1965,N_19393,N_24282);
and UO_1966 (O_1966,N_23766,N_19954);
nor UO_1967 (O_1967,N_24726,N_19697);
and UO_1968 (O_1968,N_19806,N_23878);
or UO_1969 (O_1969,N_21280,N_21410);
and UO_1970 (O_1970,N_22737,N_22224);
nor UO_1971 (O_1971,N_24311,N_21327);
nand UO_1972 (O_1972,N_21259,N_24559);
nor UO_1973 (O_1973,N_21226,N_20552);
xor UO_1974 (O_1974,N_24130,N_20350);
nor UO_1975 (O_1975,N_21209,N_23764);
or UO_1976 (O_1976,N_21884,N_19355);
nand UO_1977 (O_1977,N_21603,N_22610);
or UO_1978 (O_1978,N_21500,N_19676);
or UO_1979 (O_1979,N_20171,N_22385);
and UO_1980 (O_1980,N_22407,N_21539);
or UO_1981 (O_1981,N_20515,N_23509);
nand UO_1982 (O_1982,N_22427,N_20749);
nor UO_1983 (O_1983,N_22266,N_23115);
or UO_1984 (O_1984,N_24705,N_21373);
nand UO_1985 (O_1985,N_23195,N_24242);
and UO_1986 (O_1986,N_21861,N_24890);
nand UO_1987 (O_1987,N_23328,N_22700);
nand UO_1988 (O_1988,N_22198,N_23120);
xnor UO_1989 (O_1989,N_21414,N_20854);
nand UO_1990 (O_1990,N_24076,N_20563);
and UO_1991 (O_1991,N_23625,N_19734);
or UO_1992 (O_1992,N_22139,N_23840);
nand UO_1993 (O_1993,N_24231,N_20560);
xnor UO_1994 (O_1994,N_24047,N_19447);
nand UO_1995 (O_1995,N_24746,N_21557);
xnor UO_1996 (O_1996,N_21578,N_23260);
and UO_1997 (O_1997,N_22559,N_24971);
nor UO_1998 (O_1998,N_20246,N_22357);
nand UO_1999 (O_1999,N_23061,N_19536);
xnor UO_2000 (O_2000,N_22420,N_22184);
and UO_2001 (O_2001,N_24133,N_22254);
and UO_2002 (O_2002,N_23158,N_22641);
nor UO_2003 (O_2003,N_19649,N_22935);
or UO_2004 (O_2004,N_22251,N_23036);
or UO_2005 (O_2005,N_20659,N_23409);
nand UO_2006 (O_2006,N_22788,N_20090);
or UO_2007 (O_2007,N_19592,N_23389);
nor UO_2008 (O_2008,N_24147,N_23386);
nor UO_2009 (O_2009,N_23924,N_23668);
and UO_2010 (O_2010,N_24502,N_23814);
nor UO_2011 (O_2011,N_23863,N_24315);
or UO_2012 (O_2012,N_21678,N_24526);
xnor UO_2013 (O_2013,N_20706,N_24143);
nand UO_2014 (O_2014,N_24134,N_24179);
and UO_2015 (O_2015,N_22421,N_23926);
or UO_2016 (O_2016,N_18991,N_20172);
and UO_2017 (O_2017,N_24411,N_19021);
or UO_2018 (O_2018,N_20607,N_21411);
xnor UO_2019 (O_2019,N_19810,N_24142);
xnor UO_2020 (O_2020,N_24962,N_21974);
nor UO_2021 (O_2021,N_24985,N_22838);
nor UO_2022 (O_2022,N_20918,N_19311);
xor UO_2023 (O_2023,N_23474,N_19509);
nor UO_2024 (O_2024,N_24026,N_19759);
and UO_2025 (O_2025,N_24556,N_20757);
and UO_2026 (O_2026,N_23988,N_20569);
nand UO_2027 (O_2027,N_24114,N_24994);
and UO_2028 (O_2028,N_20295,N_22982);
and UO_2029 (O_2029,N_23437,N_21356);
nand UO_2030 (O_2030,N_22689,N_19222);
nor UO_2031 (O_2031,N_23431,N_23329);
or UO_2032 (O_2032,N_21141,N_23526);
and UO_2033 (O_2033,N_24588,N_18805);
nand UO_2034 (O_2034,N_19141,N_22380);
or UO_2035 (O_2035,N_23717,N_24883);
xor UO_2036 (O_2036,N_19891,N_20375);
nor UO_2037 (O_2037,N_23059,N_19668);
or UO_2038 (O_2038,N_24688,N_21687);
nand UO_2039 (O_2039,N_22281,N_23658);
xnor UO_2040 (O_2040,N_20836,N_22306);
or UO_2041 (O_2041,N_19198,N_22653);
xor UO_2042 (O_2042,N_24900,N_19363);
or UO_2043 (O_2043,N_23670,N_24201);
nand UO_2044 (O_2044,N_23705,N_20179);
or UO_2045 (O_2045,N_24806,N_21549);
nand UO_2046 (O_2046,N_20101,N_19792);
nor UO_2047 (O_2047,N_22463,N_21803);
nor UO_2048 (O_2048,N_19642,N_20815);
nand UO_2049 (O_2049,N_21712,N_21567);
or UO_2050 (O_2050,N_19515,N_24640);
xnor UO_2051 (O_2051,N_19726,N_23397);
and UO_2052 (O_2052,N_20595,N_23634);
nand UO_2053 (O_2053,N_22185,N_24038);
nand UO_2054 (O_2054,N_23564,N_19802);
and UO_2055 (O_2055,N_24319,N_20022);
xor UO_2056 (O_2056,N_19529,N_24686);
nor UO_2057 (O_2057,N_20681,N_24554);
and UO_2058 (O_2058,N_22651,N_22455);
nor UO_2059 (O_2059,N_22692,N_19705);
nand UO_2060 (O_2060,N_24889,N_21147);
and UO_2061 (O_2061,N_21418,N_20971);
nor UO_2062 (O_2062,N_20886,N_24423);
and UO_2063 (O_2063,N_18903,N_21510);
or UO_2064 (O_2064,N_19537,N_21508);
or UO_2065 (O_2065,N_22582,N_21611);
and UO_2066 (O_2066,N_19060,N_21890);
nor UO_2067 (O_2067,N_22095,N_21462);
nand UO_2068 (O_2068,N_19965,N_21699);
nand UO_2069 (O_2069,N_24077,N_24326);
and UO_2070 (O_2070,N_24378,N_24654);
nor UO_2071 (O_2071,N_20545,N_20535);
nand UO_2072 (O_2072,N_23335,N_20004);
nand UO_2073 (O_2073,N_19057,N_22948);
nor UO_2074 (O_2074,N_22150,N_19551);
nor UO_2075 (O_2075,N_24724,N_19616);
xnor UO_2076 (O_2076,N_23894,N_20383);
xnor UO_2077 (O_2077,N_24741,N_19046);
nand UO_2078 (O_2078,N_19316,N_24100);
xnor UO_2079 (O_2079,N_21957,N_23093);
nor UO_2080 (O_2080,N_20018,N_22570);
nand UO_2081 (O_2081,N_19522,N_23344);
nor UO_2082 (O_2082,N_23517,N_23786);
xor UO_2083 (O_2083,N_22771,N_20396);
nor UO_2084 (O_2084,N_19053,N_22488);
xnor UO_2085 (O_2085,N_24165,N_20214);
or UO_2086 (O_2086,N_22973,N_23433);
nand UO_2087 (O_2087,N_22137,N_20816);
nor UO_2088 (O_2088,N_19050,N_19320);
nand UO_2089 (O_2089,N_21628,N_21660);
nand UO_2090 (O_2090,N_22097,N_22443);
nor UO_2091 (O_2091,N_19323,N_22820);
and UO_2092 (O_2092,N_22227,N_22276);
xor UO_2093 (O_2093,N_20525,N_19347);
xor UO_2094 (O_2094,N_19687,N_23800);
xnor UO_2095 (O_2095,N_22442,N_23770);
and UO_2096 (O_2096,N_24080,N_21565);
or UO_2097 (O_2097,N_22785,N_19497);
nor UO_2098 (O_2098,N_20481,N_23868);
or UO_2099 (O_2099,N_22808,N_20151);
and UO_2100 (O_2100,N_23587,N_21752);
nor UO_2101 (O_2101,N_21465,N_19952);
nor UO_2102 (O_2102,N_22720,N_19221);
and UO_2103 (O_2103,N_18812,N_20457);
xnor UO_2104 (O_2104,N_23803,N_22657);
and UO_2105 (O_2105,N_22047,N_18778);
and UO_2106 (O_2106,N_21591,N_20794);
nor UO_2107 (O_2107,N_22856,N_24507);
nor UO_2108 (O_2108,N_22459,N_19091);
xnor UO_2109 (O_2109,N_21748,N_20916);
nor UO_2110 (O_2110,N_19219,N_20392);
nor UO_2111 (O_2111,N_20055,N_18799);
or UO_2112 (O_2112,N_18887,N_23881);
and UO_2113 (O_2113,N_19156,N_21302);
or UO_2114 (O_2114,N_19435,N_20937);
and UO_2115 (O_2115,N_23220,N_24820);
xnor UO_2116 (O_2116,N_24415,N_21107);
nor UO_2117 (O_2117,N_21637,N_23708);
or UO_2118 (O_2118,N_23363,N_19913);
xnor UO_2119 (O_2119,N_21666,N_20711);
or UO_2120 (O_2120,N_22683,N_21486);
nand UO_2121 (O_2121,N_22059,N_24469);
nand UO_2122 (O_2122,N_22485,N_19467);
nor UO_2123 (O_2123,N_18894,N_23797);
nor UO_2124 (O_2124,N_23544,N_20140);
nand UO_2125 (O_2125,N_22456,N_24341);
or UO_2126 (O_2126,N_21745,N_21577);
nor UO_2127 (O_2127,N_20379,N_20106);
xnor UO_2128 (O_2128,N_20951,N_19544);
nor UO_2129 (O_2129,N_20988,N_24486);
and UO_2130 (O_2130,N_24065,N_23045);
nor UO_2131 (O_2131,N_23756,N_22382);
and UO_2132 (O_2132,N_24372,N_21072);
or UO_2133 (O_2133,N_23374,N_22862);
xor UO_2134 (O_2134,N_24465,N_23112);
nor UO_2135 (O_2135,N_19901,N_22075);
nor UO_2136 (O_2136,N_24324,N_20874);
nand UO_2137 (O_2137,N_22742,N_20922);
nor UO_2138 (O_2138,N_19679,N_22142);
xnor UO_2139 (O_2139,N_20405,N_21198);
nand UO_2140 (O_2140,N_21116,N_21722);
nor UO_2141 (O_2141,N_22619,N_21029);
nand UO_2142 (O_2142,N_24280,N_19397);
xnor UO_2143 (O_2143,N_21201,N_21978);
or UO_2144 (O_2144,N_19955,N_24852);
xor UO_2145 (O_2145,N_24498,N_20715);
and UO_2146 (O_2146,N_19588,N_20423);
nor UO_2147 (O_2147,N_22340,N_18908);
nand UO_2148 (O_2148,N_18824,N_20974);
and UO_2149 (O_2149,N_22710,N_23266);
nand UO_2150 (O_2150,N_22083,N_19378);
and UO_2151 (O_2151,N_21214,N_21458);
and UO_2152 (O_2152,N_22128,N_23257);
or UO_2153 (O_2153,N_19145,N_21634);
xor UO_2154 (O_2154,N_19938,N_23784);
or UO_2155 (O_2155,N_20372,N_23553);
nand UO_2156 (O_2156,N_21318,N_24989);
and UO_2157 (O_2157,N_24988,N_20194);
nor UO_2158 (O_2158,N_20894,N_23017);
or UO_2159 (O_2159,N_24995,N_22515);
or UO_2160 (O_2160,N_22253,N_22806);
nand UO_2161 (O_2161,N_22642,N_20111);
or UO_2162 (O_2162,N_23233,N_22247);
nand UO_2163 (O_2163,N_23859,N_21527);
nand UO_2164 (O_2164,N_23966,N_21734);
nand UO_2165 (O_2165,N_21456,N_21375);
nand UO_2166 (O_2166,N_22975,N_22910);
nand UO_2167 (O_2167,N_22609,N_21689);
or UO_2168 (O_2168,N_18833,N_21747);
xnor UO_2169 (O_2169,N_19258,N_20252);
or UO_2170 (O_2170,N_21705,N_21263);
xnor UO_2171 (O_2171,N_22398,N_23514);
nor UO_2172 (O_2172,N_21720,N_19434);
and UO_2173 (O_2173,N_22536,N_22513);
or UO_2174 (O_2174,N_23415,N_24595);
and UO_2175 (O_2175,N_24458,N_19761);
xnor UO_2176 (O_2176,N_22676,N_21417);
xnor UO_2177 (O_2177,N_22284,N_20229);
or UO_2178 (O_2178,N_21412,N_20966);
nor UO_2179 (O_2179,N_21860,N_24865);
nor UO_2180 (O_2180,N_22881,N_24521);
or UO_2181 (O_2181,N_19657,N_23732);
xnor UO_2182 (O_2182,N_23754,N_21042);
or UO_2183 (O_2183,N_22954,N_20474);
and UO_2184 (O_2184,N_21669,N_21671);
nand UO_2185 (O_2185,N_21434,N_22950);
nor UO_2186 (O_2186,N_19713,N_21586);
and UO_2187 (O_2187,N_20553,N_19102);
nand UO_2188 (O_2188,N_24917,N_23408);
xnor UO_2189 (O_2189,N_22369,N_23400);
xnor UO_2190 (O_2190,N_18785,N_19686);
or UO_2191 (O_2191,N_19061,N_21954);
nand UO_2192 (O_2192,N_23596,N_20812);
xor UO_2193 (O_2193,N_21194,N_23826);
nand UO_2194 (O_2194,N_19163,N_24543);
nand UO_2195 (O_2195,N_22384,N_23724);
nor UO_2196 (O_2196,N_19915,N_20597);
and UO_2197 (O_2197,N_20630,N_24515);
nand UO_2198 (O_2198,N_20964,N_23561);
nor UO_2199 (O_2199,N_19382,N_24783);
or UO_2200 (O_2200,N_20724,N_23494);
xor UO_2201 (O_2201,N_19261,N_22014);
or UO_2202 (O_2202,N_23657,N_23232);
xor UO_2203 (O_2203,N_24657,N_21670);
or UO_2204 (O_2204,N_22891,N_24711);
nand UO_2205 (O_2205,N_22522,N_21389);
nand UO_2206 (O_2206,N_19576,N_24822);
and UO_2207 (O_2207,N_19962,N_22896);
nand UO_2208 (O_2208,N_23794,N_18869);
nor UO_2209 (O_2209,N_21254,N_23040);
and UO_2210 (O_2210,N_23073,N_19754);
xor UO_2211 (O_2211,N_23268,N_23703);
nor UO_2212 (O_2212,N_20760,N_23603);
or UO_2213 (O_2213,N_19344,N_21255);
nand UO_2214 (O_2214,N_23789,N_23425);
and UO_2215 (O_2215,N_21138,N_23693);
nand UO_2216 (O_2216,N_20426,N_19040);
and UO_2217 (O_2217,N_22945,N_21876);
and UO_2218 (O_2218,N_19766,N_22889);
or UO_2219 (O_2219,N_24976,N_22944);
or UO_2220 (O_2220,N_24491,N_22662);
xor UO_2221 (O_2221,N_20786,N_21334);
xnor UO_2222 (O_2222,N_22995,N_18896);
nor UO_2223 (O_2223,N_19982,N_19119);
xor UO_2224 (O_2224,N_22665,N_22770);
nor UO_2225 (O_2225,N_20708,N_22731);
xnor UO_2226 (O_2226,N_23191,N_18927);
nor UO_2227 (O_2227,N_22825,N_23726);
or UO_2228 (O_2228,N_24389,N_19346);
or UO_2229 (O_2229,N_19391,N_19921);
or UO_2230 (O_2230,N_20005,N_19875);
xnor UO_2231 (O_2231,N_21898,N_24247);
or UO_2232 (O_2232,N_20643,N_20746);
nand UO_2233 (O_2233,N_20870,N_19842);
nor UO_2234 (O_2234,N_21156,N_22293);
xor UO_2235 (O_2235,N_21127,N_20767);
and UO_2236 (O_2236,N_18818,N_22601);
nand UO_2237 (O_2237,N_20296,N_20732);
and UO_2238 (O_2238,N_23793,N_24289);
nand UO_2239 (O_2239,N_21231,N_19645);
nor UO_2240 (O_2240,N_21583,N_18758);
or UO_2241 (O_2241,N_24893,N_24223);
and UO_2242 (O_2242,N_21057,N_22118);
xnor UO_2243 (O_2243,N_23628,N_21330);
xnor UO_2244 (O_2244,N_18971,N_20852);
or UO_2245 (O_2245,N_24232,N_23327);
and UO_2246 (O_2246,N_23716,N_24717);
xnor UO_2247 (O_2247,N_20251,N_22739);
and UO_2248 (O_2248,N_21016,N_20307);
nand UO_2249 (O_2249,N_24781,N_21602);
xor UO_2250 (O_2250,N_19836,N_20530);
nand UO_2251 (O_2251,N_19280,N_20536);
nor UO_2252 (O_2252,N_23919,N_24005);
xor UO_2253 (O_2253,N_24256,N_20040);
nor UO_2254 (O_2254,N_23720,N_19727);
and UO_2255 (O_2255,N_20469,N_23338);
xnor UO_2256 (O_2256,N_22980,N_24826);
xor UO_2257 (O_2257,N_20674,N_22675);
nand UO_2258 (O_2258,N_21992,N_23844);
nand UO_2259 (O_2259,N_23609,N_20686);
nor UO_2260 (O_2260,N_20393,N_22078);
and UO_2261 (O_2261,N_24944,N_19583);
nor UO_2262 (O_2262,N_20589,N_19664);
nor UO_2263 (O_2263,N_20956,N_21985);
xnor UO_2264 (O_2264,N_24338,N_22792);
or UO_2265 (O_2265,N_23562,N_21948);
nor UO_2266 (O_2266,N_21088,N_24093);
and UO_2267 (O_2267,N_19968,N_21775);
or UO_2268 (O_2268,N_23721,N_24829);
or UO_2269 (O_2269,N_23192,N_21427);
nor UO_2270 (O_2270,N_23247,N_23482);
nand UO_2271 (O_2271,N_19354,N_24827);
nand UO_2272 (O_2272,N_22783,N_20685);
nor UO_2273 (O_2273,N_22549,N_20862);
nand UO_2274 (O_2274,N_24612,N_19274);
or UO_2275 (O_2275,N_19445,N_22865);
nor UO_2276 (O_2276,N_19123,N_21987);
or UO_2277 (O_2277,N_19278,N_21413);
and UO_2278 (O_2278,N_20654,N_21047);
or UO_2279 (O_2279,N_23149,N_21272);
nor UO_2280 (O_2280,N_23156,N_18760);
or UO_2281 (O_2281,N_22572,N_18906);
and UO_2282 (O_2282,N_21544,N_21453);
nand UO_2283 (O_2283,N_19596,N_19930);
or UO_2284 (O_2284,N_19370,N_23264);
xor UO_2285 (O_2285,N_21463,N_19704);
and UO_2286 (O_2286,N_24902,N_22733);
nor UO_2287 (O_2287,N_23929,N_24956);
or UO_2288 (O_2288,N_22446,N_19975);
xor UO_2289 (O_2289,N_22119,N_21936);
nand UO_2290 (O_2290,N_21490,N_20387);
or UO_2291 (O_2291,N_24730,N_21131);
or UO_2292 (O_2292,N_18773,N_23550);
and UO_2293 (O_2293,N_19187,N_19717);
and UO_2294 (O_2294,N_19987,N_18792);
xor UO_2295 (O_2295,N_19740,N_21594);
or UO_2296 (O_2296,N_20631,N_24755);
nand UO_2297 (O_2297,N_24557,N_20879);
xor UO_2298 (O_2298,N_22970,N_22520);
or UO_2299 (O_2299,N_22909,N_24329);
xor UO_2300 (O_2300,N_20086,N_24407);
xnor UO_2301 (O_2301,N_20158,N_23212);
nor UO_2302 (O_2302,N_22152,N_23450);
xor UO_2303 (O_2303,N_24384,N_22875);
or UO_2304 (O_2304,N_21757,N_20949);
or UO_2305 (O_2305,N_24482,N_23225);
or UO_2306 (O_2306,N_19042,N_19247);
and UO_2307 (O_2307,N_22117,N_22448);
or UO_2308 (O_2308,N_19556,N_23202);
or UO_2309 (O_2309,N_20051,N_20381);
nand UO_2310 (O_2310,N_20374,N_18808);
xnor UO_2311 (O_2311,N_21403,N_23090);
or UO_2312 (O_2312,N_19212,N_23534);
and UO_2313 (O_2313,N_21609,N_23604);
and UO_2314 (O_2314,N_22233,N_24103);
nor UO_2315 (O_2315,N_23028,N_19075);
nor UO_2316 (O_2316,N_20594,N_20077);
nand UO_2317 (O_2317,N_20506,N_22197);
nor UO_2318 (O_2318,N_24833,N_22991);
xnor UO_2319 (O_2319,N_18840,N_24774);
xor UO_2320 (O_2320,N_21176,N_19760);
nand UO_2321 (O_2321,N_20683,N_20113);
or UO_2322 (O_2322,N_23201,N_19379);
and UO_2323 (O_2323,N_21746,N_24951);
and UO_2324 (O_2324,N_20177,N_19893);
or UO_2325 (O_2325,N_23089,N_21344);
nor UO_2326 (O_2326,N_24945,N_19097);
and UO_2327 (O_2327,N_21365,N_19252);
xnor UO_2328 (O_2328,N_22449,N_23117);
nand UO_2329 (O_2329,N_23246,N_24630);
nand UO_2330 (O_2330,N_21152,N_19263);
nand UO_2331 (O_2331,N_23607,N_22173);
nand UO_2332 (O_2332,N_20107,N_20710);
nand UO_2333 (O_2333,N_22643,N_24909);
nand UO_2334 (O_2334,N_18884,N_21374);
and UO_2335 (O_2335,N_20364,N_22712);
and UO_2336 (O_2336,N_22334,N_20795);
or UO_2337 (O_2337,N_20532,N_21495);
nor UO_2338 (O_2338,N_23370,N_18816);
nor UO_2339 (O_2339,N_19593,N_22530);
or UO_2340 (O_2340,N_24784,N_20909);
nor UO_2341 (O_2341,N_19148,N_21657);
xor UO_2342 (O_2342,N_23023,N_22477);
and UO_2343 (O_2343,N_23032,N_19268);
nand UO_2344 (O_2344,N_18970,N_23095);
or UO_2345 (O_2345,N_22943,N_23558);
and UO_2346 (O_2346,N_24493,N_23179);
xnor UO_2347 (O_2347,N_19113,N_24435);
or UO_2348 (O_2348,N_21492,N_24406);
and UO_2349 (O_2349,N_21229,N_23035);
and UO_2350 (O_2350,N_21477,N_19106);
nor UO_2351 (O_2351,N_21182,N_19081);
nand UO_2352 (O_2352,N_21668,N_19725);
xor UO_2353 (O_2353,N_19673,N_24192);
and UO_2354 (O_2354,N_20445,N_19643);
nor UO_2355 (O_2355,N_20810,N_24668);
xnor UO_2356 (O_2356,N_23055,N_22997);
nor UO_2357 (O_2357,N_21467,N_24769);
and UO_2358 (O_2358,N_20411,N_18982);
and UO_2359 (O_2359,N_24478,N_21112);
xnor UO_2360 (O_2360,N_22866,N_22535);
and UO_2361 (O_2361,N_22338,N_20483);
or UO_2362 (O_2362,N_24075,N_21096);
and UO_2363 (O_2363,N_18918,N_21521);
nor UO_2364 (O_2364,N_22151,N_22373);
nor UO_2365 (O_2365,N_23317,N_23428);
and UO_2366 (O_2366,N_21739,N_19150);
and UO_2367 (O_2367,N_19270,N_23139);
nand UO_2368 (O_2368,N_21485,N_19738);
and UO_2369 (O_2369,N_21439,N_21795);
xor UO_2370 (O_2370,N_20652,N_19188);
nor UO_2371 (O_2371,N_23704,N_22043);
or UO_2372 (O_2372,N_23194,N_19105);
nor UO_2373 (O_2373,N_21036,N_21646);
and UO_2374 (O_2374,N_19465,N_24350);
nor UO_2375 (O_2375,N_22872,N_20285);
nand UO_2376 (O_2376,N_18759,N_19720);
nand UO_2377 (O_2377,N_19452,N_23804);
nand UO_2378 (O_2378,N_20056,N_20790);
nor UO_2379 (O_2379,N_21360,N_21945);
or UO_2380 (O_2380,N_20210,N_24331);
nor UO_2381 (O_2381,N_20853,N_20572);
and UO_2382 (O_2382,N_21177,N_20144);
nand UO_2383 (O_2383,N_21199,N_21807);
nor UO_2384 (O_2384,N_20738,N_21920);
nor UO_2385 (O_2385,N_22205,N_21273);
and UO_2386 (O_2386,N_24564,N_22695);
xor UO_2387 (O_2387,N_19786,N_20068);
nand UO_2388 (O_2388,N_21610,N_21346);
xnor UO_2389 (O_2389,N_21877,N_19235);
or UO_2390 (O_2390,N_21123,N_23245);
xor UO_2391 (O_2391,N_21505,N_23109);
nand UO_2392 (O_2392,N_20727,N_21819);
nand UO_2393 (O_2393,N_20373,N_21223);
and UO_2394 (O_2394,N_22750,N_24514);
xnor UO_2395 (O_2395,N_19874,N_20166);
xor UO_2396 (O_2396,N_20313,N_20402);
xnor UO_2397 (O_2397,N_23530,N_19707);
and UO_2398 (O_2398,N_23920,N_21466);
nor UO_2399 (O_2399,N_21021,N_24239);
xnor UO_2400 (O_2400,N_22041,N_19543);
or UO_2401 (O_2401,N_20528,N_23362);
nor UO_2402 (O_2402,N_19426,N_19684);
and UO_2403 (O_2403,N_23946,N_24601);
xor UO_2404 (O_2404,N_24455,N_22158);
and UO_2405 (O_2405,N_23671,N_21547);
xnor UO_2406 (O_2406,N_20947,N_20477);
or UO_2407 (O_2407,N_20260,N_23547);
xor UO_2408 (O_2408,N_19907,N_19540);
xor UO_2409 (O_2409,N_20173,N_19967);
or UO_2410 (O_2410,N_24735,N_21851);
nor UO_2411 (O_2411,N_20888,N_24703);
and UO_2412 (O_2412,N_18754,N_20924);
and UO_2413 (O_2413,N_23336,N_23320);
nand UO_2414 (O_2414,N_24227,N_21548);
and UO_2415 (O_2415,N_21014,N_21733);
xor UO_2416 (O_2416,N_21904,N_21432);
or UO_2417 (O_2417,N_21121,N_19922);
xor UO_2418 (O_2418,N_20442,N_19817);
and UO_2419 (O_2419,N_21298,N_19194);
or UO_2420 (O_2420,N_20503,N_20502);
or UO_2421 (O_2421,N_21336,N_19230);
xor UO_2422 (O_2422,N_23569,N_23442);
nand UO_2423 (O_2423,N_24481,N_20887);
nand UO_2424 (O_2424,N_20286,N_18994);
xor UO_2425 (O_2425,N_23334,N_22413);
xnor UO_2426 (O_2426,N_24765,N_20896);
nor UO_2427 (O_2427,N_23126,N_23907);
or UO_2428 (O_2428,N_22491,N_22143);
nor UO_2429 (O_2429,N_23324,N_20218);
nor UO_2430 (O_2430,N_23002,N_23504);
nand UO_2431 (O_2431,N_19372,N_24847);
nor UO_2432 (O_2432,N_19869,N_20798);
xnor UO_2433 (O_2433,N_21015,N_24509);
xnor UO_2434 (O_2434,N_20354,N_23895);
and UO_2435 (O_2435,N_20297,N_24024);
and UO_2436 (O_2436,N_19658,N_22728);
nor UO_2437 (O_2437,N_22921,N_24025);
or UO_2438 (O_2438,N_24298,N_20235);
xnor UO_2439 (O_2439,N_24128,N_23435);
or UO_2440 (O_2440,N_18972,N_19667);
or UO_2441 (O_2441,N_22409,N_19404);
nand UO_2442 (O_2442,N_19744,N_20346);
or UO_2443 (O_2443,N_19700,N_24213);
nand UO_2444 (O_2444,N_19374,N_20222);
and UO_2445 (O_2445,N_24872,N_23419);
nand UO_2446 (O_2446,N_23454,N_21631);
and UO_2447 (O_2447,N_19254,N_20306);
nor UO_2448 (O_2448,N_19456,N_20803);
or UO_2449 (O_2449,N_22052,N_23418);
or UO_2450 (O_2450,N_23644,N_19101);
nor UO_2451 (O_2451,N_19231,N_22424);
nand UO_2452 (O_2452,N_22544,N_21659);
nor UO_2453 (O_2453,N_22445,N_24837);
or UO_2454 (O_2454,N_22919,N_21516);
nor UO_2455 (O_2455,N_24821,N_24861);
nor UO_2456 (O_2456,N_23879,N_24010);
xor UO_2457 (O_2457,N_20520,N_22772);
nor UO_2458 (O_2458,N_19896,N_20384);
or UO_2459 (O_2459,N_20069,N_24650);
and UO_2460 (O_2460,N_23696,N_23958);
and UO_2461 (O_2461,N_22336,N_24751);
nor UO_2462 (O_2462,N_18931,N_19857);
or UO_2463 (O_2463,N_23555,N_21020);
or UO_2464 (O_2464,N_21232,N_21133);
and UO_2465 (O_2465,N_21283,N_23402);
nand UO_2466 (O_2466,N_21299,N_20635);
and UO_2467 (O_2467,N_19528,N_21290);
nand UO_2468 (O_2468,N_21124,N_20554);
or UO_2469 (O_2469,N_23918,N_19084);
and UO_2470 (O_2470,N_22849,N_19214);
or UO_2471 (O_2471,N_24857,N_22145);
xor UO_2472 (O_2472,N_18789,N_22514);
xnor UO_2473 (O_2473,N_22020,N_19282);
and UO_2474 (O_2474,N_24926,N_20549);
and UO_2475 (O_2475,N_20609,N_21188);
or UO_2476 (O_2476,N_20394,N_24422);
nand UO_2477 (O_2477,N_22018,N_19946);
or UO_2478 (O_2478,N_23417,N_24346);
xnor UO_2479 (O_2479,N_23321,N_24608);
and UO_2480 (O_2480,N_20664,N_24699);
and UO_2481 (O_2481,N_23570,N_19631);
or UO_2482 (O_2482,N_20747,N_23516);
nor UO_2483 (O_2483,N_21718,N_20893);
nand UO_2484 (O_2484,N_18839,N_19787);
xor UO_2485 (O_2485,N_18955,N_19703);
and UO_2486 (O_2486,N_23100,N_20998);
xnor UO_2487 (O_2487,N_20948,N_20808);
or UO_2488 (O_2488,N_22493,N_19850);
or UO_2489 (O_2489,N_24693,N_23493);
nor UO_2490 (O_2490,N_22081,N_24807);
nand UO_2491 (O_2491,N_24151,N_22839);
or UO_2492 (O_2492,N_20029,N_24918);
or UO_2493 (O_2493,N_22949,N_22101);
nand UO_2494 (O_2494,N_24758,N_23862);
nor UO_2495 (O_2495,N_20329,N_20461);
and UO_2496 (O_2496,N_23038,N_22814);
nor UO_2497 (O_2497,N_19386,N_23274);
and UO_2498 (O_2498,N_20159,N_20161);
nand UO_2499 (O_2499,N_24215,N_24689);
and UO_2500 (O_2500,N_22006,N_22375);
or UO_2501 (O_2501,N_24091,N_23578);
and UO_2502 (O_2502,N_24359,N_19737);
xor UO_2503 (O_2503,N_24261,N_19632);
and UO_2504 (O_2504,N_24919,N_24480);
or UO_2505 (O_2505,N_22057,N_20967);
and UO_2506 (O_2506,N_22800,N_19478);
or UO_2507 (O_2507,N_24460,N_18943);
nand UO_2508 (O_2508,N_24120,N_23069);
xnor UO_2509 (O_2509,N_22703,N_23373);
and UO_2510 (O_2510,N_23642,N_18957);
nor UO_2511 (O_2511,N_23042,N_21837);
or UO_2512 (O_2512,N_22761,N_24792);
nor UO_2513 (O_2513,N_20127,N_22652);
and UO_2514 (O_2514,N_18984,N_23480);
nor UO_2515 (O_2515,N_22160,N_19253);
nor UO_2516 (O_2516,N_24078,N_19392);
xor UO_2517 (O_2517,N_20627,N_21690);
and UO_2518 (O_2518,N_21451,N_19387);
and UO_2519 (O_2519,N_22153,N_24656);
or UO_2520 (O_2520,N_23133,N_23393);
and UO_2521 (O_2521,N_22809,N_21195);
xor UO_2522 (O_2522,N_21518,N_22447);
and UO_2523 (O_2523,N_24937,N_24347);
nand UO_2524 (O_2524,N_20621,N_19827);
xnor UO_2525 (O_2525,N_19303,N_23586);
and UO_2526 (O_2526,N_19591,N_23936);
xor UO_2527 (O_2527,N_23765,N_23546);
nor UO_2528 (O_2528,N_21048,N_24592);
nor UO_2529 (O_2529,N_20446,N_19142);
xnor UO_2530 (O_2530,N_19876,N_21235);
xnor UO_2531 (O_2531,N_20981,N_19597);
or UO_2532 (O_2532,N_20629,N_21284);
nor UO_2533 (O_2533,N_21759,N_22589);
and UO_2534 (O_2534,N_22965,N_19610);
nand UO_2535 (O_2535,N_24036,N_21959);
nand UO_2536 (O_2536,N_19564,N_19886);
nor UO_2537 (O_2537,N_24413,N_23063);
and UO_2538 (O_2538,N_23491,N_21856);
xor UO_2539 (O_2539,N_18875,N_23502);
and UO_2540 (O_2540,N_24495,N_23451);
or UO_2541 (O_2541,N_21004,N_21808);
nand UO_2542 (O_2542,N_21240,N_24083);
or UO_2543 (O_2543,N_21080,N_21100);
nor UO_2544 (O_2544,N_20367,N_21217);
and UO_2545 (O_2545,N_18932,N_19661);
and UO_2546 (O_2546,N_19179,N_20024);
xor UO_2547 (O_2547,N_23410,N_21813);
and UO_2548 (O_2548,N_20833,N_22555);
or UO_2549 (O_2549,N_19966,N_22576);
and UO_2550 (O_2550,N_21960,N_21504);
xor UO_2551 (O_2551,N_24064,N_19660);
or UO_2552 (O_2552,N_21833,N_22906);
nor UO_2553 (O_2553,N_21241,N_22946);
or UO_2554 (O_2554,N_21654,N_18796);
or UO_2555 (O_2555,N_18837,N_20419);
nor UO_2556 (O_2556,N_20314,N_22033);
nand UO_2557 (O_2557,N_22393,N_21656);
xnor UO_2558 (O_2558,N_24576,N_23213);
xor UO_2559 (O_2559,N_18926,N_23680);
and UO_2560 (O_2560,N_20533,N_19407);
or UO_2561 (O_2561,N_21600,N_18815);
xor UO_2562 (O_2562,N_21926,N_19916);
nor UO_2563 (O_2563,N_21472,N_20934);
and UO_2564 (O_2564,N_19132,N_19879);
nor UO_2565 (O_2565,N_21250,N_24567);
nor UO_2566 (O_2566,N_19079,N_19821);
or UO_2567 (O_2567,N_20531,N_22192);
or UO_2568 (O_2568,N_21845,N_22155);
xnor UO_2569 (O_2569,N_22640,N_21099);
xor UO_2570 (O_2570,N_24835,N_24525);
xnor UO_2571 (O_2571,N_19770,N_23010);
and UO_2572 (O_2572,N_24257,N_24531);
xnor UO_2573 (O_2573,N_23164,N_19062);
nand UO_2574 (O_2574,N_21555,N_18856);
or UO_2575 (O_2575,N_21514,N_24137);
or UO_2576 (O_2576,N_18888,N_24728);
nor UO_2577 (O_2577,N_21017,N_19711);
xor UO_2578 (O_2578,N_23690,N_21471);
nand UO_2579 (O_2579,N_21921,N_24536);
or UO_2580 (O_2580,N_20612,N_23471);
nand UO_2581 (O_2581,N_23768,N_19880);
nand UO_2582 (O_2582,N_20968,N_20590);
nand UO_2583 (O_2583,N_21384,N_23922);
xnor UO_2584 (O_2584,N_23548,N_24986);
xor UO_2585 (O_2585,N_22958,N_20268);
and UO_2586 (O_2586,N_22722,N_20376);
xor UO_2587 (O_2587,N_21997,N_21216);
xnor UO_2588 (O_2588,N_23022,N_21279);
nand UO_2589 (O_2589,N_22126,N_21684);
nor UO_2590 (O_2590,N_22730,N_22588);
or UO_2591 (O_2591,N_19479,N_24449);
xnor UO_2592 (O_2592,N_19009,N_21445);
nand UO_2593 (O_2593,N_22831,N_19000);
nor UO_2594 (O_2594,N_20455,N_19089);
nand UO_2595 (O_2595,N_24174,N_24868);
and UO_2596 (O_2596,N_23836,N_18910);
nand UO_2597 (O_2597,N_18902,N_23105);
or UO_2598 (O_2598,N_21524,N_22974);
xnor UO_2599 (O_2599,N_22092,N_21727);
and UO_2600 (O_2600,N_19457,N_21675);
and UO_2601 (O_2601,N_20219,N_22671);
nor UO_2602 (O_2602,N_23180,N_23486);
nor UO_2603 (O_2603,N_24166,N_24843);
or UO_2604 (O_2604,N_23345,N_19871);
nor UO_2605 (O_2605,N_22670,N_21847);
nor UO_2606 (O_2606,N_20639,N_20038);
nor UO_2607 (O_2607,N_21550,N_20443);
nand UO_2608 (O_2608,N_24441,N_19225);
xor UO_2609 (O_2609,N_23066,N_20855);
nand UO_2610 (O_2610,N_20463,N_20186);
and UO_2611 (O_2611,N_19910,N_22026);
and UO_2612 (O_2612,N_23277,N_20133);
nor UO_2613 (O_2613,N_22475,N_21059);
and UO_2614 (O_2614,N_24050,N_20913);
or UO_2615 (O_2615,N_19402,N_22486);
or UO_2616 (O_2616,N_20640,N_19409);
and UO_2617 (O_2617,N_22562,N_19797);
xnor UO_2618 (O_2618,N_20598,N_23084);
nand UO_2619 (O_2619,N_23616,N_24416);
nand UO_2620 (O_2620,N_24268,N_19092);
or UO_2621 (O_2621,N_21842,N_21911);
nand UO_2622 (O_2622,N_23421,N_24967);
nand UO_2623 (O_2623,N_23829,N_24236);
nor UO_2624 (O_2624,N_24457,N_22012);
nor UO_2625 (O_2625,N_23144,N_23684);
nor UO_2626 (O_2626,N_20931,N_21310);
nor UO_2627 (O_2627,N_20920,N_24371);
xor UO_2628 (O_2628,N_19937,N_19446);
and UO_2629 (O_2629,N_22744,N_22235);
or UO_2630 (O_2630,N_23841,N_20826);
nor UO_2631 (O_2631,N_21918,N_23976);
and UO_2632 (O_2632,N_20665,N_24184);
and UO_2633 (O_2633,N_19307,N_21879);
nand UO_2634 (O_2634,N_19275,N_19073);
or UO_2635 (O_2635,N_21902,N_22724);
xnor UO_2636 (O_2636,N_21115,N_19269);
xor UO_2637 (O_2637,N_23590,N_23007);
or UO_2638 (O_2638,N_23566,N_21086);
nand UO_2639 (O_2639,N_23816,N_23775);
xnor UO_2640 (O_2640,N_23188,N_23689);
nor UO_2641 (O_2641,N_19898,N_19885);
xnor UO_2642 (O_2642,N_23388,N_23667);
nor UO_2643 (O_2643,N_23969,N_24535);
xor UO_2644 (O_2644,N_21459,N_23999);
or UO_2645 (O_2645,N_19288,N_23743);
nand UO_2646 (O_2646,N_21786,N_22439);
and UO_2647 (O_2647,N_23256,N_18809);
and UO_2648 (O_2648,N_22996,N_19984);
xnor UO_2649 (O_2649,N_24146,N_20878);
and UO_2650 (O_2650,N_24404,N_24577);
and UO_2651 (O_2651,N_19892,N_23742);
and UO_2652 (O_2652,N_23492,N_22558);
xor UO_2653 (O_2653,N_19496,N_21464);
nor UO_2654 (O_2654,N_21167,N_24863);
or UO_2655 (O_2655,N_24484,N_18913);
and UO_2656 (O_2656,N_19524,N_23669);
nand UO_2657 (O_2657,N_22294,N_24269);
xnor UO_2658 (O_2658,N_21741,N_20581);
nor UO_2659 (O_2659,N_20722,N_21499);
xnor UO_2660 (O_2660,N_23326,N_20074);
xor UO_2661 (O_2661,N_21303,N_23960);
and UO_2662 (O_2662,N_24671,N_22386);
and UO_2663 (O_2663,N_24154,N_22987);
and UO_2664 (O_2664,N_23184,N_20197);
nor UO_2665 (O_2665,N_21772,N_19652);
nor UO_2666 (O_2666,N_24108,N_20473);
and UO_2667 (O_2667,N_19574,N_19884);
nand UO_2668 (O_2668,N_20012,N_19027);
nor UO_2669 (O_2669,N_20129,N_19553);
and UO_2670 (O_2670,N_24530,N_23639);
or UO_2671 (O_2671,N_24950,N_18767);
and UO_2672 (O_2672,N_19489,N_19184);
xor UO_2673 (O_2673,N_23585,N_20324);
or UO_2674 (O_2674,N_23521,N_21984);
nand UO_2675 (O_2675,N_22036,N_19001);
nand UO_2676 (O_2676,N_19935,N_20940);
nor UO_2677 (O_2677,N_21289,N_22199);
or UO_2678 (O_2678,N_21407,N_20404);
or UO_2679 (O_2679,N_19422,N_20547);
or UO_2680 (O_2680,N_21929,N_23845);
or UO_2681 (O_2681,N_22611,N_22225);
nand UO_2682 (O_2682,N_21749,N_23955);
nand UO_2683 (O_2683,N_19159,N_21027);
and UO_2684 (O_2684,N_22002,N_22347);
or UO_2685 (O_2685,N_22480,N_22087);
nor UO_2686 (O_2686,N_23102,N_21396);
xor UO_2687 (O_2687,N_22636,N_20687);
nor UO_2688 (O_2688,N_20451,N_20283);
and UO_2689 (O_2689,N_20033,N_20562);
nand UO_2690 (O_2690,N_23325,N_20185);
nand UO_2691 (O_2691,N_21092,N_24896);
xnor UO_2692 (O_2692,N_22321,N_21706);
and UO_2693 (O_2693,N_24581,N_23475);
and UO_2694 (O_2694,N_22319,N_24930);
and UO_2695 (O_2695,N_24304,N_23170);
nand UO_2696 (O_2696,N_19338,N_20456);
or UO_2697 (O_2697,N_24206,N_19862);
and UO_2698 (O_2698,N_21517,N_19530);
nor UO_2699 (O_2699,N_20721,N_20845);
nor UO_2700 (O_2700,N_20663,N_22222);
xor UO_2701 (O_2701,N_19294,N_22063);
nand UO_2702 (O_2702,N_22528,N_21242);
or UO_2703 (O_2703,N_22748,N_19063);
nor UO_2704 (O_2704,N_23119,N_21802);
nor UO_2705 (O_2705,N_23774,N_23635);
or UO_2706 (O_2706,N_20269,N_21476);
nand UO_2707 (O_2707,N_24923,N_20938);
nor UO_2708 (O_2708,N_18987,N_23481);
or UO_2709 (O_2709,N_21990,N_22539);
and UO_2710 (O_2710,N_24644,N_21025);
or UO_2711 (O_2711,N_23296,N_24743);
or UO_2712 (O_2712,N_21541,N_24279);
xnor UO_2713 (O_2713,N_21717,N_21307);
nor UO_2714 (O_2714,N_22484,N_23319);
and UO_2715 (O_2715,N_20556,N_24463);
nand UO_2716 (O_2716,N_22219,N_21002);
nand UO_2717 (O_2717,N_20688,N_20003);
or UO_2718 (O_2718,N_20537,N_23253);
and UO_2719 (O_2719,N_22406,N_21886);
and UO_2720 (O_2720,N_20337,N_20011);
xor UO_2721 (O_2721,N_24738,N_23457);
nand UO_2722 (O_2722,N_23376,N_19348);
or UO_2723 (O_2723,N_21533,N_19569);
or UO_2724 (O_2724,N_18863,N_19736);
xnor UO_2725 (O_2725,N_23101,N_19205);
and UO_2726 (O_2726,N_20108,N_24462);
nor UO_2727 (O_2727,N_21270,N_22379);
nor UO_2728 (O_2728,N_22937,N_20736);
xnor UO_2729 (O_2729,N_20825,N_19815);
and UO_2730 (O_2730,N_22553,N_23896);
nand UO_2731 (O_2731,N_21274,N_21345);
or UO_2732 (O_2732,N_23518,N_24283);
nor UO_2733 (O_2733,N_22848,N_22107);
or UO_2734 (O_2734,N_24062,N_19474);
or UO_2735 (O_2735,N_23291,N_19139);
and UO_2736 (O_2736,N_21158,N_20756);
and UO_2737 (O_2737,N_22778,N_18872);
xnor UO_2738 (O_2738,N_24939,N_21249);
xnor UO_2739 (O_2739,N_21261,N_23533);
xor UO_2740 (O_2740,N_21294,N_20926);
and UO_2741 (O_2741,N_24249,N_23857);
nor UO_2742 (O_2742,N_24017,N_22249);
nand UO_2743 (O_2743,N_20694,N_22248);
xnor UO_2744 (O_2744,N_20302,N_19867);
xor UO_2745 (O_2745,N_20579,N_21264);
and UO_2746 (O_2746,N_21878,N_21818);
nand UO_2747 (O_2747,N_23030,N_19111);
or UO_2748 (O_2748,N_24922,N_20739);
or UO_2749 (O_2749,N_21482,N_21853);
or UO_2750 (O_2750,N_24981,N_24700);
xnor UO_2751 (O_2751,N_23511,N_23272);
xnor UO_2752 (O_2752,N_20170,N_23490);
and UO_2753 (O_2753,N_20774,N_24810);
nor UO_2754 (O_2754,N_19293,N_20416);
nor UO_2755 (O_2755,N_20850,N_22004);
nand UO_2756 (O_2756,N_19087,N_24432);
xnor UO_2757 (O_2757,N_22947,N_23911);
and UO_2758 (O_2758,N_24628,N_19420);
nand UO_2759 (O_2759,N_23071,N_23823);
or UO_2760 (O_2760,N_20914,N_21083);
and UO_2761 (O_2761,N_20975,N_21319);
nand UO_2762 (O_2762,N_19799,N_20488);
and UO_2763 (O_2763,N_23287,N_19791);
xnor UO_2764 (O_2764,N_23342,N_20125);
nand UO_2765 (O_2765,N_22113,N_20840);
nand UO_2766 (O_2766,N_24795,N_20462);
nand UO_2767 (O_2767,N_24054,N_20832);
nor UO_2768 (O_2768,N_19516,N_22827);
and UO_2769 (O_2769,N_22981,N_23172);
xor UO_2770 (O_2770,N_19507,N_21046);
xor UO_2771 (O_2771,N_20600,N_24734);
nand UO_2772 (O_2772,N_24942,N_24997);
xor UO_2773 (O_2773,N_20573,N_24171);
nand UO_2774 (O_2774,N_22972,N_22388);
or UO_2775 (O_2775,N_20236,N_22904);
and UO_2776 (O_2776,N_22176,N_19662);
and UO_2777 (O_2777,N_19078,N_20900);
or UO_2778 (O_2778,N_21431,N_24306);
or UO_2779 (O_2779,N_19104,N_23824);
xor UO_2780 (O_2780,N_21075,N_22105);
xnor UO_2781 (O_2781,N_23000,N_22629);
and UO_2782 (O_2782,N_22099,N_24258);
xnor UO_2783 (O_2783,N_21994,N_23847);
xnor UO_2784 (O_2784,N_24376,N_24129);
nor UO_2785 (O_2785,N_19490,N_23016);
nor UO_2786 (O_2786,N_24874,N_20389);
xor UO_2787 (O_2787,N_22735,N_19448);
xor UO_2788 (O_2788,N_24144,N_24899);
nor UO_2789 (O_2789,N_18954,N_22366);
and UO_2790 (O_2790,N_22929,N_21910);
xnor UO_2791 (O_2791,N_22124,N_21980);
and UO_2792 (O_2792,N_22436,N_23399);
nor UO_2793 (O_2793,N_21032,N_21613);
xor UO_2794 (O_2794,N_22242,N_19985);
nand UO_2795 (O_2795,N_20752,N_21450);
or UO_2796 (O_2796,N_24487,N_18985);
or UO_2797 (O_2797,N_23631,N_24272);
and UO_2798 (O_2798,N_24906,N_23529);
or UO_2799 (O_2799,N_19250,N_24789);
nand UO_2800 (O_2800,N_21584,N_24596);
or UO_2801 (O_2801,N_24152,N_24033);
or UO_2802 (O_2802,N_19506,N_23813);
or UO_2803 (O_2803,N_24851,N_19958);
nor UO_2804 (O_2804,N_19360,N_20059);
xnor UO_2805 (O_2805,N_22923,N_24105);
or UO_2806 (O_2806,N_20943,N_20371);
or UO_2807 (O_2807,N_20017,N_21362);
nand UO_2808 (O_2808,N_20037,N_19118);
xor UO_2809 (O_2809,N_21140,N_19120);
nor UO_2810 (O_2810,N_23729,N_20963);
nor UO_2811 (O_2811,N_24210,N_20342);
nor UO_2812 (O_2812,N_19090,N_19208);
or UO_2813 (O_2813,N_24049,N_23872);
or UO_2814 (O_2814,N_21797,N_24290);
xor UO_2815 (O_2815,N_24451,N_19796);
and UO_2816 (O_2816,N_23357,N_24859);
nor UO_2817 (O_2817,N_23316,N_19986);
and UO_2818 (O_2818,N_23990,N_23584);
and UO_2819 (O_2819,N_23354,N_20309);
xnor UO_2820 (O_2820,N_23815,N_24270);
nor UO_2821 (O_2821,N_20237,N_19177);
or UO_2822 (O_2822,N_24636,N_23656);
nor UO_2823 (O_2823,N_19503,N_24669);
nand UO_2824 (O_2824,N_23467,N_22793);
and UO_2825 (O_2825,N_20164,N_19371);
nor UO_2826 (O_2826,N_20490,N_24776);
or UO_2827 (O_2827,N_21698,N_20216);
or UO_2828 (O_2828,N_23026,N_24394);
and UO_2829 (O_2829,N_20116,N_21838);
xnor UO_2830 (O_2830,N_20104,N_24427);
xor UO_2831 (O_2831,N_19213,N_24099);
xnor UO_2832 (O_2832,N_19352,N_24841);
nor UO_2833 (O_2833,N_21958,N_19246);
and UO_2834 (O_2834,N_24589,N_20167);
xnor UO_2835 (O_2835,N_21787,N_20292);
nor UO_2836 (O_2836,N_20006,N_19463);
xor UO_2837 (O_2837,N_22329,N_21399);
nand UO_2838 (O_2838,N_22775,N_22666);
or UO_2839 (O_2839,N_24913,N_23978);
and UO_2840 (O_2840,N_18820,N_20856);
or UO_2841 (O_2841,N_23702,N_24316);
xor UO_2842 (O_2842,N_19831,N_24905);
xor UO_2843 (O_2843,N_19375,N_24234);
xor UO_2844 (O_2844,N_20534,N_21102);
or UO_2845 (O_2845,N_18944,N_19002);
nand UO_2846 (O_2846,N_23515,N_21933);
or UO_2847 (O_2847,N_23860,N_23692);
and UO_2848 (O_2848,N_24158,N_23734);
xnor UO_2849 (O_2849,N_20439,N_24825);
xnor UO_2850 (O_2850,N_23951,N_20817);
nor UO_2851 (O_2851,N_21914,N_21391);
nor UO_2852 (O_2852,N_19887,N_24542);
xnor UO_2853 (O_2853,N_23254,N_20961);
nor UO_2854 (O_2854,N_20143,N_22410);
nand UO_2855 (O_2855,N_22939,N_19110);
or UO_2856 (O_2856,N_22999,N_23660);
and UO_2857 (O_2857,N_21331,N_19498);
and UO_2858 (O_2858,N_22237,N_21595);
nor UO_2859 (O_2859,N_23304,N_24661);
and UO_2860 (O_2860,N_20771,N_24297);
nor UO_2861 (O_2861,N_23169,N_19708);
and UO_2862 (O_2862,N_21368,N_24796);
nand UO_2863 (O_2863,N_19999,N_21783);
nor UO_2864 (O_2864,N_19538,N_19058);
xor UO_2865 (O_2865,N_21253,N_21774);
xnor UO_2866 (O_2866,N_19030,N_23150);
and UO_2867 (O_2867,N_21378,N_22993);
xnor UO_2868 (O_2868,N_18907,N_19829);
or UO_2869 (O_2869,N_22725,N_22206);
and UO_2870 (O_2870,N_21701,N_22658);
nor UO_2871 (O_2871,N_19977,N_20042);
nor UO_2872 (O_2872,N_20994,N_21883);
nand UO_2873 (O_2873,N_20548,N_22821);
or UO_2874 (O_2874,N_24040,N_21645);
nor UO_2875 (O_2875,N_24245,N_24600);
or UO_2876 (O_2876,N_22368,N_22717);
or UO_2877 (O_2877,N_22538,N_23403);
xor UO_2878 (O_2878,N_21172,N_19309);
nor UO_2879 (O_2879,N_24838,N_19936);
nor UO_2880 (O_2880,N_22575,N_19637);
xnor UO_2881 (O_2881,N_21444,N_21348);
nand UO_2882 (O_2882,N_19094,N_24307);
nand UO_2883 (O_2883,N_23968,N_23893);
or UO_2884 (O_2884,N_21942,N_19600);
and UO_2885 (O_2885,N_22007,N_20482);
and UO_2886 (O_2886,N_22928,N_24031);
nand UO_2887 (O_2887,N_23196,N_20420);
xnor UO_2888 (O_2888,N_24318,N_20249);
nor UO_2889 (O_2889,N_22768,N_20045);
xnor UO_2890 (O_2890,N_20428,N_21840);
and UO_2891 (O_2891,N_20120,N_18936);
nand UO_2892 (O_2892,N_20919,N_24322);
nor UO_2893 (O_2893,N_19666,N_20138);
nand UO_2894 (O_2894,N_22109,N_22323);
xor UO_2895 (O_2895,N_19500,N_19437);
or UO_2896 (O_2896,N_19028,N_23874);
or UO_2897 (O_2897,N_22894,N_24113);
xnor UO_2898 (O_2898,N_21397,N_24682);
nor UO_2899 (O_2899,N_20505,N_19056);
xor UO_2900 (O_2900,N_23429,N_18966);
nor UO_2901 (O_2901,N_23888,N_23777);
and UO_2902 (O_2902,N_21068,N_23269);
or UO_2903 (O_2903,N_23113,N_21309);
or UO_2904 (O_2904,N_22835,N_23618);
and UO_2905 (O_2905,N_21291,N_21398);
nand UO_2906 (O_2906,N_22696,N_19608);
and UO_2907 (O_2907,N_20221,N_23208);
nor UO_2908 (O_2908,N_22381,N_19065);
nand UO_2909 (O_2909,N_20670,N_21422);
nand UO_2910 (O_2910,N_20555,N_23666);
nor UO_2911 (O_2911,N_18947,N_19581);
or UO_2912 (O_2912,N_23744,N_21551);
nor UO_2913 (O_2913,N_22537,N_24362);
or UO_2914 (O_2914,N_22690,N_20819);
xor UO_2915 (O_2915,N_23817,N_24965);
and UO_2916 (O_2916,N_23750,N_20716);
or UO_2917 (O_2917,N_22573,N_24500);
nand UO_2918 (O_2918,N_24768,N_19173);
xor UO_2919 (O_2919,N_19025,N_20498);
xnor UO_2920 (O_2920,N_19400,N_21461);
or UO_2921 (O_2921,N_23162,N_19356);
or UO_2922 (O_2922,N_24199,N_21830);
nor UO_2923 (O_2923,N_22952,N_24961);
and UO_2924 (O_2924,N_24886,N_20540);
or UO_2925 (O_2925,N_22534,N_23931);
or UO_2926 (O_2926,N_23092,N_21493);
and UO_2927 (O_2927,N_21862,N_22115);
nand UO_2928 (O_2928,N_23166,N_23505);
nor UO_2929 (O_2929,N_20491,N_22901);
or UO_2930 (O_2930,N_22649,N_22560);
nor UO_2931 (O_2931,N_24391,N_19199);
nand UO_2932 (O_2932,N_20122,N_24354);
nor UO_2933 (O_2933,N_24390,N_23718);
and UO_2934 (O_2934,N_23977,N_19990);
nand UO_2935 (O_2935,N_20182,N_22441);
or UO_2936 (O_2936,N_19358,N_24004);
nor UO_2937 (O_2937,N_21030,N_21424);
or UO_2938 (O_2938,N_19165,N_22828);
xnor UO_2939 (O_2939,N_23916,N_19906);
xnor UO_2940 (O_2940,N_19133,N_21286);
and UO_2941 (O_2941,N_19318,N_19234);
nor UO_2942 (O_2942,N_23613,N_20435);
nor UO_2943 (O_2943,N_24999,N_20010);
nand UO_2944 (O_2944,N_19433,N_22685);
and UO_2945 (O_2945,N_19099,N_21849);
or UO_2946 (O_2946,N_20118,N_19421);
xnor UO_2947 (O_2947,N_23838,N_24015);
xor UO_2948 (O_2948,N_21212,N_21810);
xor UO_2949 (O_2949,N_22260,N_24501);
nand UO_2950 (O_2950,N_24264,N_19154);
nor UO_2951 (O_2951,N_18846,N_24072);
and UO_2952 (O_2952,N_19732,N_22174);
xor UO_2953 (O_2953,N_22507,N_18868);
and UO_2954 (O_2954,N_23081,N_19158);
nand UO_2955 (O_2955,N_23904,N_21737);
xor UO_2956 (O_2956,N_19174,N_18885);
nor UO_2957 (O_2957,N_18920,N_24205);
nor UO_2958 (O_2958,N_20655,N_19692);
xnor UO_2959 (O_2959,N_22810,N_23294);
nor UO_2960 (O_2960,N_21338,N_20409);
nor UO_2961 (O_2961,N_19068,N_24759);
and UO_2962 (O_2962,N_24928,N_24881);
nand UO_2963 (O_2963,N_22274,N_20906);
xor UO_2964 (O_2964,N_19991,N_21428);
or UO_2965 (O_2965,N_19908,N_21971);
nand UO_2966 (O_2966,N_22234,N_21566);
or UO_2967 (O_2967,N_21204,N_24747);
and UO_2968 (O_2968,N_24590,N_22586);
nand UO_2969 (O_2969,N_23646,N_24314);
nand UO_2970 (O_2970,N_23678,N_23343);
and UO_2971 (O_2971,N_23241,N_21262);
and UO_2972 (O_2972,N_19067,N_19200);
xnor UO_2973 (O_2973,N_22120,N_23135);
or UO_2974 (O_2974,N_23310,N_22187);
nand UO_2975 (O_2975,N_23221,N_19414);
and UO_2976 (O_2976,N_22647,N_20993);
nor UO_2977 (O_2977,N_18956,N_21596);
and UO_2978 (O_2978,N_20730,N_20395);
or UO_2979 (O_2979,N_20623,N_19450);
nand UO_2980 (O_2980,N_20580,N_18784);
xnor UO_2981 (O_2981,N_24330,N_21076);
or UO_2982 (O_2982,N_20169,N_21553);
or UO_2983 (O_2983,N_24723,N_19960);
xnor UO_2984 (O_2984,N_20871,N_23341);
nand UO_2985 (O_2985,N_24185,N_20508);
xnor UO_2986 (O_2986,N_21540,N_20075);
and UO_2987 (O_2987,N_24757,N_22361);
xnor UO_2988 (O_2988,N_24214,N_19136);
nor UO_2989 (O_2989,N_20657,N_21053);
and UO_2990 (O_2990,N_22799,N_23846);
xor UO_2991 (O_2991,N_20311,N_23124);
or UO_2992 (O_2992,N_21221,N_24742);
and UO_2993 (O_2993,N_24642,N_22330);
xor UO_2994 (O_2994,N_19683,N_21443);
xor UO_2995 (O_2995,N_21487,N_21716);
nor UO_2996 (O_2996,N_20827,N_24651);
and UO_2997 (O_2997,N_20332,N_24709);
nor UO_2998 (O_2998,N_23411,N_21627);
nand UO_2999 (O_2999,N_22048,N_19918);
endmodule