module basic_1500_15000_2000_75_levels_5xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
and U0 (N_0,In_858,In_111);
nand U1 (N_1,In_488,In_967);
or U2 (N_2,In_708,In_299);
and U3 (N_3,In_374,In_1078);
nor U4 (N_4,In_674,In_1275);
nor U5 (N_5,In_436,In_1285);
nand U6 (N_6,In_493,In_127);
nor U7 (N_7,In_1296,In_52);
nor U8 (N_8,In_54,In_514);
or U9 (N_9,In_1211,In_318);
nand U10 (N_10,In_139,In_1276);
nand U11 (N_11,In_762,In_1066);
nor U12 (N_12,In_581,In_1373);
nand U13 (N_13,In_504,In_924);
xnor U14 (N_14,In_480,In_1171);
nand U15 (N_15,In_1112,In_1083);
nor U16 (N_16,In_1011,In_198);
nor U17 (N_17,In_979,In_1407);
and U18 (N_18,In_1186,In_1352);
nand U19 (N_19,In_1201,In_178);
nor U20 (N_20,In_60,In_1333);
nor U21 (N_21,In_175,In_78);
xnor U22 (N_22,In_614,In_1154);
xnor U23 (N_23,In_471,In_664);
or U24 (N_24,In_15,In_1479);
and U25 (N_25,In_770,In_67);
nor U26 (N_26,In_756,In_499);
and U27 (N_27,In_919,In_397);
nor U28 (N_28,In_1239,In_1376);
and U29 (N_29,In_387,In_1484);
nor U30 (N_30,In_112,In_317);
nand U31 (N_31,In_1458,In_775);
nand U32 (N_32,In_264,In_752);
nor U33 (N_33,In_587,In_1172);
xnor U34 (N_34,In_974,In_865);
or U35 (N_35,In_1013,In_246);
xor U36 (N_36,In_1072,In_1055);
nor U37 (N_37,In_1430,In_764);
nand U38 (N_38,In_177,In_834);
nand U39 (N_39,In_12,In_721);
nand U40 (N_40,In_599,In_757);
and U41 (N_41,In_70,In_1393);
nand U42 (N_42,In_446,In_853);
and U43 (N_43,In_870,In_1232);
and U44 (N_44,In_204,In_972);
xor U45 (N_45,In_960,In_1203);
nand U46 (N_46,In_359,In_1104);
nand U47 (N_47,In_1018,In_1130);
or U48 (N_48,In_1400,In_107);
nand U49 (N_49,In_1480,In_569);
and U50 (N_50,In_19,In_791);
nor U51 (N_51,In_1127,In_658);
and U52 (N_52,In_63,In_1085);
or U53 (N_53,In_1418,In_975);
and U54 (N_54,In_1194,In_650);
or U55 (N_55,In_1428,In_1271);
and U56 (N_56,In_508,In_633);
and U57 (N_57,In_478,In_1037);
xnor U58 (N_58,In_273,In_1249);
and U59 (N_59,In_882,In_49);
or U60 (N_60,In_638,In_659);
or U61 (N_61,In_606,In_567);
or U62 (N_62,In_404,In_193);
nor U63 (N_63,In_1036,In_1310);
or U64 (N_64,In_460,In_794);
nor U65 (N_65,In_302,In_6);
or U66 (N_66,In_1297,In_711);
xnor U67 (N_67,In_1485,In_1354);
and U68 (N_68,In_535,In_1410);
xnor U69 (N_69,In_219,In_339);
nor U70 (N_70,In_1422,In_56);
nor U71 (N_71,In_1216,In_947);
nor U72 (N_72,In_1187,In_877);
and U73 (N_73,In_1348,In_951);
or U74 (N_74,In_1394,In_1382);
nand U75 (N_75,In_32,In_451);
and U76 (N_76,In_984,In_211);
and U77 (N_77,In_398,In_1176);
and U78 (N_78,In_630,In_83);
or U79 (N_79,In_114,In_1489);
nor U80 (N_80,In_1145,In_985);
or U81 (N_81,In_811,In_992);
nor U82 (N_82,In_701,In_1291);
or U83 (N_83,In_1375,In_513);
and U84 (N_84,In_526,In_323);
xor U85 (N_85,In_706,In_553);
nand U86 (N_86,In_242,In_1007);
and U87 (N_87,In_529,In_1160);
and U88 (N_88,In_133,In_640);
xor U89 (N_89,In_1498,In_1295);
and U90 (N_90,In_1027,In_420);
nand U91 (N_91,In_1284,In_872);
and U92 (N_92,In_332,In_199);
and U93 (N_93,In_1258,In_407);
nand U94 (N_94,In_11,In_416);
or U95 (N_95,In_1487,In_132);
nor U96 (N_96,In_1222,In_733);
nor U97 (N_97,In_1371,In_522);
nand U98 (N_98,In_86,In_266);
and U99 (N_99,In_466,In_1123);
or U100 (N_100,In_244,In_1425);
or U101 (N_101,In_572,In_1157);
nand U102 (N_102,In_682,In_169);
xor U103 (N_103,In_697,In_341);
and U104 (N_104,In_1454,In_1341);
and U105 (N_105,In_53,In_851);
nand U106 (N_106,In_1286,In_87);
nor U107 (N_107,In_176,In_262);
nor U108 (N_108,In_540,In_482);
or U109 (N_109,In_855,In_886);
nand U110 (N_110,In_863,In_1357);
nand U111 (N_111,In_0,In_1319);
nand U112 (N_112,In_1260,In_552);
nor U113 (N_113,In_425,In_1327);
or U114 (N_114,In_51,In_1469);
nor U115 (N_115,In_1241,In_1263);
or U116 (N_116,In_124,In_1240);
or U117 (N_117,In_964,In_402);
and U118 (N_118,In_427,In_996);
and U119 (N_119,In_1195,In_1220);
nor U120 (N_120,In_563,In_597);
and U121 (N_121,In_754,In_1265);
nor U122 (N_122,In_767,In_517);
xor U123 (N_123,In_1045,In_26);
and U124 (N_124,In_673,In_1251);
or U125 (N_125,In_386,In_932);
and U126 (N_126,In_1390,In_1218);
and U127 (N_127,In_434,In_278);
nor U128 (N_128,In_1046,In_1330);
nor U129 (N_129,In_1229,In_835);
xnor U130 (N_130,In_1381,In_1126);
nor U131 (N_131,In_1206,In_604);
nor U132 (N_132,In_1465,In_1403);
nand U133 (N_133,In_9,In_1169);
nor U134 (N_134,In_941,In_1438);
xor U135 (N_135,In_1415,In_1196);
or U136 (N_136,In_1064,In_761);
and U137 (N_137,In_667,In_350);
nor U138 (N_138,In_660,In_1001);
and U139 (N_139,In_376,In_953);
and U140 (N_140,In_525,In_1101);
nor U141 (N_141,In_825,In_852);
or U142 (N_142,In_342,In_443);
and U143 (N_143,In_1247,In_1017);
or U144 (N_144,In_269,In_636);
or U145 (N_145,In_691,In_934);
xor U146 (N_146,In_248,In_827);
nor U147 (N_147,In_1414,In_1308);
or U148 (N_148,In_1496,In_1050);
xnor U149 (N_149,In_605,In_785);
and U150 (N_150,In_889,In_1237);
nor U151 (N_151,In_410,In_275);
nor U152 (N_152,In_497,In_685);
nand U153 (N_153,In_698,In_27);
or U154 (N_154,In_1019,In_681);
nor U155 (N_155,In_334,In_430);
and U156 (N_156,In_356,In_362);
and U157 (N_157,In_729,In_908);
or U158 (N_158,In_710,In_1384);
nand U159 (N_159,In_120,In_1113);
nand U160 (N_160,In_654,In_705);
nor U161 (N_161,In_655,In_837);
or U162 (N_162,In_896,In_195);
nor U163 (N_163,In_530,In_1067);
nor U164 (N_164,In_1213,In_1490);
nor U165 (N_165,In_1267,In_1230);
nand U166 (N_166,In_1141,In_282);
nand U167 (N_167,In_1315,In_349);
nand U168 (N_168,In_609,In_1168);
and U169 (N_169,In_768,In_1289);
xnor U170 (N_170,In_38,In_1316);
xnor U171 (N_171,In_907,In_914);
and U172 (N_172,In_348,In_848);
or U173 (N_173,In_294,In_527);
or U174 (N_174,In_720,In_629);
xor U175 (N_175,In_40,In_1452);
nand U176 (N_176,In_329,In_208);
nor U177 (N_177,In_783,In_714);
nor U178 (N_178,In_18,In_142);
nand U179 (N_179,In_939,In_1214);
nand U180 (N_180,In_557,In_417);
and U181 (N_181,In_1069,In_122);
nand U182 (N_182,In_779,In_1223);
or U183 (N_183,In_1137,In_1132);
nand U184 (N_184,In_218,In_447);
nand U185 (N_185,In_676,In_31);
and U186 (N_186,In_1334,In_1307);
nor U187 (N_187,In_615,In_1227);
nor U188 (N_188,In_959,In_977);
and U189 (N_189,In_212,In_113);
nor U190 (N_190,In_1252,In_1235);
nor U191 (N_191,In_1389,In_73);
nor U192 (N_192,In_399,In_608);
nor U193 (N_193,In_247,In_707);
nand U194 (N_194,In_1000,In_930);
xor U195 (N_195,In_223,In_1298);
nor U196 (N_196,In_295,In_116);
and U197 (N_197,In_1099,In_744);
or U198 (N_198,In_1383,In_206);
and U199 (N_199,In_438,In_442);
and U200 (N_200,In_945,N_186);
nor U201 (N_201,In_158,In_869);
nor U202 (N_202,N_88,In_675);
or U203 (N_203,In_1362,In_841);
nand U204 (N_204,N_10,In_415);
xor U205 (N_205,In_988,In_1110);
xnor U206 (N_206,In_1379,In_566);
nor U207 (N_207,In_452,In_281);
xnor U208 (N_208,In_467,In_1444);
and U209 (N_209,In_575,In_243);
nand U210 (N_210,In_487,N_85);
nand U211 (N_211,In_1365,In_888);
nor U212 (N_212,In_732,In_36);
and U213 (N_213,In_1287,In_276);
and U214 (N_214,In_1153,N_95);
or U215 (N_215,In_821,In_766);
nand U216 (N_216,In_946,In_1256);
nand U217 (N_217,In_680,In_1329);
and U218 (N_218,In_81,In_210);
or U219 (N_219,In_47,In_1035);
nand U220 (N_220,In_1208,In_343);
nor U221 (N_221,In_782,In_815);
and U222 (N_222,In_1148,N_135);
xnor U223 (N_223,In_465,In_618);
xor U224 (N_224,In_1445,In_1059);
or U225 (N_225,In_621,In_1009);
nand U226 (N_226,In_1369,In_383);
and U227 (N_227,In_453,In_290);
nand U228 (N_228,In_289,In_700);
or U229 (N_229,In_965,N_108);
nand U230 (N_230,In_74,N_194);
nand U231 (N_231,N_40,In_1047);
nor U232 (N_232,N_31,In_33);
nand U233 (N_233,In_1156,N_53);
or U234 (N_234,In_653,In_601);
nand U235 (N_235,In_469,In_412);
nand U236 (N_236,In_1257,In_309);
and U237 (N_237,In_920,In_997);
or U238 (N_238,In_1468,In_1108);
or U239 (N_239,In_1399,In_1086);
nor U240 (N_240,In_1093,In_89);
and U241 (N_241,In_578,N_134);
nand U242 (N_242,In_82,In_335);
and U243 (N_243,N_75,In_1255);
and U244 (N_244,In_265,In_123);
or U245 (N_245,In_333,In_652);
xor U246 (N_246,N_94,In_1022);
nand U247 (N_247,In_311,In_925);
nand U248 (N_248,In_1455,In_1314);
nor U249 (N_249,In_1309,In_1277);
nand U250 (N_250,N_137,N_97);
nand U251 (N_251,In_856,In_980);
nand U252 (N_252,In_742,N_91);
nand U253 (N_253,In_331,N_106);
nor U254 (N_254,In_117,In_885);
nand U255 (N_255,In_506,In_1177);
and U256 (N_256,In_320,In_65);
xnor U257 (N_257,In_121,In_136);
xnor U258 (N_258,In_1014,In_439);
and U259 (N_259,In_91,N_0);
and U260 (N_260,N_138,In_1225);
nor U261 (N_261,In_401,N_26);
xor U262 (N_262,In_995,N_165);
or U263 (N_263,In_160,In_626);
xor U264 (N_264,In_406,In_804);
and U265 (N_265,N_49,N_67);
and U266 (N_266,In_1139,In_35);
nand U267 (N_267,In_1340,In_814);
nand U268 (N_268,N_157,In_1272);
xnor U269 (N_269,In_1170,In_695);
and U270 (N_270,In_1005,In_1401);
nand U271 (N_271,In_641,In_1446);
nor U272 (N_272,In_735,N_146);
or U273 (N_273,N_19,In_379);
and U274 (N_274,In_183,N_16);
nor U275 (N_275,In_983,In_1121);
and U276 (N_276,In_1106,In_5);
nand U277 (N_277,N_112,In_892);
and U278 (N_278,In_981,In_363);
or U279 (N_279,In_392,In_1448);
and U280 (N_280,In_923,In_725);
nand U281 (N_281,In_1424,In_1337);
nand U282 (N_282,In_890,In_125);
or U283 (N_283,N_87,In_1356);
or U284 (N_284,In_973,In_303);
xnor U285 (N_285,In_229,In_1317);
and U286 (N_286,In_1482,In_915);
nor U287 (N_287,In_1070,In_1417);
or U288 (N_288,N_158,In_1461);
and U289 (N_289,N_61,In_1450);
nor U290 (N_290,In_207,N_71);
or U291 (N_291,In_666,In_879);
nor U292 (N_292,N_188,In_291);
and U293 (N_293,In_164,In_489);
and U294 (N_294,N_11,In_1081);
xor U295 (N_295,In_153,N_96);
or U296 (N_296,In_1435,In_131);
or U297 (N_297,In_190,N_178);
nor U298 (N_298,In_1456,In_393);
and U299 (N_299,In_135,In_1486);
xor U300 (N_300,In_1494,In_267);
or U301 (N_301,In_424,In_1044);
nor U302 (N_302,In_819,In_472);
nor U303 (N_303,N_84,In_679);
nor U304 (N_304,In_632,In_95);
or U305 (N_305,N_99,In_194);
or U306 (N_306,In_1140,In_651);
nand U307 (N_307,In_272,In_1440);
nor U308 (N_308,N_51,In_1002);
or U309 (N_309,In_1060,In_554);
or U310 (N_310,In_1161,In_454);
and U311 (N_311,N_7,In_1421);
and U312 (N_312,In_481,In_1388);
and U313 (N_313,In_458,In_617);
nor U314 (N_314,In_22,In_871);
xor U315 (N_315,In_1248,N_145);
nand U316 (N_316,In_1056,In_646);
or U317 (N_317,In_357,In_507);
or U318 (N_318,In_1408,In_881);
nor U319 (N_319,In_1491,N_43);
or U320 (N_320,In_620,In_778);
or U321 (N_321,In_1398,In_1133);
or U322 (N_322,In_68,In_531);
or U323 (N_323,In_1413,In_1462);
nand U324 (N_324,In_304,In_486);
or U325 (N_325,In_1420,In_337);
nor U326 (N_326,In_585,In_790);
and U327 (N_327,In_1097,In_1473);
nand U328 (N_328,In_991,In_296);
or U329 (N_329,In_71,In_928);
or U330 (N_330,In_820,In_683);
xor U331 (N_331,N_77,In_1396);
nor U332 (N_332,N_92,In_1167);
and U333 (N_333,In_799,N_5);
nor U334 (N_334,In_798,In_186);
nor U335 (N_335,In_1025,In_986);
or U336 (N_336,In_1074,In_565);
nor U337 (N_337,N_143,In_548);
nand U338 (N_338,In_564,N_109);
nand U339 (N_339,N_192,In_1499);
or U340 (N_340,In_1320,In_1336);
nor U341 (N_341,In_812,In_222);
and U342 (N_342,In_1326,In_1439);
and U343 (N_343,In_1366,N_4);
nor U344 (N_344,In_382,In_561);
nor U345 (N_345,In_396,In_774);
nand U346 (N_346,In_1049,In_909);
or U347 (N_347,In_878,In_969);
xnor U348 (N_348,In_1301,In_631);
or U349 (N_349,In_373,N_191);
nand U350 (N_350,In_280,In_464);
nand U351 (N_351,In_904,In_255);
or U352 (N_352,In_1311,In_1135);
xor U353 (N_353,In_1449,In_101);
and U354 (N_354,In_740,In_763);
and U355 (N_355,In_105,In_976);
xor U356 (N_356,In_760,In_254);
nand U357 (N_357,In_80,In_1178);
and U358 (N_358,In_1183,In_1395);
nor U359 (N_359,In_408,In_1224);
or U360 (N_360,In_712,In_639);
and U361 (N_361,In_1463,In_583);
nand U362 (N_362,N_25,In_168);
nor U363 (N_363,N_60,In_1345);
and U364 (N_364,In_1142,N_142);
nor U365 (N_365,N_156,In_1098);
nor U366 (N_366,In_1269,N_149);
nand U367 (N_367,In_106,In_1155);
nand U368 (N_368,In_916,In_954);
nand U369 (N_369,In_839,In_780);
nand U370 (N_370,In_1210,In_1084);
nand U371 (N_371,In_927,In_1124);
nor U372 (N_372,In_665,In_477);
nor U373 (N_373,In_1350,In_419);
nor U374 (N_374,In_702,In_816);
nand U375 (N_375,In_1054,N_41);
xor U376 (N_376,In_251,In_900);
nor U377 (N_377,In_1109,In_994);
or U378 (N_378,In_786,In_543);
nand U379 (N_379,N_78,In_781);
nor U380 (N_380,In_491,In_360);
nor U381 (N_381,In_344,In_592);
or U382 (N_382,In_968,In_370);
xnor U383 (N_383,In_1058,In_1483);
or U384 (N_384,In_1434,In_1380);
nand U385 (N_385,In_1282,In_802);
or U386 (N_386,In_1219,In_1117);
nand U387 (N_387,In_1175,In_1472);
nand U388 (N_388,In_693,In_1368);
nand U389 (N_389,In_824,In_703);
and U390 (N_390,In_1377,In_388);
nand U391 (N_391,In_358,In_25);
nand U392 (N_392,In_421,In_365);
nand U393 (N_393,In_538,In_738);
or U394 (N_394,N_98,N_34);
xor U395 (N_395,In_669,In_1231);
nor U396 (N_396,In_836,In_978);
nor U397 (N_397,In_672,In_79);
nor U398 (N_398,In_542,In_1023);
nor U399 (N_399,In_509,In_428);
xnor U400 (N_400,In_233,N_361);
nand U401 (N_401,In_637,In_1071);
nor U402 (N_402,In_913,N_340);
nor U403 (N_403,In_433,In_1063);
nand U404 (N_404,In_999,N_316);
or U405 (N_405,N_330,N_128);
or U406 (N_406,In_2,In_94);
and U407 (N_407,N_246,In_1331);
nand U408 (N_408,N_235,N_327);
or U409 (N_409,In_312,N_333);
nor U410 (N_410,N_66,N_162);
and U411 (N_411,In_769,In_1464);
xnor U412 (N_412,In_745,N_254);
or U413 (N_413,In_950,In_1051);
nand U414 (N_414,N_177,In_203);
and U415 (N_415,In_474,N_351);
nand U416 (N_416,In_1385,In_643);
nor U417 (N_417,N_386,N_141);
nand U418 (N_418,In_143,In_861);
nor U419 (N_419,In_1245,In_456);
nand U420 (N_420,In_1115,N_275);
or U421 (N_421,In_1323,In_1300);
or U422 (N_422,N_306,N_369);
or U423 (N_423,N_189,In_1039);
nor U424 (N_424,In_361,N_8);
or U425 (N_425,In_1073,In_319);
or U426 (N_426,N_317,In_759);
nor U427 (N_427,N_133,In_1404);
nand U428 (N_428,N_353,N_310);
xor U429 (N_429,In_301,N_270);
nor U430 (N_430,N_181,N_394);
nor U431 (N_431,N_115,In_796);
xnor U432 (N_432,In_895,In_1259);
or U433 (N_433,In_511,N_166);
and U434 (N_434,In_805,In_724);
and U435 (N_435,In_1200,In_1033);
or U436 (N_436,In_671,N_287);
and U437 (N_437,In_34,In_1144);
nor U438 (N_438,In_1147,In_263);
nor U439 (N_439,In_730,In_1402);
nand U440 (N_440,N_116,N_121);
nor U441 (N_441,N_171,In_364);
or U442 (N_442,In_1163,In_944);
and U443 (N_443,In_1378,N_218);
and U444 (N_444,In_1409,In_1338);
and U445 (N_445,In_165,N_315);
nor U446 (N_446,In_149,In_670);
nor U447 (N_447,In_10,In_1159);
or U448 (N_448,In_822,In_1192);
and U449 (N_449,In_126,In_1152);
or U450 (N_450,In_1497,In_1467);
nor U451 (N_451,In_1433,In_1303);
nand U452 (N_452,In_613,N_379);
nand U453 (N_453,In_1181,N_104);
nand U454 (N_454,In_315,N_212);
nand U455 (N_455,In_128,In_846);
or U456 (N_456,In_515,N_349);
nand U457 (N_457,N_329,N_339);
and U458 (N_458,In_64,In_1038);
nand U459 (N_459,In_1228,In_205);
and U460 (N_460,In_1460,N_263);
and U461 (N_461,In_152,In_1416);
nor U462 (N_462,N_314,In_1191);
nor U463 (N_463,In_1205,N_389);
nand U464 (N_464,In_1335,In_518);
and U465 (N_465,N_262,In_445);
or U466 (N_466,In_536,In_550);
nand U467 (N_467,N_13,In_899);
nor U468 (N_468,In_524,N_291);
or U469 (N_469,In_297,In_906);
or U470 (N_470,In_189,In_69);
nor U471 (N_471,In_375,N_110);
nor U472 (N_472,N_341,In_298);
or U473 (N_473,In_1092,In_957);
or U474 (N_474,In_1328,In_268);
nand U475 (N_475,In_1077,N_240);
and U476 (N_476,N_324,In_832);
nor U477 (N_477,In_562,In_1114);
and U478 (N_478,In_501,In_336);
and U479 (N_479,In_1026,N_163);
xor U480 (N_480,In_1242,In_455);
nand U481 (N_481,In_505,In_103);
xnor U482 (N_482,In_1080,N_344);
and U483 (N_483,In_612,In_772);
and U484 (N_484,In_868,N_174);
nor U485 (N_485,N_23,In_926);
nand U486 (N_486,In_351,In_173);
or U487 (N_487,In_39,In_558);
or U488 (N_488,In_1179,In_305);
and U489 (N_489,N_29,In_1164);
nand U490 (N_490,N_55,N_39);
and U491 (N_491,In_118,In_731);
or U492 (N_492,N_46,In_284);
or U493 (N_493,In_849,In_75);
and U494 (N_494,N_323,In_661);
nor U495 (N_495,In_1305,N_33);
nor U496 (N_496,In_1094,In_4);
or U497 (N_497,In_476,In_338);
xor U498 (N_498,In_1016,In_624);
and U499 (N_499,N_368,In_1279);
and U500 (N_500,N_136,In_239);
nand U501 (N_501,N_86,In_854);
nand U502 (N_502,In_833,N_73);
or U503 (N_503,In_1339,In_100);
or U504 (N_504,N_155,In_1089);
xor U505 (N_505,In_145,In_1427);
nand U506 (N_506,In_635,In_391);
and U507 (N_507,In_1,N_318);
or U508 (N_508,In_547,N_366);
nand U509 (N_509,In_174,In_286);
and U510 (N_510,N_154,In_789);
or U511 (N_511,In_129,In_503);
nand U512 (N_512,In_450,In_1244);
and U513 (N_513,In_747,In_45);
xnor U514 (N_514,In_314,In_746);
and U515 (N_515,N_117,N_200);
or U516 (N_516,In_277,In_459);
or U517 (N_517,In_656,N_325);
xor U518 (N_518,In_1459,In_990);
nor U519 (N_519,In_257,In_1481);
nand U520 (N_520,N_261,In_987);
and U521 (N_521,In_1270,In_573);
or U522 (N_522,In_584,In_108);
or U523 (N_523,N_70,In_596);
nor U524 (N_524,N_187,N_197);
and U525 (N_525,In_1116,In_1392);
xnor U526 (N_526,In_324,N_207);
and U527 (N_527,In_1397,N_28);
nor U528 (N_528,N_148,In_162);
nor U529 (N_529,In_1131,In_1190);
nand U530 (N_530,In_801,In_1293);
or U531 (N_531,In_795,In_668);
or U532 (N_532,N_152,In_418);
nand U533 (N_533,In_718,In_949);
and U534 (N_534,In_227,In_1150);
and U535 (N_535,In_368,N_320);
nand U536 (N_536,N_1,N_352);
nand U537 (N_537,N_253,In_699);
or U538 (N_538,In_170,N_373);
or U539 (N_539,In_1437,In_829);
and U540 (N_540,N_204,In_866);
or U541 (N_541,In_285,In_102);
nand U542 (N_542,In_1261,N_390);
xor U543 (N_543,In_595,In_961);
or U544 (N_544,In_1364,In_1185);
nand U545 (N_545,In_340,In_260);
xnor U546 (N_546,N_126,In_1105);
nor U547 (N_547,N_328,In_1268);
and U548 (N_548,In_371,In_156);
xnor U549 (N_549,In_316,N_272);
or U550 (N_550,In_694,In_1088);
or U551 (N_551,In_66,N_144);
nor U552 (N_552,In_722,In_380);
or U553 (N_553,In_99,N_248);
or U554 (N_554,In_313,N_259);
and U555 (N_555,In_1370,In_541);
nand U556 (N_556,N_93,In_559);
xor U557 (N_557,In_1342,N_193);
and U558 (N_558,N_130,In_758);
xor U559 (N_559,In_1087,In_181);
xnor U560 (N_560,N_68,In_1004);
and U561 (N_561,In_894,N_334);
nor U562 (N_562,In_1165,In_157);
or U563 (N_563,N_113,In_119);
nand U564 (N_564,N_356,N_236);
nor U565 (N_565,In_545,In_494);
nand U566 (N_566,N_292,In_1238);
nand U567 (N_567,In_616,N_37);
or U568 (N_568,In_492,In_1361);
and U569 (N_569,In_937,N_45);
or U570 (N_570,In_234,N_132);
nand U571 (N_571,In_556,N_103);
or U572 (N_572,N_398,N_239);
nor U573 (N_573,In_577,N_357);
and U574 (N_574,In_377,In_1136);
nand U575 (N_575,In_982,In_322);
and U576 (N_576,In_912,In_441);
or U577 (N_577,In_1236,In_1166);
nor U578 (N_578,In_1441,In_955);
and U579 (N_579,In_461,N_237);
nand U580 (N_580,In_645,In_98);
nor U581 (N_581,N_294,N_83);
xor U582 (N_582,N_392,In_719);
nor U583 (N_583,In_1095,In_3);
and U584 (N_584,N_179,In_1029);
and U585 (N_585,In_1180,In_85);
or U586 (N_586,In_1367,In_918);
xor U587 (N_587,In_238,In_192);
and U588 (N_588,In_678,In_432);
nor U589 (N_589,In_838,N_335);
or U590 (N_590,N_129,In_258);
or U591 (N_591,In_602,N_256);
xnor U592 (N_592,In_1096,In_823);
or U593 (N_593,N_219,In_568);
nor U594 (N_594,In_228,N_184);
and U595 (N_595,N_210,In_771);
or U596 (N_596,In_1324,In_463);
or U597 (N_597,In_1138,In_224);
or U598 (N_598,In_1149,In_1068);
nor U599 (N_599,In_347,N_264);
nand U600 (N_600,N_426,In_55);
and U601 (N_601,N_276,N_251);
nand U602 (N_602,In_1061,In_1162);
nor U603 (N_603,N_342,N_321);
or U604 (N_604,N_411,N_388);
xnor U605 (N_605,N_111,In_751);
or U606 (N_606,In_92,In_390);
xnor U607 (N_607,In_1302,N_490);
nor U608 (N_608,In_148,In_1349);
nor U609 (N_609,N_455,In_1209);
xnor U610 (N_610,N_599,In_911);
and U611 (N_611,In_141,N_548);
and U612 (N_612,In_1273,In_696);
nand U613 (N_613,N_587,In_134);
nor U614 (N_614,In_1288,In_232);
nand U615 (N_615,N_465,In_931);
and U616 (N_616,N_561,In_1212);
or U617 (N_617,In_539,In_808);
or U618 (N_618,N_445,In_1143);
nand U619 (N_619,In_1492,In_817);
or U620 (N_620,In_426,N_568);
xnor U621 (N_621,N_370,N_397);
nor U622 (N_622,In_1347,In_748);
nor U623 (N_623,N_362,In_200);
and U624 (N_624,N_505,N_175);
nand U625 (N_625,In_546,N_150);
xnor U626 (N_626,N_407,In_859);
nor U627 (N_627,In_880,N_271);
xor U628 (N_628,N_151,In_1199);
and U629 (N_629,N_360,In_971);
nand U630 (N_630,N_580,In_1419);
or U631 (N_631,In_800,In_180);
nand U632 (N_632,In_709,N_442);
xnor U633 (N_633,In_905,In_917);
and U634 (N_634,In_1426,N_495);
or U635 (N_635,In_217,In_88);
nor U636 (N_636,N_470,In_431);
xor U637 (N_637,In_625,N_476);
nand U638 (N_638,In_196,N_387);
or U639 (N_639,In_1432,N_280);
nand U640 (N_640,In_948,In_830);
nor U641 (N_641,N_347,In_737);
and U642 (N_642,In_887,In_1477);
nand U643 (N_643,N_209,N_385);
or U644 (N_644,In_57,In_1294);
and U645 (N_645,N_9,N_242);
nand U646 (N_646,N_247,N_486);
or U647 (N_647,N_297,In_449);
nand U648 (N_648,N_422,In_138);
nand U649 (N_649,In_723,N_453);
or U650 (N_650,N_498,N_208);
or U651 (N_651,N_424,In_1006);
nand U652 (N_652,In_1412,In_649);
nand U653 (N_653,In_104,In_42);
and U654 (N_654,N_439,N_597);
nand U655 (N_655,In_187,In_741);
and U656 (N_656,In_457,In_1008);
or U657 (N_657,N_268,In_1193);
nor U658 (N_658,In_582,N_598);
nand U659 (N_659,N_124,In_498);
or U660 (N_660,In_154,N_217);
or U661 (N_661,N_199,In_619);
nand U662 (N_662,In_607,In_96);
nor U663 (N_663,N_47,In_1493);
nand U664 (N_664,N_585,In_37);
nor U665 (N_665,In_330,N_274);
and U666 (N_666,In_1436,N_474);
or U667 (N_667,N_365,N_403);
xor U668 (N_668,N_427,In_1100);
or U669 (N_669,In_826,N_577);
xnor U670 (N_670,N_444,N_170);
nand U671 (N_671,In_792,N_527);
and U672 (N_672,N_501,In_405);
nor U673 (N_673,N_562,In_140);
and U674 (N_674,In_510,In_1478);
and U675 (N_675,In_1128,In_1250);
nand U676 (N_676,N_393,In_1020);
nand U677 (N_677,In_46,N_313);
and U678 (N_678,In_803,In_1290);
xnor U679 (N_679,N_24,In_185);
and U680 (N_680,In_225,N_378);
and U681 (N_681,N_213,N_338);
nand U682 (N_682,In_580,In_739);
or U683 (N_683,In_588,In_623);
nor U684 (N_684,N_510,In_647);
xnor U685 (N_685,N_579,N_105);
or U686 (N_686,N_343,N_183);
or U687 (N_687,In_389,N_372);
and U688 (N_688,N_123,N_405);
nor U689 (N_689,N_524,In_560);
nand U690 (N_690,N_252,In_1075);
xnor U691 (N_691,In_270,In_1197);
and U692 (N_692,N_504,In_1021);
nor U693 (N_693,In_209,N_169);
xnor U694 (N_694,In_1313,N_58);
xor U695 (N_695,In_1470,N_288);
and U696 (N_696,In_381,N_250);
nand U697 (N_697,N_331,N_552);
nand U698 (N_698,In_62,In_1125);
and U699 (N_699,In_252,In_862);
nor U700 (N_700,In_28,In_1146);
and U701 (N_701,In_1129,N_534);
nand U702 (N_702,N_2,In_300);
and U703 (N_703,N_399,N_433);
nor U704 (N_704,N_122,N_273);
nor U705 (N_705,In_1040,N_588);
nand U706 (N_706,In_532,In_1233);
nand U707 (N_707,In_677,In_483);
and U708 (N_708,N_160,In_1221);
or U709 (N_709,N_266,N_195);
or U710 (N_710,N_463,N_159);
nor U711 (N_711,In_310,N_423);
nor U712 (N_712,N_447,N_435);
nand U713 (N_713,N_540,In_523);
nor U714 (N_714,In_240,In_423);
nor U715 (N_715,In_586,In_378);
nor U716 (N_716,N_15,N_284);
nand U717 (N_717,In_354,In_753);
or U718 (N_718,N_409,In_831);
nor U719 (N_719,N_583,N_211);
nand U720 (N_720,In_840,N_556);
nand U721 (N_721,In_591,In_1052);
or U722 (N_722,In_279,N_90);
xor U723 (N_723,In_1453,In_1353);
nor U724 (N_724,In_1042,N_480);
or U725 (N_725,In_293,In_151);
nor U726 (N_726,N_573,In_440);
or U727 (N_727,In_897,In_806);
and U728 (N_728,N_581,In_1010);
nor U729 (N_729,N_202,In_307);
and U730 (N_730,In_1447,In_484);
nor U731 (N_731,N_258,In_847);
nand U732 (N_732,N_220,N_482);
nor U733 (N_733,N_101,In_884);
nor U734 (N_734,N_589,In_788);
nand U735 (N_735,In_1103,N_511);
nand U736 (N_736,N_547,N_243);
nor U737 (N_737,N_441,In_14);
and U738 (N_738,N_538,In_16);
nor U739 (N_739,N_299,In_1079);
nand U740 (N_740,N_249,N_475);
and U741 (N_741,N_305,N_478);
and U742 (N_742,N_289,N_131);
nor U743 (N_743,In_520,In_1443);
or U744 (N_744,N_153,In_214);
and U745 (N_745,In_1363,N_438);
and U746 (N_746,N_309,In_1031);
and U747 (N_747,In_776,N_521);
and U748 (N_748,In_893,In_72);
nor U749 (N_749,In_860,N_322);
nor U750 (N_750,N_255,N_489);
nand U751 (N_751,In_43,In_366);
or U752 (N_752,In_213,In_435);
nand U753 (N_753,N_531,In_197);
nor U754 (N_754,N_430,N_553);
nand U755 (N_755,N_560,In_657);
and U756 (N_756,N_462,N_229);
nand U757 (N_757,In_773,In_1030);
or U758 (N_758,In_1028,N_359);
nand U759 (N_759,In_1264,In_182);
or U760 (N_760,In_253,N_383);
xor U761 (N_761,In_993,N_223);
or U762 (N_762,In_810,N_225);
or U763 (N_763,N_503,N_582);
nand U764 (N_764,In_797,In_1411);
nand U765 (N_765,N_364,N_563);
or U766 (N_766,N_38,In_437);
nor U767 (N_767,In_500,In_1280);
or U768 (N_768,N_63,N_481);
or U769 (N_769,In_395,N_185);
nor U770 (N_770,N_542,N_354);
nand U771 (N_771,In_813,N_472);
nand U772 (N_772,In_570,N_497);
nor U773 (N_773,N_436,In_828);
and U774 (N_774,In_634,In_326);
and U775 (N_775,In_167,In_179);
and U776 (N_776,N_410,N_245);
nand U777 (N_777,In_306,In_728);
xnor U778 (N_778,In_1158,N_147);
and U779 (N_779,In_485,In_901);
nor U780 (N_780,In_468,N_176);
and U781 (N_781,In_400,N_224);
xnor U782 (N_782,In_97,N_412);
or U783 (N_783,N_443,In_249);
nand U784 (N_784,N_572,In_1111);
nor U785 (N_785,N_558,In_1053);
and U786 (N_786,N_491,N_437);
and U787 (N_787,N_395,In_519);
and U788 (N_788,N_537,N_226);
or U789 (N_789,N_488,In_576);
xor U790 (N_790,In_1346,N_432);
xor U791 (N_791,In_256,In_717);
xnor U792 (N_792,N_222,In_663);
or U793 (N_793,In_30,In_20);
and U794 (N_794,N_72,In_956);
nand U795 (N_795,In_1406,In_250);
xor U796 (N_796,N_519,N_402);
or U797 (N_797,In_137,N_508);
and U798 (N_798,In_161,N_308);
xnor U799 (N_799,In_216,N_286);
nand U800 (N_800,N_278,N_302);
nand U801 (N_801,N_198,In_8);
and U802 (N_802,In_1119,In_1024);
nand U803 (N_803,N_709,In_220);
or U804 (N_804,N_682,N_792);
nor U805 (N_805,N_80,N_600);
or U806 (N_806,In_876,N_693);
nand U807 (N_807,N_690,N_216);
and U808 (N_808,N_593,In_958);
xnor U809 (N_809,N_721,In_325);
nand U810 (N_810,In_58,N_624);
and U811 (N_811,N_546,N_483);
nor U812 (N_812,In_533,In_490);
nand U813 (N_813,N_645,In_850);
nor U814 (N_814,N_787,N_479);
or U815 (N_815,In_1118,In_1120);
or U816 (N_816,N_780,In_1234);
and U817 (N_817,In_352,N_196);
nor U818 (N_818,In_1048,In_528);
nand U819 (N_819,In_1274,In_843);
and U820 (N_820,In_13,In_787);
nand U821 (N_821,In_221,In_1278);
nand U822 (N_822,N_528,In_966);
and U823 (N_823,In_17,N_710);
and U824 (N_824,N_457,N_120);
nor U825 (N_825,In_628,N_69);
nor U826 (N_826,In_159,N_536);
nand U827 (N_827,In_998,In_784);
xor U828 (N_828,N_449,In_989);
nor U829 (N_829,N_326,N_704);
or U830 (N_830,In_502,In_1312);
nand U831 (N_831,In_201,In_1189);
and U832 (N_832,N_425,In_844);
nand U833 (N_833,N_744,N_564);
nand U834 (N_834,In_610,In_600);
nand U835 (N_835,In_716,N_533);
and U836 (N_836,In_1253,N_661);
and U837 (N_837,In_1431,In_44);
xnor U838 (N_838,In_1151,N_114);
and U839 (N_839,N_567,N_520);
or U840 (N_840,N_790,In_93);
and U841 (N_841,N_367,N_452);
and U842 (N_842,In_367,In_308);
nand U843 (N_843,In_1122,N_699);
nor U844 (N_844,In_1202,N_512);
or U845 (N_845,N_269,In_818);
xnor U846 (N_846,N_750,N_675);
nand U847 (N_847,N_685,In_727);
nand U848 (N_848,N_307,In_462);
and U849 (N_849,In_689,In_7);
nand U850 (N_850,In_215,In_372);
or U851 (N_851,N_576,N_161);
or U852 (N_852,In_512,N_230);
and U853 (N_853,N_569,In_1204);
and U854 (N_854,N_724,N_789);
nor U855 (N_855,In_902,In_943);
nand U856 (N_856,N_606,N_733);
and U857 (N_857,N_571,N_44);
nand U858 (N_858,In_345,In_1003);
and U859 (N_859,In_76,N_783);
and U860 (N_860,N_784,N_652);
nor U861 (N_861,N_628,N_42);
or U862 (N_862,N_304,N_471);
nor U863 (N_863,In_755,In_549);
and U864 (N_864,N_543,N_756);
and U865 (N_865,N_118,N_663);
nor U866 (N_866,In_962,N_285);
or U867 (N_867,In_77,N_575);
xor U868 (N_868,In_1043,In_1343);
or U869 (N_869,In_144,N_522);
nor U870 (N_870,N_554,N_695);
nor U871 (N_871,N_296,N_234);
xnor U872 (N_872,N_336,N_762);
nand U873 (N_873,N_523,N_700);
or U874 (N_874,N_125,N_221);
nor U875 (N_875,In_534,N_757);
nor U876 (N_876,In_1243,In_910);
or U877 (N_877,N_760,N_257);
or U878 (N_878,N_643,In_1082);
xor U879 (N_879,N_414,N_260);
or U880 (N_880,N_20,N_346);
and U881 (N_881,In_41,N_487);
and U882 (N_882,N_610,N_772);
xnor U883 (N_883,In_644,N_778);
nand U884 (N_884,In_1474,N_391);
xnor U885 (N_885,In_1391,N_779);
and U886 (N_886,N_404,N_641);
nor U887 (N_887,N_14,In_236);
and U888 (N_888,In_1076,N_680);
or U889 (N_889,In_952,N_656);
and U890 (N_890,N_584,N_232);
nand U891 (N_891,N_716,In_1495);
nor U892 (N_892,In_475,N_782);
nand U893 (N_893,N_57,In_875);
nor U894 (N_894,N_623,N_689);
or U895 (N_895,N_301,N_771);
xor U896 (N_896,N_660,In_1299);
nor U897 (N_897,N_630,N_545);
and U898 (N_898,N_74,N_688);
nand U899 (N_899,N_290,N_674);
nor U900 (N_900,N_687,N_622);
and U901 (N_901,N_625,In_48);
nor U902 (N_902,In_328,In_235);
or U903 (N_903,N_350,N_509);
xor U904 (N_904,N_749,N_434);
or U905 (N_905,In_970,In_873);
xor U906 (N_906,N_244,In_734);
nand U907 (N_907,In_355,N_713);
nor U908 (N_908,N_634,N_603);
or U909 (N_909,In_1306,In_409);
or U910 (N_910,N_539,N_440);
xor U911 (N_911,N_746,N_735);
xnor U912 (N_912,In_188,N_698);
nor U913 (N_913,N_65,N_107);
nor U914 (N_914,In_603,In_155);
nand U915 (N_915,N_752,In_903);
nand U916 (N_916,In_403,N_459);
xnor U917 (N_917,N_420,N_319);
and U918 (N_918,In_704,N_578);
nand U919 (N_919,In_1386,N_448);
or U920 (N_920,In_551,N_332);
or U921 (N_921,N_794,N_644);
nor U922 (N_922,In_353,N_662);
nor U923 (N_923,N_456,N_139);
nand U924 (N_924,N_791,N_312);
nand U925 (N_925,N_381,In_1057);
or U926 (N_926,N_140,N_602);
and U927 (N_927,In_115,In_750);
nand U928 (N_928,N_516,N_76);
nor U929 (N_929,In_163,In_495);
nand U930 (N_930,N_56,In_938);
nand U931 (N_931,In_473,N_667);
nand U932 (N_932,N_658,In_166);
and U933 (N_933,N_703,In_662);
or U934 (N_934,In_1090,In_411);
nor U935 (N_935,N_526,N_513);
or U936 (N_936,In_736,In_1304);
and U937 (N_937,In_23,N_182);
or U938 (N_938,N_706,In_271);
nand U939 (N_939,N_728,In_172);
nor U940 (N_940,N_694,N_596);
xnor U941 (N_941,N_473,N_164);
nor U942 (N_942,In_521,In_346);
and U943 (N_943,N_35,In_777);
or U944 (N_944,In_369,In_24);
and U945 (N_945,N_81,In_1471);
and U946 (N_946,N_765,In_1198);
nand U947 (N_947,In_1372,In_642);
or U948 (N_948,N_574,N_203);
nor U949 (N_949,N_167,N_701);
and U950 (N_950,N_609,In_259);
or U951 (N_951,N_550,In_274);
nor U952 (N_952,N_785,N_267);
nor U953 (N_953,N_638,N_607);
and U954 (N_954,In_765,In_1174);
nor U955 (N_955,In_1217,N_454);
nand U956 (N_956,N_747,N_714);
or U957 (N_957,N_428,N_748);
xor U958 (N_958,In_590,N_759);
nor U959 (N_959,In_883,N_742);
nand U960 (N_960,N_477,N_377);
nor U961 (N_961,In_1476,N_758);
xnor U962 (N_962,N_494,N_493);
nor U963 (N_963,N_570,In_1281);
and U964 (N_964,In_1355,In_1321);
or U965 (N_965,N_529,In_59);
xnor U966 (N_966,In_292,In_1173);
nor U967 (N_967,In_394,In_1032);
nand U968 (N_968,N_786,N_52);
nand U969 (N_969,In_598,N_729);
or U970 (N_970,N_717,N_764);
and U971 (N_971,N_594,In_1065);
nor U972 (N_972,N_743,N_633);
and U973 (N_973,N_190,N_753);
and U974 (N_974,N_632,In_898);
nor U975 (N_975,In_230,In_935);
nor U976 (N_976,In_385,N_557);
or U977 (N_977,N_496,N_18);
nor U978 (N_978,N_775,N_6);
and U979 (N_979,N_348,In_1466);
xnor U980 (N_980,N_615,N_621);
nand U981 (N_981,N_605,In_321);
and U982 (N_982,N_781,N_468);
xor U983 (N_983,N_345,N_629);
nand U984 (N_984,N_726,In_922);
xnor U985 (N_985,In_287,N_601);
or U986 (N_986,N_777,In_593);
or U987 (N_987,In_867,In_864);
nor U988 (N_988,In_1318,N_376);
xor U989 (N_989,N_739,In_1226);
nor U990 (N_990,N_555,N_559);
nand U991 (N_991,N_102,In_84);
nand U992 (N_992,N_755,In_749);
and U993 (N_993,N_636,In_1107);
and U994 (N_994,In_684,N_22);
xor U995 (N_995,N_421,In_146);
nand U996 (N_996,N_604,N_460);
and U997 (N_997,In_845,N_774);
or U998 (N_998,N_408,In_627);
xor U999 (N_999,N_429,N_82);
nand U1000 (N_1000,N_985,N_168);
nand U1001 (N_1001,In_1292,N_892);
nor U1002 (N_1002,N_873,N_989);
nand U1003 (N_1003,N_303,N_673);
or U1004 (N_1004,N_872,In_622);
nand U1005 (N_1005,In_413,N_766);
and U1006 (N_1006,N_982,N_800);
or U1007 (N_1007,N_640,N_958);
nand U1008 (N_1008,In_1442,In_1184);
and U1009 (N_1009,N_974,N_720);
and U1010 (N_1010,N_977,N_847);
or U1011 (N_1011,N_642,N_515);
nand U1012 (N_1012,In_231,N_939);
or U1013 (N_1013,N_723,N_890);
xnor U1014 (N_1014,N_532,N_400);
and U1015 (N_1015,N_215,N_870);
nand U1016 (N_1016,N_788,N_861);
nand U1017 (N_1017,N_937,N_708);
nand U1018 (N_1018,N_863,In_1062);
or U1019 (N_1019,N_590,N_620);
or U1020 (N_1020,N_983,N_869);
or U1021 (N_1021,In_1015,N_616);
nor U1022 (N_1022,In_544,N_653);
nor U1023 (N_1023,In_963,N_371);
nor U1024 (N_1024,N_613,N_833);
or U1025 (N_1025,N_12,N_934);
nand U1026 (N_1026,N_925,N_887);
xor U1027 (N_1027,In_110,N_929);
nand U1028 (N_1028,N_964,N_671);
nand U1029 (N_1029,In_574,N_517);
or U1030 (N_1030,In_245,N_970);
nor U1031 (N_1031,N_876,In_226);
or U1032 (N_1032,N_960,In_688);
and U1033 (N_1033,N_881,N_889);
or U1034 (N_1034,N_592,N_830);
and U1035 (N_1035,N_840,N_740);
and U1036 (N_1036,In_1325,In_29);
xnor U1037 (N_1037,N_824,N_962);
and U1038 (N_1038,In_537,N_79);
nor U1039 (N_1039,N_50,N_806);
nor U1040 (N_1040,N_991,N_821);
and U1041 (N_1041,In_940,N_879);
nand U1042 (N_1042,In_516,N_898);
and U1043 (N_1043,In_1262,N_949);
or U1044 (N_1044,N_874,N_845);
nand U1045 (N_1045,N_727,In_1358);
or U1046 (N_1046,N_842,N_947);
nand U1047 (N_1047,N_891,N_910);
and U1048 (N_1048,N_923,In_288);
nor U1049 (N_1049,N_696,In_921);
nand U1050 (N_1050,N_637,In_1332);
and U1051 (N_1051,In_1254,In_715);
nand U1052 (N_1052,N_922,N_834);
nor U1053 (N_1053,N_295,In_1091);
nor U1054 (N_1054,N_948,N_619);
and U1055 (N_1055,N_231,N_839);
nand U1056 (N_1056,N_627,N_659);
xnor U1057 (N_1057,In_929,N_311);
nand U1058 (N_1058,N_672,N_804);
and U1059 (N_1059,N_849,N_595);
nor U1060 (N_1060,In_283,N_992);
and U1061 (N_1061,In_686,N_871);
nand U1062 (N_1062,N_665,N_763);
nand U1063 (N_1063,N_683,N_904);
and U1064 (N_1064,N_639,N_30);
and U1065 (N_1065,N_805,In_793);
xor U1066 (N_1066,N_648,N_883);
nand U1067 (N_1067,N_882,N_722);
nor U1068 (N_1068,In_726,In_327);
or U1069 (N_1069,In_470,In_933);
nor U1070 (N_1070,N_826,N_767);
nor U1071 (N_1071,N_751,N_707);
xnor U1072 (N_1072,N_669,N_993);
nor U1073 (N_1073,N_850,N_911);
nor U1074 (N_1074,N_626,In_50);
nor U1075 (N_1075,N_384,N_987);
or U1076 (N_1076,N_469,In_874);
nor U1077 (N_1077,N_172,N_227);
and U1078 (N_1078,N_506,In_21);
and U1079 (N_1079,N_380,N_337);
nor U1080 (N_1080,N_810,N_691);
and U1081 (N_1081,N_912,N_507);
nand U1082 (N_1082,N_666,N_358);
xor U1083 (N_1083,N_293,N_935);
nor U1084 (N_1084,N_818,N_566);
nand U1085 (N_1085,N_928,N_933);
or U1086 (N_1086,N_608,N_945);
nand U1087 (N_1087,N_936,N_813);
and U1088 (N_1088,N_451,N_959);
and U1089 (N_1089,N_967,In_611);
and U1090 (N_1090,N_829,N_896);
or U1091 (N_1091,N_544,N_916);
and U1092 (N_1092,N_990,N_884);
or U1093 (N_1093,N_877,N_100);
or U1094 (N_1094,N_893,N_363);
nand U1095 (N_1095,N_998,N_664);
xnor U1096 (N_1096,N_955,N_417);
and U1097 (N_1097,N_858,In_589);
nor U1098 (N_1098,N_951,N_89);
nand U1099 (N_1099,N_801,N_214);
xor U1100 (N_1100,N_995,In_1429);
xor U1101 (N_1101,N_901,N_802);
or U1102 (N_1102,In_1344,N_565);
or U1103 (N_1103,In_1215,In_1012);
nor U1104 (N_1104,N_586,N_737);
nor U1105 (N_1105,N_355,N_799);
nor U1106 (N_1106,N_855,N_927);
xnor U1107 (N_1107,N_484,N_612);
nor U1108 (N_1108,N_899,N_969);
and U1109 (N_1109,N_450,In_857);
nor U1110 (N_1110,N_978,N_809);
nand U1111 (N_1111,N_950,In_496);
xor U1112 (N_1112,In_579,N_732);
or U1113 (N_1113,N_968,N_201);
or U1114 (N_1114,N_238,N_827);
nand U1115 (N_1115,In_648,N_770);
or U1116 (N_1116,N_119,N_902);
nor U1117 (N_1117,N_864,In_444);
xnor U1118 (N_1118,N_678,N_618);
nand U1119 (N_1119,In_237,N_711);
and U1120 (N_1120,N_940,N_635);
nor U1121 (N_1121,N_816,N_915);
and U1122 (N_1122,N_697,N_692);
or U1123 (N_1123,N_681,In_1451);
nor U1124 (N_1124,N_396,N_908);
nand U1125 (N_1125,In_1423,N_228);
and U1126 (N_1126,N_712,N_631);
or U1127 (N_1127,N_878,N_946);
nand U1128 (N_1128,In_479,N_654);
nand U1129 (N_1129,In_1134,In_429);
nor U1130 (N_1130,N_300,N_277);
nor U1131 (N_1131,N_754,In_809);
nor U1132 (N_1132,N_525,N_500);
or U1133 (N_1133,N_614,N_909);
nand U1134 (N_1134,N_999,N_846);
nand U1135 (N_1135,N_880,N_715);
nand U1136 (N_1136,N_21,In_1207);
and U1137 (N_1137,N_535,N_731);
or U1138 (N_1138,N_868,In_1488);
xor U1139 (N_1139,In_448,N_918);
nor U1140 (N_1140,N_458,N_127);
nor U1141 (N_1141,N_943,N_825);
nand U1142 (N_1142,In_384,N_803);
and U1143 (N_1143,N_952,N_924);
xor U1144 (N_1144,N_27,N_281);
nand U1145 (N_1145,In_184,N_431);
nor U1146 (N_1146,N_986,N_920);
xnor U1147 (N_1147,In_936,N_797);
or U1148 (N_1148,N_514,N_812);
and U1149 (N_1149,N_241,N_914);
nor U1150 (N_1150,N_415,N_851);
and U1151 (N_1151,N_838,N_651);
and U1152 (N_1152,N_650,N_832);
and U1153 (N_1153,N_734,In_241);
or U1154 (N_1154,N_3,N_931);
or U1155 (N_1155,In_690,N_796);
and U1156 (N_1156,N_793,N_854);
nor U1157 (N_1157,N_705,N_298);
xor U1158 (N_1158,N_905,N_374);
nand U1159 (N_1159,N_655,N_921);
nor U1160 (N_1160,N_768,N_795);
nor U1161 (N_1161,N_903,N_180);
nand U1162 (N_1162,In_1034,N_853);
nand U1163 (N_1163,N_817,N_894);
or U1164 (N_1164,N_173,N_965);
or U1165 (N_1165,N_867,In_1246);
nor U1166 (N_1166,In_147,N_736);
or U1167 (N_1167,In_1182,N_64);
and U1168 (N_1168,In_807,N_541);
nor U1169 (N_1169,N_233,N_283);
nand U1170 (N_1170,N_492,N_932);
and U1171 (N_1171,N_282,In_942);
nor U1172 (N_1172,N_419,N_984);
nor U1173 (N_1173,N_206,N_837);
and U1174 (N_1174,In_1374,N_62);
and U1175 (N_1175,N_446,N_657);
or U1176 (N_1176,N_988,N_972);
or U1177 (N_1177,N_895,N_59);
and U1178 (N_1178,N_485,N_518);
nor U1179 (N_1179,N_36,N_900);
nand U1180 (N_1180,N_676,In_1457);
nand U1181 (N_1181,N_467,N_48);
xor U1182 (N_1182,N_930,N_773);
nor U1183 (N_1183,N_961,N_549);
nor U1184 (N_1184,N_897,N_54);
or U1185 (N_1185,N_416,N_466);
xnor U1186 (N_1186,N_971,N_702);
or U1187 (N_1187,In_1351,N_499);
nand U1188 (N_1188,N_401,N_875);
or U1189 (N_1189,N_265,N_913);
xor U1190 (N_1190,N_973,N_996);
nor U1191 (N_1191,N_807,In_743);
and U1192 (N_1192,N_502,N_843);
nand U1193 (N_1193,In_1283,N_677);
or U1194 (N_1194,N_32,N_382);
or U1195 (N_1195,In_713,N_649);
and U1196 (N_1196,N_966,N_980);
nand U1197 (N_1197,N_848,N_994);
or U1198 (N_1198,N_647,In_171);
or U1199 (N_1199,In_191,N_718);
nand U1200 (N_1200,N_1146,N_1017);
xor U1201 (N_1201,N_954,N_1178);
nor U1202 (N_1202,N_1187,In_1360);
nand U1203 (N_1203,N_1185,N_963);
nand U1204 (N_1204,N_1053,N_1130);
nand U1205 (N_1205,N_828,N_617);
or U1206 (N_1206,N_1020,N_865);
and U1207 (N_1207,N_953,N_1081);
xor U1208 (N_1208,N_1029,N_1042);
nand U1209 (N_1209,N_1176,N_997);
nor U1210 (N_1210,N_1148,N_1033);
nor U1211 (N_1211,N_1036,N_1127);
nor U1212 (N_1212,N_1090,N_1197);
or U1213 (N_1213,N_1022,N_1140);
and U1214 (N_1214,N_668,N_975);
or U1215 (N_1215,N_1145,N_857);
nand U1216 (N_1216,N_1098,N_1156);
and U1217 (N_1217,N_1094,N_1105);
and U1218 (N_1218,In_1475,N_1121);
nand U1219 (N_1219,N_1171,N_679);
nor U1220 (N_1220,In_571,N_808);
nand U1221 (N_1221,N_1128,N_1091);
nand U1222 (N_1222,N_841,N_1047);
nand U1223 (N_1223,N_375,N_1011);
or U1224 (N_1224,N_1123,N_725);
nand U1225 (N_1225,N_886,N_1037);
or U1226 (N_1226,N_1087,N_1092);
and U1227 (N_1227,N_819,N_1165);
nand U1228 (N_1228,N_1005,In_202);
nor U1229 (N_1229,N_1109,N_1074);
and U1230 (N_1230,N_1158,N_1077);
nor U1231 (N_1231,N_1058,N_1136);
and U1232 (N_1232,N_1153,N_1133);
or U1233 (N_1233,N_730,N_1186);
nor U1234 (N_1234,N_835,N_1023);
nor U1235 (N_1235,N_815,N_831);
or U1236 (N_1236,N_1082,N_1061);
xor U1237 (N_1237,N_852,N_1125);
nor U1238 (N_1238,In_1102,N_1161);
and U1239 (N_1239,N_1034,N_1159);
and U1240 (N_1240,N_1045,N_1041);
nor U1241 (N_1241,N_1184,N_823);
nand U1242 (N_1242,N_1122,N_646);
nand U1243 (N_1243,N_461,N_1038);
or U1244 (N_1244,N_1093,N_1191);
and U1245 (N_1245,N_1151,N_1007);
and U1246 (N_1246,In_90,N_1014);
nand U1247 (N_1247,N_1106,N_1144);
nand U1248 (N_1248,N_1157,N_1063);
or U1249 (N_1249,N_1084,N_1108);
nand U1250 (N_1250,N_957,N_1097);
xor U1251 (N_1251,N_719,N_1095);
and U1252 (N_1252,N_1065,In_1041);
nand U1253 (N_1253,N_591,N_1129);
nand U1254 (N_1254,N_979,N_822);
and U1255 (N_1255,In_1188,N_926);
or U1256 (N_1256,In_1322,N_1175);
xnor U1257 (N_1257,N_1001,N_464);
xor U1258 (N_1258,N_1048,N_530);
or U1259 (N_1259,N_686,N_1018);
nor U1260 (N_1260,N_1126,N_1055);
nand U1261 (N_1261,N_1078,N_1027);
or U1262 (N_1262,N_1154,N_1116);
or U1263 (N_1263,N_1013,N_1069);
nand U1264 (N_1264,N_1177,N_1030);
or U1265 (N_1265,N_611,N_418);
or U1266 (N_1266,N_738,N_1002);
nor U1267 (N_1267,N_1028,N_1166);
nand U1268 (N_1268,In_1387,In_130);
and U1269 (N_1269,N_1138,N_1194);
or U1270 (N_1270,N_885,N_1183);
nand U1271 (N_1271,N_1073,N_1179);
xor U1272 (N_1272,N_941,N_1010);
nor U1273 (N_1273,N_860,In_1405);
nand U1274 (N_1274,N_1110,N_684);
nor U1275 (N_1275,N_1174,N_1025);
and U1276 (N_1276,N_844,N_1060);
nor U1277 (N_1277,N_1003,N_1062);
and U1278 (N_1278,N_205,N_1111);
and U1279 (N_1279,N_820,N_1135);
nand U1280 (N_1280,N_1046,N_981);
and U1281 (N_1281,N_1120,In_842);
and U1282 (N_1282,N_1004,N_1075);
nand U1283 (N_1283,N_1099,N_1088);
nand U1284 (N_1284,N_745,N_1066);
or U1285 (N_1285,N_1152,N_1182);
xnor U1286 (N_1286,N_1190,N_769);
nand U1287 (N_1287,N_1195,N_1180);
nor U1288 (N_1288,N_862,N_1149);
xnor U1289 (N_1289,N_551,N_1124);
xor U1290 (N_1290,N_1119,N_1113);
xor U1291 (N_1291,N_1172,N_1137);
and U1292 (N_1292,N_1167,N_1162);
nand U1293 (N_1293,N_1056,N_1101);
nand U1294 (N_1294,N_761,In_594);
and U1295 (N_1295,N_1089,N_1096);
nand U1296 (N_1296,N_1086,N_1076);
or U1297 (N_1297,N_1131,N_1054);
nor U1298 (N_1298,N_1100,N_1169);
or U1299 (N_1299,N_1170,N_1064);
xor U1300 (N_1300,N_413,N_1142);
nand U1301 (N_1301,N_406,N_1115);
nand U1302 (N_1302,In_150,N_1079);
nor U1303 (N_1303,N_1141,N_1016);
nand U1304 (N_1304,N_17,N_1196);
and U1305 (N_1305,N_1103,N_1164);
nand U1306 (N_1306,N_1163,N_1043);
or U1307 (N_1307,N_1147,N_888);
and U1308 (N_1308,N_942,N_1188);
nor U1309 (N_1309,N_1071,In_422);
or U1310 (N_1310,N_798,N_1080);
and U1311 (N_1311,N_1189,N_1035);
and U1312 (N_1312,N_956,In_555);
and U1313 (N_1313,N_1009,N_1021);
nand U1314 (N_1314,N_1024,N_1031);
xor U1315 (N_1315,N_1112,N_741);
nand U1316 (N_1316,N_856,N_1059);
and U1317 (N_1317,N_1132,N_1192);
xor U1318 (N_1318,N_836,N_1198);
or U1319 (N_1319,N_1160,N_1072);
nor U1320 (N_1320,N_1168,N_1104);
nor U1321 (N_1321,N_1057,N_1012);
nor U1322 (N_1322,In_687,In_692);
nor U1323 (N_1323,N_1068,N_944);
nand U1324 (N_1324,N_1044,N_1050);
and U1325 (N_1325,N_1008,In_1266);
nand U1326 (N_1326,N_1118,N_1000);
nor U1327 (N_1327,N_1134,N_919);
xor U1328 (N_1328,In_261,N_1049);
nand U1329 (N_1329,N_1107,In_1359);
and U1330 (N_1330,N_776,N_859);
or U1331 (N_1331,N_906,N_1199);
and U1332 (N_1332,N_1070,N_1102);
and U1333 (N_1333,N_1026,In_61);
or U1334 (N_1334,N_1083,N_279);
nor U1335 (N_1335,N_1139,N_917);
nor U1336 (N_1336,N_1181,N_907);
nor U1337 (N_1337,N_1085,N_1006);
and U1338 (N_1338,N_1193,N_1117);
and U1339 (N_1339,N_938,N_1067);
or U1340 (N_1340,N_814,N_1040);
and U1341 (N_1341,N_1052,N_811);
or U1342 (N_1342,N_670,N_1032);
or U1343 (N_1343,N_1015,In_891);
nor U1344 (N_1344,N_1143,N_1039);
and U1345 (N_1345,N_866,N_1051);
and U1346 (N_1346,N_1173,N_1150);
nand U1347 (N_1347,N_1019,N_1114);
and U1348 (N_1348,In_109,In_414);
and U1349 (N_1349,N_1155,N_976);
and U1350 (N_1350,N_1199,N_1051);
and U1351 (N_1351,N_1104,N_1163);
nand U1352 (N_1352,In_1266,N_461);
or U1353 (N_1353,N_888,N_1127);
xor U1354 (N_1354,N_1007,N_1119);
or U1355 (N_1355,N_686,N_997);
or U1356 (N_1356,N_906,N_1098);
and U1357 (N_1357,N_1161,N_1036);
nor U1358 (N_1358,N_279,N_1023);
nand U1359 (N_1359,N_530,N_1124);
and U1360 (N_1360,N_730,N_1042);
nand U1361 (N_1361,N_1026,N_1131);
nor U1362 (N_1362,N_1101,N_942);
or U1363 (N_1363,N_1115,N_1176);
nand U1364 (N_1364,N_1025,In_594);
xnor U1365 (N_1365,N_1095,N_1130);
nand U1366 (N_1366,N_1076,N_963);
xnor U1367 (N_1367,N_1011,N_1023);
or U1368 (N_1368,In_692,N_975);
or U1369 (N_1369,N_859,N_418);
nand U1370 (N_1370,N_814,N_1182);
xnor U1371 (N_1371,In_261,In_1387);
nor U1372 (N_1372,N_1079,N_1130);
nand U1373 (N_1373,N_823,In_150);
and U1374 (N_1374,N_953,N_865);
nand U1375 (N_1375,N_1006,N_1069);
and U1376 (N_1376,N_1184,N_406);
nor U1377 (N_1377,In_692,N_1059);
nand U1378 (N_1378,N_1103,N_1171);
nand U1379 (N_1379,N_1178,In_1359);
nand U1380 (N_1380,N_1032,N_1036);
nor U1381 (N_1381,In_414,N_852);
or U1382 (N_1382,N_1153,N_1012);
and U1383 (N_1383,In_891,N_1099);
nor U1384 (N_1384,N_1131,N_1059);
nand U1385 (N_1385,N_1058,N_1102);
nor U1386 (N_1386,N_1055,N_1019);
and U1387 (N_1387,N_1136,N_1180);
xnor U1388 (N_1388,N_591,N_1039);
nand U1389 (N_1389,N_953,N_679);
nand U1390 (N_1390,N_375,N_1000);
or U1391 (N_1391,N_1145,N_617);
nand U1392 (N_1392,N_1091,N_938);
xor U1393 (N_1393,N_1121,N_1020);
nand U1394 (N_1394,N_1027,N_1196);
nor U1395 (N_1395,N_1083,N_815);
xnor U1396 (N_1396,N_1091,N_1139);
nand U1397 (N_1397,N_1175,In_555);
nand U1398 (N_1398,N_1039,N_1188);
nand U1399 (N_1399,N_886,N_1128);
or U1400 (N_1400,N_1235,N_1328);
nor U1401 (N_1401,N_1221,N_1203);
nor U1402 (N_1402,N_1352,N_1378);
nor U1403 (N_1403,N_1375,N_1242);
nor U1404 (N_1404,N_1319,N_1337);
nor U1405 (N_1405,N_1284,N_1302);
xor U1406 (N_1406,N_1315,N_1301);
xor U1407 (N_1407,N_1283,N_1345);
or U1408 (N_1408,N_1344,N_1216);
nand U1409 (N_1409,N_1397,N_1240);
and U1410 (N_1410,N_1322,N_1379);
xnor U1411 (N_1411,N_1311,N_1338);
nor U1412 (N_1412,N_1396,N_1351);
nor U1413 (N_1413,N_1326,N_1376);
and U1414 (N_1414,N_1377,N_1255);
nor U1415 (N_1415,N_1205,N_1395);
and U1416 (N_1416,N_1398,N_1295);
and U1417 (N_1417,N_1236,N_1392);
xor U1418 (N_1418,N_1321,N_1279);
nor U1419 (N_1419,N_1211,N_1366);
and U1420 (N_1420,N_1280,N_1286);
nor U1421 (N_1421,N_1316,N_1308);
and U1422 (N_1422,N_1386,N_1297);
nand U1423 (N_1423,N_1268,N_1380);
xor U1424 (N_1424,N_1265,N_1274);
nand U1425 (N_1425,N_1219,N_1259);
nand U1426 (N_1426,N_1317,N_1218);
nor U1427 (N_1427,N_1273,N_1288);
nor U1428 (N_1428,N_1239,N_1213);
or U1429 (N_1429,N_1243,N_1325);
nor U1430 (N_1430,N_1369,N_1270);
xnor U1431 (N_1431,N_1282,N_1207);
or U1432 (N_1432,N_1346,N_1383);
nor U1433 (N_1433,N_1394,N_1206);
or U1434 (N_1434,N_1313,N_1342);
nand U1435 (N_1435,N_1343,N_1226);
nor U1436 (N_1436,N_1246,N_1312);
nor U1437 (N_1437,N_1237,N_1370);
nor U1438 (N_1438,N_1341,N_1238);
and U1439 (N_1439,N_1385,N_1258);
nand U1440 (N_1440,N_1305,N_1355);
and U1441 (N_1441,N_1388,N_1271);
nor U1442 (N_1442,N_1223,N_1310);
xor U1443 (N_1443,N_1276,N_1228);
nand U1444 (N_1444,N_1290,N_1212);
xor U1445 (N_1445,N_1252,N_1220);
nand U1446 (N_1446,N_1365,N_1340);
or U1447 (N_1447,N_1281,N_1222);
nor U1448 (N_1448,N_1229,N_1289);
nand U1449 (N_1449,N_1300,N_1253);
nand U1450 (N_1450,N_1361,N_1368);
or U1451 (N_1451,N_1278,N_1225);
nand U1452 (N_1452,N_1233,N_1232);
or U1453 (N_1453,N_1353,N_1373);
or U1454 (N_1454,N_1339,N_1248);
nand U1455 (N_1455,N_1323,N_1374);
and U1456 (N_1456,N_1224,N_1269);
or U1457 (N_1457,N_1357,N_1390);
and U1458 (N_1458,N_1318,N_1363);
or U1459 (N_1459,N_1234,N_1382);
or U1460 (N_1460,N_1334,N_1251);
and U1461 (N_1461,N_1356,N_1387);
and U1462 (N_1462,N_1267,N_1299);
nor U1463 (N_1463,N_1329,N_1364);
nor U1464 (N_1464,N_1391,N_1381);
nand U1465 (N_1465,N_1320,N_1389);
and U1466 (N_1466,N_1275,N_1244);
and U1467 (N_1467,N_1359,N_1215);
nor U1468 (N_1468,N_1250,N_1347);
and U1469 (N_1469,N_1247,N_1202);
nor U1470 (N_1470,N_1204,N_1245);
or U1471 (N_1471,N_1264,N_1208);
or U1472 (N_1472,N_1335,N_1263);
nor U1473 (N_1473,N_1324,N_1257);
or U1474 (N_1474,N_1393,N_1330);
and U1475 (N_1475,N_1350,N_1231);
nor U1476 (N_1476,N_1230,N_1303);
and U1477 (N_1477,N_1200,N_1304);
xnor U1478 (N_1478,N_1261,N_1210);
or U1479 (N_1479,N_1292,N_1287);
or U1480 (N_1480,N_1358,N_1266);
or U1481 (N_1481,N_1354,N_1262);
xor U1482 (N_1482,N_1362,N_1254);
nand U1483 (N_1483,N_1296,N_1314);
nor U1484 (N_1484,N_1333,N_1367);
or U1485 (N_1485,N_1349,N_1306);
and U1486 (N_1486,N_1371,N_1214);
nand U1487 (N_1487,N_1307,N_1260);
or U1488 (N_1488,N_1249,N_1256);
and U1489 (N_1489,N_1298,N_1372);
or U1490 (N_1490,N_1293,N_1227);
or U1491 (N_1491,N_1399,N_1201);
or U1492 (N_1492,N_1291,N_1327);
and U1493 (N_1493,N_1336,N_1384);
nand U1494 (N_1494,N_1272,N_1331);
or U1495 (N_1495,N_1309,N_1277);
nor U1496 (N_1496,N_1241,N_1294);
nand U1497 (N_1497,N_1348,N_1285);
nand U1498 (N_1498,N_1332,N_1217);
or U1499 (N_1499,N_1209,N_1360);
or U1500 (N_1500,N_1275,N_1318);
nand U1501 (N_1501,N_1216,N_1205);
and U1502 (N_1502,N_1218,N_1358);
and U1503 (N_1503,N_1319,N_1216);
nand U1504 (N_1504,N_1398,N_1273);
nor U1505 (N_1505,N_1326,N_1330);
and U1506 (N_1506,N_1256,N_1380);
and U1507 (N_1507,N_1291,N_1240);
or U1508 (N_1508,N_1349,N_1223);
and U1509 (N_1509,N_1243,N_1343);
nand U1510 (N_1510,N_1256,N_1231);
nand U1511 (N_1511,N_1206,N_1302);
or U1512 (N_1512,N_1290,N_1343);
or U1513 (N_1513,N_1223,N_1393);
and U1514 (N_1514,N_1320,N_1342);
or U1515 (N_1515,N_1354,N_1307);
nor U1516 (N_1516,N_1256,N_1248);
and U1517 (N_1517,N_1283,N_1341);
or U1518 (N_1518,N_1348,N_1275);
nor U1519 (N_1519,N_1236,N_1263);
and U1520 (N_1520,N_1206,N_1312);
nor U1521 (N_1521,N_1385,N_1294);
and U1522 (N_1522,N_1269,N_1300);
and U1523 (N_1523,N_1363,N_1395);
nor U1524 (N_1524,N_1214,N_1312);
nand U1525 (N_1525,N_1234,N_1377);
or U1526 (N_1526,N_1298,N_1334);
nand U1527 (N_1527,N_1387,N_1264);
xnor U1528 (N_1528,N_1310,N_1266);
xnor U1529 (N_1529,N_1284,N_1220);
nor U1530 (N_1530,N_1382,N_1280);
nor U1531 (N_1531,N_1355,N_1200);
nor U1532 (N_1532,N_1243,N_1290);
and U1533 (N_1533,N_1341,N_1339);
nor U1534 (N_1534,N_1316,N_1368);
or U1535 (N_1535,N_1282,N_1302);
xor U1536 (N_1536,N_1280,N_1315);
xor U1537 (N_1537,N_1293,N_1374);
nand U1538 (N_1538,N_1244,N_1273);
or U1539 (N_1539,N_1327,N_1346);
or U1540 (N_1540,N_1377,N_1302);
or U1541 (N_1541,N_1231,N_1354);
and U1542 (N_1542,N_1224,N_1355);
and U1543 (N_1543,N_1326,N_1231);
nand U1544 (N_1544,N_1323,N_1260);
nand U1545 (N_1545,N_1230,N_1304);
nand U1546 (N_1546,N_1389,N_1388);
xor U1547 (N_1547,N_1328,N_1340);
nor U1548 (N_1548,N_1214,N_1217);
or U1549 (N_1549,N_1382,N_1294);
and U1550 (N_1550,N_1316,N_1251);
nand U1551 (N_1551,N_1253,N_1258);
and U1552 (N_1552,N_1318,N_1269);
and U1553 (N_1553,N_1272,N_1215);
nor U1554 (N_1554,N_1208,N_1256);
nor U1555 (N_1555,N_1273,N_1378);
or U1556 (N_1556,N_1325,N_1307);
nand U1557 (N_1557,N_1368,N_1372);
nor U1558 (N_1558,N_1277,N_1349);
nor U1559 (N_1559,N_1261,N_1392);
nand U1560 (N_1560,N_1394,N_1240);
or U1561 (N_1561,N_1341,N_1263);
xor U1562 (N_1562,N_1277,N_1286);
nor U1563 (N_1563,N_1343,N_1356);
nor U1564 (N_1564,N_1238,N_1396);
or U1565 (N_1565,N_1296,N_1266);
and U1566 (N_1566,N_1223,N_1247);
and U1567 (N_1567,N_1325,N_1245);
nor U1568 (N_1568,N_1368,N_1352);
xnor U1569 (N_1569,N_1255,N_1267);
and U1570 (N_1570,N_1276,N_1306);
nand U1571 (N_1571,N_1299,N_1388);
nor U1572 (N_1572,N_1220,N_1317);
nor U1573 (N_1573,N_1279,N_1219);
nand U1574 (N_1574,N_1342,N_1361);
and U1575 (N_1575,N_1229,N_1366);
nand U1576 (N_1576,N_1290,N_1205);
nand U1577 (N_1577,N_1378,N_1381);
nor U1578 (N_1578,N_1297,N_1378);
nor U1579 (N_1579,N_1399,N_1208);
and U1580 (N_1580,N_1204,N_1353);
xnor U1581 (N_1581,N_1369,N_1291);
or U1582 (N_1582,N_1251,N_1362);
nand U1583 (N_1583,N_1219,N_1204);
or U1584 (N_1584,N_1342,N_1243);
and U1585 (N_1585,N_1316,N_1348);
nand U1586 (N_1586,N_1309,N_1290);
xnor U1587 (N_1587,N_1345,N_1289);
or U1588 (N_1588,N_1210,N_1394);
nor U1589 (N_1589,N_1368,N_1256);
nand U1590 (N_1590,N_1219,N_1345);
xnor U1591 (N_1591,N_1220,N_1316);
or U1592 (N_1592,N_1272,N_1367);
or U1593 (N_1593,N_1375,N_1381);
or U1594 (N_1594,N_1325,N_1377);
nor U1595 (N_1595,N_1268,N_1325);
xor U1596 (N_1596,N_1383,N_1343);
or U1597 (N_1597,N_1306,N_1221);
nor U1598 (N_1598,N_1289,N_1324);
or U1599 (N_1599,N_1284,N_1218);
nor U1600 (N_1600,N_1454,N_1431);
nand U1601 (N_1601,N_1490,N_1404);
nor U1602 (N_1602,N_1553,N_1419);
nor U1603 (N_1603,N_1522,N_1421);
nand U1604 (N_1604,N_1541,N_1466);
nor U1605 (N_1605,N_1572,N_1573);
or U1606 (N_1606,N_1525,N_1401);
xnor U1607 (N_1607,N_1430,N_1532);
nand U1608 (N_1608,N_1512,N_1455);
nand U1609 (N_1609,N_1496,N_1498);
nand U1610 (N_1610,N_1445,N_1465);
nand U1611 (N_1611,N_1491,N_1479);
or U1612 (N_1612,N_1446,N_1439);
nand U1613 (N_1613,N_1552,N_1508);
nand U1614 (N_1614,N_1503,N_1457);
nor U1615 (N_1615,N_1570,N_1470);
and U1616 (N_1616,N_1580,N_1523);
nand U1617 (N_1617,N_1427,N_1544);
nor U1618 (N_1618,N_1540,N_1405);
and U1619 (N_1619,N_1548,N_1453);
nor U1620 (N_1620,N_1526,N_1534);
or U1621 (N_1621,N_1560,N_1551);
and U1622 (N_1622,N_1527,N_1422);
nand U1623 (N_1623,N_1538,N_1474);
or U1624 (N_1624,N_1585,N_1590);
nor U1625 (N_1625,N_1594,N_1500);
nand U1626 (N_1626,N_1418,N_1413);
xnor U1627 (N_1627,N_1480,N_1437);
nor U1628 (N_1628,N_1574,N_1407);
nand U1629 (N_1629,N_1459,N_1499);
nand U1630 (N_1630,N_1433,N_1494);
and U1631 (N_1631,N_1575,N_1415);
xor U1632 (N_1632,N_1542,N_1406);
nand U1633 (N_1633,N_1448,N_1428);
and U1634 (N_1634,N_1475,N_1586);
nor U1635 (N_1635,N_1472,N_1592);
or U1636 (N_1636,N_1516,N_1481);
nand U1637 (N_1637,N_1414,N_1408);
and U1638 (N_1638,N_1520,N_1409);
and U1639 (N_1639,N_1537,N_1462);
and U1640 (N_1640,N_1441,N_1420);
nor U1641 (N_1641,N_1577,N_1506);
nand U1642 (N_1642,N_1461,N_1473);
nand U1643 (N_1643,N_1443,N_1576);
nand U1644 (N_1644,N_1442,N_1438);
or U1645 (N_1645,N_1567,N_1578);
or U1646 (N_1646,N_1514,N_1564);
xnor U1647 (N_1647,N_1529,N_1556);
or U1648 (N_1648,N_1495,N_1424);
xnor U1649 (N_1649,N_1460,N_1486);
and U1650 (N_1650,N_1566,N_1571);
nand U1651 (N_1651,N_1444,N_1450);
or U1652 (N_1652,N_1563,N_1435);
or U1653 (N_1653,N_1426,N_1477);
nor U1654 (N_1654,N_1565,N_1579);
nand U1655 (N_1655,N_1416,N_1533);
or U1656 (N_1656,N_1555,N_1513);
or U1657 (N_1657,N_1501,N_1488);
nand U1658 (N_1658,N_1449,N_1561);
xnor U1659 (N_1659,N_1515,N_1589);
xor U1660 (N_1660,N_1509,N_1587);
and U1661 (N_1661,N_1543,N_1596);
nand U1662 (N_1662,N_1584,N_1468);
and U1663 (N_1663,N_1412,N_1507);
nand U1664 (N_1664,N_1536,N_1411);
and U1665 (N_1665,N_1504,N_1463);
nor U1666 (N_1666,N_1482,N_1493);
xor U1667 (N_1667,N_1489,N_1485);
and U1668 (N_1668,N_1484,N_1517);
or U1669 (N_1669,N_1557,N_1510);
and U1670 (N_1670,N_1559,N_1425);
nand U1671 (N_1671,N_1458,N_1569);
nand U1672 (N_1672,N_1434,N_1447);
nand U1673 (N_1673,N_1582,N_1524);
and U1674 (N_1674,N_1598,N_1502);
nor U1675 (N_1675,N_1558,N_1545);
or U1676 (N_1676,N_1546,N_1599);
and U1677 (N_1677,N_1432,N_1471);
nor U1678 (N_1678,N_1593,N_1531);
nand U1679 (N_1679,N_1568,N_1588);
and U1680 (N_1680,N_1451,N_1505);
or U1681 (N_1681,N_1530,N_1469);
or U1682 (N_1682,N_1476,N_1528);
nand U1683 (N_1683,N_1456,N_1429);
or U1684 (N_1684,N_1519,N_1492);
nor U1685 (N_1685,N_1583,N_1402);
and U1686 (N_1686,N_1483,N_1518);
nor U1687 (N_1687,N_1497,N_1597);
and U1688 (N_1688,N_1410,N_1539);
or U1689 (N_1689,N_1440,N_1521);
and U1690 (N_1690,N_1464,N_1562);
or U1691 (N_1691,N_1549,N_1478);
and U1692 (N_1692,N_1547,N_1436);
xnor U1693 (N_1693,N_1487,N_1595);
or U1694 (N_1694,N_1591,N_1423);
or U1695 (N_1695,N_1400,N_1452);
and U1696 (N_1696,N_1467,N_1554);
nor U1697 (N_1697,N_1511,N_1581);
and U1698 (N_1698,N_1535,N_1403);
nand U1699 (N_1699,N_1417,N_1550);
or U1700 (N_1700,N_1420,N_1423);
and U1701 (N_1701,N_1479,N_1459);
nand U1702 (N_1702,N_1482,N_1574);
nor U1703 (N_1703,N_1557,N_1576);
or U1704 (N_1704,N_1550,N_1505);
and U1705 (N_1705,N_1591,N_1493);
or U1706 (N_1706,N_1400,N_1525);
and U1707 (N_1707,N_1455,N_1500);
and U1708 (N_1708,N_1551,N_1469);
and U1709 (N_1709,N_1424,N_1471);
or U1710 (N_1710,N_1554,N_1559);
or U1711 (N_1711,N_1509,N_1554);
or U1712 (N_1712,N_1576,N_1599);
nand U1713 (N_1713,N_1587,N_1415);
or U1714 (N_1714,N_1405,N_1571);
and U1715 (N_1715,N_1565,N_1582);
nand U1716 (N_1716,N_1592,N_1471);
and U1717 (N_1717,N_1564,N_1428);
or U1718 (N_1718,N_1484,N_1469);
or U1719 (N_1719,N_1510,N_1551);
and U1720 (N_1720,N_1408,N_1593);
nor U1721 (N_1721,N_1522,N_1524);
xnor U1722 (N_1722,N_1480,N_1453);
nand U1723 (N_1723,N_1559,N_1433);
xor U1724 (N_1724,N_1547,N_1520);
nor U1725 (N_1725,N_1533,N_1451);
or U1726 (N_1726,N_1549,N_1525);
nor U1727 (N_1727,N_1571,N_1433);
nor U1728 (N_1728,N_1538,N_1522);
xnor U1729 (N_1729,N_1487,N_1532);
and U1730 (N_1730,N_1456,N_1412);
nor U1731 (N_1731,N_1418,N_1460);
xor U1732 (N_1732,N_1516,N_1435);
or U1733 (N_1733,N_1487,N_1439);
nand U1734 (N_1734,N_1539,N_1530);
nand U1735 (N_1735,N_1484,N_1551);
nor U1736 (N_1736,N_1558,N_1502);
nor U1737 (N_1737,N_1596,N_1553);
or U1738 (N_1738,N_1512,N_1514);
or U1739 (N_1739,N_1442,N_1575);
nand U1740 (N_1740,N_1452,N_1434);
xor U1741 (N_1741,N_1518,N_1599);
and U1742 (N_1742,N_1400,N_1553);
xnor U1743 (N_1743,N_1541,N_1548);
nor U1744 (N_1744,N_1548,N_1465);
xor U1745 (N_1745,N_1418,N_1513);
or U1746 (N_1746,N_1423,N_1532);
and U1747 (N_1747,N_1585,N_1577);
nand U1748 (N_1748,N_1476,N_1403);
xor U1749 (N_1749,N_1475,N_1472);
nand U1750 (N_1750,N_1469,N_1488);
or U1751 (N_1751,N_1517,N_1570);
or U1752 (N_1752,N_1513,N_1466);
and U1753 (N_1753,N_1470,N_1511);
or U1754 (N_1754,N_1545,N_1546);
or U1755 (N_1755,N_1506,N_1578);
nor U1756 (N_1756,N_1512,N_1409);
xor U1757 (N_1757,N_1520,N_1490);
nand U1758 (N_1758,N_1465,N_1530);
nand U1759 (N_1759,N_1421,N_1400);
nor U1760 (N_1760,N_1507,N_1462);
or U1761 (N_1761,N_1523,N_1558);
and U1762 (N_1762,N_1551,N_1544);
nand U1763 (N_1763,N_1493,N_1478);
nand U1764 (N_1764,N_1440,N_1461);
or U1765 (N_1765,N_1559,N_1484);
or U1766 (N_1766,N_1592,N_1413);
nand U1767 (N_1767,N_1531,N_1447);
or U1768 (N_1768,N_1540,N_1447);
nor U1769 (N_1769,N_1456,N_1490);
nand U1770 (N_1770,N_1500,N_1424);
nand U1771 (N_1771,N_1572,N_1514);
nor U1772 (N_1772,N_1461,N_1404);
nand U1773 (N_1773,N_1511,N_1404);
nor U1774 (N_1774,N_1559,N_1521);
nand U1775 (N_1775,N_1536,N_1584);
and U1776 (N_1776,N_1443,N_1445);
and U1777 (N_1777,N_1441,N_1504);
nor U1778 (N_1778,N_1485,N_1511);
nor U1779 (N_1779,N_1599,N_1584);
and U1780 (N_1780,N_1460,N_1473);
xor U1781 (N_1781,N_1563,N_1416);
or U1782 (N_1782,N_1434,N_1471);
nor U1783 (N_1783,N_1490,N_1473);
xnor U1784 (N_1784,N_1566,N_1469);
and U1785 (N_1785,N_1506,N_1415);
or U1786 (N_1786,N_1539,N_1435);
or U1787 (N_1787,N_1435,N_1417);
or U1788 (N_1788,N_1569,N_1501);
nand U1789 (N_1789,N_1426,N_1596);
and U1790 (N_1790,N_1489,N_1568);
and U1791 (N_1791,N_1588,N_1433);
and U1792 (N_1792,N_1400,N_1554);
nand U1793 (N_1793,N_1413,N_1532);
nand U1794 (N_1794,N_1555,N_1580);
and U1795 (N_1795,N_1507,N_1463);
nand U1796 (N_1796,N_1401,N_1534);
nor U1797 (N_1797,N_1439,N_1526);
nor U1798 (N_1798,N_1482,N_1587);
or U1799 (N_1799,N_1440,N_1566);
or U1800 (N_1800,N_1747,N_1778);
nor U1801 (N_1801,N_1714,N_1679);
or U1802 (N_1802,N_1697,N_1774);
nor U1803 (N_1803,N_1782,N_1637);
nor U1804 (N_1804,N_1797,N_1662);
or U1805 (N_1805,N_1645,N_1722);
xor U1806 (N_1806,N_1798,N_1687);
nor U1807 (N_1807,N_1773,N_1675);
xor U1808 (N_1808,N_1762,N_1733);
nor U1809 (N_1809,N_1757,N_1735);
nand U1810 (N_1810,N_1677,N_1781);
nand U1811 (N_1811,N_1784,N_1609);
or U1812 (N_1812,N_1776,N_1655);
nand U1813 (N_1813,N_1788,N_1616);
or U1814 (N_1814,N_1700,N_1622);
and U1815 (N_1815,N_1689,N_1644);
xnor U1816 (N_1816,N_1728,N_1795);
or U1817 (N_1817,N_1604,N_1754);
nand U1818 (N_1818,N_1794,N_1750);
or U1819 (N_1819,N_1760,N_1702);
and U1820 (N_1820,N_1764,N_1739);
xnor U1821 (N_1821,N_1650,N_1652);
nor U1822 (N_1822,N_1727,N_1752);
and U1823 (N_1823,N_1721,N_1659);
nand U1824 (N_1824,N_1611,N_1674);
xnor U1825 (N_1825,N_1631,N_1744);
nand U1826 (N_1826,N_1725,N_1691);
or U1827 (N_1827,N_1625,N_1698);
nor U1828 (N_1828,N_1623,N_1668);
or U1829 (N_1829,N_1640,N_1686);
nand U1830 (N_1830,N_1633,N_1607);
nand U1831 (N_1831,N_1756,N_1682);
nand U1832 (N_1832,N_1734,N_1710);
and U1833 (N_1833,N_1738,N_1613);
xnor U1834 (N_1834,N_1638,N_1615);
or U1835 (N_1835,N_1643,N_1660);
and U1836 (N_1836,N_1799,N_1743);
xnor U1837 (N_1837,N_1731,N_1793);
xor U1838 (N_1838,N_1765,N_1614);
and U1839 (N_1839,N_1680,N_1654);
and U1840 (N_1840,N_1639,N_1786);
or U1841 (N_1841,N_1651,N_1769);
and U1842 (N_1842,N_1635,N_1707);
nor U1843 (N_1843,N_1658,N_1605);
nor U1844 (N_1844,N_1663,N_1737);
nor U1845 (N_1845,N_1718,N_1758);
and U1846 (N_1846,N_1766,N_1742);
nor U1847 (N_1847,N_1661,N_1626);
nor U1848 (N_1848,N_1619,N_1717);
or U1849 (N_1849,N_1796,N_1775);
and U1850 (N_1850,N_1693,N_1724);
or U1851 (N_1851,N_1712,N_1627);
or U1852 (N_1852,N_1632,N_1779);
or U1853 (N_1853,N_1730,N_1706);
or U1854 (N_1854,N_1719,N_1624);
nand U1855 (N_1855,N_1629,N_1608);
nor U1856 (N_1856,N_1656,N_1705);
xor U1857 (N_1857,N_1620,N_1780);
nor U1858 (N_1858,N_1792,N_1701);
nand U1859 (N_1859,N_1732,N_1768);
nor U1860 (N_1860,N_1617,N_1603);
nand U1861 (N_1861,N_1711,N_1759);
or U1862 (N_1862,N_1669,N_1751);
nand U1863 (N_1863,N_1720,N_1741);
or U1864 (N_1864,N_1696,N_1783);
nor U1865 (N_1865,N_1777,N_1692);
or U1866 (N_1866,N_1745,N_1646);
nand U1867 (N_1867,N_1785,N_1670);
and U1868 (N_1868,N_1673,N_1685);
nand U1869 (N_1869,N_1746,N_1606);
nor U1870 (N_1870,N_1709,N_1618);
nor U1871 (N_1871,N_1749,N_1729);
nand U1872 (N_1872,N_1704,N_1601);
nand U1873 (N_1873,N_1755,N_1664);
nor U1874 (N_1874,N_1649,N_1703);
or U1875 (N_1875,N_1683,N_1684);
nand U1876 (N_1876,N_1716,N_1678);
and U1877 (N_1877,N_1708,N_1713);
nor U1878 (N_1878,N_1642,N_1695);
xnor U1879 (N_1879,N_1748,N_1761);
and U1880 (N_1880,N_1634,N_1636);
xor U1881 (N_1881,N_1647,N_1740);
and U1882 (N_1882,N_1694,N_1676);
or U1883 (N_1883,N_1681,N_1699);
xnor U1884 (N_1884,N_1736,N_1610);
nand U1885 (N_1885,N_1630,N_1648);
nor U1886 (N_1886,N_1628,N_1688);
and U1887 (N_1887,N_1787,N_1791);
and U1888 (N_1888,N_1690,N_1715);
nand U1889 (N_1889,N_1600,N_1771);
nand U1890 (N_1890,N_1621,N_1653);
nand U1891 (N_1891,N_1657,N_1602);
and U1892 (N_1892,N_1672,N_1763);
and U1893 (N_1893,N_1612,N_1723);
nand U1894 (N_1894,N_1641,N_1770);
nand U1895 (N_1895,N_1772,N_1726);
nor U1896 (N_1896,N_1665,N_1789);
nor U1897 (N_1897,N_1790,N_1767);
nor U1898 (N_1898,N_1667,N_1753);
xnor U1899 (N_1899,N_1671,N_1666);
or U1900 (N_1900,N_1764,N_1636);
nand U1901 (N_1901,N_1640,N_1631);
nor U1902 (N_1902,N_1627,N_1679);
and U1903 (N_1903,N_1616,N_1695);
and U1904 (N_1904,N_1668,N_1646);
or U1905 (N_1905,N_1647,N_1633);
nor U1906 (N_1906,N_1684,N_1647);
xnor U1907 (N_1907,N_1794,N_1641);
nand U1908 (N_1908,N_1684,N_1635);
nor U1909 (N_1909,N_1637,N_1764);
nand U1910 (N_1910,N_1651,N_1670);
or U1911 (N_1911,N_1614,N_1675);
nor U1912 (N_1912,N_1603,N_1652);
or U1913 (N_1913,N_1779,N_1680);
and U1914 (N_1914,N_1767,N_1694);
nor U1915 (N_1915,N_1713,N_1687);
nand U1916 (N_1916,N_1625,N_1687);
or U1917 (N_1917,N_1623,N_1796);
xor U1918 (N_1918,N_1715,N_1787);
and U1919 (N_1919,N_1739,N_1711);
or U1920 (N_1920,N_1713,N_1606);
nand U1921 (N_1921,N_1764,N_1772);
nor U1922 (N_1922,N_1607,N_1638);
or U1923 (N_1923,N_1665,N_1617);
xnor U1924 (N_1924,N_1793,N_1695);
nor U1925 (N_1925,N_1611,N_1789);
and U1926 (N_1926,N_1700,N_1768);
or U1927 (N_1927,N_1779,N_1698);
nor U1928 (N_1928,N_1638,N_1660);
or U1929 (N_1929,N_1789,N_1658);
or U1930 (N_1930,N_1623,N_1661);
xnor U1931 (N_1931,N_1744,N_1614);
nand U1932 (N_1932,N_1759,N_1768);
nor U1933 (N_1933,N_1776,N_1724);
xor U1934 (N_1934,N_1743,N_1673);
nor U1935 (N_1935,N_1799,N_1605);
nor U1936 (N_1936,N_1655,N_1731);
nor U1937 (N_1937,N_1704,N_1639);
nor U1938 (N_1938,N_1702,N_1788);
nand U1939 (N_1939,N_1716,N_1641);
nor U1940 (N_1940,N_1735,N_1791);
nor U1941 (N_1941,N_1766,N_1705);
nand U1942 (N_1942,N_1724,N_1631);
xnor U1943 (N_1943,N_1725,N_1622);
nand U1944 (N_1944,N_1665,N_1720);
and U1945 (N_1945,N_1699,N_1755);
or U1946 (N_1946,N_1664,N_1631);
and U1947 (N_1947,N_1706,N_1655);
xnor U1948 (N_1948,N_1726,N_1630);
nor U1949 (N_1949,N_1611,N_1629);
nor U1950 (N_1950,N_1673,N_1723);
nor U1951 (N_1951,N_1672,N_1740);
or U1952 (N_1952,N_1677,N_1630);
or U1953 (N_1953,N_1675,N_1734);
nand U1954 (N_1954,N_1743,N_1663);
nand U1955 (N_1955,N_1704,N_1663);
and U1956 (N_1956,N_1735,N_1654);
and U1957 (N_1957,N_1672,N_1617);
and U1958 (N_1958,N_1679,N_1712);
or U1959 (N_1959,N_1742,N_1782);
and U1960 (N_1960,N_1629,N_1693);
and U1961 (N_1961,N_1754,N_1653);
or U1962 (N_1962,N_1764,N_1715);
nor U1963 (N_1963,N_1722,N_1795);
nor U1964 (N_1964,N_1613,N_1697);
nand U1965 (N_1965,N_1661,N_1698);
or U1966 (N_1966,N_1622,N_1751);
nand U1967 (N_1967,N_1712,N_1647);
nand U1968 (N_1968,N_1753,N_1709);
and U1969 (N_1969,N_1655,N_1663);
and U1970 (N_1970,N_1799,N_1771);
or U1971 (N_1971,N_1704,N_1658);
nor U1972 (N_1972,N_1648,N_1720);
nor U1973 (N_1973,N_1644,N_1608);
and U1974 (N_1974,N_1685,N_1618);
or U1975 (N_1975,N_1641,N_1713);
nor U1976 (N_1976,N_1735,N_1687);
nor U1977 (N_1977,N_1760,N_1688);
and U1978 (N_1978,N_1658,N_1755);
xnor U1979 (N_1979,N_1699,N_1676);
nor U1980 (N_1980,N_1689,N_1638);
nor U1981 (N_1981,N_1740,N_1721);
nand U1982 (N_1982,N_1623,N_1721);
nand U1983 (N_1983,N_1728,N_1770);
and U1984 (N_1984,N_1655,N_1642);
nand U1985 (N_1985,N_1741,N_1615);
and U1986 (N_1986,N_1652,N_1678);
or U1987 (N_1987,N_1730,N_1625);
and U1988 (N_1988,N_1659,N_1747);
or U1989 (N_1989,N_1796,N_1753);
or U1990 (N_1990,N_1600,N_1784);
nor U1991 (N_1991,N_1705,N_1686);
nand U1992 (N_1992,N_1710,N_1754);
nand U1993 (N_1993,N_1678,N_1618);
nand U1994 (N_1994,N_1797,N_1785);
nor U1995 (N_1995,N_1776,N_1714);
or U1996 (N_1996,N_1632,N_1643);
and U1997 (N_1997,N_1738,N_1617);
nand U1998 (N_1998,N_1751,N_1723);
or U1999 (N_1999,N_1643,N_1747);
or U2000 (N_2000,N_1839,N_1824);
nand U2001 (N_2001,N_1966,N_1964);
and U2002 (N_2002,N_1812,N_1977);
nand U2003 (N_2003,N_1979,N_1858);
nor U2004 (N_2004,N_1999,N_1837);
nor U2005 (N_2005,N_1841,N_1892);
and U2006 (N_2006,N_1913,N_1942);
or U2007 (N_2007,N_1933,N_1894);
and U2008 (N_2008,N_1873,N_1822);
nand U2009 (N_2009,N_1806,N_1866);
nor U2010 (N_2010,N_1811,N_1915);
or U2011 (N_2011,N_1850,N_1876);
nand U2012 (N_2012,N_1831,N_1997);
or U2013 (N_2013,N_1846,N_1947);
or U2014 (N_2014,N_1987,N_1991);
nand U2015 (N_2015,N_1855,N_1968);
nand U2016 (N_2016,N_1814,N_1869);
and U2017 (N_2017,N_1899,N_1955);
or U2018 (N_2018,N_1874,N_1861);
and U2019 (N_2019,N_1819,N_1889);
nor U2020 (N_2020,N_1962,N_1921);
nor U2021 (N_2021,N_1941,N_1998);
and U2022 (N_2022,N_1912,N_1937);
xnor U2023 (N_2023,N_1994,N_1835);
or U2024 (N_2024,N_1978,N_1909);
xor U2025 (N_2025,N_1951,N_1905);
nor U2026 (N_2026,N_1878,N_1830);
nand U2027 (N_2027,N_1950,N_1843);
or U2028 (N_2028,N_1816,N_1976);
or U2029 (N_2029,N_1957,N_1829);
nand U2030 (N_2030,N_1840,N_1872);
or U2031 (N_2031,N_1813,N_1992);
nor U2032 (N_2032,N_1986,N_1810);
nand U2033 (N_2033,N_1936,N_1895);
xor U2034 (N_2034,N_1823,N_1862);
and U2035 (N_2035,N_1988,N_1938);
or U2036 (N_2036,N_1901,N_1900);
nand U2037 (N_2037,N_1802,N_1917);
nor U2038 (N_2038,N_1845,N_1943);
or U2039 (N_2039,N_1803,N_1825);
or U2040 (N_2040,N_1940,N_1908);
xnor U2041 (N_2041,N_1863,N_1919);
and U2042 (N_2042,N_1805,N_1877);
or U2043 (N_2043,N_1982,N_1849);
nor U2044 (N_2044,N_1907,N_1881);
nand U2045 (N_2045,N_1885,N_1800);
and U2046 (N_2046,N_1844,N_1944);
and U2047 (N_2047,N_1882,N_1854);
nand U2048 (N_2048,N_1821,N_1867);
nand U2049 (N_2049,N_1870,N_1817);
or U2050 (N_2050,N_1923,N_1856);
nor U2051 (N_2051,N_1836,N_1827);
or U2052 (N_2052,N_1970,N_1945);
or U2053 (N_2053,N_1879,N_1931);
and U2054 (N_2054,N_1851,N_1838);
nand U2055 (N_2055,N_1801,N_1902);
nor U2056 (N_2056,N_1868,N_1865);
nand U2057 (N_2057,N_1897,N_1833);
and U2058 (N_2058,N_1864,N_1848);
xor U2059 (N_2059,N_1896,N_1990);
and U2060 (N_2060,N_1949,N_1969);
xor U2061 (N_2061,N_1916,N_1929);
and U2062 (N_2062,N_1927,N_1961);
or U2063 (N_2063,N_1928,N_1884);
nor U2064 (N_2064,N_1954,N_1948);
and U2065 (N_2065,N_1807,N_1963);
or U2066 (N_2066,N_1925,N_1932);
nor U2067 (N_2067,N_1852,N_1993);
and U2068 (N_2068,N_1939,N_1967);
and U2069 (N_2069,N_1920,N_1906);
or U2070 (N_2070,N_1808,N_1888);
nand U2071 (N_2071,N_1815,N_1893);
or U2072 (N_2072,N_1887,N_1981);
and U2073 (N_2073,N_1886,N_1975);
nand U2074 (N_2074,N_1818,N_1985);
or U2075 (N_2075,N_1904,N_1804);
or U2076 (N_2076,N_1832,N_1898);
nor U2077 (N_2077,N_1847,N_1930);
nand U2078 (N_2078,N_1974,N_1809);
or U2079 (N_2079,N_1958,N_1859);
and U2080 (N_2080,N_1973,N_1959);
xor U2081 (N_2081,N_1875,N_1971);
nor U2082 (N_2082,N_1860,N_1989);
or U2083 (N_2083,N_1890,N_1926);
xor U2084 (N_2084,N_1820,N_1934);
and U2085 (N_2085,N_1891,N_1826);
nand U2086 (N_2086,N_1980,N_1903);
nor U2087 (N_2087,N_1983,N_1918);
nand U2088 (N_2088,N_1952,N_1922);
or U2089 (N_2089,N_1828,N_1996);
or U2090 (N_2090,N_1960,N_1995);
or U2091 (N_2091,N_1956,N_1871);
xor U2092 (N_2092,N_1946,N_1883);
nand U2093 (N_2093,N_1972,N_1857);
or U2094 (N_2094,N_1953,N_1965);
or U2095 (N_2095,N_1911,N_1910);
nor U2096 (N_2096,N_1935,N_1984);
xnor U2097 (N_2097,N_1880,N_1842);
nor U2098 (N_2098,N_1853,N_1834);
and U2099 (N_2099,N_1914,N_1924);
nor U2100 (N_2100,N_1898,N_1979);
nor U2101 (N_2101,N_1970,N_1914);
and U2102 (N_2102,N_1893,N_1801);
nand U2103 (N_2103,N_1874,N_1887);
nand U2104 (N_2104,N_1921,N_1843);
nand U2105 (N_2105,N_1961,N_1949);
or U2106 (N_2106,N_1971,N_1948);
nand U2107 (N_2107,N_1846,N_1970);
and U2108 (N_2108,N_1978,N_1809);
nor U2109 (N_2109,N_1994,N_1818);
or U2110 (N_2110,N_1842,N_1986);
or U2111 (N_2111,N_1918,N_1962);
and U2112 (N_2112,N_1814,N_1984);
nor U2113 (N_2113,N_1854,N_1938);
nand U2114 (N_2114,N_1926,N_1891);
and U2115 (N_2115,N_1882,N_1956);
and U2116 (N_2116,N_1941,N_1971);
nor U2117 (N_2117,N_1958,N_1957);
and U2118 (N_2118,N_1936,N_1977);
and U2119 (N_2119,N_1983,N_1998);
and U2120 (N_2120,N_1818,N_1858);
and U2121 (N_2121,N_1840,N_1882);
nand U2122 (N_2122,N_1909,N_1988);
nand U2123 (N_2123,N_1990,N_1951);
nor U2124 (N_2124,N_1887,N_1939);
xor U2125 (N_2125,N_1819,N_1858);
or U2126 (N_2126,N_1849,N_1854);
nor U2127 (N_2127,N_1801,N_1809);
and U2128 (N_2128,N_1927,N_1832);
nand U2129 (N_2129,N_1913,N_1919);
nand U2130 (N_2130,N_1931,N_1910);
nand U2131 (N_2131,N_1982,N_1871);
xor U2132 (N_2132,N_1885,N_1895);
xor U2133 (N_2133,N_1984,N_1823);
or U2134 (N_2134,N_1826,N_1877);
and U2135 (N_2135,N_1910,N_1845);
nand U2136 (N_2136,N_1869,N_1976);
or U2137 (N_2137,N_1955,N_1994);
nand U2138 (N_2138,N_1861,N_1951);
xnor U2139 (N_2139,N_1923,N_1977);
nor U2140 (N_2140,N_1926,N_1860);
or U2141 (N_2141,N_1900,N_1858);
and U2142 (N_2142,N_1907,N_1987);
xor U2143 (N_2143,N_1869,N_1874);
and U2144 (N_2144,N_1939,N_1986);
or U2145 (N_2145,N_1907,N_1802);
and U2146 (N_2146,N_1911,N_1967);
nand U2147 (N_2147,N_1806,N_1957);
nor U2148 (N_2148,N_1889,N_1986);
and U2149 (N_2149,N_1923,N_1887);
nand U2150 (N_2150,N_1860,N_1835);
and U2151 (N_2151,N_1831,N_1880);
and U2152 (N_2152,N_1995,N_1900);
nor U2153 (N_2153,N_1850,N_1973);
nor U2154 (N_2154,N_1905,N_1981);
nand U2155 (N_2155,N_1821,N_1978);
and U2156 (N_2156,N_1818,N_1874);
and U2157 (N_2157,N_1986,N_1993);
nand U2158 (N_2158,N_1991,N_1861);
or U2159 (N_2159,N_1864,N_1820);
or U2160 (N_2160,N_1932,N_1920);
nor U2161 (N_2161,N_1977,N_1876);
or U2162 (N_2162,N_1810,N_1920);
and U2163 (N_2163,N_1833,N_1826);
or U2164 (N_2164,N_1893,N_1846);
xnor U2165 (N_2165,N_1831,N_1811);
or U2166 (N_2166,N_1886,N_1942);
and U2167 (N_2167,N_1955,N_1877);
nor U2168 (N_2168,N_1999,N_1853);
and U2169 (N_2169,N_1958,N_1831);
or U2170 (N_2170,N_1898,N_1932);
and U2171 (N_2171,N_1831,N_1904);
and U2172 (N_2172,N_1809,N_1945);
and U2173 (N_2173,N_1842,N_1802);
nor U2174 (N_2174,N_1851,N_1840);
nor U2175 (N_2175,N_1820,N_1875);
nor U2176 (N_2176,N_1971,N_1966);
or U2177 (N_2177,N_1988,N_1868);
nand U2178 (N_2178,N_1966,N_1993);
nand U2179 (N_2179,N_1932,N_1955);
or U2180 (N_2180,N_1950,N_1828);
nor U2181 (N_2181,N_1889,N_1861);
nand U2182 (N_2182,N_1974,N_1977);
xor U2183 (N_2183,N_1903,N_1966);
nand U2184 (N_2184,N_1841,N_1912);
or U2185 (N_2185,N_1877,N_1956);
or U2186 (N_2186,N_1962,N_1899);
nor U2187 (N_2187,N_1901,N_1862);
and U2188 (N_2188,N_1830,N_1845);
or U2189 (N_2189,N_1940,N_1802);
or U2190 (N_2190,N_1893,N_1979);
nor U2191 (N_2191,N_1862,N_1962);
xnor U2192 (N_2192,N_1915,N_1926);
or U2193 (N_2193,N_1991,N_1970);
and U2194 (N_2194,N_1914,N_1898);
nand U2195 (N_2195,N_1843,N_1909);
and U2196 (N_2196,N_1845,N_1926);
and U2197 (N_2197,N_1861,N_1844);
and U2198 (N_2198,N_1811,N_1922);
nor U2199 (N_2199,N_1995,N_1962);
nor U2200 (N_2200,N_2074,N_2153);
or U2201 (N_2201,N_2139,N_2065);
nand U2202 (N_2202,N_2133,N_2167);
nand U2203 (N_2203,N_2147,N_2186);
xor U2204 (N_2204,N_2094,N_2113);
or U2205 (N_2205,N_2150,N_2148);
or U2206 (N_2206,N_2039,N_2028);
nor U2207 (N_2207,N_2143,N_2000);
nor U2208 (N_2208,N_2189,N_2140);
nor U2209 (N_2209,N_2125,N_2043);
nand U2210 (N_2210,N_2103,N_2062);
nand U2211 (N_2211,N_2124,N_2131);
nand U2212 (N_2212,N_2044,N_2055);
xnor U2213 (N_2213,N_2025,N_2106);
nor U2214 (N_2214,N_2076,N_2026);
nor U2215 (N_2215,N_2109,N_2061);
nand U2216 (N_2216,N_2088,N_2049);
nand U2217 (N_2217,N_2059,N_2168);
xnor U2218 (N_2218,N_2018,N_2157);
nor U2219 (N_2219,N_2081,N_2110);
nor U2220 (N_2220,N_2101,N_2117);
and U2221 (N_2221,N_2164,N_2091);
nor U2222 (N_2222,N_2116,N_2036);
or U2223 (N_2223,N_2060,N_2171);
xor U2224 (N_2224,N_2198,N_2102);
nor U2225 (N_2225,N_2086,N_2122);
and U2226 (N_2226,N_2008,N_2041);
and U2227 (N_2227,N_2134,N_2111);
nor U2228 (N_2228,N_2084,N_2033);
nor U2229 (N_2229,N_2115,N_2181);
or U2230 (N_2230,N_2191,N_2123);
nor U2231 (N_2231,N_2089,N_2172);
nor U2232 (N_2232,N_2021,N_2058);
and U2233 (N_2233,N_2146,N_2096);
nor U2234 (N_2234,N_2114,N_2112);
nand U2235 (N_2235,N_2161,N_2073);
and U2236 (N_2236,N_2010,N_2128);
and U2237 (N_2237,N_2075,N_2173);
and U2238 (N_2238,N_2022,N_2079);
and U2239 (N_2239,N_2174,N_2183);
xor U2240 (N_2240,N_2137,N_2141);
nor U2241 (N_2241,N_2035,N_2066);
nand U2242 (N_2242,N_2006,N_2046);
or U2243 (N_2243,N_2194,N_2087);
and U2244 (N_2244,N_2144,N_2014);
nand U2245 (N_2245,N_2027,N_2132);
nand U2246 (N_2246,N_2130,N_2180);
nand U2247 (N_2247,N_2188,N_2048);
nand U2248 (N_2248,N_2176,N_2121);
or U2249 (N_2249,N_2195,N_2077);
xnor U2250 (N_2250,N_2078,N_2151);
xnor U2251 (N_2251,N_2070,N_2142);
or U2252 (N_2252,N_2197,N_2024);
nand U2253 (N_2253,N_2175,N_2193);
or U2254 (N_2254,N_2119,N_2199);
nor U2255 (N_2255,N_2080,N_2162);
nor U2256 (N_2256,N_2083,N_2104);
and U2257 (N_2257,N_2145,N_2038);
nor U2258 (N_2258,N_2082,N_2013);
xor U2259 (N_2259,N_2052,N_2154);
nand U2260 (N_2260,N_2163,N_2050);
nand U2261 (N_2261,N_2057,N_2042);
xnor U2262 (N_2262,N_2129,N_2179);
or U2263 (N_2263,N_2069,N_2158);
or U2264 (N_2264,N_2085,N_2003);
xnor U2265 (N_2265,N_2100,N_2155);
nand U2266 (N_2266,N_2149,N_2092);
nand U2267 (N_2267,N_2015,N_2030);
nor U2268 (N_2268,N_2045,N_2127);
and U2269 (N_2269,N_2165,N_2063);
nor U2270 (N_2270,N_2107,N_2009);
nand U2271 (N_2271,N_2031,N_2170);
and U2272 (N_2272,N_2120,N_2185);
nor U2273 (N_2273,N_2004,N_2056);
nand U2274 (N_2274,N_2002,N_2156);
and U2275 (N_2275,N_2196,N_2054);
and U2276 (N_2276,N_2097,N_2166);
or U2277 (N_2277,N_2182,N_2053);
or U2278 (N_2278,N_2071,N_2105);
or U2279 (N_2279,N_2159,N_2034);
and U2280 (N_2280,N_2019,N_2047);
nor U2281 (N_2281,N_2192,N_2051);
nor U2282 (N_2282,N_2017,N_2072);
and U2283 (N_2283,N_2023,N_2064);
nor U2284 (N_2284,N_2005,N_2001);
or U2285 (N_2285,N_2011,N_2108);
or U2286 (N_2286,N_2169,N_2099);
and U2287 (N_2287,N_2187,N_2177);
and U2288 (N_2288,N_2098,N_2190);
nor U2289 (N_2289,N_2067,N_2037);
nor U2290 (N_2290,N_2007,N_2012);
nand U2291 (N_2291,N_2093,N_2136);
nand U2292 (N_2292,N_2135,N_2126);
nor U2293 (N_2293,N_2178,N_2152);
or U2294 (N_2294,N_2020,N_2184);
nor U2295 (N_2295,N_2160,N_2040);
and U2296 (N_2296,N_2090,N_2016);
nor U2297 (N_2297,N_2138,N_2118);
nand U2298 (N_2298,N_2029,N_2095);
and U2299 (N_2299,N_2068,N_2032);
nand U2300 (N_2300,N_2086,N_2078);
or U2301 (N_2301,N_2023,N_2042);
nand U2302 (N_2302,N_2193,N_2009);
or U2303 (N_2303,N_2008,N_2120);
or U2304 (N_2304,N_2168,N_2110);
nand U2305 (N_2305,N_2091,N_2057);
nor U2306 (N_2306,N_2002,N_2134);
nand U2307 (N_2307,N_2001,N_2029);
or U2308 (N_2308,N_2092,N_2063);
xor U2309 (N_2309,N_2098,N_2077);
or U2310 (N_2310,N_2116,N_2198);
and U2311 (N_2311,N_2121,N_2037);
or U2312 (N_2312,N_2118,N_2098);
and U2313 (N_2313,N_2173,N_2093);
nor U2314 (N_2314,N_2065,N_2037);
or U2315 (N_2315,N_2142,N_2078);
xor U2316 (N_2316,N_2092,N_2154);
nor U2317 (N_2317,N_2179,N_2027);
and U2318 (N_2318,N_2038,N_2023);
nor U2319 (N_2319,N_2112,N_2177);
nor U2320 (N_2320,N_2036,N_2014);
and U2321 (N_2321,N_2174,N_2082);
nor U2322 (N_2322,N_2185,N_2190);
and U2323 (N_2323,N_2159,N_2134);
and U2324 (N_2324,N_2058,N_2160);
and U2325 (N_2325,N_2079,N_2095);
nor U2326 (N_2326,N_2143,N_2042);
nand U2327 (N_2327,N_2131,N_2176);
and U2328 (N_2328,N_2089,N_2186);
and U2329 (N_2329,N_2092,N_2076);
nor U2330 (N_2330,N_2119,N_2138);
xnor U2331 (N_2331,N_2196,N_2129);
or U2332 (N_2332,N_2023,N_2008);
nor U2333 (N_2333,N_2103,N_2133);
or U2334 (N_2334,N_2030,N_2032);
nand U2335 (N_2335,N_2185,N_2033);
xor U2336 (N_2336,N_2148,N_2043);
xor U2337 (N_2337,N_2059,N_2005);
and U2338 (N_2338,N_2188,N_2165);
and U2339 (N_2339,N_2021,N_2032);
nor U2340 (N_2340,N_2168,N_2070);
or U2341 (N_2341,N_2115,N_2009);
nor U2342 (N_2342,N_2187,N_2120);
xnor U2343 (N_2343,N_2170,N_2054);
xor U2344 (N_2344,N_2175,N_2033);
or U2345 (N_2345,N_2195,N_2089);
nor U2346 (N_2346,N_2038,N_2143);
or U2347 (N_2347,N_2153,N_2066);
nor U2348 (N_2348,N_2011,N_2158);
and U2349 (N_2349,N_2165,N_2104);
nor U2350 (N_2350,N_2144,N_2076);
nor U2351 (N_2351,N_2168,N_2025);
xor U2352 (N_2352,N_2191,N_2177);
nand U2353 (N_2353,N_2140,N_2162);
nand U2354 (N_2354,N_2162,N_2168);
nor U2355 (N_2355,N_2137,N_2002);
nand U2356 (N_2356,N_2172,N_2173);
nand U2357 (N_2357,N_2119,N_2023);
xor U2358 (N_2358,N_2041,N_2060);
xor U2359 (N_2359,N_2114,N_2093);
nand U2360 (N_2360,N_2186,N_2160);
or U2361 (N_2361,N_2090,N_2029);
or U2362 (N_2362,N_2122,N_2022);
xor U2363 (N_2363,N_2143,N_2174);
or U2364 (N_2364,N_2072,N_2020);
or U2365 (N_2365,N_2066,N_2048);
or U2366 (N_2366,N_2000,N_2166);
nor U2367 (N_2367,N_2026,N_2023);
or U2368 (N_2368,N_2195,N_2185);
and U2369 (N_2369,N_2144,N_2057);
nor U2370 (N_2370,N_2049,N_2006);
nand U2371 (N_2371,N_2161,N_2015);
or U2372 (N_2372,N_2107,N_2142);
or U2373 (N_2373,N_2026,N_2111);
or U2374 (N_2374,N_2040,N_2044);
or U2375 (N_2375,N_2025,N_2135);
nand U2376 (N_2376,N_2188,N_2181);
or U2377 (N_2377,N_2198,N_2143);
nor U2378 (N_2378,N_2189,N_2149);
nor U2379 (N_2379,N_2189,N_2004);
nand U2380 (N_2380,N_2021,N_2035);
or U2381 (N_2381,N_2028,N_2057);
or U2382 (N_2382,N_2089,N_2059);
nand U2383 (N_2383,N_2039,N_2174);
nand U2384 (N_2384,N_2182,N_2061);
nand U2385 (N_2385,N_2068,N_2158);
and U2386 (N_2386,N_2101,N_2184);
nor U2387 (N_2387,N_2188,N_2036);
nand U2388 (N_2388,N_2004,N_2085);
xor U2389 (N_2389,N_2038,N_2040);
xor U2390 (N_2390,N_2150,N_2115);
nand U2391 (N_2391,N_2191,N_2057);
and U2392 (N_2392,N_2191,N_2146);
and U2393 (N_2393,N_2169,N_2148);
and U2394 (N_2394,N_2126,N_2006);
nor U2395 (N_2395,N_2089,N_2128);
and U2396 (N_2396,N_2103,N_2188);
nand U2397 (N_2397,N_2052,N_2144);
nand U2398 (N_2398,N_2044,N_2111);
nor U2399 (N_2399,N_2153,N_2118);
or U2400 (N_2400,N_2388,N_2323);
nor U2401 (N_2401,N_2286,N_2260);
or U2402 (N_2402,N_2233,N_2259);
or U2403 (N_2403,N_2230,N_2207);
or U2404 (N_2404,N_2270,N_2338);
nor U2405 (N_2405,N_2393,N_2303);
nand U2406 (N_2406,N_2296,N_2324);
nand U2407 (N_2407,N_2337,N_2265);
nor U2408 (N_2408,N_2316,N_2343);
xor U2409 (N_2409,N_2222,N_2390);
and U2410 (N_2410,N_2385,N_2267);
and U2411 (N_2411,N_2368,N_2225);
or U2412 (N_2412,N_2387,N_2386);
nand U2413 (N_2413,N_2301,N_2363);
nor U2414 (N_2414,N_2282,N_2320);
nand U2415 (N_2415,N_2284,N_2309);
and U2416 (N_2416,N_2208,N_2322);
nand U2417 (N_2417,N_2242,N_2354);
and U2418 (N_2418,N_2213,N_2353);
or U2419 (N_2419,N_2255,N_2352);
nand U2420 (N_2420,N_2326,N_2277);
or U2421 (N_2421,N_2399,N_2332);
or U2422 (N_2422,N_2261,N_2351);
and U2423 (N_2423,N_2330,N_2329);
nor U2424 (N_2424,N_2345,N_2218);
nor U2425 (N_2425,N_2203,N_2220);
or U2426 (N_2426,N_2310,N_2362);
or U2427 (N_2427,N_2271,N_2331);
or U2428 (N_2428,N_2238,N_2313);
or U2429 (N_2429,N_2202,N_2305);
xnor U2430 (N_2430,N_2272,N_2254);
nor U2431 (N_2431,N_2361,N_2273);
nand U2432 (N_2432,N_2283,N_2325);
nand U2433 (N_2433,N_2371,N_2302);
nand U2434 (N_2434,N_2381,N_2367);
and U2435 (N_2435,N_2299,N_2257);
nor U2436 (N_2436,N_2266,N_2221);
or U2437 (N_2437,N_2336,N_2212);
nor U2438 (N_2438,N_2344,N_2228);
xnor U2439 (N_2439,N_2375,N_2319);
nor U2440 (N_2440,N_2278,N_2364);
and U2441 (N_2441,N_2226,N_2374);
nand U2442 (N_2442,N_2245,N_2205);
and U2443 (N_2443,N_2250,N_2377);
and U2444 (N_2444,N_2223,N_2300);
and U2445 (N_2445,N_2281,N_2204);
nor U2446 (N_2446,N_2378,N_2280);
or U2447 (N_2447,N_2334,N_2392);
nor U2448 (N_2448,N_2246,N_2306);
or U2449 (N_2449,N_2297,N_2376);
nand U2450 (N_2450,N_2235,N_2335);
or U2451 (N_2451,N_2201,N_2318);
or U2452 (N_2452,N_2237,N_2360);
xor U2453 (N_2453,N_2312,N_2268);
or U2454 (N_2454,N_2210,N_2285);
nand U2455 (N_2455,N_2241,N_2249);
and U2456 (N_2456,N_2380,N_2274);
nor U2457 (N_2457,N_2216,N_2317);
xnor U2458 (N_2458,N_2311,N_2350);
or U2459 (N_2459,N_2200,N_2236);
nor U2460 (N_2460,N_2379,N_2339);
or U2461 (N_2461,N_2234,N_2397);
nand U2462 (N_2462,N_2276,N_2358);
and U2463 (N_2463,N_2215,N_2346);
and U2464 (N_2464,N_2333,N_2206);
or U2465 (N_2465,N_2369,N_2224);
and U2466 (N_2466,N_2384,N_2275);
or U2467 (N_2467,N_2217,N_2355);
and U2468 (N_2468,N_2349,N_2264);
and U2469 (N_2469,N_2227,N_2251);
or U2470 (N_2470,N_2356,N_2288);
nor U2471 (N_2471,N_2359,N_2391);
or U2472 (N_2472,N_2253,N_2294);
nor U2473 (N_2473,N_2229,N_2248);
nor U2474 (N_2474,N_2373,N_2394);
nor U2475 (N_2475,N_2366,N_2308);
or U2476 (N_2476,N_2295,N_2247);
and U2477 (N_2477,N_2342,N_2211);
and U2478 (N_2478,N_2214,N_2365);
nand U2479 (N_2479,N_2258,N_2232);
nand U2480 (N_2480,N_2348,N_2321);
xor U2481 (N_2481,N_2240,N_2279);
nor U2482 (N_2482,N_2395,N_2269);
xnor U2483 (N_2483,N_2327,N_2389);
and U2484 (N_2484,N_2370,N_2357);
nor U2485 (N_2485,N_2256,N_2287);
nand U2486 (N_2486,N_2291,N_2262);
nor U2487 (N_2487,N_2209,N_2340);
and U2488 (N_2488,N_2398,N_2307);
xnor U2489 (N_2489,N_2289,N_2382);
or U2490 (N_2490,N_2293,N_2314);
nand U2491 (N_2491,N_2252,N_2244);
nor U2492 (N_2492,N_2298,N_2304);
or U2493 (N_2493,N_2292,N_2239);
nand U2494 (N_2494,N_2347,N_2243);
nor U2495 (N_2495,N_2219,N_2341);
and U2496 (N_2496,N_2372,N_2231);
nor U2497 (N_2497,N_2396,N_2383);
and U2498 (N_2498,N_2263,N_2290);
xor U2499 (N_2499,N_2328,N_2315);
and U2500 (N_2500,N_2323,N_2350);
or U2501 (N_2501,N_2309,N_2369);
or U2502 (N_2502,N_2270,N_2354);
nand U2503 (N_2503,N_2302,N_2368);
nand U2504 (N_2504,N_2309,N_2271);
nor U2505 (N_2505,N_2243,N_2354);
nand U2506 (N_2506,N_2384,N_2246);
nor U2507 (N_2507,N_2371,N_2382);
or U2508 (N_2508,N_2320,N_2293);
nor U2509 (N_2509,N_2248,N_2375);
nor U2510 (N_2510,N_2289,N_2300);
and U2511 (N_2511,N_2254,N_2283);
and U2512 (N_2512,N_2210,N_2323);
nor U2513 (N_2513,N_2369,N_2303);
or U2514 (N_2514,N_2226,N_2350);
and U2515 (N_2515,N_2207,N_2340);
or U2516 (N_2516,N_2285,N_2325);
xnor U2517 (N_2517,N_2363,N_2390);
nand U2518 (N_2518,N_2326,N_2359);
nand U2519 (N_2519,N_2206,N_2287);
or U2520 (N_2520,N_2288,N_2269);
or U2521 (N_2521,N_2300,N_2305);
nand U2522 (N_2522,N_2345,N_2240);
xnor U2523 (N_2523,N_2291,N_2282);
xor U2524 (N_2524,N_2277,N_2376);
and U2525 (N_2525,N_2214,N_2307);
or U2526 (N_2526,N_2394,N_2313);
or U2527 (N_2527,N_2246,N_2397);
or U2528 (N_2528,N_2231,N_2360);
and U2529 (N_2529,N_2235,N_2297);
or U2530 (N_2530,N_2350,N_2293);
nor U2531 (N_2531,N_2207,N_2356);
xor U2532 (N_2532,N_2302,N_2316);
nand U2533 (N_2533,N_2239,N_2299);
and U2534 (N_2534,N_2332,N_2341);
nand U2535 (N_2535,N_2323,N_2250);
and U2536 (N_2536,N_2357,N_2220);
or U2537 (N_2537,N_2319,N_2204);
and U2538 (N_2538,N_2297,N_2320);
nor U2539 (N_2539,N_2337,N_2269);
and U2540 (N_2540,N_2309,N_2362);
nand U2541 (N_2541,N_2308,N_2262);
or U2542 (N_2542,N_2263,N_2297);
nand U2543 (N_2543,N_2214,N_2220);
xor U2544 (N_2544,N_2236,N_2354);
or U2545 (N_2545,N_2280,N_2335);
or U2546 (N_2546,N_2229,N_2235);
or U2547 (N_2547,N_2264,N_2225);
and U2548 (N_2548,N_2309,N_2214);
and U2549 (N_2549,N_2356,N_2281);
and U2550 (N_2550,N_2222,N_2287);
nand U2551 (N_2551,N_2290,N_2280);
nor U2552 (N_2552,N_2284,N_2330);
xor U2553 (N_2553,N_2237,N_2307);
nand U2554 (N_2554,N_2297,N_2330);
nor U2555 (N_2555,N_2366,N_2392);
and U2556 (N_2556,N_2205,N_2293);
xnor U2557 (N_2557,N_2369,N_2397);
nand U2558 (N_2558,N_2268,N_2348);
or U2559 (N_2559,N_2259,N_2367);
nor U2560 (N_2560,N_2274,N_2240);
nand U2561 (N_2561,N_2254,N_2291);
and U2562 (N_2562,N_2223,N_2380);
xor U2563 (N_2563,N_2218,N_2390);
or U2564 (N_2564,N_2216,N_2320);
nor U2565 (N_2565,N_2252,N_2314);
and U2566 (N_2566,N_2356,N_2395);
nor U2567 (N_2567,N_2210,N_2274);
and U2568 (N_2568,N_2271,N_2206);
or U2569 (N_2569,N_2315,N_2349);
nor U2570 (N_2570,N_2389,N_2302);
and U2571 (N_2571,N_2296,N_2384);
nand U2572 (N_2572,N_2333,N_2292);
xnor U2573 (N_2573,N_2243,N_2234);
and U2574 (N_2574,N_2250,N_2346);
nand U2575 (N_2575,N_2261,N_2290);
xnor U2576 (N_2576,N_2223,N_2399);
and U2577 (N_2577,N_2227,N_2215);
nor U2578 (N_2578,N_2280,N_2278);
and U2579 (N_2579,N_2315,N_2336);
nor U2580 (N_2580,N_2210,N_2372);
or U2581 (N_2581,N_2322,N_2306);
nor U2582 (N_2582,N_2261,N_2277);
xor U2583 (N_2583,N_2380,N_2368);
and U2584 (N_2584,N_2357,N_2260);
nand U2585 (N_2585,N_2254,N_2329);
nand U2586 (N_2586,N_2230,N_2336);
or U2587 (N_2587,N_2329,N_2252);
or U2588 (N_2588,N_2233,N_2213);
or U2589 (N_2589,N_2331,N_2239);
nor U2590 (N_2590,N_2252,N_2305);
or U2591 (N_2591,N_2231,N_2235);
or U2592 (N_2592,N_2352,N_2358);
nor U2593 (N_2593,N_2250,N_2370);
nor U2594 (N_2594,N_2315,N_2331);
xor U2595 (N_2595,N_2267,N_2213);
or U2596 (N_2596,N_2314,N_2262);
nand U2597 (N_2597,N_2365,N_2208);
or U2598 (N_2598,N_2326,N_2280);
and U2599 (N_2599,N_2247,N_2336);
nand U2600 (N_2600,N_2513,N_2512);
and U2601 (N_2601,N_2456,N_2434);
nor U2602 (N_2602,N_2482,N_2492);
xnor U2603 (N_2603,N_2465,N_2478);
nand U2604 (N_2604,N_2439,N_2497);
and U2605 (N_2605,N_2485,N_2426);
xor U2606 (N_2606,N_2444,N_2453);
nor U2607 (N_2607,N_2408,N_2584);
or U2608 (N_2608,N_2580,N_2522);
nand U2609 (N_2609,N_2582,N_2493);
or U2610 (N_2610,N_2594,N_2454);
nor U2611 (N_2611,N_2447,N_2529);
nor U2612 (N_2612,N_2515,N_2536);
and U2613 (N_2613,N_2409,N_2597);
or U2614 (N_2614,N_2587,N_2457);
xnor U2615 (N_2615,N_2468,N_2441);
xnor U2616 (N_2616,N_2538,N_2504);
nor U2617 (N_2617,N_2437,N_2541);
and U2618 (N_2618,N_2574,N_2523);
xnor U2619 (N_2619,N_2421,N_2502);
nor U2620 (N_2620,N_2476,N_2496);
and U2621 (N_2621,N_2539,N_2411);
nand U2622 (N_2622,N_2585,N_2475);
xnor U2623 (N_2623,N_2464,N_2532);
or U2624 (N_2624,N_2559,N_2481);
nor U2625 (N_2625,N_2448,N_2501);
nor U2626 (N_2626,N_2484,N_2413);
xnor U2627 (N_2627,N_2498,N_2480);
xnor U2628 (N_2628,N_2596,N_2443);
and U2629 (N_2629,N_2583,N_2568);
nand U2630 (N_2630,N_2517,N_2562);
nor U2631 (N_2631,N_2459,N_2458);
or U2632 (N_2632,N_2429,N_2570);
nand U2633 (N_2633,N_2416,N_2495);
nand U2634 (N_2634,N_2507,N_2462);
nand U2635 (N_2635,N_2543,N_2506);
and U2636 (N_2636,N_2514,N_2567);
and U2637 (N_2637,N_2440,N_2564);
nand U2638 (N_2638,N_2557,N_2436);
nand U2639 (N_2639,N_2494,N_2572);
nor U2640 (N_2640,N_2508,N_2544);
or U2641 (N_2641,N_2467,N_2450);
nor U2642 (N_2642,N_2546,N_2487);
and U2643 (N_2643,N_2591,N_2511);
nand U2644 (N_2644,N_2586,N_2460);
and U2645 (N_2645,N_2470,N_2589);
xnor U2646 (N_2646,N_2466,N_2578);
or U2647 (N_2647,N_2540,N_2535);
or U2648 (N_2648,N_2404,N_2442);
or U2649 (N_2649,N_2486,N_2431);
and U2650 (N_2650,N_2424,N_2446);
nor U2651 (N_2651,N_2577,N_2537);
and U2652 (N_2652,N_2417,N_2569);
or U2653 (N_2653,N_2520,N_2433);
and U2654 (N_2654,N_2415,N_2451);
or U2655 (N_2655,N_2549,N_2428);
or U2656 (N_2656,N_2518,N_2526);
and U2657 (N_2657,N_2412,N_2438);
nand U2658 (N_2658,N_2472,N_2531);
or U2659 (N_2659,N_2556,N_2519);
or U2660 (N_2660,N_2473,N_2547);
and U2661 (N_2661,N_2400,N_2410);
and U2662 (N_2662,N_2427,N_2505);
nor U2663 (N_2663,N_2479,N_2533);
nand U2664 (N_2664,N_2499,N_2554);
or U2665 (N_2665,N_2491,N_2405);
nand U2666 (N_2666,N_2598,N_2566);
nand U2667 (N_2667,N_2422,N_2432);
or U2668 (N_2668,N_2452,N_2555);
nor U2669 (N_2669,N_2489,N_2471);
nor U2670 (N_2670,N_2590,N_2561);
xnor U2671 (N_2671,N_2418,N_2488);
and U2672 (N_2672,N_2414,N_2402);
or U2673 (N_2673,N_2474,N_2560);
or U2674 (N_2674,N_2500,N_2469);
xnor U2675 (N_2675,N_2575,N_2563);
nand U2676 (N_2676,N_2525,N_2401);
xor U2677 (N_2677,N_2573,N_2581);
and U2678 (N_2678,N_2406,N_2524);
or U2679 (N_2679,N_2449,N_2510);
nand U2680 (N_2680,N_2551,N_2435);
xor U2681 (N_2681,N_2490,N_2419);
or U2682 (N_2682,N_2425,N_2576);
nand U2683 (N_2683,N_2552,N_2530);
nand U2684 (N_2684,N_2545,N_2579);
or U2685 (N_2685,N_2483,N_2558);
nor U2686 (N_2686,N_2423,N_2593);
or U2687 (N_2687,N_2565,N_2542);
xnor U2688 (N_2688,N_2403,N_2550);
xnor U2689 (N_2689,N_2420,N_2477);
nand U2690 (N_2690,N_2463,N_2592);
nand U2691 (N_2691,N_2528,N_2534);
nor U2692 (N_2692,N_2445,N_2509);
nand U2693 (N_2693,N_2588,N_2407);
nor U2694 (N_2694,N_2521,N_2455);
nor U2695 (N_2695,N_2461,N_2503);
or U2696 (N_2696,N_2595,N_2553);
and U2697 (N_2697,N_2599,N_2527);
or U2698 (N_2698,N_2548,N_2571);
nor U2699 (N_2699,N_2430,N_2516);
or U2700 (N_2700,N_2545,N_2521);
nand U2701 (N_2701,N_2516,N_2526);
nor U2702 (N_2702,N_2573,N_2565);
or U2703 (N_2703,N_2597,N_2580);
nor U2704 (N_2704,N_2403,N_2559);
or U2705 (N_2705,N_2575,N_2594);
xnor U2706 (N_2706,N_2442,N_2517);
and U2707 (N_2707,N_2516,N_2409);
xnor U2708 (N_2708,N_2572,N_2530);
nand U2709 (N_2709,N_2423,N_2440);
nor U2710 (N_2710,N_2502,N_2596);
nor U2711 (N_2711,N_2577,N_2410);
or U2712 (N_2712,N_2510,N_2568);
xor U2713 (N_2713,N_2403,N_2436);
nor U2714 (N_2714,N_2484,N_2477);
and U2715 (N_2715,N_2503,N_2514);
nor U2716 (N_2716,N_2432,N_2412);
or U2717 (N_2717,N_2497,N_2548);
nor U2718 (N_2718,N_2582,N_2547);
nand U2719 (N_2719,N_2581,N_2424);
and U2720 (N_2720,N_2529,N_2436);
or U2721 (N_2721,N_2548,N_2520);
nand U2722 (N_2722,N_2464,N_2567);
and U2723 (N_2723,N_2555,N_2472);
or U2724 (N_2724,N_2554,N_2565);
nor U2725 (N_2725,N_2525,N_2501);
nor U2726 (N_2726,N_2574,N_2499);
xnor U2727 (N_2727,N_2544,N_2551);
and U2728 (N_2728,N_2556,N_2462);
nor U2729 (N_2729,N_2588,N_2466);
or U2730 (N_2730,N_2568,N_2546);
and U2731 (N_2731,N_2595,N_2421);
nand U2732 (N_2732,N_2463,N_2525);
and U2733 (N_2733,N_2599,N_2511);
or U2734 (N_2734,N_2596,N_2536);
and U2735 (N_2735,N_2561,N_2489);
nand U2736 (N_2736,N_2408,N_2594);
or U2737 (N_2737,N_2418,N_2520);
and U2738 (N_2738,N_2478,N_2546);
nor U2739 (N_2739,N_2504,N_2528);
nor U2740 (N_2740,N_2447,N_2403);
xor U2741 (N_2741,N_2431,N_2437);
nand U2742 (N_2742,N_2548,N_2500);
or U2743 (N_2743,N_2405,N_2448);
nor U2744 (N_2744,N_2581,N_2478);
xnor U2745 (N_2745,N_2493,N_2412);
and U2746 (N_2746,N_2521,N_2590);
nor U2747 (N_2747,N_2496,N_2410);
nor U2748 (N_2748,N_2444,N_2507);
nor U2749 (N_2749,N_2467,N_2529);
nor U2750 (N_2750,N_2509,N_2458);
nand U2751 (N_2751,N_2535,N_2597);
nand U2752 (N_2752,N_2458,N_2477);
or U2753 (N_2753,N_2567,N_2510);
nor U2754 (N_2754,N_2586,N_2581);
or U2755 (N_2755,N_2545,N_2446);
xnor U2756 (N_2756,N_2567,N_2468);
xnor U2757 (N_2757,N_2592,N_2509);
or U2758 (N_2758,N_2463,N_2577);
nor U2759 (N_2759,N_2455,N_2571);
nor U2760 (N_2760,N_2599,N_2591);
or U2761 (N_2761,N_2573,N_2471);
and U2762 (N_2762,N_2567,N_2561);
nand U2763 (N_2763,N_2567,N_2450);
or U2764 (N_2764,N_2434,N_2494);
and U2765 (N_2765,N_2592,N_2419);
nand U2766 (N_2766,N_2488,N_2477);
and U2767 (N_2767,N_2407,N_2474);
or U2768 (N_2768,N_2433,N_2485);
nor U2769 (N_2769,N_2539,N_2416);
xor U2770 (N_2770,N_2400,N_2559);
or U2771 (N_2771,N_2486,N_2471);
and U2772 (N_2772,N_2496,N_2425);
and U2773 (N_2773,N_2515,N_2534);
nand U2774 (N_2774,N_2526,N_2426);
and U2775 (N_2775,N_2487,N_2469);
and U2776 (N_2776,N_2562,N_2534);
nor U2777 (N_2777,N_2451,N_2550);
nor U2778 (N_2778,N_2456,N_2547);
xnor U2779 (N_2779,N_2426,N_2518);
nor U2780 (N_2780,N_2418,N_2478);
or U2781 (N_2781,N_2472,N_2496);
nor U2782 (N_2782,N_2519,N_2597);
nand U2783 (N_2783,N_2536,N_2528);
and U2784 (N_2784,N_2477,N_2436);
nand U2785 (N_2785,N_2537,N_2431);
and U2786 (N_2786,N_2565,N_2547);
xor U2787 (N_2787,N_2521,N_2478);
nor U2788 (N_2788,N_2560,N_2510);
or U2789 (N_2789,N_2481,N_2422);
and U2790 (N_2790,N_2486,N_2462);
or U2791 (N_2791,N_2489,N_2582);
and U2792 (N_2792,N_2518,N_2489);
and U2793 (N_2793,N_2422,N_2498);
or U2794 (N_2794,N_2418,N_2460);
nor U2795 (N_2795,N_2459,N_2488);
nand U2796 (N_2796,N_2522,N_2468);
nand U2797 (N_2797,N_2508,N_2543);
or U2798 (N_2798,N_2563,N_2483);
nand U2799 (N_2799,N_2534,N_2574);
and U2800 (N_2800,N_2637,N_2636);
nand U2801 (N_2801,N_2694,N_2661);
and U2802 (N_2802,N_2794,N_2759);
nor U2803 (N_2803,N_2689,N_2666);
nor U2804 (N_2804,N_2798,N_2617);
and U2805 (N_2805,N_2796,N_2647);
nand U2806 (N_2806,N_2621,N_2630);
and U2807 (N_2807,N_2700,N_2656);
nand U2808 (N_2808,N_2683,N_2793);
nor U2809 (N_2809,N_2721,N_2693);
nand U2810 (N_2810,N_2601,N_2677);
xor U2811 (N_2811,N_2662,N_2745);
and U2812 (N_2812,N_2643,N_2775);
or U2813 (N_2813,N_2738,N_2633);
and U2814 (N_2814,N_2604,N_2675);
xor U2815 (N_2815,N_2697,N_2639);
and U2816 (N_2816,N_2641,N_2751);
nor U2817 (N_2817,N_2672,N_2685);
nor U2818 (N_2818,N_2783,N_2702);
and U2819 (N_2819,N_2771,N_2752);
and U2820 (N_2820,N_2781,N_2603);
xnor U2821 (N_2821,N_2784,N_2762);
nor U2822 (N_2822,N_2786,N_2717);
and U2823 (N_2823,N_2628,N_2776);
and U2824 (N_2824,N_2782,N_2620);
nor U2825 (N_2825,N_2769,N_2767);
nor U2826 (N_2826,N_2724,N_2787);
nor U2827 (N_2827,N_2734,N_2765);
nor U2828 (N_2828,N_2763,N_2692);
nand U2829 (N_2829,N_2610,N_2618);
or U2830 (N_2830,N_2723,N_2753);
and U2831 (N_2831,N_2663,N_2703);
nand U2832 (N_2832,N_2778,N_2726);
nor U2833 (N_2833,N_2736,N_2710);
nor U2834 (N_2834,N_2705,N_2695);
and U2835 (N_2835,N_2797,N_2614);
nor U2836 (N_2836,N_2606,N_2758);
and U2837 (N_2837,N_2640,N_2686);
and U2838 (N_2838,N_2788,N_2671);
or U2839 (N_2839,N_2612,N_2664);
nand U2840 (N_2840,N_2655,N_2668);
nand U2841 (N_2841,N_2725,N_2756);
or U2842 (N_2842,N_2607,N_2707);
nand U2843 (N_2843,N_2748,N_2737);
or U2844 (N_2844,N_2657,N_2605);
or U2845 (N_2845,N_2667,N_2651);
nor U2846 (N_2846,N_2709,N_2680);
nand U2847 (N_2847,N_2653,N_2619);
nand U2848 (N_2848,N_2773,N_2746);
nand U2849 (N_2849,N_2611,N_2774);
nor U2850 (N_2850,N_2760,N_2741);
xor U2851 (N_2851,N_2629,N_2730);
and U2852 (N_2852,N_2742,N_2626);
and U2853 (N_2853,N_2658,N_2799);
nand U2854 (N_2854,N_2625,N_2644);
nor U2855 (N_2855,N_2600,N_2795);
nor U2856 (N_2856,N_2708,N_2698);
xnor U2857 (N_2857,N_2659,N_2750);
nor U2858 (N_2858,N_2645,N_2650);
nand U2859 (N_2859,N_2761,N_2714);
and U2860 (N_2860,N_2669,N_2785);
or U2861 (N_2861,N_2704,N_2770);
and U2862 (N_2862,N_2648,N_2718);
or U2863 (N_2863,N_2729,N_2634);
and U2864 (N_2864,N_2711,N_2622);
or U2865 (N_2865,N_2681,N_2635);
and U2866 (N_2866,N_2732,N_2731);
and U2867 (N_2867,N_2649,N_2792);
and U2868 (N_2868,N_2768,N_2670);
nor U2869 (N_2869,N_2716,N_2757);
nor U2870 (N_2870,N_2642,N_2727);
nand U2871 (N_2871,N_2790,N_2699);
and U2872 (N_2872,N_2735,N_2713);
nor U2873 (N_2873,N_2674,N_2696);
or U2874 (N_2874,N_2632,N_2613);
and U2875 (N_2875,N_2755,N_2638);
nand U2876 (N_2876,N_2749,N_2764);
nand U2877 (N_2877,N_2766,N_2631);
nand U2878 (N_2878,N_2623,N_2646);
xor U2879 (N_2879,N_2754,N_2615);
nor U2880 (N_2880,N_2706,N_2739);
and U2881 (N_2881,N_2682,N_2609);
or U2882 (N_2882,N_2712,N_2652);
or U2883 (N_2883,N_2744,N_2720);
nand U2884 (N_2884,N_2624,N_2715);
or U2885 (N_2885,N_2777,N_2722);
nor U2886 (N_2886,N_2679,N_2602);
nor U2887 (N_2887,N_2690,N_2616);
or U2888 (N_2888,N_2780,N_2743);
or U2889 (N_2889,N_2733,N_2627);
or U2890 (N_2890,N_2779,N_2676);
and U2891 (N_2891,N_2789,N_2678);
nor U2892 (N_2892,N_2728,N_2772);
nor U2893 (N_2893,N_2654,N_2608);
and U2894 (N_2894,N_2701,N_2740);
and U2895 (N_2895,N_2688,N_2791);
or U2896 (N_2896,N_2691,N_2747);
and U2897 (N_2897,N_2719,N_2673);
nand U2898 (N_2898,N_2660,N_2687);
and U2899 (N_2899,N_2684,N_2665);
and U2900 (N_2900,N_2607,N_2687);
nand U2901 (N_2901,N_2698,N_2685);
and U2902 (N_2902,N_2713,N_2614);
nor U2903 (N_2903,N_2746,N_2614);
nor U2904 (N_2904,N_2759,N_2773);
nor U2905 (N_2905,N_2757,N_2747);
nor U2906 (N_2906,N_2678,N_2778);
nor U2907 (N_2907,N_2757,N_2793);
nor U2908 (N_2908,N_2658,N_2720);
or U2909 (N_2909,N_2705,N_2714);
and U2910 (N_2910,N_2617,N_2637);
and U2911 (N_2911,N_2747,N_2623);
nand U2912 (N_2912,N_2600,N_2783);
nand U2913 (N_2913,N_2789,N_2722);
and U2914 (N_2914,N_2696,N_2731);
and U2915 (N_2915,N_2707,N_2769);
or U2916 (N_2916,N_2795,N_2769);
nand U2917 (N_2917,N_2679,N_2656);
nor U2918 (N_2918,N_2722,N_2651);
or U2919 (N_2919,N_2687,N_2752);
or U2920 (N_2920,N_2757,N_2713);
or U2921 (N_2921,N_2720,N_2612);
and U2922 (N_2922,N_2604,N_2691);
or U2923 (N_2923,N_2794,N_2637);
and U2924 (N_2924,N_2604,N_2779);
nand U2925 (N_2925,N_2666,N_2762);
or U2926 (N_2926,N_2609,N_2789);
and U2927 (N_2927,N_2635,N_2788);
and U2928 (N_2928,N_2673,N_2676);
nand U2929 (N_2929,N_2739,N_2717);
nor U2930 (N_2930,N_2748,N_2694);
nand U2931 (N_2931,N_2755,N_2632);
or U2932 (N_2932,N_2734,N_2777);
and U2933 (N_2933,N_2727,N_2613);
nor U2934 (N_2934,N_2728,N_2691);
and U2935 (N_2935,N_2622,N_2668);
and U2936 (N_2936,N_2665,N_2786);
and U2937 (N_2937,N_2629,N_2709);
and U2938 (N_2938,N_2669,N_2627);
nand U2939 (N_2939,N_2785,N_2633);
nand U2940 (N_2940,N_2684,N_2697);
nor U2941 (N_2941,N_2783,N_2740);
or U2942 (N_2942,N_2643,N_2655);
nor U2943 (N_2943,N_2762,N_2728);
or U2944 (N_2944,N_2715,N_2752);
and U2945 (N_2945,N_2651,N_2763);
nand U2946 (N_2946,N_2747,N_2688);
and U2947 (N_2947,N_2605,N_2655);
and U2948 (N_2948,N_2656,N_2681);
or U2949 (N_2949,N_2632,N_2794);
or U2950 (N_2950,N_2763,N_2794);
nor U2951 (N_2951,N_2703,N_2604);
and U2952 (N_2952,N_2795,N_2715);
nand U2953 (N_2953,N_2659,N_2745);
or U2954 (N_2954,N_2771,N_2620);
and U2955 (N_2955,N_2685,N_2620);
or U2956 (N_2956,N_2650,N_2652);
nor U2957 (N_2957,N_2758,N_2768);
and U2958 (N_2958,N_2684,N_2644);
and U2959 (N_2959,N_2672,N_2620);
or U2960 (N_2960,N_2678,N_2700);
and U2961 (N_2961,N_2622,N_2710);
nand U2962 (N_2962,N_2616,N_2640);
or U2963 (N_2963,N_2774,N_2645);
or U2964 (N_2964,N_2621,N_2763);
nor U2965 (N_2965,N_2668,N_2695);
nor U2966 (N_2966,N_2647,N_2754);
and U2967 (N_2967,N_2606,N_2735);
xnor U2968 (N_2968,N_2740,N_2749);
xnor U2969 (N_2969,N_2714,N_2634);
nand U2970 (N_2970,N_2734,N_2610);
nand U2971 (N_2971,N_2613,N_2734);
nor U2972 (N_2972,N_2683,N_2731);
or U2973 (N_2973,N_2643,N_2708);
and U2974 (N_2974,N_2718,N_2667);
xnor U2975 (N_2975,N_2760,N_2727);
nand U2976 (N_2976,N_2687,N_2726);
nor U2977 (N_2977,N_2696,N_2699);
nor U2978 (N_2978,N_2675,N_2638);
nor U2979 (N_2979,N_2795,N_2634);
xnor U2980 (N_2980,N_2621,N_2736);
or U2981 (N_2981,N_2734,N_2788);
xor U2982 (N_2982,N_2701,N_2734);
or U2983 (N_2983,N_2757,N_2784);
nand U2984 (N_2984,N_2628,N_2710);
or U2985 (N_2985,N_2665,N_2713);
nor U2986 (N_2986,N_2693,N_2731);
nand U2987 (N_2987,N_2748,N_2662);
and U2988 (N_2988,N_2615,N_2668);
and U2989 (N_2989,N_2611,N_2646);
or U2990 (N_2990,N_2761,N_2656);
nand U2991 (N_2991,N_2609,N_2731);
nor U2992 (N_2992,N_2636,N_2747);
nor U2993 (N_2993,N_2654,N_2725);
and U2994 (N_2994,N_2763,N_2605);
and U2995 (N_2995,N_2667,N_2755);
nand U2996 (N_2996,N_2623,N_2775);
nor U2997 (N_2997,N_2688,N_2686);
xnor U2998 (N_2998,N_2640,N_2782);
or U2999 (N_2999,N_2745,N_2756);
and U3000 (N_3000,N_2947,N_2922);
nor U3001 (N_3001,N_2964,N_2814);
nand U3002 (N_3002,N_2890,N_2986);
or U3003 (N_3003,N_2999,N_2895);
xor U3004 (N_3004,N_2816,N_2841);
nor U3005 (N_3005,N_2974,N_2809);
and U3006 (N_3006,N_2845,N_2905);
nor U3007 (N_3007,N_2897,N_2908);
xnor U3008 (N_3008,N_2934,N_2998);
and U3009 (N_3009,N_2883,N_2925);
xor U3010 (N_3010,N_2924,N_2821);
or U3011 (N_3011,N_2983,N_2835);
nand U3012 (N_3012,N_2880,N_2885);
or U3013 (N_3013,N_2992,N_2965);
or U3014 (N_3014,N_2855,N_2953);
or U3015 (N_3015,N_2846,N_2938);
nand U3016 (N_3016,N_2850,N_2919);
or U3017 (N_3017,N_2881,N_2927);
or U3018 (N_3018,N_2804,N_2887);
nand U3019 (N_3019,N_2893,N_2976);
nor U3020 (N_3020,N_2932,N_2906);
nor U3021 (N_3021,N_2869,N_2987);
xnor U3022 (N_3022,N_2843,N_2854);
and U3023 (N_3023,N_2901,N_2955);
nor U3024 (N_3024,N_2871,N_2805);
nand U3025 (N_3025,N_2909,N_2904);
nor U3026 (N_3026,N_2975,N_2966);
nor U3027 (N_3027,N_2939,N_2892);
xnor U3028 (N_3028,N_2900,N_2961);
and U3029 (N_3029,N_2950,N_2811);
nand U3030 (N_3030,N_2920,N_2930);
nor U3031 (N_3031,N_2936,N_2899);
nand U3032 (N_3032,N_2954,N_2943);
and U3033 (N_3033,N_2923,N_2971);
or U3034 (N_3034,N_2826,N_2867);
or U3035 (N_3035,N_2916,N_2838);
nand U3036 (N_3036,N_2853,N_2856);
and U3037 (N_3037,N_2951,N_2870);
and U3038 (N_3038,N_2818,N_2800);
xnor U3039 (N_3039,N_2861,N_2985);
nor U3040 (N_3040,N_2839,N_2877);
nand U3041 (N_3041,N_2918,N_2865);
nor U3042 (N_3042,N_2827,N_2844);
or U3043 (N_3043,N_2913,N_2891);
nor U3044 (N_3044,N_2944,N_2902);
and U3045 (N_3045,N_2910,N_2863);
or U3046 (N_3046,N_2857,N_2847);
nand U3047 (N_3047,N_2997,N_2889);
and U3048 (N_3048,N_2832,N_2836);
nor U3049 (N_3049,N_2884,N_2833);
nand U3050 (N_3050,N_2824,N_2907);
and U3051 (N_3051,N_2803,N_2995);
and U3052 (N_3052,N_2911,N_2858);
or U3053 (N_3053,N_2878,N_2812);
nor U3054 (N_3054,N_2969,N_2852);
nand U3055 (N_3055,N_2825,N_2915);
nor U3056 (N_3056,N_2945,N_2990);
xor U3057 (N_3057,N_2848,N_2978);
nand U3058 (N_3058,N_2958,N_2942);
nand U3059 (N_3059,N_2886,N_2972);
or U3060 (N_3060,N_2866,N_2819);
or U3061 (N_3061,N_2980,N_2896);
and U3062 (N_3062,N_2921,N_2959);
xnor U3063 (N_3063,N_2875,N_2926);
nor U3064 (N_3064,N_2979,N_2973);
and U3065 (N_3065,N_2967,N_2842);
or U3066 (N_3066,N_2937,N_2837);
or U3067 (N_3067,N_2917,N_2879);
or U3068 (N_3068,N_2982,N_2807);
xnor U3069 (N_3069,N_2872,N_2948);
and U3070 (N_3070,N_2831,N_2894);
nor U3071 (N_3071,N_2956,N_2851);
nand U3072 (N_3072,N_2993,N_2876);
nand U3073 (N_3073,N_2984,N_2820);
nand U3074 (N_3074,N_2862,N_2949);
and U3075 (N_3075,N_2829,N_2888);
xnor U3076 (N_3076,N_2963,N_2914);
nand U3077 (N_3077,N_2935,N_2860);
xor U3078 (N_3078,N_2823,N_2864);
nor U3079 (N_3079,N_2977,N_2898);
nand U3080 (N_3080,N_2903,N_2989);
xor U3081 (N_3081,N_2882,N_2946);
and U3082 (N_3082,N_2840,N_2960);
or U3083 (N_3083,N_2970,N_2981);
nand U3084 (N_3084,N_2940,N_2815);
or U3085 (N_3085,N_2991,N_2933);
nand U3086 (N_3086,N_2801,N_2928);
nand U3087 (N_3087,N_2808,N_2912);
nand U3088 (N_3088,N_2810,N_2849);
nand U3089 (N_3089,N_2802,N_2868);
and U3090 (N_3090,N_2830,N_2994);
xor U3091 (N_3091,N_2828,N_2968);
and U3092 (N_3092,N_2931,N_2874);
or U3093 (N_3093,N_2957,N_2996);
nand U3094 (N_3094,N_2941,N_2834);
and U3095 (N_3095,N_2859,N_2813);
nor U3096 (N_3096,N_2873,N_2817);
nor U3097 (N_3097,N_2952,N_2822);
nor U3098 (N_3098,N_2929,N_2988);
and U3099 (N_3099,N_2806,N_2962);
or U3100 (N_3100,N_2952,N_2939);
or U3101 (N_3101,N_2871,N_2994);
or U3102 (N_3102,N_2933,N_2966);
or U3103 (N_3103,N_2939,N_2951);
nand U3104 (N_3104,N_2883,N_2923);
xor U3105 (N_3105,N_2925,N_2839);
and U3106 (N_3106,N_2908,N_2805);
nand U3107 (N_3107,N_2868,N_2909);
nand U3108 (N_3108,N_2934,N_2850);
nor U3109 (N_3109,N_2835,N_2891);
nor U3110 (N_3110,N_2894,N_2873);
or U3111 (N_3111,N_2955,N_2921);
xor U3112 (N_3112,N_2860,N_2823);
nand U3113 (N_3113,N_2819,N_2983);
and U3114 (N_3114,N_2959,N_2856);
nor U3115 (N_3115,N_2805,N_2993);
and U3116 (N_3116,N_2931,N_2900);
nand U3117 (N_3117,N_2999,N_2808);
nand U3118 (N_3118,N_2976,N_2849);
xor U3119 (N_3119,N_2818,N_2872);
and U3120 (N_3120,N_2929,N_2967);
nand U3121 (N_3121,N_2934,N_2852);
and U3122 (N_3122,N_2863,N_2902);
or U3123 (N_3123,N_2809,N_2902);
nor U3124 (N_3124,N_2941,N_2828);
or U3125 (N_3125,N_2840,N_2973);
or U3126 (N_3126,N_2905,N_2848);
nor U3127 (N_3127,N_2962,N_2921);
or U3128 (N_3128,N_2975,N_2935);
and U3129 (N_3129,N_2831,N_2860);
xor U3130 (N_3130,N_2818,N_2823);
nor U3131 (N_3131,N_2986,N_2982);
nor U3132 (N_3132,N_2804,N_2965);
nor U3133 (N_3133,N_2970,N_2915);
or U3134 (N_3134,N_2838,N_2958);
and U3135 (N_3135,N_2828,N_2988);
nand U3136 (N_3136,N_2820,N_2900);
xnor U3137 (N_3137,N_2954,N_2991);
xor U3138 (N_3138,N_2998,N_2826);
or U3139 (N_3139,N_2915,N_2826);
xor U3140 (N_3140,N_2861,N_2965);
and U3141 (N_3141,N_2847,N_2963);
nor U3142 (N_3142,N_2910,N_2874);
or U3143 (N_3143,N_2821,N_2904);
and U3144 (N_3144,N_2940,N_2937);
or U3145 (N_3145,N_2823,N_2859);
nand U3146 (N_3146,N_2910,N_2820);
or U3147 (N_3147,N_2919,N_2817);
or U3148 (N_3148,N_2804,N_2917);
nand U3149 (N_3149,N_2861,N_2882);
nor U3150 (N_3150,N_2832,N_2890);
or U3151 (N_3151,N_2927,N_2894);
nand U3152 (N_3152,N_2861,N_2869);
nand U3153 (N_3153,N_2977,N_2833);
and U3154 (N_3154,N_2905,N_2833);
nand U3155 (N_3155,N_2810,N_2895);
nor U3156 (N_3156,N_2935,N_2995);
nand U3157 (N_3157,N_2872,N_2852);
and U3158 (N_3158,N_2913,N_2825);
xor U3159 (N_3159,N_2823,N_2865);
nand U3160 (N_3160,N_2867,N_2960);
or U3161 (N_3161,N_2938,N_2852);
nand U3162 (N_3162,N_2916,N_2934);
nand U3163 (N_3163,N_2970,N_2946);
or U3164 (N_3164,N_2959,N_2973);
nand U3165 (N_3165,N_2929,N_2901);
nand U3166 (N_3166,N_2889,N_2901);
nand U3167 (N_3167,N_2897,N_2926);
nor U3168 (N_3168,N_2829,N_2959);
xnor U3169 (N_3169,N_2973,N_2937);
nor U3170 (N_3170,N_2919,N_2892);
and U3171 (N_3171,N_2830,N_2894);
and U3172 (N_3172,N_2846,N_2830);
xnor U3173 (N_3173,N_2887,N_2996);
and U3174 (N_3174,N_2848,N_2965);
nand U3175 (N_3175,N_2951,N_2925);
or U3176 (N_3176,N_2951,N_2900);
or U3177 (N_3177,N_2951,N_2957);
and U3178 (N_3178,N_2835,N_2994);
xnor U3179 (N_3179,N_2912,N_2817);
nor U3180 (N_3180,N_2904,N_2925);
nand U3181 (N_3181,N_2908,N_2836);
xor U3182 (N_3182,N_2910,N_2938);
or U3183 (N_3183,N_2938,N_2837);
or U3184 (N_3184,N_2975,N_2858);
nor U3185 (N_3185,N_2900,N_2893);
nand U3186 (N_3186,N_2910,N_2825);
and U3187 (N_3187,N_2808,N_2803);
and U3188 (N_3188,N_2888,N_2830);
or U3189 (N_3189,N_2827,N_2941);
nand U3190 (N_3190,N_2876,N_2833);
nand U3191 (N_3191,N_2927,N_2926);
or U3192 (N_3192,N_2858,N_2805);
or U3193 (N_3193,N_2978,N_2922);
nand U3194 (N_3194,N_2976,N_2802);
nand U3195 (N_3195,N_2875,N_2857);
xnor U3196 (N_3196,N_2888,N_2956);
nor U3197 (N_3197,N_2907,N_2979);
and U3198 (N_3198,N_2974,N_2902);
nand U3199 (N_3199,N_2859,N_2913);
nor U3200 (N_3200,N_3179,N_3133);
or U3201 (N_3201,N_3038,N_3043);
xor U3202 (N_3202,N_3027,N_3081);
and U3203 (N_3203,N_3055,N_3119);
xnor U3204 (N_3204,N_3028,N_3139);
nand U3205 (N_3205,N_3012,N_3091);
nand U3206 (N_3206,N_3177,N_3084);
or U3207 (N_3207,N_3068,N_3049);
nor U3208 (N_3208,N_3044,N_3198);
nand U3209 (N_3209,N_3171,N_3024);
xor U3210 (N_3210,N_3041,N_3180);
xor U3211 (N_3211,N_3196,N_3112);
or U3212 (N_3212,N_3104,N_3144);
and U3213 (N_3213,N_3037,N_3067);
and U3214 (N_3214,N_3122,N_3088);
or U3215 (N_3215,N_3064,N_3145);
nand U3216 (N_3216,N_3013,N_3129);
nor U3217 (N_3217,N_3135,N_3082);
nand U3218 (N_3218,N_3107,N_3011);
xor U3219 (N_3219,N_3142,N_3141);
or U3220 (N_3220,N_3175,N_3169);
nand U3221 (N_3221,N_3157,N_3039);
nand U3222 (N_3222,N_3158,N_3187);
and U3223 (N_3223,N_3092,N_3152);
and U3224 (N_3224,N_3020,N_3009);
or U3225 (N_3225,N_3173,N_3172);
or U3226 (N_3226,N_3190,N_3118);
nor U3227 (N_3227,N_3035,N_3188);
or U3228 (N_3228,N_3174,N_3108);
or U3229 (N_3229,N_3087,N_3083);
or U3230 (N_3230,N_3183,N_3137);
or U3231 (N_3231,N_3076,N_3094);
or U3232 (N_3232,N_3176,N_3017);
or U3233 (N_3233,N_3151,N_3033);
or U3234 (N_3234,N_3085,N_3132);
nor U3235 (N_3235,N_3052,N_3059);
nand U3236 (N_3236,N_3150,N_3022);
or U3237 (N_3237,N_3110,N_3008);
or U3238 (N_3238,N_3128,N_3078);
nor U3239 (N_3239,N_3170,N_3048);
or U3240 (N_3240,N_3154,N_3148);
nand U3241 (N_3241,N_3036,N_3073);
xnor U3242 (N_3242,N_3032,N_3195);
nor U3243 (N_3243,N_3197,N_3155);
nand U3244 (N_3244,N_3061,N_3138);
nand U3245 (N_3245,N_3004,N_3146);
and U3246 (N_3246,N_3124,N_3050);
and U3247 (N_3247,N_3072,N_3149);
nor U3248 (N_3248,N_3159,N_3106);
xnor U3249 (N_3249,N_3117,N_3095);
or U3250 (N_3250,N_3014,N_3130);
and U3251 (N_3251,N_3165,N_3160);
and U3252 (N_3252,N_3080,N_3185);
and U3253 (N_3253,N_3120,N_3053);
or U3254 (N_3254,N_3126,N_3002);
nand U3255 (N_3255,N_3105,N_3006);
and U3256 (N_3256,N_3003,N_3010);
or U3257 (N_3257,N_3075,N_3016);
nor U3258 (N_3258,N_3025,N_3168);
xnor U3259 (N_3259,N_3074,N_3161);
xor U3260 (N_3260,N_3121,N_3192);
xor U3261 (N_3261,N_3189,N_3063);
or U3262 (N_3262,N_3030,N_3089);
or U3263 (N_3263,N_3096,N_3015);
and U3264 (N_3264,N_3113,N_3090);
or U3265 (N_3265,N_3019,N_3181);
or U3266 (N_3266,N_3147,N_3062);
and U3267 (N_3267,N_3102,N_3111);
nand U3268 (N_3268,N_3060,N_3023);
xnor U3269 (N_3269,N_3057,N_3136);
or U3270 (N_3270,N_3115,N_3182);
nand U3271 (N_3271,N_3167,N_3026);
and U3272 (N_3272,N_3114,N_3191);
nor U3273 (N_3273,N_3031,N_3066);
nor U3274 (N_3274,N_3164,N_3000);
xnor U3275 (N_3275,N_3054,N_3045);
nor U3276 (N_3276,N_3140,N_3071);
or U3277 (N_3277,N_3058,N_3099);
nand U3278 (N_3278,N_3034,N_3029);
xnor U3279 (N_3279,N_3193,N_3007);
or U3280 (N_3280,N_3100,N_3046);
nand U3281 (N_3281,N_3056,N_3042);
nor U3282 (N_3282,N_3051,N_3040);
and U3283 (N_3283,N_3153,N_3021);
or U3284 (N_3284,N_3070,N_3194);
and U3285 (N_3285,N_3163,N_3156);
or U3286 (N_3286,N_3131,N_3077);
nand U3287 (N_3287,N_3186,N_3047);
nand U3288 (N_3288,N_3123,N_3134);
or U3289 (N_3289,N_3065,N_3005);
and U3290 (N_3290,N_3079,N_3018);
nand U3291 (N_3291,N_3069,N_3097);
nand U3292 (N_3292,N_3103,N_3109);
nor U3293 (N_3293,N_3184,N_3143);
nand U3294 (N_3294,N_3116,N_3093);
and U3295 (N_3295,N_3101,N_3086);
nand U3296 (N_3296,N_3127,N_3178);
nand U3297 (N_3297,N_3125,N_3001);
nand U3298 (N_3298,N_3162,N_3166);
nand U3299 (N_3299,N_3098,N_3199);
or U3300 (N_3300,N_3044,N_3186);
nand U3301 (N_3301,N_3145,N_3045);
or U3302 (N_3302,N_3163,N_3114);
and U3303 (N_3303,N_3192,N_3093);
or U3304 (N_3304,N_3092,N_3121);
nand U3305 (N_3305,N_3082,N_3113);
nand U3306 (N_3306,N_3049,N_3023);
nor U3307 (N_3307,N_3089,N_3123);
nand U3308 (N_3308,N_3026,N_3155);
xnor U3309 (N_3309,N_3100,N_3015);
or U3310 (N_3310,N_3103,N_3020);
xor U3311 (N_3311,N_3028,N_3077);
or U3312 (N_3312,N_3187,N_3162);
and U3313 (N_3313,N_3190,N_3073);
xnor U3314 (N_3314,N_3116,N_3163);
nand U3315 (N_3315,N_3106,N_3177);
and U3316 (N_3316,N_3122,N_3065);
or U3317 (N_3317,N_3117,N_3035);
and U3318 (N_3318,N_3149,N_3125);
xor U3319 (N_3319,N_3100,N_3146);
or U3320 (N_3320,N_3182,N_3069);
or U3321 (N_3321,N_3166,N_3170);
nand U3322 (N_3322,N_3071,N_3014);
or U3323 (N_3323,N_3101,N_3122);
nor U3324 (N_3324,N_3018,N_3192);
and U3325 (N_3325,N_3019,N_3143);
and U3326 (N_3326,N_3015,N_3173);
or U3327 (N_3327,N_3026,N_3077);
or U3328 (N_3328,N_3076,N_3006);
or U3329 (N_3329,N_3183,N_3136);
or U3330 (N_3330,N_3008,N_3139);
nand U3331 (N_3331,N_3027,N_3126);
xor U3332 (N_3332,N_3184,N_3064);
and U3333 (N_3333,N_3163,N_3031);
nor U3334 (N_3334,N_3108,N_3119);
or U3335 (N_3335,N_3195,N_3061);
or U3336 (N_3336,N_3030,N_3103);
nor U3337 (N_3337,N_3185,N_3189);
and U3338 (N_3338,N_3092,N_3145);
nand U3339 (N_3339,N_3163,N_3075);
and U3340 (N_3340,N_3096,N_3061);
or U3341 (N_3341,N_3130,N_3062);
and U3342 (N_3342,N_3045,N_3193);
or U3343 (N_3343,N_3128,N_3178);
nand U3344 (N_3344,N_3101,N_3053);
nand U3345 (N_3345,N_3033,N_3177);
nand U3346 (N_3346,N_3155,N_3069);
and U3347 (N_3347,N_3158,N_3063);
and U3348 (N_3348,N_3078,N_3089);
nor U3349 (N_3349,N_3021,N_3067);
nor U3350 (N_3350,N_3127,N_3092);
or U3351 (N_3351,N_3087,N_3137);
nand U3352 (N_3352,N_3070,N_3141);
nand U3353 (N_3353,N_3103,N_3029);
nor U3354 (N_3354,N_3015,N_3045);
or U3355 (N_3355,N_3013,N_3103);
and U3356 (N_3356,N_3130,N_3097);
or U3357 (N_3357,N_3196,N_3106);
nor U3358 (N_3358,N_3069,N_3140);
nor U3359 (N_3359,N_3038,N_3179);
and U3360 (N_3360,N_3026,N_3119);
nor U3361 (N_3361,N_3140,N_3055);
or U3362 (N_3362,N_3014,N_3140);
nor U3363 (N_3363,N_3107,N_3072);
nand U3364 (N_3364,N_3021,N_3096);
and U3365 (N_3365,N_3106,N_3023);
and U3366 (N_3366,N_3166,N_3003);
nor U3367 (N_3367,N_3199,N_3093);
xor U3368 (N_3368,N_3070,N_3197);
or U3369 (N_3369,N_3118,N_3180);
xnor U3370 (N_3370,N_3142,N_3111);
or U3371 (N_3371,N_3007,N_3116);
nor U3372 (N_3372,N_3106,N_3111);
or U3373 (N_3373,N_3108,N_3127);
and U3374 (N_3374,N_3001,N_3167);
or U3375 (N_3375,N_3165,N_3164);
and U3376 (N_3376,N_3135,N_3115);
nor U3377 (N_3377,N_3001,N_3130);
or U3378 (N_3378,N_3048,N_3049);
or U3379 (N_3379,N_3144,N_3081);
or U3380 (N_3380,N_3143,N_3080);
nand U3381 (N_3381,N_3054,N_3107);
nand U3382 (N_3382,N_3189,N_3191);
nor U3383 (N_3383,N_3063,N_3035);
nand U3384 (N_3384,N_3070,N_3166);
nor U3385 (N_3385,N_3058,N_3166);
nand U3386 (N_3386,N_3037,N_3024);
nand U3387 (N_3387,N_3004,N_3038);
nand U3388 (N_3388,N_3012,N_3191);
or U3389 (N_3389,N_3036,N_3050);
nand U3390 (N_3390,N_3114,N_3047);
and U3391 (N_3391,N_3082,N_3039);
nand U3392 (N_3392,N_3067,N_3154);
nand U3393 (N_3393,N_3127,N_3145);
and U3394 (N_3394,N_3173,N_3086);
or U3395 (N_3395,N_3114,N_3027);
nor U3396 (N_3396,N_3176,N_3034);
nand U3397 (N_3397,N_3083,N_3039);
nand U3398 (N_3398,N_3018,N_3139);
nor U3399 (N_3399,N_3179,N_3193);
nand U3400 (N_3400,N_3263,N_3334);
nand U3401 (N_3401,N_3286,N_3270);
or U3402 (N_3402,N_3260,N_3235);
nor U3403 (N_3403,N_3216,N_3243);
or U3404 (N_3404,N_3249,N_3329);
and U3405 (N_3405,N_3330,N_3225);
and U3406 (N_3406,N_3349,N_3383);
and U3407 (N_3407,N_3200,N_3304);
and U3408 (N_3408,N_3255,N_3232);
and U3409 (N_3409,N_3247,N_3390);
nor U3410 (N_3410,N_3236,N_3218);
xor U3411 (N_3411,N_3372,N_3266);
and U3412 (N_3412,N_3296,N_3394);
nor U3413 (N_3413,N_3326,N_3285);
xor U3414 (N_3414,N_3206,N_3250);
xnor U3415 (N_3415,N_3359,N_3233);
nand U3416 (N_3416,N_3272,N_3220);
and U3417 (N_3417,N_3358,N_3389);
and U3418 (N_3418,N_3212,N_3374);
or U3419 (N_3419,N_3340,N_3387);
nand U3420 (N_3420,N_3215,N_3360);
or U3421 (N_3421,N_3343,N_3262);
and U3422 (N_3422,N_3300,N_3397);
or U3423 (N_3423,N_3395,N_3316);
or U3424 (N_3424,N_3254,N_3258);
nor U3425 (N_3425,N_3365,N_3289);
and U3426 (N_3426,N_3347,N_3248);
nand U3427 (N_3427,N_3268,N_3208);
and U3428 (N_3428,N_3345,N_3323);
xor U3429 (N_3429,N_3307,N_3320);
nor U3430 (N_3430,N_3297,N_3338);
or U3431 (N_3431,N_3398,N_3391);
nand U3432 (N_3432,N_3325,N_3219);
or U3433 (N_3433,N_3224,N_3375);
xor U3434 (N_3434,N_3282,N_3382);
and U3435 (N_3435,N_3302,N_3203);
nand U3436 (N_3436,N_3281,N_3336);
nor U3437 (N_3437,N_3246,N_3322);
nand U3438 (N_3438,N_3321,N_3274);
nor U3439 (N_3439,N_3229,N_3284);
nor U3440 (N_3440,N_3367,N_3393);
or U3441 (N_3441,N_3292,N_3324);
and U3442 (N_3442,N_3339,N_3305);
and U3443 (N_3443,N_3279,N_3240);
nand U3444 (N_3444,N_3315,N_3384);
and U3445 (N_3445,N_3295,N_3278);
nor U3446 (N_3446,N_3265,N_3318);
and U3447 (N_3447,N_3399,N_3280);
or U3448 (N_3448,N_3207,N_3337);
nor U3449 (N_3449,N_3314,N_3201);
and U3450 (N_3450,N_3362,N_3332);
nor U3451 (N_3451,N_3237,N_3290);
xor U3452 (N_3452,N_3361,N_3275);
xnor U3453 (N_3453,N_3223,N_3303);
nor U3454 (N_3454,N_3309,N_3256);
and U3455 (N_3455,N_3351,N_3226);
xor U3456 (N_3456,N_3202,N_3344);
and U3457 (N_3457,N_3327,N_3221);
or U3458 (N_3458,N_3346,N_3230);
and U3459 (N_3459,N_3388,N_3308);
nor U3460 (N_3460,N_3228,N_3356);
nand U3461 (N_3461,N_3288,N_3353);
nand U3462 (N_3462,N_3299,N_3306);
and U3463 (N_3463,N_3373,N_3210);
nand U3464 (N_3464,N_3231,N_3317);
and U3465 (N_3465,N_3277,N_3357);
or U3466 (N_3466,N_3385,N_3355);
nand U3467 (N_3467,N_3211,N_3238);
and U3468 (N_3468,N_3205,N_3364);
nand U3469 (N_3469,N_3239,N_3381);
or U3470 (N_3470,N_3287,N_3242);
nand U3471 (N_3471,N_3209,N_3252);
xor U3472 (N_3472,N_3264,N_3386);
nor U3473 (N_3473,N_3392,N_3294);
nor U3474 (N_3474,N_3312,N_3253);
and U3475 (N_3475,N_3380,N_3271);
nor U3476 (N_3476,N_3378,N_3267);
and U3477 (N_3477,N_3227,N_3204);
nand U3478 (N_3478,N_3257,N_3313);
nand U3479 (N_3479,N_3234,N_3310);
nor U3480 (N_3480,N_3222,N_3214);
nor U3481 (N_3481,N_3213,N_3301);
nand U3482 (N_3482,N_3335,N_3244);
nand U3483 (N_3483,N_3283,N_3377);
nand U3484 (N_3484,N_3245,N_3259);
nor U3485 (N_3485,N_3369,N_3396);
xor U3486 (N_3486,N_3291,N_3328);
nor U3487 (N_3487,N_3370,N_3276);
nand U3488 (N_3488,N_3311,N_3342);
and U3489 (N_3489,N_3241,N_3261);
nor U3490 (N_3490,N_3350,N_3293);
nand U3491 (N_3491,N_3368,N_3379);
or U3492 (N_3492,N_3217,N_3352);
or U3493 (N_3493,N_3363,N_3298);
nand U3494 (N_3494,N_3376,N_3354);
or U3495 (N_3495,N_3319,N_3366);
or U3496 (N_3496,N_3371,N_3273);
or U3497 (N_3497,N_3333,N_3251);
and U3498 (N_3498,N_3269,N_3348);
nand U3499 (N_3499,N_3341,N_3331);
nand U3500 (N_3500,N_3376,N_3248);
nor U3501 (N_3501,N_3386,N_3246);
or U3502 (N_3502,N_3224,N_3273);
nor U3503 (N_3503,N_3288,N_3280);
and U3504 (N_3504,N_3248,N_3340);
and U3505 (N_3505,N_3334,N_3206);
or U3506 (N_3506,N_3371,N_3270);
nor U3507 (N_3507,N_3250,N_3288);
nor U3508 (N_3508,N_3357,N_3340);
and U3509 (N_3509,N_3390,N_3367);
nand U3510 (N_3510,N_3377,N_3307);
nor U3511 (N_3511,N_3342,N_3298);
and U3512 (N_3512,N_3327,N_3288);
nor U3513 (N_3513,N_3332,N_3323);
and U3514 (N_3514,N_3255,N_3340);
nand U3515 (N_3515,N_3258,N_3393);
nor U3516 (N_3516,N_3309,N_3239);
and U3517 (N_3517,N_3355,N_3312);
nor U3518 (N_3518,N_3386,N_3252);
or U3519 (N_3519,N_3276,N_3395);
and U3520 (N_3520,N_3335,N_3319);
and U3521 (N_3521,N_3383,N_3382);
nand U3522 (N_3522,N_3212,N_3331);
nor U3523 (N_3523,N_3235,N_3203);
and U3524 (N_3524,N_3272,N_3200);
nand U3525 (N_3525,N_3274,N_3369);
nand U3526 (N_3526,N_3207,N_3398);
or U3527 (N_3527,N_3251,N_3348);
or U3528 (N_3528,N_3240,N_3260);
and U3529 (N_3529,N_3347,N_3210);
nand U3530 (N_3530,N_3223,N_3395);
and U3531 (N_3531,N_3380,N_3314);
nor U3532 (N_3532,N_3379,N_3354);
nand U3533 (N_3533,N_3280,N_3351);
or U3534 (N_3534,N_3388,N_3398);
or U3535 (N_3535,N_3346,N_3396);
and U3536 (N_3536,N_3219,N_3252);
and U3537 (N_3537,N_3360,N_3320);
nand U3538 (N_3538,N_3350,N_3203);
or U3539 (N_3539,N_3261,N_3222);
and U3540 (N_3540,N_3261,N_3232);
nand U3541 (N_3541,N_3343,N_3384);
and U3542 (N_3542,N_3246,N_3217);
or U3543 (N_3543,N_3288,N_3268);
or U3544 (N_3544,N_3249,N_3307);
nor U3545 (N_3545,N_3302,N_3375);
or U3546 (N_3546,N_3215,N_3367);
or U3547 (N_3547,N_3306,N_3354);
or U3548 (N_3548,N_3203,N_3216);
nor U3549 (N_3549,N_3225,N_3237);
or U3550 (N_3550,N_3333,N_3289);
nand U3551 (N_3551,N_3297,N_3342);
and U3552 (N_3552,N_3312,N_3299);
and U3553 (N_3553,N_3308,N_3365);
nand U3554 (N_3554,N_3230,N_3359);
nand U3555 (N_3555,N_3302,N_3365);
nor U3556 (N_3556,N_3219,N_3343);
or U3557 (N_3557,N_3352,N_3347);
or U3558 (N_3558,N_3310,N_3337);
nand U3559 (N_3559,N_3284,N_3331);
and U3560 (N_3560,N_3279,N_3332);
or U3561 (N_3561,N_3374,N_3262);
nor U3562 (N_3562,N_3395,N_3318);
nand U3563 (N_3563,N_3348,N_3203);
or U3564 (N_3564,N_3332,N_3322);
xnor U3565 (N_3565,N_3245,N_3214);
nand U3566 (N_3566,N_3391,N_3295);
xor U3567 (N_3567,N_3205,N_3258);
xor U3568 (N_3568,N_3256,N_3245);
and U3569 (N_3569,N_3234,N_3262);
or U3570 (N_3570,N_3274,N_3295);
nand U3571 (N_3571,N_3209,N_3221);
or U3572 (N_3572,N_3391,N_3229);
nor U3573 (N_3573,N_3209,N_3393);
nand U3574 (N_3574,N_3374,N_3338);
xnor U3575 (N_3575,N_3329,N_3303);
nand U3576 (N_3576,N_3248,N_3229);
nand U3577 (N_3577,N_3271,N_3333);
and U3578 (N_3578,N_3287,N_3231);
or U3579 (N_3579,N_3318,N_3278);
nand U3580 (N_3580,N_3333,N_3203);
and U3581 (N_3581,N_3385,N_3363);
and U3582 (N_3582,N_3295,N_3325);
or U3583 (N_3583,N_3277,N_3332);
nand U3584 (N_3584,N_3305,N_3323);
xor U3585 (N_3585,N_3278,N_3232);
or U3586 (N_3586,N_3240,N_3344);
and U3587 (N_3587,N_3347,N_3259);
nor U3588 (N_3588,N_3270,N_3291);
or U3589 (N_3589,N_3373,N_3275);
nand U3590 (N_3590,N_3347,N_3253);
and U3591 (N_3591,N_3285,N_3308);
nor U3592 (N_3592,N_3281,N_3316);
or U3593 (N_3593,N_3216,N_3328);
nand U3594 (N_3594,N_3240,N_3231);
nand U3595 (N_3595,N_3347,N_3239);
nor U3596 (N_3596,N_3331,N_3278);
nor U3597 (N_3597,N_3376,N_3333);
nor U3598 (N_3598,N_3278,N_3347);
or U3599 (N_3599,N_3252,N_3302);
and U3600 (N_3600,N_3575,N_3581);
nor U3601 (N_3601,N_3458,N_3476);
nor U3602 (N_3602,N_3479,N_3452);
and U3603 (N_3603,N_3570,N_3589);
nor U3604 (N_3604,N_3577,N_3410);
and U3605 (N_3605,N_3511,N_3451);
nand U3606 (N_3606,N_3457,N_3433);
xor U3607 (N_3607,N_3468,N_3502);
and U3608 (N_3608,N_3513,N_3576);
and U3609 (N_3609,N_3426,N_3525);
and U3610 (N_3610,N_3427,N_3447);
xor U3611 (N_3611,N_3488,N_3440);
and U3612 (N_3612,N_3445,N_3551);
xnor U3613 (N_3613,N_3524,N_3541);
nor U3614 (N_3614,N_3503,N_3592);
nor U3615 (N_3615,N_3568,N_3421);
or U3616 (N_3616,N_3569,N_3456);
xor U3617 (N_3617,N_3477,N_3496);
xor U3618 (N_3618,N_3558,N_3429);
and U3619 (N_3619,N_3438,N_3544);
or U3620 (N_3620,N_3556,N_3499);
or U3621 (N_3621,N_3522,N_3453);
or U3622 (N_3622,N_3515,N_3562);
and U3623 (N_3623,N_3563,N_3587);
nor U3624 (N_3624,N_3417,N_3548);
or U3625 (N_3625,N_3439,N_3455);
nand U3626 (N_3626,N_3564,N_3425);
and U3627 (N_3627,N_3595,N_3432);
and U3628 (N_3628,N_3420,N_3549);
nand U3629 (N_3629,N_3516,N_3493);
nor U3630 (N_3630,N_3584,N_3573);
nor U3631 (N_3631,N_3550,N_3597);
or U3632 (N_3632,N_3404,N_3424);
nand U3633 (N_3633,N_3485,N_3521);
nor U3634 (N_3634,N_3506,N_3473);
nand U3635 (N_3635,N_3505,N_3475);
nor U3636 (N_3636,N_3509,N_3474);
nor U3637 (N_3637,N_3465,N_3501);
nand U3638 (N_3638,N_3442,N_3490);
and U3639 (N_3639,N_3532,N_3470);
nor U3640 (N_3640,N_3403,N_3547);
xor U3641 (N_3641,N_3593,N_3553);
or U3642 (N_3642,N_3467,N_3579);
or U3643 (N_3643,N_3406,N_3546);
nor U3644 (N_3644,N_3415,N_3400);
or U3645 (N_3645,N_3443,N_3444);
or U3646 (N_3646,N_3567,N_3537);
nand U3647 (N_3647,N_3431,N_3580);
nand U3648 (N_3648,N_3487,N_3574);
nor U3649 (N_3649,N_3566,N_3519);
and U3650 (N_3650,N_3552,N_3529);
or U3651 (N_3651,N_3586,N_3559);
nor U3652 (N_3652,N_3464,N_3540);
or U3653 (N_3653,N_3560,N_3545);
nand U3654 (N_3654,N_3497,N_3462);
or U3655 (N_3655,N_3459,N_3405);
and U3656 (N_3656,N_3555,N_3454);
and U3657 (N_3657,N_3536,N_3535);
nor U3658 (N_3658,N_3494,N_3507);
nor U3659 (N_3659,N_3542,N_3583);
or U3660 (N_3660,N_3565,N_3423);
nor U3661 (N_3661,N_3437,N_3590);
and U3662 (N_3662,N_3498,N_3594);
nand U3663 (N_3663,N_3460,N_3419);
and U3664 (N_3664,N_3518,N_3411);
and U3665 (N_3665,N_3422,N_3486);
or U3666 (N_3666,N_3534,N_3471);
nand U3667 (N_3667,N_3585,N_3500);
nor U3668 (N_3668,N_3409,N_3517);
and U3669 (N_3669,N_3450,N_3436);
xnor U3670 (N_3670,N_3480,N_3526);
nor U3671 (N_3671,N_3413,N_3401);
xor U3672 (N_3672,N_3483,N_3523);
and U3673 (N_3673,N_3448,N_3441);
nor U3674 (N_3674,N_3588,N_3598);
or U3675 (N_3675,N_3472,N_3512);
nor U3676 (N_3676,N_3402,N_3491);
nand U3677 (N_3677,N_3418,N_3531);
nor U3678 (N_3678,N_3554,N_3481);
nor U3679 (N_3679,N_3414,N_3484);
and U3680 (N_3680,N_3530,N_3538);
nor U3681 (N_3681,N_3407,N_3510);
nor U3682 (N_3682,N_3557,N_3469);
or U3683 (N_3683,N_3520,N_3495);
nand U3684 (N_3684,N_3596,N_3408);
nand U3685 (N_3685,N_3591,N_3514);
nor U3686 (N_3686,N_3482,N_3430);
nand U3687 (N_3687,N_3571,N_3463);
nand U3688 (N_3688,N_3528,N_3466);
or U3689 (N_3689,N_3416,N_3533);
or U3690 (N_3690,N_3446,N_3461);
or U3691 (N_3691,N_3478,N_3561);
nor U3692 (N_3692,N_3434,N_3449);
nand U3693 (N_3693,N_3572,N_3504);
nor U3694 (N_3694,N_3489,N_3412);
and U3695 (N_3695,N_3582,N_3543);
and U3696 (N_3696,N_3428,N_3492);
nand U3697 (N_3697,N_3539,N_3527);
nor U3698 (N_3698,N_3508,N_3599);
or U3699 (N_3699,N_3435,N_3578);
nor U3700 (N_3700,N_3535,N_3561);
nor U3701 (N_3701,N_3577,N_3485);
or U3702 (N_3702,N_3471,N_3428);
nand U3703 (N_3703,N_3411,N_3526);
or U3704 (N_3704,N_3543,N_3547);
nor U3705 (N_3705,N_3521,N_3477);
and U3706 (N_3706,N_3452,N_3430);
nor U3707 (N_3707,N_3471,N_3474);
and U3708 (N_3708,N_3432,N_3597);
and U3709 (N_3709,N_3583,N_3505);
nand U3710 (N_3710,N_3421,N_3459);
and U3711 (N_3711,N_3530,N_3439);
or U3712 (N_3712,N_3414,N_3479);
nor U3713 (N_3713,N_3469,N_3510);
and U3714 (N_3714,N_3460,N_3431);
nor U3715 (N_3715,N_3528,N_3472);
nor U3716 (N_3716,N_3582,N_3492);
nor U3717 (N_3717,N_3539,N_3517);
nor U3718 (N_3718,N_3494,N_3483);
or U3719 (N_3719,N_3576,N_3447);
and U3720 (N_3720,N_3404,N_3488);
xor U3721 (N_3721,N_3515,N_3544);
or U3722 (N_3722,N_3482,N_3503);
nor U3723 (N_3723,N_3421,N_3478);
and U3724 (N_3724,N_3467,N_3439);
and U3725 (N_3725,N_3470,N_3425);
nor U3726 (N_3726,N_3515,N_3530);
xnor U3727 (N_3727,N_3480,N_3570);
and U3728 (N_3728,N_3564,N_3574);
xnor U3729 (N_3729,N_3524,N_3451);
nor U3730 (N_3730,N_3502,N_3438);
xnor U3731 (N_3731,N_3548,N_3426);
xnor U3732 (N_3732,N_3566,N_3539);
and U3733 (N_3733,N_3554,N_3467);
nor U3734 (N_3734,N_3562,N_3480);
nor U3735 (N_3735,N_3554,N_3557);
and U3736 (N_3736,N_3443,N_3463);
nor U3737 (N_3737,N_3599,N_3569);
xor U3738 (N_3738,N_3592,N_3470);
nor U3739 (N_3739,N_3510,N_3493);
xnor U3740 (N_3740,N_3502,N_3441);
xnor U3741 (N_3741,N_3583,N_3452);
nor U3742 (N_3742,N_3574,N_3507);
nor U3743 (N_3743,N_3433,N_3524);
or U3744 (N_3744,N_3540,N_3504);
nand U3745 (N_3745,N_3593,N_3437);
nor U3746 (N_3746,N_3547,N_3536);
nand U3747 (N_3747,N_3408,N_3542);
or U3748 (N_3748,N_3496,N_3417);
nand U3749 (N_3749,N_3443,N_3473);
and U3750 (N_3750,N_3471,N_3445);
and U3751 (N_3751,N_3464,N_3594);
nand U3752 (N_3752,N_3560,N_3555);
and U3753 (N_3753,N_3577,N_3553);
or U3754 (N_3754,N_3567,N_3430);
or U3755 (N_3755,N_3493,N_3468);
and U3756 (N_3756,N_3454,N_3487);
and U3757 (N_3757,N_3574,N_3586);
nor U3758 (N_3758,N_3531,N_3557);
and U3759 (N_3759,N_3474,N_3483);
or U3760 (N_3760,N_3510,N_3441);
nor U3761 (N_3761,N_3512,N_3561);
nand U3762 (N_3762,N_3460,N_3447);
xnor U3763 (N_3763,N_3544,N_3521);
nand U3764 (N_3764,N_3427,N_3437);
or U3765 (N_3765,N_3535,N_3520);
xnor U3766 (N_3766,N_3578,N_3506);
nor U3767 (N_3767,N_3450,N_3563);
and U3768 (N_3768,N_3504,N_3428);
or U3769 (N_3769,N_3509,N_3435);
nor U3770 (N_3770,N_3412,N_3498);
nor U3771 (N_3771,N_3494,N_3593);
nor U3772 (N_3772,N_3572,N_3535);
nand U3773 (N_3773,N_3532,N_3490);
and U3774 (N_3774,N_3561,N_3596);
nor U3775 (N_3775,N_3480,N_3541);
and U3776 (N_3776,N_3450,N_3502);
nor U3777 (N_3777,N_3412,N_3415);
xnor U3778 (N_3778,N_3480,N_3507);
and U3779 (N_3779,N_3507,N_3528);
xor U3780 (N_3780,N_3514,N_3595);
nor U3781 (N_3781,N_3482,N_3457);
and U3782 (N_3782,N_3402,N_3590);
nand U3783 (N_3783,N_3586,N_3439);
and U3784 (N_3784,N_3502,N_3439);
and U3785 (N_3785,N_3547,N_3443);
nor U3786 (N_3786,N_3573,N_3433);
and U3787 (N_3787,N_3498,N_3448);
nor U3788 (N_3788,N_3523,N_3487);
and U3789 (N_3789,N_3554,N_3472);
nor U3790 (N_3790,N_3435,N_3490);
or U3791 (N_3791,N_3407,N_3545);
or U3792 (N_3792,N_3439,N_3492);
xor U3793 (N_3793,N_3567,N_3426);
and U3794 (N_3794,N_3526,N_3455);
and U3795 (N_3795,N_3469,N_3533);
nor U3796 (N_3796,N_3578,N_3426);
or U3797 (N_3797,N_3456,N_3536);
nand U3798 (N_3798,N_3502,N_3410);
or U3799 (N_3799,N_3585,N_3536);
and U3800 (N_3800,N_3680,N_3642);
and U3801 (N_3801,N_3789,N_3754);
nor U3802 (N_3802,N_3648,N_3760);
nor U3803 (N_3803,N_3695,N_3601);
or U3804 (N_3804,N_3765,N_3668);
xnor U3805 (N_3805,N_3704,N_3632);
nand U3806 (N_3806,N_3661,N_3779);
and U3807 (N_3807,N_3604,N_3702);
and U3808 (N_3808,N_3735,N_3607);
nor U3809 (N_3809,N_3685,N_3732);
nand U3810 (N_3810,N_3605,N_3781);
nand U3811 (N_3811,N_3778,N_3651);
nor U3812 (N_3812,N_3753,N_3650);
xor U3813 (N_3813,N_3646,N_3621);
nand U3814 (N_3814,N_3767,N_3701);
xnor U3815 (N_3815,N_3787,N_3707);
xnor U3816 (N_3816,N_3602,N_3688);
nor U3817 (N_3817,N_3622,N_3786);
nand U3818 (N_3818,N_3794,N_3610);
or U3819 (N_3819,N_3676,N_3798);
nor U3820 (N_3820,N_3666,N_3795);
nor U3821 (N_3821,N_3758,N_3733);
nand U3822 (N_3822,N_3641,N_3609);
nand U3823 (N_3823,N_3647,N_3736);
nand U3824 (N_3824,N_3717,N_3679);
and U3825 (N_3825,N_3708,N_3645);
nor U3826 (N_3826,N_3768,N_3674);
xor U3827 (N_3827,N_3759,N_3771);
or U3828 (N_3828,N_3729,N_3724);
nor U3829 (N_3829,N_3722,N_3744);
xnor U3830 (N_3830,N_3718,N_3792);
or U3831 (N_3831,N_3640,N_3669);
and U3832 (N_3832,N_3615,N_3629);
nor U3833 (N_3833,N_3713,N_3745);
nor U3834 (N_3834,N_3697,N_3743);
or U3835 (N_3835,N_3712,N_3737);
and U3836 (N_3836,N_3705,N_3617);
nand U3837 (N_3837,N_3700,N_3776);
and U3838 (N_3838,N_3716,N_3793);
nand U3839 (N_3839,N_3630,N_3748);
nor U3840 (N_3840,N_3764,N_3738);
nor U3841 (N_3841,N_3723,N_3638);
nand U3842 (N_3842,N_3611,N_3761);
or U3843 (N_3843,N_3710,N_3655);
nor U3844 (N_3844,N_3775,N_3720);
or U3845 (N_3845,N_3785,N_3739);
nor U3846 (N_3846,N_3692,N_3659);
nand U3847 (N_3847,N_3687,N_3624);
or U3848 (N_3848,N_3639,N_3725);
or U3849 (N_3849,N_3690,N_3634);
or U3850 (N_3850,N_3734,N_3750);
and U3851 (N_3851,N_3719,N_3625);
nor U3852 (N_3852,N_3780,N_3791);
xor U3853 (N_3853,N_3603,N_3667);
nor U3854 (N_3854,N_3671,N_3726);
and U3855 (N_3855,N_3762,N_3756);
nand U3856 (N_3856,N_3746,N_3612);
or U3857 (N_3857,N_3777,N_3799);
and U3858 (N_3858,N_3633,N_3656);
and U3859 (N_3859,N_3763,N_3643);
or U3860 (N_3860,N_3618,N_3681);
nand U3861 (N_3861,N_3749,N_3673);
xnor U3862 (N_3862,N_3698,N_3711);
or U3863 (N_3863,N_3628,N_3714);
nand U3864 (N_3864,N_3677,N_3784);
and U3865 (N_3865,N_3689,N_3727);
nand U3866 (N_3866,N_3626,N_3675);
nand U3867 (N_3867,N_3684,N_3652);
nor U3868 (N_3868,N_3686,N_3709);
nor U3869 (N_3869,N_3703,N_3730);
nand U3870 (N_3870,N_3658,N_3616);
and U3871 (N_3871,N_3678,N_3664);
nor U3872 (N_3872,N_3608,N_3774);
nand U3873 (N_3873,N_3747,N_3751);
nor U3874 (N_3874,N_3757,N_3788);
or U3875 (N_3875,N_3670,N_3654);
nor U3876 (N_3876,N_3783,N_3635);
and U3877 (N_3877,N_3797,N_3790);
and U3878 (N_3878,N_3663,N_3614);
xor U3879 (N_3879,N_3721,N_3644);
and U3880 (N_3880,N_3715,N_3660);
and U3881 (N_3881,N_3752,N_3619);
nor U3882 (N_3882,N_3620,N_3796);
or U3883 (N_3883,N_3631,N_3662);
nor U3884 (N_3884,N_3740,N_3699);
nor U3885 (N_3885,N_3766,N_3731);
and U3886 (N_3886,N_3623,N_3636);
and U3887 (N_3887,N_3782,N_3728);
xor U3888 (N_3888,N_3741,N_3769);
xor U3889 (N_3889,N_3696,N_3665);
or U3890 (N_3890,N_3627,N_3613);
xnor U3891 (N_3891,N_3606,N_3706);
and U3892 (N_3892,N_3773,N_3742);
or U3893 (N_3893,N_3755,N_3770);
nand U3894 (N_3894,N_3649,N_3637);
nand U3895 (N_3895,N_3691,N_3657);
and U3896 (N_3896,N_3653,N_3694);
xor U3897 (N_3897,N_3772,N_3682);
and U3898 (N_3898,N_3693,N_3672);
and U3899 (N_3899,N_3600,N_3683);
nor U3900 (N_3900,N_3671,N_3612);
or U3901 (N_3901,N_3694,N_3779);
or U3902 (N_3902,N_3788,N_3767);
or U3903 (N_3903,N_3730,N_3791);
xnor U3904 (N_3904,N_3619,N_3651);
and U3905 (N_3905,N_3657,N_3791);
or U3906 (N_3906,N_3638,N_3649);
nor U3907 (N_3907,N_3635,N_3786);
xnor U3908 (N_3908,N_3608,N_3642);
nand U3909 (N_3909,N_3733,N_3660);
xor U3910 (N_3910,N_3789,N_3694);
nand U3911 (N_3911,N_3739,N_3658);
and U3912 (N_3912,N_3663,N_3795);
or U3913 (N_3913,N_3645,N_3613);
nor U3914 (N_3914,N_3618,N_3793);
or U3915 (N_3915,N_3617,N_3713);
nand U3916 (N_3916,N_3630,N_3758);
nor U3917 (N_3917,N_3628,N_3635);
and U3918 (N_3918,N_3676,N_3610);
nor U3919 (N_3919,N_3759,N_3651);
nand U3920 (N_3920,N_3643,N_3634);
or U3921 (N_3921,N_3612,N_3662);
xnor U3922 (N_3922,N_3700,N_3630);
or U3923 (N_3923,N_3694,N_3732);
or U3924 (N_3924,N_3607,N_3631);
and U3925 (N_3925,N_3762,N_3783);
nor U3926 (N_3926,N_3633,N_3653);
nand U3927 (N_3927,N_3666,N_3610);
and U3928 (N_3928,N_3686,N_3666);
nand U3929 (N_3929,N_3640,N_3742);
nor U3930 (N_3930,N_3667,N_3709);
or U3931 (N_3931,N_3774,N_3794);
and U3932 (N_3932,N_3774,N_3700);
and U3933 (N_3933,N_3705,N_3713);
nor U3934 (N_3934,N_3745,N_3775);
xnor U3935 (N_3935,N_3713,N_3653);
nor U3936 (N_3936,N_3767,N_3773);
nor U3937 (N_3937,N_3717,N_3619);
nor U3938 (N_3938,N_3633,N_3764);
nor U3939 (N_3939,N_3646,N_3795);
or U3940 (N_3940,N_3758,N_3737);
nor U3941 (N_3941,N_3758,N_3654);
or U3942 (N_3942,N_3649,N_3766);
nand U3943 (N_3943,N_3616,N_3610);
nor U3944 (N_3944,N_3629,N_3670);
xor U3945 (N_3945,N_3639,N_3663);
nand U3946 (N_3946,N_3713,N_3645);
xor U3947 (N_3947,N_3628,N_3736);
xor U3948 (N_3948,N_3794,N_3629);
nor U3949 (N_3949,N_3755,N_3691);
nand U3950 (N_3950,N_3689,N_3688);
nor U3951 (N_3951,N_3797,N_3622);
and U3952 (N_3952,N_3613,N_3781);
xor U3953 (N_3953,N_3661,N_3733);
xor U3954 (N_3954,N_3748,N_3612);
nand U3955 (N_3955,N_3705,N_3673);
xor U3956 (N_3956,N_3715,N_3672);
and U3957 (N_3957,N_3750,N_3675);
or U3958 (N_3958,N_3757,N_3616);
or U3959 (N_3959,N_3604,N_3644);
nor U3960 (N_3960,N_3698,N_3625);
or U3961 (N_3961,N_3718,N_3714);
and U3962 (N_3962,N_3717,N_3608);
or U3963 (N_3963,N_3608,N_3790);
nor U3964 (N_3964,N_3758,N_3651);
nor U3965 (N_3965,N_3768,N_3777);
nor U3966 (N_3966,N_3670,N_3706);
nor U3967 (N_3967,N_3793,N_3744);
or U3968 (N_3968,N_3714,N_3694);
and U3969 (N_3969,N_3678,N_3626);
and U3970 (N_3970,N_3632,N_3641);
nor U3971 (N_3971,N_3687,N_3768);
and U3972 (N_3972,N_3721,N_3729);
nor U3973 (N_3973,N_3637,N_3770);
xor U3974 (N_3974,N_3747,N_3682);
and U3975 (N_3975,N_3664,N_3721);
nand U3976 (N_3976,N_3765,N_3711);
nand U3977 (N_3977,N_3670,N_3691);
nor U3978 (N_3978,N_3615,N_3674);
and U3979 (N_3979,N_3754,N_3755);
nand U3980 (N_3980,N_3765,N_3676);
or U3981 (N_3981,N_3734,N_3634);
nand U3982 (N_3982,N_3794,N_3630);
or U3983 (N_3983,N_3719,N_3692);
nor U3984 (N_3984,N_3781,N_3706);
or U3985 (N_3985,N_3762,N_3633);
or U3986 (N_3986,N_3763,N_3682);
nor U3987 (N_3987,N_3626,N_3724);
nor U3988 (N_3988,N_3786,N_3746);
or U3989 (N_3989,N_3743,N_3757);
or U3990 (N_3990,N_3709,N_3769);
nand U3991 (N_3991,N_3710,N_3731);
and U3992 (N_3992,N_3727,N_3657);
or U3993 (N_3993,N_3709,N_3644);
xnor U3994 (N_3994,N_3610,N_3609);
and U3995 (N_3995,N_3705,N_3613);
nor U3996 (N_3996,N_3777,N_3626);
and U3997 (N_3997,N_3753,N_3668);
and U3998 (N_3998,N_3733,N_3669);
or U3999 (N_3999,N_3785,N_3775);
xnor U4000 (N_4000,N_3834,N_3836);
nand U4001 (N_4001,N_3897,N_3964);
xor U4002 (N_4002,N_3858,N_3869);
and U4003 (N_4003,N_3935,N_3984);
nor U4004 (N_4004,N_3925,N_3977);
nand U4005 (N_4005,N_3878,N_3982);
xnor U4006 (N_4006,N_3845,N_3955);
nor U4007 (N_4007,N_3995,N_3906);
nand U4008 (N_4008,N_3861,N_3874);
nand U4009 (N_4009,N_3885,N_3952);
nor U4010 (N_4010,N_3993,N_3875);
or U4011 (N_4011,N_3828,N_3939);
nor U4012 (N_4012,N_3960,N_3871);
nor U4013 (N_4013,N_3890,N_3928);
nand U4014 (N_4014,N_3857,N_3903);
or U4015 (N_4015,N_3868,N_3812);
xnor U4016 (N_4016,N_3817,N_3986);
nor U4017 (N_4017,N_3829,N_3837);
or U4018 (N_4018,N_3902,N_3978);
nand U4019 (N_4019,N_3989,N_3922);
or U4020 (N_4020,N_3990,N_3908);
or U4021 (N_4021,N_3973,N_3974);
and U4022 (N_4022,N_3942,N_3840);
nor U4023 (N_4023,N_3929,N_3991);
nand U4024 (N_4024,N_3946,N_3898);
nand U4025 (N_4025,N_3849,N_3850);
or U4026 (N_4026,N_3801,N_3880);
nor U4027 (N_4027,N_3924,N_3821);
nand U4028 (N_4028,N_3888,N_3971);
xor U4029 (N_4029,N_3950,N_3913);
nand U4030 (N_4030,N_3987,N_3949);
nand U4031 (N_4031,N_3820,N_3816);
and U4032 (N_4032,N_3985,N_3814);
nand U4033 (N_4033,N_3915,N_3919);
or U4034 (N_4034,N_3934,N_3892);
nand U4035 (N_4035,N_3920,N_3948);
and U4036 (N_4036,N_3976,N_3853);
nor U4037 (N_4037,N_3847,N_3833);
and U4038 (N_4038,N_3962,N_3972);
nand U4039 (N_4039,N_3916,N_3927);
nand U4040 (N_4040,N_3956,N_3894);
nand U4041 (N_4041,N_3852,N_3863);
or U4042 (N_4042,N_3824,N_3806);
or U4043 (N_4043,N_3822,N_3872);
nand U4044 (N_4044,N_3926,N_3909);
or U4045 (N_4045,N_3802,N_3803);
nor U4046 (N_4046,N_3979,N_3825);
xor U4047 (N_4047,N_3889,N_3873);
or U4048 (N_4048,N_3970,N_3883);
or U4049 (N_4049,N_3996,N_3804);
nor U4050 (N_4050,N_3967,N_3818);
or U4051 (N_4051,N_3882,N_3865);
xor U4052 (N_4052,N_3937,N_3941);
nand U4053 (N_4053,N_3963,N_3831);
nor U4054 (N_4054,N_3887,N_3879);
nand U4055 (N_4055,N_3921,N_3881);
xnor U4056 (N_4056,N_3969,N_3914);
and U4057 (N_4057,N_3954,N_3811);
xor U4058 (N_4058,N_3999,N_3862);
nand U4059 (N_4059,N_3848,N_3827);
and U4060 (N_4060,N_3877,N_3912);
and U4061 (N_4061,N_3936,N_3917);
nor U4062 (N_4062,N_3886,N_3805);
xor U4063 (N_4063,N_3800,N_3867);
or U4064 (N_4064,N_3933,N_3980);
and U4065 (N_4065,N_3876,N_3893);
and U4066 (N_4066,N_3823,N_3860);
xnor U4067 (N_4067,N_3815,N_3866);
nand U4068 (N_4068,N_3911,N_3901);
and U4069 (N_4069,N_3951,N_3968);
xnor U4070 (N_4070,N_3992,N_3846);
nand U4071 (N_4071,N_3830,N_3870);
and U4072 (N_4072,N_3958,N_3988);
nor U4073 (N_4073,N_3899,N_3841);
nor U4074 (N_4074,N_3819,N_3943);
nor U4075 (N_4075,N_3932,N_3947);
nor U4076 (N_4076,N_3983,N_3851);
xnor U4077 (N_4077,N_3809,N_3854);
nor U4078 (N_4078,N_3938,N_3905);
and U4079 (N_4079,N_3891,N_3810);
xnor U4080 (N_4080,N_3856,N_3896);
nor U4081 (N_4081,N_3864,N_3855);
or U4082 (N_4082,N_3807,N_3923);
and U4083 (N_4083,N_3994,N_3931);
nand U4084 (N_4084,N_3843,N_3940);
or U4085 (N_4085,N_3838,N_3957);
xor U4086 (N_4086,N_3918,N_3998);
nand U4087 (N_4087,N_3966,N_3835);
nor U4088 (N_4088,N_3832,N_3965);
xnor U4089 (N_4089,N_3930,N_3910);
nand U4090 (N_4090,N_3959,N_3844);
or U4091 (N_4091,N_3945,N_3944);
and U4092 (N_4092,N_3842,N_3859);
nand U4093 (N_4093,N_3904,N_3826);
nor U4094 (N_4094,N_3839,N_3975);
nor U4095 (N_4095,N_3961,N_3997);
nand U4096 (N_4096,N_3981,N_3895);
or U4097 (N_4097,N_3813,N_3907);
nor U4098 (N_4098,N_3808,N_3900);
or U4099 (N_4099,N_3953,N_3884);
nor U4100 (N_4100,N_3986,N_3837);
nand U4101 (N_4101,N_3901,N_3865);
nand U4102 (N_4102,N_3901,N_3906);
nand U4103 (N_4103,N_3873,N_3832);
and U4104 (N_4104,N_3925,N_3885);
xnor U4105 (N_4105,N_3971,N_3858);
nor U4106 (N_4106,N_3969,N_3940);
and U4107 (N_4107,N_3962,N_3974);
or U4108 (N_4108,N_3824,N_3837);
nand U4109 (N_4109,N_3946,N_3900);
nor U4110 (N_4110,N_3898,N_3848);
and U4111 (N_4111,N_3916,N_3914);
nor U4112 (N_4112,N_3997,N_3905);
nor U4113 (N_4113,N_3868,N_3808);
and U4114 (N_4114,N_3858,N_3988);
nor U4115 (N_4115,N_3823,N_3976);
nor U4116 (N_4116,N_3942,N_3825);
or U4117 (N_4117,N_3883,N_3905);
nand U4118 (N_4118,N_3940,N_3881);
nor U4119 (N_4119,N_3861,N_3934);
xor U4120 (N_4120,N_3918,N_3870);
or U4121 (N_4121,N_3871,N_3837);
and U4122 (N_4122,N_3874,N_3803);
nand U4123 (N_4123,N_3806,N_3940);
xor U4124 (N_4124,N_3959,N_3926);
nor U4125 (N_4125,N_3819,N_3935);
xor U4126 (N_4126,N_3950,N_3850);
or U4127 (N_4127,N_3985,N_3902);
nand U4128 (N_4128,N_3871,N_3844);
or U4129 (N_4129,N_3942,N_3802);
nand U4130 (N_4130,N_3934,N_3974);
or U4131 (N_4131,N_3852,N_3905);
nand U4132 (N_4132,N_3874,N_3870);
and U4133 (N_4133,N_3922,N_3840);
nand U4134 (N_4134,N_3825,N_3863);
nand U4135 (N_4135,N_3860,N_3838);
or U4136 (N_4136,N_3861,N_3966);
nand U4137 (N_4137,N_3889,N_3893);
and U4138 (N_4138,N_3812,N_3807);
nand U4139 (N_4139,N_3990,N_3950);
nor U4140 (N_4140,N_3928,N_3827);
and U4141 (N_4141,N_3873,N_3939);
or U4142 (N_4142,N_3950,N_3826);
or U4143 (N_4143,N_3989,N_3982);
xor U4144 (N_4144,N_3947,N_3890);
nand U4145 (N_4145,N_3906,N_3949);
or U4146 (N_4146,N_3915,N_3852);
xnor U4147 (N_4147,N_3871,N_3895);
and U4148 (N_4148,N_3825,N_3943);
nand U4149 (N_4149,N_3925,N_3800);
and U4150 (N_4150,N_3845,N_3931);
nand U4151 (N_4151,N_3921,N_3843);
and U4152 (N_4152,N_3980,N_3976);
or U4153 (N_4153,N_3872,N_3936);
nand U4154 (N_4154,N_3924,N_3959);
nand U4155 (N_4155,N_3889,N_3860);
or U4156 (N_4156,N_3896,N_3933);
and U4157 (N_4157,N_3835,N_3857);
and U4158 (N_4158,N_3903,N_3812);
xnor U4159 (N_4159,N_3992,N_3897);
nand U4160 (N_4160,N_3847,N_3848);
nand U4161 (N_4161,N_3831,N_3903);
nand U4162 (N_4162,N_3903,N_3908);
nor U4163 (N_4163,N_3803,N_3845);
nand U4164 (N_4164,N_3809,N_3911);
and U4165 (N_4165,N_3862,N_3847);
and U4166 (N_4166,N_3907,N_3854);
and U4167 (N_4167,N_3830,N_3842);
and U4168 (N_4168,N_3951,N_3837);
nand U4169 (N_4169,N_3945,N_3864);
and U4170 (N_4170,N_3900,N_3856);
nand U4171 (N_4171,N_3922,N_3910);
nor U4172 (N_4172,N_3899,N_3923);
nand U4173 (N_4173,N_3888,N_3893);
nor U4174 (N_4174,N_3980,N_3962);
nor U4175 (N_4175,N_3986,N_3857);
nor U4176 (N_4176,N_3981,N_3908);
and U4177 (N_4177,N_3972,N_3850);
nand U4178 (N_4178,N_3844,N_3881);
nor U4179 (N_4179,N_3954,N_3929);
nand U4180 (N_4180,N_3978,N_3822);
and U4181 (N_4181,N_3849,N_3822);
or U4182 (N_4182,N_3895,N_3928);
or U4183 (N_4183,N_3836,N_3979);
or U4184 (N_4184,N_3940,N_3902);
nor U4185 (N_4185,N_3994,N_3962);
nor U4186 (N_4186,N_3870,N_3814);
nand U4187 (N_4187,N_3947,N_3877);
and U4188 (N_4188,N_3921,N_3824);
nor U4189 (N_4189,N_3876,N_3844);
nor U4190 (N_4190,N_3826,N_3967);
or U4191 (N_4191,N_3931,N_3992);
or U4192 (N_4192,N_3947,N_3892);
xnor U4193 (N_4193,N_3908,N_3920);
nand U4194 (N_4194,N_3952,N_3886);
nand U4195 (N_4195,N_3980,N_3866);
nand U4196 (N_4196,N_3968,N_3894);
and U4197 (N_4197,N_3978,N_3891);
nand U4198 (N_4198,N_3873,N_3934);
nor U4199 (N_4199,N_3916,N_3820);
nor U4200 (N_4200,N_4082,N_4007);
nand U4201 (N_4201,N_4088,N_4175);
and U4202 (N_4202,N_4026,N_4051);
and U4203 (N_4203,N_4163,N_4176);
and U4204 (N_4204,N_4152,N_4103);
xnor U4205 (N_4205,N_4135,N_4105);
and U4206 (N_4206,N_4153,N_4092);
nand U4207 (N_4207,N_4029,N_4036);
or U4208 (N_4208,N_4009,N_4011);
and U4209 (N_4209,N_4001,N_4083);
nand U4210 (N_4210,N_4032,N_4014);
or U4211 (N_4211,N_4020,N_4139);
xor U4212 (N_4212,N_4086,N_4003);
nand U4213 (N_4213,N_4084,N_4146);
nand U4214 (N_4214,N_4025,N_4089);
or U4215 (N_4215,N_4165,N_4129);
nor U4216 (N_4216,N_4170,N_4112);
xor U4217 (N_4217,N_4070,N_4085);
and U4218 (N_4218,N_4069,N_4142);
and U4219 (N_4219,N_4006,N_4094);
nor U4220 (N_4220,N_4137,N_4110);
nor U4221 (N_4221,N_4181,N_4055);
or U4222 (N_4222,N_4192,N_4038);
xnor U4223 (N_4223,N_4047,N_4194);
xor U4224 (N_4224,N_4171,N_4193);
or U4225 (N_4225,N_4002,N_4156);
nor U4226 (N_4226,N_4018,N_4075);
nor U4227 (N_4227,N_4143,N_4034);
and U4228 (N_4228,N_4107,N_4123);
and U4229 (N_4229,N_4106,N_4056);
and U4230 (N_4230,N_4172,N_4118);
nor U4231 (N_4231,N_4044,N_4049);
nor U4232 (N_4232,N_4008,N_4066);
nand U4233 (N_4233,N_4187,N_4100);
nand U4234 (N_4234,N_4188,N_4179);
nor U4235 (N_4235,N_4013,N_4154);
xor U4236 (N_4236,N_4189,N_4131);
or U4237 (N_4237,N_4198,N_4136);
nor U4238 (N_4238,N_4126,N_4149);
nand U4239 (N_4239,N_4037,N_4168);
nand U4240 (N_4240,N_4097,N_4199);
nand U4241 (N_4241,N_4160,N_4071);
or U4242 (N_4242,N_4119,N_4030);
nand U4243 (N_4243,N_4046,N_4060);
or U4244 (N_4244,N_4093,N_4130);
or U4245 (N_4245,N_4185,N_4021);
nand U4246 (N_4246,N_4104,N_4158);
and U4247 (N_4247,N_4074,N_4050);
nor U4248 (N_4248,N_4042,N_4108);
nor U4249 (N_4249,N_4040,N_4076);
nor U4250 (N_4250,N_4035,N_4031);
nand U4251 (N_4251,N_4010,N_4043);
nand U4252 (N_4252,N_4077,N_4081);
and U4253 (N_4253,N_4064,N_4065);
or U4254 (N_4254,N_4195,N_4197);
nor U4255 (N_4255,N_4079,N_4059);
nor U4256 (N_4256,N_4080,N_4161);
nand U4257 (N_4257,N_4147,N_4072);
or U4258 (N_4258,N_4053,N_4145);
nand U4259 (N_4259,N_4028,N_4144);
or U4260 (N_4260,N_4023,N_4190);
or U4261 (N_4261,N_4057,N_4166);
nand U4262 (N_4262,N_4178,N_4151);
xor U4263 (N_4263,N_4015,N_4016);
and U4264 (N_4264,N_4113,N_4196);
nor U4265 (N_4265,N_4102,N_4150);
or U4266 (N_4266,N_4121,N_4090);
nand U4267 (N_4267,N_4027,N_4164);
and U4268 (N_4268,N_4098,N_4048);
and U4269 (N_4269,N_4141,N_4067);
or U4270 (N_4270,N_4012,N_4062);
or U4271 (N_4271,N_4033,N_4122);
xnor U4272 (N_4272,N_4138,N_4114);
and U4273 (N_4273,N_4058,N_4128);
nand U4274 (N_4274,N_4182,N_4183);
or U4275 (N_4275,N_4157,N_4017);
or U4276 (N_4276,N_4120,N_4155);
nand U4277 (N_4277,N_4177,N_4101);
nand U4278 (N_4278,N_4022,N_4125);
nand U4279 (N_4279,N_4186,N_4095);
nor U4280 (N_4280,N_4162,N_4045);
or U4281 (N_4281,N_4159,N_4180);
xor U4282 (N_4282,N_4039,N_4087);
nor U4283 (N_4283,N_4054,N_4140);
nor U4284 (N_4284,N_4109,N_4174);
nand U4285 (N_4285,N_4061,N_4091);
and U4286 (N_4286,N_4005,N_4063);
nand U4287 (N_4287,N_4169,N_4000);
and U4288 (N_4288,N_4052,N_4115);
or U4289 (N_4289,N_4132,N_4184);
nand U4290 (N_4290,N_4019,N_4134);
and U4291 (N_4291,N_4073,N_4191);
and U4292 (N_4292,N_4111,N_4117);
and U4293 (N_4293,N_4099,N_4078);
or U4294 (N_4294,N_4096,N_4004);
and U4295 (N_4295,N_4148,N_4116);
and U4296 (N_4296,N_4024,N_4167);
xnor U4297 (N_4297,N_4068,N_4133);
nand U4298 (N_4298,N_4173,N_4041);
xnor U4299 (N_4299,N_4124,N_4127);
nand U4300 (N_4300,N_4013,N_4047);
or U4301 (N_4301,N_4100,N_4082);
nand U4302 (N_4302,N_4163,N_4071);
xor U4303 (N_4303,N_4196,N_4195);
and U4304 (N_4304,N_4000,N_4165);
nand U4305 (N_4305,N_4091,N_4174);
nor U4306 (N_4306,N_4020,N_4123);
nor U4307 (N_4307,N_4051,N_4121);
nand U4308 (N_4308,N_4159,N_4109);
nor U4309 (N_4309,N_4162,N_4149);
nor U4310 (N_4310,N_4091,N_4196);
nand U4311 (N_4311,N_4106,N_4034);
or U4312 (N_4312,N_4022,N_4165);
or U4313 (N_4313,N_4173,N_4120);
or U4314 (N_4314,N_4120,N_4119);
nor U4315 (N_4315,N_4006,N_4021);
or U4316 (N_4316,N_4051,N_4060);
or U4317 (N_4317,N_4120,N_4182);
nand U4318 (N_4318,N_4111,N_4011);
and U4319 (N_4319,N_4147,N_4190);
or U4320 (N_4320,N_4118,N_4006);
or U4321 (N_4321,N_4161,N_4024);
nand U4322 (N_4322,N_4004,N_4064);
nor U4323 (N_4323,N_4049,N_4109);
or U4324 (N_4324,N_4049,N_4178);
or U4325 (N_4325,N_4192,N_4118);
nor U4326 (N_4326,N_4102,N_4094);
nor U4327 (N_4327,N_4134,N_4003);
nor U4328 (N_4328,N_4172,N_4186);
xor U4329 (N_4329,N_4121,N_4021);
xor U4330 (N_4330,N_4091,N_4025);
and U4331 (N_4331,N_4015,N_4048);
or U4332 (N_4332,N_4023,N_4167);
nand U4333 (N_4333,N_4118,N_4082);
xor U4334 (N_4334,N_4075,N_4031);
nor U4335 (N_4335,N_4104,N_4199);
or U4336 (N_4336,N_4050,N_4199);
xor U4337 (N_4337,N_4131,N_4176);
nand U4338 (N_4338,N_4057,N_4157);
nor U4339 (N_4339,N_4000,N_4121);
and U4340 (N_4340,N_4067,N_4053);
and U4341 (N_4341,N_4128,N_4192);
xor U4342 (N_4342,N_4000,N_4012);
nand U4343 (N_4343,N_4032,N_4082);
xnor U4344 (N_4344,N_4156,N_4114);
nor U4345 (N_4345,N_4035,N_4097);
xnor U4346 (N_4346,N_4171,N_4152);
nor U4347 (N_4347,N_4007,N_4019);
and U4348 (N_4348,N_4020,N_4162);
nand U4349 (N_4349,N_4196,N_4146);
nor U4350 (N_4350,N_4070,N_4088);
and U4351 (N_4351,N_4140,N_4083);
and U4352 (N_4352,N_4012,N_4158);
and U4353 (N_4353,N_4075,N_4061);
nor U4354 (N_4354,N_4004,N_4147);
or U4355 (N_4355,N_4121,N_4043);
nand U4356 (N_4356,N_4156,N_4020);
nor U4357 (N_4357,N_4029,N_4016);
nand U4358 (N_4358,N_4074,N_4126);
nand U4359 (N_4359,N_4052,N_4136);
nor U4360 (N_4360,N_4045,N_4168);
or U4361 (N_4361,N_4147,N_4069);
nand U4362 (N_4362,N_4115,N_4110);
nor U4363 (N_4363,N_4188,N_4013);
or U4364 (N_4364,N_4106,N_4030);
xor U4365 (N_4365,N_4191,N_4068);
nor U4366 (N_4366,N_4180,N_4085);
nand U4367 (N_4367,N_4005,N_4187);
nor U4368 (N_4368,N_4020,N_4060);
nor U4369 (N_4369,N_4018,N_4007);
nand U4370 (N_4370,N_4107,N_4183);
or U4371 (N_4371,N_4090,N_4032);
nor U4372 (N_4372,N_4180,N_4170);
xor U4373 (N_4373,N_4101,N_4175);
nor U4374 (N_4374,N_4037,N_4012);
or U4375 (N_4375,N_4078,N_4113);
xor U4376 (N_4376,N_4097,N_4037);
nor U4377 (N_4377,N_4081,N_4159);
nand U4378 (N_4378,N_4016,N_4073);
nor U4379 (N_4379,N_4074,N_4136);
nand U4380 (N_4380,N_4172,N_4078);
nand U4381 (N_4381,N_4194,N_4065);
nor U4382 (N_4382,N_4056,N_4101);
xor U4383 (N_4383,N_4008,N_4190);
or U4384 (N_4384,N_4086,N_4030);
nand U4385 (N_4385,N_4146,N_4190);
and U4386 (N_4386,N_4132,N_4034);
nor U4387 (N_4387,N_4157,N_4115);
or U4388 (N_4388,N_4125,N_4143);
nor U4389 (N_4389,N_4103,N_4198);
nor U4390 (N_4390,N_4198,N_4171);
and U4391 (N_4391,N_4072,N_4146);
and U4392 (N_4392,N_4065,N_4102);
and U4393 (N_4393,N_4139,N_4157);
or U4394 (N_4394,N_4104,N_4112);
nor U4395 (N_4395,N_4012,N_4128);
and U4396 (N_4396,N_4110,N_4192);
nand U4397 (N_4397,N_4085,N_4122);
xor U4398 (N_4398,N_4166,N_4001);
and U4399 (N_4399,N_4123,N_4135);
or U4400 (N_4400,N_4208,N_4206);
and U4401 (N_4401,N_4288,N_4399);
or U4402 (N_4402,N_4310,N_4397);
or U4403 (N_4403,N_4358,N_4285);
and U4404 (N_4404,N_4214,N_4238);
and U4405 (N_4405,N_4356,N_4220);
and U4406 (N_4406,N_4205,N_4241);
nor U4407 (N_4407,N_4260,N_4377);
nor U4408 (N_4408,N_4343,N_4366);
nand U4409 (N_4409,N_4231,N_4264);
nor U4410 (N_4410,N_4262,N_4216);
and U4411 (N_4411,N_4368,N_4298);
or U4412 (N_4412,N_4332,N_4270);
and U4413 (N_4413,N_4211,N_4280);
or U4414 (N_4414,N_4226,N_4396);
nor U4415 (N_4415,N_4307,N_4318);
and U4416 (N_4416,N_4225,N_4251);
and U4417 (N_4417,N_4393,N_4229);
nor U4418 (N_4418,N_4242,N_4248);
and U4419 (N_4419,N_4323,N_4247);
or U4420 (N_4420,N_4266,N_4376);
xnor U4421 (N_4421,N_4304,N_4256);
or U4422 (N_4422,N_4339,N_4255);
nor U4423 (N_4423,N_4379,N_4244);
and U4424 (N_4424,N_4201,N_4227);
and U4425 (N_4425,N_4233,N_4268);
xor U4426 (N_4426,N_4375,N_4367);
nand U4427 (N_4427,N_4346,N_4301);
nor U4428 (N_4428,N_4328,N_4364);
and U4429 (N_4429,N_4232,N_4378);
or U4430 (N_4430,N_4355,N_4352);
xnor U4431 (N_4431,N_4273,N_4371);
nor U4432 (N_4432,N_4240,N_4385);
or U4433 (N_4433,N_4363,N_4391);
and U4434 (N_4434,N_4327,N_4223);
nand U4435 (N_4435,N_4258,N_4299);
or U4436 (N_4436,N_4249,N_4274);
nand U4437 (N_4437,N_4284,N_4372);
or U4438 (N_4438,N_4338,N_4265);
nor U4439 (N_4439,N_4263,N_4315);
nand U4440 (N_4440,N_4336,N_4321);
nand U4441 (N_4441,N_4259,N_4219);
and U4442 (N_4442,N_4362,N_4294);
nor U4443 (N_4443,N_4330,N_4390);
or U4444 (N_4444,N_4302,N_4373);
nor U4445 (N_4445,N_4235,N_4221);
and U4446 (N_4446,N_4287,N_4337);
or U4447 (N_4447,N_4218,N_4341);
nor U4448 (N_4448,N_4292,N_4334);
or U4449 (N_4449,N_4269,N_4388);
nand U4450 (N_4450,N_4389,N_4217);
nor U4451 (N_4451,N_4359,N_4215);
or U4452 (N_4452,N_4275,N_4278);
or U4453 (N_4453,N_4289,N_4369);
nor U4454 (N_4454,N_4326,N_4281);
nand U4455 (N_4455,N_4212,N_4222);
and U4456 (N_4456,N_4322,N_4236);
or U4457 (N_4457,N_4279,N_4202);
and U4458 (N_4458,N_4335,N_4353);
nand U4459 (N_4459,N_4345,N_4230);
nor U4460 (N_4460,N_4380,N_4300);
nand U4461 (N_4461,N_4209,N_4224);
nor U4462 (N_4462,N_4344,N_4213);
or U4463 (N_4463,N_4348,N_4210);
nor U4464 (N_4464,N_4374,N_4387);
nor U4465 (N_4465,N_4257,N_4200);
and U4466 (N_4466,N_4316,N_4272);
nand U4467 (N_4467,N_4350,N_4324);
nand U4468 (N_4468,N_4250,N_4290);
nor U4469 (N_4469,N_4311,N_4320);
or U4470 (N_4470,N_4237,N_4297);
nor U4471 (N_4471,N_4384,N_4354);
nor U4472 (N_4472,N_4382,N_4361);
nor U4473 (N_4473,N_4351,N_4398);
nand U4474 (N_4474,N_4204,N_4296);
nor U4475 (N_4475,N_4267,N_4314);
and U4476 (N_4476,N_4291,N_4277);
nand U4477 (N_4477,N_4394,N_4357);
nand U4478 (N_4478,N_4395,N_4333);
nand U4479 (N_4479,N_4286,N_4386);
or U4480 (N_4480,N_4239,N_4234);
nor U4481 (N_4481,N_4283,N_4313);
nand U4482 (N_4482,N_4392,N_4295);
nand U4483 (N_4483,N_4271,N_4370);
or U4484 (N_4484,N_4293,N_4276);
and U4485 (N_4485,N_4261,N_4245);
and U4486 (N_4486,N_4319,N_4312);
nor U4487 (N_4487,N_4308,N_4246);
and U4488 (N_4488,N_4383,N_4228);
or U4489 (N_4489,N_4329,N_4349);
nand U4490 (N_4490,N_4303,N_4306);
or U4491 (N_4491,N_4317,N_4254);
nand U4492 (N_4492,N_4340,N_4342);
nor U4493 (N_4493,N_4381,N_4252);
nand U4494 (N_4494,N_4331,N_4325);
or U4495 (N_4495,N_4207,N_4243);
and U4496 (N_4496,N_4347,N_4305);
nand U4497 (N_4497,N_4282,N_4309);
nor U4498 (N_4498,N_4203,N_4360);
xor U4499 (N_4499,N_4365,N_4253);
nor U4500 (N_4500,N_4212,N_4332);
and U4501 (N_4501,N_4278,N_4374);
nand U4502 (N_4502,N_4399,N_4242);
and U4503 (N_4503,N_4343,N_4395);
nand U4504 (N_4504,N_4281,N_4368);
or U4505 (N_4505,N_4380,N_4223);
nor U4506 (N_4506,N_4310,N_4274);
nand U4507 (N_4507,N_4292,N_4281);
or U4508 (N_4508,N_4359,N_4300);
nor U4509 (N_4509,N_4340,N_4359);
and U4510 (N_4510,N_4387,N_4341);
nor U4511 (N_4511,N_4312,N_4235);
or U4512 (N_4512,N_4293,N_4324);
and U4513 (N_4513,N_4381,N_4327);
nand U4514 (N_4514,N_4231,N_4217);
xor U4515 (N_4515,N_4326,N_4391);
and U4516 (N_4516,N_4263,N_4347);
and U4517 (N_4517,N_4205,N_4246);
or U4518 (N_4518,N_4373,N_4241);
nor U4519 (N_4519,N_4224,N_4358);
or U4520 (N_4520,N_4226,N_4397);
nand U4521 (N_4521,N_4396,N_4241);
xnor U4522 (N_4522,N_4360,N_4394);
nand U4523 (N_4523,N_4361,N_4224);
nor U4524 (N_4524,N_4307,N_4323);
or U4525 (N_4525,N_4206,N_4225);
or U4526 (N_4526,N_4305,N_4254);
or U4527 (N_4527,N_4264,N_4327);
nor U4528 (N_4528,N_4259,N_4353);
nor U4529 (N_4529,N_4281,N_4273);
or U4530 (N_4530,N_4244,N_4375);
nand U4531 (N_4531,N_4388,N_4266);
nor U4532 (N_4532,N_4326,N_4365);
and U4533 (N_4533,N_4251,N_4220);
nor U4534 (N_4534,N_4236,N_4224);
nand U4535 (N_4535,N_4378,N_4272);
and U4536 (N_4536,N_4247,N_4342);
and U4537 (N_4537,N_4394,N_4388);
nand U4538 (N_4538,N_4219,N_4330);
nor U4539 (N_4539,N_4220,N_4291);
nor U4540 (N_4540,N_4396,N_4246);
or U4541 (N_4541,N_4392,N_4346);
nor U4542 (N_4542,N_4309,N_4367);
or U4543 (N_4543,N_4378,N_4314);
nor U4544 (N_4544,N_4392,N_4271);
and U4545 (N_4545,N_4261,N_4292);
nor U4546 (N_4546,N_4301,N_4316);
nand U4547 (N_4547,N_4345,N_4394);
nor U4548 (N_4548,N_4307,N_4299);
xor U4549 (N_4549,N_4339,N_4331);
nor U4550 (N_4550,N_4226,N_4212);
xnor U4551 (N_4551,N_4369,N_4306);
xnor U4552 (N_4552,N_4319,N_4317);
and U4553 (N_4553,N_4288,N_4214);
or U4554 (N_4554,N_4388,N_4300);
and U4555 (N_4555,N_4248,N_4221);
and U4556 (N_4556,N_4233,N_4340);
or U4557 (N_4557,N_4200,N_4309);
xor U4558 (N_4558,N_4213,N_4332);
and U4559 (N_4559,N_4200,N_4364);
or U4560 (N_4560,N_4309,N_4340);
or U4561 (N_4561,N_4300,N_4298);
and U4562 (N_4562,N_4392,N_4263);
nand U4563 (N_4563,N_4221,N_4362);
nand U4564 (N_4564,N_4289,N_4383);
nor U4565 (N_4565,N_4250,N_4312);
xnor U4566 (N_4566,N_4212,N_4243);
nor U4567 (N_4567,N_4375,N_4352);
nor U4568 (N_4568,N_4298,N_4211);
nor U4569 (N_4569,N_4206,N_4335);
nand U4570 (N_4570,N_4236,N_4213);
xor U4571 (N_4571,N_4247,N_4272);
nor U4572 (N_4572,N_4218,N_4391);
or U4573 (N_4573,N_4399,N_4392);
and U4574 (N_4574,N_4258,N_4260);
nor U4575 (N_4575,N_4240,N_4362);
or U4576 (N_4576,N_4366,N_4306);
nand U4577 (N_4577,N_4378,N_4224);
and U4578 (N_4578,N_4295,N_4297);
or U4579 (N_4579,N_4231,N_4330);
nor U4580 (N_4580,N_4210,N_4217);
nor U4581 (N_4581,N_4292,N_4212);
nand U4582 (N_4582,N_4304,N_4202);
or U4583 (N_4583,N_4393,N_4280);
nand U4584 (N_4584,N_4213,N_4226);
nor U4585 (N_4585,N_4365,N_4204);
nand U4586 (N_4586,N_4292,N_4270);
nand U4587 (N_4587,N_4250,N_4240);
nand U4588 (N_4588,N_4314,N_4248);
or U4589 (N_4589,N_4274,N_4394);
nor U4590 (N_4590,N_4303,N_4201);
or U4591 (N_4591,N_4371,N_4262);
and U4592 (N_4592,N_4390,N_4241);
or U4593 (N_4593,N_4283,N_4364);
nor U4594 (N_4594,N_4226,N_4340);
nor U4595 (N_4595,N_4296,N_4372);
nor U4596 (N_4596,N_4264,N_4209);
or U4597 (N_4597,N_4270,N_4260);
or U4598 (N_4598,N_4353,N_4347);
and U4599 (N_4599,N_4253,N_4220);
nor U4600 (N_4600,N_4581,N_4465);
xor U4601 (N_4601,N_4573,N_4531);
and U4602 (N_4602,N_4453,N_4556);
nor U4603 (N_4603,N_4414,N_4549);
and U4604 (N_4604,N_4506,N_4517);
nor U4605 (N_4605,N_4534,N_4522);
or U4606 (N_4606,N_4539,N_4508);
and U4607 (N_4607,N_4553,N_4408);
nand U4608 (N_4608,N_4528,N_4463);
or U4609 (N_4609,N_4430,N_4524);
nor U4610 (N_4610,N_4477,N_4546);
nor U4611 (N_4611,N_4419,N_4564);
and U4612 (N_4612,N_4421,N_4501);
or U4613 (N_4613,N_4472,N_4409);
nor U4614 (N_4614,N_4505,N_4586);
nand U4615 (N_4615,N_4494,N_4563);
xnor U4616 (N_4616,N_4545,N_4535);
nand U4617 (N_4617,N_4441,N_4440);
nor U4618 (N_4618,N_4500,N_4540);
or U4619 (N_4619,N_4491,N_4555);
nor U4620 (N_4620,N_4589,N_4541);
nand U4621 (N_4621,N_4562,N_4485);
nand U4622 (N_4622,N_4426,N_4410);
nor U4623 (N_4623,N_4418,N_4436);
and U4624 (N_4624,N_4442,N_4484);
or U4625 (N_4625,N_4527,N_4544);
and U4626 (N_4626,N_4515,N_4425);
and U4627 (N_4627,N_4446,N_4497);
nand U4628 (N_4628,N_4449,N_4483);
nand U4629 (N_4629,N_4424,N_4513);
nand U4630 (N_4630,N_4478,N_4413);
nand U4631 (N_4631,N_4536,N_4530);
or U4632 (N_4632,N_4594,N_4575);
nor U4633 (N_4633,N_4595,N_4512);
nor U4634 (N_4634,N_4474,N_4403);
or U4635 (N_4635,N_4554,N_4489);
nor U4636 (N_4636,N_4407,N_4533);
xnor U4637 (N_4637,N_4591,N_4572);
and U4638 (N_4638,N_4461,N_4538);
or U4639 (N_4639,N_4420,N_4401);
nor U4640 (N_4640,N_4509,N_4570);
nand U4641 (N_4641,N_4473,N_4510);
or U4642 (N_4642,N_4558,N_4495);
nand U4643 (N_4643,N_4415,N_4464);
nor U4644 (N_4644,N_4499,N_4592);
nand U4645 (N_4645,N_4585,N_4435);
nor U4646 (N_4646,N_4576,N_4571);
nor U4647 (N_4647,N_4525,N_4526);
xnor U4648 (N_4648,N_4588,N_4561);
nand U4649 (N_4649,N_4577,N_4458);
or U4650 (N_4650,N_4565,N_4502);
xnor U4651 (N_4651,N_4516,N_4411);
or U4652 (N_4652,N_4537,N_4490);
xnor U4653 (N_4653,N_4593,N_4496);
nor U4654 (N_4654,N_4404,N_4569);
and U4655 (N_4655,N_4559,N_4479);
and U4656 (N_4656,N_4417,N_4429);
or U4657 (N_4657,N_4596,N_4583);
and U4658 (N_4658,N_4460,N_4574);
or U4659 (N_4659,N_4511,N_4462);
and U4660 (N_4660,N_4590,N_4523);
and U4661 (N_4661,N_4437,N_4503);
and U4662 (N_4662,N_4599,N_4434);
nand U4663 (N_4663,N_4433,N_4514);
and U4664 (N_4664,N_4551,N_4492);
nand U4665 (N_4665,N_4470,N_4456);
or U4666 (N_4666,N_4468,N_4486);
nor U4667 (N_4667,N_4582,N_4480);
or U4668 (N_4668,N_4432,N_4439);
xor U4669 (N_4669,N_4469,N_4405);
nand U4670 (N_4670,N_4457,N_4428);
or U4671 (N_4671,N_4507,N_4493);
nand U4672 (N_4672,N_4459,N_4438);
nor U4673 (N_4673,N_4443,N_4482);
nand U4674 (N_4674,N_4447,N_4452);
and U4675 (N_4675,N_4542,N_4498);
nor U4676 (N_4676,N_4520,N_4579);
nand U4677 (N_4677,N_4552,N_4543);
nor U4678 (N_4678,N_4548,N_4597);
xnor U4679 (N_4679,N_4475,N_4444);
or U4680 (N_4680,N_4578,N_4402);
and U4681 (N_4681,N_4532,N_4406);
and U4682 (N_4682,N_4400,N_4566);
nor U4683 (N_4683,N_4451,N_4547);
or U4684 (N_4684,N_4454,N_4450);
and U4685 (N_4685,N_4567,N_4557);
and U4686 (N_4686,N_4445,N_4521);
and U4687 (N_4687,N_4584,N_4431);
and U4688 (N_4688,N_4423,N_4568);
nor U4689 (N_4689,N_4427,N_4481);
nand U4690 (N_4690,N_4560,N_4504);
nor U4691 (N_4691,N_4580,N_4448);
nor U4692 (N_4692,N_4412,N_4471);
nor U4693 (N_4693,N_4467,N_4488);
or U4694 (N_4694,N_4587,N_4455);
nand U4695 (N_4695,N_4519,N_4487);
nor U4696 (N_4696,N_4598,N_4550);
nor U4697 (N_4697,N_4422,N_4466);
or U4698 (N_4698,N_4518,N_4476);
nor U4699 (N_4699,N_4529,N_4416);
xnor U4700 (N_4700,N_4524,N_4461);
and U4701 (N_4701,N_4430,N_4506);
and U4702 (N_4702,N_4567,N_4527);
xor U4703 (N_4703,N_4433,N_4415);
and U4704 (N_4704,N_4560,N_4432);
xnor U4705 (N_4705,N_4574,N_4554);
xor U4706 (N_4706,N_4437,N_4495);
nor U4707 (N_4707,N_4483,N_4447);
nor U4708 (N_4708,N_4498,N_4480);
or U4709 (N_4709,N_4534,N_4495);
nand U4710 (N_4710,N_4502,N_4559);
or U4711 (N_4711,N_4467,N_4588);
or U4712 (N_4712,N_4506,N_4509);
and U4713 (N_4713,N_4474,N_4426);
or U4714 (N_4714,N_4529,N_4571);
or U4715 (N_4715,N_4466,N_4495);
nand U4716 (N_4716,N_4404,N_4431);
or U4717 (N_4717,N_4581,N_4506);
nor U4718 (N_4718,N_4476,N_4578);
and U4719 (N_4719,N_4531,N_4517);
or U4720 (N_4720,N_4591,N_4461);
xor U4721 (N_4721,N_4492,N_4488);
nand U4722 (N_4722,N_4444,N_4429);
and U4723 (N_4723,N_4402,N_4585);
or U4724 (N_4724,N_4555,N_4437);
nand U4725 (N_4725,N_4480,N_4465);
and U4726 (N_4726,N_4452,N_4443);
xor U4727 (N_4727,N_4588,N_4446);
nor U4728 (N_4728,N_4584,N_4593);
nor U4729 (N_4729,N_4443,N_4490);
nor U4730 (N_4730,N_4499,N_4549);
nor U4731 (N_4731,N_4550,N_4485);
nor U4732 (N_4732,N_4408,N_4496);
nor U4733 (N_4733,N_4569,N_4555);
and U4734 (N_4734,N_4557,N_4508);
nand U4735 (N_4735,N_4494,N_4502);
xor U4736 (N_4736,N_4582,N_4521);
and U4737 (N_4737,N_4483,N_4563);
and U4738 (N_4738,N_4414,N_4473);
nor U4739 (N_4739,N_4579,N_4495);
or U4740 (N_4740,N_4549,N_4538);
nand U4741 (N_4741,N_4472,N_4504);
nand U4742 (N_4742,N_4591,N_4449);
and U4743 (N_4743,N_4533,N_4517);
nand U4744 (N_4744,N_4552,N_4536);
and U4745 (N_4745,N_4525,N_4409);
and U4746 (N_4746,N_4430,N_4456);
or U4747 (N_4747,N_4543,N_4590);
and U4748 (N_4748,N_4489,N_4563);
and U4749 (N_4749,N_4453,N_4588);
or U4750 (N_4750,N_4586,N_4442);
xnor U4751 (N_4751,N_4458,N_4566);
nor U4752 (N_4752,N_4533,N_4585);
and U4753 (N_4753,N_4401,N_4596);
and U4754 (N_4754,N_4510,N_4409);
nor U4755 (N_4755,N_4522,N_4549);
xor U4756 (N_4756,N_4473,N_4519);
or U4757 (N_4757,N_4511,N_4425);
nor U4758 (N_4758,N_4410,N_4445);
xor U4759 (N_4759,N_4548,N_4537);
xor U4760 (N_4760,N_4563,N_4559);
or U4761 (N_4761,N_4587,N_4579);
nand U4762 (N_4762,N_4454,N_4536);
or U4763 (N_4763,N_4478,N_4546);
nand U4764 (N_4764,N_4430,N_4481);
or U4765 (N_4765,N_4468,N_4496);
and U4766 (N_4766,N_4473,N_4406);
or U4767 (N_4767,N_4481,N_4574);
and U4768 (N_4768,N_4567,N_4442);
or U4769 (N_4769,N_4504,N_4576);
xnor U4770 (N_4770,N_4475,N_4428);
or U4771 (N_4771,N_4466,N_4594);
nor U4772 (N_4772,N_4417,N_4557);
nand U4773 (N_4773,N_4434,N_4530);
nand U4774 (N_4774,N_4598,N_4437);
and U4775 (N_4775,N_4447,N_4485);
xnor U4776 (N_4776,N_4412,N_4510);
nand U4777 (N_4777,N_4448,N_4483);
and U4778 (N_4778,N_4435,N_4416);
nor U4779 (N_4779,N_4586,N_4407);
nand U4780 (N_4780,N_4505,N_4424);
nor U4781 (N_4781,N_4475,N_4483);
or U4782 (N_4782,N_4406,N_4552);
nor U4783 (N_4783,N_4487,N_4498);
nand U4784 (N_4784,N_4416,N_4542);
and U4785 (N_4785,N_4475,N_4548);
and U4786 (N_4786,N_4590,N_4495);
nand U4787 (N_4787,N_4491,N_4564);
and U4788 (N_4788,N_4473,N_4514);
or U4789 (N_4789,N_4597,N_4425);
and U4790 (N_4790,N_4496,N_4461);
or U4791 (N_4791,N_4564,N_4426);
nand U4792 (N_4792,N_4430,N_4421);
and U4793 (N_4793,N_4480,N_4441);
or U4794 (N_4794,N_4480,N_4504);
nor U4795 (N_4795,N_4567,N_4475);
nand U4796 (N_4796,N_4516,N_4598);
nor U4797 (N_4797,N_4482,N_4413);
nand U4798 (N_4798,N_4457,N_4590);
nand U4799 (N_4799,N_4462,N_4580);
nor U4800 (N_4800,N_4767,N_4725);
and U4801 (N_4801,N_4620,N_4710);
or U4802 (N_4802,N_4751,N_4785);
and U4803 (N_4803,N_4789,N_4649);
nand U4804 (N_4804,N_4614,N_4708);
nor U4805 (N_4805,N_4702,N_4713);
nand U4806 (N_4806,N_4752,N_4659);
nand U4807 (N_4807,N_4731,N_4775);
nand U4808 (N_4808,N_4791,N_4683);
and U4809 (N_4809,N_4719,N_4703);
and U4810 (N_4810,N_4625,N_4726);
and U4811 (N_4811,N_4691,N_4641);
nand U4812 (N_4812,N_4743,N_4681);
nand U4813 (N_4813,N_4701,N_4788);
or U4814 (N_4814,N_4632,N_4772);
or U4815 (N_4815,N_4796,N_4643);
nand U4816 (N_4816,N_4697,N_4766);
xnor U4817 (N_4817,N_4673,N_4768);
nor U4818 (N_4818,N_4685,N_4780);
nor U4819 (N_4819,N_4642,N_4727);
and U4820 (N_4820,N_4795,N_4774);
or U4821 (N_4821,N_4686,N_4636);
and U4822 (N_4822,N_4630,N_4600);
nand U4823 (N_4823,N_4656,N_4604);
nor U4824 (N_4824,N_4711,N_4737);
and U4825 (N_4825,N_4682,N_4666);
and U4826 (N_4826,N_4793,N_4650);
and U4827 (N_4827,N_4669,N_4709);
nand U4828 (N_4828,N_4657,N_4733);
or U4829 (N_4829,N_4741,N_4618);
and U4830 (N_4830,N_4738,N_4615);
or U4831 (N_4831,N_4716,N_4704);
nand U4832 (N_4832,N_4748,N_4706);
nor U4833 (N_4833,N_4693,N_4621);
or U4834 (N_4834,N_4779,N_4690);
nor U4835 (N_4835,N_4714,N_4728);
nand U4836 (N_4836,N_4646,N_4660);
nor U4837 (N_4837,N_4663,N_4652);
and U4838 (N_4838,N_4707,N_4696);
or U4839 (N_4839,N_4611,N_4603);
or U4840 (N_4840,N_4765,N_4665);
xnor U4841 (N_4841,N_4626,N_4799);
and U4842 (N_4842,N_4648,N_4721);
or U4843 (N_4843,N_4671,N_4672);
nand U4844 (N_4844,N_4638,N_4722);
or U4845 (N_4845,N_4602,N_4645);
nand U4846 (N_4846,N_4678,N_4605);
or U4847 (N_4847,N_4684,N_4769);
or U4848 (N_4848,N_4732,N_4613);
or U4849 (N_4849,N_4745,N_4736);
nand U4850 (N_4850,N_4616,N_4631);
or U4851 (N_4851,N_4670,N_4720);
nand U4852 (N_4852,N_4633,N_4667);
nor U4853 (N_4853,N_4723,N_4661);
or U4854 (N_4854,N_4692,N_4781);
nor U4855 (N_4855,N_4609,N_4755);
and U4856 (N_4856,N_4792,N_4607);
nand U4857 (N_4857,N_4759,N_4662);
nor U4858 (N_4858,N_4730,N_4658);
and U4859 (N_4859,N_4762,N_4651);
and U4860 (N_4860,N_4610,N_4601);
or U4861 (N_4861,N_4689,N_4778);
nand U4862 (N_4862,N_4739,N_4655);
and U4863 (N_4863,N_4680,N_4699);
nor U4864 (N_4864,N_4623,N_4757);
nor U4865 (N_4865,N_4679,N_4771);
nand U4866 (N_4866,N_4634,N_4617);
nor U4867 (N_4867,N_4742,N_4787);
nor U4868 (N_4868,N_4606,N_4729);
nor U4869 (N_4869,N_4746,N_4770);
and U4870 (N_4870,N_4694,N_4777);
nand U4871 (N_4871,N_4763,N_4676);
nor U4872 (N_4872,N_4627,N_4744);
nor U4873 (N_4873,N_4688,N_4776);
nor U4874 (N_4874,N_4717,N_4760);
nor U4875 (N_4875,N_4794,N_4654);
xnor U4876 (N_4876,N_4647,N_4644);
nand U4877 (N_4877,N_4653,N_4756);
or U4878 (N_4878,N_4718,N_4750);
and U4879 (N_4879,N_4734,N_4624);
or U4880 (N_4880,N_4687,N_4747);
or U4881 (N_4881,N_4764,N_4783);
xnor U4882 (N_4882,N_4675,N_4677);
or U4883 (N_4883,N_4619,N_4705);
or U4884 (N_4884,N_4754,N_4640);
nand U4885 (N_4885,N_4695,N_4790);
or U4886 (N_4886,N_4761,N_4668);
and U4887 (N_4887,N_4608,N_4715);
nand U4888 (N_4888,N_4622,N_4664);
nor U4889 (N_4889,N_4637,N_4782);
and U4890 (N_4890,N_4773,N_4639);
nor U4891 (N_4891,N_4628,N_4629);
and U4892 (N_4892,N_4698,N_4724);
and U4893 (N_4893,N_4735,N_4612);
xnor U4894 (N_4894,N_4749,N_4797);
and U4895 (N_4895,N_4798,N_4635);
nor U4896 (N_4896,N_4674,N_4784);
xnor U4897 (N_4897,N_4712,N_4786);
and U4898 (N_4898,N_4700,N_4740);
and U4899 (N_4899,N_4758,N_4753);
nand U4900 (N_4900,N_4685,N_4777);
and U4901 (N_4901,N_4664,N_4797);
and U4902 (N_4902,N_4744,N_4628);
nand U4903 (N_4903,N_4649,N_4627);
or U4904 (N_4904,N_4785,N_4711);
nand U4905 (N_4905,N_4741,N_4787);
and U4906 (N_4906,N_4771,N_4621);
xnor U4907 (N_4907,N_4762,N_4721);
nand U4908 (N_4908,N_4701,N_4601);
nor U4909 (N_4909,N_4635,N_4759);
and U4910 (N_4910,N_4771,N_4675);
or U4911 (N_4911,N_4603,N_4794);
nor U4912 (N_4912,N_4715,N_4732);
nand U4913 (N_4913,N_4652,N_4759);
or U4914 (N_4914,N_4611,N_4758);
or U4915 (N_4915,N_4624,N_4744);
nor U4916 (N_4916,N_4677,N_4763);
nor U4917 (N_4917,N_4768,N_4722);
or U4918 (N_4918,N_4651,N_4698);
nand U4919 (N_4919,N_4646,N_4689);
or U4920 (N_4920,N_4739,N_4787);
or U4921 (N_4921,N_4648,N_4602);
nand U4922 (N_4922,N_4778,N_4638);
nand U4923 (N_4923,N_4755,N_4669);
and U4924 (N_4924,N_4766,N_4643);
nor U4925 (N_4925,N_4739,N_4659);
or U4926 (N_4926,N_4702,N_4645);
nand U4927 (N_4927,N_4673,N_4742);
xor U4928 (N_4928,N_4789,N_4700);
nor U4929 (N_4929,N_4620,N_4689);
or U4930 (N_4930,N_4789,N_4659);
xnor U4931 (N_4931,N_4610,N_4707);
or U4932 (N_4932,N_4755,N_4654);
and U4933 (N_4933,N_4697,N_4765);
and U4934 (N_4934,N_4743,N_4706);
nor U4935 (N_4935,N_4765,N_4768);
and U4936 (N_4936,N_4604,N_4715);
and U4937 (N_4937,N_4624,N_4720);
nor U4938 (N_4938,N_4677,N_4793);
and U4939 (N_4939,N_4789,N_4776);
xnor U4940 (N_4940,N_4720,N_4740);
and U4941 (N_4941,N_4636,N_4764);
nand U4942 (N_4942,N_4771,N_4781);
or U4943 (N_4943,N_4689,N_4619);
xnor U4944 (N_4944,N_4776,N_4738);
nand U4945 (N_4945,N_4723,N_4707);
or U4946 (N_4946,N_4780,N_4686);
and U4947 (N_4947,N_4616,N_4716);
nor U4948 (N_4948,N_4786,N_4738);
nand U4949 (N_4949,N_4782,N_4781);
or U4950 (N_4950,N_4740,N_4625);
or U4951 (N_4951,N_4755,N_4744);
or U4952 (N_4952,N_4739,N_4785);
and U4953 (N_4953,N_4653,N_4749);
and U4954 (N_4954,N_4628,N_4793);
nor U4955 (N_4955,N_4754,N_4631);
or U4956 (N_4956,N_4762,N_4772);
xor U4957 (N_4957,N_4639,N_4665);
and U4958 (N_4958,N_4710,N_4680);
or U4959 (N_4959,N_4672,N_4616);
nand U4960 (N_4960,N_4737,N_4708);
and U4961 (N_4961,N_4769,N_4763);
or U4962 (N_4962,N_4702,N_4609);
xor U4963 (N_4963,N_4741,N_4687);
nand U4964 (N_4964,N_4764,N_4799);
or U4965 (N_4965,N_4728,N_4668);
nor U4966 (N_4966,N_4715,N_4666);
or U4967 (N_4967,N_4650,N_4679);
nor U4968 (N_4968,N_4615,N_4621);
or U4969 (N_4969,N_4675,N_4725);
and U4970 (N_4970,N_4606,N_4616);
nor U4971 (N_4971,N_4777,N_4788);
nor U4972 (N_4972,N_4740,N_4656);
xor U4973 (N_4973,N_4669,N_4620);
xnor U4974 (N_4974,N_4667,N_4768);
or U4975 (N_4975,N_4628,N_4697);
nor U4976 (N_4976,N_4764,N_4781);
nand U4977 (N_4977,N_4779,N_4684);
nor U4978 (N_4978,N_4759,N_4624);
nand U4979 (N_4979,N_4763,N_4709);
or U4980 (N_4980,N_4748,N_4776);
xnor U4981 (N_4981,N_4742,N_4609);
xor U4982 (N_4982,N_4741,N_4701);
xnor U4983 (N_4983,N_4650,N_4798);
nand U4984 (N_4984,N_4723,N_4677);
and U4985 (N_4985,N_4607,N_4699);
nand U4986 (N_4986,N_4708,N_4679);
and U4987 (N_4987,N_4736,N_4784);
or U4988 (N_4988,N_4763,N_4631);
and U4989 (N_4989,N_4668,N_4741);
nand U4990 (N_4990,N_4682,N_4795);
or U4991 (N_4991,N_4743,N_4679);
and U4992 (N_4992,N_4751,N_4735);
nor U4993 (N_4993,N_4670,N_4623);
and U4994 (N_4994,N_4732,N_4669);
or U4995 (N_4995,N_4747,N_4658);
nor U4996 (N_4996,N_4715,N_4672);
and U4997 (N_4997,N_4797,N_4630);
and U4998 (N_4998,N_4603,N_4651);
nand U4999 (N_4999,N_4783,N_4639);
nand U5000 (N_5000,N_4959,N_4981);
nand U5001 (N_5001,N_4936,N_4993);
and U5002 (N_5002,N_4968,N_4962);
or U5003 (N_5003,N_4848,N_4886);
nor U5004 (N_5004,N_4902,N_4854);
nand U5005 (N_5005,N_4914,N_4892);
nor U5006 (N_5006,N_4957,N_4916);
and U5007 (N_5007,N_4982,N_4844);
and U5008 (N_5008,N_4926,N_4950);
and U5009 (N_5009,N_4822,N_4846);
nor U5010 (N_5010,N_4823,N_4992);
nand U5011 (N_5011,N_4937,N_4866);
nand U5012 (N_5012,N_4975,N_4842);
or U5013 (N_5013,N_4881,N_4988);
or U5014 (N_5014,N_4915,N_4999);
or U5015 (N_5015,N_4851,N_4969);
or U5016 (N_5016,N_4889,N_4845);
or U5017 (N_5017,N_4973,N_4820);
and U5018 (N_5018,N_4928,N_4977);
and U5019 (N_5019,N_4841,N_4879);
and U5020 (N_5020,N_4805,N_4954);
nor U5021 (N_5021,N_4939,N_4890);
nand U5022 (N_5022,N_4813,N_4903);
nor U5023 (N_5023,N_4897,N_4898);
or U5024 (N_5024,N_4967,N_4861);
or U5025 (N_5025,N_4933,N_4833);
nor U5026 (N_5026,N_4945,N_4989);
xnor U5027 (N_5027,N_4900,N_4987);
nor U5028 (N_5028,N_4811,N_4994);
nand U5029 (N_5029,N_4852,N_4877);
and U5030 (N_5030,N_4932,N_4971);
nand U5031 (N_5031,N_4834,N_4947);
or U5032 (N_5032,N_4893,N_4955);
nand U5033 (N_5033,N_4850,N_4864);
nor U5034 (N_5034,N_4995,N_4817);
or U5035 (N_5035,N_4983,N_4942);
nor U5036 (N_5036,N_4878,N_4929);
nor U5037 (N_5037,N_4944,N_4910);
and U5038 (N_5038,N_4904,N_4906);
nand U5039 (N_5039,N_4899,N_4991);
and U5040 (N_5040,N_4818,N_4888);
or U5041 (N_5041,N_4951,N_4857);
nor U5042 (N_5042,N_4940,N_4908);
or U5043 (N_5043,N_4815,N_4853);
nand U5044 (N_5044,N_4804,N_4816);
xor U5045 (N_5045,N_4997,N_4985);
and U5046 (N_5046,N_4913,N_4812);
nor U5047 (N_5047,N_4838,N_4880);
nor U5048 (N_5048,N_4986,N_4839);
nand U5049 (N_5049,N_4927,N_4948);
and U5050 (N_5050,N_4949,N_4867);
nor U5051 (N_5051,N_4829,N_4996);
nand U5052 (N_5052,N_4882,N_4855);
xor U5053 (N_5053,N_4966,N_4843);
and U5054 (N_5054,N_4935,N_4911);
xnor U5055 (N_5055,N_4946,N_4847);
nor U5056 (N_5056,N_4980,N_4970);
nor U5057 (N_5057,N_4923,N_4802);
nor U5058 (N_5058,N_4919,N_4803);
nor U5059 (N_5059,N_4896,N_4930);
and U5060 (N_5060,N_4891,N_4874);
or U5061 (N_5061,N_4840,N_4974);
nor U5062 (N_5062,N_4863,N_4821);
or U5063 (N_5063,N_4826,N_4810);
nand U5064 (N_5064,N_4998,N_4885);
or U5065 (N_5065,N_4871,N_4809);
nor U5066 (N_5066,N_4835,N_4963);
nor U5067 (N_5067,N_4827,N_4984);
nand U5068 (N_5068,N_4925,N_4979);
and U5069 (N_5069,N_4934,N_4894);
nor U5070 (N_5070,N_4941,N_4917);
and U5071 (N_5071,N_4859,N_4868);
or U5072 (N_5072,N_4953,N_4924);
or U5073 (N_5073,N_4832,N_4865);
nand U5074 (N_5074,N_4901,N_4800);
nand U5075 (N_5075,N_4907,N_4801);
nand U5076 (N_5076,N_4976,N_4828);
nor U5077 (N_5077,N_4819,N_4884);
nand U5078 (N_5078,N_4912,N_4836);
and U5079 (N_5079,N_4860,N_4808);
nor U5080 (N_5080,N_4825,N_4943);
nand U5081 (N_5081,N_4831,N_4869);
nor U5082 (N_5082,N_4883,N_4972);
nor U5083 (N_5083,N_4876,N_4921);
or U5084 (N_5084,N_4920,N_4870);
and U5085 (N_5085,N_4958,N_4887);
nor U5086 (N_5086,N_4806,N_4814);
or U5087 (N_5087,N_4849,N_4978);
nand U5088 (N_5088,N_4918,N_4938);
and U5089 (N_5089,N_4895,N_4965);
xnor U5090 (N_5090,N_4961,N_4830);
and U5091 (N_5091,N_4824,N_4909);
nor U5092 (N_5092,N_4875,N_4931);
and U5093 (N_5093,N_4858,N_4873);
nand U5094 (N_5094,N_4872,N_4837);
nand U5095 (N_5095,N_4922,N_4964);
nor U5096 (N_5096,N_4990,N_4960);
and U5097 (N_5097,N_4905,N_4952);
nand U5098 (N_5098,N_4856,N_4862);
nor U5099 (N_5099,N_4807,N_4956);
xor U5100 (N_5100,N_4818,N_4932);
or U5101 (N_5101,N_4851,N_4870);
and U5102 (N_5102,N_4824,N_4865);
or U5103 (N_5103,N_4953,N_4853);
nand U5104 (N_5104,N_4925,N_4816);
and U5105 (N_5105,N_4970,N_4820);
or U5106 (N_5106,N_4925,N_4827);
nor U5107 (N_5107,N_4935,N_4907);
nor U5108 (N_5108,N_4872,N_4980);
nor U5109 (N_5109,N_4879,N_4898);
nand U5110 (N_5110,N_4854,N_4827);
or U5111 (N_5111,N_4958,N_4944);
and U5112 (N_5112,N_4891,N_4862);
or U5113 (N_5113,N_4982,N_4911);
or U5114 (N_5114,N_4990,N_4974);
nand U5115 (N_5115,N_4846,N_4939);
nand U5116 (N_5116,N_4809,N_4963);
nor U5117 (N_5117,N_4854,N_4844);
nand U5118 (N_5118,N_4946,N_4899);
or U5119 (N_5119,N_4907,N_4967);
nand U5120 (N_5120,N_4876,N_4882);
or U5121 (N_5121,N_4914,N_4961);
and U5122 (N_5122,N_4988,N_4800);
xor U5123 (N_5123,N_4963,N_4889);
nand U5124 (N_5124,N_4992,N_4876);
or U5125 (N_5125,N_4869,N_4990);
nor U5126 (N_5126,N_4896,N_4817);
or U5127 (N_5127,N_4874,N_4984);
and U5128 (N_5128,N_4993,N_4921);
nand U5129 (N_5129,N_4966,N_4838);
nor U5130 (N_5130,N_4992,N_4919);
nor U5131 (N_5131,N_4853,N_4835);
or U5132 (N_5132,N_4883,N_4897);
or U5133 (N_5133,N_4920,N_4975);
or U5134 (N_5134,N_4933,N_4907);
xnor U5135 (N_5135,N_4935,N_4849);
nand U5136 (N_5136,N_4876,N_4875);
or U5137 (N_5137,N_4820,N_4829);
and U5138 (N_5138,N_4889,N_4936);
or U5139 (N_5139,N_4962,N_4891);
and U5140 (N_5140,N_4844,N_4826);
nor U5141 (N_5141,N_4915,N_4930);
or U5142 (N_5142,N_4862,N_4879);
or U5143 (N_5143,N_4944,N_4891);
xor U5144 (N_5144,N_4886,N_4889);
or U5145 (N_5145,N_4829,N_4846);
and U5146 (N_5146,N_4999,N_4913);
nor U5147 (N_5147,N_4945,N_4850);
xnor U5148 (N_5148,N_4953,N_4914);
nand U5149 (N_5149,N_4925,N_4813);
and U5150 (N_5150,N_4856,N_4814);
xor U5151 (N_5151,N_4884,N_4964);
nand U5152 (N_5152,N_4973,N_4924);
xor U5153 (N_5153,N_4936,N_4864);
nand U5154 (N_5154,N_4917,N_4832);
or U5155 (N_5155,N_4991,N_4907);
xnor U5156 (N_5156,N_4810,N_4941);
nand U5157 (N_5157,N_4990,N_4910);
nand U5158 (N_5158,N_4879,N_4840);
or U5159 (N_5159,N_4964,N_4890);
or U5160 (N_5160,N_4836,N_4801);
nand U5161 (N_5161,N_4915,N_4929);
and U5162 (N_5162,N_4927,N_4956);
or U5163 (N_5163,N_4961,N_4978);
or U5164 (N_5164,N_4839,N_4925);
or U5165 (N_5165,N_4860,N_4930);
nor U5166 (N_5166,N_4970,N_4808);
nand U5167 (N_5167,N_4983,N_4988);
xor U5168 (N_5168,N_4844,N_4913);
xnor U5169 (N_5169,N_4899,N_4873);
nand U5170 (N_5170,N_4954,N_4925);
or U5171 (N_5171,N_4900,N_4831);
xor U5172 (N_5172,N_4854,N_4814);
or U5173 (N_5173,N_4854,N_4845);
nand U5174 (N_5174,N_4959,N_4829);
nand U5175 (N_5175,N_4996,N_4897);
and U5176 (N_5176,N_4873,N_4814);
and U5177 (N_5177,N_4968,N_4808);
or U5178 (N_5178,N_4851,N_4976);
or U5179 (N_5179,N_4905,N_4813);
or U5180 (N_5180,N_4928,N_4872);
or U5181 (N_5181,N_4822,N_4860);
and U5182 (N_5182,N_4922,N_4800);
or U5183 (N_5183,N_4911,N_4960);
nand U5184 (N_5184,N_4976,N_4819);
xnor U5185 (N_5185,N_4844,N_4882);
nor U5186 (N_5186,N_4814,N_4878);
or U5187 (N_5187,N_4834,N_4833);
and U5188 (N_5188,N_4968,N_4993);
and U5189 (N_5189,N_4828,N_4923);
xnor U5190 (N_5190,N_4943,N_4809);
and U5191 (N_5191,N_4937,N_4930);
nor U5192 (N_5192,N_4988,N_4878);
or U5193 (N_5193,N_4828,N_4857);
or U5194 (N_5194,N_4983,N_4944);
or U5195 (N_5195,N_4877,N_4840);
or U5196 (N_5196,N_4930,N_4859);
nor U5197 (N_5197,N_4883,N_4870);
nand U5198 (N_5198,N_4814,N_4963);
and U5199 (N_5199,N_4865,N_4976);
or U5200 (N_5200,N_5177,N_5156);
and U5201 (N_5201,N_5101,N_5066);
xor U5202 (N_5202,N_5144,N_5055);
nand U5203 (N_5203,N_5172,N_5143);
nand U5204 (N_5204,N_5104,N_5054);
nor U5205 (N_5205,N_5031,N_5073);
or U5206 (N_5206,N_5078,N_5019);
and U5207 (N_5207,N_5111,N_5180);
nand U5208 (N_5208,N_5158,N_5120);
or U5209 (N_5209,N_5110,N_5133);
and U5210 (N_5210,N_5174,N_5035);
and U5211 (N_5211,N_5163,N_5027);
nor U5212 (N_5212,N_5012,N_5173);
or U5213 (N_5213,N_5011,N_5103);
and U5214 (N_5214,N_5091,N_5128);
nand U5215 (N_5215,N_5152,N_5094);
and U5216 (N_5216,N_5171,N_5096);
nand U5217 (N_5217,N_5041,N_5070);
or U5218 (N_5218,N_5001,N_5068);
nor U5219 (N_5219,N_5048,N_5183);
nand U5220 (N_5220,N_5033,N_5131);
nor U5221 (N_5221,N_5017,N_5176);
nor U5222 (N_5222,N_5190,N_5112);
nor U5223 (N_5223,N_5077,N_5024);
nor U5224 (N_5224,N_5197,N_5058);
nor U5225 (N_5225,N_5010,N_5164);
nand U5226 (N_5226,N_5137,N_5045);
or U5227 (N_5227,N_5130,N_5123);
nand U5228 (N_5228,N_5006,N_5184);
or U5229 (N_5229,N_5047,N_5021);
and U5230 (N_5230,N_5149,N_5038);
nand U5231 (N_5231,N_5194,N_5060);
nand U5232 (N_5232,N_5052,N_5026);
or U5233 (N_5233,N_5046,N_5007);
nor U5234 (N_5234,N_5166,N_5051);
nor U5235 (N_5235,N_5132,N_5037);
nand U5236 (N_5236,N_5099,N_5134);
xor U5237 (N_5237,N_5022,N_5115);
or U5238 (N_5238,N_5072,N_5074);
nor U5239 (N_5239,N_5141,N_5168);
and U5240 (N_5240,N_5023,N_5125);
xor U5241 (N_5241,N_5043,N_5151);
xor U5242 (N_5242,N_5092,N_5015);
xnor U5243 (N_5243,N_5114,N_5162);
nand U5244 (N_5244,N_5097,N_5036);
or U5245 (N_5245,N_5161,N_5193);
nor U5246 (N_5246,N_5062,N_5109);
nand U5247 (N_5247,N_5185,N_5170);
nor U5248 (N_5248,N_5159,N_5102);
xnor U5249 (N_5249,N_5199,N_5155);
nand U5250 (N_5250,N_5080,N_5087);
nand U5251 (N_5251,N_5084,N_5121);
nand U5252 (N_5252,N_5067,N_5098);
or U5253 (N_5253,N_5196,N_5076);
nor U5254 (N_5254,N_5032,N_5028);
nand U5255 (N_5255,N_5086,N_5085);
and U5256 (N_5256,N_5083,N_5005);
xnor U5257 (N_5257,N_5105,N_5153);
or U5258 (N_5258,N_5139,N_5146);
nand U5259 (N_5259,N_5191,N_5082);
xnor U5260 (N_5260,N_5009,N_5063);
or U5261 (N_5261,N_5018,N_5142);
nor U5262 (N_5262,N_5044,N_5089);
or U5263 (N_5263,N_5020,N_5136);
nand U5264 (N_5264,N_5118,N_5002);
and U5265 (N_5265,N_5050,N_5004);
nand U5266 (N_5266,N_5056,N_5029);
nor U5267 (N_5267,N_5075,N_5003);
or U5268 (N_5268,N_5182,N_5117);
nor U5269 (N_5269,N_5129,N_5165);
nor U5270 (N_5270,N_5160,N_5100);
or U5271 (N_5271,N_5088,N_5138);
or U5272 (N_5272,N_5025,N_5127);
nor U5273 (N_5273,N_5154,N_5124);
or U5274 (N_5274,N_5049,N_5106);
or U5275 (N_5275,N_5040,N_5057);
or U5276 (N_5276,N_5065,N_5008);
nand U5277 (N_5277,N_5122,N_5150);
xnor U5278 (N_5278,N_5140,N_5169);
nand U5279 (N_5279,N_5187,N_5175);
nand U5280 (N_5280,N_5016,N_5167);
or U5281 (N_5281,N_5147,N_5192);
nand U5282 (N_5282,N_5116,N_5198);
nor U5283 (N_5283,N_5000,N_5108);
or U5284 (N_5284,N_5090,N_5178);
or U5285 (N_5285,N_5042,N_5093);
or U5286 (N_5286,N_5119,N_5030);
and U5287 (N_5287,N_5107,N_5081);
nand U5288 (N_5288,N_5079,N_5195);
and U5289 (N_5289,N_5059,N_5039);
nand U5290 (N_5290,N_5189,N_5095);
and U5291 (N_5291,N_5113,N_5013);
nand U5292 (N_5292,N_5064,N_5188);
nand U5293 (N_5293,N_5014,N_5157);
or U5294 (N_5294,N_5053,N_5135);
xnor U5295 (N_5295,N_5186,N_5061);
and U5296 (N_5296,N_5126,N_5181);
nor U5297 (N_5297,N_5069,N_5145);
xor U5298 (N_5298,N_5034,N_5179);
nand U5299 (N_5299,N_5071,N_5148);
nand U5300 (N_5300,N_5178,N_5022);
nor U5301 (N_5301,N_5082,N_5031);
or U5302 (N_5302,N_5171,N_5061);
nand U5303 (N_5303,N_5190,N_5099);
or U5304 (N_5304,N_5104,N_5138);
nor U5305 (N_5305,N_5075,N_5018);
nor U5306 (N_5306,N_5129,N_5154);
or U5307 (N_5307,N_5148,N_5193);
or U5308 (N_5308,N_5159,N_5145);
or U5309 (N_5309,N_5023,N_5019);
and U5310 (N_5310,N_5170,N_5088);
xor U5311 (N_5311,N_5075,N_5016);
nor U5312 (N_5312,N_5154,N_5033);
nand U5313 (N_5313,N_5090,N_5144);
nor U5314 (N_5314,N_5016,N_5039);
nor U5315 (N_5315,N_5013,N_5017);
and U5316 (N_5316,N_5164,N_5091);
nor U5317 (N_5317,N_5017,N_5022);
nand U5318 (N_5318,N_5003,N_5152);
nand U5319 (N_5319,N_5064,N_5075);
or U5320 (N_5320,N_5109,N_5174);
nand U5321 (N_5321,N_5146,N_5181);
nand U5322 (N_5322,N_5118,N_5053);
nand U5323 (N_5323,N_5152,N_5165);
nor U5324 (N_5324,N_5052,N_5015);
or U5325 (N_5325,N_5126,N_5043);
nand U5326 (N_5326,N_5004,N_5065);
nand U5327 (N_5327,N_5013,N_5063);
nor U5328 (N_5328,N_5140,N_5016);
or U5329 (N_5329,N_5191,N_5050);
or U5330 (N_5330,N_5191,N_5158);
nand U5331 (N_5331,N_5064,N_5082);
nand U5332 (N_5332,N_5162,N_5175);
or U5333 (N_5333,N_5185,N_5025);
nor U5334 (N_5334,N_5056,N_5184);
nor U5335 (N_5335,N_5103,N_5072);
or U5336 (N_5336,N_5057,N_5153);
nor U5337 (N_5337,N_5044,N_5031);
and U5338 (N_5338,N_5152,N_5101);
nor U5339 (N_5339,N_5065,N_5105);
or U5340 (N_5340,N_5098,N_5045);
nor U5341 (N_5341,N_5125,N_5155);
and U5342 (N_5342,N_5086,N_5189);
and U5343 (N_5343,N_5063,N_5131);
or U5344 (N_5344,N_5074,N_5080);
nor U5345 (N_5345,N_5106,N_5063);
and U5346 (N_5346,N_5140,N_5114);
and U5347 (N_5347,N_5035,N_5193);
nand U5348 (N_5348,N_5115,N_5068);
nand U5349 (N_5349,N_5107,N_5034);
and U5350 (N_5350,N_5048,N_5182);
xnor U5351 (N_5351,N_5069,N_5118);
or U5352 (N_5352,N_5022,N_5113);
and U5353 (N_5353,N_5165,N_5157);
and U5354 (N_5354,N_5193,N_5064);
nor U5355 (N_5355,N_5165,N_5134);
nor U5356 (N_5356,N_5184,N_5158);
nor U5357 (N_5357,N_5075,N_5162);
or U5358 (N_5358,N_5042,N_5113);
nor U5359 (N_5359,N_5042,N_5049);
xnor U5360 (N_5360,N_5013,N_5119);
nor U5361 (N_5361,N_5052,N_5180);
or U5362 (N_5362,N_5152,N_5064);
and U5363 (N_5363,N_5126,N_5069);
nor U5364 (N_5364,N_5058,N_5008);
xor U5365 (N_5365,N_5112,N_5024);
or U5366 (N_5366,N_5091,N_5176);
nand U5367 (N_5367,N_5183,N_5058);
and U5368 (N_5368,N_5023,N_5184);
and U5369 (N_5369,N_5034,N_5172);
xor U5370 (N_5370,N_5003,N_5100);
nand U5371 (N_5371,N_5010,N_5039);
or U5372 (N_5372,N_5034,N_5058);
or U5373 (N_5373,N_5094,N_5028);
nand U5374 (N_5374,N_5151,N_5069);
nor U5375 (N_5375,N_5166,N_5071);
and U5376 (N_5376,N_5173,N_5089);
nor U5377 (N_5377,N_5166,N_5043);
and U5378 (N_5378,N_5075,N_5180);
and U5379 (N_5379,N_5170,N_5142);
and U5380 (N_5380,N_5101,N_5029);
nor U5381 (N_5381,N_5133,N_5022);
and U5382 (N_5382,N_5060,N_5098);
nor U5383 (N_5383,N_5090,N_5075);
nand U5384 (N_5384,N_5080,N_5015);
nor U5385 (N_5385,N_5038,N_5188);
nand U5386 (N_5386,N_5107,N_5135);
xor U5387 (N_5387,N_5107,N_5037);
or U5388 (N_5388,N_5152,N_5016);
and U5389 (N_5389,N_5066,N_5166);
or U5390 (N_5390,N_5079,N_5108);
nor U5391 (N_5391,N_5093,N_5091);
and U5392 (N_5392,N_5099,N_5022);
nor U5393 (N_5393,N_5011,N_5055);
xnor U5394 (N_5394,N_5170,N_5076);
and U5395 (N_5395,N_5092,N_5058);
nand U5396 (N_5396,N_5171,N_5195);
and U5397 (N_5397,N_5020,N_5051);
nand U5398 (N_5398,N_5065,N_5000);
nand U5399 (N_5399,N_5123,N_5074);
or U5400 (N_5400,N_5207,N_5248);
and U5401 (N_5401,N_5283,N_5295);
nor U5402 (N_5402,N_5272,N_5377);
and U5403 (N_5403,N_5256,N_5341);
xnor U5404 (N_5404,N_5356,N_5331);
nand U5405 (N_5405,N_5355,N_5278);
nand U5406 (N_5406,N_5261,N_5378);
or U5407 (N_5407,N_5232,N_5359);
and U5408 (N_5408,N_5229,N_5345);
nand U5409 (N_5409,N_5399,N_5227);
and U5410 (N_5410,N_5326,N_5223);
xnor U5411 (N_5411,N_5205,N_5389);
nand U5412 (N_5412,N_5246,N_5307);
nand U5413 (N_5413,N_5308,N_5357);
or U5414 (N_5414,N_5323,N_5259);
and U5415 (N_5415,N_5228,N_5328);
or U5416 (N_5416,N_5215,N_5358);
nor U5417 (N_5417,N_5230,N_5234);
nor U5418 (N_5418,N_5243,N_5244);
nand U5419 (N_5419,N_5201,N_5262);
nor U5420 (N_5420,N_5263,N_5347);
nor U5421 (N_5421,N_5206,N_5382);
nor U5422 (N_5422,N_5363,N_5318);
and U5423 (N_5423,N_5216,N_5361);
nand U5424 (N_5424,N_5374,N_5375);
or U5425 (N_5425,N_5214,N_5224);
xor U5426 (N_5426,N_5366,N_5335);
xor U5427 (N_5427,N_5360,N_5371);
nor U5428 (N_5428,N_5293,N_5238);
or U5429 (N_5429,N_5280,N_5383);
xnor U5430 (N_5430,N_5219,N_5247);
or U5431 (N_5431,N_5306,N_5217);
nand U5432 (N_5432,N_5320,N_5297);
nand U5433 (N_5433,N_5364,N_5393);
nor U5434 (N_5434,N_5354,N_5202);
and U5435 (N_5435,N_5309,N_5290);
or U5436 (N_5436,N_5252,N_5314);
nor U5437 (N_5437,N_5342,N_5231);
or U5438 (N_5438,N_5332,N_5222);
nand U5439 (N_5439,N_5220,N_5316);
nand U5440 (N_5440,N_5255,N_5395);
and U5441 (N_5441,N_5233,N_5221);
nand U5442 (N_5442,N_5239,N_5250);
and U5443 (N_5443,N_5349,N_5277);
or U5444 (N_5444,N_5271,N_5373);
or U5445 (N_5445,N_5386,N_5203);
or U5446 (N_5446,N_5209,N_5264);
nor U5447 (N_5447,N_5321,N_5379);
nor U5448 (N_5448,N_5236,N_5289);
xor U5449 (N_5449,N_5284,N_5305);
and U5450 (N_5450,N_5322,N_5388);
or U5451 (N_5451,N_5267,N_5368);
and U5452 (N_5452,N_5372,N_5208);
and U5453 (N_5453,N_5212,N_5300);
or U5454 (N_5454,N_5291,N_5376);
xor U5455 (N_5455,N_5338,N_5313);
nand U5456 (N_5456,N_5294,N_5398);
or U5457 (N_5457,N_5237,N_5339);
and U5458 (N_5458,N_5310,N_5235);
or U5459 (N_5459,N_5218,N_5288);
nor U5460 (N_5460,N_5241,N_5390);
or U5461 (N_5461,N_5292,N_5275);
nor U5462 (N_5462,N_5317,N_5258);
and U5463 (N_5463,N_5242,N_5325);
nor U5464 (N_5464,N_5394,N_5269);
or U5465 (N_5465,N_5319,N_5337);
xnor U5466 (N_5466,N_5381,N_5350);
and U5467 (N_5467,N_5260,N_5298);
or U5468 (N_5468,N_5273,N_5200);
nor U5469 (N_5469,N_5226,N_5303);
nand U5470 (N_5470,N_5346,N_5340);
or U5471 (N_5471,N_5396,N_5324);
or U5472 (N_5472,N_5385,N_5365);
and U5473 (N_5473,N_5287,N_5334);
and U5474 (N_5474,N_5387,N_5352);
xor U5475 (N_5475,N_5391,N_5279);
xor U5476 (N_5476,N_5211,N_5370);
or U5477 (N_5477,N_5329,N_5344);
nor U5478 (N_5478,N_5274,N_5240);
xor U5479 (N_5479,N_5367,N_5251);
nor U5480 (N_5480,N_5380,N_5286);
or U5481 (N_5481,N_5348,N_5265);
xor U5482 (N_5482,N_5204,N_5210);
xor U5483 (N_5483,N_5384,N_5296);
nor U5484 (N_5484,N_5330,N_5225);
or U5485 (N_5485,N_5254,N_5392);
and U5486 (N_5486,N_5397,N_5362);
nor U5487 (N_5487,N_5304,N_5245);
or U5488 (N_5488,N_5343,N_5266);
and U5489 (N_5489,N_5301,N_5333);
or U5490 (N_5490,N_5253,N_5268);
xor U5491 (N_5491,N_5351,N_5336);
or U5492 (N_5492,N_5327,N_5285);
nand U5493 (N_5493,N_5249,N_5302);
nand U5494 (N_5494,N_5282,N_5281);
xnor U5495 (N_5495,N_5312,N_5276);
or U5496 (N_5496,N_5257,N_5213);
or U5497 (N_5497,N_5315,N_5311);
or U5498 (N_5498,N_5353,N_5270);
or U5499 (N_5499,N_5299,N_5369);
or U5500 (N_5500,N_5275,N_5366);
and U5501 (N_5501,N_5299,N_5315);
nand U5502 (N_5502,N_5258,N_5262);
nand U5503 (N_5503,N_5269,N_5383);
nor U5504 (N_5504,N_5242,N_5374);
or U5505 (N_5505,N_5239,N_5255);
and U5506 (N_5506,N_5386,N_5247);
nor U5507 (N_5507,N_5352,N_5381);
or U5508 (N_5508,N_5264,N_5375);
and U5509 (N_5509,N_5235,N_5399);
nor U5510 (N_5510,N_5295,N_5247);
and U5511 (N_5511,N_5228,N_5375);
or U5512 (N_5512,N_5213,N_5252);
or U5513 (N_5513,N_5268,N_5335);
nor U5514 (N_5514,N_5335,N_5367);
xor U5515 (N_5515,N_5311,N_5360);
and U5516 (N_5516,N_5211,N_5302);
nand U5517 (N_5517,N_5238,N_5351);
nand U5518 (N_5518,N_5351,N_5282);
nor U5519 (N_5519,N_5316,N_5336);
xnor U5520 (N_5520,N_5391,N_5346);
nor U5521 (N_5521,N_5261,N_5292);
nor U5522 (N_5522,N_5363,N_5229);
nor U5523 (N_5523,N_5351,N_5247);
xor U5524 (N_5524,N_5343,N_5381);
nor U5525 (N_5525,N_5394,N_5228);
nand U5526 (N_5526,N_5224,N_5215);
and U5527 (N_5527,N_5328,N_5399);
nor U5528 (N_5528,N_5347,N_5392);
nor U5529 (N_5529,N_5251,N_5364);
xor U5530 (N_5530,N_5363,N_5248);
nor U5531 (N_5531,N_5395,N_5321);
nand U5532 (N_5532,N_5257,N_5366);
or U5533 (N_5533,N_5397,N_5257);
nor U5534 (N_5534,N_5390,N_5345);
nor U5535 (N_5535,N_5338,N_5394);
or U5536 (N_5536,N_5363,N_5239);
or U5537 (N_5537,N_5293,N_5359);
or U5538 (N_5538,N_5218,N_5327);
nor U5539 (N_5539,N_5232,N_5253);
or U5540 (N_5540,N_5396,N_5212);
or U5541 (N_5541,N_5219,N_5336);
nand U5542 (N_5542,N_5399,N_5300);
xor U5543 (N_5543,N_5201,N_5325);
or U5544 (N_5544,N_5373,N_5346);
nand U5545 (N_5545,N_5370,N_5383);
and U5546 (N_5546,N_5383,N_5322);
nor U5547 (N_5547,N_5306,N_5377);
xor U5548 (N_5548,N_5341,N_5347);
nor U5549 (N_5549,N_5393,N_5354);
nand U5550 (N_5550,N_5212,N_5226);
and U5551 (N_5551,N_5342,N_5267);
or U5552 (N_5552,N_5230,N_5341);
nor U5553 (N_5553,N_5265,N_5377);
xor U5554 (N_5554,N_5305,N_5336);
nand U5555 (N_5555,N_5279,N_5323);
nor U5556 (N_5556,N_5239,N_5234);
nand U5557 (N_5557,N_5209,N_5330);
and U5558 (N_5558,N_5270,N_5378);
nor U5559 (N_5559,N_5368,N_5292);
nand U5560 (N_5560,N_5349,N_5300);
or U5561 (N_5561,N_5365,N_5268);
or U5562 (N_5562,N_5255,N_5269);
nand U5563 (N_5563,N_5296,N_5339);
nand U5564 (N_5564,N_5209,N_5366);
or U5565 (N_5565,N_5396,N_5384);
or U5566 (N_5566,N_5359,N_5285);
and U5567 (N_5567,N_5365,N_5225);
xor U5568 (N_5568,N_5392,N_5325);
nand U5569 (N_5569,N_5303,N_5387);
xor U5570 (N_5570,N_5243,N_5284);
nand U5571 (N_5571,N_5342,N_5255);
xor U5572 (N_5572,N_5298,N_5258);
xnor U5573 (N_5573,N_5260,N_5210);
and U5574 (N_5574,N_5222,N_5311);
and U5575 (N_5575,N_5203,N_5290);
nor U5576 (N_5576,N_5379,N_5242);
nand U5577 (N_5577,N_5342,N_5343);
xnor U5578 (N_5578,N_5231,N_5337);
and U5579 (N_5579,N_5276,N_5362);
xnor U5580 (N_5580,N_5265,N_5380);
nand U5581 (N_5581,N_5289,N_5287);
or U5582 (N_5582,N_5291,N_5333);
and U5583 (N_5583,N_5209,N_5358);
nand U5584 (N_5584,N_5202,N_5246);
or U5585 (N_5585,N_5294,N_5368);
xnor U5586 (N_5586,N_5399,N_5287);
nor U5587 (N_5587,N_5341,N_5311);
or U5588 (N_5588,N_5259,N_5270);
nand U5589 (N_5589,N_5323,N_5303);
nand U5590 (N_5590,N_5371,N_5304);
nor U5591 (N_5591,N_5373,N_5320);
or U5592 (N_5592,N_5382,N_5293);
or U5593 (N_5593,N_5346,N_5274);
nand U5594 (N_5594,N_5368,N_5337);
nor U5595 (N_5595,N_5200,N_5202);
nand U5596 (N_5596,N_5353,N_5254);
or U5597 (N_5597,N_5226,N_5261);
or U5598 (N_5598,N_5245,N_5312);
and U5599 (N_5599,N_5328,N_5264);
or U5600 (N_5600,N_5435,N_5434);
or U5601 (N_5601,N_5411,N_5529);
nand U5602 (N_5602,N_5452,N_5420);
nand U5603 (N_5603,N_5578,N_5559);
or U5604 (N_5604,N_5426,N_5493);
nor U5605 (N_5605,N_5568,N_5561);
or U5606 (N_5606,N_5507,N_5583);
and U5607 (N_5607,N_5488,N_5535);
nand U5608 (N_5608,N_5436,N_5525);
and U5609 (N_5609,N_5431,N_5487);
or U5610 (N_5610,N_5400,N_5503);
and U5611 (N_5611,N_5425,N_5589);
nand U5612 (N_5612,N_5497,N_5410);
nor U5613 (N_5613,N_5473,N_5586);
nand U5614 (N_5614,N_5422,N_5567);
and U5615 (N_5615,N_5536,N_5490);
and U5616 (N_5616,N_5492,N_5415);
xnor U5617 (N_5617,N_5403,N_5482);
or U5618 (N_5618,N_5484,N_5542);
nor U5619 (N_5619,N_5514,N_5527);
nand U5620 (N_5620,N_5506,N_5595);
nor U5621 (N_5621,N_5518,N_5590);
and U5622 (N_5622,N_5512,N_5458);
or U5623 (N_5623,N_5523,N_5537);
and U5624 (N_5624,N_5584,N_5448);
xor U5625 (N_5625,N_5481,N_5453);
nand U5626 (N_5626,N_5534,N_5547);
nor U5627 (N_5627,N_5580,N_5456);
or U5628 (N_5628,N_5549,N_5408);
and U5629 (N_5629,N_5418,N_5405);
and U5630 (N_5630,N_5413,N_5552);
xnor U5631 (N_5631,N_5548,N_5588);
nor U5632 (N_5632,N_5432,N_5466);
nor U5633 (N_5633,N_5558,N_5597);
or U5634 (N_5634,N_5572,N_5457);
nand U5635 (N_5635,N_5499,N_5504);
nand U5636 (N_5636,N_5433,N_5520);
xor U5637 (N_5637,N_5569,N_5599);
and U5638 (N_5638,N_5546,N_5449);
nor U5639 (N_5639,N_5511,N_5553);
nor U5640 (N_5640,N_5485,N_5424);
nor U5641 (N_5641,N_5554,N_5587);
or U5642 (N_5642,N_5563,N_5528);
and U5643 (N_5643,N_5416,N_5522);
and U5644 (N_5644,N_5469,N_5489);
nand U5645 (N_5645,N_5521,N_5519);
nand U5646 (N_5646,N_5442,N_5401);
or U5647 (N_5647,N_5510,N_5596);
nand U5648 (N_5648,N_5406,N_5429);
or U5649 (N_5649,N_5545,N_5491);
nor U5650 (N_5650,N_5474,N_5470);
nand U5651 (N_5651,N_5441,N_5508);
or U5652 (N_5652,N_5582,N_5409);
or U5653 (N_5653,N_5478,N_5476);
or U5654 (N_5654,N_5532,N_5557);
nor U5655 (N_5655,N_5496,N_5560);
nor U5656 (N_5656,N_5598,N_5550);
nand U5657 (N_5657,N_5467,N_5585);
and U5658 (N_5658,N_5501,N_5423);
xor U5659 (N_5659,N_5573,N_5459);
nor U5660 (N_5660,N_5444,N_5556);
and U5661 (N_5661,N_5575,N_5571);
nor U5662 (N_5662,N_5517,N_5570);
or U5663 (N_5663,N_5579,N_5412);
or U5664 (N_5664,N_5428,N_5464);
or U5665 (N_5665,N_5477,N_5446);
nand U5666 (N_5666,N_5454,N_5594);
and U5667 (N_5667,N_5451,N_5465);
xor U5668 (N_5668,N_5516,N_5439);
and U5669 (N_5669,N_5417,N_5515);
nand U5670 (N_5670,N_5471,N_5562);
nor U5671 (N_5671,N_5544,N_5483);
nor U5672 (N_5672,N_5502,N_5540);
and U5673 (N_5673,N_5513,N_5468);
nand U5674 (N_5674,N_5494,N_5591);
xor U5675 (N_5675,N_5566,N_5463);
or U5676 (N_5676,N_5437,N_5564);
and U5677 (N_5677,N_5565,N_5475);
nor U5678 (N_5678,N_5438,N_5593);
or U5679 (N_5679,N_5526,N_5445);
or U5680 (N_5680,N_5447,N_5524);
or U5681 (N_5681,N_5576,N_5495);
nor U5682 (N_5682,N_5505,N_5480);
or U5683 (N_5683,N_5430,N_5402);
and U5684 (N_5684,N_5479,N_5509);
nand U5685 (N_5685,N_5427,N_5462);
or U5686 (N_5686,N_5450,N_5555);
nor U5687 (N_5687,N_5500,N_5543);
nor U5688 (N_5688,N_5581,N_5443);
nand U5689 (N_5689,N_5460,N_5530);
and U5690 (N_5690,N_5498,N_5461);
nor U5691 (N_5691,N_5541,N_5455);
nand U5692 (N_5692,N_5419,N_5551);
and U5693 (N_5693,N_5533,N_5472);
nor U5694 (N_5694,N_5486,N_5404);
xnor U5695 (N_5695,N_5421,N_5592);
nand U5696 (N_5696,N_5539,N_5574);
xnor U5697 (N_5697,N_5407,N_5577);
nand U5698 (N_5698,N_5538,N_5414);
nor U5699 (N_5699,N_5440,N_5531);
xor U5700 (N_5700,N_5499,N_5584);
nor U5701 (N_5701,N_5476,N_5590);
xor U5702 (N_5702,N_5483,N_5538);
nand U5703 (N_5703,N_5535,N_5503);
nand U5704 (N_5704,N_5467,N_5599);
xor U5705 (N_5705,N_5542,N_5593);
xor U5706 (N_5706,N_5561,N_5525);
and U5707 (N_5707,N_5494,N_5558);
nand U5708 (N_5708,N_5528,N_5438);
nand U5709 (N_5709,N_5472,N_5515);
or U5710 (N_5710,N_5523,N_5585);
and U5711 (N_5711,N_5509,N_5560);
and U5712 (N_5712,N_5509,N_5448);
and U5713 (N_5713,N_5419,N_5517);
and U5714 (N_5714,N_5423,N_5431);
or U5715 (N_5715,N_5443,N_5525);
and U5716 (N_5716,N_5520,N_5486);
nand U5717 (N_5717,N_5492,N_5518);
nand U5718 (N_5718,N_5536,N_5487);
nor U5719 (N_5719,N_5543,N_5569);
or U5720 (N_5720,N_5454,N_5524);
nor U5721 (N_5721,N_5498,N_5447);
nor U5722 (N_5722,N_5554,N_5477);
nor U5723 (N_5723,N_5428,N_5484);
nor U5724 (N_5724,N_5493,N_5533);
or U5725 (N_5725,N_5528,N_5405);
or U5726 (N_5726,N_5434,N_5598);
xor U5727 (N_5727,N_5511,N_5512);
nand U5728 (N_5728,N_5566,N_5496);
and U5729 (N_5729,N_5498,N_5569);
and U5730 (N_5730,N_5466,N_5442);
or U5731 (N_5731,N_5539,N_5577);
or U5732 (N_5732,N_5598,N_5590);
or U5733 (N_5733,N_5590,N_5461);
nand U5734 (N_5734,N_5470,N_5433);
and U5735 (N_5735,N_5490,N_5455);
or U5736 (N_5736,N_5530,N_5570);
xor U5737 (N_5737,N_5487,N_5449);
nand U5738 (N_5738,N_5425,N_5559);
or U5739 (N_5739,N_5527,N_5499);
nor U5740 (N_5740,N_5512,N_5561);
or U5741 (N_5741,N_5497,N_5477);
and U5742 (N_5742,N_5445,N_5485);
nand U5743 (N_5743,N_5410,N_5458);
and U5744 (N_5744,N_5556,N_5469);
and U5745 (N_5745,N_5470,N_5594);
nor U5746 (N_5746,N_5444,N_5596);
nand U5747 (N_5747,N_5546,N_5432);
nand U5748 (N_5748,N_5562,N_5530);
nor U5749 (N_5749,N_5574,N_5444);
and U5750 (N_5750,N_5446,N_5538);
nor U5751 (N_5751,N_5558,N_5484);
xnor U5752 (N_5752,N_5478,N_5475);
xor U5753 (N_5753,N_5439,N_5451);
and U5754 (N_5754,N_5429,N_5480);
xor U5755 (N_5755,N_5409,N_5470);
xor U5756 (N_5756,N_5482,N_5546);
nor U5757 (N_5757,N_5478,N_5408);
and U5758 (N_5758,N_5522,N_5593);
nand U5759 (N_5759,N_5444,N_5515);
nand U5760 (N_5760,N_5429,N_5467);
nand U5761 (N_5761,N_5426,N_5473);
and U5762 (N_5762,N_5447,N_5491);
and U5763 (N_5763,N_5570,N_5462);
nor U5764 (N_5764,N_5532,N_5536);
nand U5765 (N_5765,N_5475,N_5515);
nand U5766 (N_5766,N_5423,N_5464);
nand U5767 (N_5767,N_5575,N_5451);
nand U5768 (N_5768,N_5416,N_5505);
or U5769 (N_5769,N_5410,N_5489);
or U5770 (N_5770,N_5465,N_5504);
or U5771 (N_5771,N_5552,N_5425);
or U5772 (N_5772,N_5441,N_5491);
nor U5773 (N_5773,N_5499,N_5538);
nand U5774 (N_5774,N_5502,N_5519);
nor U5775 (N_5775,N_5564,N_5449);
nor U5776 (N_5776,N_5534,N_5598);
and U5777 (N_5777,N_5483,N_5413);
nor U5778 (N_5778,N_5472,N_5585);
or U5779 (N_5779,N_5494,N_5472);
and U5780 (N_5780,N_5543,N_5552);
nand U5781 (N_5781,N_5485,N_5537);
nand U5782 (N_5782,N_5553,N_5509);
and U5783 (N_5783,N_5530,N_5490);
or U5784 (N_5784,N_5586,N_5493);
nand U5785 (N_5785,N_5425,N_5418);
nand U5786 (N_5786,N_5563,N_5412);
nor U5787 (N_5787,N_5463,N_5409);
nand U5788 (N_5788,N_5545,N_5409);
nor U5789 (N_5789,N_5424,N_5544);
or U5790 (N_5790,N_5585,N_5450);
or U5791 (N_5791,N_5486,N_5493);
or U5792 (N_5792,N_5594,N_5403);
or U5793 (N_5793,N_5401,N_5570);
and U5794 (N_5794,N_5411,N_5458);
or U5795 (N_5795,N_5571,N_5402);
nor U5796 (N_5796,N_5577,N_5479);
nor U5797 (N_5797,N_5429,N_5594);
or U5798 (N_5798,N_5525,N_5471);
or U5799 (N_5799,N_5447,N_5440);
xor U5800 (N_5800,N_5760,N_5765);
nand U5801 (N_5801,N_5735,N_5716);
or U5802 (N_5802,N_5781,N_5691);
and U5803 (N_5803,N_5692,N_5669);
and U5804 (N_5804,N_5699,N_5745);
or U5805 (N_5805,N_5720,N_5793);
or U5806 (N_5806,N_5618,N_5619);
or U5807 (N_5807,N_5648,N_5630);
nand U5808 (N_5808,N_5631,N_5626);
nor U5809 (N_5809,N_5732,N_5799);
nand U5810 (N_5810,N_5776,N_5796);
and U5811 (N_5811,N_5752,N_5607);
and U5812 (N_5812,N_5700,N_5647);
or U5813 (N_5813,N_5778,N_5780);
xnor U5814 (N_5814,N_5612,N_5712);
nor U5815 (N_5815,N_5623,N_5683);
nand U5816 (N_5816,N_5763,N_5670);
nor U5817 (N_5817,N_5688,N_5707);
and U5818 (N_5818,N_5746,N_5788);
nor U5819 (N_5819,N_5636,N_5655);
xor U5820 (N_5820,N_5704,N_5798);
and U5821 (N_5821,N_5654,N_5741);
or U5822 (N_5822,N_5603,N_5690);
and U5823 (N_5823,N_5650,N_5785);
or U5824 (N_5824,N_5681,N_5770);
nand U5825 (N_5825,N_5666,N_5661);
and U5826 (N_5826,N_5671,N_5621);
nor U5827 (N_5827,N_5774,N_5672);
or U5828 (N_5828,N_5701,N_5693);
nand U5829 (N_5829,N_5660,N_5769);
or U5830 (N_5830,N_5668,N_5751);
or U5831 (N_5831,N_5784,N_5729);
and U5832 (N_5832,N_5656,N_5742);
nor U5833 (N_5833,N_5719,N_5674);
or U5834 (N_5834,N_5721,N_5740);
nor U5835 (N_5835,N_5767,N_5791);
xnor U5836 (N_5836,N_5768,N_5724);
nor U5837 (N_5837,N_5676,N_5698);
nor U5838 (N_5838,N_5609,N_5675);
or U5839 (N_5839,N_5726,N_5787);
or U5840 (N_5840,N_5758,N_5628);
nand U5841 (N_5841,N_5749,N_5703);
xor U5842 (N_5842,N_5708,N_5795);
nor U5843 (N_5843,N_5715,N_5773);
nor U5844 (N_5844,N_5632,N_5757);
or U5845 (N_5845,N_5738,N_5682);
nand U5846 (N_5846,N_5622,N_5739);
or U5847 (N_5847,N_5646,N_5772);
and U5848 (N_5848,N_5652,N_5615);
nand U5849 (N_5849,N_5792,N_5734);
and U5850 (N_5850,N_5642,N_5685);
nor U5851 (N_5851,N_5737,N_5635);
or U5852 (N_5852,N_5783,N_5673);
nand U5853 (N_5853,N_5779,N_5702);
and U5854 (N_5854,N_5625,N_5633);
or U5855 (N_5855,N_5696,N_5640);
nor U5856 (N_5856,N_5736,N_5651);
nor U5857 (N_5857,N_5687,N_5717);
or U5858 (N_5858,N_5747,N_5750);
nand U5859 (N_5859,N_5748,N_5761);
nor U5860 (N_5860,N_5608,N_5727);
or U5861 (N_5861,N_5600,N_5777);
and U5862 (N_5862,N_5706,N_5602);
and U5863 (N_5863,N_5710,N_5766);
or U5864 (N_5864,N_5634,N_5718);
xnor U5865 (N_5865,N_5601,N_5677);
nor U5866 (N_5866,N_5709,N_5658);
and U5867 (N_5867,N_5753,N_5756);
nor U5868 (N_5868,N_5782,N_5762);
nor U5869 (N_5869,N_5723,N_5794);
or U5870 (N_5870,N_5733,N_5644);
and U5871 (N_5871,N_5629,N_5680);
and U5872 (N_5872,N_5725,N_5638);
or U5873 (N_5873,N_5789,N_5662);
nor U5874 (N_5874,N_5653,N_5754);
nand U5875 (N_5875,N_5667,N_5610);
or U5876 (N_5876,N_5614,N_5713);
or U5877 (N_5877,N_5722,N_5743);
nand U5878 (N_5878,N_5771,N_5606);
or U5879 (N_5879,N_5711,N_5694);
and U5880 (N_5880,N_5649,N_5665);
nand U5881 (N_5881,N_5678,N_5643);
nor U5882 (N_5882,N_5620,N_5624);
nor U5883 (N_5883,N_5705,N_5689);
or U5884 (N_5884,N_5786,N_5686);
nand U5885 (N_5885,N_5744,N_5639);
xor U5886 (N_5886,N_5790,N_5637);
nand U5887 (N_5887,N_5728,N_5679);
and U5888 (N_5888,N_5641,N_5659);
nor U5889 (N_5889,N_5605,N_5764);
and U5890 (N_5890,N_5759,N_5663);
nor U5891 (N_5891,N_5730,N_5657);
and U5892 (N_5892,N_5627,N_5604);
nor U5893 (N_5893,N_5697,N_5797);
or U5894 (N_5894,N_5684,N_5664);
or U5895 (N_5895,N_5695,N_5611);
nor U5896 (N_5896,N_5645,N_5731);
and U5897 (N_5897,N_5613,N_5755);
nor U5898 (N_5898,N_5617,N_5714);
nand U5899 (N_5899,N_5616,N_5775);
or U5900 (N_5900,N_5679,N_5683);
xnor U5901 (N_5901,N_5682,N_5692);
or U5902 (N_5902,N_5720,N_5794);
nor U5903 (N_5903,N_5649,N_5780);
nor U5904 (N_5904,N_5663,N_5792);
and U5905 (N_5905,N_5792,N_5716);
xor U5906 (N_5906,N_5646,N_5641);
xnor U5907 (N_5907,N_5656,N_5626);
and U5908 (N_5908,N_5721,N_5762);
xor U5909 (N_5909,N_5602,N_5612);
or U5910 (N_5910,N_5621,N_5718);
and U5911 (N_5911,N_5709,N_5712);
xor U5912 (N_5912,N_5768,N_5662);
or U5913 (N_5913,N_5762,N_5691);
or U5914 (N_5914,N_5794,N_5635);
nor U5915 (N_5915,N_5790,N_5737);
nor U5916 (N_5916,N_5739,N_5742);
nor U5917 (N_5917,N_5627,N_5652);
and U5918 (N_5918,N_5734,N_5771);
nor U5919 (N_5919,N_5751,N_5759);
and U5920 (N_5920,N_5659,N_5777);
or U5921 (N_5921,N_5613,N_5734);
and U5922 (N_5922,N_5665,N_5629);
or U5923 (N_5923,N_5756,N_5784);
nor U5924 (N_5924,N_5710,N_5682);
or U5925 (N_5925,N_5634,N_5626);
nor U5926 (N_5926,N_5699,N_5651);
xor U5927 (N_5927,N_5667,N_5763);
nand U5928 (N_5928,N_5779,N_5786);
or U5929 (N_5929,N_5757,N_5621);
nor U5930 (N_5930,N_5764,N_5759);
and U5931 (N_5931,N_5753,N_5674);
or U5932 (N_5932,N_5797,N_5762);
or U5933 (N_5933,N_5614,N_5643);
nand U5934 (N_5934,N_5623,N_5797);
nor U5935 (N_5935,N_5663,N_5691);
nand U5936 (N_5936,N_5757,N_5744);
and U5937 (N_5937,N_5608,N_5653);
and U5938 (N_5938,N_5646,N_5625);
or U5939 (N_5939,N_5774,N_5640);
and U5940 (N_5940,N_5671,N_5665);
and U5941 (N_5941,N_5706,N_5736);
and U5942 (N_5942,N_5608,N_5685);
xor U5943 (N_5943,N_5731,N_5749);
xor U5944 (N_5944,N_5668,N_5620);
nand U5945 (N_5945,N_5736,N_5743);
and U5946 (N_5946,N_5636,N_5777);
or U5947 (N_5947,N_5681,N_5675);
and U5948 (N_5948,N_5760,N_5690);
and U5949 (N_5949,N_5707,N_5611);
and U5950 (N_5950,N_5644,N_5601);
and U5951 (N_5951,N_5652,N_5628);
or U5952 (N_5952,N_5643,N_5651);
nand U5953 (N_5953,N_5703,N_5657);
and U5954 (N_5954,N_5789,N_5639);
xnor U5955 (N_5955,N_5796,N_5613);
or U5956 (N_5956,N_5750,N_5719);
and U5957 (N_5957,N_5757,N_5776);
nand U5958 (N_5958,N_5630,N_5704);
nor U5959 (N_5959,N_5683,N_5605);
nand U5960 (N_5960,N_5791,N_5641);
xor U5961 (N_5961,N_5645,N_5610);
and U5962 (N_5962,N_5661,N_5676);
nor U5963 (N_5963,N_5638,N_5603);
or U5964 (N_5964,N_5777,N_5637);
nor U5965 (N_5965,N_5725,N_5710);
nor U5966 (N_5966,N_5788,N_5720);
nor U5967 (N_5967,N_5703,N_5600);
nand U5968 (N_5968,N_5766,N_5605);
and U5969 (N_5969,N_5635,N_5752);
nor U5970 (N_5970,N_5747,N_5648);
nor U5971 (N_5971,N_5730,N_5746);
or U5972 (N_5972,N_5643,N_5702);
and U5973 (N_5973,N_5796,N_5761);
or U5974 (N_5974,N_5715,N_5790);
and U5975 (N_5975,N_5739,N_5687);
xor U5976 (N_5976,N_5791,N_5683);
xor U5977 (N_5977,N_5794,N_5623);
nor U5978 (N_5978,N_5654,N_5767);
nor U5979 (N_5979,N_5665,N_5788);
or U5980 (N_5980,N_5753,N_5767);
nand U5981 (N_5981,N_5676,N_5639);
and U5982 (N_5982,N_5690,N_5753);
and U5983 (N_5983,N_5673,N_5724);
and U5984 (N_5984,N_5716,N_5772);
xnor U5985 (N_5985,N_5673,N_5721);
nor U5986 (N_5986,N_5709,N_5681);
or U5987 (N_5987,N_5609,N_5711);
nand U5988 (N_5988,N_5650,N_5601);
or U5989 (N_5989,N_5648,N_5779);
nor U5990 (N_5990,N_5601,N_5636);
or U5991 (N_5991,N_5792,N_5677);
xnor U5992 (N_5992,N_5681,N_5654);
nor U5993 (N_5993,N_5798,N_5764);
nor U5994 (N_5994,N_5608,N_5738);
nor U5995 (N_5995,N_5699,N_5760);
and U5996 (N_5996,N_5729,N_5618);
nand U5997 (N_5997,N_5699,N_5662);
nor U5998 (N_5998,N_5609,N_5620);
xnor U5999 (N_5999,N_5766,N_5741);
or U6000 (N_6000,N_5844,N_5949);
or U6001 (N_6001,N_5986,N_5943);
nand U6002 (N_6002,N_5954,N_5992);
xnor U6003 (N_6003,N_5831,N_5916);
and U6004 (N_6004,N_5969,N_5937);
nand U6005 (N_6005,N_5920,N_5854);
nor U6006 (N_6006,N_5863,N_5967);
nor U6007 (N_6007,N_5883,N_5962);
or U6008 (N_6008,N_5830,N_5833);
nor U6009 (N_6009,N_5834,N_5934);
nor U6010 (N_6010,N_5936,N_5953);
nand U6011 (N_6011,N_5886,N_5930);
or U6012 (N_6012,N_5882,N_5887);
nor U6013 (N_6013,N_5956,N_5881);
or U6014 (N_6014,N_5976,N_5980);
or U6015 (N_6015,N_5957,N_5987);
nand U6016 (N_6016,N_5868,N_5919);
nor U6017 (N_6017,N_5802,N_5900);
nor U6018 (N_6018,N_5924,N_5869);
or U6019 (N_6019,N_5837,N_5932);
nand U6020 (N_6020,N_5832,N_5896);
nand U6021 (N_6021,N_5878,N_5984);
nand U6022 (N_6022,N_5893,N_5905);
xor U6023 (N_6023,N_5917,N_5996);
nor U6024 (N_6024,N_5860,N_5985);
or U6025 (N_6025,N_5885,N_5897);
or U6026 (N_6026,N_5904,N_5908);
and U6027 (N_6027,N_5861,N_5931);
or U6028 (N_6028,N_5872,N_5981);
and U6029 (N_6029,N_5983,N_5915);
or U6030 (N_6030,N_5903,N_5940);
and U6031 (N_6031,N_5907,N_5909);
xnor U6032 (N_6032,N_5906,N_5952);
nor U6033 (N_6033,N_5825,N_5978);
nand U6034 (N_6034,N_5811,N_5829);
nand U6035 (N_6035,N_5975,N_5808);
nand U6036 (N_6036,N_5828,N_5859);
nand U6037 (N_6037,N_5990,N_5911);
or U6038 (N_6038,N_5852,N_5968);
nand U6039 (N_6039,N_5815,N_5877);
or U6040 (N_6040,N_5840,N_5880);
or U6041 (N_6041,N_5855,N_5923);
and U6042 (N_6042,N_5958,N_5901);
nand U6043 (N_6043,N_5847,N_5888);
and U6044 (N_6044,N_5870,N_5827);
nor U6045 (N_6045,N_5876,N_5944);
nor U6046 (N_6046,N_5902,N_5913);
or U6047 (N_6047,N_5974,N_5850);
or U6048 (N_6048,N_5942,N_5977);
nand U6049 (N_6049,N_5822,N_5960);
nor U6050 (N_6050,N_5951,N_5812);
and U6051 (N_6051,N_5971,N_5973);
or U6052 (N_6052,N_5826,N_5889);
nor U6053 (N_6053,N_5820,N_5921);
or U6054 (N_6054,N_5864,N_5867);
and U6055 (N_6055,N_5991,N_5843);
or U6056 (N_6056,N_5899,N_5972);
or U6057 (N_6057,N_5819,N_5862);
xnor U6058 (N_6058,N_5946,N_5959);
nor U6059 (N_6059,N_5965,N_5806);
and U6060 (N_6060,N_5963,N_5925);
or U6061 (N_6061,N_5857,N_5873);
xor U6062 (N_6062,N_5851,N_5821);
or U6063 (N_6063,N_5848,N_5874);
or U6064 (N_6064,N_5966,N_5928);
or U6065 (N_6065,N_5918,N_5804);
nor U6066 (N_6066,N_5997,N_5884);
and U6067 (N_6067,N_5853,N_5818);
and U6068 (N_6068,N_5890,N_5922);
and U6069 (N_6069,N_5933,N_5964);
or U6070 (N_6070,N_5988,N_5865);
and U6071 (N_6071,N_5871,N_5935);
and U6072 (N_6072,N_5961,N_5948);
nand U6073 (N_6073,N_5817,N_5970);
and U6074 (N_6074,N_5912,N_5835);
or U6075 (N_6075,N_5982,N_5939);
nand U6076 (N_6076,N_5816,N_5910);
nand U6077 (N_6077,N_5994,N_5895);
nand U6078 (N_6078,N_5866,N_5998);
nor U6079 (N_6079,N_5824,N_5800);
nor U6080 (N_6080,N_5894,N_5813);
and U6081 (N_6081,N_5879,N_5845);
nand U6082 (N_6082,N_5945,N_5849);
or U6083 (N_6083,N_5898,N_5842);
nand U6084 (N_6084,N_5979,N_5858);
nor U6085 (N_6085,N_5989,N_5807);
nand U6086 (N_6086,N_5836,N_5814);
or U6087 (N_6087,N_5941,N_5999);
and U6088 (N_6088,N_5955,N_5995);
nand U6089 (N_6089,N_5927,N_5926);
nand U6090 (N_6090,N_5838,N_5801);
nor U6091 (N_6091,N_5891,N_5993);
nand U6092 (N_6092,N_5875,N_5950);
nand U6093 (N_6093,N_5841,N_5823);
and U6094 (N_6094,N_5810,N_5809);
nand U6095 (N_6095,N_5805,N_5947);
nor U6096 (N_6096,N_5892,N_5803);
nand U6097 (N_6097,N_5929,N_5938);
or U6098 (N_6098,N_5856,N_5914);
xnor U6099 (N_6099,N_5839,N_5846);
and U6100 (N_6100,N_5899,N_5966);
and U6101 (N_6101,N_5827,N_5866);
or U6102 (N_6102,N_5945,N_5942);
or U6103 (N_6103,N_5999,N_5826);
and U6104 (N_6104,N_5834,N_5884);
or U6105 (N_6105,N_5939,N_5951);
nor U6106 (N_6106,N_5962,N_5874);
xnor U6107 (N_6107,N_5903,N_5854);
xnor U6108 (N_6108,N_5902,N_5989);
nand U6109 (N_6109,N_5914,N_5956);
or U6110 (N_6110,N_5823,N_5807);
xnor U6111 (N_6111,N_5912,N_5983);
nor U6112 (N_6112,N_5919,N_5891);
nand U6113 (N_6113,N_5901,N_5939);
or U6114 (N_6114,N_5862,N_5827);
or U6115 (N_6115,N_5934,N_5962);
nand U6116 (N_6116,N_5811,N_5845);
or U6117 (N_6117,N_5873,N_5966);
and U6118 (N_6118,N_5811,N_5968);
or U6119 (N_6119,N_5866,N_5967);
xnor U6120 (N_6120,N_5811,N_5942);
or U6121 (N_6121,N_5972,N_5837);
nor U6122 (N_6122,N_5821,N_5965);
nand U6123 (N_6123,N_5889,N_5921);
nor U6124 (N_6124,N_5882,N_5980);
nor U6125 (N_6125,N_5840,N_5869);
xor U6126 (N_6126,N_5993,N_5995);
nor U6127 (N_6127,N_5943,N_5865);
xnor U6128 (N_6128,N_5809,N_5817);
and U6129 (N_6129,N_5905,N_5800);
nand U6130 (N_6130,N_5991,N_5900);
nor U6131 (N_6131,N_5823,N_5990);
and U6132 (N_6132,N_5824,N_5895);
or U6133 (N_6133,N_5950,N_5825);
and U6134 (N_6134,N_5961,N_5999);
and U6135 (N_6135,N_5887,N_5846);
or U6136 (N_6136,N_5903,N_5846);
xnor U6137 (N_6137,N_5983,N_5949);
and U6138 (N_6138,N_5813,N_5805);
nand U6139 (N_6139,N_5997,N_5934);
nand U6140 (N_6140,N_5861,N_5950);
and U6141 (N_6141,N_5910,N_5897);
or U6142 (N_6142,N_5803,N_5918);
and U6143 (N_6143,N_5914,N_5915);
and U6144 (N_6144,N_5957,N_5820);
or U6145 (N_6145,N_5888,N_5880);
nand U6146 (N_6146,N_5977,N_5993);
and U6147 (N_6147,N_5847,N_5981);
nand U6148 (N_6148,N_5928,N_5977);
or U6149 (N_6149,N_5991,N_5920);
nor U6150 (N_6150,N_5956,N_5863);
xnor U6151 (N_6151,N_5896,N_5909);
or U6152 (N_6152,N_5979,N_5822);
nor U6153 (N_6153,N_5881,N_5868);
xor U6154 (N_6154,N_5922,N_5999);
or U6155 (N_6155,N_5918,N_5837);
nor U6156 (N_6156,N_5872,N_5969);
or U6157 (N_6157,N_5925,N_5839);
nor U6158 (N_6158,N_5872,N_5989);
nor U6159 (N_6159,N_5844,N_5864);
or U6160 (N_6160,N_5902,N_5969);
nor U6161 (N_6161,N_5924,N_5969);
and U6162 (N_6162,N_5840,N_5872);
or U6163 (N_6163,N_5967,N_5952);
nor U6164 (N_6164,N_5956,N_5912);
or U6165 (N_6165,N_5810,N_5921);
nand U6166 (N_6166,N_5965,N_5854);
and U6167 (N_6167,N_5872,N_5937);
nand U6168 (N_6168,N_5887,N_5929);
xnor U6169 (N_6169,N_5920,N_5822);
nand U6170 (N_6170,N_5897,N_5887);
nor U6171 (N_6171,N_5984,N_5954);
or U6172 (N_6172,N_5979,N_5812);
nor U6173 (N_6173,N_5903,N_5984);
nand U6174 (N_6174,N_5920,N_5812);
and U6175 (N_6175,N_5943,N_5954);
nand U6176 (N_6176,N_5957,N_5938);
nor U6177 (N_6177,N_5857,N_5855);
and U6178 (N_6178,N_5875,N_5917);
and U6179 (N_6179,N_5946,N_5988);
nor U6180 (N_6180,N_5830,N_5939);
nand U6181 (N_6181,N_5892,N_5969);
or U6182 (N_6182,N_5987,N_5955);
xnor U6183 (N_6183,N_5885,N_5975);
and U6184 (N_6184,N_5956,N_5993);
or U6185 (N_6185,N_5836,N_5987);
nor U6186 (N_6186,N_5847,N_5983);
nor U6187 (N_6187,N_5816,N_5977);
xor U6188 (N_6188,N_5871,N_5988);
nand U6189 (N_6189,N_5925,N_5989);
xor U6190 (N_6190,N_5960,N_5845);
or U6191 (N_6191,N_5877,N_5977);
or U6192 (N_6192,N_5865,N_5861);
nand U6193 (N_6193,N_5946,N_5977);
or U6194 (N_6194,N_5839,N_5922);
and U6195 (N_6195,N_5845,N_5824);
nand U6196 (N_6196,N_5923,N_5943);
nand U6197 (N_6197,N_5928,N_5922);
nor U6198 (N_6198,N_5862,N_5857);
or U6199 (N_6199,N_5882,N_5919);
or U6200 (N_6200,N_6112,N_6013);
xor U6201 (N_6201,N_6075,N_6158);
and U6202 (N_6202,N_6019,N_6094);
and U6203 (N_6203,N_6135,N_6194);
xor U6204 (N_6204,N_6118,N_6017);
and U6205 (N_6205,N_6160,N_6035);
nor U6206 (N_6206,N_6026,N_6055);
nor U6207 (N_6207,N_6061,N_6077);
and U6208 (N_6208,N_6111,N_6159);
nor U6209 (N_6209,N_6018,N_6126);
or U6210 (N_6210,N_6009,N_6027);
nor U6211 (N_6211,N_6070,N_6151);
and U6212 (N_6212,N_6167,N_6106);
or U6213 (N_6213,N_6054,N_6191);
and U6214 (N_6214,N_6195,N_6034);
nand U6215 (N_6215,N_6095,N_6044);
nor U6216 (N_6216,N_6175,N_6028);
xor U6217 (N_6217,N_6101,N_6000);
and U6218 (N_6218,N_6108,N_6093);
or U6219 (N_6219,N_6153,N_6192);
nor U6220 (N_6220,N_6004,N_6076);
and U6221 (N_6221,N_6022,N_6138);
nand U6222 (N_6222,N_6127,N_6064);
xnor U6223 (N_6223,N_6168,N_6120);
nor U6224 (N_6224,N_6199,N_6079);
or U6225 (N_6225,N_6130,N_6186);
and U6226 (N_6226,N_6178,N_6110);
nand U6227 (N_6227,N_6050,N_6128);
nand U6228 (N_6228,N_6053,N_6190);
nand U6229 (N_6229,N_6173,N_6060);
or U6230 (N_6230,N_6176,N_6097);
nor U6231 (N_6231,N_6081,N_6072);
xnor U6232 (N_6232,N_6152,N_6136);
and U6233 (N_6233,N_6189,N_6002);
and U6234 (N_6234,N_6091,N_6031);
nor U6235 (N_6235,N_6123,N_6085);
and U6236 (N_6236,N_6051,N_6185);
nor U6237 (N_6237,N_6132,N_6144);
nor U6238 (N_6238,N_6184,N_6080);
and U6239 (N_6239,N_6150,N_6121);
nand U6240 (N_6240,N_6103,N_6179);
and U6241 (N_6241,N_6193,N_6030);
nor U6242 (N_6242,N_6043,N_6165);
nand U6243 (N_6243,N_6142,N_6041);
or U6244 (N_6244,N_6197,N_6088);
or U6245 (N_6245,N_6102,N_6032);
or U6246 (N_6246,N_6114,N_6164);
or U6247 (N_6247,N_6058,N_6001);
xor U6248 (N_6248,N_6162,N_6014);
or U6249 (N_6249,N_6147,N_6023);
or U6250 (N_6250,N_6096,N_6171);
or U6251 (N_6251,N_6090,N_6166);
nand U6252 (N_6252,N_6119,N_6078);
nor U6253 (N_6253,N_6169,N_6146);
nor U6254 (N_6254,N_6016,N_6065);
nand U6255 (N_6255,N_6122,N_6149);
and U6256 (N_6256,N_6105,N_6115);
xor U6257 (N_6257,N_6036,N_6154);
nand U6258 (N_6258,N_6145,N_6182);
nor U6259 (N_6259,N_6008,N_6015);
nand U6260 (N_6260,N_6198,N_6083);
or U6261 (N_6261,N_6048,N_6038);
or U6262 (N_6262,N_6082,N_6170);
nand U6263 (N_6263,N_6057,N_6116);
nand U6264 (N_6264,N_6117,N_6141);
and U6265 (N_6265,N_6137,N_6140);
xor U6266 (N_6266,N_6183,N_6020);
nand U6267 (N_6267,N_6039,N_6069);
xnor U6268 (N_6268,N_6133,N_6040);
or U6269 (N_6269,N_6196,N_6180);
and U6270 (N_6270,N_6047,N_6073);
nand U6271 (N_6271,N_6177,N_6187);
and U6272 (N_6272,N_6042,N_6188);
or U6273 (N_6273,N_6046,N_6157);
or U6274 (N_6274,N_6139,N_6109);
and U6275 (N_6275,N_6056,N_6163);
and U6276 (N_6276,N_6033,N_6087);
nand U6277 (N_6277,N_6007,N_6131);
nand U6278 (N_6278,N_6156,N_6005);
nand U6279 (N_6279,N_6011,N_6143);
nand U6280 (N_6280,N_6124,N_6021);
or U6281 (N_6281,N_6010,N_6174);
nor U6282 (N_6282,N_6063,N_6049);
and U6283 (N_6283,N_6107,N_6084);
or U6284 (N_6284,N_6052,N_6098);
and U6285 (N_6285,N_6100,N_6025);
and U6286 (N_6286,N_6059,N_6037);
and U6287 (N_6287,N_6125,N_6074);
nor U6288 (N_6288,N_6012,N_6092);
nand U6289 (N_6289,N_6006,N_6181);
nand U6290 (N_6290,N_6062,N_6086);
nand U6291 (N_6291,N_6099,N_6148);
or U6292 (N_6292,N_6029,N_6024);
and U6293 (N_6293,N_6161,N_6066);
and U6294 (N_6294,N_6129,N_6071);
xnor U6295 (N_6295,N_6134,N_6067);
xnor U6296 (N_6296,N_6089,N_6104);
xor U6297 (N_6297,N_6068,N_6113);
nor U6298 (N_6298,N_6155,N_6045);
and U6299 (N_6299,N_6003,N_6172);
nand U6300 (N_6300,N_6068,N_6141);
nand U6301 (N_6301,N_6018,N_6169);
nor U6302 (N_6302,N_6067,N_6001);
and U6303 (N_6303,N_6025,N_6121);
and U6304 (N_6304,N_6041,N_6124);
or U6305 (N_6305,N_6043,N_6179);
nand U6306 (N_6306,N_6180,N_6085);
nand U6307 (N_6307,N_6108,N_6078);
nand U6308 (N_6308,N_6151,N_6029);
nand U6309 (N_6309,N_6123,N_6061);
nor U6310 (N_6310,N_6068,N_6114);
and U6311 (N_6311,N_6073,N_6029);
nand U6312 (N_6312,N_6058,N_6130);
xnor U6313 (N_6313,N_6096,N_6066);
xor U6314 (N_6314,N_6127,N_6084);
or U6315 (N_6315,N_6069,N_6020);
nor U6316 (N_6316,N_6008,N_6053);
or U6317 (N_6317,N_6130,N_6015);
and U6318 (N_6318,N_6093,N_6074);
or U6319 (N_6319,N_6183,N_6058);
or U6320 (N_6320,N_6081,N_6039);
or U6321 (N_6321,N_6115,N_6081);
nand U6322 (N_6322,N_6090,N_6086);
or U6323 (N_6323,N_6127,N_6163);
xnor U6324 (N_6324,N_6044,N_6071);
nand U6325 (N_6325,N_6047,N_6046);
or U6326 (N_6326,N_6116,N_6131);
and U6327 (N_6327,N_6013,N_6000);
and U6328 (N_6328,N_6055,N_6159);
nor U6329 (N_6329,N_6120,N_6184);
nand U6330 (N_6330,N_6081,N_6182);
nand U6331 (N_6331,N_6090,N_6145);
or U6332 (N_6332,N_6056,N_6065);
or U6333 (N_6333,N_6020,N_6010);
nand U6334 (N_6334,N_6007,N_6197);
and U6335 (N_6335,N_6020,N_6152);
nand U6336 (N_6336,N_6092,N_6131);
nand U6337 (N_6337,N_6133,N_6131);
or U6338 (N_6338,N_6044,N_6175);
nand U6339 (N_6339,N_6119,N_6173);
xor U6340 (N_6340,N_6051,N_6163);
xnor U6341 (N_6341,N_6070,N_6169);
and U6342 (N_6342,N_6181,N_6137);
xor U6343 (N_6343,N_6014,N_6026);
nor U6344 (N_6344,N_6100,N_6102);
nand U6345 (N_6345,N_6024,N_6066);
and U6346 (N_6346,N_6115,N_6059);
or U6347 (N_6347,N_6137,N_6032);
or U6348 (N_6348,N_6118,N_6154);
or U6349 (N_6349,N_6091,N_6131);
or U6350 (N_6350,N_6148,N_6041);
nor U6351 (N_6351,N_6056,N_6073);
or U6352 (N_6352,N_6112,N_6162);
nand U6353 (N_6353,N_6163,N_6189);
nand U6354 (N_6354,N_6012,N_6014);
and U6355 (N_6355,N_6112,N_6066);
xnor U6356 (N_6356,N_6074,N_6170);
xor U6357 (N_6357,N_6037,N_6062);
or U6358 (N_6358,N_6184,N_6119);
and U6359 (N_6359,N_6118,N_6018);
or U6360 (N_6360,N_6065,N_6005);
nor U6361 (N_6361,N_6162,N_6089);
or U6362 (N_6362,N_6037,N_6085);
xor U6363 (N_6363,N_6048,N_6073);
and U6364 (N_6364,N_6008,N_6098);
or U6365 (N_6365,N_6166,N_6183);
nand U6366 (N_6366,N_6134,N_6032);
nor U6367 (N_6367,N_6139,N_6048);
or U6368 (N_6368,N_6126,N_6014);
or U6369 (N_6369,N_6155,N_6019);
or U6370 (N_6370,N_6140,N_6098);
and U6371 (N_6371,N_6079,N_6154);
nor U6372 (N_6372,N_6047,N_6008);
nor U6373 (N_6373,N_6103,N_6020);
and U6374 (N_6374,N_6071,N_6048);
or U6375 (N_6375,N_6111,N_6027);
nor U6376 (N_6376,N_6136,N_6014);
or U6377 (N_6377,N_6006,N_6113);
or U6378 (N_6378,N_6178,N_6002);
xor U6379 (N_6379,N_6084,N_6099);
and U6380 (N_6380,N_6173,N_6188);
and U6381 (N_6381,N_6106,N_6100);
and U6382 (N_6382,N_6175,N_6052);
nor U6383 (N_6383,N_6199,N_6180);
nor U6384 (N_6384,N_6003,N_6032);
xor U6385 (N_6385,N_6191,N_6194);
nor U6386 (N_6386,N_6189,N_6155);
nor U6387 (N_6387,N_6152,N_6038);
or U6388 (N_6388,N_6015,N_6020);
nor U6389 (N_6389,N_6138,N_6193);
or U6390 (N_6390,N_6010,N_6177);
nor U6391 (N_6391,N_6123,N_6005);
and U6392 (N_6392,N_6060,N_6165);
nand U6393 (N_6393,N_6135,N_6073);
or U6394 (N_6394,N_6111,N_6015);
nor U6395 (N_6395,N_6185,N_6183);
nor U6396 (N_6396,N_6160,N_6170);
nand U6397 (N_6397,N_6140,N_6164);
nor U6398 (N_6398,N_6010,N_6007);
nor U6399 (N_6399,N_6113,N_6066);
nor U6400 (N_6400,N_6371,N_6307);
or U6401 (N_6401,N_6380,N_6385);
and U6402 (N_6402,N_6368,N_6315);
and U6403 (N_6403,N_6340,N_6369);
nor U6404 (N_6404,N_6292,N_6324);
and U6405 (N_6405,N_6258,N_6393);
or U6406 (N_6406,N_6354,N_6257);
nand U6407 (N_6407,N_6282,N_6314);
xor U6408 (N_6408,N_6271,N_6212);
and U6409 (N_6409,N_6215,N_6364);
nor U6410 (N_6410,N_6219,N_6376);
and U6411 (N_6411,N_6217,N_6275);
nand U6412 (N_6412,N_6317,N_6254);
nor U6413 (N_6413,N_6398,N_6229);
nand U6414 (N_6414,N_6206,N_6333);
xor U6415 (N_6415,N_6350,N_6337);
xor U6416 (N_6416,N_6200,N_6331);
nor U6417 (N_6417,N_6244,N_6285);
nor U6418 (N_6418,N_6280,N_6290);
nand U6419 (N_6419,N_6230,N_6234);
nor U6420 (N_6420,N_6353,N_6309);
nor U6421 (N_6421,N_6249,N_6363);
nand U6422 (N_6422,N_6298,N_6205);
or U6423 (N_6423,N_6239,N_6281);
nor U6424 (N_6424,N_6302,N_6240);
nand U6425 (N_6425,N_6318,N_6365);
and U6426 (N_6426,N_6295,N_6387);
or U6427 (N_6427,N_6265,N_6236);
nand U6428 (N_6428,N_6359,N_6394);
and U6429 (N_6429,N_6341,N_6242);
or U6430 (N_6430,N_6381,N_6300);
or U6431 (N_6431,N_6372,N_6322);
nand U6432 (N_6432,N_6326,N_6320);
and U6433 (N_6433,N_6374,N_6276);
nor U6434 (N_6434,N_6362,N_6202);
nand U6435 (N_6435,N_6347,N_6390);
or U6436 (N_6436,N_6223,N_6349);
xnor U6437 (N_6437,N_6253,N_6266);
and U6438 (N_6438,N_6251,N_6301);
nor U6439 (N_6439,N_6283,N_6335);
nor U6440 (N_6440,N_6312,N_6308);
xor U6441 (N_6441,N_6248,N_6262);
or U6442 (N_6442,N_6222,N_6386);
and U6443 (N_6443,N_6220,N_6216);
or U6444 (N_6444,N_6210,N_6332);
or U6445 (N_6445,N_6201,N_6299);
xor U6446 (N_6446,N_6306,N_6246);
or U6447 (N_6447,N_6228,N_6218);
nor U6448 (N_6448,N_6238,N_6329);
or U6449 (N_6449,N_6392,N_6391);
nand U6450 (N_6450,N_6395,N_6310);
or U6451 (N_6451,N_6227,N_6296);
and U6452 (N_6452,N_6224,N_6334);
or U6453 (N_6453,N_6278,N_6264);
nand U6454 (N_6454,N_6336,N_6203);
or U6455 (N_6455,N_6245,N_6370);
and U6456 (N_6456,N_6346,N_6288);
nand U6457 (N_6457,N_6361,N_6382);
xnor U6458 (N_6458,N_6396,N_6297);
and U6459 (N_6459,N_6343,N_6311);
nand U6460 (N_6460,N_6232,N_6286);
xor U6461 (N_6461,N_6397,N_6367);
nor U6462 (N_6462,N_6211,N_6221);
and U6463 (N_6463,N_6399,N_6384);
nor U6464 (N_6464,N_6213,N_6304);
and U6465 (N_6465,N_6233,N_6339);
or U6466 (N_6466,N_6388,N_6268);
nand U6467 (N_6467,N_6328,N_6325);
and U6468 (N_6468,N_6208,N_6273);
nor U6469 (N_6469,N_6291,N_6204);
nand U6470 (N_6470,N_6226,N_6277);
nor U6471 (N_6471,N_6250,N_6231);
and U6472 (N_6472,N_6256,N_6261);
or U6473 (N_6473,N_6342,N_6366);
nor U6474 (N_6474,N_6293,N_6383);
and U6475 (N_6475,N_6378,N_6351);
nor U6476 (N_6476,N_6243,N_6303);
or U6477 (N_6477,N_6269,N_6345);
nand U6478 (N_6478,N_6348,N_6355);
xnor U6479 (N_6479,N_6235,N_6294);
or U6480 (N_6480,N_6289,N_6255);
nand U6481 (N_6481,N_6344,N_6321);
or U6482 (N_6482,N_6305,N_6247);
nor U6483 (N_6483,N_6375,N_6237);
xnor U6484 (N_6484,N_6252,N_6272);
xnor U6485 (N_6485,N_6316,N_6356);
xor U6486 (N_6486,N_6225,N_6313);
or U6487 (N_6487,N_6330,N_6360);
nand U6488 (N_6488,N_6214,N_6377);
and U6489 (N_6489,N_6327,N_6352);
and U6490 (N_6490,N_6274,N_6319);
or U6491 (N_6491,N_6357,N_6389);
or U6492 (N_6492,N_6279,N_6207);
nand U6493 (N_6493,N_6241,N_6284);
or U6494 (N_6494,N_6260,N_6287);
or U6495 (N_6495,N_6270,N_6358);
or U6496 (N_6496,N_6338,N_6379);
nor U6497 (N_6497,N_6373,N_6209);
nor U6498 (N_6498,N_6263,N_6323);
or U6499 (N_6499,N_6267,N_6259);
or U6500 (N_6500,N_6319,N_6391);
or U6501 (N_6501,N_6213,N_6379);
nor U6502 (N_6502,N_6240,N_6315);
and U6503 (N_6503,N_6319,N_6272);
nand U6504 (N_6504,N_6338,N_6263);
nor U6505 (N_6505,N_6348,N_6222);
or U6506 (N_6506,N_6366,N_6376);
or U6507 (N_6507,N_6267,N_6304);
xnor U6508 (N_6508,N_6305,N_6245);
nand U6509 (N_6509,N_6325,N_6370);
nor U6510 (N_6510,N_6317,N_6369);
and U6511 (N_6511,N_6258,N_6337);
nand U6512 (N_6512,N_6379,N_6301);
nand U6513 (N_6513,N_6267,N_6273);
or U6514 (N_6514,N_6265,N_6226);
and U6515 (N_6515,N_6284,N_6399);
or U6516 (N_6516,N_6334,N_6379);
xor U6517 (N_6517,N_6220,N_6269);
or U6518 (N_6518,N_6396,N_6321);
nor U6519 (N_6519,N_6367,N_6209);
nor U6520 (N_6520,N_6375,N_6320);
or U6521 (N_6521,N_6250,N_6388);
and U6522 (N_6522,N_6293,N_6347);
or U6523 (N_6523,N_6369,N_6267);
and U6524 (N_6524,N_6261,N_6372);
nor U6525 (N_6525,N_6234,N_6388);
or U6526 (N_6526,N_6241,N_6380);
or U6527 (N_6527,N_6231,N_6249);
nor U6528 (N_6528,N_6306,N_6278);
nand U6529 (N_6529,N_6340,N_6334);
nor U6530 (N_6530,N_6225,N_6290);
nand U6531 (N_6531,N_6264,N_6295);
and U6532 (N_6532,N_6246,N_6354);
nand U6533 (N_6533,N_6272,N_6221);
xor U6534 (N_6534,N_6218,N_6280);
xnor U6535 (N_6535,N_6358,N_6277);
xor U6536 (N_6536,N_6313,N_6309);
nor U6537 (N_6537,N_6248,N_6325);
and U6538 (N_6538,N_6248,N_6251);
nand U6539 (N_6539,N_6201,N_6326);
or U6540 (N_6540,N_6301,N_6398);
or U6541 (N_6541,N_6205,N_6327);
or U6542 (N_6542,N_6263,N_6216);
or U6543 (N_6543,N_6358,N_6217);
xor U6544 (N_6544,N_6340,N_6207);
and U6545 (N_6545,N_6369,N_6292);
nor U6546 (N_6546,N_6219,N_6323);
or U6547 (N_6547,N_6369,N_6259);
or U6548 (N_6548,N_6277,N_6242);
or U6549 (N_6549,N_6253,N_6259);
and U6550 (N_6550,N_6269,N_6260);
xnor U6551 (N_6551,N_6222,N_6252);
or U6552 (N_6552,N_6327,N_6337);
xnor U6553 (N_6553,N_6355,N_6235);
nor U6554 (N_6554,N_6219,N_6294);
and U6555 (N_6555,N_6235,N_6307);
nor U6556 (N_6556,N_6357,N_6296);
or U6557 (N_6557,N_6321,N_6354);
nand U6558 (N_6558,N_6207,N_6355);
xnor U6559 (N_6559,N_6294,N_6289);
and U6560 (N_6560,N_6213,N_6268);
nor U6561 (N_6561,N_6381,N_6278);
nand U6562 (N_6562,N_6339,N_6251);
xor U6563 (N_6563,N_6387,N_6315);
nand U6564 (N_6564,N_6377,N_6398);
and U6565 (N_6565,N_6265,N_6335);
xor U6566 (N_6566,N_6273,N_6233);
xor U6567 (N_6567,N_6208,N_6354);
xor U6568 (N_6568,N_6220,N_6302);
nor U6569 (N_6569,N_6328,N_6238);
xnor U6570 (N_6570,N_6259,N_6281);
nor U6571 (N_6571,N_6398,N_6321);
or U6572 (N_6572,N_6333,N_6256);
nand U6573 (N_6573,N_6270,N_6240);
and U6574 (N_6574,N_6303,N_6366);
nor U6575 (N_6575,N_6257,N_6291);
nor U6576 (N_6576,N_6332,N_6236);
xor U6577 (N_6577,N_6288,N_6381);
and U6578 (N_6578,N_6270,N_6360);
or U6579 (N_6579,N_6302,N_6260);
and U6580 (N_6580,N_6297,N_6223);
nand U6581 (N_6581,N_6235,N_6207);
nand U6582 (N_6582,N_6267,N_6297);
or U6583 (N_6583,N_6340,N_6240);
or U6584 (N_6584,N_6364,N_6230);
and U6585 (N_6585,N_6212,N_6370);
and U6586 (N_6586,N_6213,N_6218);
or U6587 (N_6587,N_6262,N_6276);
nand U6588 (N_6588,N_6201,N_6203);
xor U6589 (N_6589,N_6268,N_6217);
nand U6590 (N_6590,N_6237,N_6338);
or U6591 (N_6591,N_6259,N_6289);
or U6592 (N_6592,N_6215,N_6272);
nor U6593 (N_6593,N_6392,N_6261);
xor U6594 (N_6594,N_6331,N_6317);
nor U6595 (N_6595,N_6243,N_6330);
or U6596 (N_6596,N_6250,N_6253);
xnor U6597 (N_6597,N_6272,N_6237);
and U6598 (N_6598,N_6320,N_6386);
and U6599 (N_6599,N_6226,N_6325);
or U6600 (N_6600,N_6521,N_6401);
nand U6601 (N_6601,N_6512,N_6449);
and U6602 (N_6602,N_6487,N_6404);
nor U6603 (N_6603,N_6540,N_6410);
nand U6604 (N_6604,N_6571,N_6480);
or U6605 (N_6605,N_6585,N_6425);
and U6606 (N_6606,N_6453,N_6447);
nor U6607 (N_6607,N_6539,N_6586);
nand U6608 (N_6608,N_6541,N_6436);
nand U6609 (N_6609,N_6456,N_6478);
or U6610 (N_6610,N_6488,N_6444);
nor U6611 (N_6611,N_6473,N_6483);
xor U6612 (N_6612,N_6424,N_6454);
or U6613 (N_6613,N_6426,N_6467);
nor U6614 (N_6614,N_6529,N_6402);
and U6615 (N_6615,N_6418,N_6505);
nand U6616 (N_6616,N_6591,N_6500);
nor U6617 (N_6617,N_6552,N_6573);
nand U6618 (N_6618,N_6497,N_6469);
and U6619 (N_6619,N_6545,N_6550);
nor U6620 (N_6620,N_6577,N_6407);
nand U6621 (N_6621,N_6531,N_6493);
nand U6622 (N_6622,N_6459,N_6440);
nor U6623 (N_6623,N_6414,N_6455);
and U6624 (N_6624,N_6406,N_6439);
nor U6625 (N_6625,N_6594,N_6518);
or U6626 (N_6626,N_6504,N_6429);
or U6627 (N_6627,N_6448,N_6522);
nor U6628 (N_6628,N_6560,N_6567);
or U6629 (N_6629,N_6554,N_6432);
and U6630 (N_6630,N_6547,N_6598);
nor U6631 (N_6631,N_6462,N_6514);
or U6632 (N_6632,N_6517,N_6451);
or U6633 (N_6633,N_6470,N_6437);
nor U6634 (N_6634,N_6513,N_6568);
and U6635 (N_6635,N_6544,N_6533);
or U6636 (N_6636,N_6492,N_6403);
and U6637 (N_6637,N_6419,N_6572);
or U6638 (N_6638,N_6475,N_6490);
nor U6639 (N_6639,N_6408,N_6570);
nor U6640 (N_6640,N_6515,N_6535);
nand U6641 (N_6641,N_6576,N_6468);
nor U6642 (N_6642,N_6536,N_6516);
or U6643 (N_6643,N_6489,N_6564);
or U6644 (N_6644,N_6430,N_6460);
and U6645 (N_6645,N_6509,N_6481);
nand U6646 (N_6646,N_6413,N_6421);
or U6647 (N_6647,N_6511,N_6443);
and U6648 (N_6648,N_6428,N_6485);
and U6649 (N_6649,N_6441,N_6530);
nor U6650 (N_6650,N_6415,N_6476);
nand U6651 (N_6651,N_6555,N_6581);
nand U6652 (N_6652,N_6528,N_6546);
nand U6653 (N_6653,N_6534,N_6596);
nor U6654 (N_6654,N_6538,N_6597);
nor U6655 (N_6655,N_6486,N_6508);
xor U6656 (N_6656,N_6558,N_6543);
and U6657 (N_6657,N_6434,N_6556);
nand U6658 (N_6658,N_6464,N_6400);
or U6659 (N_6659,N_6563,N_6471);
or U6660 (N_6660,N_6506,N_6507);
nor U6661 (N_6661,N_6501,N_6435);
or U6662 (N_6662,N_6433,N_6412);
nor U6663 (N_6663,N_6450,N_6431);
nand U6664 (N_6664,N_6491,N_6599);
nand U6665 (N_6665,N_6519,N_6474);
or U6666 (N_6666,N_6405,N_6463);
xnor U6667 (N_6667,N_6502,N_6446);
and U6668 (N_6668,N_6565,N_6498);
and U6669 (N_6669,N_6582,N_6542);
and U6670 (N_6670,N_6575,N_6482);
nor U6671 (N_6671,N_6562,N_6549);
or U6672 (N_6672,N_6445,N_6579);
nand U6673 (N_6673,N_6574,N_6561);
nand U6674 (N_6674,N_6411,N_6589);
and U6675 (N_6675,N_6495,N_6525);
nor U6676 (N_6676,N_6527,N_6422);
and U6677 (N_6677,N_6420,N_6524);
nand U6678 (N_6678,N_6496,N_6466);
and U6679 (N_6679,N_6442,N_6417);
and U6680 (N_6680,N_6457,N_6588);
and U6681 (N_6681,N_6569,N_6472);
or U6682 (N_6682,N_6499,N_6438);
xnor U6683 (N_6683,N_6583,N_6503);
or U6684 (N_6684,N_6510,N_6553);
or U6685 (N_6685,N_6477,N_6578);
xnor U6686 (N_6686,N_6494,N_6584);
nor U6687 (N_6687,N_6551,N_6523);
or U6688 (N_6688,N_6590,N_6537);
or U6689 (N_6689,N_6409,N_6484);
and U6690 (N_6690,N_6592,N_6580);
or U6691 (N_6691,N_6427,N_6520);
and U6692 (N_6692,N_6479,N_6593);
and U6693 (N_6693,N_6595,N_6452);
nor U6694 (N_6694,N_6559,N_6548);
and U6695 (N_6695,N_6557,N_6465);
nand U6696 (N_6696,N_6532,N_6458);
nand U6697 (N_6697,N_6461,N_6566);
nand U6698 (N_6698,N_6423,N_6526);
nand U6699 (N_6699,N_6587,N_6416);
nand U6700 (N_6700,N_6495,N_6502);
nand U6701 (N_6701,N_6562,N_6593);
nand U6702 (N_6702,N_6402,N_6423);
nor U6703 (N_6703,N_6516,N_6510);
nand U6704 (N_6704,N_6462,N_6579);
or U6705 (N_6705,N_6437,N_6587);
nor U6706 (N_6706,N_6512,N_6470);
xnor U6707 (N_6707,N_6581,N_6455);
or U6708 (N_6708,N_6547,N_6585);
nor U6709 (N_6709,N_6508,N_6586);
or U6710 (N_6710,N_6422,N_6572);
and U6711 (N_6711,N_6448,N_6573);
xor U6712 (N_6712,N_6566,N_6588);
nand U6713 (N_6713,N_6582,N_6527);
nand U6714 (N_6714,N_6544,N_6449);
and U6715 (N_6715,N_6468,N_6465);
or U6716 (N_6716,N_6469,N_6580);
and U6717 (N_6717,N_6439,N_6502);
nor U6718 (N_6718,N_6566,N_6451);
and U6719 (N_6719,N_6534,N_6496);
nor U6720 (N_6720,N_6512,N_6565);
and U6721 (N_6721,N_6485,N_6476);
xor U6722 (N_6722,N_6540,N_6430);
nor U6723 (N_6723,N_6467,N_6529);
or U6724 (N_6724,N_6550,N_6464);
or U6725 (N_6725,N_6589,N_6568);
nor U6726 (N_6726,N_6527,N_6419);
nand U6727 (N_6727,N_6574,N_6467);
nor U6728 (N_6728,N_6571,N_6507);
xnor U6729 (N_6729,N_6409,N_6433);
and U6730 (N_6730,N_6437,N_6436);
nor U6731 (N_6731,N_6581,N_6425);
nor U6732 (N_6732,N_6515,N_6593);
nand U6733 (N_6733,N_6485,N_6545);
nor U6734 (N_6734,N_6462,N_6561);
nand U6735 (N_6735,N_6590,N_6404);
and U6736 (N_6736,N_6541,N_6560);
and U6737 (N_6737,N_6493,N_6452);
or U6738 (N_6738,N_6431,N_6557);
or U6739 (N_6739,N_6436,N_6473);
nand U6740 (N_6740,N_6565,N_6462);
or U6741 (N_6741,N_6516,N_6532);
and U6742 (N_6742,N_6588,N_6444);
and U6743 (N_6743,N_6587,N_6577);
nor U6744 (N_6744,N_6456,N_6423);
xor U6745 (N_6745,N_6449,N_6542);
nor U6746 (N_6746,N_6554,N_6551);
nand U6747 (N_6747,N_6466,N_6502);
nor U6748 (N_6748,N_6554,N_6473);
nand U6749 (N_6749,N_6514,N_6585);
nand U6750 (N_6750,N_6479,N_6528);
nand U6751 (N_6751,N_6569,N_6521);
nor U6752 (N_6752,N_6543,N_6549);
or U6753 (N_6753,N_6475,N_6569);
nand U6754 (N_6754,N_6541,N_6536);
nor U6755 (N_6755,N_6510,N_6519);
and U6756 (N_6756,N_6566,N_6520);
and U6757 (N_6757,N_6539,N_6427);
nor U6758 (N_6758,N_6480,N_6478);
and U6759 (N_6759,N_6416,N_6536);
and U6760 (N_6760,N_6418,N_6499);
nor U6761 (N_6761,N_6457,N_6570);
xnor U6762 (N_6762,N_6447,N_6425);
or U6763 (N_6763,N_6574,N_6420);
or U6764 (N_6764,N_6516,N_6442);
or U6765 (N_6765,N_6524,N_6530);
and U6766 (N_6766,N_6488,N_6514);
and U6767 (N_6767,N_6570,N_6517);
nor U6768 (N_6768,N_6421,N_6554);
nor U6769 (N_6769,N_6479,N_6561);
nand U6770 (N_6770,N_6521,N_6420);
and U6771 (N_6771,N_6486,N_6454);
and U6772 (N_6772,N_6508,N_6460);
and U6773 (N_6773,N_6552,N_6562);
nand U6774 (N_6774,N_6425,N_6504);
and U6775 (N_6775,N_6428,N_6527);
nand U6776 (N_6776,N_6479,N_6526);
nor U6777 (N_6777,N_6586,N_6457);
nor U6778 (N_6778,N_6409,N_6592);
or U6779 (N_6779,N_6454,N_6529);
or U6780 (N_6780,N_6543,N_6417);
and U6781 (N_6781,N_6519,N_6408);
xnor U6782 (N_6782,N_6498,N_6484);
nand U6783 (N_6783,N_6489,N_6415);
and U6784 (N_6784,N_6543,N_6452);
xor U6785 (N_6785,N_6487,N_6576);
nand U6786 (N_6786,N_6444,N_6409);
or U6787 (N_6787,N_6450,N_6477);
or U6788 (N_6788,N_6410,N_6429);
nand U6789 (N_6789,N_6575,N_6409);
xnor U6790 (N_6790,N_6456,N_6400);
nor U6791 (N_6791,N_6459,N_6586);
nand U6792 (N_6792,N_6467,N_6573);
and U6793 (N_6793,N_6452,N_6517);
xor U6794 (N_6794,N_6537,N_6492);
nor U6795 (N_6795,N_6444,N_6441);
and U6796 (N_6796,N_6438,N_6526);
nor U6797 (N_6797,N_6550,N_6425);
nand U6798 (N_6798,N_6436,N_6435);
nand U6799 (N_6799,N_6574,N_6548);
nor U6800 (N_6800,N_6652,N_6702);
or U6801 (N_6801,N_6760,N_6694);
nand U6802 (N_6802,N_6755,N_6769);
nor U6803 (N_6803,N_6637,N_6780);
nand U6804 (N_6804,N_6645,N_6748);
nor U6805 (N_6805,N_6624,N_6794);
and U6806 (N_6806,N_6677,N_6703);
nor U6807 (N_6807,N_6697,N_6707);
nand U6808 (N_6808,N_6632,N_6753);
and U6809 (N_6809,N_6715,N_6732);
and U6810 (N_6810,N_6616,N_6785);
or U6811 (N_6811,N_6681,N_6695);
nand U6812 (N_6812,N_6669,N_6743);
and U6813 (N_6813,N_6655,N_6754);
or U6814 (N_6814,N_6604,N_6670);
nand U6815 (N_6815,N_6619,N_6767);
nand U6816 (N_6816,N_6724,N_6607);
nand U6817 (N_6817,N_6706,N_6720);
and U6818 (N_6818,N_6602,N_6723);
nand U6819 (N_6819,N_6745,N_6691);
and U6820 (N_6820,N_6777,N_6644);
nand U6821 (N_6821,N_6678,N_6718);
nor U6822 (N_6822,N_6689,N_6609);
nand U6823 (N_6823,N_6698,N_6658);
or U6824 (N_6824,N_6662,N_6630);
and U6825 (N_6825,N_6742,N_6731);
nand U6826 (N_6826,N_6699,N_6640);
nor U6827 (N_6827,N_6727,N_6617);
and U6828 (N_6828,N_6618,N_6651);
or U6829 (N_6829,N_6711,N_6773);
and U6830 (N_6830,N_6749,N_6759);
nor U6831 (N_6831,N_6710,N_6659);
nor U6832 (N_6832,N_6735,N_6763);
nand U6833 (N_6833,N_6793,N_6775);
nor U6834 (N_6834,N_6601,N_6721);
and U6835 (N_6835,N_6643,N_6782);
nor U6836 (N_6836,N_6653,N_6730);
xnor U6837 (N_6837,N_6642,N_6622);
and U6838 (N_6838,N_6791,N_6781);
or U6839 (N_6839,N_6668,N_6631);
nand U6840 (N_6840,N_6674,N_6722);
nand U6841 (N_6841,N_6633,N_6686);
nand U6842 (N_6842,N_6679,N_6747);
or U6843 (N_6843,N_6627,N_6704);
or U6844 (N_6844,N_6746,N_6744);
nand U6845 (N_6845,N_6621,N_6614);
nor U6846 (N_6846,N_6673,N_6600);
and U6847 (N_6847,N_6661,N_6638);
nand U6848 (N_6848,N_6650,N_6737);
and U6849 (N_6849,N_6740,N_6615);
or U6850 (N_6850,N_6714,N_6636);
nand U6851 (N_6851,N_6776,N_6639);
or U6852 (N_6852,N_6774,N_6738);
or U6853 (N_6853,N_6693,N_6770);
or U6854 (N_6854,N_6716,N_6797);
and U6855 (N_6855,N_6603,N_6717);
and U6856 (N_6856,N_6733,N_6647);
and U6857 (N_6857,N_6729,N_6708);
and U6858 (N_6858,N_6783,N_6613);
and U6859 (N_6859,N_6726,N_6682);
and U6860 (N_6860,N_6771,N_6758);
xor U6861 (N_6861,N_6709,N_6750);
nor U6862 (N_6862,N_6646,N_6795);
nand U6863 (N_6863,N_6656,N_6687);
or U6864 (N_6864,N_6765,N_6696);
and U6865 (N_6865,N_6685,N_6611);
nor U6866 (N_6866,N_6728,N_6665);
nand U6867 (N_6867,N_6788,N_6768);
nand U6868 (N_6868,N_6736,N_6734);
nor U6869 (N_6869,N_6798,N_6700);
and U6870 (N_6870,N_6756,N_6787);
nor U6871 (N_6871,N_6666,N_6641);
or U6872 (N_6872,N_6751,N_6684);
xor U6873 (N_6873,N_6626,N_6725);
or U6874 (N_6874,N_6792,N_6649);
nand U6875 (N_6875,N_6690,N_6676);
or U6876 (N_6876,N_6796,N_6784);
nor U6877 (N_6877,N_6623,N_6635);
xor U6878 (N_6878,N_6608,N_6790);
nand U6879 (N_6879,N_6772,N_6789);
or U6880 (N_6880,N_6692,N_6683);
or U6881 (N_6881,N_6663,N_6766);
and U6882 (N_6882,N_6680,N_6705);
and U6883 (N_6883,N_6712,N_6628);
nand U6884 (N_6884,N_6620,N_6648);
nand U6885 (N_6885,N_6660,N_6713);
or U6886 (N_6886,N_6761,N_6606);
and U6887 (N_6887,N_6757,N_6752);
and U6888 (N_6888,N_6786,N_6612);
nor U6889 (N_6889,N_6667,N_6762);
and U6890 (N_6890,N_6779,N_6625);
or U6891 (N_6891,N_6672,N_6629);
nand U6892 (N_6892,N_6764,N_6605);
nand U6893 (N_6893,N_6675,N_6657);
and U6894 (N_6894,N_6671,N_6741);
nor U6895 (N_6895,N_6664,N_6701);
nand U6896 (N_6896,N_6688,N_6719);
and U6897 (N_6897,N_6778,N_6654);
or U6898 (N_6898,N_6739,N_6634);
nand U6899 (N_6899,N_6799,N_6610);
nand U6900 (N_6900,N_6658,N_6682);
or U6901 (N_6901,N_6708,N_6794);
xor U6902 (N_6902,N_6773,N_6653);
and U6903 (N_6903,N_6712,N_6608);
or U6904 (N_6904,N_6710,N_6706);
nor U6905 (N_6905,N_6639,N_6789);
or U6906 (N_6906,N_6760,N_6705);
nand U6907 (N_6907,N_6714,N_6795);
xor U6908 (N_6908,N_6698,N_6608);
or U6909 (N_6909,N_6619,N_6616);
xnor U6910 (N_6910,N_6691,N_6767);
nand U6911 (N_6911,N_6676,N_6706);
or U6912 (N_6912,N_6689,N_6665);
nor U6913 (N_6913,N_6691,N_6617);
and U6914 (N_6914,N_6650,N_6628);
nand U6915 (N_6915,N_6684,N_6678);
and U6916 (N_6916,N_6791,N_6722);
and U6917 (N_6917,N_6651,N_6602);
nor U6918 (N_6918,N_6667,N_6681);
nand U6919 (N_6919,N_6770,N_6744);
xnor U6920 (N_6920,N_6631,N_6636);
or U6921 (N_6921,N_6646,N_6715);
nor U6922 (N_6922,N_6629,N_6715);
or U6923 (N_6923,N_6618,N_6740);
xnor U6924 (N_6924,N_6641,N_6734);
and U6925 (N_6925,N_6649,N_6602);
nand U6926 (N_6926,N_6784,N_6772);
and U6927 (N_6927,N_6770,N_6761);
and U6928 (N_6928,N_6744,N_6700);
nor U6929 (N_6929,N_6704,N_6623);
or U6930 (N_6930,N_6723,N_6765);
xor U6931 (N_6931,N_6673,N_6780);
xnor U6932 (N_6932,N_6707,N_6797);
or U6933 (N_6933,N_6743,N_6691);
or U6934 (N_6934,N_6620,N_6639);
and U6935 (N_6935,N_6614,N_6722);
nand U6936 (N_6936,N_6675,N_6724);
nor U6937 (N_6937,N_6764,N_6750);
and U6938 (N_6938,N_6779,N_6773);
nand U6939 (N_6939,N_6691,N_6703);
or U6940 (N_6940,N_6791,N_6636);
xnor U6941 (N_6941,N_6768,N_6758);
nand U6942 (N_6942,N_6664,N_6658);
nor U6943 (N_6943,N_6621,N_6644);
nor U6944 (N_6944,N_6608,N_6615);
and U6945 (N_6945,N_6755,N_6759);
nor U6946 (N_6946,N_6755,N_6735);
nand U6947 (N_6947,N_6774,N_6739);
nand U6948 (N_6948,N_6645,N_6730);
xnor U6949 (N_6949,N_6764,N_6627);
nor U6950 (N_6950,N_6728,N_6623);
nand U6951 (N_6951,N_6780,N_6764);
or U6952 (N_6952,N_6784,N_6617);
and U6953 (N_6953,N_6686,N_6663);
or U6954 (N_6954,N_6766,N_6673);
and U6955 (N_6955,N_6681,N_6701);
or U6956 (N_6956,N_6774,N_6735);
and U6957 (N_6957,N_6689,N_6765);
or U6958 (N_6958,N_6628,N_6748);
or U6959 (N_6959,N_6736,N_6705);
nor U6960 (N_6960,N_6632,N_6792);
or U6961 (N_6961,N_6678,N_6782);
or U6962 (N_6962,N_6741,N_6712);
and U6963 (N_6963,N_6604,N_6699);
nand U6964 (N_6964,N_6669,N_6709);
nor U6965 (N_6965,N_6746,N_6704);
nor U6966 (N_6966,N_6796,N_6702);
nand U6967 (N_6967,N_6767,N_6785);
nand U6968 (N_6968,N_6728,N_6771);
or U6969 (N_6969,N_6610,N_6795);
or U6970 (N_6970,N_6733,N_6600);
nor U6971 (N_6971,N_6767,N_6751);
nand U6972 (N_6972,N_6657,N_6654);
and U6973 (N_6973,N_6770,N_6692);
nor U6974 (N_6974,N_6747,N_6652);
nor U6975 (N_6975,N_6606,N_6742);
and U6976 (N_6976,N_6712,N_6690);
nand U6977 (N_6977,N_6639,N_6645);
and U6978 (N_6978,N_6767,N_6739);
nand U6979 (N_6979,N_6625,N_6644);
nor U6980 (N_6980,N_6715,N_6687);
nand U6981 (N_6981,N_6791,N_6729);
nand U6982 (N_6982,N_6695,N_6610);
nand U6983 (N_6983,N_6761,N_6631);
nor U6984 (N_6984,N_6668,N_6618);
nand U6985 (N_6985,N_6696,N_6656);
and U6986 (N_6986,N_6734,N_6780);
or U6987 (N_6987,N_6760,N_6726);
nor U6988 (N_6988,N_6716,N_6631);
and U6989 (N_6989,N_6778,N_6685);
or U6990 (N_6990,N_6783,N_6775);
or U6991 (N_6991,N_6687,N_6757);
nor U6992 (N_6992,N_6715,N_6640);
xor U6993 (N_6993,N_6766,N_6652);
or U6994 (N_6994,N_6774,N_6713);
nor U6995 (N_6995,N_6757,N_6692);
and U6996 (N_6996,N_6785,N_6733);
and U6997 (N_6997,N_6771,N_6703);
and U6998 (N_6998,N_6722,N_6679);
and U6999 (N_6999,N_6765,N_6789);
and U7000 (N_7000,N_6933,N_6852);
and U7001 (N_7001,N_6866,N_6984);
nor U7002 (N_7002,N_6966,N_6974);
nand U7003 (N_7003,N_6897,N_6952);
or U7004 (N_7004,N_6929,N_6905);
nand U7005 (N_7005,N_6987,N_6881);
nand U7006 (N_7006,N_6926,N_6802);
or U7007 (N_7007,N_6873,N_6836);
or U7008 (N_7008,N_6908,N_6997);
nor U7009 (N_7009,N_6972,N_6869);
nor U7010 (N_7010,N_6875,N_6843);
nor U7011 (N_7011,N_6943,N_6989);
or U7012 (N_7012,N_6932,N_6892);
xnor U7013 (N_7013,N_6807,N_6857);
and U7014 (N_7014,N_6982,N_6870);
nor U7015 (N_7015,N_6887,N_6898);
nand U7016 (N_7016,N_6981,N_6941);
or U7017 (N_7017,N_6853,N_6900);
nor U7018 (N_7018,N_6819,N_6928);
and U7019 (N_7019,N_6842,N_6803);
nor U7020 (N_7020,N_6838,N_6823);
nand U7021 (N_7021,N_6874,N_6922);
xnor U7022 (N_7022,N_6812,N_6851);
nor U7023 (N_7023,N_6890,N_6940);
or U7024 (N_7024,N_6994,N_6855);
or U7025 (N_7025,N_6945,N_6828);
nor U7026 (N_7026,N_6862,N_6831);
or U7027 (N_7027,N_6957,N_6854);
nand U7028 (N_7028,N_6814,N_6833);
nand U7029 (N_7029,N_6899,N_6906);
nor U7030 (N_7030,N_6985,N_6834);
and U7031 (N_7031,N_6930,N_6979);
or U7032 (N_7032,N_6811,N_6888);
xnor U7033 (N_7033,N_6889,N_6924);
and U7034 (N_7034,N_6856,N_6968);
nand U7035 (N_7035,N_6992,N_6969);
and U7036 (N_7036,N_6810,N_6849);
nand U7037 (N_7037,N_6965,N_6931);
nand U7038 (N_7038,N_6885,N_6896);
xor U7039 (N_7039,N_6953,N_6850);
nand U7040 (N_7040,N_6872,N_6996);
or U7041 (N_7041,N_6827,N_6805);
and U7042 (N_7042,N_6914,N_6806);
xnor U7043 (N_7043,N_6884,N_6944);
and U7044 (N_7044,N_6871,N_6882);
nor U7045 (N_7045,N_6858,N_6835);
nand U7046 (N_7046,N_6848,N_6891);
and U7047 (N_7047,N_6917,N_6859);
or U7048 (N_7048,N_6956,N_6864);
nor U7049 (N_7049,N_6936,N_6955);
nand U7050 (N_7050,N_6967,N_6877);
xor U7051 (N_7051,N_6977,N_6947);
or U7052 (N_7052,N_6837,N_6867);
and U7053 (N_7053,N_6949,N_6844);
nor U7054 (N_7054,N_6970,N_6880);
or U7055 (N_7055,N_6841,N_6993);
or U7056 (N_7056,N_6948,N_6845);
or U7057 (N_7057,N_6911,N_6920);
nand U7058 (N_7058,N_6907,N_6904);
nor U7059 (N_7059,N_6808,N_6815);
nor U7060 (N_7060,N_6818,N_6801);
or U7061 (N_7061,N_6962,N_6895);
and U7062 (N_7062,N_6826,N_6951);
and U7063 (N_7063,N_6804,N_6916);
and U7064 (N_7064,N_6991,N_6942);
or U7065 (N_7065,N_6937,N_6986);
nor U7066 (N_7066,N_6865,N_6902);
xor U7067 (N_7067,N_6813,N_6910);
nor U7068 (N_7068,N_6923,N_6868);
nor U7069 (N_7069,N_6839,N_6950);
or U7070 (N_7070,N_6976,N_6903);
nand U7071 (N_7071,N_6958,N_6961);
nand U7072 (N_7072,N_6861,N_6988);
and U7073 (N_7073,N_6830,N_6846);
and U7074 (N_7074,N_6840,N_6800);
nand U7075 (N_7075,N_6954,N_6939);
or U7076 (N_7076,N_6817,N_6816);
nand U7077 (N_7077,N_6925,N_6894);
or U7078 (N_7078,N_6971,N_6963);
xnor U7079 (N_7079,N_6978,N_6822);
nor U7080 (N_7080,N_6915,N_6934);
nor U7081 (N_7081,N_6964,N_6878);
xnor U7082 (N_7082,N_6995,N_6909);
xnor U7083 (N_7083,N_6935,N_6847);
and U7084 (N_7084,N_6959,N_6809);
and U7085 (N_7085,N_6927,N_6921);
and U7086 (N_7086,N_6825,N_6879);
or U7087 (N_7087,N_6829,N_6919);
and U7088 (N_7088,N_6999,N_6901);
nor U7089 (N_7089,N_6946,N_6913);
nand U7090 (N_7090,N_6990,N_6980);
nor U7091 (N_7091,N_6876,N_6883);
or U7092 (N_7092,N_6983,N_6973);
and U7093 (N_7093,N_6820,N_6886);
nor U7094 (N_7094,N_6912,N_6960);
nor U7095 (N_7095,N_6863,N_6998);
nor U7096 (N_7096,N_6821,N_6832);
or U7097 (N_7097,N_6918,N_6938);
nor U7098 (N_7098,N_6860,N_6975);
nor U7099 (N_7099,N_6824,N_6893);
nor U7100 (N_7100,N_6850,N_6915);
and U7101 (N_7101,N_6993,N_6930);
or U7102 (N_7102,N_6943,N_6825);
or U7103 (N_7103,N_6843,N_6833);
nor U7104 (N_7104,N_6905,N_6981);
xnor U7105 (N_7105,N_6916,N_6986);
nand U7106 (N_7106,N_6898,N_6914);
and U7107 (N_7107,N_6850,N_6913);
and U7108 (N_7108,N_6822,N_6852);
and U7109 (N_7109,N_6858,N_6874);
nand U7110 (N_7110,N_6949,N_6898);
or U7111 (N_7111,N_6828,N_6950);
and U7112 (N_7112,N_6982,N_6850);
and U7113 (N_7113,N_6869,N_6929);
or U7114 (N_7114,N_6845,N_6931);
or U7115 (N_7115,N_6834,N_6994);
nor U7116 (N_7116,N_6848,N_6860);
nand U7117 (N_7117,N_6951,N_6890);
nor U7118 (N_7118,N_6806,N_6822);
nand U7119 (N_7119,N_6836,N_6963);
and U7120 (N_7120,N_6854,N_6838);
nor U7121 (N_7121,N_6954,N_6999);
nand U7122 (N_7122,N_6825,N_6819);
nand U7123 (N_7123,N_6938,N_6990);
nand U7124 (N_7124,N_6871,N_6962);
nand U7125 (N_7125,N_6891,N_6896);
or U7126 (N_7126,N_6942,N_6826);
nor U7127 (N_7127,N_6819,N_6907);
nand U7128 (N_7128,N_6810,N_6934);
nor U7129 (N_7129,N_6810,N_6899);
nor U7130 (N_7130,N_6925,N_6959);
nor U7131 (N_7131,N_6954,N_6981);
xor U7132 (N_7132,N_6942,N_6960);
or U7133 (N_7133,N_6901,N_6973);
nor U7134 (N_7134,N_6834,N_6840);
and U7135 (N_7135,N_6885,N_6878);
nand U7136 (N_7136,N_6924,N_6969);
xor U7137 (N_7137,N_6992,N_6944);
or U7138 (N_7138,N_6891,N_6998);
and U7139 (N_7139,N_6970,N_6922);
and U7140 (N_7140,N_6908,N_6823);
nand U7141 (N_7141,N_6842,N_6801);
nand U7142 (N_7142,N_6831,N_6863);
nor U7143 (N_7143,N_6810,N_6996);
and U7144 (N_7144,N_6971,N_6857);
xnor U7145 (N_7145,N_6980,N_6987);
or U7146 (N_7146,N_6939,N_6995);
and U7147 (N_7147,N_6941,N_6800);
and U7148 (N_7148,N_6960,N_6990);
and U7149 (N_7149,N_6883,N_6845);
nor U7150 (N_7150,N_6987,N_6853);
xnor U7151 (N_7151,N_6841,N_6888);
nor U7152 (N_7152,N_6990,N_6914);
or U7153 (N_7153,N_6811,N_6849);
nand U7154 (N_7154,N_6845,N_6983);
or U7155 (N_7155,N_6859,N_6977);
and U7156 (N_7156,N_6982,N_6981);
nor U7157 (N_7157,N_6839,N_6801);
nor U7158 (N_7158,N_6859,N_6903);
nand U7159 (N_7159,N_6806,N_6865);
nor U7160 (N_7160,N_6993,N_6939);
nand U7161 (N_7161,N_6945,N_6888);
nand U7162 (N_7162,N_6989,N_6909);
or U7163 (N_7163,N_6860,N_6928);
and U7164 (N_7164,N_6866,N_6948);
or U7165 (N_7165,N_6836,N_6834);
and U7166 (N_7166,N_6820,N_6892);
nand U7167 (N_7167,N_6896,N_6955);
and U7168 (N_7168,N_6986,N_6855);
nor U7169 (N_7169,N_6800,N_6822);
nor U7170 (N_7170,N_6810,N_6815);
and U7171 (N_7171,N_6996,N_6935);
and U7172 (N_7172,N_6868,N_6900);
nor U7173 (N_7173,N_6900,N_6908);
or U7174 (N_7174,N_6815,N_6872);
xor U7175 (N_7175,N_6949,N_6899);
nand U7176 (N_7176,N_6878,N_6899);
nand U7177 (N_7177,N_6968,N_6999);
or U7178 (N_7178,N_6839,N_6911);
nor U7179 (N_7179,N_6835,N_6941);
nand U7180 (N_7180,N_6804,N_6952);
or U7181 (N_7181,N_6961,N_6897);
and U7182 (N_7182,N_6927,N_6968);
nand U7183 (N_7183,N_6948,N_6978);
nand U7184 (N_7184,N_6816,N_6981);
nand U7185 (N_7185,N_6981,N_6817);
and U7186 (N_7186,N_6879,N_6925);
nand U7187 (N_7187,N_6885,N_6866);
and U7188 (N_7188,N_6820,N_6993);
and U7189 (N_7189,N_6993,N_6833);
xor U7190 (N_7190,N_6891,N_6890);
xnor U7191 (N_7191,N_6944,N_6923);
xnor U7192 (N_7192,N_6861,N_6897);
xnor U7193 (N_7193,N_6800,N_6934);
and U7194 (N_7194,N_6945,N_6906);
or U7195 (N_7195,N_6802,N_6852);
nor U7196 (N_7196,N_6917,N_6998);
or U7197 (N_7197,N_6899,N_6821);
or U7198 (N_7198,N_6873,N_6904);
and U7199 (N_7199,N_6822,N_6932);
nor U7200 (N_7200,N_7173,N_7134);
and U7201 (N_7201,N_7120,N_7090);
or U7202 (N_7202,N_7130,N_7060);
or U7203 (N_7203,N_7071,N_7153);
nor U7204 (N_7204,N_7026,N_7199);
and U7205 (N_7205,N_7020,N_7183);
and U7206 (N_7206,N_7049,N_7172);
xnor U7207 (N_7207,N_7063,N_7073);
nor U7208 (N_7208,N_7150,N_7149);
nand U7209 (N_7209,N_7121,N_7167);
and U7210 (N_7210,N_7054,N_7115);
and U7211 (N_7211,N_7089,N_7044);
and U7212 (N_7212,N_7087,N_7059);
nor U7213 (N_7213,N_7056,N_7021);
and U7214 (N_7214,N_7097,N_7031);
or U7215 (N_7215,N_7076,N_7040);
nor U7216 (N_7216,N_7064,N_7003);
nand U7217 (N_7217,N_7085,N_7123);
nor U7218 (N_7218,N_7142,N_7039);
or U7219 (N_7219,N_7010,N_7161);
nand U7220 (N_7220,N_7111,N_7081);
xor U7221 (N_7221,N_7198,N_7112);
nand U7222 (N_7222,N_7058,N_7029);
or U7223 (N_7223,N_7037,N_7061);
nand U7224 (N_7224,N_7125,N_7051);
or U7225 (N_7225,N_7147,N_7146);
or U7226 (N_7226,N_7138,N_7067);
nand U7227 (N_7227,N_7139,N_7107);
and U7228 (N_7228,N_7065,N_7100);
nand U7229 (N_7229,N_7177,N_7022);
nor U7230 (N_7230,N_7116,N_7184);
xor U7231 (N_7231,N_7109,N_7050);
nand U7232 (N_7232,N_7160,N_7137);
or U7233 (N_7233,N_7195,N_7178);
and U7234 (N_7234,N_7118,N_7091);
or U7235 (N_7235,N_7086,N_7175);
or U7236 (N_7236,N_7028,N_7001);
nor U7237 (N_7237,N_7135,N_7093);
nand U7238 (N_7238,N_7144,N_7033);
nor U7239 (N_7239,N_7114,N_7075);
nor U7240 (N_7240,N_7154,N_7008);
xnor U7241 (N_7241,N_7038,N_7053);
and U7242 (N_7242,N_7155,N_7068);
xnor U7243 (N_7243,N_7131,N_7062);
or U7244 (N_7244,N_7048,N_7084);
and U7245 (N_7245,N_7152,N_7192);
or U7246 (N_7246,N_7196,N_7126);
or U7247 (N_7247,N_7069,N_7129);
or U7248 (N_7248,N_7019,N_7074);
or U7249 (N_7249,N_7043,N_7151);
nand U7250 (N_7250,N_7124,N_7136);
or U7251 (N_7251,N_7018,N_7077);
or U7252 (N_7252,N_7055,N_7009);
nand U7253 (N_7253,N_7042,N_7013);
and U7254 (N_7254,N_7148,N_7041);
nor U7255 (N_7255,N_7141,N_7176);
nor U7256 (N_7256,N_7095,N_7108);
and U7257 (N_7257,N_7005,N_7023);
nand U7258 (N_7258,N_7163,N_7104);
nand U7259 (N_7259,N_7000,N_7015);
nand U7260 (N_7260,N_7016,N_7078);
or U7261 (N_7261,N_7159,N_7004);
nand U7262 (N_7262,N_7162,N_7165);
and U7263 (N_7263,N_7186,N_7185);
xnor U7264 (N_7264,N_7174,N_7194);
nor U7265 (N_7265,N_7007,N_7158);
nor U7266 (N_7266,N_7113,N_7024);
nand U7267 (N_7267,N_7170,N_7046);
and U7268 (N_7268,N_7017,N_7182);
nor U7269 (N_7269,N_7101,N_7080);
nand U7270 (N_7270,N_7197,N_7143);
and U7271 (N_7271,N_7190,N_7094);
nor U7272 (N_7272,N_7187,N_7070);
and U7273 (N_7273,N_7096,N_7025);
nand U7274 (N_7274,N_7191,N_7128);
nand U7275 (N_7275,N_7132,N_7032);
nand U7276 (N_7276,N_7157,N_7066);
nor U7277 (N_7277,N_7188,N_7156);
nand U7278 (N_7278,N_7140,N_7180);
or U7279 (N_7279,N_7171,N_7027);
nand U7280 (N_7280,N_7168,N_7006);
and U7281 (N_7281,N_7088,N_7164);
and U7282 (N_7282,N_7047,N_7181);
and U7283 (N_7283,N_7110,N_7102);
or U7284 (N_7284,N_7103,N_7169);
nor U7285 (N_7285,N_7014,N_7133);
nand U7286 (N_7286,N_7105,N_7045);
and U7287 (N_7287,N_7030,N_7179);
nand U7288 (N_7288,N_7034,N_7011);
nor U7289 (N_7289,N_7083,N_7035);
xor U7290 (N_7290,N_7057,N_7052);
or U7291 (N_7291,N_7122,N_7127);
xnor U7292 (N_7292,N_7036,N_7012);
nand U7293 (N_7293,N_7002,N_7072);
or U7294 (N_7294,N_7166,N_7119);
and U7295 (N_7295,N_7106,N_7079);
or U7296 (N_7296,N_7189,N_7092);
xor U7297 (N_7297,N_7082,N_7098);
or U7298 (N_7298,N_7193,N_7099);
nor U7299 (N_7299,N_7117,N_7145);
nor U7300 (N_7300,N_7047,N_7149);
or U7301 (N_7301,N_7014,N_7146);
or U7302 (N_7302,N_7192,N_7059);
nand U7303 (N_7303,N_7061,N_7079);
xnor U7304 (N_7304,N_7004,N_7142);
and U7305 (N_7305,N_7067,N_7036);
nor U7306 (N_7306,N_7013,N_7090);
nor U7307 (N_7307,N_7120,N_7181);
or U7308 (N_7308,N_7006,N_7042);
or U7309 (N_7309,N_7109,N_7055);
nand U7310 (N_7310,N_7129,N_7189);
and U7311 (N_7311,N_7059,N_7161);
and U7312 (N_7312,N_7183,N_7012);
nor U7313 (N_7313,N_7069,N_7070);
xnor U7314 (N_7314,N_7016,N_7004);
nor U7315 (N_7315,N_7090,N_7102);
and U7316 (N_7316,N_7083,N_7118);
or U7317 (N_7317,N_7046,N_7163);
and U7318 (N_7318,N_7199,N_7158);
xor U7319 (N_7319,N_7036,N_7169);
and U7320 (N_7320,N_7195,N_7189);
and U7321 (N_7321,N_7092,N_7008);
nor U7322 (N_7322,N_7071,N_7015);
or U7323 (N_7323,N_7132,N_7053);
xor U7324 (N_7324,N_7182,N_7020);
and U7325 (N_7325,N_7132,N_7176);
or U7326 (N_7326,N_7186,N_7111);
or U7327 (N_7327,N_7179,N_7019);
or U7328 (N_7328,N_7096,N_7137);
and U7329 (N_7329,N_7013,N_7040);
or U7330 (N_7330,N_7041,N_7177);
nor U7331 (N_7331,N_7131,N_7172);
and U7332 (N_7332,N_7101,N_7097);
nand U7333 (N_7333,N_7132,N_7013);
nand U7334 (N_7334,N_7142,N_7092);
nand U7335 (N_7335,N_7094,N_7087);
nor U7336 (N_7336,N_7186,N_7198);
nand U7337 (N_7337,N_7134,N_7043);
xnor U7338 (N_7338,N_7014,N_7137);
nor U7339 (N_7339,N_7165,N_7134);
nand U7340 (N_7340,N_7174,N_7140);
nand U7341 (N_7341,N_7094,N_7027);
and U7342 (N_7342,N_7010,N_7129);
and U7343 (N_7343,N_7161,N_7056);
nand U7344 (N_7344,N_7141,N_7063);
nor U7345 (N_7345,N_7044,N_7029);
and U7346 (N_7346,N_7031,N_7024);
and U7347 (N_7347,N_7004,N_7165);
or U7348 (N_7348,N_7087,N_7052);
nand U7349 (N_7349,N_7131,N_7103);
xor U7350 (N_7350,N_7189,N_7085);
or U7351 (N_7351,N_7188,N_7079);
nor U7352 (N_7352,N_7190,N_7000);
nand U7353 (N_7353,N_7077,N_7199);
and U7354 (N_7354,N_7171,N_7084);
nor U7355 (N_7355,N_7026,N_7191);
and U7356 (N_7356,N_7092,N_7084);
or U7357 (N_7357,N_7163,N_7120);
and U7358 (N_7358,N_7001,N_7032);
nor U7359 (N_7359,N_7155,N_7122);
xnor U7360 (N_7360,N_7066,N_7015);
nor U7361 (N_7361,N_7012,N_7116);
nand U7362 (N_7362,N_7098,N_7103);
nor U7363 (N_7363,N_7024,N_7105);
nor U7364 (N_7364,N_7111,N_7097);
or U7365 (N_7365,N_7002,N_7190);
or U7366 (N_7366,N_7170,N_7017);
and U7367 (N_7367,N_7122,N_7147);
or U7368 (N_7368,N_7145,N_7022);
and U7369 (N_7369,N_7198,N_7085);
nor U7370 (N_7370,N_7150,N_7133);
nor U7371 (N_7371,N_7043,N_7176);
or U7372 (N_7372,N_7165,N_7065);
or U7373 (N_7373,N_7096,N_7001);
nor U7374 (N_7374,N_7142,N_7099);
and U7375 (N_7375,N_7109,N_7059);
nand U7376 (N_7376,N_7093,N_7126);
and U7377 (N_7377,N_7172,N_7119);
nand U7378 (N_7378,N_7096,N_7014);
nor U7379 (N_7379,N_7025,N_7038);
and U7380 (N_7380,N_7182,N_7025);
xnor U7381 (N_7381,N_7132,N_7172);
nor U7382 (N_7382,N_7013,N_7136);
xor U7383 (N_7383,N_7199,N_7168);
and U7384 (N_7384,N_7106,N_7190);
and U7385 (N_7385,N_7195,N_7155);
and U7386 (N_7386,N_7011,N_7092);
or U7387 (N_7387,N_7100,N_7118);
and U7388 (N_7388,N_7026,N_7101);
xnor U7389 (N_7389,N_7055,N_7019);
xor U7390 (N_7390,N_7125,N_7073);
and U7391 (N_7391,N_7105,N_7120);
and U7392 (N_7392,N_7076,N_7191);
or U7393 (N_7393,N_7186,N_7071);
and U7394 (N_7394,N_7108,N_7190);
xor U7395 (N_7395,N_7100,N_7148);
nand U7396 (N_7396,N_7025,N_7185);
nand U7397 (N_7397,N_7015,N_7031);
or U7398 (N_7398,N_7060,N_7169);
and U7399 (N_7399,N_7051,N_7022);
xor U7400 (N_7400,N_7395,N_7252);
or U7401 (N_7401,N_7243,N_7345);
or U7402 (N_7402,N_7256,N_7202);
nand U7403 (N_7403,N_7232,N_7367);
nor U7404 (N_7404,N_7330,N_7348);
and U7405 (N_7405,N_7351,N_7397);
nor U7406 (N_7406,N_7249,N_7304);
or U7407 (N_7407,N_7390,N_7388);
or U7408 (N_7408,N_7372,N_7343);
nand U7409 (N_7409,N_7214,N_7242);
nand U7410 (N_7410,N_7258,N_7262);
xor U7411 (N_7411,N_7282,N_7327);
and U7412 (N_7412,N_7361,N_7329);
nor U7413 (N_7413,N_7350,N_7230);
nand U7414 (N_7414,N_7245,N_7339);
nor U7415 (N_7415,N_7307,N_7385);
or U7416 (N_7416,N_7324,N_7200);
and U7417 (N_7417,N_7320,N_7222);
or U7418 (N_7418,N_7254,N_7284);
nand U7419 (N_7419,N_7301,N_7399);
nor U7420 (N_7420,N_7267,N_7346);
nor U7421 (N_7421,N_7318,N_7341);
and U7422 (N_7422,N_7208,N_7263);
or U7423 (N_7423,N_7279,N_7357);
or U7424 (N_7424,N_7360,N_7336);
nand U7425 (N_7425,N_7277,N_7261);
nand U7426 (N_7426,N_7280,N_7212);
or U7427 (N_7427,N_7389,N_7270);
or U7428 (N_7428,N_7364,N_7334);
nand U7429 (N_7429,N_7325,N_7305);
or U7430 (N_7430,N_7313,N_7323);
or U7431 (N_7431,N_7275,N_7228);
or U7432 (N_7432,N_7237,N_7347);
or U7433 (N_7433,N_7315,N_7306);
and U7434 (N_7434,N_7335,N_7290);
or U7435 (N_7435,N_7303,N_7294);
and U7436 (N_7436,N_7209,N_7268);
nor U7437 (N_7437,N_7331,N_7226);
and U7438 (N_7438,N_7308,N_7251);
or U7439 (N_7439,N_7260,N_7356);
and U7440 (N_7440,N_7373,N_7281);
nand U7441 (N_7441,N_7398,N_7238);
and U7442 (N_7442,N_7394,N_7312);
or U7443 (N_7443,N_7358,N_7241);
nand U7444 (N_7444,N_7297,N_7298);
nor U7445 (N_7445,N_7381,N_7382);
or U7446 (N_7446,N_7366,N_7264);
and U7447 (N_7447,N_7362,N_7219);
nand U7448 (N_7448,N_7393,N_7266);
nor U7449 (N_7449,N_7383,N_7338);
xnor U7450 (N_7450,N_7310,N_7291);
xor U7451 (N_7451,N_7231,N_7253);
nand U7452 (N_7452,N_7218,N_7234);
nor U7453 (N_7453,N_7326,N_7201);
or U7454 (N_7454,N_7283,N_7371);
nand U7455 (N_7455,N_7272,N_7309);
and U7456 (N_7456,N_7288,N_7299);
nand U7457 (N_7457,N_7375,N_7206);
and U7458 (N_7458,N_7207,N_7225);
and U7459 (N_7459,N_7380,N_7352);
nor U7460 (N_7460,N_7392,N_7365);
or U7461 (N_7461,N_7235,N_7316);
nand U7462 (N_7462,N_7227,N_7257);
and U7463 (N_7463,N_7205,N_7217);
nand U7464 (N_7464,N_7379,N_7319);
nand U7465 (N_7465,N_7293,N_7376);
and U7466 (N_7466,N_7224,N_7285);
nor U7467 (N_7467,N_7387,N_7370);
and U7468 (N_7468,N_7354,N_7378);
xor U7469 (N_7469,N_7273,N_7344);
or U7470 (N_7470,N_7384,N_7216);
nand U7471 (N_7471,N_7233,N_7322);
xnor U7472 (N_7472,N_7321,N_7374);
nor U7473 (N_7473,N_7215,N_7289);
or U7474 (N_7474,N_7340,N_7342);
or U7475 (N_7475,N_7287,N_7278);
or U7476 (N_7476,N_7244,N_7302);
or U7477 (N_7477,N_7391,N_7349);
nand U7478 (N_7478,N_7210,N_7274);
xnor U7479 (N_7479,N_7236,N_7213);
and U7480 (N_7480,N_7296,N_7259);
and U7481 (N_7481,N_7265,N_7332);
nor U7482 (N_7482,N_7221,N_7203);
or U7483 (N_7483,N_7246,N_7353);
and U7484 (N_7484,N_7271,N_7368);
nand U7485 (N_7485,N_7223,N_7328);
xnor U7486 (N_7486,N_7333,N_7295);
and U7487 (N_7487,N_7250,N_7311);
and U7488 (N_7488,N_7276,N_7292);
nand U7489 (N_7489,N_7314,N_7355);
and U7490 (N_7490,N_7255,N_7386);
and U7491 (N_7491,N_7220,N_7337);
nand U7492 (N_7492,N_7239,N_7377);
nor U7493 (N_7493,N_7317,N_7363);
nand U7494 (N_7494,N_7286,N_7300);
and U7495 (N_7495,N_7396,N_7269);
nand U7496 (N_7496,N_7229,N_7211);
and U7497 (N_7497,N_7240,N_7247);
and U7498 (N_7498,N_7359,N_7369);
and U7499 (N_7499,N_7204,N_7248);
nand U7500 (N_7500,N_7385,N_7227);
or U7501 (N_7501,N_7382,N_7306);
and U7502 (N_7502,N_7276,N_7380);
or U7503 (N_7503,N_7204,N_7330);
or U7504 (N_7504,N_7380,N_7325);
and U7505 (N_7505,N_7222,N_7302);
nor U7506 (N_7506,N_7390,N_7378);
nor U7507 (N_7507,N_7260,N_7391);
or U7508 (N_7508,N_7392,N_7257);
or U7509 (N_7509,N_7374,N_7339);
nor U7510 (N_7510,N_7219,N_7359);
or U7511 (N_7511,N_7387,N_7272);
nor U7512 (N_7512,N_7212,N_7291);
nand U7513 (N_7513,N_7236,N_7235);
and U7514 (N_7514,N_7264,N_7207);
and U7515 (N_7515,N_7376,N_7349);
or U7516 (N_7516,N_7288,N_7220);
nand U7517 (N_7517,N_7376,N_7310);
and U7518 (N_7518,N_7391,N_7229);
and U7519 (N_7519,N_7284,N_7268);
or U7520 (N_7520,N_7326,N_7363);
nor U7521 (N_7521,N_7211,N_7261);
or U7522 (N_7522,N_7346,N_7316);
nor U7523 (N_7523,N_7310,N_7211);
nor U7524 (N_7524,N_7269,N_7392);
and U7525 (N_7525,N_7365,N_7327);
xor U7526 (N_7526,N_7282,N_7298);
xnor U7527 (N_7527,N_7372,N_7291);
xnor U7528 (N_7528,N_7283,N_7205);
nand U7529 (N_7529,N_7276,N_7395);
nand U7530 (N_7530,N_7276,N_7259);
nand U7531 (N_7531,N_7341,N_7245);
or U7532 (N_7532,N_7267,N_7247);
nor U7533 (N_7533,N_7222,N_7207);
nand U7534 (N_7534,N_7215,N_7353);
nand U7535 (N_7535,N_7287,N_7391);
xnor U7536 (N_7536,N_7282,N_7200);
and U7537 (N_7537,N_7385,N_7279);
nand U7538 (N_7538,N_7366,N_7203);
nand U7539 (N_7539,N_7307,N_7322);
and U7540 (N_7540,N_7376,N_7281);
nor U7541 (N_7541,N_7231,N_7242);
or U7542 (N_7542,N_7333,N_7200);
nor U7543 (N_7543,N_7386,N_7245);
or U7544 (N_7544,N_7207,N_7236);
nor U7545 (N_7545,N_7299,N_7334);
or U7546 (N_7546,N_7324,N_7348);
nand U7547 (N_7547,N_7272,N_7210);
nor U7548 (N_7548,N_7391,N_7269);
and U7549 (N_7549,N_7245,N_7205);
or U7550 (N_7550,N_7371,N_7369);
xor U7551 (N_7551,N_7316,N_7374);
nand U7552 (N_7552,N_7259,N_7324);
nand U7553 (N_7553,N_7254,N_7343);
and U7554 (N_7554,N_7287,N_7353);
xnor U7555 (N_7555,N_7286,N_7389);
or U7556 (N_7556,N_7350,N_7390);
nor U7557 (N_7557,N_7305,N_7238);
nor U7558 (N_7558,N_7330,N_7243);
xor U7559 (N_7559,N_7346,N_7310);
nor U7560 (N_7560,N_7270,N_7395);
nand U7561 (N_7561,N_7304,N_7265);
xnor U7562 (N_7562,N_7229,N_7293);
or U7563 (N_7563,N_7325,N_7373);
xor U7564 (N_7564,N_7311,N_7276);
nor U7565 (N_7565,N_7339,N_7284);
or U7566 (N_7566,N_7265,N_7212);
and U7567 (N_7567,N_7305,N_7377);
nor U7568 (N_7568,N_7309,N_7335);
nand U7569 (N_7569,N_7316,N_7370);
nor U7570 (N_7570,N_7376,N_7246);
or U7571 (N_7571,N_7367,N_7248);
and U7572 (N_7572,N_7260,N_7230);
or U7573 (N_7573,N_7362,N_7360);
nor U7574 (N_7574,N_7249,N_7262);
and U7575 (N_7575,N_7348,N_7375);
and U7576 (N_7576,N_7330,N_7340);
nand U7577 (N_7577,N_7385,N_7309);
or U7578 (N_7578,N_7257,N_7354);
nand U7579 (N_7579,N_7323,N_7229);
nor U7580 (N_7580,N_7220,N_7261);
nor U7581 (N_7581,N_7209,N_7318);
and U7582 (N_7582,N_7241,N_7349);
and U7583 (N_7583,N_7261,N_7278);
nor U7584 (N_7584,N_7371,N_7236);
or U7585 (N_7585,N_7222,N_7339);
xnor U7586 (N_7586,N_7290,N_7209);
or U7587 (N_7587,N_7317,N_7259);
nor U7588 (N_7588,N_7374,N_7330);
or U7589 (N_7589,N_7318,N_7202);
xnor U7590 (N_7590,N_7343,N_7202);
nand U7591 (N_7591,N_7316,N_7283);
or U7592 (N_7592,N_7237,N_7303);
nand U7593 (N_7593,N_7293,N_7385);
xnor U7594 (N_7594,N_7280,N_7399);
xnor U7595 (N_7595,N_7301,N_7318);
and U7596 (N_7596,N_7379,N_7337);
nor U7597 (N_7597,N_7338,N_7201);
and U7598 (N_7598,N_7259,N_7267);
and U7599 (N_7599,N_7296,N_7394);
or U7600 (N_7600,N_7494,N_7489);
xnor U7601 (N_7601,N_7443,N_7560);
nor U7602 (N_7602,N_7552,N_7536);
nand U7603 (N_7603,N_7546,N_7408);
nor U7604 (N_7604,N_7400,N_7428);
nor U7605 (N_7605,N_7592,N_7468);
nor U7606 (N_7606,N_7455,N_7557);
or U7607 (N_7607,N_7480,N_7532);
or U7608 (N_7608,N_7487,N_7451);
nor U7609 (N_7609,N_7527,N_7572);
and U7610 (N_7610,N_7598,N_7472);
nand U7611 (N_7611,N_7515,N_7407);
and U7612 (N_7612,N_7485,N_7435);
and U7613 (N_7613,N_7461,N_7488);
nor U7614 (N_7614,N_7475,N_7594);
nand U7615 (N_7615,N_7433,N_7492);
and U7616 (N_7616,N_7458,N_7574);
and U7617 (N_7617,N_7464,N_7459);
and U7618 (N_7618,N_7550,N_7521);
and U7619 (N_7619,N_7440,N_7434);
nand U7620 (N_7620,N_7441,N_7448);
and U7621 (N_7621,N_7576,N_7577);
nand U7622 (N_7622,N_7409,N_7497);
and U7623 (N_7623,N_7418,N_7549);
nand U7624 (N_7624,N_7539,N_7582);
and U7625 (N_7625,N_7584,N_7562);
xnor U7626 (N_7626,N_7529,N_7477);
or U7627 (N_7627,N_7419,N_7450);
nand U7628 (N_7628,N_7482,N_7597);
nor U7629 (N_7629,N_7474,N_7495);
nor U7630 (N_7630,N_7411,N_7432);
and U7631 (N_7631,N_7438,N_7462);
and U7632 (N_7632,N_7523,N_7454);
or U7633 (N_7633,N_7504,N_7535);
nor U7634 (N_7634,N_7556,N_7564);
nor U7635 (N_7635,N_7514,N_7404);
xor U7636 (N_7636,N_7561,N_7573);
nor U7637 (N_7637,N_7402,N_7406);
or U7638 (N_7638,N_7509,N_7412);
xor U7639 (N_7639,N_7421,N_7534);
xnor U7640 (N_7640,N_7569,N_7442);
nand U7641 (N_7641,N_7566,N_7479);
nor U7642 (N_7642,N_7586,N_7568);
nand U7643 (N_7643,N_7538,N_7583);
nor U7644 (N_7644,N_7465,N_7496);
nand U7645 (N_7645,N_7498,N_7415);
or U7646 (N_7646,N_7429,N_7500);
or U7647 (N_7647,N_7427,N_7518);
nand U7648 (N_7648,N_7571,N_7512);
nand U7649 (N_7649,N_7519,N_7516);
nor U7650 (N_7650,N_7444,N_7491);
and U7651 (N_7651,N_7417,N_7528);
and U7652 (N_7652,N_7548,N_7416);
nor U7653 (N_7653,N_7525,N_7445);
or U7654 (N_7654,N_7547,N_7587);
or U7655 (N_7655,N_7467,N_7414);
and U7656 (N_7656,N_7478,N_7542);
or U7657 (N_7657,N_7531,N_7511);
and U7658 (N_7658,N_7508,N_7540);
nor U7659 (N_7659,N_7555,N_7581);
and U7660 (N_7660,N_7589,N_7503);
or U7661 (N_7661,N_7513,N_7520);
or U7662 (N_7662,N_7570,N_7460);
and U7663 (N_7663,N_7410,N_7524);
nor U7664 (N_7664,N_7483,N_7431);
or U7665 (N_7665,N_7558,N_7575);
xor U7666 (N_7666,N_7473,N_7426);
or U7667 (N_7667,N_7490,N_7522);
nor U7668 (N_7668,N_7551,N_7413);
nand U7669 (N_7669,N_7510,N_7502);
nand U7670 (N_7670,N_7424,N_7563);
and U7671 (N_7671,N_7526,N_7437);
nor U7672 (N_7672,N_7423,N_7567);
nor U7673 (N_7673,N_7590,N_7541);
and U7674 (N_7674,N_7446,N_7466);
xnor U7675 (N_7675,N_7585,N_7470);
and U7676 (N_7676,N_7507,N_7505);
nand U7677 (N_7677,N_7457,N_7599);
and U7678 (N_7678,N_7544,N_7506);
nor U7679 (N_7679,N_7493,N_7486);
nand U7680 (N_7680,N_7452,N_7501);
and U7681 (N_7681,N_7553,N_7554);
or U7682 (N_7682,N_7543,N_7481);
nor U7683 (N_7683,N_7565,N_7545);
nand U7684 (N_7684,N_7593,N_7579);
and U7685 (N_7685,N_7559,N_7578);
or U7686 (N_7686,N_7517,N_7499);
nand U7687 (N_7687,N_7401,N_7580);
nor U7688 (N_7688,N_7484,N_7591);
or U7689 (N_7689,N_7422,N_7463);
and U7690 (N_7690,N_7456,N_7430);
or U7691 (N_7691,N_7476,N_7595);
and U7692 (N_7692,N_7425,N_7471);
nand U7693 (N_7693,N_7588,N_7533);
nor U7694 (N_7694,N_7403,N_7596);
or U7695 (N_7695,N_7530,N_7537);
nor U7696 (N_7696,N_7449,N_7447);
or U7697 (N_7697,N_7420,N_7439);
and U7698 (N_7698,N_7469,N_7405);
and U7699 (N_7699,N_7453,N_7436);
nand U7700 (N_7700,N_7588,N_7560);
nand U7701 (N_7701,N_7533,N_7474);
and U7702 (N_7702,N_7570,N_7505);
nor U7703 (N_7703,N_7516,N_7561);
or U7704 (N_7704,N_7571,N_7464);
nand U7705 (N_7705,N_7483,N_7569);
nand U7706 (N_7706,N_7487,N_7404);
nand U7707 (N_7707,N_7486,N_7472);
or U7708 (N_7708,N_7534,N_7462);
nand U7709 (N_7709,N_7443,N_7513);
or U7710 (N_7710,N_7518,N_7510);
and U7711 (N_7711,N_7462,N_7543);
xor U7712 (N_7712,N_7546,N_7499);
and U7713 (N_7713,N_7482,N_7544);
nor U7714 (N_7714,N_7476,N_7515);
nand U7715 (N_7715,N_7592,N_7513);
and U7716 (N_7716,N_7544,N_7522);
nand U7717 (N_7717,N_7503,N_7597);
nor U7718 (N_7718,N_7503,N_7439);
xor U7719 (N_7719,N_7478,N_7432);
nor U7720 (N_7720,N_7538,N_7400);
nor U7721 (N_7721,N_7513,N_7420);
nand U7722 (N_7722,N_7547,N_7403);
and U7723 (N_7723,N_7455,N_7482);
nor U7724 (N_7724,N_7405,N_7482);
and U7725 (N_7725,N_7521,N_7434);
nor U7726 (N_7726,N_7586,N_7587);
nand U7727 (N_7727,N_7523,N_7459);
xnor U7728 (N_7728,N_7513,N_7562);
and U7729 (N_7729,N_7556,N_7465);
xor U7730 (N_7730,N_7543,N_7557);
xnor U7731 (N_7731,N_7562,N_7444);
xnor U7732 (N_7732,N_7485,N_7572);
and U7733 (N_7733,N_7490,N_7428);
nor U7734 (N_7734,N_7449,N_7573);
or U7735 (N_7735,N_7466,N_7543);
xor U7736 (N_7736,N_7466,N_7462);
and U7737 (N_7737,N_7441,N_7586);
xnor U7738 (N_7738,N_7431,N_7400);
nand U7739 (N_7739,N_7449,N_7455);
nor U7740 (N_7740,N_7408,N_7513);
or U7741 (N_7741,N_7504,N_7417);
and U7742 (N_7742,N_7582,N_7495);
xnor U7743 (N_7743,N_7412,N_7426);
nor U7744 (N_7744,N_7567,N_7553);
or U7745 (N_7745,N_7485,N_7591);
or U7746 (N_7746,N_7499,N_7539);
nand U7747 (N_7747,N_7472,N_7425);
nor U7748 (N_7748,N_7494,N_7490);
nor U7749 (N_7749,N_7547,N_7456);
nand U7750 (N_7750,N_7447,N_7437);
nand U7751 (N_7751,N_7563,N_7406);
and U7752 (N_7752,N_7440,N_7517);
nor U7753 (N_7753,N_7422,N_7556);
nand U7754 (N_7754,N_7412,N_7401);
nand U7755 (N_7755,N_7461,N_7517);
or U7756 (N_7756,N_7551,N_7485);
nand U7757 (N_7757,N_7477,N_7567);
nand U7758 (N_7758,N_7400,N_7565);
xnor U7759 (N_7759,N_7543,N_7521);
nor U7760 (N_7760,N_7583,N_7438);
and U7761 (N_7761,N_7534,N_7560);
and U7762 (N_7762,N_7521,N_7546);
nor U7763 (N_7763,N_7452,N_7588);
or U7764 (N_7764,N_7531,N_7515);
nand U7765 (N_7765,N_7478,N_7450);
or U7766 (N_7766,N_7558,N_7543);
or U7767 (N_7767,N_7421,N_7554);
nand U7768 (N_7768,N_7498,N_7523);
xnor U7769 (N_7769,N_7562,N_7561);
and U7770 (N_7770,N_7587,N_7428);
or U7771 (N_7771,N_7515,N_7574);
and U7772 (N_7772,N_7421,N_7485);
nand U7773 (N_7773,N_7505,N_7553);
or U7774 (N_7774,N_7528,N_7547);
nand U7775 (N_7775,N_7519,N_7425);
and U7776 (N_7776,N_7443,N_7476);
and U7777 (N_7777,N_7414,N_7508);
and U7778 (N_7778,N_7467,N_7429);
and U7779 (N_7779,N_7560,N_7417);
nor U7780 (N_7780,N_7564,N_7522);
or U7781 (N_7781,N_7434,N_7578);
and U7782 (N_7782,N_7459,N_7547);
xor U7783 (N_7783,N_7580,N_7560);
and U7784 (N_7784,N_7535,N_7575);
nor U7785 (N_7785,N_7482,N_7545);
nand U7786 (N_7786,N_7485,N_7481);
and U7787 (N_7787,N_7450,N_7540);
or U7788 (N_7788,N_7525,N_7545);
nand U7789 (N_7789,N_7565,N_7590);
and U7790 (N_7790,N_7576,N_7518);
or U7791 (N_7791,N_7553,N_7506);
nand U7792 (N_7792,N_7514,N_7508);
nand U7793 (N_7793,N_7583,N_7507);
nand U7794 (N_7794,N_7462,N_7478);
or U7795 (N_7795,N_7502,N_7447);
or U7796 (N_7796,N_7415,N_7459);
and U7797 (N_7797,N_7532,N_7498);
or U7798 (N_7798,N_7553,N_7478);
xor U7799 (N_7799,N_7517,N_7575);
or U7800 (N_7800,N_7643,N_7641);
or U7801 (N_7801,N_7763,N_7628);
nand U7802 (N_7802,N_7634,N_7609);
nor U7803 (N_7803,N_7780,N_7756);
and U7804 (N_7804,N_7759,N_7608);
and U7805 (N_7805,N_7657,N_7750);
nor U7806 (N_7806,N_7775,N_7732);
or U7807 (N_7807,N_7760,N_7639);
nand U7808 (N_7808,N_7681,N_7709);
nor U7809 (N_7809,N_7768,N_7623);
xnor U7810 (N_7810,N_7695,N_7617);
or U7811 (N_7811,N_7770,N_7795);
and U7812 (N_7812,N_7683,N_7751);
nand U7813 (N_7813,N_7700,N_7726);
nor U7814 (N_7814,N_7610,N_7682);
nor U7815 (N_7815,N_7616,N_7607);
nand U7816 (N_7816,N_7633,N_7799);
or U7817 (N_7817,N_7653,N_7785);
and U7818 (N_7818,N_7711,N_7757);
nand U7819 (N_7819,N_7745,N_7696);
nor U7820 (N_7820,N_7739,N_7753);
or U7821 (N_7821,N_7729,N_7779);
nand U7822 (N_7822,N_7767,N_7670);
nor U7823 (N_7823,N_7725,N_7788);
nand U7824 (N_7824,N_7638,N_7606);
nand U7825 (N_7825,N_7662,N_7783);
and U7826 (N_7826,N_7667,N_7733);
xor U7827 (N_7827,N_7621,N_7744);
nand U7828 (N_7828,N_7714,N_7717);
nand U7829 (N_7829,N_7650,N_7743);
nor U7830 (N_7830,N_7747,N_7784);
nor U7831 (N_7831,N_7630,N_7720);
nand U7832 (N_7832,N_7647,N_7635);
or U7833 (N_7833,N_7656,N_7602);
xor U7834 (N_7834,N_7731,N_7673);
and U7835 (N_7835,N_7614,N_7772);
xor U7836 (N_7836,N_7624,N_7605);
nor U7837 (N_7837,N_7613,N_7705);
nor U7838 (N_7838,N_7790,N_7737);
and U7839 (N_7839,N_7663,N_7664);
or U7840 (N_7840,N_7652,N_7707);
nor U7841 (N_7841,N_7690,N_7694);
or U7842 (N_7842,N_7715,N_7658);
or U7843 (N_7843,N_7674,N_7766);
nor U7844 (N_7844,N_7644,N_7651);
and U7845 (N_7845,N_7769,N_7771);
nor U7846 (N_7846,N_7713,N_7716);
or U7847 (N_7847,N_7789,N_7741);
nor U7848 (N_7848,N_7693,N_7679);
and U7849 (N_7849,N_7734,N_7797);
or U7850 (N_7850,N_7740,N_7773);
or U7851 (N_7851,N_7728,N_7710);
nor U7852 (N_7852,N_7661,N_7697);
nor U7853 (N_7853,N_7601,N_7631);
or U7854 (N_7854,N_7618,N_7724);
nor U7855 (N_7855,N_7615,N_7738);
nand U7856 (N_7856,N_7698,N_7604);
xnor U7857 (N_7857,N_7686,N_7781);
and U7858 (N_7858,N_7689,N_7794);
nor U7859 (N_7859,N_7676,N_7622);
nand U7860 (N_7860,N_7612,N_7701);
or U7861 (N_7861,N_7712,N_7688);
nand U7862 (N_7862,N_7774,N_7672);
or U7863 (N_7863,N_7629,N_7762);
nand U7864 (N_7864,N_7671,N_7678);
nand U7865 (N_7865,N_7619,N_7782);
nor U7866 (N_7866,N_7675,N_7666);
xor U7867 (N_7867,N_7748,N_7702);
nor U7868 (N_7868,N_7684,N_7765);
xnor U7869 (N_7869,N_7600,N_7777);
nand U7870 (N_7870,N_7755,N_7746);
nand U7871 (N_7871,N_7626,N_7754);
nand U7872 (N_7872,N_7721,N_7636);
nand U7873 (N_7873,N_7632,N_7718);
nor U7874 (N_7874,N_7719,N_7659);
and U7875 (N_7875,N_7708,N_7620);
nor U7876 (N_7876,N_7786,N_7723);
nand U7877 (N_7877,N_7742,N_7692);
nand U7878 (N_7878,N_7699,N_7798);
or U7879 (N_7879,N_7704,N_7691);
nor U7880 (N_7880,N_7749,N_7776);
nand U7881 (N_7881,N_7796,N_7646);
nand U7882 (N_7882,N_7752,N_7703);
xnor U7883 (N_7883,N_7791,N_7687);
or U7884 (N_7884,N_7787,N_7677);
xor U7885 (N_7885,N_7625,N_7627);
nand U7886 (N_7886,N_7680,N_7665);
nand U7887 (N_7887,N_7706,N_7735);
nand U7888 (N_7888,N_7764,N_7640);
and U7889 (N_7889,N_7778,N_7603);
nand U7890 (N_7890,N_7761,N_7649);
xor U7891 (N_7891,N_7637,N_7685);
or U7892 (N_7892,N_7642,N_7793);
nor U7893 (N_7893,N_7660,N_7730);
and U7894 (N_7894,N_7648,N_7736);
nor U7895 (N_7895,N_7722,N_7669);
and U7896 (N_7896,N_7655,N_7758);
nand U7897 (N_7897,N_7668,N_7727);
or U7898 (N_7898,N_7645,N_7654);
nor U7899 (N_7899,N_7611,N_7792);
or U7900 (N_7900,N_7752,N_7739);
nor U7901 (N_7901,N_7774,N_7653);
nor U7902 (N_7902,N_7641,N_7650);
or U7903 (N_7903,N_7747,N_7699);
nor U7904 (N_7904,N_7647,N_7615);
and U7905 (N_7905,N_7794,N_7772);
and U7906 (N_7906,N_7671,N_7665);
and U7907 (N_7907,N_7747,N_7743);
xnor U7908 (N_7908,N_7783,N_7683);
or U7909 (N_7909,N_7701,N_7725);
nor U7910 (N_7910,N_7670,N_7761);
and U7911 (N_7911,N_7661,N_7632);
nand U7912 (N_7912,N_7692,N_7638);
nor U7913 (N_7913,N_7699,N_7602);
or U7914 (N_7914,N_7662,N_7712);
nand U7915 (N_7915,N_7755,N_7603);
xor U7916 (N_7916,N_7789,N_7723);
xor U7917 (N_7917,N_7659,N_7673);
or U7918 (N_7918,N_7612,N_7756);
and U7919 (N_7919,N_7767,N_7601);
nor U7920 (N_7920,N_7658,N_7659);
xnor U7921 (N_7921,N_7651,N_7682);
and U7922 (N_7922,N_7746,N_7717);
or U7923 (N_7923,N_7671,N_7661);
xnor U7924 (N_7924,N_7739,N_7754);
and U7925 (N_7925,N_7689,N_7630);
and U7926 (N_7926,N_7769,N_7785);
or U7927 (N_7927,N_7683,N_7638);
or U7928 (N_7928,N_7645,N_7758);
or U7929 (N_7929,N_7680,N_7796);
xor U7930 (N_7930,N_7722,N_7719);
nand U7931 (N_7931,N_7695,N_7619);
nand U7932 (N_7932,N_7603,N_7674);
or U7933 (N_7933,N_7761,N_7722);
nand U7934 (N_7934,N_7763,N_7714);
and U7935 (N_7935,N_7743,N_7701);
and U7936 (N_7936,N_7771,N_7726);
nor U7937 (N_7937,N_7751,N_7709);
and U7938 (N_7938,N_7654,N_7717);
and U7939 (N_7939,N_7735,N_7654);
and U7940 (N_7940,N_7711,N_7724);
xnor U7941 (N_7941,N_7785,N_7767);
nand U7942 (N_7942,N_7628,N_7776);
nor U7943 (N_7943,N_7716,N_7676);
nand U7944 (N_7944,N_7776,N_7747);
nor U7945 (N_7945,N_7656,N_7641);
nor U7946 (N_7946,N_7621,N_7717);
and U7947 (N_7947,N_7682,N_7716);
nand U7948 (N_7948,N_7611,N_7630);
nand U7949 (N_7949,N_7751,N_7656);
and U7950 (N_7950,N_7663,N_7616);
nor U7951 (N_7951,N_7661,N_7685);
nor U7952 (N_7952,N_7621,N_7714);
or U7953 (N_7953,N_7703,N_7674);
nand U7954 (N_7954,N_7789,N_7772);
and U7955 (N_7955,N_7673,N_7635);
or U7956 (N_7956,N_7601,N_7787);
xnor U7957 (N_7957,N_7755,N_7748);
nor U7958 (N_7958,N_7764,N_7768);
and U7959 (N_7959,N_7668,N_7782);
and U7960 (N_7960,N_7738,N_7647);
xnor U7961 (N_7961,N_7723,N_7717);
nor U7962 (N_7962,N_7610,N_7768);
nor U7963 (N_7963,N_7645,N_7757);
nand U7964 (N_7964,N_7724,N_7735);
nor U7965 (N_7965,N_7648,N_7734);
nor U7966 (N_7966,N_7655,N_7731);
or U7967 (N_7967,N_7669,N_7730);
and U7968 (N_7968,N_7709,N_7682);
or U7969 (N_7969,N_7729,N_7675);
or U7970 (N_7970,N_7720,N_7758);
nand U7971 (N_7971,N_7655,N_7739);
or U7972 (N_7972,N_7788,N_7649);
and U7973 (N_7973,N_7728,N_7669);
xnor U7974 (N_7974,N_7681,N_7776);
nor U7975 (N_7975,N_7684,N_7628);
nand U7976 (N_7976,N_7663,N_7727);
and U7977 (N_7977,N_7738,N_7748);
and U7978 (N_7978,N_7756,N_7727);
nor U7979 (N_7979,N_7672,N_7613);
and U7980 (N_7980,N_7704,N_7619);
nor U7981 (N_7981,N_7748,N_7666);
and U7982 (N_7982,N_7769,N_7760);
nor U7983 (N_7983,N_7785,N_7646);
and U7984 (N_7984,N_7601,N_7692);
or U7985 (N_7985,N_7764,N_7680);
or U7986 (N_7986,N_7690,N_7732);
nand U7987 (N_7987,N_7738,N_7779);
or U7988 (N_7988,N_7681,N_7695);
or U7989 (N_7989,N_7620,N_7723);
and U7990 (N_7990,N_7770,N_7646);
nand U7991 (N_7991,N_7620,N_7724);
nor U7992 (N_7992,N_7725,N_7610);
xor U7993 (N_7993,N_7720,N_7738);
or U7994 (N_7994,N_7759,N_7735);
and U7995 (N_7995,N_7654,N_7614);
nor U7996 (N_7996,N_7710,N_7664);
xor U7997 (N_7997,N_7769,N_7693);
and U7998 (N_7998,N_7650,N_7638);
and U7999 (N_7999,N_7709,N_7640);
nand U8000 (N_8000,N_7900,N_7833);
nand U8001 (N_8001,N_7902,N_7838);
nor U8002 (N_8002,N_7867,N_7849);
nor U8003 (N_8003,N_7827,N_7869);
nor U8004 (N_8004,N_7977,N_7870);
or U8005 (N_8005,N_7897,N_7801);
nor U8006 (N_8006,N_7852,N_7837);
and U8007 (N_8007,N_7924,N_7800);
or U8008 (N_8008,N_7996,N_7915);
nor U8009 (N_8009,N_7885,N_7840);
and U8010 (N_8010,N_7925,N_7811);
and U8011 (N_8011,N_7803,N_7904);
nor U8012 (N_8012,N_7936,N_7958);
or U8013 (N_8013,N_7814,N_7985);
or U8014 (N_8014,N_7922,N_7993);
nor U8015 (N_8015,N_7937,N_7964);
or U8016 (N_8016,N_7911,N_7995);
or U8017 (N_8017,N_7947,N_7920);
nand U8018 (N_8018,N_7868,N_7820);
nor U8019 (N_8019,N_7826,N_7966);
or U8020 (N_8020,N_7836,N_7975);
nand U8021 (N_8021,N_7974,N_7898);
or U8022 (N_8022,N_7971,N_7851);
nand U8023 (N_8023,N_7857,N_7878);
nand U8024 (N_8024,N_7862,N_7972);
and U8025 (N_8025,N_7889,N_7956);
or U8026 (N_8026,N_7832,N_7808);
xnor U8027 (N_8027,N_7927,N_7951);
or U8028 (N_8028,N_7860,N_7874);
or U8029 (N_8029,N_7965,N_7893);
or U8030 (N_8030,N_7979,N_7976);
and U8031 (N_8031,N_7845,N_7962);
nand U8032 (N_8032,N_7831,N_7987);
or U8033 (N_8033,N_7994,N_7984);
nand U8034 (N_8034,N_7968,N_7846);
and U8035 (N_8035,N_7998,N_7855);
nor U8036 (N_8036,N_7821,N_7992);
nor U8037 (N_8037,N_7986,N_7918);
nand U8038 (N_8038,N_7969,N_7844);
xor U8039 (N_8039,N_7932,N_7933);
or U8040 (N_8040,N_7901,N_7948);
xnor U8041 (N_8041,N_7883,N_7828);
nand U8042 (N_8042,N_7890,N_7907);
and U8043 (N_8043,N_7818,N_7912);
nor U8044 (N_8044,N_7963,N_7863);
or U8045 (N_8045,N_7879,N_7812);
nand U8046 (N_8046,N_7978,N_7815);
and U8047 (N_8047,N_7980,N_7873);
and U8048 (N_8048,N_7991,N_7949);
nor U8049 (N_8049,N_7824,N_7944);
xnor U8050 (N_8050,N_7950,N_7959);
and U8051 (N_8051,N_7946,N_7960);
or U8052 (N_8052,N_7871,N_7967);
xnor U8053 (N_8053,N_7955,N_7886);
or U8054 (N_8054,N_7858,N_7806);
and U8055 (N_8055,N_7940,N_7953);
nand U8056 (N_8056,N_7938,N_7903);
and U8057 (N_8057,N_7850,N_7854);
nor U8058 (N_8058,N_7807,N_7997);
nor U8059 (N_8059,N_7926,N_7847);
nand U8060 (N_8060,N_7872,N_7892);
nor U8061 (N_8061,N_7919,N_7817);
nor U8062 (N_8062,N_7822,N_7896);
xor U8063 (N_8063,N_7954,N_7864);
xnor U8064 (N_8064,N_7819,N_7887);
or U8065 (N_8065,N_7983,N_7923);
nor U8066 (N_8066,N_7835,N_7816);
nand U8067 (N_8067,N_7899,N_7880);
nor U8068 (N_8068,N_7877,N_7804);
and U8069 (N_8069,N_7961,N_7908);
and U8070 (N_8070,N_7884,N_7842);
nand U8071 (N_8071,N_7982,N_7830);
nand U8072 (N_8072,N_7888,N_7823);
or U8073 (N_8073,N_7917,N_7859);
and U8074 (N_8074,N_7945,N_7999);
nand U8075 (N_8075,N_7894,N_7825);
nand U8076 (N_8076,N_7876,N_7906);
nand U8077 (N_8077,N_7990,N_7853);
nand U8078 (N_8078,N_7909,N_7802);
or U8079 (N_8079,N_7866,N_7813);
nor U8080 (N_8080,N_7856,N_7848);
nand U8081 (N_8081,N_7935,N_7952);
nand U8082 (N_8082,N_7910,N_7881);
xnor U8083 (N_8083,N_7973,N_7921);
xnor U8084 (N_8084,N_7916,N_7834);
nand U8085 (N_8085,N_7809,N_7829);
nand U8086 (N_8086,N_7841,N_7970);
or U8087 (N_8087,N_7989,N_7805);
and U8088 (N_8088,N_7934,N_7913);
and U8089 (N_8089,N_7865,N_7843);
nand U8090 (N_8090,N_7981,N_7810);
and U8091 (N_8091,N_7939,N_7988);
nor U8092 (N_8092,N_7882,N_7941);
or U8093 (N_8093,N_7930,N_7931);
nor U8094 (N_8094,N_7928,N_7914);
nor U8095 (N_8095,N_7839,N_7943);
nand U8096 (N_8096,N_7942,N_7957);
or U8097 (N_8097,N_7929,N_7875);
nand U8098 (N_8098,N_7861,N_7891);
or U8099 (N_8099,N_7895,N_7905);
nand U8100 (N_8100,N_7806,N_7869);
or U8101 (N_8101,N_7888,N_7805);
nand U8102 (N_8102,N_7862,N_7864);
nor U8103 (N_8103,N_7908,N_7906);
and U8104 (N_8104,N_7923,N_7966);
or U8105 (N_8105,N_7950,N_7817);
nand U8106 (N_8106,N_7936,N_7856);
nand U8107 (N_8107,N_7906,N_7828);
or U8108 (N_8108,N_7945,N_7935);
nand U8109 (N_8109,N_7898,N_7987);
and U8110 (N_8110,N_7804,N_7861);
xor U8111 (N_8111,N_7944,N_7981);
or U8112 (N_8112,N_7906,N_7800);
nand U8113 (N_8113,N_7950,N_7857);
nand U8114 (N_8114,N_7837,N_7873);
xor U8115 (N_8115,N_7857,N_7931);
or U8116 (N_8116,N_7893,N_7933);
or U8117 (N_8117,N_7810,N_7964);
nand U8118 (N_8118,N_7800,N_7976);
nand U8119 (N_8119,N_7870,N_7805);
nor U8120 (N_8120,N_7918,N_7960);
and U8121 (N_8121,N_7974,N_7903);
and U8122 (N_8122,N_7984,N_7839);
nand U8123 (N_8123,N_7994,N_7860);
or U8124 (N_8124,N_7932,N_7901);
nor U8125 (N_8125,N_7922,N_7900);
or U8126 (N_8126,N_7983,N_7907);
nand U8127 (N_8127,N_7987,N_7951);
nor U8128 (N_8128,N_7930,N_7947);
nand U8129 (N_8129,N_7980,N_7906);
nand U8130 (N_8130,N_7880,N_7904);
nor U8131 (N_8131,N_7971,N_7999);
and U8132 (N_8132,N_7988,N_7963);
nand U8133 (N_8133,N_7926,N_7928);
nand U8134 (N_8134,N_7829,N_7950);
nor U8135 (N_8135,N_7958,N_7992);
nand U8136 (N_8136,N_7926,N_7857);
and U8137 (N_8137,N_7930,N_7906);
and U8138 (N_8138,N_7803,N_7946);
or U8139 (N_8139,N_7997,N_7931);
or U8140 (N_8140,N_7883,N_7903);
and U8141 (N_8141,N_7816,N_7826);
nor U8142 (N_8142,N_7967,N_7850);
and U8143 (N_8143,N_7876,N_7817);
nor U8144 (N_8144,N_7879,N_7885);
nor U8145 (N_8145,N_7889,N_7832);
nor U8146 (N_8146,N_7903,N_7870);
nand U8147 (N_8147,N_7841,N_7969);
nor U8148 (N_8148,N_7997,N_7851);
or U8149 (N_8149,N_7982,N_7857);
nand U8150 (N_8150,N_7856,N_7905);
or U8151 (N_8151,N_7820,N_7858);
nor U8152 (N_8152,N_7804,N_7983);
or U8153 (N_8153,N_7832,N_7994);
and U8154 (N_8154,N_7829,N_7996);
nand U8155 (N_8155,N_7909,N_7956);
nor U8156 (N_8156,N_7835,N_7860);
nor U8157 (N_8157,N_7913,N_7852);
and U8158 (N_8158,N_7950,N_7984);
xnor U8159 (N_8159,N_7888,N_7845);
xor U8160 (N_8160,N_7879,N_7960);
nor U8161 (N_8161,N_7867,N_7984);
and U8162 (N_8162,N_7823,N_7884);
nand U8163 (N_8163,N_7946,N_7991);
xor U8164 (N_8164,N_7901,N_7946);
nor U8165 (N_8165,N_7960,N_7844);
nor U8166 (N_8166,N_7943,N_7908);
nor U8167 (N_8167,N_7876,N_7838);
nor U8168 (N_8168,N_7947,N_7978);
nor U8169 (N_8169,N_7817,N_7941);
nor U8170 (N_8170,N_7975,N_7921);
or U8171 (N_8171,N_7978,N_7980);
nand U8172 (N_8172,N_7950,N_7847);
or U8173 (N_8173,N_7906,N_7842);
or U8174 (N_8174,N_7911,N_7807);
xnor U8175 (N_8175,N_7908,N_7917);
nand U8176 (N_8176,N_7941,N_7950);
nand U8177 (N_8177,N_7998,N_7980);
or U8178 (N_8178,N_7869,N_7804);
nand U8179 (N_8179,N_7852,N_7962);
or U8180 (N_8180,N_7902,N_7960);
nor U8181 (N_8181,N_7853,N_7983);
nor U8182 (N_8182,N_7909,N_7815);
or U8183 (N_8183,N_7938,N_7850);
nand U8184 (N_8184,N_7815,N_7828);
nand U8185 (N_8185,N_7968,N_7855);
nand U8186 (N_8186,N_7989,N_7818);
or U8187 (N_8187,N_7871,N_7985);
nor U8188 (N_8188,N_7961,N_7800);
and U8189 (N_8189,N_7884,N_7948);
or U8190 (N_8190,N_7881,N_7825);
or U8191 (N_8191,N_7936,N_7815);
nor U8192 (N_8192,N_7959,N_7848);
or U8193 (N_8193,N_7857,N_7920);
or U8194 (N_8194,N_7886,N_7923);
nand U8195 (N_8195,N_7858,N_7879);
nor U8196 (N_8196,N_7943,N_7829);
and U8197 (N_8197,N_7920,N_7820);
nor U8198 (N_8198,N_7991,N_7886);
and U8199 (N_8199,N_7860,N_7886);
and U8200 (N_8200,N_8187,N_8104);
or U8201 (N_8201,N_8129,N_8126);
nor U8202 (N_8202,N_8184,N_8109);
nand U8203 (N_8203,N_8085,N_8152);
nor U8204 (N_8204,N_8175,N_8174);
and U8205 (N_8205,N_8067,N_8038);
or U8206 (N_8206,N_8043,N_8015);
nand U8207 (N_8207,N_8058,N_8191);
or U8208 (N_8208,N_8132,N_8177);
nor U8209 (N_8209,N_8195,N_8074);
nor U8210 (N_8210,N_8091,N_8116);
nor U8211 (N_8211,N_8061,N_8054);
nor U8212 (N_8212,N_8030,N_8083);
and U8213 (N_8213,N_8036,N_8135);
or U8214 (N_8214,N_8045,N_8055);
nor U8215 (N_8215,N_8044,N_8107);
or U8216 (N_8216,N_8170,N_8034);
and U8217 (N_8217,N_8014,N_8183);
nor U8218 (N_8218,N_8039,N_8007);
nor U8219 (N_8219,N_8008,N_8047);
nand U8220 (N_8220,N_8062,N_8118);
and U8221 (N_8221,N_8105,N_8141);
and U8222 (N_8222,N_8026,N_8179);
and U8223 (N_8223,N_8082,N_8143);
and U8224 (N_8224,N_8169,N_8134);
nor U8225 (N_8225,N_8000,N_8124);
xnor U8226 (N_8226,N_8128,N_8136);
nand U8227 (N_8227,N_8110,N_8076);
or U8228 (N_8228,N_8188,N_8147);
nand U8229 (N_8229,N_8005,N_8053);
or U8230 (N_8230,N_8086,N_8078);
and U8231 (N_8231,N_8160,N_8114);
or U8232 (N_8232,N_8139,N_8165);
nor U8233 (N_8233,N_8130,N_8112);
and U8234 (N_8234,N_8075,N_8190);
nand U8235 (N_8235,N_8042,N_8090);
nand U8236 (N_8236,N_8099,N_8144);
nor U8237 (N_8237,N_8020,N_8092);
nor U8238 (N_8238,N_8154,N_8193);
nor U8239 (N_8239,N_8133,N_8021);
or U8240 (N_8240,N_8117,N_8159);
xor U8241 (N_8241,N_8029,N_8089);
xnor U8242 (N_8242,N_8097,N_8010);
or U8243 (N_8243,N_8064,N_8155);
nor U8244 (N_8244,N_8120,N_8172);
and U8245 (N_8245,N_8140,N_8071);
or U8246 (N_8246,N_8138,N_8024);
nand U8247 (N_8247,N_8011,N_8153);
nor U8248 (N_8248,N_8066,N_8013);
or U8249 (N_8249,N_8173,N_8150);
or U8250 (N_8250,N_8131,N_8145);
nor U8251 (N_8251,N_8101,N_8103);
nand U8252 (N_8252,N_8027,N_8046);
and U8253 (N_8253,N_8088,N_8166);
and U8254 (N_8254,N_8148,N_8146);
nand U8255 (N_8255,N_8196,N_8186);
nand U8256 (N_8256,N_8069,N_8102);
nand U8257 (N_8257,N_8137,N_8068);
and U8258 (N_8258,N_8072,N_8163);
nand U8259 (N_8259,N_8040,N_8035);
and U8260 (N_8260,N_8079,N_8168);
and U8261 (N_8261,N_8002,N_8051);
and U8262 (N_8262,N_8050,N_8185);
nor U8263 (N_8263,N_8041,N_8158);
nor U8264 (N_8264,N_8176,N_8199);
xnor U8265 (N_8265,N_8115,N_8113);
xor U8266 (N_8266,N_8119,N_8161);
nand U8267 (N_8267,N_8031,N_8023);
nor U8268 (N_8268,N_8181,N_8077);
or U8269 (N_8269,N_8003,N_8001);
and U8270 (N_8270,N_8197,N_8096);
or U8271 (N_8271,N_8009,N_8025);
and U8272 (N_8272,N_8149,N_8022);
or U8273 (N_8273,N_8081,N_8070);
and U8274 (N_8274,N_8056,N_8095);
nand U8275 (N_8275,N_8033,N_8032);
xor U8276 (N_8276,N_8182,N_8059);
or U8277 (N_8277,N_8052,N_8048);
nand U8278 (N_8278,N_8004,N_8125);
and U8279 (N_8279,N_8189,N_8164);
or U8280 (N_8280,N_8121,N_8156);
nor U8281 (N_8281,N_8122,N_8012);
nand U8282 (N_8282,N_8060,N_8087);
or U8283 (N_8283,N_8106,N_8093);
nand U8284 (N_8284,N_8162,N_8180);
and U8285 (N_8285,N_8192,N_8111);
and U8286 (N_8286,N_8151,N_8157);
nor U8287 (N_8287,N_8028,N_8019);
and U8288 (N_8288,N_8065,N_8080);
and U8289 (N_8289,N_8108,N_8017);
nand U8290 (N_8290,N_8084,N_8171);
nor U8291 (N_8291,N_8049,N_8057);
and U8292 (N_8292,N_8100,N_8006);
or U8293 (N_8293,N_8178,N_8037);
nand U8294 (N_8294,N_8167,N_8098);
and U8295 (N_8295,N_8194,N_8198);
or U8296 (N_8296,N_8073,N_8127);
xor U8297 (N_8297,N_8018,N_8094);
nor U8298 (N_8298,N_8123,N_8016);
nor U8299 (N_8299,N_8063,N_8142);
nand U8300 (N_8300,N_8043,N_8129);
nand U8301 (N_8301,N_8140,N_8118);
and U8302 (N_8302,N_8001,N_8020);
or U8303 (N_8303,N_8099,N_8048);
nand U8304 (N_8304,N_8068,N_8060);
and U8305 (N_8305,N_8198,N_8167);
and U8306 (N_8306,N_8096,N_8110);
nand U8307 (N_8307,N_8184,N_8003);
nor U8308 (N_8308,N_8148,N_8197);
or U8309 (N_8309,N_8039,N_8138);
nor U8310 (N_8310,N_8030,N_8190);
xor U8311 (N_8311,N_8075,N_8076);
or U8312 (N_8312,N_8175,N_8162);
and U8313 (N_8313,N_8070,N_8158);
xnor U8314 (N_8314,N_8049,N_8136);
or U8315 (N_8315,N_8052,N_8056);
xor U8316 (N_8316,N_8181,N_8094);
xnor U8317 (N_8317,N_8131,N_8123);
and U8318 (N_8318,N_8042,N_8076);
nand U8319 (N_8319,N_8187,N_8194);
nor U8320 (N_8320,N_8024,N_8132);
and U8321 (N_8321,N_8012,N_8026);
nor U8322 (N_8322,N_8113,N_8182);
xor U8323 (N_8323,N_8075,N_8126);
nor U8324 (N_8324,N_8075,N_8187);
nor U8325 (N_8325,N_8130,N_8100);
or U8326 (N_8326,N_8107,N_8132);
nor U8327 (N_8327,N_8113,N_8045);
or U8328 (N_8328,N_8008,N_8155);
and U8329 (N_8329,N_8127,N_8116);
or U8330 (N_8330,N_8023,N_8020);
or U8331 (N_8331,N_8163,N_8086);
and U8332 (N_8332,N_8105,N_8051);
or U8333 (N_8333,N_8011,N_8185);
nand U8334 (N_8334,N_8188,N_8044);
nor U8335 (N_8335,N_8146,N_8112);
and U8336 (N_8336,N_8029,N_8126);
or U8337 (N_8337,N_8192,N_8070);
nor U8338 (N_8338,N_8192,N_8154);
nand U8339 (N_8339,N_8033,N_8072);
or U8340 (N_8340,N_8180,N_8126);
nand U8341 (N_8341,N_8008,N_8132);
xor U8342 (N_8342,N_8163,N_8159);
and U8343 (N_8343,N_8175,N_8097);
nor U8344 (N_8344,N_8092,N_8191);
nand U8345 (N_8345,N_8154,N_8068);
and U8346 (N_8346,N_8134,N_8085);
xnor U8347 (N_8347,N_8140,N_8197);
nor U8348 (N_8348,N_8193,N_8096);
and U8349 (N_8349,N_8158,N_8047);
and U8350 (N_8350,N_8160,N_8093);
and U8351 (N_8351,N_8069,N_8128);
xor U8352 (N_8352,N_8089,N_8170);
nand U8353 (N_8353,N_8161,N_8060);
and U8354 (N_8354,N_8184,N_8168);
nor U8355 (N_8355,N_8038,N_8174);
xnor U8356 (N_8356,N_8114,N_8029);
or U8357 (N_8357,N_8093,N_8048);
xnor U8358 (N_8358,N_8079,N_8127);
or U8359 (N_8359,N_8086,N_8167);
and U8360 (N_8360,N_8030,N_8127);
or U8361 (N_8361,N_8094,N_8040);
or U8362 (N_8362,N_8186,N_8031);
or U8363 (N_8363,N_8085,N_8057);
nor U8364 (N_8364,N_8188,N_8005);
nand U8365 (N_8365,N_8026,N_8099);
and U8366 (N_8366,N_8193,N_8007);
nor U8367 (N_8367,N_8115,N_8120);
xor U8368 (N_8368,N_8180,N_8025);
nor U8369 (N_8369,N_8175,N_8196);
and U8370 (N_8370,N_8198,N_8127);
or U8371 (N_8371,N_8011,N_8065);
and U8372 (N_8372,N_8038,N_8006);
xor U8373 (N_8373,N_8146,N_8000);
or U8374 (N_8374,N_8045,N_8175);
xor U8375 (N_8375,N_8011,N_8095);
or U8376 (N_8376,N_8109,N_8150);
nand U8377 (N_8377,N_8098,N_8152);
nand U8378 (N_8378,N_8064,N_8060);
nor U8379 (N_8379,N_8130,N_8069);
nor U8380 (N_8380,N_8106,N_8123);
or U8381 (N_8381,N_8065,N_8035);
nor U8382 (N_8382,N_8021,N_8167);
xnor U8383 (N_8383,N_8082,N_8076);
nand U8384 (N_8384,N_8023,N_8080);
and U8385 (N_8385,N_8086,N_8041);
or U8386 (N_8386,N_8066,N_8144);
and U8387 (N_8387,N_8048,N_8100);
and U8388 (N_8388,N_8046,N_8023);
nand U8389 (N_8389,N_8084,N_8111);
and U8390 (N_8390,N_8130,N_8050);
nand U8391 (N_8391,N_8132,N_8180);
and U8392 (N_8392,N_8168,N_8191);
or U8393 (N_8393,N_8026,N_8091);
and U8394 (N_8394,N_8053,N_8059);
nand U8395 (N_8395,N_8070,N_8124);
or U8396 (N_8396,N_8066,N_8065);
nor U8397 (N_8397,N_8072,N_8066);
nor U8398 (N_8398,N_8154,N_8108);
nor U8399 (N_8399,N_8198,N_8055);
nand U8400 (N_8400,N_8381,N_8248);
nand U8401 (N_8401,N_8373,N_8286);
or U8402 (N_8402,N_8244,N_8347);
nand U8403 (N_8403,N_8226,N_8210);
and U8404 (N_8404,N_8321,N_8219);
and U8405 (N_8405,N_8380,N_8229);
xor U8406 (N_8406,N_8383,N_8280);
or U8407 (N_8407,N_8310,N_8395);
or U8408 (N_8408,N_8379,N_8333);
and U8409 (N_8409,N_8334,N_8369);
nand U8410 (N_8410,N_8370,N_8367);
nand U8411 (N_8411,N_8218,N_8304);
and U8412 (N_8412,N_8261,N_8258);
nor U8413 (N_8413,N_8339,N_8275);
nor U8414 (N_8414,N_8313,N_8257);
or U8415 (N_8415,N_8223,N_8217);
and U8416 (N_8416,N_8213,N_8341);
or U8417 (N_8417,N_8228,N_8282);
nand U8418 (N_8418,N_8396,N_8366);
xor U8419 (N_8419,N_8355,N_8338);
or U8420 (N_8420,N_8300,N_8352);
or U8421 (N_8421,N_8279,N_8284);
nand U8422 (N_8422,N_8269,N_8377);
or U8423 (N_8423,N_8225,N_8245);
or U8424 (N_8424,N_8259,N_8351);
and U8425 (N_8425,N_8212,N_8320);
and U8426 (N_8426,N_8289,N_8220);
or U8427 (N_8427,N_8357,N_8332);
xor U8428 (N_8428,N_8281,N_8241);
xnor U8429 (N_8429,N_8208,N_8363);
or U8430 (N_8430,N_8246,N_8233);
or U8431 (N_8431,N_8323,N_8202);
nor U8432 (N_8432,N_8267,N_8205);
or U8433 (N_8433,N_8335,N_8372);
xnor U8434 (N_8434,N_8353,N_8316);
nor U8435 (N_8435,N_8359,N_8388);
or U8436 (N_8436,N_8287,N_8399);
or U8437 (N_8437,N_8387,N_8361);
nand U8438 (N_8438,N_8243,N_8266);
nor U8439 (N_8439,N_8262,N_8356);
nor U8440 (N_8440,N_8371,N_8293);
nand U8441 (N_8441,N_8238,N_8348);
or U8442 (N_8442,N_8260,N_8382);
nand U8443 (N_8443,N_8346,N_8354);
or U8444 (N_8444,N_8274,N_8368);
or U8445 (N_8445,N_8285,N_8214);
and U8446 (N_8446,N_8206,N_8365);
or U8447 (N_8447,N_8394,N_8340);
nor U8448 (N_8448,N_8236,N_8215);
nand U8449 (N_8449,N_8314,N_8331);
or U8450 (N_8450,N_8299,N_8325);
and U8451 (N_8451,N_8291,N_8242);
nor U8452 (N_8452,N_8294,N_8398);
nor U8453 (N_8453,N_8328,N_8270);
and U8454 (N_8454,N_8318,N_8337);
nor U8455 (N_8455,N_8374,N_8230);
and U8456 (N_8456,N_8385,N_8319);
nor U8457 (N_8457,N_8364,N_8397);
nor U8458 (N_8458,N_8303,N_8342);
or U8459 (N_8459,N_8297,N_8204);
and U8460 (N_8460,N_8386,N_8256);
nor U8461 (N_8461,N_8330,N_8298);
nor U8462 (N_8462,N_8278,N_8311);
or U8463 (N_8463,N_8222,N_8211);
or U8464 (N_8464,N_8322,N_8307);
xor U8465 (N_8465,N_8315,N_8272);
nand U8466 (N_8466,N_8263,N_8251);
nand U8467 (N_8467,N_8358,N_8306);
nor U8468 (N_8468,N_8255,N_8253);
xnor U8469 (N_8469,N_8290,N_8209);
and U8470 (N_8470,N_8265,N_8232);
or U8471 (N_8471,N_8239,N_8305);
nand U8472 (N_8472,N_8201,N_8390);
nor U8473 (N_8473,N_8324,N_8329);
or U8474 (N_8474,N_8231,N_8203);
and U8475 (N_8475,N_8277,N_8234);
or U8476 (N_8476,N_8237,N_8224);
nor U8477 (N_8477,N_8344,N_8292);
nor U8478 (N_8478,N_8249,N_8283);
nand U8479 (N_8479,N_8221,N_8227);
nor U8480 (N_8480,N_8216,N_8378);
xor U8481 (N_8481,N_8250,N_8302);
nand U8482 (N_8482,N_8247,N_8200);
and U8483 (N_8483,N_8391,N_8271);
xor U8484 (N_8484,N_8360,N_8375);
nand U8485 (N_8485,N_8389,N_8309);
nand U8486 (N_8486,N_8264,N_8240);
and U8487 (N_8487,N_8268,N_8295);
or U8488 (N_8488,N_8207,N_8376);
nand U8489 (N_8489,N_8362,N_8350);
and U8490 (N_8490,N_8308,N_8345);
or U8491 (N_8491,N_8317,N_8301);
and U8492 (N_8492,N_8288,N_8326);
and U8493 (N_8493,N_8349,N_8312);
or U8494 (N_8494,N_8327,N_8343);
or U8495 (N_8495,N_8392,N_8273);
nor U8496 (N_8496,N_8393,N_8384);
or U8497 (N_8497,N_8336,N_8254);
and U8498 (N_8498,N_8276,N_8235);
or U8499 (N_8499,N_8252,N_8296);
or U8500 (N_8500,N_8343,N_8286);
and U8501 (N_8501,N_8369,N_8263);
xnor U8502 (N_8502,N_8384,N_8395);
nor U8503 (N_8503,N_8262,N_8306);
nor U8504 (N_8504,N_8245,N_8390);
and U8505 (N_8505,N_8325,N_8318);
xor U8506 (N_8506,N_8350,N_8370);
nand U8507 (N_8507,N_8335,N_8297);
and U8508 (N_8508,N_8282,N_8240);
nor U8509 (N_8509,N_8226,N_8205);
and U8510 (N_8510,N_8246,N_8362);
and U8511 (N_8511,N_8209,N_8257);
xor U8512 (N_8512,N_8210,N_8235);
and U8513 (N_8513,N_8315,N_8264);
or U8514 (N_8514,N_8309,N_8333);
or U8515 (N_8515,N_8344,N_8264);
nor U8516 (N_8516,N_8292,N_8265);
nand U8517 (N_8517,N_8296,N_8284);
nand U8518 (N_8518,N_8349,N_8306);
xor U8519 (N_8519,N_8381,N_8259);
and U8520 (N_8520,N_8390,N_8346);
xnor U8521 (N_8521,N_8341,N_8389);
nand U8522 (N_8522,N_8398,N_8303);
or U8523 (N_8523,N_8268,N_8253);
nor U8524 (N_8524,N_8293,N_8207);
or U8525 (N_8525,N_8217,N_8371);
nand U8526 (N_8526,N_8399,N_8337);
nor U8527 (N_8527,N_8331,N_8253);
nand U8528 (N_8528,N_8356,N_8238);
nand U8529 (N_8529,N_8354,N_8389);
or U8530 (N_8530,N_8240,N_8211);
nand U8531 (N_8531,N_8377,N_8319);
nand U8532 (N_8532,N_8289,N_8368);
nor U8533 (N_8533,N_8318,N_8290);
or U8534 (N_8534,N_8344,N_8224);
or U8535 (N_8535,N_8292,N_8368);
nor U8536 (N_8536,N_8325,N_8397);
xnor U8537 (N_8537,N_8329,N_8264);
or U8538 (N_8538,N_8309,N_8384);
or U8539 (N_8539,N_8376,N_8250);
nor U8540 (N_8540,N_8295,N_8255);
and U8541 (N_8541,N_8295,N_8298);
and U8542 (N_8542,N_8253,N_8295);
and U8543 (N_8543,N_8349,N_8333);
and U8544 (N_8544,N_8200,N_8236);
xnor U8545 (N_8545,N_8296,N_8351);
or U8546 (N_8546,N_8308,N_8332);
nand U8547 (N_8547,N_8350,N_8334);
or U8548 (N_8548,N_8336,N_8218);
or U8549 (N_8549,N_8244,N_8200);
nor U8550 (N_8550,N_8373,N_8289);
nand U8551 (N_8551,N_8223,N_8359);
xor U8552 (N_8552,N_8271,N_8265);
nand U8553 (N_8553,N_8316,N_8282);
or U8554 (N_8554,N_8389,N_8328);
or U8555 (N_8555,N_8342,N_8253);
xnor U8556 (N_8556,N_8326,N_8385);
nor U8557 (N_8557,N_8319,N_8282);
xnor U8558 (N_8558,N_8264,N_8396);
nor U8559 (N_8559,N_8329,N_8318);
xnor U8560 (N_8560,N_8243,N_8329);
or U8561 (N_8561,N_8387,N_8243);
nor U8562 (N_8562,N_8231,N_8228);
nand U8563 (N_8563,N_8320,N_8295);
nor U8564 (N_8564,N_8272,N_8386);
nor U8565 (N_8565,N_8345,N_8233);
nor U8566 (N_8566,N_8394,N_8206);
nand U8567 (N_8567,N_8294,N_8306);
xnor U8568 (N_8568,N_8207,N_8362);
nand U8569 (N_8569,N_8283,N_8208);
nor U8570 (N_8570,N_8243,N_8364);
nand U8571 (N_8571,N_8234,N_8307);
nor U8572 (N_8572,N_8219,N_8338);
or U8573 (N_8573,N_8294,N_8230);
or U8574 (N_8574,N_8279,N_8330);
nor U8575 (N_8575,N_8394,N_8389);
nand U8576 (N_8576,N_8359,N_8302);
nand U8577 (N_8577,N_8304,N_8307);
or U8578 (N_8578,N_8235,N_8297);
nor U8579 (N_8579,N_8234,N_8272);
or U8580 (N_8580,N_8322,N_8230);
and U8581 (N_8581,N_8224,N_8232);
nor U8582 (N_8582,N_8290,N_8355);
and U8583 (N_8583,N_8349,N_8364);
or U8584 (N_8584,N_8373,N_8360);
xnor U8585 (N_8585,N_8375,N_8288);
or U8586 (N_8586,N_8291,N_8323);
and U8587 (N_8587,N_8357,N_8293);
and U8588 (N_8588,N_8387,N_8244);
nand U8589 (N_8589,N_8368,N_8313);
nand U8590 (N_8590,N_8296,N_8260);
xnor U8591 (N_8591,N_8374,N_8291);
or U8592 (N_8592,N_8285,N_8368);
nor U8593 (N_8593,N_8347,N_8270);
and U8594 (N_8594,N_8392,N_8209);
nand U8595 (N_8595,N_8305,N_8333);
or U8596 (N_8596,N_8378,N_8270);
or U8597 (N_8597,N_8388,N_8368);
nand U8598 (N_8598,N_8398,N_8237);
and U8599 (N_8599,N_8395,N_8342);
or U8600 (N_8600,N_8558,N_8403);
xor U8601 (N_8601,N_8549,N_8500);
nand U8602 (N_8602,N_8589,N_8406);
and U8603 (N_8603,N_8465,N_8409);
nand U8604 (N_8604,N_8433,N_8529);
nand U8605 (N_8605,N_8469,N_8437);
or U8606 (N_8606,N_8509,N_8568);
or U8607 (N_8607,N_8517,N_8514);
and U8608 (N_8608,N_8490,N_8575);
nor U8609 (N_8609,N_8519,N_8561);
nor U8610 (N_8610,N_8489,N_8539);
or U8611 (N_8611,N_8476,N_8594);
nand U8612 (N_8612,N_8516,N_8559);
or U8613 (N_8613,N_8477,N_8591);
nand U8614 (N_8614,N_8446,N_8571);
nor U8615 (N_8615,N_8416,N_8435);
and U8616 (N_8616,N_8598,N_8551);
and U8617 (N_8617,N_8494,N_8468);
nor U8618 (N_8618,N_8544,N_8426);
and U8619 (N_8619,N_8515,N_8581);
nor U8620 (N_8620,N_8506,N_8419);
or U8621 (N_8621,N_8505,N_8497);
nand U8622 (N_8622,N_8560,N_8548);
or U8623 (N_8623,N_8556,N_8481);
nand U8624 (N_8624,N_8498,N_8460);
nor U8625 (N_8625,N_8570,N_8553);
nand U8626 (N_8626,N_8520,N_8586);
xnor U8627 (N_8627,N_8532,N_8486);
nand U8628 (N_8628,N_8522,N_8564);
or U8629 (N_8629,N_8455,N_8474);
nor U8630 (N_8630,N_8488,N_8493);
nor U8631 (N_8631,N_8495,N_8577);
xor U8632 (N_8632,N_8457,N_8540);
nand U8633 (N_8633,N_8580,N_8450);
or U8634 (N_8634,N_8464,N_8443);
nor U8635 (N_8635,N_8459,N_8547);
nor U8636 (N_8636,N_8579,N_8537);
and U8637 (N_8637,N_8438,N_8587);
nand U8638 (N_8638,N_8496,N_8550);
nor U8639 (N_8639,N_8415,N_8422);
and U8640 (N_8640,N_8541,N_8472);
or U8641 (N_8641,N_8456,N_8499);
and U8642 (N_8642,N_8471,N_8595);
or U8643 (N_8643,N_8504,N_8585);
or U8644 (N_8644,N_8428,N_8404);
xor U8645 (N_8645,N_8593,N_8400);
or U8646 (N_8646,N_8508,N_8573);
xnor U8647 (N_8647,N_8533,N_8451);
nor U8648 (N_8648,N_8507,N_8427);
or U8649 (N_8649,N_8442,N_8590);
xor U8650 (N_8650,N_8431,N_8430);
nor U8651 (N_8651,N_8420,N_8411);
nand U8652 (N_8652,N_8424,N_8536);
or U8653 (N_8653,N_8578,N_8449);
and U8654 (N_8654,N_8535,N_8583);
or U8655 (N_8655,N_8531,N_8557);
nor U8656 (N_8656,N_8487,N_8475);
and U8657 (N_8657,N_8574,N_8596);
xnor U8658 (N_8658,N_8597,N_8480);
or U8659 (N_8659,N_8562,N_8521);
and U8660 (N_8660,N_8552,N_8513);
nor U8661 (N_8661,N_8413,N_8524);
nor U8662 (N_8662,N_8418,N_8408);
nand U8663 (N_8663,N_8492,N_8491);
or U8664 (N_8664,N_8458,N_8410);
and U8665 (N_8665,N_8510,N_8432);
xnor U8666 (N_8666,N_8402,N_8523);
nand U8667 (N_8667,N_8441,N_8576);
or U8668 (N_8668,N_8545,N_8423);
nor U8669 (N_8669,N_8599,N_8445);
xnor U8670 (N_8670,N_8567,N_8582);
nor U8671 (N_8671,N_8592,N_8542);
nand U8672 (N_8672,N_8440,N_8452);
and U8673 (N_8673,N_8518,N_8565);
and U8674 (N_8674,N_8526,N_8543);
nand U8675 (N_8675,N_8530,N_8525);
or U8676 (N_8676,N_8478,N_8546);
and U8677 (N_8677,N_8461,N_8528);
nand U8678 (N_8678,N_8483,N_8566);
or U8679 (N_8679,N_8425,N_8588);
xnor U8680 (N_8680,N_8563,N_8470);
nand U8681 (N_8681,N_8473,N_8463);
and U8682 (N_8682,N_8534,N_8569);
or U8683 (N_8683,N_8405,N_8447);
nor U8684 (N_8684,N_8444,N_8453);
xor U8685 (N_8685,N_8434,N_8555);
nor U8686 (N_8686,N_8538,N_8572);
or U8687 (N_8687,N_8436,N_8448);
nand U8688 (N_8688,N_8439,N_8502);
and U8689 (N_8689,N_8407,N_8401);
and U8690 (N_8690,N_8417,N_8462);
or U8691 (N_8691,N_8467,N_8554);
nand U8692 (N_8692,N_8511,N_8484);
and U8693 (N_8693,N_8503,N_8412);
nor U8694 (N_8694,N_8429,N_8466);
and U8695 (N_8695,N_8421,N_8512);
nor U8696 (N_8696,N_8501,N_8482);
xnor U8697 (N_8697,N_8485,N_8527);
nand U8698 (N_8698,N_8414,N_8479);
nand U8699 (N_8699,N_8584,N_8454);
nor U8700 (N_8700,N_8496,N_8457);
and U8701 (N_8701,N_8580,N_8525);
or U8702 (N_8702,N_8455,N_8491);
or U8703 (N_8703,N_8564,N_8416);
xor U8704 (N_8704,N_8593,N_8598);
nand U8705 (N_8705,N_8491,N_8501);
nor U8706 (N_8706,N_8433,N_8480);
or U8707 (N_8707,N_8472,N_8473);
and U8708 (N_8708,N_8543,N_8434);
nor U8709 (N_8709,N_8446,N_8529);
or U8710 (N_8710,N_8484,N_8409);
xnor U8711 (N_8711,N_8409,N_8433);
or U8712 (N_8712,N_8471,N_8550);
nor U8713 (N_8713,N_8522,N_8512);
nand U8714 (N_8714,N_8470,N_8522);
nand U8715 (N_8715,N_8470,N_8585);
and U8716 (N_8716,N_8520,N_8400);
nand U8717 (N_8717,N_8565,N_8575);
and U8718 (N_8718,N_8593,N_8421);
and U8719 (N_8719,N_8464,N_8575);
nand U8720 (N_8720,N_8591,N_8465);
nand U8721 (N_8721,N_8526,N_8458);
xnor U8722 (N_8722,N_8491,N_8493);
and U8723 (N_8723,N_8468,N_8436);
and U8724 (N_8724,N_8476,N_8409);
nor U8725 (N_8725,N_8530,N_8404);
and U8726 (N_8726,N_8549,N_8580);
or U8727 (N_8727,N_8479,N_8488);
nor U8728 (N_8728,N_8467,N_8528);
xnor U8729 (N_8729,N_8567,N_8495);
and U8730 (N_8730,N_8510,N_8549);
nand U8731 (N_8731,N_8572,N_8569);
and U8732 (N_8732,N_8457,N_8475);
or U8733 (N_8733,N_8463,N_8431);
xor U8734 (N_8734,N_8528,N_8415);
nor U8735 (N_8735,N_8558,N_8538);
nand U8736 (N_8736,N_8426,N_8510);
nor U8737 (N_8737,N_8424,N_8573);
and U8738 (N_8738,N_8599,N_8409);
and U8739 (N_8739,N_8509,N_8516);
nor U8740 (N_8740,N_8553,N_8547);
and U8741 (N_8741,N_8550,N_8515);
nor U8742 (N_8742,N_8414,N_8410);
xnor U8743 (N_8743,N_8561,N_8459);
nor U8744 (N_8744,N_8505,N_8476);
or U8745 (N_8745,N_8435,N_8427);
nand U8746 (N_8746,N_8582,N_8407);
and U8747 (N_8747,N_8428,N_8537);
nand U8748 (N_8748,N_8525,N_8546);
and U8749 (N_8749,N_8497,N_8582);
nor U8750 (N_8750,N_8590,N_8582);
and U8751 (N_8751,N_8579,N_8500);
or U8752 (N_8752,N_8442,N_8463);
or U8753 (N_8753,N_8465,N_8538);
nand U8754 (N_8754,N_8581,N_8437);
nor U8755 (N_8755,N_8532,N_8564);
and U8756 (N_8756,N_8554,N_8489);
and U8757 (N_8757,N_8573,N_8556);
or U8758 (N_8758,N_8422,N_8492);
nor U8759 (N_8759,N_8403,N_8598);
or U8760 (N_8760,N_8444,N_8525);
and U8761 (N_8761,N_8569,N_8551);
or U8762 (N_8762,N_8447,N_8448);
nand U8763 (N_8763,N_8460,N_8437);
nand U8764 (N_8764,N_8440,N_8505);
or U8765 (N_8765,N_8472,N_8417);
and U8766 (N_8766,N_8439,N_8453);
nor U8767 (N_8767,N_8569,N_8420);
and U8768 (N_8768,N_8528,N_8565);
and U8769 (N_8769,N_8550,N_8523);
or U8770 (N_8770,N_8580,N_8425);
and U8771 (N_8771,N_8475,N_8596);
and U8772 (N_8772,N_8481,N_8450);
nor U8773 (N_8773,N_8549,N_8456);
nor U8774 (N_8774,N_8505,N_8557);
or U8775 (N_8775,N_8477,N_8539);
nor U8776 (N_8776,N_8434,N_8502);
nand U8777 (N_8777,N_8577,N_8424);
or U8778 (N_8778,N_8522,N_8517);
nor U8779 (N_8779,N_8592,N_8533);
or U8780 (N_8780,N_8501,N_8471);
nand U8781 (N_8781,N_8427,N_8526);
and U8782 (N_8782,N_8503,N_8479);
xnor U8783 (N_8783,N_8488,N_8515);
and U8784 (N_8784,N_8543,N_8429);
nor U8785 (N_8785,N_8474,N_8401);
or U8786 (N_8786,N_8454,N_8559);
nor U8787 (N_8787,N_8596,N_8447);
and U8788 (N_8788,N_8495,N_8440);
or U8789 (N_8789,N_8420,N_8578);
nor U8790 (N_8790,N_8527,N_8551);
and U8791 (N_8791,N_8517,N_8507);
or U8792 (N_8792,N_8434,N_8512);
or U8793 (N_8793,N_8534,N_8478);
or U8794 (N_8794,N_8523,N_8476);
nor U8795 (N_8795,N_8508,N_8475);
or U8796 (N_8796,N_8569,N_8452);
or U8797 (N_8797,N_8584,N_8417);
nor U8798 (N_8798,N_8428,N_8527);
and U8799 (N_8799,N_8423,N_8589);
nand U8800 (N_8800,N_8669,N_8716);
or U8801 (N_8801,N_8625,N_8696);
or U8802 (N_8802,N_8712,N_8624);
nand U8803 (N_8803,N_8730,N_8648);
xnor U8804 (N_8804,N_8715,N_8787);
and U8805 (N_8805,N_8740,N_8731);
nor U8806 (N_8806,N_8620,N_8656);
or U8807 (N_8807,N_8738,N_8788);
and U8808 (N_8808,N_8641,N_8630);
and U8809 (N_8809,N_8707,N_8644);
nor U8810 (N_8810,N_8632,N_8617);
or U8811 (N_8811,N_8703,N_8640);
and U8812 (N_8812,N_8764,N_8623);
nand U8813 (N_8813,N_8627,N_8643);
nor U8814 (N_8814,N_8766,N_8743);
xnor U8815 (N_8815,N_8756,N_8762);
nor U8816 (N_8816,N_8718,N_8774);
nor U8817 (N_8817,N_8609,N_8659);
or U8818 (N_8818,N_8747,N_8708);
or U8819 (N_8819,N_8688,N_8631);
and U8820 (N_8820,N_8654,N_8770);
nor U8821 (N_8821,N_8767,N_8606);
and U8822 (N_8822,N_8755,N_8645);
xnor U8823 (N_8823,N_8786,N_8634);
nor U8824 (N_8824,N_8795,N_8773);
or U8825 (N_8825,N_8678,N_8721);
and U8826 (N_8826,N_8646,N_8761);
nor U8827 (N_8827,N_8799,N_8649);
or U8828 (N_8828,N_8750,N_8769);
xor U8829 (N_8829,N_8790,N_8724);
nor U8830 (N_8830,N_8791,N_8725);
or U8831 (N_8831,N_8663,N_8779);
or U8832 (N_8832,N_8727,N_8768);
and U8833 (N_8833,N_8616,N_8601);
xor U8834 (N_8834,N_8600,N_8670);
xnor U8835 (N_8835,N_8772,N_8677);
nor U8836 (N_8836,N_8763,N_8642);
xor U8837 (N_8837,N_8783,N_8662);
nor U8838 (N_8838,N_8776,N_8660);
nor U8839 (N_8839,N_8621,N_8690);
nor U8840 (N_8840,N_8733,N_8650);
nor U8841 (N_8841,N_8757,N_8753);
or U8842 (N_8842,N_8680,N_8658);
xnor U8843 (N_8843,N_8666,N_8639);
nand U8844 (N_8844,N_8636,N_8711);
or U8845 (N_8845,N_8647,N_8653);
and U8846 (N_8846,N_8612,N_8661);
nand U8847 (N_8847,N_8635,N_8760);
and U8848 (N_8848,N_8734,N_8693);
nand U8849 (N_8849,N_8792,N_8668);
or U8850 (N_8850,N_8604,N_8726);
or U8851 (N_8851,N_8687,N_8744);
nand U8852 (N_8852,N_8782,N_8793);
or U8853 (N_8853,N_8602,N_8697);
or U8854 (N_8854,N_8603,N_8619);
nor U8855 (N_8855,N_8723,N_8710);
or U8856 (N_8856,N_8665,N_8780);
nor U8857 (N_8857,N_8682,N_8695);
nand U8858 (N_8858,N_8615,N_8797);
xnor U8859 (N_8859,N_8657,N_8671);
nand U8860 (N_8860,N_8796,N_8720);
or U8861 (N_8861,N_8737,N_8789);
and U8862 (N_8862,N_8667,N_8626);
and U8863 (N_8863,N_8675,N_8709);
or U8864 (N_8864,N_8638,N_8702);
nand U8865 (N_8865,N_8637,N_8729);
and U8866 (N_8866,N_8691,N_8664);
nor U8867 (N_8867,N_8605,N_8722);
xnor U8868 (N_8868,N_8689,N_8701);
or U8869 (N_8869,N_8674,N_8785);
xnor U8870 (N_8870,N_8683,N_8633);
or U8871 (N_8871,N_8681,N_8749);
nor U8872 (N_8872,N_8714,N_8794);
nor U8873 (N_8873,N_8751,N_8742);
and U8874 (N_8874,N_8704,N_8758);
nor U8875 (N_8875,N_8611,N_8685);
or U8876 (N_8876,N_8652,N_8706);
or U8877 (N_8877,N_8699,N_8651);
nor U8878 (N_8878,N_8613,N_8673);
and U8879 (N_8879,N_8614,N_8781);
and U8880 (N_8880,N_8700,N_8607);
and U8881 (N_8881,N_8746,N_8655);
and U8882 (N_8882,N_8694,N_8610);
nand U8883 (N_8883,N_8777,N_8752);
and U8884 (N_8884,N_8748,N_8717);
xor U8885 (N_8885,N_8739,N_8745);
nor U8886 (N_8886,N_8732,N_8759);
or U8887 (N_8887,N_8754,N_8728);
nand U8888 (N_8888,N_8735,N_8618);
nand U8889 (N_8889,N_8705,N_8679);
and U8890 (N_8890,N_8608,N_8686);
and U8891 (N_8891,N_8778,N_8629);
or U8892 (N_8892,N_8672,N_8798);
or U8893 (N_8893,N_8741,N_8771);
nor U8894 (N_8894,N_8719,N_8684);
or U8895 (N_8895,N_8622,N_8692);
nand U8896 (N_8896,N_8775,N_8765);
or U8897 (N_8897,N_8736,N_8698);
nor U8898 (N_8898,N_8676,N_8628);
nor U8899 (N_8899,N_8713,N_8784);
and U8900 (N_8900,N_8752,N_8622);
and U8901 (N_8901,N_8781,N_8636);
nand U8902 (N_8902,N_8736,N_8657);
or U8903 (N_8903,N_8681,N_8698);
nor U8904 (N_8904,N_8762,N_8634);
or U8905 (N_8905,N_8655,N_8677);
nand U8906 (N_8906,N_8774,N_8768);
xnor U8907 (N_8907,N_8681,N_8605);
or U8908 (N_8908,N_8677,N_8627);
xor U8909 (N_8909,N_8626,N_8685);
nor U8910 (N_8910,N_8753,N_8681);
nand U8911 (N_8911,N_8668,N_8771);
nor U8912 (N_8912,N_8736,N_8691);
xnor U8913 (N_8913,N_8732,N_8641);
or U8914 (N_8914,N_8778,N_8754);
or U8915 (N_8915,N_8753,N_8677);
or U8916 (N_8916,N_8785,N_8630);
and U8917 (N_8917,N_8702,N_8620);
nor U8918 (N_8918,N_8632,N_8710);
nand U8919 (N_8919,N_8623,N_8699);
and U8920 (N_8920,N_8639,N_8787);
nor U8921 (N_8921,N_8682,N_8734);
nand U8922 (N_8922,N_8694,N_8751);
or U8923 (N_8923,N_8651,N_8696);
and U8924 (N_8924,N_8710,N_8725);
xor U8925 (N_8925,N_8612,N_8741);
nand U8926 (N_8926,N_8603,N_8676);
nor U8927 (N_8927,N_8742,N_8661);
nor U8928 (N_8928,N_8604,N_8746);
nand U8929 (N_8929,N_8647,N_8652);
and U8930 (N_8930,N_8787,N_8712);
nand U8931 (N_8931,N_8750,N_8679);
nand U8932 (N_8932,N_8704,N_8736);
nand U8933 (N_8933,N_8613,N_8697);
nor U8934 (N_8934,N_8629,N_8796);
xor U8935 (N_8935,N_8607,N_8647);
nor U8936 (N_8936,N_8762,N_8610);
or U8937 (N_8937,N_8740,N_8706);
and U8938 (N_8938,N_8650,N_8707);
or U8939 (N_8939,N_8632,N_8657);
nand U8940 (N_8940,N_8644,N_8732);
and U8941 (N_8941,N_8749,N_8652);
nand U8942 (N_8942,N_8645,N_8705);
nand U8943 (N_8943,N_8698,N_8642);
nand U8944 (N_8944,N_8689,N_8705);
and U8945 (N_8945,N_8730,N_8653);
nand U8946 (N_8946,N_8668,N_8644);
nor U8947 (N_8947,N_8757,N_8775);
and U8948 (N_8948,N_8644,N_8692);
xnor U8949 (N_8949,N_8700,N_8656);
and U8950 (N_8950,N_8659,N_8662);
and U8951 (N_8951,N_8799,N_8627);
or U8952 (N_8952,N_8717,N_8639);
and U8953 (N_8953,N_8704,N_8695);
nor U8954 (N_8954,N_8668,N_8614);
or U8955 (N_8955,N_8658,N_8684);
or U8956 (N_8956,N_8795,N_8615);
nor U8957 (N_8957,N_8667,N_8777);
and U8958 (N_8958,N_8764,N_8670);
and U8959 (N_8959,N_8669,N_8684);
or U8960 (N_8960,N_8729,N_8780);
or U8961 (N_8961,N_8703,N_8694);
nand U8962 (N_8962,N_8793,N_8780);
nor U8963 (N_8963,N_8622,N_8784);
or U8964 (N_8964,N_8609,N_8759);
and U8965 (N_8965,N_8696,N_8644);
xor U8966 (N_8966,N_8724,N_8689);
or U8967 (N_8967,N_8649,N_8706);
nand U8968 (N_8968,N_8763,N_8795);
nand U8969 (N_8969,N_8602,N_8796);
xnor U8970 (N_8970,N_8751,N_8701);
or U8971 (N_8971,N_8768,N_8751);
nor U8972 (N_8972,N_8721,N_8796);
or U8973 (N_8973,N_8695,N_8699);
nor U8974 (N_8974,N_8793,N_8614);
nand U8975 (N_8975,N_8782,N_8690);
nand U8976 (N_8976,N_8666,N_8755);
or U8977 (N_8977,N_8789,N_8651);
nand U8978 (N_8978,N_8636,N_8763);
nand U8979 (N_8979,N_8715,N_8733);
and U8980 (N_8980,N_8641,N_8779);
nand U8981 (N_8981,N_8604,N_8615);
nor U8982 (N_8982,N_8642,N_8726);
nor U8983 (N_8983,N_8733,N_8664);
or U8984 (N_8984,N_8705,N_8690);
and U8985 (N_8985,N_8630,N_8629);
or U8986 (N_8986,N_8681,N_8772);
and U8987 (N_8987,N_8674,N_8721);
and U8988 (N_8988,N_8734,N_8660);
nor U8989 (N_8989,N_8630,N_8719);
xor U8990 (N_8990,N_8799,N_8768);
or U8991 (N_8991,N_8669,N_8739);
and U8992 (N_8992,N_8797,N_8714);
or U8993 (N_8993,N_8751,N_8667);
nor U8994 (N_8994,N_8636,N_8638);
nand U8995 (N_8995,N_8610,N_8703);
or U8996 (N_8996,N_8712,N_8728);
nand U8997 (N_8997,N_8742,N_8715);
and U8998 (N_8998,N_8705,N_8713);
or U8999 (N_8999,N_8601,N_8787);
and U9000 (N_9000,N_8845,N_8956);
and U9001 (N_9001,N_8869,N_8808);
and U9002 (N_9002,N_8885,N_8862);
nand U9003 (N_9003,N_8897,N_8918);
and U9004 (N_9004,N_8855,N_8815);
xor U9005 (N_9005,N_8863,N_8802);
nand U9006 (N_9006,N_8858,N_8824);
and U9007 (N_9007,N_8905,N_8881);
and U9008 (N_9008,N_8819,N_8989);
nand U9009 (N_9009,N_8821,N_8875);
and U9010 (N_9010,N_8866,N_8960);
or U9011 (N_9011,N_8859,N_8830);
or U9012 (N_9012,N_8831,N_8916);
xnor U9013 (N_9013,N_8964,N_8877);
nor U9014 (N_9014,N_8857,N_8913);
nand U9015 (N_9015,N_8952,N_8828);
nor U9016 (N_9016,N_8986,N_8843);
or U9017 (N_9017,N_8864,N_8974);
nor U9018 (N_9018,N_8870,N_8871);
nor U9019 (N_9019,N_8908,N_8966);
nor U9020 (N_9020,N_8838,N_8963);
and U9021 (N_9021,N_8832,N_8940);
nand U9022 (N_9022,N_8874,N_8826);
or U9023 (N_9023,N_8879,N_8817);
nand U9024 (N_9024,N_8903,N_8933);
and U9025 (N_9025,N_8810,N_8853);
nand U9026 (N_9026,N_8997,N_8920);
or U9027 (N_9027,N_8892,N_8809);
or U9028 (N_9028,N_8948,N_8803);
nand U9029 (N_9029,N_8900,N_8910);
xor U9030 (N_9030,N_8833,N_8822);
and U9031 (N_9031,N_8856,N_8927);
and U9032 (N_9032,N_8851,N_8829);
and U9033 (N_9033,N_8827,N_8931);
or U9034 (N_9034,N_8939,N_8899);
nand U9035 (N_9035,N_8949,N_8847);
and U9036 (N_9036,N_8812,N_8806);
nor U9037 (N_9037,N_8891,N_8995);
and U9038 (N_9038,N_8898,N_8893);
nand U9039 (N_9039,N_8981,N_8975);
or U9040 (N_9040,N_8965,N_8996);
and U9041 (N_9041,N_8932,N_8991);
or U9042 (N_9042,N_8883,N_8912);
nand U9043 (N_9043,N_8800,N_8902);
nand U9044 (N_9044,N_8816,N_8923);
or U9045 (N_9045,N_8985,N_8814);
nor U9046 (N_9046,N_8841,N_8839);
and U9047 (N_9047,N_8994,N_8926);
nand U9048 (N_9048,N_8867,N_8888);
and U9049 (N_9049,N_8872,N_8961);
and U9050 (N_9050,N_8970,N_8811);
nor U9051 (N_9051,N_8894,N_8852);
and U9052 (N_9052,N_8942,N_8895);
nand U9053 (N_9053,N_8880,N_8835);
nor U9054 (N_9054,N_8917,N_8947);
xnor U9055 (N_9055,N_8825,N_8954);
nand U9056 (N_9056,N_8882,N_8876);
or U9057 (N_9057,N_8924,N_8935);
or U9058 (N_9058,N_8983,N_8951);
or U9059 (N_9059,N_8909,N_8848);
nor U9060 (N_9060,N_8896,N_8907);
and U9061 (N_9061,N_8801,N_8890);
or U9062 (N_9062,N_8937,N_8849);
nor U9063 (N_9063,N_8968,N_8976);
or U9064 (N_9064,N_8837,N_8958);
or U9065 (N_9065,N_8805,N_8928);
xor U9066 (N_9066,N_8915,N_8930);
or U9067 (N_9067,N_8969,N_8868);
or U9068 (N_9068,N_8984,N_8988);
nor U9069 (N_9069,N_8906,N_8934);
nand U9070 (N_9070,N_8914,N_8901);
nand U9071 (N_9071,N_8955,N_8804);
nand U9072 (N_9072,N_8818,N_8998);
nand U9073 (N_9073,N_8943,N_8921);
nor U9074 (N_9074,N_8938,N_8957);
and U9075 (N_9075,N_8945,N_8950);
or U9076 (N_9076,N_8944,N_8844);
and U9077 (N_9077,N_8846,N_8865);
and U9078 (N_9078,N_8886,N_8962);
nor U9079 (N_9079,N_8953,N_8959);
nand U9080 (N_9080,N_8823,N_8836);
or U9081 (N_9081,N_8904,N_8990);
nand U9082 (N_9082,N_8929,N_8987);
nor U9083 (N_9083,N_8925,N_8861);
xor U9084 (N_9084,N_8941,N_8873);
nand U9085 (N_9085,N_8993,N_8911);
xnor U9086 (N_9086,N_8889,N_8936);
or U9087 (N_9087,N_8813,N_8967);
nand U9088 (N_9088,N_8834,N_8887);
or U9089 (N_9089,N_8946,N_8884);
and U9090 (N_9090,N_8878,N_8854);
nor U9091 (N_9091,N_8978,N_8979);
and U9092 (N_9092,N_8977,N_8842);
nor U9093 (N_9093,N_8973,N_8999);
nand U9094 (N_9094,N_8807,N_8992);
nand U9095 (N_9095,N_8980,N_8840);
nor U9096 (N_9096,N_8850,N_8972);
nor U9097 (N_9097,N_8860,N_8820);
and U9098 (N_9098,N_8922,N_8982);
nor U9099 (N_9099,N_8971,N_8919);
nor U9100 (N_9100,N_8949,N_8839);
or U9101 (N_9101,N_8864,N_8885);
or U9102 (N_9102,N_8902,N_8823);
and U9103 (N_9103,N_8862,N_8894);
and U9104 (N_9104,N_8999,N_8941);
nor U9105 (N_9105,N_8974,N_8861);
or U9106 (N_9106,N_8877,N_8933);
xnor U9107 (N_9107,N_8927,N_8954);
xnor U9108 (N_9108,N_8977,N_8865);
or U9109 (N_9109,N_8859,N_8974);
or U9110 (N_9110,N_8905,N_8945);
or U9111 (N_9111,N_8997,N_8885);
nand U9112 (N_9112,N_8814,N_8876);
nor U9113 (N_9113,N_8994,N_8921);
nor U9114 (N_9114,N_8946,N_8939);
or U9115 (N_9115,N_8808,N_8862);
nand U9116 (N_9116,N_8982,N_8938);
nor U9117 (N_9117,N_8899,N_8968);
and U9118 (N_9118,N_8825,N_8987);
nand U9119 (N_9119,N_8975,N_8927);
nor U9120 (N_9120,N_8848,N_8925);
nand U9121 (N_9121,N_8900,N_8849);
and U9122 (N_9122,N_8805,N_8821);
and U9123 (N_9123,N_8988,N_8800);
and U9124 (N_9124,N_8950,N_8941);
or U9125 (N_9125,N_8820,N_8958);
or U9126 (N_9126,N_8853,N_8824);
and U9127 (N_9127,N_8887,N_8906);
or U9128 (N_9128,N_8984,N_8925);
xnor U9129 (N_9129,N_8930,N_8926);
nor U9130 (N_9130,N_8818,N_8857);
or U9131 (N_9131,N_8814,N_8800);
xor U9132 (N_9132,N_8921,N_8898);
and U9133 (N_9133,N_8825,N_8958);
nor U9134 (N_9134,N_8817,N_8807);
nand U9135 (N_9135,N_8886,N_8905);
nand U9136 (N_9136,N_8884,N_8849);
nor U9137 (N_9137,N_8902,N_8947);
or U9138 (N_9138,N_8801,N_8903);
nand U9139 (N_9139,N_8909,N_8979);
nand U9140 (N_9140,N_8985,N_8839);
nor U9141 (N_9141,N_8817,N_8928);
nand U9142 (N_9142,N_8841,N_8855);
and U9143 (N_9143,N_8980,N_8995);
nor U9144 (N_9144,N_8822,N_8930);
nor U9145 (N_9145,N_8826,N_8829);
and U9146 (N_9146,N_8985,N_8943);
or U9147 (N_9147,N_8816,N_8821);
and U9148 (N_9148,N_8823,N_8934);
nand U9149 (N_9149,N_8858,N_8831);
nand U9150 (N_9150,N_8862,N_8961);
nand U9151 (N_9151,N_8942,N_8866);
nand U9152 (N_9152,N_8807,N_8943);
nand U9153 (N_9153,N_8899,N_8813);
or U9154 (N_9154,N_8991,N_8931);
nor U9155 (N_9155,N_8849,N_8847);
or U9156 (N_9156,N_8859,N_8994);
nor U9157 (N_9157,N_8984,N_8869);
or U9158 (N_9158,N_8814,N_8865);
nand U9159 (N_9159,N_8839,N_8886);
nand U9160 (N_9160,N_8875,N_8995);
nand U9161 (N_9161,N_8923,N_8992);
and U9162 (N_9162,N_8927,N_8895);
or U9163 (N_9163,N_8867,N_8881);
or U9164 (N_9164,N_8944,N_8875);
nor U9165 (N_9165,N_8998,N_8967);
nand U9166 (N_9166,N_8898,N_8900);
and U9167 (N_9167,N_8800,N_8970);
and U9168 (N_9168,N_8904,N_8975);
and U9169 (N_9169,N_8979,N_8995);
nor U9170 (N_9170,N_8993,N_8826);
and U9171 (N_9171,N_8922,N_8928);
nor U9172 (N_9172,N_8851,N_8807);
and U9173 (N_9173,N_8950,N_8983);
nand U9174 (N_9174,N_8823,N_8983);
or U9175 (N_9175,N_8995,N_8925);
and U9176 (N_9176,N_8915,N_8981);
nor U9177 (N_9177,N_8980,N_8941);
nand U9178 (N_9178,N_8991,N_8921);
or U9179 (N_9179,N_8897,N_8863);
or U9180 (N_9180,N_8887,N_8886);
nand U9181 (N_9181,N_8879,N_8901);
nor U9182 (N_9182,N_8955,N_8886);
or U9183 (N_9183,N_8848,N_8946);
and U9184 (N_9184,N_8875,N_8878);
nor U9185 (N_9185,N_8976,N_8902);
and U9186 (N_9186,N_8922,N_8947);
and U9187 (N_9187,N_8981,N_8873);
and U9188 (N_9188,N_8861,N_8990);
and U9189 (N_9189,N_8908,N_8881);
and U9190 (N_9190,N_8903,N_8958);
or U9191 (N_9191,N_8835,N_8969);
or U9192 (N_9192,N_8852,N_8990);
and U9193 (N_9193,N_8996,N_8832);
xor U9194 (N_9194,N_8848,N_8921);
nand U9195 (N_9195,N_8830,N_8874);
nand U9196 (N_9196,N_8877,N_8996);
xnor U9197 (N_9197,N_8913,N_8936);
and U9198 (N_9198,N_8895,N_8821);
or U9199 (N_9199,N_8962,N_8915);
nand U9200 (N_9200,N_9077,N_9060);
nor U9201 (N_9201,N_9174,N_9169);
or U9202 (N_9202,N_9190,N_9115);
nor U9203 (N_9203,N_9170,N_9024);
nor U9204 (N_9204,N_9092,N_9029);
and U9205 (N_9205,N_9026,N_9096);
and U9206 (N_9206,N_9013,N_9117);
or U9207 (N_9207,N_9030,N_9078);
nand U9208 (N_9208,N_9059,N_9016);
nor U9209 (N_9209,N_9017,N_9146);
xor U9210 (N_9210,N_9104,N_9116);
nor U9211 (N_9211,N_9139,N_9186);
or U9212 (N_9212,N_9152,N_9006);
nor U9213 (N_9213,N_9185,N_9130);
or U9214 (N_9214,N_9121,N_9122);
or U9215 (N_9215,N_9074,N_9001);
or U9216 (N_9216,N_9015,N_9157);
nand U9217 (N_9217,N_9008,N_9133);
nor U9218 (N_9218,N_9011,N_9056);
nand U9219 (N_9219,N_9173,N_9064);
nor U9220 (N_9220,N_9176,N_9161);
nand U9221 (N_9221,N_9098,N_9093);
or U9222 (N_9222,N_9196,N_9166);
and U9223 (N_9223,N_9079,N_9076);
and U9224 (N_9224,N_9073,N_9182);
nand U9225 (N_9225,N_9109,N_9007);
xor U9226 (N_9226,N_9118,N_9183);
and U9227 (N_9227,N_9087,N_9199);
and U9228 (N_9228,N_9113,N_9034);
nor U9229 (N_9229,N_9036,N_9031);
and U9230 (N_9230,N_9153,N_9102);
or U9231 (N_9231,N_9197,N_9151);
and U9232 (N_9232,N_9163,N_9108);
nand U9233 (N_9233,N_9189,N_9136);
or U9234 (N_9234,N_9179,N_9148);
or U9235 (N_9235,N_9042,N_9062);
or U9236 (N_9236,N_9039,N_9123);
and U9237 (N_9237,N_9090,N_9019);
nand U9238 (N_9238,N_9167,N_9111);
and U9239 (N_9239,N_9072,N_9050);
or U9240 (N_9240,N_9069,N_9014);
nand U9241 (N_9241,N_9112,N_9103);
xor U9242 (N_9242,N_9131,N_9054);
or U9243 (N_9243,N_9192,N_9106);
xor U9244 (N_9244,N_9178,N_9175);
or U9245 (N_9245,N_9184,N_9158);
and U9246 (N_9246,N_9028,N_9124);
and U9247 (N_9247,N_9127,N_9048);
nand U9248 (N_9248,N_9097,N_9162);
nor U9249 (N_9249,N_9101,N_9081);
nor U9250 (N_9250,N_9140,N_9107);
and U9251 (N_9251,N_9128,N_9126);
nand U9252 (N_9252,N_9181,N_9145);
nand U9253 (N_9253,N_9149,N_9177);
nand U9254 (N_9254,N_9194,N_9114);
and U9255 (N_9255,N_9000,N_9047);
and U9256 (N_9256,N_9100,N_9094);
nor U9257 (N_9257,N_9082,N_9105);
and U9258 (N_9258,N_9044,N_9010);
nor U9259 (N_9259,N_9053,N_9080);
xor U9260 (N_9260,N_9052,N_9132);
or U9261 (N_9261,N_9003,N_9041);
nor U9262 (N_9262,N_9051,N_9049);
nand U9263 (N_9263,N_9119,N_9063);
nor U9264 (N_9264,N_9020,N_9091);
and U9265 (N_9265,N_9023,N_9171);
and U9266 (N_9266,N_9075,N_9004);
or U9267 (N_9267,N_9055,N_9156);
nor U9268 (N_9268,N_9038,N_9138);
or U9269 (N_9269,N_9022,N_9160);
or U9270 (N_9270,N_9021,N_9180);
or U9271 (N_9271,N_9095,N_9187);
and U9272 (N_9272,N_9089,N_9099);
nor U9273 (N_9273,N_9012,N_9172);
and U9274 (N_9274,N_9033,N_9058);
or U9275 (N_9275,N_9110,N_9065);
and U9276 (N_9276,N_9088,N_9046);
nor U9277 (N_9277,N_9134,N_9195);
and U9278 (N_9278,N_9129,N_9018);
and U9279 (N_9279,N_9120,N_9085);
nand U9280 (N_9280,N_9198,N_9070);
nand U9281 (N_9281,N_9040,N_9043);
or U9282 (N_9282,N_9168,N_9150);
nand U9283 (N_9283,N_9188,N_9032);
nand U9284 (N_9284,N_9141,N_9057);
nand U9285 (N_9285,N_9035,N_9191);
and U9286 (N_9286,N_9002,N_9027);
and U9287 (N_9287,N_9193,N_9135);
and U9288 (N_9288,N_9045,N_9083);
and U9289 (N_9289,N_9067,N_9009);
nor U9290 (N_9290,N_9165,N_9142);
or U9291 (N_9291,N_9005,N_9143);
and U9292 (N_9292,N_9086,N_9137);
nand U9293 (N_9293,N_9154,N_9144);
or U9294 (N_9294,N_9084,N_9125);
and U9295 (N_9295,N_9061,N_9155);
and U9296 (N_9296,N_9159,N_9164);
or U9297 (N_9297,N_9068,N_9025);
nor U9298 (N_9298,N_9071,N_9037);
nor U9299 (N_9299,N_9147,N_9066);
xor U9300 (N_9300,N_9188,N_9162);
nor U9301 (N_9301,N_9163,N_9151);
nor U9302 (N_9302,N_9073,N_9009);
or U9303 (N_9303,N_9196,N_9064);
xnor U9304 (N_9304,N_9189,N_9110);
nor U9305 (N_9305,N_9153,N_9049);
and U9306 (N_9306,N_9124,N_9056);
or U9307 (N_9307,N_9001,N_9136);
or U9308 (N_9308,N_9066,N_9035);
or U9309 (N_9309,N_9018,N_9062);
nand U9310 (N_9310,N_9117,N_9054);
nor U9311 (N_9311,N_9179,N_9015);
or U9312 (N_9312,N_9163,N_9158);
nand U9313 (N_9313,N_9093,N_9060);
or U9314 (N_9314,N_9161,N_9194);
and U9315 (N_9315,N_9075,N_9118);
xor U9316 (N_9316,N_9055,N_9128);
and U9317 (N_9317,N_9054,N_9114);
nand U9318 (N_9318,N_9028,N_9022);
or U9319 (N_9319,N_9192,N_9008);
nor U9320 (N_9320,N_9175,N_9112);
and U9321 (N_9321,N_9095,N_9171);
nor U9322 (N_9322,N_9093,N_9089);
nor U9323 (N_9323,N_9009,N_9011);
or U9324 (N_9324,N_9141,N_9166);
xor U9325 (N_9325,N_9080,N_9079);
and U9326 (N_9326,N_9095,N_9088);
xnor U9327 (N_9327,N_9060,N_9053);
nand U9328 (N_9328,N_9105,N_9150);
and U9329 (N_9329,N_9165,N_9164);
nand U9330 (N_9330,N_9151,N_9031);
nand U9331 (N_9331,N_9146,N_9071);
nand U9332 (N_9332,N_9171,N_9112);
or U9333 (N_9333,N_9153,N_9175);
or U9334 (N_9334,N_9090,N_9031);
or U9335 (N_9335,N_9041,N_9105);
and U9336 (N_9336,N_9148,N_9047);
nand U9337 (N_9337,N_9017,N_9057);
nor U9338 (N_9338,N_9196,N_9090);
nor U9339 (N_9339,N_9031,N_9042);
or U9340 (N_9340,N_9100,N_9189);
nor U9341 (N_9341,N_9135,N_9011);
and U9342 (N_9342,N_9046,N_9064);
nor U9343 (N_9343,N_9192,N_9060);
or U9344 (N_9344,N_9110,N_9179);
or U9345 (N_9345,N_9076,N_9120);
nand U9346 (N_9346,N_9052,N_9144);
and U9347 (N_9347,N_9113,N_9155);
nand U9348 (N_9348,N_9027,N_9150);
and U9349 (N_9349,N_9170,N_9138);
or U9350 (N_9350,N_9089,N_9155);
nand U9351 (N_9351,N_9092,N_9182);
and U9352 (N_9352,N_9096,N_9186);
nand U9353 (N_9353,N_9027,N_9095);
nand U9354 (N_9354,N_9003,N_9044);
nor U9355 (N_9355,N_9006,N_9033);
and U9356 (N_9356,N_9099,N_9034);
nand U9357 (N_9357,N_9172,N_9074);
xor U9358 (N_9358,N_9156,N_9036);
or U9359 (N_9359,N_9107,N_9169);
and U9360 (N_9360,N_9046,N_9087);
nand U9361 (N_9361,N_9144,N_9177);
nor U9362 (N_9362,N_9158,N_9077);
and U9363 (N_9363,N_9119,N_9076);
and U9364 (N_9364,N_9169,N_9081);
nand U9365 (N_9365,N_9194,N_9186);
or U9366 (N_9366,N_9014,N_9094);
xnor U9367 (N_9367,N_9123,N_9076);
or U9368 (N_9368,N_9053,N_9158);
nand U9369 (N_9369,N_9141,N_9104);
nand U9370 (N_9370,N_9097,N_9058);
nor U9371 (N_9371,N_9170,N_9142);
xnor U9372 (N_9372,N_9166,N_9165);
xnor U9373 (N_9373,N_9133,N_9018);
nand U9374 (N_9374,N_9162,N_9019);
nor U9375 (N_9375,N_9171,N_9137);
or U9376 (N_9376,N_9120,N_9083);
xor U9377 (N_9377,N_9093,N_9189);
nor U9378 (N_9378,N_9046,N_9152);
and U9379 (N_9379,N_9156,N_9048);
or U9380 (N_9380,N_9028,N_9130);
xnor U9381 (N_9381,N_9053,N_9097);
and U9382 (N_9382,N_9020,N_9118);
or U9383 (N_9383,N_9092,N_9181);
and U9384 (N_9384,N_9097,N_9018);
and U9385 (N_9385,N_9192,N_9139);
and U9386 (N_9386,N_9155,N_9002);
xor U9387 (N_9387,N_9157,N_9050);
nor U9388 (N_9388,N_9030,N_9149);
nand U9389 (N_9389,N_9100,N_9084);
nor U9390 (N_9390,N_9052,N_9187);
nand U9391 (N_9391,N_9084,N_9115);
nand U9392 (N_9392,N_9172,N_9083);
or U9393 (N_9393,N_9175,N_9090);
nor U9394 (N_9394,N_9194,N_9043);
and U9395 (N_9395,N_9133,N_9140);
and U9396 (N_9396,N_9104,N_9053);
nor U9397 (N_9397,N_9016,N_9055);
and U9398 (N_9398,N_9173,N_9038);
xor U9399 (N_9399,N_9124,N_9022);
nand U9400 (N_9400,N_9340,N_9285);
nor U9401 (N_9401,N_9282,N_9249);
nor U9402 (N_9402,N_9217,N_9225);
or U9403 (N_9403,N_9355,N_9316);
and U9404 (N_9404,N_9378,N_9286);
nor U9405 (N_9405,N_9243,N_9254);
nand U9406 (N_9406,N_9326,N_9364);
and U9407 (N_9407,N_9374,N_9244);
and U9408 (N_9408,N_9226,N_9229);
or U9409 (N_9409,N_9222,N_9291);
nand U9410 (N_9410,N_9308,N_9256);
or U9411 (N_9411,N_9344,N_9269);
nand U9412 (N_9412,N_9330,N_9230);
nor U9413 (N_9413,N_9359,N_9204);
nor U9414 (N_9414,N_9306,N_9370);
or U9415 (N_9415,N_9305,N_9303);
xnor U9416 (N_9416,N_9311,N_9373);
and U9417 (N_9417,N_9283,N_9358);
nor U9418 (N_9418,N_9208,N_9383);
nor U9419 (N_9419,N_9272,N_9346);
and U9420 (N_9420,N_9251,N_9267);
and U9421 (N_9421,N_9264,N_9381);
and U9422 (N_9422,N_9270,N_9260);
nor U9423 (N_9423,N_9376,N_9337);
xnor U9424 (N_9424,N_9266,N_9261);
xor U9425 (N_9425,N_9362,N_9331);
or U9426 (N_9426,N_9221,N_9371);
nor U9427 (N_9427,N_9307,N_9312);
or U9428 (N_9428,N_9388,N_9257);
and U9429 (N_9429,N_9333,N_9252);
nor U9430 (N_9430,N_9369,N_9295);
nor U9431 (N_9431,N_9253,N_9367);
nand U9432 (N_9432,N_9321,N_9339);
nor U9433 (N_9433,N_9353,N_9209);
nor U9434 (N_9434,N_9350,N_9317);
and U9435 (N_9435,N_9259,N_9396);
or U9436 (N_9436,N_9268,N_9345);
and U9437 (N_9437,N_9386,N_9233);
nor U9438 (N_9438,N_9223,N_9352);
nand U9439 (N_9439,N_9319,N_9245);
nand U9440 (N_9440,N_9284,N_9368);
or U9441 (N_9441,N_9384,N_9277);
xnor U9442 (N_9442,N_9336,N_9275);
nor U9443 (N_9443,N_9310,N_9382);
nor U9444 (N_9444,N_9315,N_9292);
or U9445 (N_9445,N_9356,N_9335);
and U9446 (N_9446,N_9342,N_9318);
xor U9447 (N_9447,N_9372,N_9273);
nand U9448 (N_9448,N_9296,N_9361);
nand U9449 (N_9449,N_9320,N_9328);
nand U9450 (N_9450,N_9236,N_9322);
or U9451 (N_9451,N_9218,N_9231);
and U9452 (N_9452,N_9325,N_9232);
nand U9453 (N_9453,N_9343,N_9302);
or U9454 (N_9454,N_9366,N_9389);
nor U9455 (N_9455,N_9250,N_9262);
and U9456 (N_9456,N_9215,N_9280);
and U9457 (N_9457,N_9298,N_9324);
and U9458 (N_9458,N_9313,N_9309);
nor U9459 (N_9459,N_9246,N_9347);
nand U9460 (N_9460,N_9348,N_9294);
and U9461 (N_9461,N_9227,N_9274);
and U9462 (N_9462,N_9379,N_9341);
nand U9463 (N_9463,N_9203,N_9354);
nand U9464 (N_9464,N_9293,N_9220);
nand U9465 (N_9465,N_9202,N_9242);
xnor U9466 (N_9466,N_9357,N_9281);
nor U9467 (N_9467,N_9216,N_9332);
or U9468 (N_9468,N_9210,N_9394);
xnor U9469 (N_9469,N_9314,N_9228);
nand U9470 (N_9470,N_9327,N_9391);
nand U9471 (N_9471,N_9237,N_9329);
and U9472 (N_9472,N_9206,N_9279);
xor U9473 (N_9473,N_9290,N_9397);
or U9474 (N_9474,N_9239,N_9399);
nand U9475 (N_9475,N_9240,N_9258);
nor U9476 (N_9476,N_9301,N_9271);
nor U9477 (N_9477,N_9392,N_9263);
or U9478 (N_9478,N_9289,N_9234);
nand U9479 (N_9479,N_9213,N_9377);
nand U9480 (N_9480,N_9276,N_9360);
nor U9481 (N_9481,N_9255,N_9211);
or U9482 (N_9482,N_9287,N_9398);
and U9483 (N_9483,N_9200,N_9390);
or U9484 (N_9484,N_9395,N_9238);
and U9485 (N_9485,N_9365,N_9393);
or U9486 (N_9486,N_9334,N_9278);
and U9487 (N_9487,N_9380,N_9338);
or U9488 (N_9488,N_9349,N_9385);
or U9489 (N_9489,N_9205,N_9299);
nor U9490 (N_9490,N_9304,N_9300);
or U9491 (N_9491,N_9224,N_9248);
nand U9492 (N_9492,N_9235,N_9323);
nand U9493 (N_9493,N_9207,N_9297);
or U9494 (N_9494,N_9212,N_9219);
nor U9495 (N_9495,N_9201,N_9375);
and U9496 (N_9496,N_9351,N_9288);
nand U9497 (N_9497,N_9214,N_9363);
and U9498 (N_9498,N_9241,N_9247);
and U9499 (N_9499,N_9387,N_9265);
or U9500 (N_9500,N_9396,N_9319);
nand U9501 (N_9501,N_9322,N_9345);
or U9502 (N_9502,N_9354,N_9396);
nand U9503 (N_9503,N_9228,N_9208);
nor U9504 (N_9504,N_9322,N_9203);
or U9505 (N_9505,N_9279,N_9231);
nor U9506 (N_9506,N_9295,N_9236);
and U9507 (N_9507,N_9381,N_9272);
nor U9508 (N_9508,N_9324,N_9218);
or U9509 (N_9509,N_9367,N_9249);
or U9510 (N_9510,N_9242,N_9232);
or U9511 (N_9511,N_9217,N_9356);
nor U9512 (N_9512,N_9357,N_9256);
nand U9513 (N_9513,N_9209,N_9264);
or U9514 (N_9514,N_9202,N_9393);
nand U9515 (N_9515,N_9227,N_9264);
nand U9516 (N_9516,N_9300,N_9213);
or U9517 (N_9517,N_9360,N_9271);
or U9518 (N_9518,N_9294,N_9253);
and U9519 (N_9519,N_9276,N_9329);
xnor U9520 (N_9520,N_9246,N_9292);
nand U9521 (N_9521,N_9346,N_9292);
nor U9522 (N_9522,N_9323,N_9204);
and U9523 (N_9523,N_9272,N_9212);
nor U9524 (N_9524,N_9334,N_9229);
or U9525 (N_9525,N_9203,N_9358);
nand U9526 (N_9526,N_9377,N_9274);
nor U9527 (N_9527,N_9297,N_9261);
and U9528 (N_9528,N_9297,N_9396);
and U9529 (N_9529,N_9330,N_9342);
nand U9530 (N_9530,N_9271,N_9366);
or U9531 (N_9531,N_9317,N_9336);
and U9532 (N_9532,N_9342,N_9258);
nand U9533 (N_9533,N_9257,N_9334);
or U9534 (N_9534,N_9308,N_9392);
nand U9535 (N_9535,N_9368,N_9209);
or U9536 (N_9536,N_9359,N_9298);
nor U9537 (N_9537,N_9315,N_9205);
or U9538 (N_9538,N_9216,N_9380);
and U9539 (N_9539,N_9335,N_9299);
nand U9540 (N_9540,N_9396,N_9272);
nand U9541 (N_9541,N_9245,N_9296);
nor U9542 (N_9542,N_9213,N_9256);
nor U9543 (N_9543,N_9222,N_9282);
nand U9544 (N_9544,N_9279,N_9275);
and U9545 (N_9545,N_9265,N_9257);
xor U9546 (N_9546,N_9286,N_9335);
nand U9547 (N_9547,N_9365,N_9355);
or U9548 (N_9548,N_9368,N_9355);
and U9549 (N_9549,N_9271,N_9270);
nand U9550 (N_9550,N_9240,N_9318);
xor U9551 (N_9551,N_9307,N_9241);
xnor U9552 (N_9552,N_9323,N_9389);
nand U9553 (N_9553,N_9341,N_9303);
and U9554 (N_9554,N_9251,N_9338);
nand U9555 (N_9555,N_9354,N_9243);
and U9556 (N_9556,N_9363,N_9212);
xor U9557 (N_9557,N_9311,N_9366);
nand U9558 (N_9558,N_9349,N_9381);
or U9559 (N_9559,N_9293,N_9258);
or U9560 (N_9560,N_9226,N_9315);
nand U9561 (N_9561,N_9247,N_9244);
nand U9562 (N_9562,N_9392,N_9209);
nor U9563 (N_9563,N_9212,N_9283);
or U9564 (N_9564,N_9324,N_9313);
or U9565 (N_9565,N_9213,N_9313);
or U9566 (N_9566,N_9309,N_9391);
nand U9567 (N_9567,N_9369,N_9269);
and U9568 (N_9568,N_9257,N_9360);
or U9569 (N_9569,N_9374,N_9352);
nor U9570 (N_9570,N_9276,N_9283);
nor U9571 (N_9571,N_9249,N_9372);
or U9572 (N_9572,N_9202,N_9318);
or U9573 (N_9573,N_9297,N_9282);
nor U9574 (N_9574,N_9329,N_9397);
nand U9575 (N_9575,N_9314,N_9307);
xnor U9576 (N_9576,N_9370,N_9389);
nand U9577 (N_9577,N_9369,N_9312);
or U9578 (N_9578,N_9269,N_9382);
and U9579 (N_9579,N_9357,N_9311);
or U9580 (N_9580,N_9210,N_9267);
nor U9581 (N_9581,N_9234,N_9219);
nand U9582 (N_9582,N_9316,N_9328);
nor U9583 (N_9583,N_9257,N_9339);
nand U9584 (N_9584,N_9398,N_9302);
nor U9585 (N_9585,N_9242,N_9341);
and U9586 (N_9586,N_9245,N_9264);
or U9587 (N_9587,N_9284,N_9321);
nand U9588 (N_9588,N_9207,N_9284);
or U9589 (N_9589,N_9264,N_9260);
nor U9590 (N_9590,N_9342,N_9227);
nor U9591 (N_9591,N_9238,N_9333);
and U9592 (N_9592,N_9312,N_9334);
and U9593 (N_9593,N_9371,N_9249);
nand U9594 (N_9594,N_9241,N_9311);
nor U9595 (N_9595,N_9244,N_9390);
nor U9596 (N_9596,N_9201,N_9335);
nor U9597 (N_9597,N_9311,N_9276);
xnor U9598 (N_9598,N_9223,N_9380);
or U9599 (N_9599,N_9252,N_9215);
and U9600 (N_9600,N_9446,N_9453);
nor U9601 (N_9601,N_9445,N_9413);
nand U9602 (N_9602,N_9555,N_9546);
xnor U9603 (N_9603,N_9507,N_9571);
nand U9604 (N_9604,N_9545,N_9462);
nand U9605 (N_9605,N_9414,N_9549);
nand U9606 (N_9606,N_9557,N_9518);
and U9607 (N_9607,N_9538,N_9592);
and U9608 (N_9608,N_9455,N_9520);
and U9609 (N_9609,N_9466,N_9457);
and U9610 (N_9610,N_9500,N_9512);
nand U9611 (N_9611,N_9409,N_9437);
and U9612 (N_9612,N_9493,N_9495);
and U9613 (N_9613,N_9450,N_9548);
nand U9614 (N_9614,N_9406,N_9532);
and U9615 (N_9615,N_9432,N_9528);
nor U9616 (N_9616,N_9465,N_9519);
nand U9617 (N_9617,N_9561,N_9496);
and U9618 (N_9618,N_9475,N_9584);
nand U9619 (N_9619,N_9476,N_9568);
or U9620 (N_9620,N_9580,N_9436);
xnor U9621 (N_9621,N_9504,N_9411);
and U9622 (N_9622,N_9408,N_9425);
or U9623 (N_9623,N_9560,N_9422);
and U9624 (N_9624,N_9569,N_9575);
or U9625 (N_9625,N_9439,N_9481);
nor U9626 (N_9626,N_9535,N_9435);
nand U9627 (N_9627,N_9442,N_9428);
nor U9628 (N_9628,N_9407,N_9487);
xnor U9629 (N_9629,N_9521,N_9524);
nand U9630 (N_9630,N_9451,N_9485);
nor U9631 (N_9631,N_9574,N_9567);
and U9632 (N_9632,N_9576,N_9539);
or U9633 (N_9633,N_9597,N_9591);
and U9634 (N_9634,N_9492,N_9410);
or U9635 (N_9635,N_9426,N_9564);
nand U9636 (N_9636,N_9404,N_9563);
and U9637 (N_9637,N_9578,N_9460);
and U9638 (N_9638,N_9582,N_9506);
nand U9639 (N_9639,N_9483,N_9478);
or U9640 (N_9640,N_9551,N_9447);
or U9641 (N_9641,N_9470,N_9438);
nor U9642 (N_9642,N_9531,N_9522);
nor U9643 (N_9643,N_9468,N_9456);
nand U9644 (N_9644,N_9565,N_9527);
and U9645 (N_9645,N_9441,N_9430);
and U9646 (N_9646,N_9431,N_9523);
nor U9647 (N_9647,N_9547,N_9402);
nand U9648 (N_9648,N_9590,N_9572);
and U9649 (N_9649,N_9443,N_9554);
nor U9650 (N_9650,N_9508,N_9467);
nor U9651 (N_9651,N_9585,N_9544);
nand U9652 (N_9652,N_9513,N_9434);
or U9653 (N_9653,N_9530,N_9461);
and U9654 (N_9654,N_9577,N_9490);
or U9655 (N_9655,N_9494,N_9525);
nor U9656 (N_9656,N_9593,N_9499);
or U9657 (N_9657,N_9403,N_9594);
nand U9658 (N_9658,N_9526,N_9503);
nor U9659 (N_9659,N_9480,N_9579);
nor U9660 (N_9660,N_9598,N_9473);
or U9661 (N_9661,N_9484,N_9449);
nand U9662 (N_9662,N_9540,N_9553);
and U9663 (N_9663,N_9558,N_9536);
or U9664 (N_9664,N_9501,N_9587);
or U9665 (N_9665,N_9534,N_9550);
or U9666 (N_9666,N_9542,N_9562);
nor U9667 (N_9667,N_9418,N_9498);
or U9668 (N_9668,N_9415,N_9529);
or U9669 (N_9669,N_9433,N_9488);
nand U9670 (N_9670,N_9589,N_9463);
and U9671 (N_9671,N_9416,N_9505);
xor U9672 (N_9672,N_9458,N_9552);
nor U9673 (N_9673,N_9556,N_9472);
or U9674 (N_9674,N_9595,N_9448);
or U9675 (N_9675,N_9429,N_9417);
nand U9676 (N_9676,N_9444,N_9452);
and U9677 (N_9677,N_9405,N_9479);
and U9678 (N_9678,N_9482,N_9516);
or U9679 (N_9679,N_9583,N_9537);
or U9680 (N_9680,N_9420,N_9454);
or U9681 (N_9681,N_9566,N_9486);
or U9682 (N_9682,N_9400,N_9497);
or U9683 (N_9683,N_9510,N_9427);
nand U9684 (N_9684,N_9533,N_9459);
nor U9685 (N_9685,N_9491,N_9509);
and U9686 (N_9686,N_9514,N_9401);
and U9687 (N_9687,N_9515,N_9517);
and U9688 (N_9688,N_9419,N_9421);
nand U9689 (N_9689,N_9502,N_9541);
nor U9690 (N_9690,N_9570,N_9596);
xnor U9691 (N_9691,N_9474,N_9412);
and U9692 (N_9692,N_9599,N_9588);
nor U9693 (N_9693,N_9489,N_9543);
and U9694 (N_9694,N_9559,N_9464);
nand U9695 (N_9695,N_9424,N_9581);
nor U9696 (N_9696,N_9573,N_9471);
nand U9697 (N_9697,N_9469,N_9423);
nand U9698 (N_9698,N_9586,N_9477);
xor U9699 (N_9699,N_9511,N_9440);
and U9700 (N_9700,N_9567,N_9441);
nand U9701 (N_9701,N_9554,N_9405);
and U9702 (N_9702,N_9447,N_9549);
xnor U9703 (N_9703,N_9492,N_9512);
and U9704 (N_9704,N_9590,N_9587);
and U9705 (N_9705,N_9549,N_9592);
nand U9706 (N_9706,N_9593,N_9592);
nand U9707 (N_9707,N_9471,N_9599);
xor U9708 (N_9708,N_9401,N_9490);
and U9709 (N_9709,N_9404,N_9519);
nand U9710 (N_9710,N_9510,N_9416);
and U9711 (N_9711,N_9402,N_9540);
nand U9712 (N_9712,N_9479,N_9473);
nand U9713 (N_9713,N_9528,N_9472);
nand U9714 (N_9714,N_9489,N_9556);
or U9715 (N_9715,N_9499,N_9469);
nor U9716 (N_9716,N_9531,N_9594);
nor U9717 (N_9717,N_9552,N_9403);
and U9718 (N_9718,N_9593,N_9536);
nand U9719 (N_9719,N_9483,N_9447);
nand U9720 (N_9720,N_9567,N_9402);
nor U9721 (N_9721,N_9508,N_9505);
and U9722 (N_9722,N_9412,N_9552);
nor U9723 (N_9723,N_9452,N_9526);
or U9724 (N_9724,N_9570,N_9405);
nor U9725 (N_9725,N_9408,N_9491);
nor U9726 (N_9726,N_9538,N_9517);
nor U9727 (N_9727,N_9556,N_9513);
and U9728 (N_9728,N_9568,N_9589);
and U9729 (N_9729,N_9571,N_9508);
nor U9730 (N_9730,N_9452,N_9484);
or U9731 (N_9731,N_9589,N_9515);
nand U9732 (N_9732,N_9419,N_9503);
nor U9733 (N_9733,N_9552,N_9487);
nor U9734 (N_9734,N_9486,N_9419);
xnor U9735 (N_9735,N_9597,N_9474);
or U9736 (N_9736,N_9422,N_9547);
or U9737 (N_9737,N_9451,N_9456);
or U9738 (N_9738,N_9538,N_9569);
or U9739 (N_9739,N_9454,N_9479);
and U9740 (N_9740,N_9553,N_9556);
and U9741 (N_9741,N_9561,N_9459);
and U9742 (N_9742,N_9496,N_9442);
and U9743 (N_9743,N_9581,N_9550);
and U9744 (N_9744,N_9400,N_9493);
nand U9745 (N_9745,N_9456,N_9462);
and U9746 (N_9746,N_9590,N_9529);
nand U9747 (N_9747,N_9556,N_9554);
xnor U9748 (N_9748,N_9582,N_9552);
or U9749 (N_9749,N_9460,N_9510);
nor U9750 (N_9750,N_9595,N_9493);
nor U9751 (N_9751,N_9458,N_9545);
nand U9752 (N_9752,N_9414,N_9506);
and U9753 (N_9753,N_9526,N_9552);
and U9754 (N_9754,N_9477,N_9551);
nor U9755 (N_9755,N_9546,N_9405);
or U9756 (N_9756,N_9526,N_9450);
or U9757 (N_9757,N_9490,N_9463);
or U9758 (N_9758,N_9516,N_9427);
xnor U9759 (N_9759,N_9550,N_9566);
and U9760 (N_9760,N_9535,N_9484);
xor U9761 (N_9761,N_9573,N_9579);
or U9762 (N_9762,N_9597,N_9463);
and U9763 (N_9763,N_9463,N_9549);
nor U9764 (N_9764,N_9504,N_9400);
nor U9765 (N_9765,N_9439,N_9530);
and U9766 (N_9766,N_9549,N_9542);
or U9767 (N_9767,N_9598,N_9453);
or U9768 (N_9768,N_9564,N_9581);
or U9769 (N_9769,N_9562,N_9521);
or U9770 (N_9770,N_9580,N_9472);
nand U9771 (N_9771,N_9584,N_9455);
and U9772 (N_9772,N_9573,N_9475);
nand U9773 (N_9773,N_9525,N_9438);
nor U9774 (N_9774,N_9515,N_9487);
nor U9775 (N_9775,N_9445,N_9584);
nand U9776 (N_9776,N_9453,N_9521);
nor U9777 (N_9777,N_9471,N_9437);
xnor U9778 (N_9778,N_9495,N_9426);
or U9779 (N_9779,N_9597,N_9418);
nor U9780 (N_9780,N_9463,N_9587);
or U9781 (N_9781,N_9510,N_9455);
or U9782 (N_9782,N_9432,N_9414);
xnor U9783 (N_9783,N_9560,N_9446);
xor U9784 (N_9784,N_9490,N_9473);
or U9785 (N_9785,N_9407,N_9554);
nor U9786 (N_9786,N_9413,N_9571);
nor U9787 (N_9787,N_9537,N_9529);
nand U9788 (N_9788,N_9568,N_9506);
xor U9789 (N_9789,N_9452,N_9553);
nand U9790 (N_9790,N_9541,N_9505);
nor U9791 (N_9791,N_9421,N_9550);
and U9792 (N_9792,N_9532,N_9480);
and U9793 (N_9793,N_9538,N_9593);
and U9794 (N_9794,N_9471,N_9485);
and U9795 (N_9795,N_9515,N_9406);
xor U9796 (N_9796,N_9491,N_9592);
or U9797 (N_9797,N_9519,N_9576);
nand U9798 (N_9798,N_9552,N_9459);
and U9799 (N_9799,N_9509,N_9577);
nand U9800 (N_9800,N_9793,N_9622);
or U9801 (N_9801,N_9672,N_9777);
nand U9802 (N_9802,N_9710,N_9664);
nor U9803 (N_9803,N_9612,N_9776);
or U9804 (N_9804,N_9707,N_9633);
nand U9805 (N_9805,N_9685,N_9603);
nor U9806 (N_9806,N_9607,N_9682);
or U9807 (N_9807,N_9683,N_9732);
or U9808 (N_9808,N_9613,N_9722);
nand U9809 (N_9809,N_9688,N_9698);
and U9810 (N_9810,N_9785,N_9624);
nand U9811 (N_9811,N_9733,N_9640);
or U9812 (N_9812,N_9704,N_9714);
nand U9813 (N_9813,N_9773,N_9711);
xor U9814 (N_9814,N_9638,N_9716);
nand U9815 (N_9815,N_9620,N_9792);
and U9816 (N_9816,N_9650,N_9771);
nand U9817 (N_9817,N_9621,N_9751);
nand U9818 (N_9818,N_9798,N_9794);
and U9819 (N_9819,N_9750,N_9634);
nor U9820 (N_9820,N_9632,N_9699);
nand U9821 (N_9821,N_9791,N_9696);
nor U9822 (N_9822,N_9646,N_9656);
or U9823 (N_9823,N_9759,N_9774);
and U9824 (N_9824,N_9743,N_9770);
or U9825 (N_9825,N_9605,N_9731);
nor U9826 (N_9826,N_9604,N_9687);
nand U9827 (N_9827,N_9693,N_9655);
or U9828 (N_9828,N_9667,N_9764);
nor U9829 (N_9829,N_9601,N_9691);
nand U9830 (N_9830,N_9659,N_9629);
and U9831 (N_9831,N_9709,N_9727);
and U9832 (N_9832,N_9639,N_9738);
nand U9833 (N_9833,N_9643,N_9670);
or U9834 (N_9834,N_9676,N_9679);
nor U9835 (N_9835,N_9627,N_9781);
or U9836 (N_9836,N_9675,N_9726);
xnor U9837 (N_9837,N_9662,N_9702);
and U9838 (N_9838,N_9649,N_9749);
and U9839 (N_9839,N_9723,N_9712);
xor U9840 (N_9840,N_9737,N_9626);
nand U9841 (N_9841,N_9706,N_9784);
nor U9842 (N_9842,N_9769,N_9747);
nor U9843 (N_9843,N_9684,N_9772);
or U9844 (N_9844,N_9775,N_9677);
nand U9845 (N_9845,N_9758,N_9782);
nor U9846 (N_9846,N_9680,N_9739);
and U9847 (N_9847,N_9705,N_9674);
xor U9848 (N_9848,N_9665,N_9615);
and U9849 (N_9849,N_9745,N_9761);
nor U9850 (N_9850,N_9763,N_9618);
nand U9851 (N_9851,N_9609,N_9729);
nand U9852 (N_9852,N_9623,N_9795);
nor U9853 (N_9853,N_9668,N_9600);
nand U9854 (N_9854,N_9602,N_9721);
or U9855 (N_9855,N_9637,N_9689);
nor U9856 (N_9856,N_9720,N_9779);
nor U9857 (N_9857,N_9760,N_9753);
nand U9858 (N_9858,N_9715,N_9631);
and U9859 (N_9859,N_9625,N_9799);
and U9860 (N_9860,N_9740,N_9628);
or U9861 (N_9861,N_9756,N_9783);
nor U9862 (N_9862,N_9766,N_9614);
and U9863 (N_9863,N_9703,N_9719);
and U9864 (N_9864,N_9744,N_9741);
or U9865 (N_9865,N_9630,N_9717);
or U9866 (N_9866,N_9635,N_9641);
nand U9867 (N_9867,N_9658,N_9697);
and U9868 (N_9868,N_9786,N_9701);
nand U9869 (N_9869,N_9736,N_9700);
and U9870 (N_9870,N_9654,N_9718);
and U9871 (N_9871,N_9765,N_9694);
or U9872 (N_9872,N_9644,N_9671);
and U9873 (N_9873,N_9748,N_9610);
and U9874 (N_9874,N_9796,N_9619);
nand U9875 (N_9875,N_9663,N_9606);
and U9876 (N_9876,N_9787,N_9746);
or U9877 (N_9877,N_9754,N_9728);
nand U9878 (N_9878,N_9725,N_9616);
nand U9879 (N_9879,N_9788,N_9780);
or U9880 (N_9880,N_9617,N_9657);
and U9881 (N_9881,N_9742,N_9611);
and U9882 (N_9882,N_9647,N_9790);
nand U9883 (N_9883,N_9636,N_9648);
or U9884 (N_9884,N_9724,N_9695);
or U9885 (N_9885,N_9669,N_9767);
and U9886 (N_9886,N_9692,N_9681);
and U9887 (N_9887,N_9673,N_9757);
nand U9888 (N_9888,N_9678,N_9652);
xnor U9889 (N_9889,N_9651,N_9645);
or U9890 (N_9890,N_9734,N_9660);
nand U9891 (N_9891,N_9713,N_9642);
nand U9892 (N_9892,N_9778,N_9686);
nand U9893 (N_9893,N_9768,N_9608);
or U9894 (N_9894,N_9797,N_9752);
nor U9895 (N_9895,N_9730,N_9661);
nand U9896 (N_9896,N_9789,N_9690);
or U9897 (N_9897,N_9735,N_9762);
and U9898 (N_9898,N_9666,N_9708);
nand U9899 (N_9899,N_9653,N_9755);
nor U9900 (N_9900,N_9660,N_9718);
nor U9901 (N_9901,N_9756,N_9712);
nand U9902 (N_9902,N_9634,N_9767);
nand U9903 (N_9903,N_9622,N_9720);
or U9904 (N_9904,N_9665,N_9625);
and U9905 (N_9905,N_9626,N_9681);
or U9906 (N_9906,N_9789,N_9627);
and U9907 (N_9907,N_9644,N_9615);
and U9908 (N_9908,N_9638,N_9618);
or U9909 (N_9909,N_9600,N_9741);
nor U9910 (N_9910,N_9757,N_9754);
or U9911 (N_9911,N_9612,N_9673);
nand U9912 (N_9912,N_9717,N_9646);
or U9913 (N_9913,N_9787,N_9607);
or U9914 (N_9914,N_9607,N_9654);
or U9915 (N_9915,N_9625,N_9635);
and U9916 (N_9916,N_9786,N_9686);
and U9917 (N_9917,N_9613,N_9742);
nand U9918 (N_9918,N_9786,N_9634);
nand U9919 (N_9919,N_9665,N_9725);
or U9920 (N_9920,N_9650,N_9609);
or U9921 (N_9921,N_9727,N_9615);
or U9922 (N_9922,N_9650,N_9789);
or U9923 (N_9923,N_9717,N_9677);
and U9924 (N_9924,N_9721,N_9775);
nand U9925 (N_9925,N_9649,N_9760);
nand U9926 (N_9926,N_9793,N_9655);
nand U9927 (N_9927,N_9798,N_9621);
nand U9928 (N_9928,N_9779,N_9663);
and U9929 (N_9929,N_9767,N_9602);
nand U9930 (N_9930,N_9619,N_9683);
or U9931 (N_9931,N_9663,N_9785);
and U9932 (N_9932,N_9755,N_9742);
nand U9933 (N_9933,N_9648,N_9754);
xnor U9934 (N_9934,N_9625,N_9604);
and U9935 (N_9935,N_9709,N_9664);
and U9936 (N_9936,N_9714,N_9614);
nand U9937 (N_9937,N_9791,N_9728);
nand U9938 (N_9938,N_9774,N_9616);
nor U9939 (N_9939,N_9797,N_9685);
xor U9940 (N_9940,N_9727,N_9744);
nor U9941 (N_9941,N_9787,N_9638);
nor U9942 (N_9942,N_9727,N_9607);
or U9943 (N_9943,N_9735,N_9767);
nor U9944 (N_9944,N_9635,N_9664);
nor U9945 (N_9945,N_9613,N_9689);
and U9946 (N_9946,N_9728,N_9610);
nor U9947 (N_9947,N_9794,N_9747);
xor U9948 (N_9948,N_9639,N_9632);
xnor U9949 (N_9949,N_9624,N_9744);
nor U9950 (N_9950,N_9709,N_9683);
and U9951 (N_9951,N_9716,N_9700);
xor U9952 (N_9952,N_9700,N_9649);
nand U9953 (N_9953,N_9762,N_9695);
xnor U9954 (N_9954,N_9644,N_9647);
nor U9955 (N_9955,N_9660,N_9618);
nor U9956 (N_9956,N_9745,N_9784);
and U9957 (N_9957,N_9623,N_9668);
nand U9958 (N_9958,N_9696,N_9734);
xnor U9959 (N_9959,N_9710,N_9737);
and U9960 (N_9960,N_9708,N_9704);
xor U9961 (N_9961,N_9704,N_9735);
and U9962 (N_9962,N_9789,N_9733);
and U9963 (N_9963,N_9734,N_9742);
and U9964 (N_9964,N_9763,N_9652);
nand U9965 (N_9965,N_9603,N_9697);
and U9966 (N_9966,N_9785,N_9672);
nand U9967 (N_9967,N_9658,N_9729);
or U9968 (N_9968,N_9625,N_9739);
nor U9969 (N_9969,N_9602,N_9664);
and U9970 (N_9970,N_9744,N_9792);
or U9971 (N_9971,N_9611,N_9713);
or U9972 (N_9972,N_9620,N_9671);
and U9973 (N_9973,N_9642,N_9603);
nor U9974 (N_9974,N_9642,N_9636);
or U9975 (N_9975,N_9763,N_9663);
or U9976 (N_9976,N_9658,N_9667);
or U9977 (N_9977,N_9726,N_9687);
or U9978 (N_9978,N_9631,N_9694);
or U9979 (N_9979,N_9690,N_9729);
or U9980 (N_9980,N_9613,N_9705);
or U9981 (N_9981,N_9612,N_9605);
or U9982 (N_9982,N_9687,N_9651);
and U9983 (N_9983,N_9643,N_9676);
and U9984 (N_9984,N_9751,N_9786);
and U9985 (N_9985,N_9704,N_9737);
nor U9986 (N_9986,N_9721,N_9733);
nor U9987 (N_9987,N_9727,N_9799);
or U9988 (N_9988,N_9758,N_9761);
or U9989 (N_9989,N_9750,N_9796);
nor U9990 (N_9990,N_9740,N_9786);
nor U9991 (N_9991,N_9651,N_9780);
and U9992 (N_9992,N_9671,N_9769);
and U9993 (N_9993,N_9654,N_9739);
nor U9994 (N_9994,N_9699,N_9760);
xor U9995 (N_9995,N_9789,N_9638);
and U9996 (N_9996,N_9675,N_9788);
or U9997 (N_9997,N_9666,N_9728);
nand U9998 (N_9998,N_9742,N_9664);
nor U9999 (N_9999,N_9615,N_9681);
nor U10000 (N_10000,N_9809,N_9838);
and U10001 (N_10001,N_9991,N_9942);
or U10002 (N_10002,N_9817,N_9971);
nand U10003 (N_10003,N_9891,N_9924);
or U10004 (N_10004,N_9970,N_9888);
nor U10005 (N_10005,N_9807,N_9922);
and U10006 (N_10006,N_9901,N_9806);
nor U10007 (N_10007,N_9816,N_9859);
xnor U10008 (N_10008,N_9897,N_9883);
xor U10009 (N_10009,N_9907,N_9915);
and U10010 (N_10010,N_9962,N_9905);
or U10011 (N_10011,N_9958,N_9840);
nor U10012 (N_10012,N_9974,N_9882);
and U10013 (N_10013,N_9821,N_9870);
nor U10014 (N_10014,N_9815,N_9895);
xor U10015 (N_10015,N_9823,N_9914);
nor U10016 (N_10016,N_9873,N_9956);
and U10017 (N_10017,N_9878,N_9802);
or U10018 (N_10018,N_9953,N_9803);
xnor U10019 (N_10019,N_9844,N_9919);
or U10020 (N_10020,N_9811,N_9909);
and U10021 (N_10021,N_9975,N_9952);
and U10022 (N_10022,N_9865,N_9862);
nor U10023 (N_10023,N_9973,N_9810);
nand U10024 (N_10024,N_9886,N_9856);
nand U10025 (N_10025,N_9997,N_9880);
or U10026 (N_10026,N_9985,N_9853);
nor U10027 (N_10027,N_9904,N_9872);
and U10028 (N_10028,N_9874,N_9800);
nand U10029 (N_10029,N_9913,N_9935);
and U10030 (N_10030,N_9871,N_9881);
or U10031 (N_10031,N_9827,N_9959);
and U10032 (N_10032,N_9968,N_9887);
nand U10033 (N_10033,N_9834,N_9890);
nand U10034 (N_10034,N_9825,N_9930);
nor U10035 (N_10035,N_9885,N_9858);
or U10036 (N_10036,N_9948,N_9855);
xor U10037 (N_10037,N_9812,N_9999);
or U10038 (N_10038,N_9993,N_9826);
nor U10039 (N_10039,N_9900,N_9955);
and U10040 (N_10040,N_9896,N_9884);
or U10041 (N_10041,N_9851,N_9943);
xnor U10042 (N_10042,N_9839,N_9967);
nand U10043 (N_10043,N_9928,N_9921);
nand U10044 (N_10044,N_9863,N_9845);
nand U10045 (N_10045,N_9992,N_9960);
nand U10046 (N_10046,N_9941,N_9950);
nor U10047 (N_10047,N_9964,N_9898);
and U10048 (N_10048,N_9932,N_9824);
and U10049 (N_10049,N_9831,N_9920);
xnor U10050 (N_10050,N_9814,N_9938);
nand U10051 (N_10051,N_9850,N_9829);
nor U10052 (N_10052,N_9848,N_9830);
nand U10053 (N_10053,N_9983,N_9899);
xnor U10054 (N_10054,N_9804,N_9929);
nor U10055 (N_10055,N_9987,N_9923);
nor U10056 (N_10056,N_9966,N_9903);
nand U10057 (N_10057,N_9828,N_9989);
or U10058 (N_10058,N_9910,N_9918);
and U10059 (N_10059,N_9980,N_9965);
and U10060 (N_10060,N_9902,N_9925);
or U10061 (N_10061,N_9820,N_9944);
nand U10062 (N_10062,N_9990,N_9951);
and U10063 (N_10063,N_9861,N_9996);
nand U10064 (N_10064,N_9911,N_9933);
and U10065 (N_10065,N_9946,N_9867);
nand U10066 (N_10066,N_9852,N_9988);
nand U10067 (N_10067,N_9846,N_9876);
and U10068 (N_10068,N_9912,N_9866);
nor U10069 (N_10069,N_9860,N_9864);
and U10070 (N_10070,N_9949,N_9875);
nand U10071 (N_10071,N_9995,N_9813);
xor U10072 (N_10072,N_9893,N_9843);
or U10073 (N_10073,N_9857,N_9934);
and U10074 (N_10074,N_9917,N_9981);
nor U10075 (N_10075,N_9847,N_9936);
nor U10076 (N_10076,N_9889,N_9849);
nand U10077 (N_10077,N_9836,N_9908);
nor U10078 (N_10078,N_9805,N_9894);
or U10079 (N_10079,N_9931,N_9854);
or U10080 (N_10080,N_9998,N_9940);
nand U10081 (N_10081,N_9927,N_9822);
nor U10082 (N_10082,N_9947,N_9833);
and U10083 (N_10083,N_9954,N_9961);
or U10084 (N_10084,N_9978,N_9842);
and U10085 (N_10085,N_9986,N_9979);
or U10086 (N_10086,N_9945,N_9984);
or U10087 (N_10087,N_9906,N_9994);
nor U10088 (N_10088,N_9869,N_9835);
and U10089 (N_10089,N_9868,N_9801);
nand U10090 (N_10090,N_9808,N_9916);
nand U10091 (N_10091,N_9977,N_9832);
nor U10092 (N_10092,N_9972,N_9818);
nor U10093 (N_10093,N_9937,N_9976);
nor U10094 (N_10094,N_9819,N_9982);
nor U10095 (N_10095,N_9837,N_9963);
or U10096 (N_10096,N_9841,N_9957);
or U10097 (N_10097,N_9926,N_9877);
nor U10098 (N_10098,N_9969,N_9892);
or U10099 (N_10099,N_9939,N_9879);
xor U10100 (N_10100,N_9862,N_9892);
and U10101 (N_10101,N_9855,N_9967);
nor U10102 (N_10102,N_9857,N_9961);
nand U10103 (N_10103,N_9973,N_9848);
or U10104 (N_10104,N_9998,N_9884);
nand U10105 (N_10105,N_9877,N_9814);
nor U10106 (N_10106,N_9804,N_9950);
and U10107 (N_10107,N_9998,N_9881);
and U10108 (N_10108,N_9881,N_9829);
or U10109 (N_10109,N_9842,N_9888);
or U10110 (N_10110,N_9853,N_9849);
xor U10111 (N_10111,N_9837,N_9885);
and U10112 (N_10112,N_9800,N_9985);
nor U10113 (N_10113,N_9913,N_9974);
xor U10114 (N_10114,N_9910,N_9885);
or U10115 (N_10115,N_9928,N_9949);
and U10116 (N_10116,N_9926,N_9893);
xnor U10117 (N_10117,N_9801,N_9952);
or U10118 (N_10118,N_9900,N_9947);
or U10119 (N_10119,N_9869,N_9830);
xor U10120 (N_10120,N_9804,N_9948);
nand U10121 (N_10121,N_9920,N_9812);
nand U10122 (N_10122,N_9949,N_9948);
and U10123 (N_10123,N_9944,N_9922);
nor U10124 (N_10124,N_9879,N_9860);
xor U10125 (N_10125,N_9939,N_9828);
and U10126 (N_10126,N_9955,N_9880);
nor U10127 (N_10127,N_9918,N_9922);
nand U10128 (N_10128,N_9930,N_9931);
nor U10129 (N_10129,N_9825,N_9990);
xor U10130 (N_10130,N_9840,N_9896);
or U10131 (N_10131,N_9829,N_9952);
and U10132 (N_10132,N_9898,N_9844);
and U10133 (N_10133,N_9955,N_9927);
nand U10134 (N_10134,N_9814,N_9843);
nand U10135 (N_10135,N_9918,N_9907);
nor U10136 (N_10136,N_9933,N_9903);
or U10137 (N_10137,N_9882,N_9962);
nor U10138 (N_10138,N_9939,N_9898);
nor U10139 (N_10139,N_9900,N_9953);
xor U10140 (N_10140,N_9867,N_9840);
nor U10141 (N_10141,N_9944,N_9991);
or U10142 (N_10142,N_9870,N_9936);
and U10143 (N_10143,N_9823,N_9998);
nor U10144 (N_10144,N_9876,N_9911);
or U10145 (N_10145,N_9968,N_9857);
and U10146 (N_10146,N_9957,N_9930);
nor U10147 (N_10147,N_9991,N_9964);
nor U10148 (N_10148,N_9872,N_9974);
or U10149 (N_10149,N_9861,N_9898);
and U10150 (N_10150,N_9872,N_9973);
and U10151 (N_10151,N_9878,N_9965);
nor U10152 (N_10152,N_9819,N_9862);
nor U10153 (N_10153,N_9928,N_9847);
and U10154 (N_10154,N_9986,N_9804);
nand U10155 (N_10155,N_9932,N_9803);
xor U10156 (N_10156,N_9947,N_9804);
nor U10157 (N_10157,N_9963,N_9980);
nor U10158 (N_10158,N_9880,N_9992);
xnor U10159 (N_10159,N_9828,N_9927);
and U10160 (N_10160,N_9957,N_9824);
nor U10161 (N_10161,N_9946,N_9829);
or U10162 (N_10162,N_9806,N_9988);
nand U10163 (N_10163,N_9891,N_9969);
nand U10164 (N_10164,N_9858,N_9867);
xor U10165 (N_10165,N_9979,N_9812);
and U10166 (N_10166,N_9907,N_9948);
nor U10167 (N_10167,N_9953,N_9835);
nand U10168 (N_10168,N_9981,N_9994);
and U10169 (N_10169,N_9953,N_9917);
nand U10170 (N_10170,N_9828,N_9879);
and U10171 (N_10171,N_9871,N_9969);
or U10172 (N_10172,N_9988,N_9860);
xnor U10173 (N_10173,N_9950,N_9898);
nor U10174 (N_10174,N_9938,N_9816);
and U10175 (N_10175,N_9977,N_9902);
nand U10176 (N_10176,N_9907,N_9851);
nor U10177 (N_10177,N_9951,N_9868);
nand U10178 (N_10178,N_9938,N_9865);
xor U10179 (N_10179,N_9953,N_9887);
nand U10180 (N_10180,N_9963,N_9800);
or U10181 (N_10181,N_9823,N_9927);
nand U10182 (N_10182,N_9875,N_9915);
nor U10183 (N_10183,N_9909,N_9839);
and U10184 (N_10184,N_9929,N_9925);
nor U10185 (N_10185,N_9982,N_9812);
and U10186 (N_10186,N_9840,N_9861);
nor U10187 (N_10187,N_9879,N_9914);
nor U10188 (N_10188,N_9959,N_9803);
or U10189 (N_10189,N_9939,N_9835);
nand U10190 (N_10190,N_9925,N_9815);
or U10191 (N_10191,N_9815,N_9941);
nor U10192 (N_10192,N_9982,N_9863);
or U10193 (N_10193,N_9917,N_9857);
nand U10194 (N_10194,N_9891,N_9850);
nor U10195 (N_10195,N_9822,N_9881);
and U10196 (N_10196,N_9972,N_9821);
nand U10197 (N_10197,N_9888,N_9872);
xnor U10198 (N_10198,N_9821,N_9867);
xnor U10199 (N_10199,N_9824,N_9833);
or U10200 (N_10200,N_10060,N_10116);
nor U10201 (N_10201,N_10190,N_10183);
xnor U10202 (N_10202,N_10155,N_10140);
or U10203 (N_10203,N_10144,N_10036);
nor U10204 (N_10204,N_10139,N_10147);
nand U10205 (N_10205,N_10187,N_10051);
nor U10206 (N_10206,N_10006,N_10143);
or U10207 (N_10207,N_10089,N_10101);
and U10208 (N_10208,N_10088,N_10065);
and U10209 (N_10209,N_10160,N_10017);
and U10210 (N_10210,N_10098,N_10104);
and U10211 (N_10211,N_10199,N_10039);
xor U10212 (N_10212,N_10063,N_10015);
xnor U10213 (N_10213,N_10166,N_10177);
and U10214 (N_10214,N_10188,N_10020);
nand U10215 (N_10215,N_10007,N_10107);
nand U10216 (N_10216,N_10138,N_10081);
nand U10217 (N_10217,N_10168,N_10167);
nand U10218 (N_10218,N_10161,N_10057);
or U10219 (N_10219,N_10103,N_10146);
nor U10220 (N_10220,N_10040,N_10151);
nor U10221 (N_10221,N_10096,N_10001);
nor U10222 (N_10222,N_10087,N_10179);
or U10223 (N_10223,N_10084,N_10186);
nand U10224 (N_10224,N_10148,N_10111);
or U10225 (N_10225,N_10061,N_10184);
or U10226 (N_10226,N_10134,N_10198);
nand U10227 (N_10227,N_10128,N_10112);
nand U10228 (N_10228,N_10086,N_10054);
nor U10229 (N_10229,N_10085,N_10047);
or U10230 (N_10230,N_10176,N_10008);
nand U10231 (N_10231,N_10091,N_10082);
or U10232 (N_10232,N_10123,N_10074);
nor U10233 (N_10233,N_10126,N_10153);
nor U10234 (N_10234,N_10165,N_10191);
nor U10235 (N_10235,N_10083,N_10178);
or U10236 (N_10236,N_10108,N_10070);
and U10237 (N_10237,N_10130,N_10080);
nand U10238 (N_10238,N_10012,N_10196);
nor U10239 (N_10239,N_10005,N_10052);
and U10240 (N_10240,N_10124,N_10050);
or U10241 (N_10241,N_10189,N_10113);
and U10242 (N_10242,N_10000,N_10014);
or U10243 (N_10243,N_10182,N_10023);
nor U10244 (N_10244,N_10021,N_10055);
and U10245 (N_10245,N_10154,N_10046);
and U10246 (N_10246,N_10171,N_10169);
nor U10247 (N_10247,N_10044,N_10035);
nor U10248 (N_10248,N_10117,N_10135);
and U10249 (N_10249,N_10159,N_10094);
xor U10250 (N_10250,N_10068,N_10025);
and U10251 (N_10251,N_10129,N_10100);
xor U10252 (N_10252,N_10106,N_10033);
nand U10253 (N_10253,N_10152,N_10149);
and U10254 (N_10254,N_10192,N_10018);
nand U10255 (N_10255,N_10019,N_10120);
or U10256 (N_10256,N_10145,N_10181);
nor U10257 (N_10257,N_10141,N_10026);
nor U10258 (N_10258,N_10099,N_10058);
or U10259 (N_10259,N_10136,N_10158);
xnor U10260 (N_10260,N_10133,N_10121);
nor U10261 (N_10261,N_10062,N_10180);
nand U10262 (N_10262,N_10027,N_10043);
and U10263 (N_10263,N_10024,N_10110);
nor U10264 (N_10264,N_10131,N_10079);
nand U10265 (N_10265,N_10185,N_10078);
xor U10266 (N_10266,N_10009,N_10115);
or U10267 (N_10267,N_10105,N_10045);
and U10268 (N_10268,N_10175,N_10072);
or U10269 (N_10269,N_10071,N_10157);
or U10270 (N_10270,N_10150,N_10197);
nand U10271 (N_10271,N_10193,N_10194);
xnor U10272 (N_10272,N_10059,N_10142);
or U10273 (N_10273,N_10114,N_10002);
or U10274 (N_10274,N_10031,N_10064);
or U10275 (N_10275,N_10042,N_10092);
or U10276 (N_10276,N_10003,N_10156);
nand U10277 (N_10277,N_10075,N_10016);
xnor U10278 (N_10278,N_10049,N_10125);
nand U10279 (N_10279,N_10034,N_10048);
or U10280 (N_10280,N_10119,N_10022);
or U10281 (N_10281,N_10132,N_10073);
xnor U10282 (N_10282,N_10077,N_10004);
or U10283 (N_10283,N_10037,N_10164);
nor U10284 (N_10284,N_10053,N_10056);
nor U10285 (N_10285,N_10029,N_10067);
or U10286 (N_10286,N_10013,N_10032);
or U10287 (N_10287,N_10011,N_10069);
nor U10288 (N_10288,N_10163,N_10066);
or U10289 (N_10289,N_10162,N_10102);
or U10290 (N_10290,N_10174,N_10195);
nor U10291 (N_10291,N_10093,N_10030);
or U10292 (N_10292,N_10173,N_10170);
or U10293 (N_10293,N_10010,N_10172);
nand U10294 (N_10294,N_10041,N_10109);
nand U10295 (N_10295,N_10137,N_10118);
xnor U10296 (N_10296,N_10097,N_10038);
nand U10297 (N_10297,N_10076,N_10095);
or U10298 (N_10298,N_10122,N_10127);
nor U10299 (N_10299,N_10028,N_10090);
and U10300 (N_10300,N_10084,N_10027);
nand U10301 (N_10301,N_10056,N_10076);
or U10302 (N_10302,N_10084,N_10139);
xor U10303 (N_10303,N_10184,N_10093);
or U10304 (N_10304,N_10072,N_10036);
xor U10305 (N_10305,N_10114,N_10031);
nor U10306 (N_10306,N_10162,N_10130);
and U10307 (N_10307,N_10094,N_10057);
and U10308 (N_10308,N_10124,N_10115);
nor U10309 (N_10309,N_10024,N_10050);
and U10310 (N_10310,N_10028,N_10072);
or U10311 (N_10311,N_10131,N_10154);
nand U10312 (N_10312,N_10182,N_10139);
and U10313 (N_10313,N_10180,N_10002);
and U10314 (N_10314,N_10048,N_10035);
or U10315 (N_10315,N_10044,N_10144);
and U10316 (N_10316,N_10039,N_10136);
or U10317 (N_10317,N_10100,N_10041);
and U10318 (N_10318,N_10099,N_10032);
nor U10319 (N_10319,N_10191,N_10105);
nor U10320 (N_10320,N_10134,N_10074);
and U10321 (N_10321,N_10045,N_10198);
and U10322 (N_10322,N_10019,N_10030);
or U10323 (N_10323,N_10040,N_10033);
nor U10324 (N_10324,N_10185,N_10178);
and U10325 (N_10325,N_10019,N_10076);
and U10326 (N_10326,N_10073,N_10142);
nand U10327 (N_10327,N_10187,N_10071);
nor U10328 (N_10328,N_10027,N_10015);
and U10329 (N_10329,N_10031,N_10066);
nand U10330 (N_10330,N_10141,N_10128);
or U10331 (N_10331,N_10058,N_10007);
or U10332 (N_10332,N_10105,N_10035);
or U10333 (N_10333,N_10063,N_10089);
nand U10334 (N_10334,N_10019,N_10026);
or U10335 (N_10335,N_10013,N_10161);
nand U10336 (N_10336,N_10046,N_10091);
and U10337 (N_10337,N_10177,N_10122);
or U10338 (N_10338,N_10037,N_10090);
and U10339 (N_10339,N_10166,N_10098);
and U10340 (N_10340,N_10125,N_10129);
nor U10341 (N_10341,N_10062,N_10044);
xor U10342 (N_10342,N_10119,N_10057);
nand U10343 (N_10343,N_10113,N_10032);
nand U10344 (N_10344,N_10147,N_10163);
and U10345 (N_10345,N_10131,N_10095);
or U10346 (N_10346,N_10181,N_10046);
and U10347 (N_10347,N_10163,N_10167);
nor U10348 (N_10348,N_10002,N_10018);
nand U10349 (N_10349,N_10003,N_10177);
and U10350 (N_10350,N_10162,N_10022);
and U10351 (N_10351,N_10021,N_10006);
and U10352 (N_10352,N_10072,N_10193);
nand U10353 (N_10353,N_10015,N_10139);
or U10354 (N_10354,N_10146,N_10118);
or U10355 (N_10355,N_10079,N_10191);
nor U10356 (N_10356,N_10127,N_10148);
and U10357 (N_10357,N_10169,N_10097);
and U10358 (N_10358,N_10066,N_10072);
and U10359 (N_10359,N_10055,N_10069);
nor U10360 (N_10360,N_10019,N_10189);
nor U10361 (N_10361,N_10046,N_10198);
nor U10362 (N_10362,N_10050,N_10059);
nand U10363 (N_10363,N_10169,N_10004);
nand U10364 (N_10364,N_10063,N_10192);
nor U10365 (N_10365,N_10087,N_10052);
or U10366 (N_10366,N_10010,N_10055);
and U10367 (N_10367,N_10030,N_10076);
nor U10368 (N_10368,N_10181,N_10131);
nand U10369 (N_10369,N_10060,N_10008);
xor U10370 (N_10370,N_10116,N_10115);
or U10371 (N_10371,N_10116,N_10187);
and U10372 (N_10372,N_10001,N_10102);
xor U10373 (N_10373,N_10009,N_10143);
nor U10374 (N_10374,N_10019,N_10046);
nand U10375 (N_10375,N_10042,N_10045);
and U10376 (N_10376,N_10150,N_10088);
nor U10377 (N_10377,N_10183,N_10025);
and U10378 (N_10378,N_10015,N_10189);
nand U10379 (N_10379,N_10085,N_10174);
and U10380 (N_10380,N_10071,N_10186);
nor U10381 (N_10381,N_10190,N_10153);
or U10382 (N_10382,N_10043,N_10151);
or U10383 (N_10383,N_10130,N_10116);
xor U10384 (N_10384,N_10121,N_10103);
or U10385 (N_10385,N_10166,N_10073);
nand U10386 (N_10386,N_10062,N_10164);
or U10387 (N_10387,N_10082,N_10040);
nand U10388 (N_10388,N_10004,N_10181);
nor U10389 (N_10389,N_10188,N_10125);
nand U10390 (N_10390,N_10134,N_10106);
and U10391 (N_10391,N_10143,N_10116);
nor U10392 (N_10392,N_10006,N_10076);
nand U10393 (N_10393,N_10167,N_10118);
and U10394 (N_10394,N_10115,N_10023);
and U10395 (N_10395,N_10022,N_10171);
nand U10396 (N_10396,N_10086,N_10081);
and U10397 (N_10397,N_10152,N_10090);
or U10398 (N_10398,N_10033,N_10005);
nand U10399 (N_10399,N_10100,N_10127);
nand U10400 (N_10400,N_10362,N_10281);
and U10401 (N_10401,N_10257,N_10284);
and U10402 (N_10402,N_10241,N_10220);
and U10403 (N_10403,N_10256,N_10309);
nor U10404 (N_10404,N_10370,N_10270);
and U10405 (N_10405,N_10260,N_10391);
or U10406 (N_10406,N_10317,N_10338);
nor U10407 (N_10407,N_10264,N_10352);
or U10408 (N_10408,N_10226,N_10332);
and U10409 (N_10409,N_10319,N_10335);
or U10410 (N_10410,N_10393,N_10327);
nand U10411 (N_10411,N_10214,N_10377);
nor U10412 (N_10412,N_10245,N_10240);
nor U10413 (N_10413,N_10367,N_10231);
and U10414 (N_10414,N_10348,N_10325);
or U10415 (N_10415,N_10273,N_10349);
nand U10416 (N_10416,N_10254,N_10301);
nand U10417 (N_10417,N_10251,N_10266);
and U10418 (N_10418,N_10380,N_10218);
nor U10419 (N_10419,N_10372,N_10295);
xor U10420 (N_10420,N_10347,N_10246);
nor U10421 (N_10421,N_10308,N_10290);
or U10422 (N_10422,N_10376,N_10344);
or U10423 (N_10423,N_10207,N_10351);
xor U10424 (N_10424,N_10313,N_10353);
or U10425 (N_10425,N_10209,N_10250);
nor U10426 (N_10426,N_10244,N_10329);
nand U10427 (N_10427,N_10236,N_10314);
and U10428 (N_10428,N_10228,N_10343);
xnor U10429 (N_10429,N_10396,N_10390);
nor U10430 (N_10430,N_10263,N_10326);
and U10431 (N_10431,N_10235,N_10334);
or U10432 (N_10432,N_10224,N_10269);
and U10433 (N_10433,N_10365,N_10321);
nand U10434 (N_10434,N_10356,N_10294);
nor U10435 (N_10435,N_10300,N_10275);
nor U10436 (N_10436,N_10350,N_10303);
or U10437 (N_10437,N_10296,N_10346);
nor U10438 (N_10438,N_10213,N_10259);
nand U10439 (N_10439,N_10238,N_10305);
nand U10440 (N_10440,N_10312,N_10201);
nand U10441 (N_10441,N_10291,N_10381);
xor U10442 (N_10442,N_10359,N_10292);
or U10443 (N_10443,N_10252,N_10271);
xor U10444 (N_10444,N_10331,N_10375);
nand U10445 (N_10445,N_10366,N_10200);
and U10446 (N_10446,N_10210,N_10399);
nor U10447 (N_10447,N_10223,N_10341);
nand U10448 (N_10448,N_10289,N_10274);
nand U10449 (N_10449,N_10222,N_10398);
nand U10450 (N_10450,N_10282,N_10297);
nand U10451 (N_10451,N_10387,N_10310);
nor U10452 (N_10452,N_10371,N_10330);
and U10453 (N_10453,N_10299,N_10225);
and U10454 (N_10454,N_10361,N_10287);
nand U10455 (N_10455,N_10204,N_10219);
nor U10456 (N_10456,N_10262,N_10358);
xor U10457 (N_10457,N_10316,N_10221);
or U10458 (N_10458,N_10357,N_10395);
nor U10459 (N_10459,N_10217,N_10234);
and U10460 (N_10460,N_10258,N_10386);
and U10461 (N_10461,N_10208,N_10267);
nor U10462 (N_10462,N_10337,N_10322);
and U10463 (N_10463,N_10247,N_10354);
and U10464 (N_10464,N_10339,N_10379);
or U10465 (N_10465,N_10277,N_10323);
and U10466 (N_10466,N_10206,N_10383);
and U10467 (N_10467,N_10374,N_10268);
or U10468 (N_10468,N_10363,N_10232);
or U10469 (N_10469,N_10388,N_10285);
nand U10470 (N_10470,N_10394,N_10255);
nor U10471 (N_10471,N_10288,N_10205);
or U10472 (N_10472,N_10318,N_10243);
and U10473 (N_10473,N_10272,N_10239);
or U10474 (N_10474,N_10306,N_10382);
or U10475 (N_10475,N_10283,N_10265);
nand U10476 (N_10476,N_10384,N_10307);
nand U10477 (N_10477,N_10360,N_10355);
and U10478 (N_10478,N_10324,N_10242);
nor U10479 (N_10479,N_10342,N_10397);
nor U10480 (N_10480,N_10216,N_10389);
and U10481 (N_10481,N_10211,N_10237);
nor U10482 (N_10482,N_10280,N_10278);
nor U10483 (N_10483,N_10202,N_10315);
nand U10484 (N_10484,N_10212,N_10328);
and U10485 (N_10485,N_10233,N_10261);
nand U10486 (N_10486,N_10279,N_10340);
or U10487 (N_10487,N_10333,N_10248);
or U10488 (N_10488,N_10368,N_10203);
xnor U10489 (N_10489,N_10276,N_10227);
or U10490 (N_10490,N_10320,N_10378);
nor U10491 (N_10491,N_10229,N_10230);
nand U10492 (N_10492,N_10311,N_10298);
xor U10493 (N_10493,N_10304,N_10336);
xnor U10494 (N_10494,N_10345,N_10215);
or U10495 (N_10495,N_10385,N_10373);
xnor U10496 (N_10496,N_10302,N_10369);
nor U10497 (N_10497,N_10364,N_10293);
nand U10498 (N_10498,N_10286,N_10392);
and U10499 (N_10499,N_10253,N_10249);
nor U10500 (N_10500,N_10322,N_10245);
or U10501 (N_10501,N_10275,N_10393);
nor U10502 (N_10502,N_10254,N_10208);
and U10503 (N_10503,N_10249,N_10332);
nand U10504 (N_10504,N_10247,N_10321);
and U10505 (N_10505,N_10366,N_10343);
or U10506 (N_10506,N_10292,N_10274);
or U10507 (N_10507,N_10227,N_10349);
and U10508 (N_10508,N_10250,N_10296);
nand U10509 (N_10509,N_10202,N_10234);
or U10510 (N_10510,N_10338,N_10243);
or U10511 (N_10511,N_10345,N_10296);
nor U10512 (N_10512,N_10376,N_10238);
nand U10513 (N_10513,N_10262,N_10345);
or U10514 (N_10514,N_10263,N_10257);
nand U10515 (N_10515,N_10246,N_10227);
xor U10516 (N_10516,N_10228,N_10201);
and U10517 (N_10517,N_10273,N_10294);
nor U10518 (N_10518,N_10249,N_10243);
or U10519 (N_10519,N_10392,N_10381);
nand U10520 (N_10520,N_10370,N_10201);
nor U10521 (N_10521,N_10218,N_10394);
and U10522 (N_10522,N_10309,N_10221);
and U10523 (N_10523,N_10356,N_10381);
nand U10524 (N_10524,N_10218,N_10229);
nand U10525 (N_10525,N_10227,N_10264);
nand U10526 (N_10526,N_10360,N_10260);
nor U10527 (N_10527,N_10261,N_10310);
nor U10528 (N_10528,N_10208,N_10253);
or U10529 (N_10529,N_10397,N_10364);
and U10530 (N_10530,N_10220,N_10316);
nand U10531 (N_10531,N_10263,N_10237);
xnor U10532 (N_10532,N_10398,N_10213);
or U10533 (N_10533,N_10239,N_10303);
nor U10534 (N_10534,N_10355,N_10245);
and U10535 (N_10535,N_10336,N_10291);
and U10536 (N_10536,N_10397,N_10247);
xor U10537 (N_10537,N_10316,N_10302);
or U10538 (N_10538,N_10327,N_10275);
xor U10539 (N_10539,N_10321,N_10209);
xor U10540 (N_10540,N_10332,N_10306);
or U10541 (N_10541,N_10345,N_10346);
and U10542 (N_10542,N_10370,N_10379);
nand U10543 (N_10543,N_10256,N_10303);
and U10544 (N_10544,N_10374,N_10309);
xor U10545 (N_10545,N_10336,N_10361);
xor U10546 (N_10546,N_10381,N_10301);
nor U10547 (N_10547,N_10328,N_10216);
and U10548 (N_10548,N_10383,N_10399);
nor U10549 (N_10549,N_10338,N_10354);
nor U10550 (N_10550,N_10279,N_10253);
nor U10551 (N_10551,N_10385,N_10267);
and U10552 (N_10552,N_10275,N_10363);
and U10553 (N_10553,N_10280,N_10217);
nor U10554 (N_10554,N_10243,N_10218);
nand U10555 (N_10555,N_10352,N_10269);
xor U10556 (N_10556,N_10279,N_10351);
and U10557 (N_10557,N_10289,N_10257);
or U10558 (N_10558,N_10380,N_10354);
nand U10559 (N_10559,N_10338,N_10225);
and U10560 (N_10560,N_10265,N_10396);
or U10561 (N_10561,N_10286,N_10226);
xor U10562 (N_10562,N_10252,N_10379);
nor U10563 (N_10563,N_10340,N_10390);
or U10564 (N_10564,N_10362,N_10297);
nor U10565 (N_10565,N_10312,N_10387);
nand U10566 (N_10566,N_10352,N_10294);
nor U10567 (N_10567,N_10277,N_10369);
xor U10568 (N_10568,N_10261,N_10333);
nor U10569 (N_10569,N_10341,N_10280);
nand U10570 (N_10570,N_10293,N_10211);
nor U10571 (N_10571,N_10312,N_10234);
nand U10572 (N_10572,N_10313,N_10384);
and U10573 (N_10573,N_10318,N_10214);
nand U10574 (N_10574,N_10268,N_10296);
nand U10575 (N_10575,N_10327,N_10249);
and U10576 (N_10576,N_10200,N_10330);
or U10577 (N_10577,N_10229,N_10387);
or U10578 (N_10578,N_10216,N_10277);
and U10579 (N_10579,N_10270,N_10219);
or U10580 (N_10580,N_10273,N_10314);
nor U10581 (N_10581,N_10221,N_10288);
nor U10582 (N_10582,N_10231,N_10245);
nand U10583 (N_10583,N_10349,N_10288);
xnor U10584 (N_10584,N_10276,N_10201);
nand U10585 (N_10585,N_10392,N_10236);
and U10586 (N_10586,N_10384,N_10378);
nor U10587 (N_10587,N_10213,N_10349);
nor U10588 (N_10588,N_10200,N_10272);
nor U10589 (N_10589,N_10376,N_10310);
and U10590 (N_10590,N_10307,N_10387);
and U10591 (N_10591,N_10221,N_10273);
xnor U10592 (N_10592,N_10239,N_10373);
or U10593 (N_10593,N_10259,N_10322);
xor U10594 (N_10594,N_10366,N_10324);
nand U10595 (N_10595,N_10200,N_10326);
or U10596 (N_10596,N_10276,N_10389);
xor U10597 (N_10597,N_10269,N_10208);
or U10598 (N_10598,N_10283,N_10334);
nor U10599 (N_10599,N_10273,N_10352);
and U10600 (N_10600,N_10400,N_10423);
and U10601 (N_10601,N_10419,N_10584);
nand U10602 (N_10602,N_10441,N_10598);
xor U10603 (N_10603,N_10413,N_10477);
nor U10604 (N_10604,N_10556,N_10575);
nand U10605 (N_10605,N_10593,N_10469);
nor U10606 (N_10606,N_10591,N_10425);
or U10607 (N_10607,N_10481,N_10555);
nand U10608 (N_10608,N_10544,N_10523);
or U10609 (N_10609,N_10527,N_10572);
nor U10610 (N_10610,N_10532,N_10518);
nand U10611 (N_10611,N_10447,N_10459);
nand U10612 (N_10612,N_10581,N_10507);
nand U10613 (N_10613,N_10424,N_10466);
and U10614 (N_10614,N_10467,N_10534);
nand U10615 (N_10615,N_10512,N_10509);
or U10616 (N_10616,N_10434,N_10546);
xor U10617 (N_10617,N_10588,N_10574);
nand U10618 (N_10618,N_10548,N_10498);
xor U10619 (N_10619,N_10590,N_10449);
and U10620 (N_10620,N_10409,N_10420);
or U10621 (N_10621,N_10484,N_10433);
nand U10622 (N_10622,N_10554,N_10583);
nor U10623 (N_10623,N_10442,N_10472);
or U10624 (N_10624,N_10489,N_10520);
or U10625 (N_10625,N_10460,N_10525);
nand U10626 (N_10626,N_10547,N_10476);
and U10627 (N_10627,N_10511,N_10402);
nand U10628 (N_10628,N_10506,N_10415);
and U10629 (N_10629,N_10505,N_10437);
xnor U10630 (N_10630,N_10439,N_10464);
nand U10631 (N_10631,N_10465,N_10570);
and U10632 (N_10632,N_10566,N_10474);
nor U10633 (N_10633,N_10597,N_10430);
nand U10634 (N_10634,N_10411,N_10488);
and U10635 (N_10635,N_10595,N_10564);
and U10636 (N_10636,N_10542,N_10559);
nor U10637 (N_10637,N_10526,N_10568);
or U10638 (N_10638,N_10428,N_10475);
nand U10639 (N_10639,N_10596,N_10443);
nor U10640 (N_10640,N_10471,N_10516);
and U10641 (N_10641,N_10500,N_10426);
and U10642 (N_10642,N_10578,N_10462);
nor U10643 (N_10643,N_10470,N_10493);
and U10644 (N_10644,N_10579,N_10448);
and U10645 (N_10645,N_10401,N_10435);
nand U10646 (N_10646,N_10478,N_10536);
nor U10647 (N_10647,N_10504,N_10586);
nand U10648 (N_10648,N_10561,N_10533);
or U10649 (N_10649,N_10514,N_10582);
and U10650 (N_10650,N_10496,N_10427);
and U10651 (N_10651,N_10454,N_10497);
nor U10652 (N_10652,N_10589,N_10529);
nor U10653 (N_10653,N_10412,N_10416);
or U10654 (N_10654,N_10531,N_10524);
and U10655 (N_10655,N_10587,N_10408);
or U10656 (N_10656,N_10431,N_10456);
or U10657 (N_10657,N_10539,N_10557);
nor U10658 (N_10658,N_10594,N_10445);
nor U10659 (N_10659,N_10510,N_10545);
or U10660 (N_10660,N_10501,N_10487);
nor U10661 (N_10661,N_10499,N_10463);
and U10662 (N_10662,N_10453,N_10440);
nand U10663 (N_10663,N_10451,N_10490);
and U10664 (N_10664,N_10502,N_10492);
nand U10665 (N_10665,N_10418,N_10436);
and U10666 (N_10666,N_10558,N_10535);
nor U10667 (N_10667,N_10513,N_10553);
or U10668 (N_10668,N_10521,N_10452);
nor U10669 (N_10669,N_10563,N_10414);
nor U10670 (N_10670,N_10551,N_10486);
nand U10671 (N_10671,N_10599,N_10543);
nor U10672 (N_10672,N_10494,N_10585);
nor U10673 (N_10673,N_10483,N_10573);
nor U10674 (N_10674,N_10468,N_10491);
nand U10675 (N_10675,N_10580,N_10571);
and U10676 (N_10676,N_10576,N_10519);
and U10677 (N_10677,N_10417,N_10495);
nand U10678 (N_10678,N_10549,N_10565);
and U10679 (N_10679,N_10405,N_10569);
or U10680 (N_10680,N_10457,N_10567);
or U10681 (N_10681,N_10410,N_10403);
nor U10682 (N_10682,N_10530,N_10482);
or U10683 (N_10683,N_10577,N_10480);
nor U10684 (N_10684,N_10517,N_10446);
or U10685 (N_10685,N_10528,N_10508);
and U10686 (N_10686,N_10406,N_10438);
nor U10687 (N_10687,N_10429,N_10540);
and U10688 (N_10688,N_10404,N_10538);
nand U10689 (N_10689,N_10422,N_10562);
nor U10690 (N_10690,N_10421,N_10485);
nor U10691 (N_10691,N_10473,N_10515);
or U10692 (N_10692,N_10503,N_10541);
and U10693 (N_10693,N_10444,N_10560);
xnor U10694 (N_10694,N_10537,N_10552);
nand U10695 (N_10695,N_10432,N_10458);
xor U10696 (N_10696,N_10550,N_10461);
nand U10697 (N_10697,N_10450,N_10455);
nand U10698 (N_10698,N_10522,N_10592);
or U10699 (N_10699,N_10407,N_10479);
and U10700 (N_10700,N_10511,N_10573);
and U10701 (N_10701,N_10508,N_10599);
xnor U10702 (N_10702,N_10530,N_10571);
xnor U10703 (N_10703,N_10510,N_10448);
nand U10704 (N_10704,N_10542,N_10480);
and U10705 (N_10705,N_10473,N_10456);
or U10706 (N_10706,N_10422,N_10528);
or U10707 (N_10707,N_10500,N_10458);
nand U10708 (N_10708,N_10473,N_10508);
nand U10709 (N_10709,N_10410,N_10412);
and U10710 (N_10710,N_10596,N_10590);
nand U10711 (N_10711,N_10592,N_10486);
or U10712 (N_10712,N_10539,N_10568);
and U10713 (N_10713,N_10493,N_10590);
xnor U10714 (N_10714,N_10507,N_10555);
nor U10715 (N_10715,N_10452,N_10538);
or U10716 (N_10716,N_10460,N_10487);
or U10717 (N_10717,N_10445,N_10415);
and U10718 (N_10718,N_10567,N_10494);
or U10719 (N_10719,N_10557,N_10444);
or U10720 (N_10720,N_10595,N_10447);
or U10721 (N_10721,N_10404,N_10425);
nor U10722 (N_10722,N_10556,N_10573);
and U10723 (N_10723,N_10582,N_10578);
and U10724 (N_10724,N_10530,N_10465);
nand U10725 (N_10725,N_10410,N_10451);
nor U10726 (N_10726,N_10431,N_10586);
and U10727 (N_10727,N_10531,N_10400);
nand U10728 (N_10728,N_10481,N_10540);
or U10729 (N_10729,N_10539,N_10453);
nand U10730 (N_10730,N_10483,N_10418);
xor U10731 (N_10731,N_10577,N_10542);
nand U10732 (N_10732,N_10512,N_10470);
or U10733 (N_10733,N_10577,N_10475);
nand U10734 (N_10734,N_10585,N_10450);
xor U10735 (N_10735,N_10457,N_10418);
or U10736 (N_10736,N_10571,N_10406);
or U10737 (N_10737,N_10538,N_10565);
nor U10738 (N_10738,N_10412,N_10531);
and U10739 (N_10739,N_10580,N_10425);
and U10740 (N_10740,N_10538,N_10557);
xor U10741 (N_10741,N_10444,N_10518);
nor U10742 (N_10742,N_10571,N_10557);
nand U10743 (N_10743,N_10575,N_10510);
xnor U10744 (N_10744,N_10477,N_10447);
and U10745 (N_10745,N_10404,N_10598);
nand U10746 (N_10746,N_10423,N_10430);
nor U10747 (N_10747,N_10492,N_10501);
or U10748 (N_10748,N_10438,N_10533);
nor U10749 (N_10749,N_10501,N_10491);
xnor U10750 (N_10750,N_10418,N_10515);
or U10751 (N_10751,N_10558,N_10427);
and U10752 (N_10752,N_10560,N_10528);
and U10753 (N_10753,N_10450,N_10476);
nor U10754 (N_10754,N_10572,N_10403);
or U10755 (N_10755,N_10566,N_10596);
or U10756 (N_10756,N_10429,N_10418);
nor U10757 (N_10757,N_10531,N_10573);
nor U10758 (N_10758,N_10593,N_10559);
nor U10759 (N_10759,N_10413,N_10587);
xor U10760 (N_10760,N_10465,N_10406);
and U10761 (N_10761,N_10556,N_10433);
and U10762 (N_10762,N_10428,N_10404);
nand U10763 (N_10763,N_10417,N_10420);
nor U10764 (N_10764,N_10488,N_10472);
nor U10765 (N_10765,N_10529,N_10448);
and U10766 (N_10766,N_10592,N_10524);
or U10767 (N_10767,N_10584,N_10427);
and U10768 (N_10768,N_10441,N_10582);
nand U10769 (N_10769,N_10440,N_10441);
or U10770 (N_10770,N_10514,N_10442);
nor U10771 (N_10771,N_10422,N_10522);
and U10772 (N_10772,N_10421,N_10588);
nor U10773 (N_10773,N_10562,N_10470);
or U10774 (N_10774,N_10433,N_10515);
nor U10775 (N_10775,N_10581,N_10583);
and U10776 (N_10776,N_10502,N_10554);
nand U10777 (N_10777,N_10575,N_10555);
xnor U10778 (N_10778,N_10561,N_10598);
nand U10779 (N_10779,N_10450,N_10459);
nor U10780 (N_10780,N_10480,N_10567);
nor U10781 (N_10781,N_10533,N_10593);
and U10782 (N_10782,N_10481,N_10580);
nor U10783 (N_10783,N_10416,N_10508);
nor U10784 (N_10784,N_10518,N_10421);
nand U10785 (N_10785,N_10546,N_10509);
or U10786 (N_10786,N_10546,N_10584);
and U10787 (N_10787,N_10546,N_10409);
nand U10788 (N_10788,N_10422,N_10456);
or U10789 (N_10789,N_10538,N_10471);
or U10790 (N_10790,N_10457,N_10557);
xor U10791 (N_10791,N_10483,N_10441);
and U10792 (N_10792,N_10462,N_10487);
and U10793 (N_10793,N_10576,N_10588);
and U10794 (N_10794,N_10435,N_10428);
nand U10795 (N_10795,N_10481,N_10419);
nand U10796 (N_10796,N_10452,N_10472);
nor U10797 (N_10797,N_10593,N_10445);
xor U10798 (N_10798,N_10524,N_10445);
or U10799 (N_10799,N_10513,N_10463);
nor U10800 (N_10800,N_10782,N_10742);
and U10801 (N_10801,N_10746,N_10606);
nor U10802 (N_10802,N_10763,N_10664);
nor U10803 (N_10803,N_10766,N_10645);
nand U10804 (N_10804,N_10699,N_10663);
or U10805 (N_10805,N_10736,N_10604);
or U10806 (N_10806,N_10776,N_10647);
nor U10807 (N_10807,N_10637,N_10760);
nor U10808 (N_10808,N_10773,N_10695);
nor U10809 (N_10809,N_10761,N_10702);
or U10810 (N_10810,N_10709,N_10780);
nand U10811 (N_10811,N_10603,N_10779);
nand U10812 (N_10812,N_10751,N_10651);
nand U10813 (N_10813,N_10687,N_10667);
xor U10814 (N_10814,N_10798,N_10661);
xnor U10815 (N_10815,N_10639,N_10697);
nand U10816 (N_10816,N_10731,N_10660);
nand U10817 (N_10817,N_10656,N_10605);
and U10818 (N_10818,N_10655,N_10725);
or U10819 (N_10819,N_10619,N_10690);
nor U10820 (N_10820,N_10646,N_10648);
nand U10821 (N_10821,N_10737,N_10629);
nand U10822 (N_10822,N_10719,N_10749);
nand U10823 (N_10823,N_10640,N_10723);
nand U10824 (N_10824,N_10627,N_10630);
and U10825 (N_10825,N_10633,N_10693);
nor U10826 (N_10826,N_10700,N_10724);
or U10827 (N_10827,N_10718,N_10613);
nor U10828 (N_10828,N_10675,N_10673);
and U10829 (N_10829,N_10621,N_10715);
nand U10830 (N_10830,N_10796,N_10712);
or U10831 (N_10831,N_10786,N_10743);
nand U10832 (N_10832,N_10741,N_10703);
nor U10833 (N_10833,N_10623,N_10626);
or U10834 (N_10834,N_10711,N_10602);
and U10835 (N_10835,N_10654,N_10767);
nand U10836 (N_10836,N_10642,N_10608);
nor U10837 (N_10837,N_10616,N_10735);
and U10838 (N_10838,N_10748,N_10789);
nor U10839 (N_10839,N_10634,N_10682);
nand U10840 (N_10840,N_10686,N_10730);
and U10841 (N_10841,N_10706,N_10607);
and U10842 (N_10842,N_10618,N_10774);
xor U10843 (N_10843,N_10681,N_10657);
and U10844 (N_10844,N_10745,N_10747);
xnor U10845 (N_10845,N_10768,N_10707);
nand U10846 (N_10846,N_10732,N_10728);
nor U10847 (N_10847,N_10775,N_10729);
or U10848 (N_10848,N_10635,N_10674);
nor U10849 (N_10849,N_10788,N_10609);
nand U10850 (N_10850,N_10678,N_10722);
and U10851 (N_10851,N_10636,N_10754);
and U10852 (N_10852,N_10644,N_10666);
or U10853 (N_10853,N_10701,N_10600);
or U10854 (N_10854,N_10791,N_10790);
xor U10855 (N_10855,N_10787,N_10772);
or U10856 (N_10856,N_10659,N_10755);
or U10857 (N_10857,N_10759,N_10658);
nor U10858 (N_10858,N_10739,N_10713);
nor U10859 (N_10859,N_10727,N_10710);
or U10860 (N_10860,N_10696,N_10641);
nor U10861 (N_10861,N_10676,N_10677);
nand U10862 (N_10862,N_10762,N_10714);
xor U10863 (N_10863,N_10781,N_10670);
nor U10864 (N_10864,N_10794,N_10669);
or U10865 (N_10865,N_10643,N_10756);
or U10866 (N_10866,N_10601,N_10679);
xnor U10867 (N_10867,N_10705,N_10784);
nor U10868 (N_10868,N_10716,N_10615);
nand U10869 (N_10869,N_10769,N_10620);
nand U10870 (N_10870,N_10720,N_10684);
nand U10871 (N_10871,N_10792,N_10622);
or U10872 (N_10872,N_10764,N_10752);
nor U10873 (N_10873,N_10708,N_10691);
nand U10874 (N_10874,N_10785,N_10704);
or U10875 (N_10875,N_10793,N_10628);
xnor U10876 (N_10876,N_10611,N_10738);
or U10877 (N_10877,N_10668,N_10653);
nand U10878 (N_10878,N_10649,N_10744);
and U10879 (N_10879,N_10617,N_10631);
and U10880 (N_10880,N_10650,N_10770);
xor U10881 (N_10881,N_10671,N_10777);
and U10882 (N_10882,N_10689,N_10758);
nand U10883 (N_10883,N_10688,N_10625);
nor U10884 (N_10884,N_10624,N_10638);
and U10885 (N_10885,N_10717,N_10614);
nand U10886 (N_10886,N_10795,N_10778);
nand U10887 (N_10887,N_10610,N_10721);
nor U10888 (N_10888,N_10652,N_10632);
or U10889 (N_10889,N_10680,N_10683);
and U10890 (N_10890,N_10692,N_10797);
xor U10891 (N_10891,N_10662,N_10665);
nor U10892 (N_10892,N_10733,N_10734);
xnor U10893 (N_10893,N_10765,N_10771);
nor U10894 (N_10894,N_10740,N_10750);
or U10895 (N_10895,N_10685,N_10757);
nand U10896 (N_10896,N_10612,N_10783);
or U10897 (N_10897,N_10694,N_10672);
and U10898 (N_10898,N_10726,N_10698);
and U10899 (N_10899,N_10753,N_10799);
nor U10900 (N_10900,N_10775,N_10713);
or U10901 (N_10901,N_10638,N_10659);
and U10902 (N_10902,N_10703,N_10641);
nand U10903 (N_10903,N_10678,N_10681);
or U10904 (N_10904,N_10744,N_10701);
nor U10905 (N_10905,N_10644,N_10693);
nor U10906 (N_10906,N_10641,N_10631);
or U10907 (N_10907,N_10745,N_10689);
or U10908 (N_10908,N_10645,N_10719);
nand U10909 (N_10909,N_10717,N_10709);
and U10910 (N_10910,N_10780,N_10696);
nor U10911 (N_10911,N_10729,N_10606);
xnor U10912 (N_10912,N_10767,N_10677);
nand U10913 (N_10913,N_10784,N_10683);
or U10914 (N_10914,N_10705,N_10771);
nor U10915 (N_10915,N_10670,N_10630);
nand U10916 (N_10916,N_10678,N_10714);
or U10917 (N_10917,N_10786,N_10639);
or U10918 (N_10918,N_10691,N_10783);
and U10919 (N_10919,N_10708,N_10744);
nand U10920 (N_10920,N_10695,N_10689);
nand U10921 (N_10921,N_10753,N_10685);
nand U10922 (N_10922,N_10666,N_10675);
nand U10923 (N_10923,N_10663,N_10636);
nor U10924 (N_10924,N_10619,N_10705);
nand U10925 (N_10925,N_10709,N_10600);
xor U10926 (N_10926,N_10752,N_10661);
and U10927 (N_10927,N_10715,N_10641);
nor U10928 (N_10928,N_10752,N_10686);
or U10929 (N_10929,N_10749,N_10720);
nor U10930 (N_10930,N_10732,N_10719);
nor U10931 (N_10931,N_10719,N_10726);
xnor U10932 (N_10932,N_10775,N_10787);
or U10933 (N_10933,N_10600,N_10637);
and U10934 (N_10934,N_10618,N_10788);
nand U10935 (N_10935,N_10748,N_10700);
and U10936 (N_10936,N_10681,N_10621);
nor U10937 (N_10937,N_10625,N_10779);
nand U10938 (N_10938,N_10640,N_10776);
nand U10939 (N_10939,N_10752,N_10727);
nor U10940 (N_10940,N_10672,N_10760);
or U10941 (N_10941,N_10794,N_10632);
xnor U10942 (N_10942,N_10747,N_10751);
and U10943 (N_10943,N_10781,N_10700);
and U10944 (N_10944,N_10749,N_10751);
and U10945 (N_10945,N_10705,N_10675);
and U10946 (N_10946,N_10716,N_10641);
nand U10947 (N_10947,N_10628,N_10712);
nor U10948 (N_10948,N_10632,N_10763);
nor U10949 (N_10949,N_10660,N_10753);
xnor U10950 (N_10950,N_10758,N_10757);
xnor U10951 (N_10951,N_10751,N_10786);
or U10952 (N_10952,N_10787,N_10736);
or U10953 (N_10953,N_10656,N_10611);
nand U10954 (N_10954,N_10679,N_10796);
and U10955 (N_10955,N_10712,N_10692);
and U10956 (N_10956,N_10718,N_10654);
or U10957 (N_10957,N_10649,N_10717);
xnor U10958 (N_10958,N_10635,N_10784);
and U10959 (N_10959,N_10607,N_10630);
xnor U10960 (N_10960,N_10763,N_10658);
nand U10961 (N_10961,N_10678,N_10676);
or U10962 (N_10962,N_10686,N_10609);
nand U10963 (N_10963,N_10706,N_10700);
or U10964 (N_10964,N_10754,N_10669);
nor U10965 (N_10965,N_10796,N_10657);
and U10966 (N_10966,N_10736,N_10716);
or U10967 (N_10967,N_10764,N_10775);
and U10968 (N_10968,N_10752,N_10636);
and U10969 (N_10969,N_10622,N_10692);
nand U10970 (N_10970,N_10734,N_10621);
or U10971 (N_10971,N_10784,N_10704);
nor U10972 (N_10972,N_10693,N_10722);
or U10973 (N_10973,N_10700,N_10622);
xor U10974 (N_10974,N_10686,N_10646);
or U10975 (N_10975,N_10789,N_10626);
nor U10976 (N_10976,N_10768,N_10687);
or U10977 (N_10977,N_10760,N_10617);
or U10978 (N_10978,N_10673,N_10758);
and U10979 (N_10979,N_10790,N_10617);
nand U10980 (N_10980,N_10732,N_10620);
nand U10981 (N_10981,N_10671,N_10709);
nor U10982 (N_10982,N_10641,N_10785);
or U10983 (N_10983,N_10693,N_10636);
nand U10984 (N_10984,N_10703,N_10797);
nand U10985 (N_10985,N_10767,N_10700);
and U10986 (N_10986,N_10648,N_10604);
nor U10987 (N_10987,N_10636,N_10686);
nand U10988 (N_10988,N_10715,N_10763);
and U10989 (N_10989,N_10744,N_10700);
or U10990 (N_10990,N_10751,N_10788);
and U10991 (N_10991,N_10656,N_10703);
nand U10992 (N_10992,N_10681,N_10622);
and U10993 (N_10993,N_10755,N_10741);
nand U10994 (N_10994,N_10739,N_10775);
and U10995 (N_10995,N_10779,N_10792);
nand U10996 (N_10996,N_10728,N_10775);
and U10997 (N_10997,N_10753,N_10698);
or U10998 (N_10998,N_10784,N_10644);
nor U10999 (N_10999,N_10770,N_10649);
nand U11000 (N_11000,N_10955,N_10968);
nor U11001 (N_11001,N_10857,N_10874);
or U11002 (N_11002,N_10837,N_10861);
xnor U11003 (N_11003,N_10970,N_10981);
and U11004 (N_11004,N_10890,N_10954);
and U11005 (N_11005,N_10994,N_10905);
xor U11006 (N_11006,N_10871,N_10953);
or U11007 (N_11007,N_10863,N_10891);
or U11008 (N_11008,N_10928,N_10849);
or U11009 (N_11009,N_10851,N_10864);
or U11010 (N_11010,N_10895,N_10937);
or U11011 (N_11011,N_10848,N_10836);
xnor U11012 (N_11012,N_10920,N_10912);
nor U11013 (N_11013,N_10831,N_10972);
or U11014 (N_11014,N_10971,N_10870);
nand U11015 (N_11015,N_10974,N_10804);
nand U11016 (N_11016,N_10860,N_10850);
nand U11017 (N_11017,N_10923,N_10884);
and U11018 (N_11018,N_10975,N_10980);
xnor U11019 (N_11019,N_10946,N_10852);
or U11020 (N_11020,N_10883,N_10840);
or U11021 (N_11021,N_10800,N_10957);
or U11022 (N_11022,N_10872,N_10993);
xor U11023 (N_11023,N_10992,N_10806);
and U11024 (N_11024,N_10940,N_10941);
and U11025 (N_11025,N_10931,N_10896);
or U11026 (N_11026,N_10939,N_10904);
or U11027 (N_11027,N_10906,N_10965);
or U11028 (N_11028,N_10911,N_10832);
nand U11029 (N_11029,N_10997,N_10828);
or U11030 (N_11030,N_10844,N_10914);
nor U11031 (N_11031,N_10983,N_10805);
nand U11032 (N_11032,N_10926,N_10976);
nor U11033 (N_11033,N_10986,N_10809);
or U11034 (N_11034,N_10846,N_10973);
xnor U11035 (N_11035,N_10877,N_10936);
xnor U11036 (N_11036,N_10990,N_10902);
and U11037 (N_11037,N_10982,N_10934);
or U11038 (N_11038,N_10803,N_10922);
nor U11039 (N_11039,N_10819,N_10995);
nand U11040 (N_11040,N_10996,N_10894);
xor U11041 (N_11041,N_10862,N_10908);
nor U11042 (N_11042,N_10897,N_10878);
and U11043 (N_11043,N_10948,N_10901);
and U11044 (N_11044,N_10821,N_10917);
nor U11045 (N_11045,N_10817,N_10930);
xor U11046 (N_11046,N_10873,N_10811);
or U11047 (N_11047,N_10845,N_10825);
nor U11048 (N_11048,N_10885,N_10909);
nor U11049 (N_11049,N_10812,N_10814);
and U11050 (N_11050,N_10964,N_10918);
or U11051 (N_11051,N_10867,N_10991);
nor U11052 (N_11052,N_10869,N_10838);
nand U11053 (N_11053,N_10888,N_10855);
and U11054 (N_11054,N_10924,N_10898);
or U11055 (N_11055,N_10858,N_10969);
or U11056 (N_11056,N_10932,N_10816);
nor U11057 (N_11057,N_10903,N_10960);
and U11058 (N_11058,N_10900,N_10826);
and U11059 (N_11059,N_10835,N_10985);
nand U11060 (N_11060,N_10886,N_10933);
and U11061 (N_11061,N_10944,N_10829);
and U11062 (N_11062,N_10843,N_10979);
and U11063 (N_11063,N_10899,N_10802);
nand U11064 (N_11064,N_10929,N_10810);
or U11065 (N_11065,N_10833,N_10892);
nand U11066 (N_11066,N_10988,N_10967);
nand U11067 (N_11067,N_10998,N_10868);
xnor U11068 (N_11068,N_10919,N_10824);
nand U11069 (N_11069,N_10882,N_10977);
or U11070 (N_11070,N_10916,N_10949);
and U11071 (N_11071,N_10818,N_10910);
xnor U11072 (N_11072,N_10854,N_10841);
or U11073 (N_11073,N_10842,N_10875);
and U11074 (N_11074,N_10834,N_10925);
or U11075 (N_11075,N_10952,N_10889);
and U11076 (N_11076,N_10856,N_10943);
nand U11077 (N_11077,N_10963,N_10915);
or U11078 (N_11078,N_10820,N_10950);
or U11079 (N_11079,N_10847,N_10879);
and U11080 (N_11080,N_10999,N_10853);
nand U11081 (N_11081,N_10951,N_10815);
nand U11082 (N_11082,N_10984,N_10830);
and U11083 (N_11083,N_10987,N_10876);
or U11084 (N_11084,N_10813,N_10959);
nor U11085 (N_11085,N_10989,N_10801);
or U11086 (N_11086,N_10807,N_10822);
nand U11087 (N_11087,N_10827,N_10956);
xor U11088 (N_11088,N_10887,N_10938);
and U11089 (N_11089,N_10913,N_10966);
and U11090 (N_11090,N_10893,N_10927);
and U11091 (N_11091,N_10942,N_10958);
or U11092 (N_11092,N_10961,N_10823);
nand U11093 (N_11093,N_10880,N_10865);
and U11094 (N_11094,N_10808,N_10859);
nor U11095 (N_11095,N_10947,N_10839);
nor U11096 (N_11096,N_10945,N_10935);
nand U11097 (N_11097,N_10962,N_10907);
or U11098 (N_11098,N_10881,N_10978);
nor U11099 (N_11099,N_10866,N_10921);
nor U11100 (N_11100,N_10819,N_10987);
nor U11101 (N_11101,N_10911,N_10881);
or U11102 (N_11102,N_10952,N_10804);
and U11103 (N_11103,N_10971,N_10898);
nand U11104 (N_11104,N_10952,N_10956);
xnor U11105 (N_11105,N_10843,N_10900);
nor U11106 (N_11106,N_10935,N_10883);
nand U11107 (N_11107,N_10962,N_10979);
xnor U11108 (N_11108,N_10978,N_10951);
xnor U11109 (N_11109,N_10917,N_10822);
nand U11110 (N_11110,N_10844,N_10865);
nand U11111 (N_11111,N_10812,N_10872);
and U11112 (N_11112,N_10846,N_10912);
or U11113 (N_11113,N_10869,N_10848);
and U11114 (N_11114,N_10987,N_10887);
and U11115 (N_11115,N_10861,N_10852);
xnor U11116 (N_11116,N_10822,N_10804);
or U11117 (N_11117,N_10832,N_10876);
or U11118 (N_11118,N_10874,N_10839);
nand U11119 (N_11119,N_10876,N_10846);
nand U11120 (N_11120,N_10886,N_10917);
nor U11121 (N_11121,N_10916,N_10802);
xnor U11122 (N_11122,N_10853,N_10973);
nor U11123 (N_11123,N_10872,N_10867);
and U11124 (N_11124,N_10874,N_10966);
nand U11125 (N_11125,N_10990,N_10822);
nand U11126 (N_11126,N_10908,N_10851);
or U11127 (N_11127,N_10863,N_10879);
nor U11128 (N_11128,N_10845,N_10831);
and U11129 (N_11129,N_10831,N_10852);
or U11130 (N_11130,N_10849,N_10942);
nor U11131 (N_11131,N_10932,N_10943);
or U11132 (N_11132,N_10832,N_10857);
nand U11133 (N_11133,N_10908,N_10932);
and U11134 (N_11134,N_10834,N_10923);
xnor U11135 (N_11135,N_10842,N_10938);
nor U11136 (N_11136,N_10861,N_10882);
xor U11137 (N_11137,N_10855,N_10816);
or U11138 (N_11138,N_10828,N_10870);
and U11139 (N_11139,N_10929,N_10934);
and U11140 (N_11140,N_10918,N_10881);
nor U11141 (N_11141,N_10859,N_10992);
nor U11142 (N_11142,N_10827,N_10990);
or U11143 (N_11143,N_10856,N_10908);
and U11144 (N_11144,N_10918,N_10939);
xor U11145 (N_11145,N_10955,N_10986);
nand U11146 (N_11146,N_10984,N_10966);
and U11147 (N_11147,N_10937,N_10865);
and U11148 (N_11148,N_10898,N_10982);
and U11149 (N_11149,N_10925,N_10895);
nand U11150 (N_11150,N_10855,N_10806);
or U11151 (N_11151,N_10931,N_10997);
nand U11152 (N_11152,N_10815,N_10835);
nor U11153 (N_11153,N_10864,N_10872);
nand U11154 (N_11154,N_10995,N_10999);
nor U11155 (N_11155,N_10871,N_10982);
and U11156 (N_11156,N_10843,N_10941);
or U11157 (N_11157,N_10874,N_10908);
nor U11158 (N_11158,N_10958,N_10820);
nand U11159 (N_11159,N_10884,N_10811);
nand U11160 (N_11160,N_10912,N_10976);
nand U11161 (N_11161,N_10907,N_10812);
and U11162 (N_11162,N_10924,N_10879);
nor U11163 (N_11163,N_10979,N_10828);
nand U11164 (N_11164,N_10827,N_10811);
and U11165 (N_11165,N_10819,N_10806);
or U11166 (N_11166,N_10990,N_10905);
or U11167 (N_11167,N_10956,N_10866);
and U11168 (N_11168,N_10939,N_10943);
nand U11169 (N_11169,N_10936,N_10896);
nand U11170 (N_11170,N_10972,N_10886);
and U11171 (N_11171,N_10816,N_10891);
or U11172 (N_11172,N_10888,N_10865);
or U11173 (N_11173,N_10838,N_10866);
and U11174 (N_11174,N_10803,N_10956);
xor U11175 (N_11175,N_10946,N_10949);
nand U11176 (N_11176,N_10835,N_10851);
nor U11177 (N_11177,N_10829,N_10903);
and U11178 (N_11178,N_10913,N_10919);
and U11179 (N_11179,N_10982,N_10821);
nor U11180 (N_11180,N_10909,N_10907);
nand U11181 (N_11181,N_10944,N_10940);
nand U11182 (N_11182,N_10896,N_10993);
nand U11183 (N_11183,N_10953,N_10838);
nand U11184 (N_11184,N_10899,N_10876);
or U11185 (N_11185,N_10956,N_10985);
xnor U11186 (N_11186,N_10953,N_10969);
nor U11187 (N_11187,N_10835,N_10859);
xnor U11188 (N_11188,N_10966,N_10959);
or U11189 (N_11189,N_10850,N_10830);
or U11190 (N_11190,N_10848,N_10855);
xor U11191 (N_11191,N_10856,N_10845);
xnor U11192 (N_11192,N_10929,N_10831);
and U11193 (N_11193,N_10867,N_10965);
nor U11194 (N_11194,N_10930,N_10889);
and U11195 (N_11195,N_10813,N_10968);
nand U11196 (N_11196,N_10947,N_10973);
nand U11197 (N_11197,N_10857,N_10815);
or U11198 (N_11198,N_10972,N_10871);
xor U11199 (N_11199,N_10832,N_10870);
and U11200 (N_11200,N_11097,N_11027);
xnor U11201 (N_11201,N_11089,N_11045);
nor U11202 (N_11202,N_11128,N_11121);
nand U11203 (N_11203,N_11088,N_11002);
nor U11204 (N_11204,N_11197,N_11174);
nor U11205 (N_11205,N_11050,N_11185);
and U11206 (N_11206,N_11099,N_11077);
and U11207 (N_11207,N_11102,N_11169);
nor U11208 (N_11208,N_11084,N_11113);
or U11209 (N_11209,N_11031,N_11017);
xnor U11210 (N_11210,N_11042,N_11131);
and U11211 (N_11211,N_11104,N_11076);
nor U11212 (N_11212,N_11028,N_11044);
and U11213 (N_11213,N_11082,N_11153);
nand U11214 (N_11214,N_11091,N_11090);
nand U11215 (N_11215,N_11190,N_11086);
nand U11216 (N_11216,N_11036,N_11168);
nor U11217 (N_11217,N_11160,N_11046);
and U11218 (N_11218,N_11182,N_11196);
or U11219 (N_11219,N_11134,N_11101);
xnor U11220 (N_11220,N_11054,N_11038);
or U11221 (N_11221,N_11195,N_11058);
and U11222 (N_11222,N_11126,N_11175);
and U11223 (N_11223,N_11110,N_11149);
nand U11224 (N_11224,N_11093,N_11188);
and U11225 (N_11225,N_11192,N_11105);
nor U11226 (N_11226,N_11194,N_11062);
nor U11227 (N_11227,N_11164,N_11114);
nand U11228 (N_11228,N_11103,N_11141);
nand U11229 (N_11229,N_11096,N_11193);
nand U11230 (N_11230,N_11095,N_11001);
nor U11231 (N_11231,N_11184,N_11008);
or U11232 (N_11232,N_11063,N_11068);
and U11233 (N_11233,N_11013,N_11030);
or U11234 (N_11234,N_11047,N_11145);
xnor U11235 (N_11235,N_11150,N_11041);
or U11236 (N_11236,N_11180,N_11032);
and U11237 (N_11237,N_11158,N_11018);
and U11238 (N_11238,N_11007,N_11163);
nand U11239 (N_11239,N_11187,N_11039);
and U11240 (N_11240,N_11026,N_11181);
and U11241 (N_11241,N_11074,N_11019);
or U11242 (N_11242,N_11132,N_11155);
and U11243 (N_11243,N_11080,N_11087);
nor U11244 (N_11244,N_11052,N_11198);
xor U11245 (N_11245,N_11170,N_11122);
nor U11246 (N_11246,N_11014,N_11064);
and U11247 (N_11247,N_11120,N_11067);
nand U11248 (N_11248,N_11124,N_11078);
and U11249 (N_11249,N_11159,N_11100);
or U11250 (N_11250,N_11025,N_11156);
or U11251 (N_11251,N_11112,N_11173);
nand U11252 (N_11252,N_11178,N_11119);
or U11253 (N_11253,N_11161,N_11053);
nor U11254 (N_11254,N_11075,N_11020);
or U11255 (N_11255,N_11094,N_11116);
or U11256 (N_11256,N_11006,N_11092);
and U11257 (N_11257,N_11166,N_11011);
or U11258 (N_11258,N_11154,N_11098);
nor U11259 (N_11259,N_11051,N_11033);
or U11260 (N_11260,N_11060,N_11136);
and U11261 (N_11261,N_11069,N_11133);
or U11262 (N_11262,N_11079,N_11171);
and U11263 (N_11263,N_11056,N_11138);
or U11264 (N_11264,N_11189,N_11143);
nor U11265 (N_11265,N_11117,N_11130);
or U11266 (N_11266,N_11003,N_11172);
xnor U11267 (N_11267,N_11123,N_11157);
nand U11268 (N_11268,N_11016,N_11043);
xor U11269 (N_11269,N_11035,N_11059);
nand U11270 (N_11270,N_11147,N_11081);
nand U11271 (N_11271,N_11167,N_11073);
or U11272 (N_11272,N_11176,N_11012);
nand U11273 (N_11273,N_11144,N_11024);
nand U11274 (N_11274,N_11152,N_11107);
or U11275 (N_11275,N_11106,N_11179);
and U11276 (N_11276,N_11040,N_11165);
xnor U11277 (N_11277,N_11135,N_11055);
and U11278 (N_11278,N_11191,N_11127);
nand U11279 (N_11279,N_11022,N_11111);
and U11280 (N_11280,N_11140,N_11009);
nand U11281 (N_11281,N_11139,N_11049);
or U11282 (N_11282,N_11129,N_11071);
and U11283 (N_11283,N_11072,N_11000);
or U11284 (N_11284,N_11186,N_11162);
nand U11285 (N_11285,N_11183,N_11057);
xor U11286 (N_11286,N_11065,N_11115);
and U11287 (N_11287,N_11021,N_11048);
nor U11288 (N_11288,N_11108,N_11137);
nor U11289 (N_11289,N_11085,N_11015);
and U11290 (N_11290,N_11109,N_11177);
nand U11291 (N_11291,N_11004,N_11034);
or U11292 (N_11292,N_11061,N_11010);
nor U11293 (N_11293,N_11151,N_11083);
nor U11294 (N_11294,N_11066,N_11070);
and U11295 (N_11295,N_11029,N_11148);
nor U11296 (N_11296,N_11125,N_11118);
nor U11297 (N_11297,N_11146,N_11005);
nor U11298 (N_11298,N_11037,N_11023);
nor U11299 (N_11299,N_11142,N_11199);
or U11300 (N_11300,N_11190,N_11029);
or U11301 (N_11301,N_11027,N_11015);
xor U11302 (N_11302,N_11017,N_11094);
xnor U11303 (N_11303,N_11028,N_11083);
nor U11304 (N_11304,N_11155,N_11147);
nor U11305 (N_11305,N_11123,N_11122);
xnor U11306 (N_11306,N_11062,N_11168);
or U11307 (N_11307,N_11125,N_11107);
nand U11308 (N_11308,N_11024,N_11109);
xor U11309 (N_11309,N_11184,N_11039);
and U11310 (N_11310,N_11010,N_11046);
nand U11311 (N_11311,N_11011,N_11152);
nand U11312 (N_11312,N_11088,N_11145);
and U11313 (N_11313,N_11059,N_11140);
and U11314 (N_11314,N_11089,N_11081);
nor U11315 (N_11315,N_11036,N_11054);
and U11316 (N_11316,N_11042,N_11023);
nor U11317 (N_11317,N_11178,N_11114);
nor U11318 (N_11318,N_11032,N_11060);
and U11319 (N_11319,N_11192,N_11125);
nor U11320 (N_11320,N_11164,N_11157);
or U11321 (N_11321,N_11014,N_11182);
nor U11322 (N_11322,N_11125,N_11018);
or U11323 (N_11323,N_11040,N_11176);
or U11324 (N_11324,N_11125,N_11157);
and U11325 (N_11325,N_11101,N_11000);
and U11326 (N_11326,N_11196,N_11066);
or U11327 (N_11327,N_11052,N_11089);
or U11328 (N_11328,N_11022,N_11152);
nand U11329 (N_11329,N_11158,N_11166);
nand U11330 (N_11330,N_11052,N_11154);
and U11331 (N_11331,N_11010,N_11066);
nand U11332 (N_11332,N_11195,N_11048);
nand U11333 (N_11333,N_11061,N_11139);
and U11334 (N_11334,N_11166,N_11027);
nor U11335 (N_11335,N_11015,N_11133);
and U11336 (N_11336,N_11055,N_11102);
and U11337 (N_11337,N_11072,N_11054);
xnor U11338 (N_11338,N_11197,N_11132);
nand U11339 (N_11339,N_11077,N_11034);
nand U11340 (N_11340,N_11092,N_11054);
and U11341 (N_11341,N_11067,N_11155);
nor U11342 (N_11342,N_11019,N_11041);
and U11343 (N_11343,N_11168,N_11012);
nor U11344 (N_11344,N_11159,N_11076);
nor U11345 (N_11345,N_11194,N_11013);
nand U11346 (N_11346,N_11134,N_11033);
nand U11347 (N_11347,N_11003,N_11110);
or U11348 (N_11348,N_11154,N_11119);
nand U11349 (N_11349,N_11030,N_11115);
xnor U11350 (N_11350,N_11124,N_11191);
nand U11351 (N_11351,N_11190,N_11163);
nor U11352 (N_11352,N_11109,N_11032);
xnor U11353 (N_11353,N_11115,N_11061);
and U11354 (N_11354,N_11140,N_11050);
nor U11355 (N_11355,N_11036,N_11047);
nor U11356 (N_11356,N_11001,N_11019);
and U11357 (N_11357,N_11089,N_11014);
and U11358 (N_11358,N_11103,N_11076);
nand U11359 (N_11359,N_11045,N_11193);
nor U11360 (N_11360,N_11194,N_11073);
and U11361 (N_11361,N_11137,N_11089);
nor U11362 (N_11362,N_11094,N_11097);
or U11363 (N_11363,N_11107,N_11157);
nand U11364 (N_11364,N_11161,N_11099);
nand U11365 (N_11365,N_11043,N_11179);
nand U11366 (N_11366,N_11058,N_11194);
and U11367 (N_11367,N_11134,N_11069);
or U11368 (N_11368,N_11099,N_11069);
or U11369 (N_11369,N_11111,N_11103);
or U11370 (N_11370,N_11151,N_11154);
nand U11371 (N_11371,N_11183,N_11181);
or U11372 (N_11372,N_11104,N_11162);
nand U11373 (N_11373,N_11081,N_11047);
nand U11374 (N_11374,N_11184,N_11139);
xnor U11375 (N_11375,N_11134,N_11110);
nand U11376 (N_11376,N_11082,N_11189);
xnor U11377 (N_11377,N_11193,N_11053);
nand U11378 (N_11378,N_11017,N_11168);
or U11379 (N_11379,N_11144,N_11081);
and U11380 (N_11380,N_11185,N_11016);
or U11381 (N_11381,N_11009,N_11157);
and U11382 (N_11382,N_11167,N_11054);
nand U11383 (N_11383,N_11187,N_11022);
nand U11384 (N_11384,N_11057,N_11096);
or U11385 (N_11385,N_11069,N_11025);
nand U11386 (N_11386,N_11130,N_11036);
or U11387 (N_11387,N_11170,N_11031);
nand U11388 (N_11388,N_11020,N_11097);
nor U11389 (N_11389,N_11061,N_11028);
or U11390 (N_11390,N_11097,N_11015);
and U11391 (N_11391,N_11044,N_11148);
nor U11392 (N_11392,N_11183,N_11192);
or U11393 (N_11393,N_11152,N_11190);
and U11394 (N_11394,N_11136,N_11077);
and U11395 (N_11395,N_11111,N_11015);
xor U11396 (N_11396,N_11135,N_11137);
xnor U11397 (N_11397,N_11026,N_11049);
and U11398 (N_11398,N_11139,N_11156);
or U11399 (N_11399,N_11082,N_11148);
and U11400 (N_11400,N_11258,N_11361);
nor U11401 (N_11401,N_11207,N_11319);
nand U11402 (N_11402,N_11392,N_11205);
xnor U11403 (N_11403,N_11275,N_11313);
nand U11404 (N_11404,N_11238,N_11263);
nor U11405 (N_11405,N_11375,N_11329);
or U11406 (N_11406,N_11236,N_11311);
xnor U11407 (N_11407,N_11269,N_11277);
and U11408 (N_11408,N_11298,N_11260);
nor U11409 (N_11409,N_11248,N_11334);
or U11410 (N_11410,N_11376,N_11374);
nor U11411 (N_11411,N_11208,N_11378);
and U11412 (N_11412,N_11367,N_11391);
xor U11413 (N_11413,N_11373,N_11371);
and U11414 (N_11414,N_11396,N_11237);
nand U11415 (N_11415,N_11301,N_11253);
or U11416 (N_11416,N_11251,N_11398);
or U11417 (N_11417,N_11384,N_11203);
nor U11418 (N_11418,N_11273,N_11234);
and U11419 (N_11419,N_11235,N_11302);
or U11420 (N_11420,N_11349,N_11315);
nor U11421 (N_11421,N_11383,N_11387);
and U11422 (N_11422,N_11330,N_11286);
and U11423 (N_11423,N_11229,N_11347);
nor U11424 (N_11424,N_11216,N_11249);
nor U11425 (N_11425,N_11252,N_11303);
or U11426 (N_11426,N_11210,N_11246);
and U11427 (N_11427,N_11346,N_11261);
or U11428 (N_11428,N_11356,N_11389);
or U11429 (N_11429,N_11395,N_11222);
xor U11430 (N_11430,N_11254,N_11358);
and U11431 (N_11431,N_11350,N_11285);
xor U11432 (N_11432,N_11227,N_11233);
nor U11433 (N_11433,N_11215,N_11245);
or U11434 (N_11434,N_11214,N_11368);
nor U11435 (N_11435,N_11364,N_11281);
xnor U11436 (N_11436,N_11316,N_11318);
and U11437 (N_11437,N_11354,N_11393);
nor U11438 (N_11438,N_11326,N_11381);
xor U11439 (N_11439,N_11306,N_11331);
and U11440 (N_11440,N_11265,N_11341);
and U11441 (N_11441,N_11336,N_11268);
nand U11442 (N_11442,N_11292,N_11217);
or U11443 (N_11443,N_11372,N_11399);
nor U11444 (N_11444,N_11266,N_11380);
or U11445 (N_11445,N_11325,N_11293);
and U11446 (N_11446,N_11312,N_11332);
or U11447 (N_11447,N_11212,N_11259);
xor U11448 (N_11448,N_11338,N_11213);
or U11449 (N_11449,N_11337,N_11239);
and U11450 (N_11450,N_11345,N_11369);
nand U11451 (N_11451,N_11230,N_11370);
nor U11452 (N_11452,N_11304,N_11226);
xor U11453 (N_11453,N_11328,N_11257);
nor U11454 (N_11454,N_11323,N_11224);
xnor U11455 (N_11455,N_11202,N_11355);
nand U11456 (N_11456,N_11225,N_11267);
nand U11457 (N_11457,N_11362,N_11218);
xor U11458 (N_11458,N_11223,N_11397);
nand U11459 (N_11459,N_11333,N_11282);
nand U11460 (N_11460,N_11250,N_11385);
and U11461 (N_11461,N_11348,N_11321);
nand U11462 (N_11462,N_11291,N_11296);
nor U11463 (N_11463,N_11324,N_11278);
or U11464 (N_11464,N_11309,N_11359);
xnor U11465 (N_11465,N_11287,N_11290);
nand U11466 (N_11466,N_11221,N_11271);
and U11467 (N_11467,N_11322,N_11240);
nor U11468 (N_11468,N_11360,N_11388);
or U11469 (N_11469,N_11289,N_11310);
and U11470 (N_11470,N_11283,N_11357);
or U11471 (N_11471,N_11200,N_11351);
nand U11472 (N_11472,N_11220,N_11307);
and U11473 (N_11473,N_11377,N_11294);
nand U11474 (N_11474,N_11255,N_11270);
and U11475 (N_11475,N_11242,N_11327);
nor U11476 (N_11476,N_11232,N_11305);
nand U11477 (N_11477,N_11386,N_11209);
and U11478 (N_11478,N_11335,N_11342);
or U11479 (N_11479,N_11264,N_11295);
or U11480 (N_11480,N_11276,N_11231);
nor U11481 (N_11481,N_11297,N_11272);
nand U11482 (N_11482,N_11344,N_11340);
and U11483 (N_11483,N_11320,N_11206);
nand U11484 (N_11484,N_11390,N_11274);
or U11485 (N_11485,N_11279,N_11314);
and U11486 (N_11486,N_11262,N_11204);
xor U11487 (N_11487,N_11299,N_11241);
xnor U11488 (N_11488,N_11382,N_11308);
nor U11489 (N_11489,N_11243,N_11363);
xor U11490 (N_11490,N_11366,N_11211);
or U11491 (N_11491,N_11244,N_11247);
nor U11492 (N_11492,N_11352,N_11394);
nand U11493 (N_11493,N_11280,N_11339);
xor U11494 (N_11494,N_11317,N_11379);
nand U11495 (N_11495,N_11219,N_11284);
nor U11496 (N_11496,N_11300,N_11343);
and U11497 (N_11497,N_11228,N_11353);
and U11498 (N_11498,N_11256,N_11288);
and U11499 (N_11499,N_11201,N_11365);
and U11500 (N_11500,N_11386,N_11298);
nand U11501 (N_11501,N_11227,N_11313);
and U11502 (N_11502,N_11343,N_11213);
xnor U11503 (N_11503,N_11372,N_11363);
and U11504 (N_11504,N_11235,N_11288);
and U11505 (N_11505,N_11324,N_11347);
or U11506 (N_11506,N_11276,N_11385);
and U11507 (N_11507,N_11285,N_11325);
nor U11508 (N_11508,N_11259,N_11272);
or U11509 (N_11509,N_11325,N_11284);
or U11510 (N_11510,N_11296,N_11216);
nor U11511 (N_11511,N_11268,N_11360);
and U11512 (N_11512,N_11313,N_11240);
xor U11513 (N_11513,N_11333,N_11287);
xnor U11514 (N_11514,N_11206,N_11279);
nand U11515 (N_11515,N_11354,N_11325);
and U11516 (N_11516,N_11337,N_11368);
or U11517 (N_11517,N_11332,N_11220);
or U11518 (N_11518,N_11290,N_11399);
nand U11519 (N_11519,N_11272,N_11273);
and U11520 (N_11520,N_11330,N_11321);
and U11521 (N_11521,N_11219,N_11389);
and U11522 (N_11522,N_11204,N_11336);
or U11523 (N_11523,N_11252,N_11316);
xor U11524 (N_11524,N_11285,N_11389);
and U11525 (N_11525,N_11270,N_11215);
nor U11526 (N_11526,N_11353,N_11234);
nor U11527 (N_11527,N_11212,N_11381);
nor U11528 (N_11528,N_11278,N_11379);
or U11529 (N_11529,N_11243,N_11258);
or U11530 (N_11530,N_11215,N_11274);
nand U11531 (N_11531,N_11273,N_11357);
and U11532 (N_11532,N_11286,N_11243);
nor U11533 (N_11533,N_11255,N_11242);
nand U11534 (N_11534,N_11319,N_11246);
or U11535 (N_11535,N_11358,N_11245);
xor U11536 (N_11536,N_11235,N_11202);
nand U11537 (N_11537,N_11202,N_11335);
nor U11538 (N_11538,N_11327,N_11307);
and U11539 (N_11539,N_11334,N_11201);
nand U11540 (N_11540,N_11311,N_11379);
nand U11541 (N_11541,N_11214,N_11309);
nand U11542 (N_11542,N_11329,N_11269);
nor U11543 (N_11543,N_11212,N_11210);
nor U11544 (N_11544,N_11281,N_11341);
or U11545 (N_11545,N_11385,N_11217);
nand U11546 (N_11546,N_11311,N_11368);
nor U11547 (N_11547,N_11250,N_11340);
or U11548 (N_11548,N_11224,N_11312);
nand U11549 (N_11549,N_11245,N_11314);
and U11550 (N_11550,N_11335,N_11262);
and U11551 (N_11551,N_11204,N_11341);
or U11552 (N_11552,N_11304,N_11376);
or U11553 (N_11553,N_11377,N_11251);
nor U11554 (N_11554,N_11206,N_11200);
and U11555 (N_11555,N_11394,N_11310);
and U11556 (N_11556,N_11340,N_11335);
and U11557 (N_11557,N_11260,N_11277);
nor U11558 (N_11558,N_11306,N_11232);
or U11559 (N_11559,N_11260,N_11379);
nor U11560 (N_11560,N_11361,N_11209);
nand U11561 (N_11561,N_11328,N_11363);
and U11562 (N_11562,N_11396,N_11231);
nand U11563 (N_11563,N_11239,N_11220);
and U11564 (N_11564,N_11386,N_11330);
nand U11565 (N_11565,N_11213,N_11291);
or U11566 (N_11566,N_11271,N_11269);
nand U11567 (N_11567,N_11234,N_11318);
and U11568 (N_11568,N_11366,N_11293);
and U11569 (N_11569,N_11256,N_11354);
or U11570 (N_11570,N_11234,N_11289);
nand U11571 (N_11571,N_11332,N_11314);
nand U11572 (N_11572,N_11200,N_11387);
nor U11573 (N_11573,N_11220,N_11218);
nor U11574 (N_11574,N_11363,N_11246);
and U11575 (N_11575,N_11282,N_11372);
and U11576 (N_11576,N_11259,N_11322);
nand U11577 (N_11577,N_11284,N_11336);
nand U11578 (N_11578,N_11354,N_11326);
nor U11579 (N_11579,N_11213,N_11257);
or U11580 (N_11580,N_11314,N_11274);
or U11581 (N_11581,N_11281,N_11309);
and U11582 (N_11582,N_11302,N_11234);
nor U11583 (N_11583,N_11322,N_11302);
xnor U11584 (N_11584,N_11372,N_11394);
xor U11585 (N_11585,N_11233,N_11202);
nor U11586 (N_11586,N_11346,N_11339);
nand U11587 (N_11587,N_11250,N_11260);
nand U11588 (N_11588,N_11284,N_11227);
and U11589 (N_11589,N_11290,N_11371);
and U11590 (N_11590,N_11254,N_11303);
nand U11591 (N_11591,N_11379,N_11240);
and U11592 (N_11592,N_11354,N_11226);
nor U11593 (N_11593,N_11292,N_11274);
and U11594 (N_11594,N_11374,N_11288);
xnor U11595 (N_11595,N_11372,N_11246);
xnor U11596 (N_11596,N_11327,N_11350);
nor U11597 (N_11597,N_11278,N_11320);
or U11598 (N_11598,N_11335,N_11303);
nor U11599 (N_11599,N_11380,N_11288);
nor U11600 (N_11600,N_11527,N_11422);
and U11601 (N_11601,N_11562,N_11403);
nor U11602 (N_11602,N_11560,N_11592);
nand U11603 (N_11603,N_11449,N_11453);
xor U11604 (N_11604,N_11400,N_11471);
nor U11605 (N_11605,N_11524,N_11401);
and U11606 (N_11606,N_11547,N_11561);
or U11607 (N_11607,N_11454,N_11450);
or U11608 (N_11608,N_11540,N_11529);
and U11609 (N_11609,N_11525,N_11459);
or U11610 (N_11610,N_11416,N_11576);
nor U11611 (N_11611,N_11478,N_11485);
and U11612 (N_11612,N_11555,N_11439);
nor U11613 (N_11613,N_11499,N_11544);
nand U11614 (N_11614,N_11519,N_11408);
and U11615 (N_11615,N_11533,N_11427);
and U11616 (N_11616,N_11558,N_11426);
nand U11617 (N_11617,N_11553,N_11411);
or U11618 (N_11618,N_11467,N_11438);
xor U11619 (N_11619,N_11483,N_11535);
or U11620 (N_11620,N_11473,N_11462);
xnor U11621 (N_11621,N_11491,N_11490);
nor U11622 (N_11622,N_11404,N_11494);
nor U11623 (N_11623,N_11460,N_11418);
xnor U11624 (N_11624,N_11407,N_11442);
or U11625 (N_11625,N_11406,N_11586);
nand U11626 (N_11626,N_11534,N_11564);
and U11627 (N_11627,N_11474,N_11433);
and U11628 (N_11628,N_11549,N_11530);
and U11629 (N_11629,N_11476,N_11573);
xor U11630 (N_11630,N_11511,N_11580);
nor U11631 (N_11631,N_11466,N_11456);
nand U11632 (N_11632,N_11415,N_11516);
or U11633 (N_11633,N_11568,N_11579);
nand U11634 (N_11634,N_11598,N_11597);
nand U11635 (N_11635,N_11548,N_11566);
and U11636 (N_11636,N_11497,N_11585);
or U11637 (N_11637,N_11463,N_11507);
nor U11638 (N_11638,N_11414,N_11596);
xor U11639 (N_11639,N_11412,N_11495);
or U11640 (N_11640,N_11417,N_11437);
nor U11641 (N_11641,N_11569,N_11577);
nand U11642 (N_11642,N_11531,N_11588);
nor U11643 (N_11643,N_11594,N_11452);
or U11644 (N_11644,N_11526,N_11424);
or U11645 (N_11645,N_11436,N_11582);
nor U11646 (N_11646,N_11480,N_11444);
or U11647 (N_11647,N_11479,N_11559);
nor U11648 (N_11648,N_11468,N_11539);
nor U11649 (N_11649,N_11506,N_11419);
nand U11650 (N_11650,N_11570,N_11420);
nand U11651 (N_11651,N_11554,N_11441);
nor U11652 (N_11652,N_11574,N_11445);
xnor U11653 (N_11653,N_11477,N_11593);
or U11654 (N_11654,N_11472,N_11551);
and U11655 (N_11655,N_11521,N_11509);
xor U11656 (N_11656,N_11517,N_11546);
nand U11657 (N_11657,N_11440,N_11410);
or U11658 (N_11658,N_11556,N_11402);
or U11659 (N_11659,N_11518,N_11487);
or U11660 (N_11660,N_11435,N_11508);
nand U11661 (N_11661,N_11421,N_11470);
or U11662 (N_11662,N_11489,N_11457);
and U11663 (N_11663,N_11541,N_11475);
or U11664 (N_11664,N_11505,N_11557);
nand U11665 (N_11665,N_11434,N_11552);
nand U11666 (N_11666,N_11584,N_11514);
and U11667 (N_11667,N_11581,N_11448);
or U11668 (N_11668,N_11500,N_11563);
nor U11669 (N_11669,N_11578,N_11432);
xor U11670 (N_11670,N_11536,N_11504);
nor U11671 (N_11671,N_11591,N_11486);
nor U11672 (N_11672,N_11455,N_11513);
nand U11673 (N_11673,N_11496,N_11590);
nand U11674 (N_11674,N_11575,N_11589);
nand U11675 (N_11675,N_11522,N_11595);
or U11676 (N_11676,N_11482,N_11484);
nor U11677 (N_11677,N_11431,N_11587);
nor U11678 (N_11678,N_11565,N_11572);
xnor U11679 (N_11679,N_11501,N_11430);
nand U11680 (N_11680,N_11537,N_11515);
nand U11681 (N_11681,N_11423,N_11461);
nand U11682 (N_11682,N_11443,N_11523);
or U11683 (N_11683,N_11458,N_11545);
or U11684 (N_11684,N_11583,N_11571);
and U11685 (N_11685,N_11429,N_11512);
nand U11686 (N_11686,N_11503,N_11510);
nor U11687 (N_11687,N_11550,N_11599);
nand U11688 (N_11688,N_11447,N_11481);
nor U11689 (N_11689,N_11567,N_11465);
and U11690 (N_11690,N_11528,N_11538);
and U11691 (N_11691,N_11520,N_11498);
xor U11692 (N_11692,N_11543,N_11469);
nor U11693 (N_11693,N_11493,N_11492);
or U11694 (N_11694,N_11425,N_11446);
and U11695 (N_11695,N_11451,N_11405);
nand U11696 (N_11696,N_11409,N_11413);
nor U11697 (N_11697,N_11532,N_11502);
nand U11698 (N_11698,N_11464,N_11428);
nor U11699 (N_11699,N_11488,N_11542);
and U11700 (N_11700,N_11584,N_11544);
xnor U11701 (N_11701,N_11581,N_11403);
xor U11702 (N_11702,N_11503,N_11573);
nand U11703 (N_11703,N_11457,N_11428);
and U11704 (N_11704,N_11576,N_11464);
nand U11705 (N_11705,N_11493,N_11561);
nand U11706 (N_11706,N_11460,N_11472);
nand U11707 (N_11707,N_11537,N_11555);
or U11708 (N_11708,N_11533,N_11501);
or U11709 (N_11709,N_11494,N_11469);
and U11710 (N_11710,N_11564,N_11500);
and U11711 (N_11711,N_11506,N_11466);
or U11712 (N_11712,N_11569,N_11534);
or U11713 (N_11713,N_11497,N_11535);
and U11714 (N_11714,N_11570,N_11531);
or U11715 (N_11715,N_11479,N_11587);
nor U11716 (N_11716,N_11590,N_11501);
nor U11717 (N_11717,N_11493,N_11448);
and U11718 (N_11718,N_11572,N_11540);
nor U11719 (N_11719,N_11590,N_11463);
nand U11720 (N_11720,N_11452,N_11479);
nor U11721 (N_11721,N_11429,N_11547);
nor U11722 (N_11722,N_11516,N_11560);
and U11723 (N_11723,N_11531,N_11445);
and U11724 (N_11724,N_11408,N_11510);
nor U11725 (N_11725,N_11523,N_11474);
nand U11726 (N_11726,N_11419,N_11594);
nand U11727 (N_11727,N_11579,N_11557);
xnor U11728 (N_11728,N_11418,N_11511);
nand U11729 (N_11729,N_11492,N_11407);
and U11730 (N_11730,N_11501,N_11542);
and U11731 (N_11731,N_11488,N_11411);
and U11732 (N_11732,N_11596,N_11529);
and U11733 (N_11733,N_11575,N_11569);
or U11734 (N_11734,N_11490,N_11489);
nor U11735 (N_11735,N_11422,N_11473);
nand U11736 (N_11736,N_11480,N_11572);
and U11737 (N_11737,N_11498,N_11556);
nand U11738 (N_11738,N_11519,N_11486);
and U11739 (N_11739,N_11521,N_11466);
nand U11740 (N_11740,N_11456,N_11408);
nand U11741 (N_11741,N_11540,N_11545);
nor U11742 (N_11742,N_11493,N_11569);
nor U11743 (N_11743,N_11552,N_11489);
or U11744 (N_11744,N_11511,N_11415);
nand U11745 (N_11745,N_11489,N_11402);
or U11746 (N_11746,N_11525,N_11552);
xnor U11747 (N_11747,N_11550,N_11488);
nand U11748 (N_11748,N_11423,N_11402);
and U11749 (N_11749,N_11493,N_11571);
or U11750 (N_11750,N_11551,N_11542);
nand U11751 (N_11751,N_11466,N_11519);
nor U11752 (N_11752,N_11591,N_11593);
or U11753 (N_11753,N_11557,N_11498);
nand U11754 (N_11754,N_11464,N_11424);
nand U11755 (N_11755,N_11576,N_11584);
or U11756 (N_11756,N_11438,N_11585);
nor U11757 (N_11757,N_11541,N_11498);
nand U11758 (N_11758,N_11524,N_11443);
and U11759 (N_11759,N_11592,N_11563);
nor U11760 (N_11760,N_11512,N_11463);
nand U11761 (N_11761,N_11473,N_11493);
or U11762 (N_11762,N_11552,N_11463);
nand U11763 (N_11763,N_11468,N_11491);
and U11764 (N_11764,N_11431,N_11451);
or U11765 (N_11765,N_11486,N_11427);
and U11766 (N_11766,N_11562,N_11434);
nand U11767 (N_11767,N_11439,N_11438);
nor U11768 (N_11768,N_11500,N_11411);
or U11769 (N_11769,N_11495,N_11478);
and U11770 (N_11770,N_11420,N_11571);
nor U11771 (N_11771,N_11597,N_11541);
or U11772 (N_11772,N_11439,N_11572);
nor U11773 (N_11773,N_11453,N_11447);
or U11774 (N_11774,N_11478,N_11584);
nand U11775 (N_11775,N_11520,N_11526);
nand U11776 (N_11776,N_11407,N_11494);
nor U11777 (N_11777,N_11418,N_11512);
or U11778 (N_11778,N_11487,N_11434);
and U11779 (N_11779,N_11431,N_11516);
and U11780 (N_11780,N_11589,N_11462);
or U11781 (N_11781,N_11442,N_11570);
xnor U11782 (N_11782,N_11441,N_11476);
nand U11783 (N_11783,N_11484,N_11452);
and U11784 (N_11784,N_11467,N_11522);
nand U11785 (N_11785,N_11405,N_11431);
and U11786 (N_11786,N_11497,N_11495);
nor U11787 (N_11787,N_11475,N_11574);
and U11788 (N_11788,N_11406,N_11515);
nor U11789 (N_11789,N_11447,N_11442);
nor U11790 (N_11790,N_11515,N_11452);
xnor U11791 (N_11791,N_11409,N_11412);
and U11792 (N_11792,N_11531,N_11452);
nor U11793 (N_11793,N_11442,N_11449);
nor U11794 (N_11794,N_11513,N_11543);
and U11795 (N_11795,N_11463,N_11541);
and U11796 (N_11796,N_11434,N_11477);
and U11797 (N_11797,N_11475,N_11571);
xor U11798 (N_11798,N_11568,N_11576);
nor U11799 (N_11799,N_11489,N_11430);
nor U11800 (N_11800,N_11663,N_11623);
and U11801 (N_11801,N_11717,N_11744);
nand U11802 (N_11802,N_11657,N_11654);
nor U11803 (N_11803,N_11601,N_11671);
nand U11804 (N_11804,N_11768,N_11765);
or U11805 (N_11805,N_11763,N_11600);
xor U11806 (N_11806,N_11707,N_11726);
nand U11807 (N_11807,N_11751,N_11645);
or U11808 (N_11808,N_11697,N_11652);
or U11809 (N_11809,N_11708,N_11703);
nor U11810 (N_11810,N_11670,N_11784);
and U11811 (N_11811,N_11612,N_11642);
or U11812 (N_11812,N_11653,N_11626);
nand U11813 (N_11813,N_11676,N_11710);
or U11814 (N_11814,N_11790,N_11699);
nor U11815 (N_11815,N_11683,N_11721);
nand U11816 (N_11816,N_11621,N_11741);
or U11817 (N_11817,N_11732,N_11687);
nand U11818 (N_11818,N_11791,N_11675);
xnor U11819 (N_11819,N_11793,N_11633);
xnor U11820 (N_11820,N_11735,N_11605);
or U11821 (N_11821,N_11616,N_11719);
nor U11822 (N_11822,N_11713,N_11760);
nand U11823 (N_11823,N_11783,N_11720);
nand U11824 (N_11824,N_11706,N_11775);
or U11825 (N_11825,N_11694,N_11648);
nor U11826 (N_11826,N_11607,N_11702);
nand U11827 (N_11827,N_11769,N_11754);
or U11828 (N_11828,N_11677,N_11602);
nor U11829 (N_11829,N_11746,N_11682);
nand U11830 (N_11830,N_11636,N_11611);
nor U11831 (N_11831,N_11739,N_11684);
or U11832 (N_11832,N_11701,N_11651);
or U11833 (N_11833,N_11729,N_11704);
or U11834 (N_11834,N_11705,N_11680);
or U11835 (N_11835,N_11620,N_11716);
nor U11836 (N_11836,N_11692,N_11777);
nor U11837 (N_11837,N_11672,N_11617);
or U11838 (N_11838,N_11722,N_11691);
nor U11839 (N_11839,N_11650,N_11641);
or U11840 (N_11840,N_11622,N_11759);
nor U11841 (N_11841,N_11627,N_11731);
nand U11842 (N_11842,N_11625,N_11678);
or U11843 (N_11843,N_11757,N_11718);
or U11844 (N_11844,N_11660,N_11798);
nor U11845 (N_11845,N_11655,N_11635);
or U11846 (N_11846,N_11733,N_11690);
nand U11847 (N_11847,N_11662,N_11770);
xnor U11848 (N_11848,N_11795,N_11630);
nand U11849 (N_11849,N_11646,N_11725);
and U11850 (N_11850,N_11679,N_11778);
xor U11851 (N_11851,N_11738,N_11797);
nand U11852 (N_11852,N_11737,N_11724);
nor U11853 (N_11853,N_11644,N_11714);
nor U11854 (N_11854,N_11674,N_11748);
nand U11855 (N_11855,N_11698,N_11693);
nand U11856 (N_11856,N_11764,N_11668);
nand U11857 (N_11857,N_11734,N_11700);
nor U11858 (N_11858,N_11758,N_11643);
and U11859 (N_11859,N_11673,N_11709);
or U11860 (N_11860,N_11728,N_11661);
nor U11861 (N_11861,N_11615,N_11624);
nand U11862 (N_11862,N_11613,N_11799);
and U11863 (N_11863,N_11781,N_11666);
nand U11864 (N_11864,N_11740,N_11730);
nor U11865 (N_11865,N_11785,N_11685);
nor U11866 (N_11866,N_11727,N_11776);
xor U11867 (N_11867,N_11736,N_11796);
or U11868 (N_11868,N_11632,N_11792);
nand U11869 (N_11869,N_11743,N_11665);
nor U11870 (N_11870,N_11686,N_11639);
and U11871 (N_11871,N_11656,N_11649);
nand U11872 (N_11872,N_11745,N_11695);
or U11873 (N_11873,N_11782,N_11640);
and U11874 (N_11874,N_11774,N_11773);
or U11875 (N_11875,N_11609,N_11762);
and U11876 (N_11876,N_11788,N_11742);
and U11877 (N_11877,N_11767,N_11638);
nor U11878 (N_11878,N_11628,N_11772);
nor U11879 (N_11879,N_11787,N_11634);
xor U11880 (N_11880,N_11711,N_11780);
and U11881 (N_11881,N_11669,N_11752);
or U11882 (N_11882,N_11618,N_11658);
nand U11883 (N_11883,N_11610,N_11603);
nor U11884 (N_11884,N_11712,N_11794);
nor U11885 (N_11885,N_11766,N_11659);
nand U11886 (N_11886,N_11681,N_11779);
nor U11887 (N_11887,N_11664,N_11786);
nor U11888 (N_11888,N_11606,N_11614);
and U11889 (N_11889,N_11629,N_11696);
or U11890 (N_11890,N_11723,N_11631);
and U11891 (N_11891,N_11647,N_11608);
and U11892 (N_11892,N_11688,N_11619);
or U11893 (N_11893,N_11755,N_11747);
nand U11894 (N_11894,N_11749,N_11750);
nand U11895 (N_11895,N_11771,N_11761);
nand U11896 (N_11896,N_11689,N_11604);
and U11897 (N_11897,N_11637,N_11756);
or U11898 (N_11898,N_11753,N_11715);
xnor U11899 (N_11899,N_11667,N_11789);
or U11900 (N_11900,N_11633,N_11670);
nor U11901 (N_11901,N_11658,N_11779);
and U11902 (N_11902,N_11789,N_11649);
and U11903 (N_11903,N_11647,N_11668);
nand U11904 (N_11904,N_11649,N_11760);
nand U11905 (N_11905,N_11611,N_11650);
or U11906 (N_11906,N_11702,N_11635);
and U11907 (N_11907,N_11767,N_11745);
xnor U11908 (N_11908,N_11758,N_11652);
nor U11909 (N_11909,N_11786,N_11605);
and U11910 (N_11910,N_11655,N_11794);
nand U11911 (N_11911,N_11640,N_11763);
and U11912 (N_11912,N_11673,N_11681);
nor U11913 (N_11913,N_11650,N_11796);
nor U11914 (N_11914,N_11723,N_11681);
nand U11915 (N_11915,N_11670,N_11720);
nand U11916 (N_11916,N_11775,N_11748);
or U11917 (N_11917,N_11605,N_11741);
and U11918 (N_11918,N_11771,N_11753);
or U11919 (N_11919,N_11627,N_11682);
nand U11920 (N_11920,N_11611,N_11614);
nand U11921 (N_11921,N_11615,N_11758);
nor U11922 (N_11922,N_11641,N_11753);
nand U11923 (N_11923,N_11683,N_11739);
or U11924 (N_11924,N_11795,N_11733);
nor U11925 (N_11925,N_11755,N_11691);
or U11926 (N_11926,N_11628,N_11662);
nor U11927 (N_11927,N_11700,N_11723);
or U11928 (N_11928,N_11623,N_11716);
and U11929 (N_11929,N_11707,N_11712);
and U11930 (N_11930,N_11774,N_11676);
nor U11931 (N_11931,N_11616,N_11669);
nand U11932 (N_11932,N_11728,N_11696);
xnor U11933 (N_11933,N_11731,N_11719);
nand U11934 (N_11934,N_11696,N_11699);
nor U11935 (N_11935,N_11686,N_11663);
nand U11936 (N_11936,N_11752,N_11716);
or U11937 (N_11937,N_11726,N_11675);
nor U11938 (N_11938,N_11626,N_11663);
or U11939 (N_11939,N_11696,N_11602);
nand U11940 (N_11940,N_11702,N_11748);
nor U11941 (N_11941,N_11610,N_11617);
or U11942 (N_11942,N_11637,N_11618);
nand U11943 (N_11943,N_11608,N_11742);
or U11944 (N_11944,N_11609,N_11623);
or U11945 (N_11945,N_11738,N_11758);
nand U11946 (N_11946,N_11796,N_11640);
nand U11947 (N_11947,N_11651,N_11687);
nor U11948 (N_11948,N_11652,N_11628);
or U11949 (N_11949,N_11603,N_11704);
nand U11950 (N_11950,N_11742,N_11789);
nand U11951 (N_11951,N_11732,N_11781);
nor U11952 (N_11952,N_11773,N_11799);
and U11953 (N_11953,N_11740,N_11612);
or U11954 (N_11954,N_11606,N_11723);
and U11955 (N_11955,N_11655,N_11734);
xnor U11956 (N_11956,N_11661,N_11713);
nand U11957 (N_11957,N_11641,N_11788);
nor U11958 (N_11958,N_11705,N_11611);
and U11959 (N_11959,N_11769,N_11602);
or U11960 (N_11960,N_11668,N_11690);
nor U11961 (N_11961,N_11778,N_11727);
nor U11962 (N_11962,N_11737,N_11759);
nand U11963 (N_11963,N_11734,N_11616);
and U11964 (N_11964,N_11711,N_11648);
or U11965 (N_11965,N_11796,N_11601);
nor U11966 (N_11966,N_11744,N_11769);
nand U11967 (N_11967,N_11768,N_11602);
nor U11968 (N_11968,N_11632,N_11774);
nand U11969 (N_11969,N_11607,N_11650);
nor U11970 (N_11970,N_11655,N_11699);
nand U11971 (N_11971,N_11788,N_11790);
or U11972 (N_11972,N_11789,N_11733);
and U11973 (N_11973,N_11694,N_11631);
nor U11974 (N_11974,N_11711,N_11650);
nor U11975 (N_11975,N_11706,N_11621);
nand U11976 (N_11976,N_11686,N_11731);
and U11977 (N_11977,N_11679,N_11626);
nand U11978 (N_11978,N_11639,N_11754);
or U11979 (N_11979,N_11621,N_11724);
nor U11980 (N_11980,N_11644,N_11676);
or U11981 (N_11981,N_11747,N_11667);
nand U11982 (N_11982,N_11668,N_11741);
xor U11983 (N_11983,N_11791,N_11676);
and U11984 (N_11984,N_11732,N_11663);
nand U11985 (N_11985,N_11662,N_11778);
nand U11986 (N_11986,N_11793,N_11682);
nor U11987 (N_11987,N_11628,N_11749);
and U11988 (N_11988,N_11783,N_11609);
and U11989 (N_11989,N_11612,N_11735);
nor U11990 (N_11990,N_11624,N_11616);
nand U11991 (N_11991,N_11717,N_11657);
and U11992 (N_11992,N_11661,N_11779);
nand U11993 (N_11993,N_11664,N_11793);
nand U11994 (N_11994,N_11720,N_11633);
and U11995 (N_11995,N_11698,N_11766);
or U11996 (N_11996,N_11739,N_11666);
or U11997 (N_11997,N_11653,N_11760);
or U11998 (N_11998,N_11606,N_11625);
nand U11999 (N_11999,N_11654,N_11772);
or U12000 (N_12000,N_11991,N_11947);
and U12001 (N_12001,N_11904,N_11956);
nor U12002 (N_12002,N_11847,N_11915);
and U12003 (N_12003,N_11872,N_11914);
nor U12004 (N_12004,N_11878,N_11884);
nor U12005 (N_12005,N_11963,N_11845);
xnor U12006 (N_12006,N_11870,N_11826);
nor U12007 (N_12007,N_11889,N_11842);
nor U12008 (N_12008,N_11906,N_11873);
nor U12009 (N_12009,N_11919,N_11824);
or U12010 (N_12010,N_11863,N_11858);
or U12011 (N_12011,N_11905,N_11818);
xnor U12012 (N_12012,N_11838,N_11867);
nor U12013 (N_12013,N_11973,N_11950);
nand U12014 (N_12014,N_11933,N_11971);
and U12015 (N_12015,N_11869,N_11948);
or U12016 (N_12016,N_11806,N_11935);
nand U12017 (N_12017,N_11939,N_11891);
and U12018 (N_12018,N_11982,N_11892);
nor U12019 (N_12019,N_11890,N_11999);
and U12020 (N_12020,N_11940,N_11898);
xor U12021 (N_12021,N_11822,N_11909);
or U12022 (N_12022,N_11900,N_11804);
nand U12023 (N_12023,N_11981,N_11849);
or U12024 (N_12024,N_11925,N_11916);
nor U12025 (N_12025,N_11841,N_11880);
and U12026 (N_12026,N_11876,N_11848);
and U12027 (N_12027,N_11859,N_11882);
nand U12028 (N_12028,N_11951,N_11812);
and U12029 (N_12029,N_11929,N_11819);
nor U12030 (N_12030,N_11985,N_11946);
and U12031 (N_12031,N_11801,N_11907);
nand U12032 (N_12032,N_11836,N_11886);
nor U12033 (N_12033,N_11928,N_11839);
nand U12034 (N_12034,N_11988,N_11958);
and U12035 (N_12035,N_11962,N_11883);
xnor U12036 (N_12036,N_11972,N_11930);
nand U12037 (N_12037,N_11866,N_11918);
nand U12038 (N_12038,N_11885,N_11923);
and U12039 (N_12039,N_11984,N_11854);
xor U12040 (N_12040,N_11857,N_11899);
nor U12041 (N_12041,N_11980,N_11881);
and U12042 (N_12042,N_11827,N_11910);
xnor U12043 (N_12043,N_11830,N_11911);
or U12044 (N_12044,N_11860,N_11871);
nand U12045 (N_12045,N_11993,N_11868);
and U12046 (N_12046,N_11913,N_11957);
xnor U12047 (N_12047,N_11896,N_11995);
or U12048 (N_12048,N_11851,N_11924);
or U12049 (N_12049,N_11989,N_11979);
or U12050 (N_12050,N_11877,N_11810);
and U12051 (N_12051,N_11862,N_11887);
or U12052 (N_12052,N_11879,N_11986);
or U12053 (N_12053,N_11959,N_11941);
and U12054 (N_12054,N_11825,N_11844);
nor U12055 (N_12055,N_11966,N_11893);
and U12056 (N_12056,N_11996,N_11920);
or U12057 (N_12057,N_11931,N_11977);
or U12058 (N_12058,N_11921,N_11908);
nor U12059 (N_12059,N_11821,N_11955);
or U12060 (N_12060,N_11994,N_11846);
or U12061 (N_12061,N_11865,N_11843);
nand U12062 (N_12062,N_11856,N_11897);
and U12063 (N_12063,N_11937,N_11820);
and U12064 (N_12064,N_11945,N_11990);
nand U12065 (N_12065,N_11805,N_11901);
nand U12066 (N_12066,N_11927,N_11954);
nand U12067 (N_12067,N_11975,N_11834);
nor U12068 (N_12068,N_11936,N_11864);
or U12069 (N_12069,N_11942,N_11850);
nor U12070 (N_12070,N_11894,N_11852);
nand U12071 (N_12071,N_11817,N_11875);
nor U12072 (N_12072,N_11938,N_11813);
and U12073 (N_12073,N_11987,N_11902);
or U12074 (N_12074,N_11803,N_11926);
or U12075 (N_12075,N_11960,N_11802);
or U12076 (N_12076,N_11814,N_11823);
nand U12077 (N_12077,N_11829,N_11998);
or U12078 (N_12078,N_11983,N_11964);
nor U12079 (N_12079,N_11961,N_11932);
nor U12080 (N_12080,N_11944,N_11800);
or U12081 (N_12081,N_11968,N_11974);
nor U12082 (N_12082,N_11828,N_11815);
nor U12083 (N_12083,N_11969,N_11903);
or U12084 (N_12084,N_11917,N_11807);
and U12085 (N_12085,N_11953,N_11853);
nor U12086 (N_12086,N_11997,N_11970);
or U12087 (N_12087,N_11808,N_11835);
nor U12088 (N_12088,N_11831,N_11943);
and U12089 (N_12089,N_11976,N_11832);
or U12090 (N_12090,N_11816,N_11861);
or U12091 (N_12091,N_11837,N_11895);
nand U12092 (N_12092,N_11949,N_11811);
and U12093 (N_12093,N_11855,N_11874);
or U12094 (N_12094,N_11840,N_11809);
nor U12095 (N_12095,N_11888,N_11912);
nor U12096 (N_12096,N_11965,N_11978);
or U12097 (N_12097,N_11934,N_11967);
and U12098 (N_12098,N_11952,N_11922);
and U12099 (N_12099,N_11833,N_11992);
and U12100 (N_12100,N_11803,N_11813);
nand U12101 (N_12101,N_11892,N_11817);
or U12102 (N_12102,N_11977,N_11820);
and U12103 (N_12103,N_11917,N_11847);
nand U12104 (N_12104,N_11899,N_11938);
nand U12105 (N_12105,N_11997,N_11824);
nor U12106 (N_12106,N_11960,N_11948);
and U12107 (N_12107,N_11925,N_11942);
nand U12108 (N_12108,N_11861,N_11933);
and U12109 (N_12109,N_11931,N_11983);
nor U12110 (N_12110,N_11946,N_11876);
xnor U12111 (N_12111,N_11810,N_11868);
and U12112 (N_12112,N_11976,N_11908);
nand U12113 (N_12113,N_11940,N_11999);
nand U12114 (N_12114,N_11862,N_11816);
and U12115 (N_12115,N_11868,N_11892);
nor U12116 (N_12116,N_11949,N_11899);
nor U12117 (N_12117,N_11951,N_11987);
nand U12118 (N_12118,N_11911,N_11984);
and U12119 (N_12119,N_11951,N_11999);
nand U12120 (N_12120,N_11967,N_11959);
nand U12121 (N_12121,N_11882,N_11941);
nor U12122 (N_12122,N_11906,N_11834);
and U12123 (N_12123,N_11931,N_11803);
and U12124 (N_12124,N_11956,N_11962);
and U12125 (N_12125,N_11885,N_11924);
nor U12126 (N_12126,N_11920,N_11835);
nand U12127 (N_12127,N_11859,N_11956);
nor U12128 (N_12128,N_11854,N_11806);
nor U12129 (N_12129,N_11905,N_11902);
or U12130 (N_12130,N_11955,N_11908);
and U12131 (N_12131,N_11987,N_11942);
or U12132 (N_12132,N_11942,N_11926);
or U12133 (N_12133,N_11834,N_11859);
and U12134 (N_12134,N_11820,N_11982);
and U12135 (N_12135,N_11803,N_11872);
and U12136 (N_12136,N_11973,N_11970);
nand U12137 (N_12137,N_11920,N_11917);
and U12138 (N_12138,N_11872,N_11860);
or U12139 (N_12139,N_11826,N_11828);
or U12140 (N_12140,N_11927,N_11926);
nand U12141 (N_12141,N_11819,N_11909);
nor U12142 (N_12142,N_11801,N_11979);
nor U12143 (N_12143,N_11856,N_11830);
and U12144 (N_12144,N_11950,N_11841);
and U12145 (N_12145,N_11861,N_11994);
or U12146 (N_12146,N_11990,N_11804);
and U12147 (N_12147,N_11940,N_11951);
or U12148 (N_12148,N_11982,N_11833);
nand U12149 (N_12149,N_11991,N_11920);
and U12150 (N_12150,N_11848,N_11917);
nor U12151 (N_12151,N_11826,N_11978);
xor U12152 (N_12152,N_11879,N_11832);
nor U12153 (N_12153,N_11975,N_11980);
nand U12154 (N_12154,N_11910,N_11915);
and U12155 (N_12155,N_11905,N_11839);
and U12156 (N_12156,N_11872,N_11806);
and U12157 (N_12157,N_11878,N_11845);
nor U12158 (N_12158,N_11865,N_11820);
and U12159 (N_12159,N_11993,N_11803);
nand U12160 (N_12160,N_11916,N_11868);
and U12161 (N_12161,N_11809,N_11914);
and U12162 (N_12162,N_11926,N_11869);
xor U12163 (N_12163,N_11968,N_11814);
nand U12164 (N_12164,N_11921,N_11811);
nor U12165 (N_12165,N_11888,N_11808);
nand U12166 (N_12166,N_11889,N_11858);
or U12167 (N_12167,N_11956,N_11908);
nand U12168 (N_12168,N_11812,N_11819);
and U12169 (N_12169,N_11940,N_11942);
or U12170 (N_12170,N_11948,N_11892);
or U12171 (N_12171,N_11947,N_11882);
and U12172 (N_12172,N_11889,N_11860);
and U12173 (N_12173,N_11991,N_11805);
xnor U12174 (N_12174,N_11922,N_11854);
xnor U12175 (N_12175,N_11844,N_11938);
nand U12176 (N_12176,N_11978,N_11979);
or U12177 (N_12177,N_11816,N_11904);
or U12178 (N_12178,N_11947,N_11941);
and U12179 (N_12179,N_11944,N_11872);
and U12180 (N_12180,N_11895,N_11940);
and U12181 (N_12181,N_11827,N_11966);
nor U12182 (N_12182,N_11936,N_11926);
nor U12183 (N_12183,N_11889,N_11947);
nor U12184 (N_12184,N_11972,N_11978);
nor U12185 (N_12185,N_11838,N_11969);
or U12186 (N_12186,N_11940,N_11968);
xnor U12187 (N_12187,N_11914,N_11856);
nor U12188 (N_12188,N_11821,N_11944);
and U12189 (N_12189,N_11922,N_11800);
and U12190 (N_12190,N_11939,N_11825);
nor U12191 (N_12191,N_11856,N_11809);
or U12192 (N_12192,N_11986,N_11935);
and U12193 (N_12193,N_11901,N_11957);
and U12194 (N_12194,N_11880,N_11931);
nand U12195 (N_12195,N_11951,N_11880);
or U12196 (N_12196,N_11896,N_11809);
or U12197 (N_12197,N_11843,N_11940);
nand U12198 (N_12198,N_11901,N_11909);
or U12199 (N_12199,N_11966,N_11873);
or U12200 (N_12200,N_12082,N_12050);
nand U12201 (N_12201,N_12101,N_12197);
nor U12202 (N_12202,N_12019,N_12027);
and U12203 (N_12203,N_12161,N_12017);
or U12204 (N_12204,N_12004,N_12039);
and U12205 (N_12205,N_12041,N_12015);
or U12206 (N_12206,N_12046,N_12144);
or U12207 (N_12207,N_12010,N_12185);
and U12208 (N_12208,N_12131,N_12178);
and U12209 (N_12209,N_12100,N_12164);
or U12210 (N_12210,N_12024,N_12135);
nor U12211 (N_12211,N_12180,N_12083);
nand U12212 (N_12212,N_12189,N_12081);
and U12213 (N_12213,N_12124,N_12057);
nor U12214 (N_12214,N_12110,N_12145);
or U12215 (N_12215,N_12003,N_12097);
nand U12216 (N_12216,N_12078,N_12018);
nand U12217 (N_12217,N_12179,N_12045);
xnor U12218 (N_12218,N_12030,N_12187);
nand U12219 (N_12219,N_12048,N_12064);
and U12220 (N_12220,N_12021,N_12198);
nor U12221 (N_12221,N_12159,N_12062);
or U12222 (N_12222,N_12075,N_12183);
xnor U12223 (N_12223,N_12169,N_12121);
nand U12224 (N_12224,N_12166,N_12001);
and U12225 (N_12225,N_12089,N_12091);
and U12226 (N_12226,N_12170,N_12171);
nand U12227 (N_12227,N_12053,N_12199);
nor U12228 (N_12228,N_12026,N_12037);
nand U12229 (N_12229,N_12051,N_12073);
or U12230 (N_12230,N_12005,N_12065);
and U12231 (N_12231,N_12142,N_12040);
nor U12232 (N_12232,N_12134,N_12071);
nand U12233 (N_12233,N_12147,N_12123);
nand U12234 (N_12234,N_12196,N_12036);
nor U12235 (N_12235,N_12141,N_12028);
nand U12236 (N_12236,N_12140,N_12193);
xnor U12237 (N_12237,N_12116,N_12129);
nand U12238 (N_12238,N_12059,N_12072);
or U12239 (N_12239,N_12126,N_12025);
nand U12240 (N_12240,N_12150,N_12022);
nor U12241 (N_12241,N_12084,N_12168);
or U12242 (N_12242,N_12099,N_12054);
nand U12243 (N_12243,N_12137,N_12176);
nor U12244 (N_12244,N_12095,N_12151);
or U12245 (N_12245,N_12104,N_12108);
xor U12246 (N_12246,N_12103,N_12080);
and U12247 (N_12247,N_12006,N_12152);
xnor U12248 (N_12248,N_12098,N_12011);
or U12249 (N_12249,N_12014,N_12031);
nand U12250 (N_12250,N_12192,N_12013);
nand U12251 (N_12251,N_12069,N_12138);
or U12252 (N_12252,N_12077,N_12125);
nor U12253 (N_12253,N_12132,N_12186);
xor U12254 (N_12254,N_12154,N_12191);
or U12255 (N_12255,N_12092,N_12130);
and U12256 (N_12256,N_12023,N_12063);
or U12257 (N_12257,N_12087,N_12115);
nor U12258 (N_12258,N_12167,N_12085);
nand U12259 (N_12259,N_12032,N_12000);
or U12260 (N_12260,N_12143,N_12184);
nor U12261 (N_12261,N_12181,N_12086);
nand U12262 (N_12262,N_12034,N_12160);
and U12263 (N_12263,N_12060,N_12066);
nand U12264 (N_12264,N_12173,N_12044);
nor U12265 (N_12265,N_12002,N_12043);
nand U12266 (N_12266,N_12007,N_12111);
and U12267 (N_12267,N_12029,N_12153);
nand U12268 (N_12268,N_12118,N_12107);
nor U12269 (N_12269,N_12148,N_12052);
nand U12270 (N_12270,N_12033,N_12035);
xor U12271 (N_12271,N_12068,N_12106);
and U12272 (N_12272,N_12113,N_12093);
nor U12273 (N_12273,N_12061,N_12076);
nor U12274 (N_12274,N_12195,N_12175);
nor U12275 (N_12275,N_12122,N_12155);
nand U12276 (N_12276,N_12070,N_12038);
nor U12277 (N_12277,N_12109,N_12120);
nand U12278 (N_12278,N_12177,N_12174);
or U12279 (N_12279,N_12146,N_12139);
nand U12280 (N_12280,N_12049,N_12055);
or U12281 (N_12281,N_12047,N_12156);
nor U12282 (N_12282,N_12194,N_12067);
nand U12283 (N_12283,N_12149,N_12117);
nand U12284 (N_12284,N_12058,N_12009);
nor U12285 (N_12285,N_12119,N_12094);
nand U12286 (N_12286,N_12090,N_12182);
or U12287 (N_12287,N_12074,N_12096);
xnor U12288 (N_12288,N_12127,N_12008);
nand U12289 (N_12289,N_12163,N_12016);
or U12290 (N_12290,N_12128,N_12165);
nor U12291 (N_12291,N_12102,N_12136);
and U12292 (N_12292,N_12012,N_12157);
or U12293 (N_12293,N_12056,N_12088);
or U12294 (N_12294,N_12158,N_12105);
nor U12295 (N_12295,N_12020,N_12114);
nand U12296 (N_12296,N_12042,N_12172);
and U12297 (N_12297,N_12190,N_12188);
xor U12298 (N_12298,N_12112,N_12162);
nand U12299 (N_12299,N_12133,N_12079);
nand U12300 (N_12300,N_12117,N_12185);
or U12301 (N_12301,N_12157,N_12126);
and U12302 (N_12302,N_12068,N_12197);
nand U12303 (N_12303,N_12098,N_12151);
nand U12304 (N_12304,N_12135,N_12025);
and U12305 (N_12305,N_12108,N_12055);
nor U12306 (N_12306,N_12094,N_12182);
xor U12307 (N_12307,N_12199,N_12049);
nor U12308 (N_12308,N_12139,N_12099);
nand U12309 (N_12309,N_12029,N_12198);
nor U12310 (N_12310,N_12146,N_12188);
nand U12311 (N_12311,N_12136,N_12132);
and U12312 (N_12312,N_12125,N_12188);
or U12313 (N_12313,N_12143,N_12105);
and U12314 (N_12314,N_12017,N_12183);
nor U12315 (N_12315,N_12106,N_12097);
nand U12316 (N_12316,N_12009,N_12129);
or U12317 (N_12317,N_12055,N_12146);
and U12318 (N_12318,N_12158,N_12192);
nor U12319 (N_12319,N_12063,N_12050);
xnor U12320 (N_12320,N_12151,N_12082);
nor U12321 (N_12321,N_12086,N_12058);
or U12322 (N_12322,N_12121,N_12159);
nand U12323 (N_12323,N_12041,N_12112);
or U12324 (N_12324,N_12179,N_12197);
and U12325 (N_12325,N_12192,N_12169);
or U12326 (N_12326,N_12018,N_12033);
and U12327 (N_12327,N_12112,N_12185);
and U12328 (N_12328,N_12182,N_12191);
and U12329 (N_12329,N_12092,N_12065);
and U12330 (N_12330,N_12017,N_12146);
xor U12331 (N_12331,N_12038,N_12155);
and U12332 (N_12332,N_12042,N_12095);
or U12333 (N_12333,N_12054,N_12135);
nor U12334 (N_12334,N_12029,N_12056);
nand U12335 (N_12335,N_12177,N_12106);
xnor U12336 (N_12336,N_12111,N_12098);
nand U12337 (N_12337,N_12025,N_12028);
nor U12338 (N_12338,N_12063,N_12143);
and U12339 (N_12339,N_12086,N_12134);
xnor U12340 (N_12340,N_12145,N_12048);
nand U12341 (N_12341,N_12112,N_12128);
nor U12342 (N_12342,N_12010,N_12162);
nor U12343 (N_12343,N_12170,N_12115);
nor U12344 (N_12344,N_12051,N_12182);
and U12345 (N_12345,N_12026,N_12125);
nor U12346 (N_12346,N_12142,N_12129);
nor U12347 (N_12347,N_12026,N_12071);
or U12348 (N_12348,N_12150,N_12154);
nand U12349 (N_12349,N_12125,N_12140);
and U12350 (N_12350,N_12110,N_12010);
or U12351 (N_12351,N_12101,N_12150);
or U12352 (N_12352,N_12070,N_12146);
and U12353 (N_12353,N_12074,N_12009);
and U12354 (N_12354,N_12172,N_12112);
or U12355 (N_12355,N_12085,N_12138);
nor U12356 (N_12356,N_12093,N_12138);
nor U12357 (N_12357,N_12107,N_12152);
nand U12358 (N_12358,N_12193,N_12093);
nor U12359 (N_12359,N_12119,N_12010);
xnor U12360 (N_12360,N_12156,N_12171);
nand U12361 (N_12361,N_12103,N_12147);
nor U12362 (N_12362,N_12125,N_12099);
xnor U12363 (N_12363,N_12055,N_12046);
nor U12364 (N_12364,N_12069,N_12076);
xnor U12365 (N_12365,N_12106,N_12123);
xnor U12366 (N_12366,N_12029,N_12075);
and U12367 (N_12367,N_12112,N_12105);
and U12368 (N_12368,N_12036,N_12167);
or U12369 (N_12369,N_12081,N_12103);
or U12370 (N_12370,N_12060,N_12101);
nor U12371 (N_12371,N_12089,N_12025);
nor U12372 (N_12372,N_12026,N_12041);
nand U12373 (N_12373,N_12079,N_12102);
nand U12374 (N_12374,N_12004,N_12100);
nand U12375 (N_12375,N_12039,N_12136);
xnor U12376 (N_12376,N_12033,N_12134);
nor U12377 (N_12377,N_12002,N_12197);
nor U12378 (N_12378,N_12106,N_12113);
nor U12379 (N_12379,N_12072,N_12140);
or U12380 (N_12380,N_12192,N_12095);
and U12381 (N_12381,N_12035,N_12123);
or U12382 (N_12382,N_12006,N_12064);
nand U12383 (N_12383,N_12138,N_12198);
and U12384 (N_12384,N_12060,N_12086);
xnor U12385 (N_12385,N_12017,N_12007);
nand U12386 (N_12386,N_12050,N_12127);
nor U12387 (N_12387,N_12074,N_12023);
xor U12388 (N_12388,N_12145,N_12171);
nor U12389 (N_12389,N_12029,N_12039);
nand U12390 (N_12390,N_12057,N_12116);
or U12391 (N_12391,N_12136,N_12104);
and U12392 (N_12392,N_12074,N_12175);
and U12393 (N_12393,N_12104,N_12064);
nand U12394 (N_12394,N_12128,N_12022);
and U12395 (N_12395,N_12033,N_12184);
and U12396 (N_12396,N_12189,N_12124);
and U12397 (N_12397,N_12054,N_12096);
and U12398 (N_12398,N_12066,N_12175);
nand U12399 (N_12399,N_12180,N_12043);
xnor U12400 (N_12400,N_12256,N_12212);
nand U12401 (N_12401,N_12364,N_12239);
nor U12402 (N_12402,N_12230,N_12234);
nor U12403 (N_12403,N_12281,N_12302);
nor U12404 (N_12404,N_12251,N_12263);
nand U12405 (N_12405,N_12326,N_12201);
or U12406 (N_12406,N_12397,N_12386);
nand U12407 (N_12407,N_12345,N_12250);
nor U12408 (N_12408,N_12357,N_12210);
or U12409 (N_12409,N_12282,N_12334);
nor U12410 (N_12410,N_12280,N_12283);
and U12411 (N_12411,N_12394,N_12306);
nand U12412 (N_12412,N_12399,N_12307);
nor U12413 (N_12413,N_12314,N_12347);
nand U12414 (N_12414,N_12265,N_12366);
or U12415 (N_12415,N_12241,N_12275);
nor U12416 (N_12416,N_12367,N_12342);
and U12417 (N_12417,N_12365,N_12226);
nand U12418 (N_12418,N_12258,N_12341);
nand U12419 (N_12419,N_12264,N_12233);
nand U12420 (N_12420,N_12247,N_12296);
and U12421 (N_12421,N_12348,N_12203);
nor U12422 (N_12422,N_12242,N_12354);
or U12423 (N_12423,N_12317,N_12236);
and U12424 (N_12424,N_12385,N_12297);
nand U12425 (N_12425,N_12325,N_12391);
nand U12426 (N_12426,N_12315,N_12245);
nor U12427 (N_12427,N_12253,N_12299);
nand U12428 (N_12428,N_12272,N_12387);
nor U12429 (N_12429,N_12327,N_12329);
xnor U12430 (N_12430,N_12255,N_12309);
nand U12431 (N_12431,N_12262,N_12398);
nand U12432 (N_12432,N_12376,N_12213);
nor U12433 (N_12433,N_12286,N_12249);
and U12434 (N_12434,N_12279,N_12240);
nand U12435 (N_12435,N_12287,N_12211);
or U12436 (N_12436,N_12353,N_12337);
nand U12437 (N_12437,N_12328,N_12206);
nand U12438 (N_12438,N_12207,N_12349);
or U12439 (N_12439,N_12260,N_12300);
nor U12440 (N_12440,N_12323,N_12209);
and U12441 (N_12441,N_12316,N_12359);
or U12442 (N_12442,N_12295,N_12333);
nor U12443 (N_12443,N_12244,N_12267);
and U12444 (N_12444,N_12224,N_12340);
or U12445 (N_12445,N_12219,N_12202);
nand U12446 (N_12446,N_12285,N_12322);
and U12447 (N_12447,N_12220,N_12257);
and U12448 (N_12448,N_12273,N_12266);
and U12449 (N_12449,N_12370,N_12293);
nor U12450 (N_12450,N_12393,N_12392);
and U12451 (N_12451,N_12380,N_12320);
and U12452 (N_12452,N_12214,N_12311);
or U12453 (N_12453,N_12379,N_12248);
nand U12454 (N_12454,N_12259,N_12396);
or U12455 (N_12455,N_12352,N_12388);
or U12456 (N_12456,N_12355,N_12303);
nand U12457 (N_12457,N_12304,N_12301);
nor U12458 (N_12458,N_12390,N_12284);
nand U12459 (N_12459,N_12373,N_12338);
or U12460 (N_12460,N_12384,N_12344);
or U12461 (N_12461,N_12290,N_12254);
nor U12462 (N_12462,N_12288,N_12268);
and U12463 (N_12463,N_12270,N_12375);
and U12464 (N_12464,N_12318,N_12223);
or U12465 (N_12465,N_12368,N_12246);
nand U12466 (N_12466,N_12321,N_12332);
and U12467 (N_12467,N_12336,N_12389);
or U12468 (N_12468,N_12319,N_12271);
or U12469 (N_12469,N_12346,N_12229);
nand U12470 (N_12470,N_12363,N_12289);
nor U12471 (N_12471,N_12313,N_12330);
nand U12472 (N_12472,N_12217,N_12227);
or U12473 (N_12473,N_12231,N_12205);
nand U12474 (N_12474,N_12208,N_12204);
and U12475 (N_12475,N_12252,N_12228);
or U12476 (N_12476,N_12310,N_12222);
or U12477 (N_12477,N_12377,N_12351);
nand U12478 (N_12478,N_12274,N_12261);
nor U12479 (N_12479,N_12308,N_12324);
nand U12480 (N_12480,N_12361,N_12237);
nand U12481 (N_12481,N_12358,N_12360);
xnor U12482 (N_12482,N_12235,N_12294);
or U12483 (N_12483,N_12356,N_12298);
or U12484 (N_12484,N_12369,N_12362);
xnor U12485 (N_12485,N_12232,N_12383);
or U12486 (N_12486,N_12312,N_12292);
nand U12487 (N_12487,N_12350,N_12276);
or U12488 (N_12488,N_12200,N_12378);
nand U12489 (N_12489,N_12277,N_12225);
and U12490 (N_12490,N_12343,N_12305);
nor U12491 (N_12491,N_12291,N_12335);
nand U12492 (N_12492,N_12371,N_12374);
or U12493 (N_12493,N_12269,N_12243);
nand U12494 (N_12494,N_12278,N_12381);
or U12495 (N_12495,N_12216,N_12218);
nor U12496 (N_12496,N_12339,N_12372);
and U12497 (N_12497,N_12215,N_12221);
nand U12498 (N_12498,N_12238,N_12331);
xnor U12499 (N_12499,N_12395,N_12382);
nand U12500 (N_12500,N_12209,N_12285);
or U12501 (N_12501,N_12340,N_12373);
nor U12502 (N_12502,N_12236,N_12370);
nor U12503 (N_12503,N_12229,N_12260);
nor U12504 (N_12504,N_12285,N_12393);
nand U12505 (N_12505,N_12387,N_12228);
or U12506 (N_12506,N_12253,N_12214);
nand U12507 (N_12507,N_12225,N_12307);
nor U12508 (N_12508,N_12375,N_12307);
and U12509 (N_12509,N_12254,N_12364);
or U12510 (N_12510,N_12223,N_12267);
and U12511 (N_12511,N_12272,N_12371);
xnor U12512 (N_12512,N_12213,N_12340);
nand U12513 (N_12513,N_12357,N_12393);
or U12514 (N_12514,N_12274,N_12358);
or U12515 (N_12515,N_12244,N_12208);
nand U12516 (N_12516,N_12327,N_12363);
or U12517 (N_12517,N_12230,N_12266);
nand U12518 (N_12518,N_12295,N_12246);
nor U12519 (N_12519,N_12312,N_12296);
and U12520 (N_12520,N_12254,N_12347);
xor U12521 (N_12521,N_12361,N_12362);
or U12522 (N_12522,N_12342,N_12216);
or U12523 (N_12523,N_12366,N_12324);
or U12524 (N_12524,N_12338,N_12378);
xor U12525 (N_12525,N_12217,N_12222);
or U12526 (N_12526,N_12334,N_12274);
nand U12527 (N_12527,N_12227,N_12292);
nor U12528 (N_12528,N_12215,N_12225);
and U12529 (N_12529,N_12217,N_12308);
and U12530 (N_12530,N_12380,N_12328);
or U12531 (N_12531,N_12325,N_12320);
or U12532 (N_12532,N_12316,N_12243);
or U12533 (N_12533,N_12276,N_12207);
nor U12534 (N_12534,N_12200,N_12304);
nand U12535 (N_12535,N_12386,N_12362);
xnor U12536 (N_12536,N_12363,N_12309);
nand U12537 (N_12537,N_12396,N_12302);
nand U12538 (N_12538,N_12256,N_12298);
and U12539 (N_12539,N_12232,N_12272);
xor U12540 (N_12540,N_12318,N_12254);
nand U12541 (N_12541,N_12252,N_12333);
and U12542 (N_12542,N_12312,N_12261);
xor U12543 (N_12543,N_12392,N_12253);
nor U12544 (N_12544,N_12389,N_12276);
and U12545 (N_12545,N_12228,N_12367);
and U12546 (N_12546,N_12314,N_12238);
xor U12547 (N_12547,N_12266,N_12325);
and U12548 (N_12548,N_12307,N_12290);
nor U12549 (N_12549,N_12203,N_12261);
and U12550 (N_12550,N_12382,N_12346);
xor U12551 (N_12551,N_12278,N_12251);
or U12552 (N_12552,N_12361,N_12385);
or U12553 (N_12553,N_12247,N_12219);
nor U12554 (N_12554,N_12266,N_12241);
or U12555 (N_12555,N_12226,N_12319);
nand U12556 (N_12556,N_12304,N_12394);
and U12557 (N_12557,N_12355,N_12353);
and U12558 (N_12558,N_12349,N_12262);
nand U12559 (N_12559,N_12309,N_12384);
or U12560 (N_12560,N_12301,N_12225);
nor U12561 (N_12561,N_12216,N_12274);
or U12562 (N_12562,N_12385,N_12281);
or U12563 (N_12563,N_12346,N_12354);
or U12564 (N_12564,N_12388,N_12373);
xor U12565 (N_12565,N_12282,N_12359);
nor U12566 (N_12566,N_12264,N_12342);
nand U12567 (N_12567,N_12353,N_12285);
xnor U12568 (N_12568,N_12280,N_12239);
or U12569 (N_12569,N_12307,N_12391);
and U12570 (N_12570,N_12229,N_12302);
nand U12571 (N_12571,N_12386,N_12338);
or U12572 (N_12572,N_12294,N_12334);
and U12573 (N_12573,N_12337,N_12203);
nor U12574 (N_12574,N_12364,N_12217);
or U12575 (N_12575,N_12249,N_12232);
and U12576 (N_12576,N_12319,N_12213);
nor U12577 (N_12577,N_12321,N_12208);
or U12578 (N_12578,N_12368,N_12280);
xnor U12579 (N_12579,N_12276,N_12298);
nand U12580 (N_12580,N_12390,N_12279);
and U12581 (N_12581,N_12294,N_12248);
or U12582 (N_12582,N_12355,N_12270);
nor U12583 (N_12583,N_12228,N_12230);
and U12584 (N_12584,N_12376,N_12397);
and U12585 (N_12585,N_12214,N_12251);
nor U12586 (N_12586,N_12231,N_12366);
and U12587 (N_12587,N_12229,N_12287);
and U12588 (N_12588,N_12330,N_12302);
nand U12589 (N_12589,N_12239,N_12275);
and U12590 (N_12590,N_12213,N_12298);
or U12591 (N_12591,N_12262,N_12273);
nand U12592 (N_12592,N_12317,N_12318);
and U12593 (N_12593,N_12355,N_12279);
nor U12594 (N_12594,N_12395,N_12303);
nor U12595 (N_12595,N_12227,N_12238);
nor U12596 (N_12596,N_12381,N_12366);
or U12597 (N_12597,N_12240,N_12395);
and U12598 (N_12598,N_12398,N_12327);
nand U12599 (N_12599,N_12312,N_12367);
and U12600 (N_12600,N_12497,N_12585);
and U12601 (N_12601,N_12501,N_12413);
and U12602 (N_12602,N_12534,N_12402);
nand U12603 (N_12603,N_12547,N_12579);
xnor U12604 (N_12604,N_12480,N_12594);
and U12605 (N_12605,N_12537,N_12505);
and U12606 (N_12606,N_12464,N_12493);
or U12607 (N_12607,N_12460,N_12409);
and U12608 (N_12608,N_12449,N_12439);
and U12609 (N_12609,N_12452,N_12580);
nand U12610 (N_12610,N_12471,N_12578);
xnor U12611 (N_12611,N_12477,N_12442);
or U12612 (N_12612,N_12473,N_12592);
nand U12613 (N_12613,N_12433,N_12516);
nand U12614 (N_12614,N_12487,N_12444);
xnor U12615 (N_12615,N_12500,N_12559);
nor U12616 (N_12616,N_12535,N_12539);
and U12617 (N_12617,N_12568,N_12434);
nand U12618 (N_12618,N_12507,N_12514);
nand U12619 (N_12619,N_12446,N_12510);
nand U12620 (N_12620,N_12408,N_12426);
nand U12621 (N_12621,N_12599,N_12575);
xor U12622 (N_12622,N_12572,N_12486);
or U12623 (N_12623,N_12489,N_12569);
nand U12624 (N_12624,N_12561,N_12520);
nand U12625 (N_12625,N_12437,N_12483);
and U12626 (N_12626,N_12523,N_12427);
and U12627 (N_12627,N_12590,N_12411);
nand U12628 (N_12628,N_12525,N_12588);
or U12629 (N_12629,N_12491,N_12546);
or U12630 (N_12630,N_12541,N_12492);
or U12631 (N_12631,N_12574,N_12414);
or U12632 (N_12632,N_12416,N_12481);
xor U12633 (N_12633,N_12531,N_12404);
nor U12634 (N_12634,N_12456,N_12478);
or U12635 (N_12635,N_12540,N_12519);
nand U12636 (N_12636,N_12528,N_12401);
or U12637 (N_12637,N_12428,N_12445);
and U12638 (N_12638,N_12403,N_12530);
and U12639 (N_12639,N_12515,N_12584);
nor U12640 (N_12640,N_12593,N_12412);
or U12641 (N_12641,N_12479,N_12508);
and U12642 (N_12642,N_12533,N_12443);
nor U12643 (N_12643,N_12474,N_12488);
nor U12644 (N_12644,N_12462,N_12415);
nor U12645 (N_12645,N_12577,N_12564);
or U12646 (N_12646,N_12591,N_12556);
and U12647 (N_12647,N_12466,N_12495);
and U12648 (N_12648,N_12566,N_12406);
or U12649 (N_12649,N_12405,N_12562);
nor U12650 (N_12650,N_12467,N_12576);
nand U12651 (N_12651,N_12513,N_12551);
and U12652 (N_12652,N_12554,N_12450);
xor U12653 (N_12653,N_12553,N_12423);
nor U12654 (N_12654,N_12490,N_12407);
or U12655 (N_12655,N_12598,N_12506);
nor U12656 (N_12656,N_12532,N_12430);
nor U12657 (N_12657,N_12472,N_12476);
nand U12658 (N_12658,N_12435,N_12499);
or U12659 (N_12659,N_12461,N_12468);
nor U12660 (N_12660,N_12571,N_12438);
nor U12661 (N_12661,N_12587,N_12498);
nand U12662 (N_12662,N_12440,N_12447);
or U12663 (N_12663,N_12589,N_12453);
and U12664 (N_12664,N_12543,N_12454);
or U12665 (N_12665,N_12545,N_12536);
nand U12666 (N_12666,N_12521,N_12470);
nor U12667 (N_12667,N_12418,N_12563);
xor U12668 (N_12668,N_12511,N_12573);
nand U12669 (N_12669,N_12496,N_12529);
and U12670 (N_12670,N_12421,N_12560);
nor U12671 (N_12671,N_12484,N_12522);
xnor U12672 (N_12672,N_12552,N_12567);
nor U12673 (N_12673,N_12595,N_12597);
nand U12674 (N_12674,N_12526,N_12596);
nor U12675 (N_12675,N_12517,N_12429);
xnor U12676 (N_12676,N_12544,N_12441);
and U12677 (N_12677,N_12548,N_12581);
or U12678 (N_12678,N_12512,N_12503);
or U12679 (N_12679,N_12457,N_12459);
and U12680 (N_12680,N_12419,N_12422);
xnor U12681 (N_12681,N_12518,N_12420);
nand U12682 (N_12682,N_12475,N_12425);
nand U12683 (N_12683,N_12504,N_12469);
and U12684 (N_12684,N_12570,N_12558);
nor U12685 (N_12685,N_12550,N_12400);
or U12686 (N_12686,N_12494,N_12527);
xnor U12687 (N_12687,N_12538,N_12482);
and U12688 (N_12688,N_12583,N_12485);
and U12689 (N_12689,N_12431,N_12542);
nor U12690 (N_12690,N_12451,N_12436);
nand U12691 (N_12691,N_12502,N_12458);
or U12692 (N_12692,N_12509,N_12565);
nand U12693 (N_12693,N_12582,N_12455);
and U12694 (N_12694,N_12424,N_12555);
nand U12695 (N_12695,N_12557,N_12417);
or U12696 (N_12696,N_12448,N_12410);
or U12697 (N_12697,N_12465,N_12432);
nor U12698 (N_12698,N_12586,N_12524);
nor U12699 (N_12699,N_12549,N_12463);
nand U12700 (N_12700,N_12479,N_12501);
xor U12701 (N_12701,N_12571,N_12545);
nand U12702 (N_12702,N_12564,N_12486);
nand U12703 (N_12703,N_12527,N_12537);
nand U12704 (N_12704,N_12416,N_12471);
or U12705 (N_12705,N_12535,N_12413);
and U12706 (N_12706,N_12552,N_12557);
or U12707 (N_12707,N_12553,N_12457);
xnor U12708 (N_12708,N_12513,N_12488);
nand U12709 (N_12709,N_12505,N_12568);
or U12710 (N_12710,N_12413,N_12537);
or U12711 (N_12711,N_12520,N_12593);
xnor U12712 (N_12712,N_12431,N_12539);
and U12713 (N_12713,N_12407,N_12418);
nand U12714 (N_12714,N_12531,N_12532);
nand U12715 (N_12715,N_12591,N_12540);
and U12716 (N_12716,N_12526,N_12404);
xor U12717 (N_12717,N_12583,N_12472);
and U12718 (N_12718,N_12437,N_12579);
nand U12719 (N_12719,N_12446,N_12498);
and U12720 (N_12720,N_12586,N_12474);
and U12721 (N_12721,N_12476,N_12416);
nand U12722 (N_12722,N_12541,N_12418);
and U12723 (N_12723,N_12426,N_12500);
or U12724 (N_12724,N_12468,N_12568);
or U12725 (N_12725,N_12545,N_12404);
nor U12726 (N_12726,N_12432,N_12438);
or U12727 (N_12727,N_12562,N_12433);
nor U12728 (N_12728,N_12506,N_12586);
and U12729 (N_12729,N_12411,N_12505);
nor U12730 (N_12730,N_12461,N_12400);
nor U12731 (N_12731,N_12485,N_12565);
nor U12732 (N_12732,N_12515,N_12599);
or U12733 (N_12733,N_12570,N_12490);
nor U12734 (N_12734,N_12565,N_12407);
nor U12735 (N_12735,N_12485,N_12466);
and U12736 (N_12736,N_12427,N_12434);
and U12737 (N_12737,N_12574,N_12553);
nor U12738 (N_12738,N_12486,N_12546);
or U12739 (N_12739,N_12501,N_12596);
nor U12740 (N_12740,N_12502,N_12477);
and U12741 (N_12741,N_12408,N_12513);
nand U12742 (N_12742,N_12588,N_12478);
nand U12743 (N_12743,N_12589,N_12563);
nand U12744 (N_12744,N_12495,N_12490);
nand U12745 (N_12745,N_12488,N_12572);
nor U12746 (N_12746,N_12549,N_12448);
xor U12747 (N_12747,N_12519,N_12535);
nand U12748 (N_12748,N_12429,N_12586);
or U12749 (N_12749,N_12514,N_12408);
and U12750 (N_12750,N_12455,N_12523);
nor U12751 (N_12751,N_12532,N_12526);
xor U12752 (N_12752,N_12510,N_12593);
nand U12753 (N_12753,N_12562,N_12484);
or U12754 (N_12754,N_12483,N_12449);
or U12755 (N_12755,N_12401,N_12556);
nor U12756 (N_12756,N_12517,N_12574);
nand U12757 (N_12757,N_12538,N_12567);
or U12758 (N_12758,N_12452,N_12409);
xor U12759 (N_12759,N_12412,N_12536);
and U12760 (N_12760,N_12482,N_12444);
or U12761 (N_12761,N_12431,N_12447);
and U12762 (N_12762,N_12523,N_12513);
xor U12763 (N_12763,N_12460,N_12540);
or U12764 (N_12764,N_12576,N_12505);
nor U12765 (N_12765,N_12479,N_12596);
nor U12766 (N_12766,N_12530,N_12519);
nor U12767 (N_12767,N_12505,N_12416);
nand U12768 (N_12768,N_12497,N_12467);
and U12769 (N_12769,N_12594,N_12408);
nor U12770 (N_12770,N_12440,N_12505);
nor U12771 (N_12771,N_12413,N_12432);
nand U12772 (N_12772,N_12521,N_12515);
or U12773 (N_12773,N_12538,N_12421);
or U12774 (N_12774,N_12400,N_12532);
and U12775 (N_12775,N_12581,N_12410);
and U12776 (N_12776,N_12567,N_12432);
nand U12777 (N_12777,N_12427,N_12452);
nor U12778 (N_12778,N_12477,N_12511);
xor U12779 (N_12779,N_12467,N_12438);
xnor U12780 (N_12780,N_12590,N_12596);
nand U12781 (N_12781,N_12557,N_12424);
and U12782 (N_12782,N_12552,N_12455);
nor U12783 (N_12783,N_12502,N_12532);
and U12784 (N_12784,N_12497,N_12514);
or U12785 (N_12785,N_12407,N_12434);
nand U12786 (N_12786,N_12419,N_12509);
nand U12787 (N_12787,N_12540,N_12512);
xnor U12788 (N_12788,N_12503,N_12581);
nand U12789 (N_12789,N_12465,N_12544);
and U12790 (N_12790,N_12573,N_12472);
and U12791 (N_12791,N_12430,N_12404);
or U12792 (N_12792,N_12565,N_12544);
xor U12793 (N_12793,N_12417,N_12500);
nor U12794 (N_12794,N_12486,N_12475);
xor U12795 (N_12795,N_12505,N_12535);
and U12796 (N_12796,N_12505,N_12585);
or U12797 (N_12797,N_12469,N_12465);
nor U12798 (N_12798,N_12523,N_12526);
and U12799 (N_12799,N_12498,N_12415);
xor U12800 (N_12800,N_12719,N_12705);
nand U12801 (N_12801,N_12750,N_12709);
and U12802 (N_12802,N_12734,N_12736);
and U12803 (N_12803,N_12692,N_12783);
and U12804 (N_12804,N_12745,N_12754);
nand U12805 (N_12805,N_12796,N_12684);
and U12806 (N_12806,N_12603,N_12649);
nor U12807 (N_12807,N_12704,N_12670);
nor U12808 (N_12808,N_12673,N_12730);
or U12809 (N_12809,N_12729,N_12635);
or U12810 (N_12810,N_12721,N_12623);
nor U12811 (N_12811,N_12767,N_12795);
nand U12812 (N_12812,N_12689,N_12791);
nand U12813 (N_12813,N_12798,N_12607);
xor U12814 (N_12814,N_12661,N_12696);
nor U12815 (N_12815,N_12768,N_12714);
xor U12816 (N_12816,N_12735,N_12782);
nor U12817 (N_12817,N_12794,N_12604);
or U12818 (N_12818,N_12761,N_12668);
nor U12819 (N_12819,N_12606,N_12618);
and U12820 (N_12820,N_12741,N_12781);
nor U12821 (N_12821,N_12642,N_12631);
and U12822 (N_12822,N_12720,N_12609);
nand U12823 (N_12823,N_12725,N_12713);
xnor U12824 (N_12824,N_12742,N_12625);
nand U12825 (N_12825,N_12777,N_12667);
nand U12826 (N_12826,N_12664,N_12722);
and U12827 (N_12827,N_12680,N_12724);
nand U12828 (N_12828,N_12715,N_12786);
nor U12829 (N_12829,N_12691,N_12651);
and U12830 (N_12830,N_12697,N_12608);
or U12831 (N_12831,N_12706,N_12634);
or U12832 (N_12832,N_12656,N_12749);
nand U12833 (N_12833,N_12797,N_12646);
nand U12834 (N_12834,N_12717,N_12698);
xnor U12835 (N_12835,N_12764,N_12601);
nand U12836 (N_12836,N_12622,N_12650);
nor U12837 (N_12837,N_12658,N_12732);
and U12838 (N_12838,N_12748,N_12645);
nand U12839 (N_12839,N_12653,N_12716);
nor U12840 (N_12840,N_12612,N_12637);
or U12841 (N_12841,N_12702,N_12699);
and U12842 (N_12842,N_12688,N_12703);
nor U12843 (N_12843,N_12752,N_12681);
nand U12844 (N_12844,N_12652,N_12683);
nor U12845 (N_12845,N_12687,N_12643);
or U12846 (N_12846,N_12627,N_12787);
nor U12847 (N_12847,N_12677,N_12740);
or U12848 (N_12848,N_12780,N_12682);
and U12849 (N_12849,N_12640,N_12728);
nor U12850 (N_12850,N_12785,N_12778);
nor U12851 (N_12851,N_12753,N_12774);
and U12852 (N_12852,N_12723,N_12746);
and U12853 (N_12853,N_12769,N_12611);
and U12854 (N_12854,N_12657,N_12685);
nand U12855 (N_12855,N_12737,N_12636);
nand U12856 (N_12856,N_12788,N_12708);
or U12857 (N_12857,N_12617,N_12600);
nand U12858 (N_12858,N_12676,N_12632);
xor U12859 (N_12859,N_12765,N_12789);
or U12860 (N_12860,N_12662,N_12647);
and U12861 (N_12861,N_12638,N_12710);
nor U12862 (N_12862,N_12763,N_12672);
xor U12863 (N_12863,N_12610,N_12629);
nand U12864 (N_12864,N_12744,N_12621);
nand U12865 (N_12865,N_12731,N_12700);
nand U12866 (N_12866,N_12613,N_12678);
nand U12867 (N_12867,N_12711,N_12799);
nand U12868 (N_12868,N_12679,N_12747);
nor U12869 (N_12869,N_12790,N_12760);
nor U12870 (N_12870,N_12644,N_12766);
nor U12871 (N_12871,N_12793,N_12686);
or U12872 (N_12872,N_12639,N_12619);
nand U12873 (N_12873,N_12771,N_12701);
nor U12874 (N_12874,N_12773,N_12733);
nand U12875 (N_12875,N_12671,N_12762);
and U12876 (N_12876,N_12675,N_12620);
and U12877 (N_12877,N_12690,N_12712);
or U12878 (N_12878,N_12738,N_12695);
and U12879 (N_12879,N_12630,N_12674);
nor U12880 (N_12880,N_12772,N_12726);
xnor U12881 (N_12881,N_12663,N_12779);
nor U12882 (N_12882,N_12624,N_12707);
nand U12883 (N_12883,N_12693,N_12633);
nand U12884 (N_12884,N_12665,N_12784);
or U12885 (N_12885,N_12605,N_12614);
nand U12886 (N_12886,N_12641,N_12770);
xor U12887 (N_12887,N_12739,N_12757);
or U12888 (N_12888,N_12756,N_12755);
xor U12889 (N_12889,N_12743,N_12602);
and U12890 (N_12890,N_12727,N_12669);
or U12891 (N_12891,N_12666,N_12775);
and U12892 (N_12892,N_12616,N_12615);
nor U12893 (N_12893,N_12751,N_12792);
or U12894 (N_12894,N_12626,N_12758);
nor U12895 (N_12895,N_12654,N_12659);
nor U12896 (N_12896,N_12718,N_12655);
nand U12897 (N_12897,N_12648,N_12759);
nor U12898 (N_12898,N_12776,N_12660);
and U12899 (N_12899,N_12694,N_12628);
and U12900 (N_12900,N_12607,N_12678);
nor U12901 (N_12901,N_12768,N_12724);
or U12902 (N_12902,N_12751,N_12704);
xor U12903 (N_12903,N_12649,N_12690);
and U12904 (N_12904,N_12726,N_12799);
and U12905 (N_12905,N_12677,N_12625);
nor U12906 (N_12906,N_12619,N_12704);
or U12907 (N_12907,N_12791,N_12668);
nor U12908 (N_12908,N_12775,N_12675);
nand U12909 (N_12909,N_12682,N_12645);
or U12910 (N_12910,N_12692,N_12702);
nand U12911 (N_12911,N_12791,N_12601);
and U12912 (N_12912,N_12628,N_12793);
or U12913 (N_12913,N_12687,N_12770);
or U12914 (N_12914,N_12694,N_12631);
or U12915 (N_12915,N_12750,N_12677);
and U12916 (N_12916,N_12776,N_12756);
or U12917 (N_12917,N_12647,N_12714);
nor U12918 (N_12918,N_12650,N_12694);
and U12919 (N_12919,N_12768,N_12754);
nor U12920 (N_12920,N_12733,N_12707);
and U12921 (N_12921,N_12765,N_12714);
and U12922 (N_12922,N_12604,N_12762);
nor U12923 (N_12923,N_12619,N_12680);
xor U12924 (N_12924,N_12633,N_12727);
and U12925 (N_12925,N_12612,N_12794);
nand U12926 (N_12926,N_12703,N_12750);
nand U12927 (N_12927,N_12744,N_12628);
nor U12928 (N_12928,N_12655,N_12773);
nor U12929 (N_12929,N_12691,N_12661);
and U12930 (N_12930,N_12792,N_12678);
or U12931 (N_12931,N_12662,N_12785);
nand U12932 (N_12932,N_12702,N_12729);
nor U12933 (N_12933,N_12722,N_12610);
or U12934 (N_12934,N_12625,N_12741);
and U12935 (N_12935,N_12732,N_12617);
nand U12936 (N_12936,N_12793,N_12674);
xor U12937 (N_12937,N_12613,N_12755);
or U12938 (N_12938,N_12760,N_12617);
and U12939 (N_12939,N_12767,N_12675);
or U12940 (N_12940,N_12603,N_12783);
or U12941 (N_12941,N_12705,N_12615);
xnor U12942 (N_12942,N_12723,N_12740);
nor U12943 (N_12943,N_12739,N_12795);
and U12944 (N_12944,N_12635,N_12706);
or U12945 (N_12945,N_12619,N_12762);
or U12946 (N_12946,N_12633,N_12630);
nand U12947 (N_12947,N_12665,N_12799);
nand U12948 (N_12948,N_12785,N_12660);
nand U12949 (N_12949,N_12657,N_12656);
or U12950 (N_12950,N_12664,N_12709);
nand U12951 (N_12951,N_12614,N_12641);
or U12952 (N_12952,N_12697,N_12609);
and U12953 (N_12953,N_12614,N_12679);
nand U12954 (N_12954,N_12644,N_12601);
nand U12955 (N_12955,N_12740,N_12689);
xor U12956 (N_12956,N_12727,N_12705);
or U12957 (N_12957,N_12792,N_12630);
nor U12958 (N_12958,N_12729,N_12732);
and U12959 (N_12959,N_12758,N_12643);
nor U12960 (N_12960,N_12727,N_12608);
and U12961 (N_12961,N_12777,N_12789);
or U12962 (N_12962,N_12712,N_12672);
and U12963 (N_12963,N_12695,N_12658);
or U12964 (N_12964,N_12663,N_12713);
xor U12965 (N_12965,N_12641,N_12696);
or U12966 (N_12966,N_12776,N_12757);
or U12967 (N_12967,N_12732,N_12627);
or U12968 (N_12968,N_12725,N_12778);
and U12969 (N_12969,N_12626,N_12780);
nor U12970 (N_12970,N_12781,N_12698);
nor U12971 (N_12971,N_12624,N_12685);
nand U12972 (N_12972,N_12682,N_12738);
nand U12973 (N_12973,N_12691,N_12757);
nor U12974 (N_12974,N_12658,N_12659);
nor U12975 (N_12975,N_12649,N_12778);
nor U12976 (N_12976,N_12718,N_12778);
or U12977 (N_12977,N_12775,N_12674);
nor U12978 (N_12978,N_12685,N_12687);
and U12979 (N_12979,N_12722,N_12715);
or U12980 (N_12980,N_12697,N_12619);
or U12981 (N_12981,N_12684,N_12741);
and U12982 (N_12982,N_12608,N_12712);
nor U12983 (N_12983,N_12676,N_12761);
xor U12984 (N_12984,N_12786,N_12692);
and U12985 (N_12985,N_12668,N_12679);
xnor U12986 (N_12986,N_12650,N_12767);
or U12987 (N_12987,N_12669,N_12705);
nand U12988 (N_12988,N_12719,N_12779);
nand U12989 (N_12989,N_12717,N_12739);
and U12990 (N_12990,N_12787,N_12727);
and U12991 (N_12991,N_12744,N_12720);
or U12992 (N_12992,N_12605,N_12728);
or U12993 (N_12993,N_12622,N_12743);
or U12994 (N_12994,N_12775,N_12694);
and U12995 (N_12995,N_12672,N_12644);
nor U12996 (N_12996,N_12609,N_12649);
nand U12997 (N_12997,N_12792,N_12672);
and U12998 (N_12998,N_12636,N_12648);
nor U12999 (N_12999,N_12664,N_12686);
and U13000 (N_13000,N_12825,N_12914);
or U13001 (N_13001,N_12916,N_12814);
and U13002 (N_13002,N_12919,N_12805);
and U13003 (N_13003,N_12828,N_12834);
nor U13004 (N_13004,N_12965,N_12820);
or U13005 (N_13005,N_12842,N_12878);
or U13006 (N_13006,N_12997,N_12956);
nor U13007 (N_13007,N_12909,N_12926);
nor U13008 (N_13008,N_12801,N_12806);
or U13009 (N_13009,N_12959,N_12870);
and U13010 (N_13010,N_12984,N_12857);
nand U13011 (N_13011,N_12838,N_12999);
and U13012 (N_13012,N_12970,N_12827);
xnor U13013 (N_13013,N_12837,N_12949);
nand U13014 (N_13014,N_12951,N_12869);
nand U13015 (N_13015,N_12811,N_12867);
nand U13016 (N_13016,N_12856,N_12860);
nor U13017 (N_13017,N_12912,N_12808);
xnor U13018 (N_13018,N_12928,N_12908);
xor U13019 (N_13019,N_12897,N_12843);
and U13020 (N_13020,N_12937,N_12985);
or U13021 (N_13021,N_12812,N_12960);
nor U13022 (N_13022,N_12891,N_12952);
nand U13023 (N_13023,N_12854,N_12815);
nand U13024 (N_13024,N_12818,N_12849);
or U13025 (N_13025,N_12941,N_12976);
xnor U13026 (N_13026,N_12879,N_12865);
nor U13027 (N_13027,N_12872,N_12836);
nand U13028 (N_13028,N_12800,N_12840);
and U13029 (N_13029,N_12992,N_12925);
xnor U13030 (N_13030,N_12807,N_12968);
and U13031 (N_13031,N_12957,N_12998);
and U13032 (N_13032,N_12917,N_12927);
nand U13033 (N_13033,N_12948,N_12933);
and U13034 (N_13034,N_12996,N_12905);
nand U13035 (N_13035,N_12884,N_12893);
nand U13036 (N_13036,N_12974,N_12923);
nand U13037 (N_13037,N_12846,N_12841);
and U13038 (N_13038,N_12946,N_12902);
nor U13039 (N_13039,N_12901,N_12889);
or U13040 (N_13040,N_12866,N_12898);
and U13041 (N_13041,N_12953,N_12848);
nand U13042 (N_13042,N_12899,N_12903);
or U13043 (N_13043,N_12862,N_12940);
or U13044 (N_13044,N_12881,N_12822);
and U13045 (N_13045,N_12904,N_12887);
nor U13046 (N_13046,N_12935,N_12880);
and U13047 (N_13047,N_12885,N_12924);
nor U13048 (N_13048,N_12971,N_12829);
nand U13049 (N_13049,N_12873,N_12930);
nand U13050 (N_13050,N_12906,N_12876);
xnor U13051 (N_13051,N_12844,N_12890);
and U13052 (N_13052,N_12810,N_12910);
nor U13053 (N_13053,N_12804,N_12967);
nor U13054 (N_13054,N_12934,N_12817);
nand U13055 (N_13055,N_12882,N_12803);
and U13056 (N_13056,N_12947,N_12877);
and U13057 (N_13057,N_12875,N_12955);
nor U13058 (N_13058,N_12987,N_12830);
nand U13059 (N_13059,N_12921,N_12826);
or U13060 (N_13060,N_12961,N_12942);
nand U13061 (N_13061,N_12858,N_12945);
nor U13062 (N_13062,N_12993,N_12964);
and U13063 (N_13063,N_12939,N_12943);
or U13064 (N_13064,N_12809,N_12991);
nand U13065 (N_13065,N_12832,N_12819);
and U13066 (N_13066,N_12978,N_12894);
or U13067 (N_13067,N_12833,N_12977);
nor U13068 (N_13068,N_12835,N_12831);
nand U13069 (N_13069,N_12938,N_12975);
nor U13070 (N_13070,N_12918,N_12915);
and U13071 (N_13071,N_12845,N_12907);
and U13072 (N_13072,N_12864,N_12980);
xor U13073 (N_13073,N_12802,N_12913);
or U13074 (N_13074,N_12981,N_12958);
or U13075 (N_13075,N_12839,N_12994);
and U13076 (N_13076,N_12895,N_12989);
or U13077 (N_13077,N_12813,N_12954);
nand U13078 (N_13078,N_12972,N_12896);
xnor U13079 (N_13079,N_12986,N_12868);
xnor U13080 (N_13080,N_12911,N_12932);
nand U13081 (N_13081,N_12874,N_12886);
or U13082 (N_13082,N_12821,N_12861);
nor U13083 (N_13083,N_12892,N_12859);
and U13084 (N_13084,N_12969,N_12847);
nand U13085 (N_13085,N_12853,N_12963);
nor U13086 (N_13086,N_12823,N_12900);
nand U13087 (N_13087,N_12995,N_12855);
xor U13088 (N_13088,N_12950,N_12922);
or U13089 (N_13089,N_12990,N_12888);
and U13090 (N_13090,N_12824,N_12816);
and U13091 (N_13091,N_12920,N_12871);
and U13092 (N_13092,N_12944,N_12988);
nor U13093 (N_13093,N_12962,N_12863);
or U13094 (N_13094,N_12982,N_12852);
or U13095 (N_13095,N_12883,N_12966);
or U13096 (N_13096,N_12973,N_12931);
or U13097 (N_13097,N_12850,N_12851);
and U13098 (N_13098,N_12929,N_12983);
and U13099 (N_13099,N_12979,N_12936);
or U13100 (N_13100,N_12912,N_12942);
nor U13101 (N_13101,N_12887,N_12998);
xor U13102 (N_13102,N_12920,N_12937);
nand U13103 (N_13103,N_12856,N_12830);
or U13104 (N_13104,N_12897,N_12905);
nor U13105 (N_13105,N_12869,N_12905);
and U13106 (N_13106,N_12885,N_12858);
xnor U13107 (N_13107,N_12973,N_12907);
nor U13108 (N_13108,N_12803,N_12844);
nor U13109 (N_13109,N_12876,N_12904);
nand U13110 (N_13110,N_12959,N_12836);
nor U13111 (N_13111,N_12815,N_12969);
nand U13112 (N_13112,N_12856,N_12816);
and U13113 (N_13113,N_12998,N_12918);
nor U13114 (N_13114,N_12832,N_12887);
nand U13115 (N_13115,N_12887,N_12804);
nand U13116 (N_13116,N_12984,N_12821);
and U13117 (N_13117,N_12891,N_12846);
or U13118 (N_13118,N_12811,N_12919);
and U13119 (N_13119,N_12996,N_12824);
nor U13120 (N_13120,N_12911,N_12841);
and U13121 (N_13121,N_12863,N_12927);
nand U13122 (N_13122,N_12853,N_12996);
or U13123 (N_13123,N_12849,N_12815);
nor U13124 (N_13124,N_12857,N_12981);
nand U13125 (N_13125,N_12806,N_12951);
nand U13126 (N_13126,N_12872,N_12966);
or U13127 (N_13127,N_12826,N_12842);
xnor U13128 (N_13128,N_12934,N_12991);
and U13129 (N_13129,N_12850,N_12891);
nand U13130 (N_13130,N_12880,N_12996);
and U13131 (N_13131,N_12871,N_12893);
and U13132 (N_13132,N_12886,N_12967);
nor U13133 (N_13133,N_12986,N_12969);
nand U13134 (N_13134,N_12981,N_12903);
and U13135 (N_13135,N_12942,N_12849);
and U13136 (N_13136,N_12834,N_12925);
and U13137 (N_13137,N_12946,N_12898);
xor U13138 (N_13138,N_12977,N_12837);
xnor U13139 (N_13139,N_12952,N_12842);
nand U13140 (N_13140,N_12971,N_12974);
nand U13141 (N_13141,N_12971,N_12929);
or U13142 (N_13142,N_12956,N_12941);
nor U13143 (N_13143,N_12914,N_12927);
and U13144 (N_13144,N_12808,N_12950);
nor U13145 (N_13145,N_12859,N_12978);
nand U13146 (N_13146,N_12952,N_12887);
nor U13147 (N_13147,N_12817,N_12868);
or U13148 (N_13148,N_12903,N_12907);
and U13149 (N_13149,N_12894,N_12917);
xor U13150 (N_13150,N_12839,N_12939);
or U13151 (N_13151,N_12934,N_12953);
or U13152 (N_13152,N_12823,N_12968);
nand U13153 (N_13153,N_12943,N_12970);
or U13154 (N_13154,N_12845,N_12834);
or U13155 (N_13155,N_12983,N_12837);
xnor U13156 (N_13156,N_12929,N_12950);
xnor U13157 (N_13157,N_12924,N_12804);
nor U13158 (N_13158,N_12924,N_12997);
nor U13159 (N_13159,N_12998,N_12883);
xor U13160 (N_13160,N_12828,N_12808);
nand U13161 (N_13161,N_12931,N_12949);
nor U13162 (N_13162,N_12814,N_12915);
xnor U13163 (N_13163,N_12872,N_12983);
and U13164 (N_13164,N_12981,N_12990);
or U13165 (N_13165,N_12806,N_12917);
nand U13166 (N_13166,N_12999,N_12988);
nor U13167 (N_13167,N_12930,N_12866);
and U13168 (N_13168,N_12931,N_12960);
nand U13169 (N_13169,N_12943,N_12911);
or U13170 (N_13170,N_12905,N_12834);
xor U13171 (N_13171,N_12820,N_12968);
nand U13172 (N_13172,N_12992,N_12885);
and U13173 (N_13173,N_12827,N_12908);
nor U13174 (N_13174,N_12817,N_12906);
and U13175 (N_13175,N_12845,N_12935);
or U13176 (N_13176,N_12813,N_12897);
or U13177 (N_13177,N_12813,N_12957);
nor U13178 (N_13178,N_12912,N_12867);
nand U13179 (N_13179,N_12893,N_12973);
nor U13180 (N_13180,N_12909,N_12920);
and U13181 (N_13181,N_12964,N_12846);
xnor U13182 (N_13182,N_12915,N_12951);
nand U13183 (N_13183,N_12823,N_12990);
or U13184 (N_13184,N_12952,N_12816);
nor U13185 (N_13185,N_12803,N_12832);
nor U13186 (N_13186,N_12821,N_12871);
nor U13187 (N_13187,N_12919,N_12860);
nand U13188 (N_13188,N_12975,N_12929);
and U13189 (N_13189,N_12954,N_12855);
xnor U13190 (N_13190,N_12903,N_12876);
nand U13191 (N_13191,N_12938,N_12857);
nor U13192 (N_13192,N_12964,N_12978);
nand U13193 (N_13193,N_12972,N_12876);
or U13194 (N_13194,N_12814,N_12870);
xor U13195 (N_13195,N_12841,N_12905);
nor U13196 (N_13196,N_12950,N_12869);
nand U13197 (N_13197,N_12925,N_12960);
nor U13198 (N_13198,N_12832,N_12864);
and U13199 (N_13199,N_12852,N_12907);
and U13200 (N_13200,N_13077,N_13087);
and U13201 (N_13201,N_13140,N_13106);
and U13202 (N_13202,N_13167,N_13161);
xnor U13203 (N_13203,N_13086,N_13107);
xor U13204 (N_13204,N_13160,N_13147);
or U13205 (N_13205,N_13164,N_13048);
or U13206 (N_13206,N_13036,N_13184);
or U13207 (N_13207,N_13119,N_13025);
xnor U13208 (N_13208,N_13121,N_13054);
nor U13209 (N_13209,N_13096,N_13033);
and U13210 (N_13210,N_13139,N_13020);
nor U13211 (N_13211,N_13064,N_13116);
nand U13212 (N_13212,N_13075,N_13098);
or U13213 (N_13213,N_13009,N_13059);
nand U13214 (N_13214,N_13056,N_13028);
nand U13215 (N_13215,N_13100,N_13132);
xor U13216 (N_13216,N_13127,N_13101);
and U13217 (N_13217,N_13170,N_13102);
nand U13218 (N_13218,N_13191,N_13148);
or U13219 (N_13219,N_13122,N_13030);
or U13220 (N_13220,N_13017,N_13003);
nand U13221 (N_13221,N_13179,N_13136);
or U13222 (N_13222,N_13112,N_13097);
or U13223 (N_13223,N_13111,N_13151);
and U13224 (N_13224,N_13195,N_13123);
or U13225 (N_13225,N_13149,N_13150);
xor U13226 (N_13226,N_13176,N_13006);
or U13227 (N_13227,N_13004,N_13031);
nand U13228 (N_13228,N_13072,N_13007);
or U13229 (N_13229,N_13157,N_13068);
xor U13230 (N_13230,N_13037,N_13042);
and U13231 (N_13231,N_13193,N_13019);
nor U13232 (N_13232,N_13070,N_13095);
and U13233 (N_13233,N_13115,N_13069);
nand U13234 (N_13234,N_13197,N_13051);
nand U13235 (N_13235,N_13002,N_13016);
and U13236 (N_13236,N_13171,N_13175);
or U13237 (N_13237,N_13000,N_13022);
and U13238 (N_13238,N_13074,N_13125);
nand U13239 (N_13239,N_13142,N_13135);
or U13240 (N_13240,N_13152,N_13049);
and U13241 (N_13241,N_13105,N_13084);
xnor U13242 (N_13242,N_13013,N_13034);
and U13243 (N_13243,N_13192,N_13108);
and U13244 (N_13244,N_13026,N_13081);
or U13245 (N_13245,N_13082,N_13154);
or U13246 (N_13246,N_13113,N_13126);
or U13247 (N_13247,N_13027,N_13010);
xor U13248 (N_13248,N_13090,N_13029);
nand U13249 (N_13249,N_13186,N_13089);
or U13250 (N_13250,N_13021,N_13146);
nor U13251 (N_13251,N_13177,N_13032);
nor U13252 (N_13252,N_13180,N_13188);
or U13253 (N_13253,N_13083,N_13093);
or U13254 (N_13254,N_13073,N_13050);
and U13255 (N_13255,N_13014,N_13061);
nand U13256 (N_13256,N_13045,N_13076);
or U13257 (N_13257,N_13196,N_13023);
or U13258 (N_13258,N_13066,N_13015);
and U13259 (N_13259,N_13174,N_13008);
and U13260 (N_13260,N_13162,N_13062);
and U13261 (N_13261,N_13118,N_13185);
and U13262 (N_13262,N_13156,N_13158);
nor U13263 (N_13263,N_13114,N_13005);
nor U13264 (N_13264,N_13078,N_13052);
xor U13265 (N_13265,N_13190,N_13138);
and U13266 (N_13266,N_13043,N_13166);
nand U13267 (N_13267,N_13039,N_13079);
and U13268 (N_13268,N_13131,N_13153);
nand U13269 (N_13269,N_13024,N_13058);
xnor U13270 (N_13270,N_13104,N_13094);
xnor U13271 (N_13271,N_13133,N_13109);
nand U13272 (N_13272,N_13053,N_13046);
and U13273 (N_13273,N_13194,N_13099);
and U13274 (N_13274,N_13044,N_13040);
nor U13275 (N_13275,N_13011,N_13041);
nor U13276 (N_13276,N_13199,N_13071);
and U13277 (N_13277,N_13141,N_13137);
nand U13278 (N_13278,N_13182,N_13143);
or U13279 (N_13279,N_13134,N_13088);
and U13280 (N_13280,N_13055,N_13155);
nor U13281 (N_13281,N_13001,N_13144);
nand U13282 (N_13282,N_13189,N_13165);
or U13283 (N_13283,N_13187,N_13063);
nand U13284 (N_13284,N_13173,N_13085);
and U13285 (N_13285,N_13035,N_13159);
nand U13286 (N_13286,N_13038,N_13047);
nor U13287 (N_13287,N_13128,N_13198);
nand U13288 (N_13288,N_13012,N_13065);
nand U13289 (N_13289,N_13057,N_13110);
and U13290 (N_13290,N_13145,N_13091);
and U13291 (N_13291,N_13120,N_13181);
and U13292 (N_13292,N_13169,N_13168);
nand U13293 (N_13293,N_13060,N_13183);
and U13294 (N_13294,N_13129,N_13103);
nor U13295 (N_13295,N_13018,N_13080);
nor U13296 (N_13296,N_13178,N_13117);
nand U13297 (N_13297,N_13124,N_13067);
and U13298 (N_13298,N_13172,N_13130);
xor U13299 (N_13299,N_13163,N_13092);
nor U13300 (N_13300,N_13089,N_13113);
nand U13301 (N_13301,N_13055,N_13149);
nor U13302 (N_13302,N_13023,N_13107);
xnor U13303 (N_13303,N_13083,N_13054);
and U13304 (N_13304,N_13133,N_13198);
nor U13305 (N_13305,N_13016,N_13147);
nor U13306 (N_13306,N_13138,N_13178);
and U13307 (N_13307,N_13015,N_13016);
nand U13308 (N_13308,N_13158,N_13022);
nand U13309 (N_13309,N_13032,N_13158);
and U13310 (N_13310,N_13138,N_13106);
nand U13311 (N_13311,N_13151,N_13022);
xnor U13312 (N_13312,N_13076,N_13182);
nor U13313 (N_13313,N_13031,N_13166);
or U13314 (N_13314,N_13091,N_13079);
or U13315 (N_13315,N_13196,N_13155);
nor U13316 (N_13316,N_13015,N_13134);
and U13317 (N_13317,N_13000,N_13112);
nand U13318 (N_13318,N_13049,N_13073);
and U13319 (N_13319,N_13161,N_13112);
and U13320 (N_13320,N_13167,N_13134);
and U13321 (N_13321,N_13088,N_13169);
nor U13322 (N_13322,N_13100,N_13033);
and U13323 (N_13323,N_13127,N_13199);
nand U13324 (N_13324,N_13197,N_13071);
nand U13325 (N_13325,N_13000,N_13156);
nor U13326 (N_13326,N_13076,N_13067);
nor U13327 (N_13327,N_13097,N_13061);
and U13328 (N_13328,N_13140,N_13150);
nor U13329 (N_13329,N_13092,N_13002);
xor U13330 (N_13330,N_13018,N_13176);
nand U13331 (N_13331,N_13032,N_13016);
and U13332 (N_13332,N_13061,N_13082);
and U13333 (N_13333,N_13030,N_13079);
or U13334 (N_13334,N_13046,N_13122);
nand U13335 (N_13335,N_13068,N_13011);
and U13336 (N_13336,N_13073,N_13186);
and U13337 (N_13337,N_13041,N_13107);
nand U13338 (N_13338,N_13059,N_13152);
xor U13339 (N_13339,N_13121,N_13177);
or U13340 (N_13340,N_13084,N_13037);
xor U13341 (N_13341,N_13011,N_13178);
nor U13342 (N_13342,N_13022,N_13119);
or U13343 (N_13343,N_13116,N_13136);
or U13344 (N_13344,N_13124,N_13135);
or U13345 (N_13345,N_13039,N_13042);
and U13346 (N_13346,N_13137,N_13036);
nand U13347 (N_13347,N_13180,N_13072);
or U13348 (N_13348,N_13197,N_13182);
nand U13349 (N_13349,N_13000,N_13036);
nor U13350 (N_13350,N_13180,N_13064);
and U13351 (N_13351,N_13141,N_13033);
nor U13352 (N_13352,N_13171,N_13063);
or U13353 (N_13353,N_13064,N_13104);
nor U13354 (N_13354,N_13102,N_13183);
nor U13355 (N_13355,N_13122,N_13025);
nor U13356 (N_13356,N_13118,N_13144);
or U13357 (N_13357,N_13028,N_13029);
and U13358 (N_13358,N_13022,N_13159);
and U13359 (N_13359,N_13038,N_13027);
nor U13360 (N_13360,N_13060,N_13031);
nand U13361 (N_13361,N_13024,N_13064);
nor U13362 (N_13362,N_13077,N_13053);
nand U13363 (N_13363,N_13189,N_13083);
or U13364 (N_13364,N_13066,N_13130);
nand U13365 (N_13365,N_13005,N_13007);
or U13366 (N_13366,N_13162,N_13130);
or U13367 (N_13367,N_13043,N_13091);
or U13368 (N_13368,N_13042,N_13112);
nand U13369 (N_13369,N_13027,N_13102);
nand U13370 (N_13370,N_13073,N_13030);
and U13371 (N_13371,N_13007,N_13020);
and U13372 (N_13372,N_13009,N_13062);
nand U13373 (N_13373,N_13147,N_13135);
or U13374 (N_13374,N_13186,N_13151);
nand U13375 (N_13375,N_13086,N_13084);
or U13376 (N_13376,N_13123,N_13141);
or U13377 (N_13377,N_13080,N_13185);
xnor U13378 (N_13378,N_13041,N_13199);
nand U13379 (N_13379,N_13054,N_13139);
and U13380 (N_13380,N_13191,N_13084);
xor U13381 (N_13381,N_13172,N_13167);
or U13382 (N_13382,N_13109,N_13092);
and U13383 (N_13383,N_13153,N_13095);
xor U13384 (N_13384,N_13183,N_13157);
and U13385 (N_13385,N_13089,N_13155);
nand U13386 (N_13386,N_13102,N_13094);
nor U13387 (N_13387,N_13054,N_13184);
or U13388 (N_13388,N_13024,N_13177);
nor U13389 (N_13389,N_13067,N_13162);
nand U13390 (N_13390,N_13142,N_13132);
xnor U13391 (N_13391,N_13147,N_13010);
or U13392 (N_13392,N_13067,N_13084);
or U13393 (N_13393,N_13199,N_13192);
nor U13394 (N_13394,N_13067,N_13029);
nand U13395 (N_13395,N_13073,N_13017);
nor U13396 (N_13396,N_13016,N_13189);
or U13397 (N_13397,N_13185,N_13138);
and U13398 (N_13398,N_13058,N_13134);
or U13399 (N_13399,N_13143,N_13181);
and U13400 (N_13400,N_13338,N_13381);
and U13401 (N_13401,N_13232,N_13330);
nand U13402 (N_13402,N_13393,N_13342);
nor U13403 (N_13403,N_13269,N_13335);
nand U13404 (N_13404,N_13340,N_13222);
xor U13405 (N_13405,N_13253,N_13270);
nor U13406 (N_13406,N_13395,N_13271);
nand U13407 (N_13407,N_13392,N_13208);
or U13408 (N_13408,N_13298,N_13220);
nor U13409 (N_13409,N_13239,N_13315);
and U13410 (N_13410,N_13390,N_13313);
nor U13411 (N_13411,N_13397,N_13287);
nand U13412 (N_13412,N_13305,N_13260);
nor U13413 (N_13413,N_13375,N_13245);
nor U13414 (N_13414,N_13265,N_13310);
and U13415 (N_13415,N_13295,N_13250);
nor U13416 (N_13416,N_13333,N_13227);
nand U13417 (N_13417,N_13344,N_13299);
nor U13418 (N_13418,N_13230,N_13215);
xnor U13419 (N_13419,N_13296,N_13293);
nor U13420 (N_13420,N_13329,N_13307);
nor U13421 (N_13421,N_13206,N_13274);
xnor U13422 (N_13422,N_13308,N_13289);
xnor U13423 (N_13423,N_13384,N_13218);
and U13424 (N_13424,N_13263,N_13272);
or U13425 (N_13425,N_13280,N_13292);
xnor U13426 (N_13426,N_13261,N_13337);
xor U13427 (N_13427,N_13216,N_13377);
and U13428 (N_13428,N_13275,N_13366);
nand U13429 (N_13429,N_13279,N_13318);
or U13430 (N_13430,N_13290,N_13378);
or U13431 (N_13431,N_13389,N_13256);
or U13432 (N_13432,N_13352,N_13251);
or U13433 (N_13433,N_13359,N_13383);
or U13434 (N_13434,N_13210,N_13213);
and U13435 (N_13435,N_13309,N_13328);
or U13436 (N_13436,N_13300,N_13234);
and U13437 (N_13437,N_13365,N_13268);
xnor U13438 (N_13438,N_13396,N_13224);
and U13439 (N_13439,N_13354,N_13254);
or U13440 (N_13440,N_13368,N_13212);
nor U13441 (N_13441,N_13353,N_13398);
nor U13442 (N_13442,N_13262,N_13363);
or U13443 (N_13443,N_13372,N_13355);
and U13444 (N_13444,N_13219,N_13200);
nor U13445 (N_13445,N_13399,N_13282);
nor U13446 (N_13446,N_13229,N_13369);
or U13447 (N_13447,N_13386,N_13209);
or U13448 (N_13448,N_13350,N_13336);
and U13449 (N_13449,N_13345,N_13346);
nor U13450 (N_13450,N_13370,N_13217);
nand U13451 (N_13451,N_13285,N_13388);
nand U13452 (N_13452,N_13273,N_13228);
nor U13453 (N_13453,N_13325,N_13348);
or U13454 (N_13454,N_13214,N_13225);
and U13455 (N_13455,N_13276,N_13321);
and U13456 (N_13456,N_13294,N_13376);
nand U13457 (N_13457,N_13252,N_13238);
and U13458 (N_13458,N_13326,N_13231);
xnor U13459 (N_13459,N_13266,N_13284);
xnor U13460 (N_13460,N_13316,N_13205);
nand U13461 (N_13461,N_13255,N_13259);
and U13462 (N_13462,N_13235,N_13286);
nor U13463 (N_13463,N_13391,N_13242);
or U13464 (N_13464,N_13358,N_13324);
xor U13465 (N_13465,N_13360,N_13297);
and U13466 (N_13466,N_13247,N_13322);
xor U13467 (N_13467,N_13201,N_13323);
or U13468 (N_13468,N_13211,N_13204);
or U13469 (N_13469,N_13226,N_13221);
nand U13470 (N_13470,N_13278,N_13382);
xor U13471 (N_13471,N_13237,N_13306);
or U13472 (N_13472,N_13267,N_13302);
and U13473 (N_13473,N_13240,N_13332);
nor U13474 (N_13474,N_13233,N_13347);
nand U13475 (N_13475,N_13202,N_13277);
and U13476 (N_13476,N_13320,N_13367);
nand U13477 (N_13477,N_13258,N_13246);
xor U13478 (N_13478,N_13357,N_13394);
nor U13479 (N_13479,N_13361,N_13351);
nand U13480 (N_13480,N_13349,N_13303);
xor U13481 (N_13481,N_13203,N_13314);
nand U13482 (N_13482,N_13281,N_13223);
nand U13483 (N_13483,N_13331,N_13385);
or U13484 (N_13484,N_13243,N_13207);
nor U13485 (N_13485,N_13356,N_13249);
nand U13486 (N_13486,N_13374,N_13317);
and U13487 (N_13487,N_13364,N_13291);
xor U13488 (N_13488,N_13373,N_13311);
and U13489 (N_13489,N_13327,N_13380);
nor U13490 (N_13490,N_13248,N_13339);
and U13491 (N_13491,N_13288,N_13244);
nand U13492 (N_13492,N_13236,N_13283);
or U13493 (N_13493,N_13312,N_13301);
nand U13494 (N_13494,N_13387,N_13334);
or U13495 (N_13495,N_13257,N_13343);
or U13496 (N_13496,N_13319,N_13379);
nor U13497 (N_13497,N_13264,N_13241);
nand U13498 (N_13498,N_13341,N_13304);
nor U13499 (N_13499,N_13362,N_13371);
or U13500 (N_13500,N_13363,N_13214);
or U13501 (N_13501,N_13242,N_13363);
nand U13502 (N_13502,N_13316,N_13229);
nor U13503 (N_13503,N_13301,N_13303);
xnor U13504 (N_13504,N_13274,N_13301);
or U13505 (N_13505,N_13330,N_13218);
nand U13506 (N_13506,N_13267,N_13200);
and U13507 (N_13507,N_13276,N_13358);
xor U13508 (N_13508,N_13323,N_13328);
or U13509 (N_13509,N_13397,N_13291);
and U13510 (N_13510,N_13226,N_13399);
nor U13511 (N_13511,N_13322,N_13375);
nand U13512 (N_13512,N_13392,N_13316);
nor U13513 (N_13513,N_13363,N_13265);
or U13514 (N_13514,N_13370,N_13266);
or U13515 (N_13515,N_13350,N_13319);
or U13516 (N_13516,N_13292,N_13397);
nor U13517 (N_13517,N_13380,N_13210);
nor U13518 (N_13518,N_13341,N_13328);
nor U13519 (N_13519,N_13360,N_13334);
or U13520 (N_13520,N_13275,N_13208);
nand U13521 (N_13521,N_13299,N_13291);
nand U13522 (N_13522,N_13395,N_13397);
and U13523 (N_13523,N_13236,N_13354);
or U13524 (N_13524,N_13205,N_13221);
and U13525 (N_13525,N_13290,N_13358);
or U13526 (N_13526,N_13367,N_13298);
nand U13527 (N_13527,N_13313,N_13289);
or U13528 (N_13528,N_13204,N_13288);
or U13529 (N_13529,N_13346,N_13261);
nor U13530 (N_13530,N_13386,N_13325);
nor U13531 (N_13531,N_13349,N_13304);
nand U13532 (N_13532,N_13345,N_13205);
and U13533 (N_13533,N_13222,N_13361);
or U13534 (N_13534,N_13232,N_13274);
and U13535 (N_13535,N_13396,N_13210);
nand U13536 (N_13536,N_13227,N_13374);
xnor U13537 (N_13537,N_13354,N_13239);
nand U13538 (N_13538,N_13220,N_13228);
or U13539 (N_13539,N_13388,N_13385);
nand U13540 (N_13540,N_13226,N_13211);
nor U13541 (N_13541,N_13318,N_13275);
and U13542 (N_13542,N_13210,N_13378);
and U13543 (N_13543,N_13201,N_13293);
nand U13544 (N_13544,N_13271,N_13386);
and U13545 (N_13545,N_13274,N_13287);
nand U13546 (N_13546,N_13376,N_13388);
and U13547 (N_13547,N_13222,N_13238);
and U13548 (N_13548,N_13296,N_13233);
xor U13549 (N_13549,N_13313,N_13387);
nor U13550 (N_13550,N_13243,N_13310);
nand U13551 (N_13551,N_13228,N_13301);
and U13552 (N_13552,N_13288,N_13245);
nor U13553 (N_13553,N_13282,N_13248);
xnor U13554 (N_13554,N_13384,N_13246);
and U13555 (N_13555,N_13327,N_13390);
nor U13556 (N_13556,N_13258,N_13298);
nand U13557 (N_13557,N_13282,N_13229);
or U13558 (N_13558,N_13305,N_13367);
nand U13559 (N_13559,N_13314,N_13346);
nand U13560 (N_13560,N_13333,N_13305);
nand U13561 (N_13561,N_13228,N_13308);
nand U13562 (N_13562,N_13233,N_13256);
and U13563 (N_13563,N_13241,N_13239);
nand U13564 (N_13564,N_13397,N_13374);
and U13565 (N_13565,N_13334,N_13226);
nand U13566 (N_13566,N_13341,N_13298);
and U13567 (N_13567,N_13297,N_13259);
nand U13568 (N_13568,N_13239,N_13249);
nor U13569 (N_13569,N_13242,N_13370);
or U13570 (N_13570,N_13284,N_13293);
or U13571 (N_13571,N_13333,N_13313);
and U13572 (N_13572,N_13272,N_13216);
nor U13573 (N_13573,N_13337,N_13349);
nor U13574 (N_13574,N_13394,N_13243);
or U13575 (N_13575,N_13376,N_13281);
nand U13576 (N_13576,N_13381,N_13305);
and U13577 (N_13577,N_13280,N_13282);
or U13578 (N_13578,N_13342,N_13212);
or U13579 (N_13579,N_13384,N_13232);
nand U13580 (N_13580,N_13368,N_13397);
or U13581 (N_13581,N_13214,N_13397);
nor U13582 (N_13582,N_13391,N_13234);
nand U13583 (N_13583,N_13235,N_13340);
and U13584 (N_13584,N_13245,N_13392);
or U13585 (N_13585,N_13295,N_13259);
nor U13586 (N_13586,N_13264,N_13287);
nand U13587 (N_13587,N_13303,N_13309);
and U13588 (N_13588,N_13266,N_13335);
nor U13589 (N_13589,N_13298,N_13304);
xnor U13590 (N_13590,N_13216,N_13288);
xor U13591 (N_13591,N_13206,N_13271);
xnor U13592 (N_13592,N_13219,N_13255);
nand U13593 (N_13593,N_13369,N_13368);
nand U13594 (N_13594,N_13393,N_13380);
nor U13595 (N_13595,N_13292,N_13329);
nor U13596 (N_13596,N_13331,N_13343);
nand U13597 (N_13597,N_13272,N_13321);
nand U13598 (N_13598,N_13222,N_13369);
xor U13599 (N_13599,N_13201,N_13254);
nor U13600 (N_13600,N_13480,N_13577);
or U13601 (N_13601,N_13400,N_13567);
or U13602 (N_13602,N_13563,N_13465);
nand U13603 (N_13603,N_13481,N_13452);
and U13604 (N_13604,N_13502,N_13471);
or U13605 (N_13605,N_13537,N_13512);
nand U13606 (N_13606,N_13441,N_13503);
nand U13607 (N_13607,N_13489,N_13504);
and U13608 (N_13608,N_13597,N_13491);
or U13609 (N_13609,N_13490,N_13442);
and U13610 (N_13610,N_13543,N_13520);
nand U13611 (N_13611,N_13409,N_13429);
and U13612 (N_13612,N_13474,N_13595);
or U13613 (N_13613,N_13405,N_13403);
and U13614 (N_13614,N_13410,N_13433);
nor U13615 (N_13615,N_13517,N_13562);
nand U13616 (N_13616,N_13523,N_13586);
nor U13617 (N_13617,N_13402,N_13440);
nand U13618 (N_13618,N_13580,N_13588);
xnor U13619 (N_13619,N_13482,N_13487);
nor U13620 (N_13620,N_13421,N_13492);
nor U13621 (N_13621,N_13579,N_13498);
or U13622 (N_13622,N_13493,N_13591);
xor U13623 (N_13623,N_13509,N_13594);
nand U13624 (N_13624,N_13553,N_13547);
or U13625 (N_13625,N_13404,N_13443);
nor U13626 (N_13626,N_13526,N_13420);
xor U13627 (N_13627,N_13436,N_13448);
or U13628 (N_13628,N_13434,N_13450);
nor U13629 (N_13629,N_13497,N_13447);
nor U13630 (N_13630,N_13554,N_13499);
and U13631 (N_13631,N_13593,N_13453);
nand U13632 (N_13632,N_13483,N_13590);
nor U13633 (N_13633,N_13510,N_13406);
and U13634 (N_13634,N_13576,N_13524);
and U13635 (N_13635,N_13539,N_13521);
nand U13636 (N_13636,N_13559,N_13513);
nand U13637 (N_13637,N_13444,N_13438);
nand U13638 (N_13638,N_13564,N_13578);
nor U13639 (N_13639,N_13519,N_13467);
nand U13640 (N_13640,N_13466,N_13449);
xor U13641 (N_13641,N_13476,N_13459);
xor U13642 (N_13642,N_13548,N_13516);
and U13643 (N_13643,N_13460,N_13424);
or U13644 (N_13644,N_13583,N_13506);
nor U13645 (N_13645,N_13592,N_13430);
or U13646 (N_13646,N_13435,N_13589);
and U13647 (N_13647,N_13418,N_13461);
nand U13648 (N_13648,N_13536,N_13426);
and U13649 (N_13649,N_13570,N_13598);
nand U13650 (N_13650,N_13571,N_13557);
or U13651 (N_13651,N_13488,N_13596);
xnor U13652 (N_13652,N_13556,N_13525);
nand U13653 (N_13653,N_13468,N_13412);
nor U13654 (N_13654,N_13538,N_13462);
and U13655 (N_13655,N_13451,N_13561);
or U13656 (N_13656,N_13582,N_13584);
or U13657 (N_13657,N_13500,N_13549);
nor U13658 (N_13658,N_13533,N_13469);
and U13659 (N_13659,N_13425,N_13565);
nand U13660 (N_13660,N_13495,N_13475);
nand U13661 (N_13661,N_13535,N_13446);
xnor U13662 (N_13662,N_13585,N_13531);
or U13663 (N_13663,N_13530,N_13457);
and U13664 (N_13664,N_13454,N_13514);
or U13665 (N_13665,N_13401,N_13477);
or U13666 (N_13666,N_13463,N_13542);
nor U13667 (N_13667,N_13507,N_13464);
nand U13668 (N_13668,N_13522,N_13540);
and U13669 (N_13669,N_13573,N_13574);
nand U13670 (N_13670,N_13431,N_13416);
or U13671 (N_13671,N_13422,N_13550);
nand U13672 (N_13672,N_13528,N_13445);
xnor U13673 (N_13673,N_13575,N_13437);
or U13674 (N_13674,N_13432,N_13413);
nand U13675 (N_13675,N_13566,N_13439);
nor U13676 (N_13676,N_13532,N_13423);
and U13677 (N_13677,N_13545,N_13534);
xor U13678 (N_13678,N_13546,N_13552);
and U13679 (N_13679,N_13496,N_13414);
nand U13680 (N_13680,N_13455,N_13558);
nor U13681 (N_13681,N_13470,N_13473);
and U13682 (N_13682,N_13544,N_13485);
and U13683 (N_13683,N_13551,N_13415);
xnor U13684 (N_13684,N_13560,N_13427);
and U13685 (N_13685,N_13508,N_13456);
and U13686 (N_13686,N_13458,N_13472);
nand U13687 (N_13687,N_13518,N_13555);
and U13688 (N_13688,N_13494,N_13484);
and U13689 (N_13689,N_13411,N_13501);
and U13690 (N_13690,N_13417,N_13581);
or U13691 (N_13691,N_13428,N_13529);
nor U13692 (N_13692,N_13599,N_13527);
and U13693 (N_13693,N_13515,N_13505);
nand U13694 (N_13694,N_13587,N_13541);
nand U13695 (N_13695,N_13486,N_13407);
nand U13696 (N_13696,N_13408,N_13569);
nor U13697 (N_13697,N_13568,N_13479);
nand U13698 (N_13698,N_13478,N_13572);
and U13699 (N_13699,N_13419,N_13511);
or U13700 (N_13700,N_13525,N_13550);
nand U13701 (N_13701,N_13544,N_13570);
or U13702 (N_13702,N_13566,N_13508);
or U13703 (N_13703,N_13590,N_13564);
nand U13704 (N_13704,N_13543,N_13550);
and U13705 (N_13705,N_13523,N_13580);
and U13706 (N_13706,N_13563,N_13572);
xor U13707 (N_13707,N_13490,N_13463);
xor U13708 (N_13708,N_13427,N_13528);
nand U13709 (N_13709,N_13411,N_13520);
nor U13710 (N_13710,N_13551,N_13573);
and U13711 (N_13711,N_13565,N_13518);
and U13712 (N_13712,N_13461,N_13430);
and U13713 (N_13713,N_13415,N_13594);
nor U13714 (N_13714,N_13594,N_13478);
and U13715 (N_13715,N_13549,N_13535);
and U13716 (N_13716,N_13424,N_13438);
nor U13717 (N_13717,N_13572,N_13596);
nand U13718 (N_13718,N_13558,N_13493);
or U13719 (N_13719,N_13557,N_13521);
nand U13720 (N_13720,N_13508,N_13550);
nor U13721 (N_13721,N_13567,N_13492);
or U13722 (N_13722,N_13445,N_13475);
or U13723 (N_13723,N_13526,N_13400);
nand U13724 (N_13724,N_13579,N_13581);
and U13725 (N_13725,N_13552,N_13443);
or U13726 (N_13726,N_13580,N_13568);
and U13727 (N_13727,N_13500,N_13458);
or U13728 (N_13728,N_13504,N_13525);
or U13729 (N_13729,N_13461,N_13476);
and U13730 (N_13730,N_13440,N_13523);
nand U13731 (N_13731,N_13495,N_13443);
or U13732 (N_13732,N_13527,N_13408);
and U13733 (N_13733,N_13514,N_13463);
and U13734 (N_13734,N_13478,N_13495);
and U13735 (N_13735,N_13544,N_13459);
or U13736 (N_13736,N_13572,N_13420);
or U13737 (N_13737,N_13443,N_13531);
nor U13738 (N_13738,N_13403,N_13457);
and U13739 (N_13739,N_13507,N_13519);
or U13740 (N_13740,N_13546,N_13507);
nor U13741 (N_13741,N_13524,N_13411);
or U13742 (N_13742,N_13501,N_13400);
or U13743 (N_13743,N_13554,N_13514);
nand U13744 (N_13744,N_13463,N_13568);
nand U13745 (N_13745,N_13437,N_13588);
or U13746 (N_13746,N_13468,N_13528);
nand U13747 (N_13747,N_13555,N_13560);
or U13748 (N_13748,N_13500,N_13401);
or U13749 (N_13749,N_13500,N_13463);
nand U13750 (N_13750,N_13515,N_13420);
nor U13751 (N_13751,N_13509,N_13512);
nand U13752 (N_13752,N_13437,N_13514);
nor U13753 (N_13753,N_13598,N_13475);
and U13754 (N_13754,N_13435,N_13405);
nand U13755 (N_13755,N_13410,N_13485);
xor U13756 (N_13756,N_13450,N_13543);
xor U13757 (N_13757,N_13403,N_13538);
and U13758 (N_13758,N_13551,N_13599);
and U13759 (N_13759,N_13459,N_13549);
nand U13760 (N_13760,N_13540,N_13544);
nand U13761 (N_13761,N_13506,N_13454);
nor U13762 (N_13762,N_13430,N_13409);
and U13763 (N_13763,N_13511,N_13595);
and U13764 (N_13764,N_13532,N_13564);
or U13765 (N_13765,N_13486,N_13556);
nor U13766 (N_13766,N_13585,N_13487);
nor U13767 (N_13767,N_13496,N_13436);
nor U13768 (N_13768,N_13463,N_13449);
and U13769 (N_13769,N_13458,N_13488);
nor U13770 (N_13770,N_13417,N_13505);
nor U13771 (N_13771,N_13548,N_13406);
nand U13772 (N_13772,N_13463,N_13570);
nand U13773 (N_13773,N_13575,N_13566);
nand U13774 (N_13774,N_13558,N_13547);
or U13775 (N_13775,N_13464,N_13499);
nand U13776 (N_13776,N_13570,N_13430);
or U13777 (N_13777,N_13401,N_13536);
and U13778 (N_13778,N_13599,N_13572);
nand U13779 (N_13779,N_13415,N_13533);
nand U13780 (N_13780,N_13446,N_13586);
or U13781 (N_13781,N_13578,N_13520);
xor U13782 (N_13782,N_13441,N_13584);
xor U13783 (N_13783,N_13583,N_13586);
and U13784 (N_13784,N_13547,N_13541);
or U13785 (N_13785,N_13597,N_13530);
nor U13786 (N_13786,N_13401,N_13556);
and U13787 (N_13787,N_13495,N_13427);
and U13788 (N_13788,N_13417,N_13504);
nand U13789 (N_13789,N_13554,N_13540);
xor U13790 (N_13790,N_13418,N_13582);
nor U13791 (N_13791,N_13413,N_13489);
or U13792 (N_13792,N_13456,N_13416);
or U13793 (N_13793,N_13504,N_13410);
nand U13794 (N_13794,N_13530,N_13598);
nor U13795 (N_13795,N_13561,N_13569);
or U13796 (N_13796,N_13590,N_13490);
and U13797 (N_13797,N_13466,N_13533);
and U13798 (N_13798,N_13434,N_13497);
and U13799 (N_13799,N_13517,N_13463);
nand U13800 (N_13800,N_13768,N_13675);
xnor U13801 (N_13801,N_13780,N_13747);
nand U13802 (N_13802,N_13659,N_13703);
nor U13803 (N_13803,N_13712,N_13602);
nand U13804 (N_13804,N_13706,N_13762);
and U13805 (N_13805,N_13689,N_13621);
nor U13806 (N_13806,N_13651,N_13781);
nand U13807 (N_13807,N_13797,N_13707);
nand U13808 (N_13808,N_13719,N_13615);
nor U13809 (N_13809,N_13711,N_13656);
nand U13810 (N_13810,N_13616,N_13605);
nand U13811 (N_13811,N_13695,N_13640);
nand U13812 (N_13812,N_13697,N_13693);
nand U13813 (N_13813,N_13754,N_13676);
nor U13814 (N_13814,N_13738,N_13677);
or U13815 (N_13815,N_13700,N_13641);
nand U13816 (N_13816,N_13679,N_13652);
and U13817 (N_13817,N_13773,N_13649);
or U13818 (N_13818,N_13756,N_13708);
and U13819 (N_13819,N_13654,N_13715);
or U13820 (N_13820,N_13767,N_13776);
or U13821 (N_13821,N_13786,N_13655);
nor U13822 (N_13822,N_13682,N_13774);
nor U13823 (N_13823,N_13729,N_13643);
nor U13824 (N_13824,N_13753,N_13704);
or U13825 (N_13825,N_13670,N_13680);
and U13826 (N_13826,N_13720,N_13751);
and U13827 (N_13827,N_13765,N_13785);
and U13828 (N_13828,N_13645,N_13789);
nor U13829 (N_13829,N_13790,N_13600);
nand U13830 (N_13830,N_13736,N_13716);
and U13831 (N_13831,N_13604,N_13788);
nand U13832 (N_13832,N_13687,N_13690);
xnor U13833 (N_13833,N_13783,N_13717);
xnor U13834 (N_13834,N_13726,N_13694);
xnor U13835 (N_13835,N_13669,N_13723);
xor U13836 (N_13836,N_13667,N_13761);
nor U13837 (N_13837,N_13784,N_13671);
or U13838 (N_13838,N_13743,N_13763);
and U13839 (N_13839,N_13623,N_13793);
and U13840 (N_13840,N_13684,N_13627);
nor U13841 (N_13841,N_13660,N_13779);
or U13842 (N_13842,N_13744,N_13755);
nand U13843 (N_13843,N_13666,N_13759);
nand U13844 (N_13844,N_13688,N_13624);
or U13845 (N_13845,N_13618,N_13725);
nand U13846 (N_13846,N_13610,N_13657);
and U13847 (N_13847,N_13639,N_13798);
or U13848 (N_13848,N_13737,N_13620);
or U13849 (N_13849,N_13668,N_13638);
or U13850 (N_13850,N_13609,N_13607);
nand U13851 (N_13851,N_13702,N_13733);
nand U13852 (N_13852,N_13672,N_13746);
and U13853 (N_13853,N_13709,N_13752);
nor U13854 (N_13854,N_13792,N_13614);
or U13855 (N_13855,N_13772,N_13778);
and U13856 (N_13856,N_13777,N_13705);
nand U13857 (N_13857,N_13757,N_13769);
nor U13858 (N_13858,N_13748,N_13644);
nand U13859 (N_13859,N_13612,N_13724);
and U13860 (N_13860,N_13760,N_13745);
and U13861 (N_13861,N_13633,N_13673);
nand U13862 (N_13862,N_13625,N_13735);
or U13863 (N_13863,N_13750,N_13661);
or U13864 (N_13864,N_13713,N_13611);
or U13865 (N_13865,N_13642,N_13739);
nor U13866 (N_13866,N_13650,N_13758);
nand U13867 (N_13867,N_13663,N_13692);
and U13868 (N_13868,N_13795,N_13617);
nor U13869 (N_13869,N_13636,N_13791);
and U13870 (N_13870,N_13603,N_13648);
and U13871 (N_13871,N_13727,N_13787);
nor U13872 (N_13872,N_13698,N_13678);
nand U13873 (N_13873,N_13782,N_13630);
and U13874 (N_13874,N_13731,N_13658);
xnor U13875 (N_13875,N_13699,N_13628);
nor U13876 (N_13876,N_13665,N_13646);
nor U13877 (N_13877,N_13771,N_13629);
nand U13878 (N_13878,N_13732,N_13686);
nand U13879 (N_13879,N_13696,N_13613);
xor U13880 (N_13880,N_13742,N_13601);
or U13881 (N_13881,N_13794,N_13647);
nor U13882 (N_13882,N_13691,N_13775);
nor U13883 (N_13883,N_13722,N_13674);
xor U13884 (N_13884,N_13749,N_13740);
and U13885 (N_13885,N_13764,N_13766);
nand U13886 (N_13886,N_13710,N_13632);
nor U13887 (N_13887,N_13701,N_13664);
xnor U13888 (N_13888,N_13662,N_13606);
nand U13889 (N_13889,N_13626,N_13681);
nor U13890 (N_13890,N_13653,N_13622);
and U13891 (N_13891,N_13714,N_13637);
nor U13892 (N_13892,N_13728,N_13718);
and U13893 (N_13893,N_13796,N_13608);
nand U13894 (N_13894,N_13619,N_13685);
or U13895 (N_13895,N_13799,N_13730);
and U13896 (N_13896,N_13635,N_13634);
xor U13897 (N_13897,N_13734,N_13721);
or U13898 (N_13898,N_13741,N_13770);
nand U13899 (N_13899,N_13631,N_13683);
or U13900 (N_13900,N_13786,N_13727);
or U13901 (N_13901,N_13797,N_13786);
or U13902 (N_13902,N_13685,N_13730);
nand U13903 (N_13903,N_13607,N_13764);
and U13904 (N_13904,N_13616,N_13740);
or U13905 (N_13905,N_13753,N_13662);
nand U13906 (N_13906,N_13624,N_13722);
and U13907 (N_13907,N_13759,N_13799);
or U13908 (N_13908,N_13600,N_13711);
and U13909 (N_13909,N_13652,N_13671);
nand U13910 (N_13910,N_13620,N_13765);
and U13911 (N_13911,N_13679,N_13727);
and U13912 (N_13912,N_13771,N_13622);
nor U13913 (N_13913,N_13746,N_13615);
nand U13914 (N_13914,N_13717,N_13681);
and U13915 (N_13915,N_13788,N_13791);
or U13916 (N_13916,N_13746,N_13750);
xnor U13917 (N_13917,N_13789,N_13608);
nand U13918 (N_13918,N_13793,N_13786);
nor U13919 (N_13919,N_13617,N_13773);
and U13920 (N_13920,N_13611,N_13736);
nor U13921 (N_13921,N_13683,N_13655);
nand U13922 (N_13922,N_13603,N_13754);
nand U13923 (N_13923,N_13759,N_13697);
nor U13924 (N_13924,N_13654,N_13716);
nor U13925 (N_13925,N_13759,N_13764);
nor U13926 (N_13926,N_13624,N_13711);
or U13927 (N_13927,N_13795,N_13681);
and U13928 (N_13928,N_13700,N_13682);
nand U13929 (N_13929,N_13636,N_13705);
xor U13930 (N_13930,N_13767,N_13606);
xnor U13931 (N_13931,N_13627,N_13643);
xnor U13932 (N_13932,N_13615,N_13652);
nor U13933 (N_13933,N_13732,N_13601);
and U13934 (N_13934,N_13712,N_13670);
or U13935 (N_13935,N_13658,N_13672);
nand U13936 (N_13936,N_13656,N_13792);
nand U13937 (N_13937,N_13760,N_13798);
nand U13938 (N_13938,N_13637,N_13780);
or U13939 (N_13939,N_13645,N_13611);
nor U13940 (N_13940,N_13674,N_13602);
or U13941 (N_13941,N_13705,N_13794);
and U13942 (N_13942,N_13700,N_13720);
nand U13943 (N_13943,N_13729,N_13629);
nand U13944 (N_13944,N_13764,N_13722);
xor U13945 (N_13945,N_13767,N_13729);
and U13946 (N_13946,N_13636,N_13641);
nand U13947 (N_13947,N_13613,N_13624);
nand U13948 (N_13948,N_13646,N_13638);
or U13949 (N_13949,N_13743,N_13637);
xor U13950 (N_13950,N_13778,N_13650);
nand U13951 (N_13951,N_13706,N_13704);
nor U13952 (N_13952,N_13690,N_13768);
nor U13953 (N_13953,N_13674,N_13734);
or U13954 (N_13954,N_13777,N_13640);
and U13955 (N_13955,N_13687,N_13715);
nor U13956 (N_13956,N_13698,N_13712);
nor U13957 (N_13957,N_13741,N_13785);
nand U13958 (N_13958,N_13698,N_13746);
nand U13959 (N_13959,N_13663,N_13742);
nor U13960 (N_13960,N_13757,N_13610);
and U13961 (N_13961,N_13799,N_13762);
nand U13962 (N_13962,N_13782,N_13729);
and U13963 (N_13963,N_13778,N_13689);
or U13964 (N_13964,N_13681,N_13738);
nor U13965 (N_13965,N_13659,N_13681);
nor U13966 (N_13966,N_13608,N_13618);
nor U13967 (N_13967,N_13607,N_13665);
nand U13968 (N_13968,N_13709,N_13604);
nor U13969 (N_13969,N_13706,N_13660);
and U13970 (N_13970,N_13610,N_13747);
or U13971 (N_13971,N_13624,N_13731);
or U13972 (N_13972,N_13747,N_13635);
nand U13973 (N_13973,N_13710,N_13695);
or U13974 (N_13974,N_13797,N_13782);
and U13975 (N_13975,N_13782,N_13614);
or U13976 (N_13976,N_13739,N_13620);
nor U13977 (N_13977,N_13722,N_13751);
or U13978 (N_13978,N_13691,N_13601);
xor U13979 (N_13979,N_13693,N_13641);
nand U13980 (N_13980,N_13641,N_13618);
and U13981 (N_13981,N_13763,N_13631);
or U13982 (N_13982,N_13799,N_13795);
or U13983 (N_13983,N_13694,N_13628);
nand U13984 (N_13984,N_13650,N_13611);
xor U13985 (N_13985,N_13761,N_13607);
nand U13986 (N_13986,N_13730,N_13768);
and U13987 (N_13987,N_13780,N_13618);
nor U13988 (N_13988,N_13798,N_13771);
nor U13989 (N_13989,N_13710,N_13788);
and U13990 (N_13990,N_13724,N_13632);
nand U13991 (N_13991,N_13716,N_13668);
and U13992 (N_13992,N_13715,N_13635);
and U13993 (N_13993,N_13698,N_13737);
and U13994 (N_13994,N_13791,N_13794);
or U13995 (N_13995,N_13637,N_13695);
or U13996 (N_13996,N_13779,N_13639);
and U13997 (N_13997,N_13662,N_13768);
nor U13998 (N_13998,N_13704,N_13655);
nand U13999 (N_13999,N_13674,N_13708);
nand U14000 (N_14000,N_13972,N_13945);
nor U14001 (N_14001,N_13971,N_13915);
and U14002 (N_14002,N_13892,N_13897);
xnor U14003 (N_14003,N_13988,N_13855);
or U14004 (N_14004,N_13916,N_13837);
or U14005 (N_14005,N_13808,N_13857);
nand U14006 (N_14006,N_13999,N_13849);
nor U14007 (N_14007,N_13978,N_13856);
nor U14008 (N_14008,N_13844,N_13828);
nand U14009 (N_14009,N_13974,N_13902);
nor U14010 (N_14010,N_13879,N_13961);
nand U14011 (N_14011,N_13968,N_13917);
nand U14012 (N_14012,N_13838,N_13913);
or U14013 (N_14013,N_13829,N_13835);
and U14014 (N_14014,N_13967,N_13993);
and U14015 (N_14015,N_13951,N_13994);
or U14016 (N_14016,N_13890,N_13943);
nor U14017 (N_14017,N_13919,N_13927);
or U14018 (N_14018,N_13990,N_13893);
nor U14019 (N_14019,N_13870,N_13823);
xnor U14020 (N_14020,N_13941,N_13956);
and U14021 (N_14021,N_13886,N_13960);
and U14022 (N_14022,N_13975,N_13981);
nand U14023 (N_14023,N_13965,N_13964);
and U14024 (N_14024,N_13803,N_13819);
nand U14025 (N_14025,N_13843,N_13959);
nor U14026 (N_14026,N_13818,N_13806);
nor U14027 (N_14027,N_13896,N_13992);
and U14028 (N_14028,N_13839,N_13942);
xor U14029 (N_14029,N_13813,N_13987);
nor U14030 (N_14030,N_13833,N_13810);
nand U14031 (N_14031,N_13832,N_13875);
and U14032 (N_14032,N_13904,N_13957);
nand U14033 (N_14033,N_13908,N_13841);
xor U14034 (N_14034,N_13977,N_13934);
xor U14035 (N_14035,N_13817,N_13858);
or U14036 (N_14036,N_13936,N_13851);
and U14037 (N_14037,N_13926,N_13871);
or U14038 (N_14038,N_13863,N_13885);
nor U14039 (N_14039,N_13912,N_13937);
nor U14040 (N_14040,N_13903,N_13814);
nand U14041 (N_14041,N_13888,N_13962);
nand U14042 (N_14042,N_13931,N_13824);
or U14043 (N_14043,N_13869,N_13900);
nand U14044 (N_14044,N_13920,N_13939);
xor U14045 (N_14045,N_13815,N_13947);
xnor U14046 (N_14046,N_13980,N_13949);
nand U14047 (N_14047,N_13963,N_13830);
xnor U14048 (N_14048,N_13929,N_13985);
xnor U14049 (N_14049,N_13802,N_13880);
nand U14050 (N_14050,N_13807,N_13848);
nor U14051 (N_14051,N_13969,N_13840);
nor U14052 (N_14052,N_13878,N_13846);
or U14053 (N_14053,N_13928,N_13862);
or U14054 (N_14054,N_13921,N_13935);
nor U14055 (N_14055,N_13914,N_13860);
nor U14056 (N_14056,N_13873,N_13909);
or U14057 (N_14057,N_13997,N_13811);
xnor U14058 (N_14058,N_13989,N_13991);
nand U14059 (N_14059,N_13982,N_13874);
nand U14060 (N_14060,N_13923,N_13865);
nand U14061 (N_14061,N_13867,N_13852);
nand U14062 (N_14062,N_13933,N_13922);
nor U14063 (N_14063,N_13866,N_13950);
nor U14064 (N_14064,N_13809,N_13812);
nand U14065 (N_14065,N_13948,N_13996);
or U14066 (N_14066,N_13944,N_13911);
or U14067 (N_14067,N_13821,N_13816);
and U14068 (N_14068,N_13845,N_13930);
nand U14069 (N_14069,N_13894,N_13976);
nand U14070 (N_14070,N_13973,N_13979);
nor U14071 (N_14071,N_13876,N_13984);
or U14072 (N_14072,N_13905,N_13899);
xnor U14073 (N_14073,N_13953,N_13827);
and U14074 (N_14074,N_13884,N_13877);
nor U14075 (N_14075,N_13966,N_13925);
or U14076 (N_14076,N_13826,N_13801);
or U14077 (N_14077,N_13898,N_13954);
nor U14078 (N_14078,N_13834,N_13970);
or U14079 (N_14079,N_13924,N_13881);
nor U14080 (N_14080,N_13872,N_13940);
and U14081 (N_14081,N_13906,N_13932);
nand U14082 (N_14082,N_13861,N_13891);
or U14083 (N_14083,N_13889,N_13804);
and U14084 (N_14084,N_13946,N_13847);
nand U14085 (N_14085,N_13958,N_13910);
nor U14086 (N_14086,N_13883,N_13805);
nor U14087 (N_14087,N_13842,N_13859);
nand U14088 (N_14088,N_13820,N_13853);
nand U14089 (N_14089,N_13864,N_13998);
nand U14090 (N_14090,N_13822,N_13918);
or U14091 (N_14091,N_13887,N_13800);
and U14092 (N_14092,N_13882,N_13901);
nor U14093 (N_14093,N_13986,N_13952);
nand U14094 (N_14094,N_13836,N_13983);
or U14095 (N_14095,N_13831,N_13895);
and U14096 (N_14096,N_13825,N_13907);
nor U14097 (N_14097,N_13854,N_13955);
nor U14098 (N_14098,N_13938,N_13868);
nand U14099 (N_14099,N_13850,N_13995);
or U14100 (N_14100,N_13809,N_13818);
nand U14101 (N_14101,N_13893,N_13875);
nor U14102 (N_14102,N_13998,N_13858);
nor U14103 (N_14103,N_13963,N_13814);
or U14104 (N_14104,N_13936,N_13896);
nor U14105 (N_14105,N_13894,N_13895);
nand U14106 (N_14106,N_13838,N_13975);
nand U14107 (N_14107,N_13849,N_13888);
and U14108 (N_14108,N_13939,N_13931);
or U14109 (N_14109,N_13880,N_13966);
or U14110 (N_14110,N_13905,N_13953);
nand U14111 (N_14111,N_13994,N_13909);
and U14112 (N_14112,N_13821,N_13950);
nand U14113 (N_14113,N_13902,N_13866);
and U14114 (N_14114,N_13869,N_13933);
nand U14115 (N_14115,N_13896,N_13942);
xnor U14116 (N_14116,N_13824,N_13928);
nor U14117 (N_14117,N_13827,N_13961);
nand U14118 (N_14118,N_13951,N_13946);
xor U14119 (N_14119,N_13924,N_13866);
nor U14120 (N_14120,N_13980,N_13948);
or U14121 (N_14121,N_13840,N_13963);
nor U14122 (N_14122,N_13883,N_13811);
or U14123 (N_14123,N_13818,N_13928);
nand U14124 (N_14124,N_13970,N_13946);
and U14125 (N_14125,N_13851,N_13866);
or U14126 (N_14126,N_13847,N_13950);
nor U14127 (N_14127,N_13991,N_13911);
nand U14128 (N_14128,N_13987,N_13914);
nor U14129 (N_14129,N_13987,N_13964);
and U14130 (N_14130,N_13854,N_13940);
or U14131 (N_14131,N_13973,N_13838);
nor U14132 (N_14132,N_13930,N_13904);
and U14133 (N_14133,N_13834,N_13894);
nand U14134 (N_14134,N_13809,N_13853);
and U14135 (N_14135,N_13907,N_13814);
nor U14136 (N_14136,N_13992,N_13966);
and U14137 (N_14137,N_13818,N_13988);
nor U14138 (N_14138,N_13831,N_13823);
and U14139 (N_14139,N_13857,N_13972);
or U14140 (N_14140,N_13917,N_13819);
and U14141 (N_14141,N_13931,N_13865);
nand U14142 (N_14142,N_13852,N_13801);
nand U14143 (N_14143,N_13815,N_13911);
nor U14144 (N_14144,N_13938,N_13900);
nand U14145 (N_14145,N_13897,N_13990);
or U14146 (N_14146,N_13938,N_13864);
nor U14147 (N_14147,N_13842,N_13997);
nor U14148 (N_14148,N_13935,N_13865);
nor U14149 (N_14149,N_13970,N_13982);
or U14150 (N_14150,N_13907,N_13830);
nor U14151 (N_14151,N_13842,N_13998);
nand U14152 (N_14152,N_13845,N_13927);
or U14153 (N_14153,N_13814,N_13871);
or U14154 (N_14154,N_13991,N_13893);
nor U14155 (N_14155,N_13939,N_13890);
nor U14156 (N_14156,N_13982,N_13988);
and U14157 (N_14157,N_13957,N_13969);
or U14158 (N_14158,N_13817,N_13958);
or U14159 (N_14159,N_13891,N_13812);
or U14160 (N_14160,N_13930,N_13913);
or U14161 (N_14161,N_13852,N_13924);
nor U14162 (N_14162,N_13909,N_13818);
nand U14163 (N_14163,N_13966,N_13977);
nand U14164 (N_14164,N_13984,N_13807);
or U14165 (N_14165,N_13948,N_13848);
nand U14166 (N_14166,N_13998,N_13958);
nand U14167 (N_14167,N_13934,N_13865);
or U14168 (N_14168,N_13831,N_13981);
nor U14169 (N_14169,N_13954,N_13871);
or U14170 (N_14170,N_13820,N_13849);
xor U14171 (N_14171,N_13845,N_13818);
or U14172 (N_14172,N_13815,N_13998);
nand U14173 (N_14173,N_13940,N_13915);
nor U14174 (N_14174,N_13874,N_13839);
nand U14175 (N_14175,N_13973,N_13937);
and U14176 (N_14176,N_13884,N_13940);
nor U14177 (N_14177,N_13896,N_13855);
or U14178 (N_14178,N_13840,N_13914);
nand U14179 (N_14179,N_13993,N_13803);
nor U14180 (N_14180,N_13974,N_13873);
xor U14181 (N_14181,N_13931,N_13823);
or U14182 (N_14182,N_13977,N_13833);
xnor U14183 (N_14183,N_13862,N_13945);
or U14184 (N_14184,N_13900,N_13833);
and U14185 (N_14185,N_13894,N_13929);
or U14186 (N_14186,N_13967,N_13858);
nand U14187 (N_14187,N_13896,N_13809);
nand U14188 (N_14188,N_13847,N_13919);
or U14189 (N_14189,N_13959,N_13810);
nor U14190 (N_14190,N_13910,N_13834);
or U14191 (N_14191,N_13813,N_13922);
nand U14192 (N_14192,N_13844,N_13826);
nand U14193 (N_14193,N_13877,N_13969);
or U14194 (N_14194,N_13861,N_13901);
and U14195 (N_14195,N_13801,N_13902);
or U14196 (N_14196,N_13843,N_13963);
and U14197 (N_14197,N_13813,N_13887);
and U14198 (N_14198,N_13826,N_13916);
or U14199 (N_14199,N_13853,N_13939);
or U14200 (N_14200,N_14014,N_14178);
nand U14201 (N_14201,N_14146,N_14118);
and U14202 (N_14202,N_14016,N_14011);
nor U14203 (N_14203,N_14051,N_14122);
nor U14204 (N_14204,N_14023,N_14001);
and U14205 (N_14205,N_14002,N_14083);
or U14206 (N_14206,N_14187,N_14056);
nand U14207 (N_14207,N_14152,N_14113);
or U14208 (N_14208,N_14165,N_14010);
nand U14209 (N_14209,N_14167,N_14192);
or U14210 (N_14210,N_14163,N_14173);
nand U14211 (N_14211,N_14093,N_14097);
nand U14212 (N_14212,N_14112,N_14139);
xor U14213 (N_14213,N_14191,N_14190);
xor U14214 (N_14214,N_14041,N_14168);
xnor U14215 (N_14215,N_14107,N_14099);
nor U14216 (N_14216,N_14132,N_14183);
or U14217 (N_14217,N_14071,N_14094);
or U14218 (N_14218,N_14111,N_14038);
nor U14219 (N_14219,N_14176,N_14170);
xnor U14220 (N_14220,N_14162,N_14159);
or U14221 (N_14221,N_14196,N_14156);
nor U14222 (N_14222,N_14120,N_14096);
nand U14223 (N_14223,N_14089,N_14064);
nor U14224 (N_14224,N_14047,N_14019);
or U14225 (N_14225,N_14022,N_14189);
and U14226 (N_14226,N_14007,N_14151);
or U14227 (N_14227,N_14172,N_14069);
nand U14228 (N_14228,N_14033,N_14029);
nand U14229 (N_14229,N_14150,N_14091);
nand U14230 (N_14230,N_14013,N_14055);
xor U14231 (N_14231,N_14021,N_14050);
and U14232 (N_14232,N_14067,N_14034);
or U14233 (N_14233,N_14006,N_14017);
xnor U14234 (N_14234,N_14004,N_14144);
nand U14235 (N_14235,N_14043,N_14155);
and U14236 (N_14236,N_14018,N_14053);
and U14237 (N_14237,N_14110,N_14186);
nor U14238 (N_14238,N_14081,N_14130);
xor U14239 (N_14239,N_14161,N_14092);
or U14240 (N_14240,N_14135,N_14049);
nor U14241 (N_14241,N_14009,N_14140);
nor U14242 (N_14242,N_14199,N_14102);
and U14243 (N_14243,N_14076,N_14119);
and U14244 (N_14244,N_14020,N_14160);
nor U14245 (N_14245,N_14166,N_14042);
nand U14246 (N_14246,N_14116,N_14154);
or U14247 (N_14247,N_14141,N_14101);
and U14248 (N_14248,N_14149,N_14126);
nand U14249 (N_14249,N_14039,N_14164);
nor U14250 (N_14250,N_14078,N_14195);
nand U14251 (N_14251,N_14036,N_14185);
nand U14252 (N_14252,N_14142,N_14012);
nor U14253 (N_14253,N_14157,N_14075);
or U14254 (N_14254,N_14068,N_14114);
and U14255 (N_14255,N_14052,N_14123);
nor U14256 (N_14256,N_14087,N_14105);
and U14257 (N_14257,N_14058,N_14045);
nor U14258 (N_14258,N_14025,N_14082);
xor U14259 (N_14259,N_14090,N_14184);
or U14260 (N_14260,N_14040,N_14100);
nand U14261 (N_14261,N_14054,N_14134);
nor U14262 (N_14262,N_14037,N_14061);
or U14263 (N_14263,N_14117,N_14198);
nand U14264 (N_14264,N_14084,N_14026);
and U14265 (N_14265,N_14133,N_14153);
nand U14266 (N_14266,N_14148,N_14145);
and U14267 (N_14267,N_14070,N_14085);
nor U14268 (N_14268,N_14115,N_14024);
nand U14269 (N_14269,N_14175,N_14169);
xor U14270 (N_14270,N_14137,N_14138);
and U14271 (N_14271,N_14103,N_14181);
or U14272 (N_14272,N_14106,N_14127);
xnor U14273 (N_14273,N_14060,N_14108);
and U14274 (N_14274,N_14000,N_14073);
or U14275 (N_14275,N_14077,N_14059);
nor U14276 (N_14276,N_14158,N_14080);
and U14277 (N_14277,N_14028,N_14086);
and U14278 (N_14278,N_14174,N_14182);
nor U14279 (N_14279,N_14032,N_14057);
and U14280 (N_14280,N_14088,N_14095);
nand U14281 (N_14281,N_14194,N_14027);
and U14282 (N_14282,N_14063,N_14136);
xor U14283 (N_14283,N_14177,N_14193);
nor U14284 (N_14284,N_14143,N_14074);
or U14285 (N_14285,N_14046,N_14131);
nor U14286 (N_14286,N_14031,N_14005);
nor U14287 (N_14287,N_14129,N_14121);
or U14288 (N_14288,N_14098,N_14008);
xor U14289 (N_14289,N_14125,N_14124);
or U14290 (N_14290,N_14104,N_14079);
xor U14291 (N_14291,N_14048,N_14179);
or U14292 (N_14292,N_14015,N_14147);
nor U14293 (N_14293,N_14044,N_14003);
nand U14294 (N_14294,N_14072,N_14171);
nand U14295 (N_14295,N_14197,N_14188);
and U14296 (N_14296,N_14180,N_14065);
nor U14297 (N_14297,N_14128,N_14066);
nor U14298 (N_14298,N_14030,N_14109);
and U14299 (N_14299,N_14062,N_14035);
and U14300 (N_14300,N_14081,N_14004);
xor U14301 (N_14301,N_14148,N_14012);
and U14302 (N_14302,N_14103,N_14119);
and U14303 (N_14303,N_14014,N_14098);
or U14304 (N_14304,N_14186,N_14044);
and U14305 (N_14305,N_14125,N_14040);
xnor U14306 (N_14306,N_14027,N_14120);
nor U14307 (N_14307,N_14155,N_14099);
or U14308 (N_14308,N_14191,N_14014);
or U14309 (N_14309,N_14008,N_14120);
or U14310 (N_14310,N_14010,N_14071);
nand U14311 (N_14311,N_14008,N_14087);
nor U14312 (N_14312,N_14117,N_14069);
or U14313 (N_14313,N_14086,N_14119);
nor U14314 (N_14314,N_14049,N_14096);
and U14315 (N_14315,N_14131,N_14169);
or U14316 (N_14316,N_14013,N_14052);
nor U14317 (N_14317,N_14084,N_14117);
nand U14318 (N_14318,N_14092,N_14078);
nand U14319 (N_14319,N_14047,N_14115);
nor U14320 (N_14320,N_14193,N_14047);
or U14321 (N_14321,N_14048,N_14037);
nand U14322 (N_14322,N_14054,N_14188);
or U14323 (N_14323,N_14023,N_14171);
nor U14324 (N_14324,N_14042,N_14181);
nand U14325 (N_14325,N_14130,N_14124);
nor U14326 (N_14326,N_14198,N_14174);
or U14327 (N_14327,N_14188,N_14156);
nor U14328 (N_14328,N_14091,N_14049);
or U14329 (N_14329,N_14120,N_14019);
xnor U14330 (N_14330,N_14123,N_14197);
nand U14331 (N_14331,N_14069,N_14066);
or U14332 (N_14332,N_14095,N_14069);
nand U14333 (N_14333,N_14097,N_14150);
nand U14334 (N_14334,N_14148,N_14089);
nor U14335 (N_14335,N_14027,N_14007);
and U14336 (N_14336,N_14088,N_14173);
and U14337 (N_14337,N_14064,N_14189);
nand U14338 (N_14338,N_14176,N_14190);
nor U14339 (N_14339,N_14044,N_14033);
and U14340 (N_14340,N_14124,N_14053);
nor U14341 (N_14341,N_14150,N_14180);
or U14342 (N_14342,N_14110,N_14046);
and U14343 (N_14343,N_14056,N_14162);
xor U14344 (N_14344,N_14122,N_14113);
nand U14345 (N_14345,N_14045,N_14197);
nor U14346 (N_14346,N_14084,N_14166);
and U14347 (N_14347,N_14095,N_14047);
nor U14348 (N_14348,N_14050,N_14020);
or U14349 (N_14349,N_14098,N_14110);
nor U14350 (N_14350,N_14009,N_14199);
xnor U14351 (N_14351,N_14174,N_14073);
or U14352 (N_14352,N_14039,N_14110);
nor U14353 (N_14353,N_14126,N_14181);
and U14354 (N_14354,N_14020,N_14057);
nor U14355 (N_14355,N_14092,N_14116);
or U14356 (N_14356,N_14109,N_14090);
or U14357 (N_14357,N_14092,N_14170);
or U14358 (N_14358,N_14118,N_14096);
or U14359 (N_14359,N_14169,N_14089);
xor U14360 (N_14360,N_14180,N_14169);
nand U14361 (N_14361,N_14192,N_14035);
nor U14362 (N_14362,N_14144,N_14099);
nand U14363 (N_14363,N_14154,N_14009);
nand U14364 (N_14364,N_14017,N_14023);
nand U14365 (N_14365,N_14028,N_14040);
nand U14366 (N_14366,N_14129,N_14061);
nand U14367 (N_14367,N_14196,N_14097);
nor U14368 (N_14368,N_14129,N_14081);
nand U14369 (N_14369,N_14154,N_14141);
and U14370 (N_14370,N_14033,N_14147);
nand U14371 (N_14371,N_14087,N_14084);
and U14372 (N_14372,N_14025,N_14188);
nor U14373 (N_14373,N_14032,N_14113);
xnor U14374 (N_14374,N_14092,N_14182);
nand U14375 (N_14375,N_14083,N_14189);
nand U14376 (N_14376,N_14160,N_14174);
xnor U14377 (N_14377,N_14113,N_14153);
nor U14378 (N_14378,N_14192,N_14152);
and U14379 (N_14379,N_14058,N_14032);
nor U14380 (N_14380,N_14134,N_14053);
nand U14381 (N_14381,N_14038,N_14098);
xnor U14382 (N_14382,N_14177,N_14099);
or U14383 (N_14383,N_14168,N_14021);
nand U14384 (N_14384,N_14153,N_14124);
xor U14385 (N_14385,N_14009,N_14030);
nor U14386 (N_14386,N_14126,N_14075);
xnor U14387 (N_14387,N_14149,N_14084);
or U14388 (N_14388,N_14101,N_14090);
or U14389 (N_14389,N_14044,N_14016);
and U14390 (N_14390,N_14051,N_14111);
or U14391 (N_14391,N_14144,N_14164);
or U14392 (N_14392,N_14142,N_14071);
nand U14393 (N_14393,N_14026,N_14195);
xor U14394 (N_14394,N_14182,N_14150);
nand U14395 (N_14395,N_14077,N_14038);
and U14396 (N_14396,N_14129,N_14055);
nand U14397 (N_14397,N_14000,N_14089);
and U14398 (N_14398,N_14148,N_14072);
or U14399 (N_14399,N_14029,N_14162);
nand U14400 (N_14400,N_14263,N_14238);
or U14401 (N_14401,N_14388,N_14274);
and U14402 (N_14402,N_14213,N_14314);
nand U14403 (N_14403,N_14209,N_14331);
or U14404 (N_14404,N_14351,N_14342);
and U14405 (N_14405,N_14299,N_14223);
and U14406 (N_14406,N_14229,N_14217);
nand U14407 (N_14407,N_14369,N_14211);
and U14408 (N_14408,N_14260,N_14309);
xor U14409 (N_14409,N_14358,N_14287);
nand U14410 (N_14410,N_14333,N_14216);
nand U14411 (N_14411,N_14231,N_14389);
nand U14412 (N_14412,N_14203,N_14234);
and U14413 (N_14413,N_14256,N_14355);
nand U14414 (N_14414,N_14367,N_14200);
nand U14415 (N_14415,N_14214,N_14207);
xnor U14416 (N_14416,N_14360,N_14265);
nand U14417 (N_14417,N_14377,N_14357);
or U14418 (N_14418,N_14324,N_14396);
and U14419 (N_14419,N_14390,N_14264);
nand U14420 (N_14420,N_14364,N_14359);
and U14421 (N_14421,N_14399,N_14218);
nand U14422 (N_14422,N_14278,N_14329);
nor U14423 (N_14423,N_14334,N_14255);
xor U14424 (N_14424,N_14322,N_14286);
or U14425 (N_14425,N_14325,N_14373);
xor U14426 (N_14426,N_14391,N_14280);
or U14427 (N_14427,N_14226,N_14227);
or U14428 (N_14428,N_14305,N_14266);
nand U14429 (N_14429,N_14340,N_14210);
nand U14430 (N_14430,N_14247,N_14252);
nand U14431 (N_14431,N_14318,N_14354);
nand U14432 (N_14432,N_14307,N_14328);
xnor U14433 (N_14433,N_14288,N_14366);
xor U14434 (N_14434,N_14381,N_14346);
or U14435 (N_14435,N_14387,N_14356);
nor U14436 (N_14436,N_14230,N_14393);
nor U14437 (N_14437,N_14250,N_14277);
or U14438 (N_14438,N_14253,N_14370);
nor U14439 (N_14439,N_14303,N_14332);
nand U14440 (N_14440,N_14383,N_14348);
and U14441 (N_14441,N_14310,N_14323);
nor U14442 (N_14442,N_14352,N_14371);
or U14443 (N_14443,N_14361,N_14241);
or U14444 (N_14444,N_14285,N_14363);
and U14445 (N_14445,N_14254,N_14271);
nor U14446 (N_14446,N_14344,N_14315);
nand U14447 (N_14447,N_14335,N_14395);
nand U14448 (N_14448,N_14304,N_14242);
and U14449 (N_14449,N_14205,N_14374);
nor U14450 (N_14450,N_14341,N_14269);
or U14451 (N_14451,N_14385,N_14275);
nand U14452 (N_14452,N_14248,N_14257);
nor U14453 (N_14453,N_14239,N_14273);
nor U14454 (N_14454,N_14221,N_14379);
or U14455 (N_14455,N_14397,N_14368);
nor U14456 (N_14456,N_14394,N_14330);
and U14457 (N_14457,N_14282,N_14312);
or U14458 (N_14458,N_14353,N_14372);
nand U14459 (N_14459,N_14289,N_14249);
nor U14460 (N_14460,N_14327,N_14306);
and U14461 (N_14461,N_14233,N_14380);
or U14462 (N_14462,N_14228,N_14224);
or U14463 (N_14463,N_14345,N_14212);
or U14464 (N_14464,N_14343,N_14300);
xor U14465 (N_14465,N_14201,N_14298);
or U14466 (N_14466,N_14290,N_14259);
xnor U14467 (N_14467,N_14319,N_14326);
nor U14468 (N_14468,N_14398,N_14279);
nand U14469 (N_14469,N_14302,N_14336);
nand U14470 (N_14470,N_14313,N_14320);
nor U14471 (N_14471,N_14208,N_14362);
and U14472 (N_14472,N_14276,N_14347);
nor U14473 (N_14473,N_14204,N_14283);
nand U14474 (N_14474,N_14294,N_14281);
nand U14475 (N_14475,N_14232,N_14258);
and U14476 (N_14476,N_14350,N_14292);
nand U14477 (N_14477,N_14225,N_14386);
or U14478 (N_14478,N_14261,N_14235);
and U14479 (N_14479,N_14321,N_14267);
nand U14480 (N_14480,N_14237,N_14236);
or U14481 (N_14481,N_14206,N_14376);
nor U14482 (N_14482,N_14297,N_14384);
or U14483 (N_14483,N_14316,N_14246);
nor U14484 (N_14484,N_14244,N_14349);
or U14485 (N_14485,N_14311,N_14284);
or U14486 (N_14486,N_14338,N_14337);
nor U14487 (N_14487,N_14296,N_14243);
and U14488 (N_14488,N_14293,N_14262);
or U14489 (N_14489,N_14382,N_14375);
and U14490 (N_14490,N_14308,N_14222);
and U14491 (N_14491,N_14220,N_14392);
and U14492 (N_14492,N_14215,N_14378);
and U14493 (N_14493,N_14219,N_14272);
nor U14494 (N_14494,N_14339,N_14301);
or U14495 (N_14495,N_14202,N_14251);
and U14496 (N_14496,N_14365,N_14268);
and U14497 (N_14497,N_14245,N_14240);
and U14498 (N_14498,N_14295,N_14270);
and U14499 (N_14499,N_14317,N_14291);
nor U14500 (N_14500,N_14217,N_14346);
and U14501 (N_14501,N_14314,N_14258);
nor U14502 (N_14502,N_14229,N_14249);
or U14503 (N_14503,N_14226,N_14223);
or U14504 (N_14504,N_14261,N_14391);
nor U14505 (N_14505,N_14232,N_14277);
nor U14506 (N_14506,N_14206,N_14388);
xnor U14507 (N_14507,N_14264,N_14291);
nor U14508 (N_14508,N_14291,N_14379);
and U14509 (N_14509,N_14360,N_14340);
and U14510 (N_14510,N_14278,N_14300);
nand U14511 (N_14511,N_14357,N_14265);
xnor U14512 (N_14512,N_14323,N_14206);
and U14513 (N_14513,N_14239,N_14354);
and U14514 (N_14514,N_14357,N_14299);
or U14515 (N_14515,N_14359,N_14360);
and U14516 (N_14516,N_14370,N_14212);
and U14517 (N_14517,N_14225,N_14260);
or U14518 (N_14518,N_14246,N_14297);
and U14519 (N_14519,N_14375,N_14224);
nand U14520 (N_14520,N_14291,N_14386);
and U14521 (N_14521,N_14381,N_14225);
and U14522 (N_14522,N_14289,N_14322);
and U14523 (N_14523,N_14323,N_14383);
and U14524 (N_14524,N_14275,N_14317);
nand U14525 (N_14525,N_14379,N_14243);
and U14526 (N_14526,N_14251,N_14236);
nor U14527 (N_14527,N_14237,N_14355);
nand U14528 (N_14528,N_14236,N_14370);
nand U14529 (N_14529,N_14211,N_14296);
and U14530 (N_14530,N_14261,N_14354);
nor U14531 (N_14531,N_14386,N_14346);
or U14532 (N_14532,N_14375,N_14264);
and U14533 (N_14533,N_14240,N_14302);
nor U14534 (N_14534,N_14289,N_14330);
or U14535 (N_14535,N_14262,N_14349);
nor U14536 (N_14536,N_14387,N_14283);
and U14537 (N_14537,N_14219,N_14359);
and U14538 (N_14538,N_14214,N_14315);
or U14539 (N_14539,N_14309,N_14265);
xnor U14540 (N_14540,N_14287,N_14399);
or U14541 (N_14541,N_14317,N_14349);
or U14542 (N_14542,N_14263,N_14393);
or U14543 (N_14543,N_14394,N_14310);
or U14544 (N_14544,N_14262,N_14216);
or U14545 (N_14545,N_14253,N_14278);
and U14546 (N_14546,N_14240,N_14238);
nand U14547 (N_14547,N_14311,N_14200);
and U14548 (N_14548,N_14290,N_14287);
or U14549 (N_14549,N_14250,N_14383);
nand U14550 (N_14550,N_14322,N_14378);
or U14551 (N_14551,N_14324,N_14387);
and U14552 (N_14552,N_14354,N_14245);
nand U14553 (N_14553,N_14247,N_14368);
or U14554 (N_14554,N_14249,N_14318);
nand U14555 (N_14555,N_14274,N_14354);
and U14556 (N_14556,N_14287,N_14258);
nor U14557 (N_14557,N_14250,N_14223);
and U14558 (N_14558,N_14284,N_14344);
nor U14559 (N_14559,N_14291,N_14221);
and U14560 (N_14560,N_14353,N_14325);
and U14561 (N_14561,N_14310,N_14333);
nor U14562 (N_14562,N_14351,N_14369);
nor U14563 (N_14563,N_14226,N_14361);
nor U14564 (N_14564,N_14379,N_14380);
xor U14565 (N_14565,N_14364,N_14229);
nand U14566 (N_14566,N_14309,N_14324);
xor U14567 (N_14567,N_14325,N_14274);
and U14568 (N_14568,N_14325,N_14331);
nand U14569 (N_14569,N_14392,N_14270);
or U14570 (N_14570,N_14332,N_14217);
or U14571 (N_14571,N_14220,N_14344);
nand U14572 (N_14572,N_14320,N_14229);
nand U14573 (N_14573,N_14207,N_14263);
nor U14574 (N_14574,N_14254,N_14220);
nor U14575 (N_14575,N_14358,N_14391);
nand U14576 (N_14576,N_14284,N_14273);
and U14577 (N_14577,N_14291,N_14384);
nor U14578 (N_14578,N_14352,N_14384);
nor U14579 (N_14579,N_14360,N_14352);
and U14580 (N_14580,N_14374,N_14367);
and U14581 (N_14581,N_14331,N_14207);
xor U14582 (N_14582,N_14397,N_14223);
and U14583 (N_14583,N_14247,N_14391);
xor U14584 (N_14584,N_14306,N_14338);
xor U14585 (N_14585,N_14202,N_14275);
nor U14586 (N_14586,N_14339,N_14279);
or U14587 (N_14587,N_14231,N_14296);
nor U14588 (N_14588,N_14384,N_14372);
and U14589 (N_14589,N_14378,N_14210);
and U14590 (N_14590,N_14290,N_14248);
and U14591 (N_14591,N_14378,N_14303);
or U14592 (N_14592,N_14221,N_14308);
nand U14593 (N_14593,N_14267,N_14337);
nand U14594 (N_14594,N_14310,N_14216);
nor U14595 (N_14595,N_14360,N_14308);
nor U14596 (N_14596,N_14257,N_14335);
or U14597 (N_14597,N_14319,N_14357);
nor U14598 (N_14598,N_14238,N_14264);
nand U14599 (N_14599,N_14283,N_14322);
nand U14600 (N_14600,N_14561,N_14510);
or U14601 (N_14601,N_14579,N_14419);
xor U14602 (N_14602,N_14493,N_14438);
or U14603 (N_14603,N_14573,N_14422);
nor U14604 (N_14604,N_14440,N_14566);
xor U14605 (N_14605,N_14410,N_14456);
or U14606 (N_14606,N_14484,N_14401);
nand U14607 (N_14607,N_14454,N_14504);
or U14608 (N_14608,N_14408,N_14525);
and U14609 (N_14609,N_14433,N_14558);
nand U14610 (N_14610,N_14567,N_14500);
or U14611 (N_14611,N_14596,N_14444);
or U14612 (N_14612,N_14439,N_14520);
or U14613 (N_14613,N_14513,N_14551);
and U14614 (N_14614,N_14588,N_14404);
or U14615 (N_14615,N_14432,N_14589);
nand U14616 (N_14616,N_14443,N_14515);
or U14617 (N_14617,N_14505,N_14564);
nand U14618 (N_14618,N_14570,N_14402);
xor U14619 (N_14619,N_14495,N_14425);
or U14620 (N_14620,N_14571,N_14494);
or U14621 (N_14621,N_14580,N_14575);
nand U14622 (N_14622,N_14529,N_14538);
nor U14623 (N_14623,N_14523,N_14437);
or U14624 (N_14624,N_14599,N_14507);
or U14625 (N_14625,N_14569,N_14465);
nand U14626 (N_14626,N_14423,N_14470);
and U14627 (N_14627,N_14591,N_14453);
xor U14628 (N_14628,N_14446,N_14597);
or U14629 (N_14629,N_14536,N_14594);
xnor U14630 (N_14630,N_14543,N_14428);
or U14631 (N_14631,N_14553,N_14539);
nand U14632 (N_14632,N_14481,N_14458);
or U14633 (N_14633,N_14563,N_14487);
and U14634 (N_14634,N_14461,N_14473);
xnor U14635 (N_14635,N_14577,N_14518);
nand U14636 (N_14636,N_14595,N_14431);
and U14637 (N_14637,N_14581,N_14450);
nor U14638 (N_14638,N_14545,N_14424);
nand U14639 (N_14639,N_14441,N_14414);
nor U14640 (N_14640,N_14593,N_14436);
nand U14641 (N_14641,N_14405,N_14560);
nand U14642 (N_14642,N_14530,N_14565);
nor U14643 (N_14643,N_14485,N_14497);
xnor U14644 (N_14644,N_14476,N_14598);
or U14645 (N_14645,N_14512,N_14421);
or U14646 (N_14646,N_14528,N_14413);
and U14647 (N_14647,N_14435,N_14502);
nand U14648 (N_14648,N_14469,N_14556);
or U14649 (N_14649,N_14409,N_14585);
nand U14650 (N_14650,N_14420,N_14445);
nand U14651 (N_14651,N_14482,N_14480);
and U14652 (N_14652,N_14537,N_14514);
nand U14653 (N_14653,N_14568,N_14496);
nand U14654 (N_14654,N_14474,N_14407);
or U14655 (N_14655,N_14448,N_14426);
or U14656 (N_14656,N_14531,N_14455);
nand U14657 (N_14657,N_14509,N_14459);
nor U14658 (N_14658,N_14491,N_14462);
nor U14659 (N_14659,N_14449,N_14478);
xor U14660 (N_14660,N_14427,N_14521);
nor U14661 (N_14661,N_14488,N_14519);
nand U14662 (N_14662,N_14486,N_14429);
or U14663 (N_14663,N_14540,N_14503);
nor U14664 (N_14664,N_14406,N_14535);
xor U14665 (N_14665,N_14590,N_14501);
and U14666 (N_14666,N_14584,N_14550);
or U14667 (N_14667,N_14574,N_14434);
nand U14668 (N_14668,N_14583,N_14552);
nor U14669 (N_14669,N_14554,N_14452);
or U14670 (N_14670,N_14541,N_14549);
or U14671 (N_14671,N_14516,N_14508);
nor U14672 (N_14672,N_14411,N_14403);
nor U14673 (N_14673,N_14412,N_14471);
nand U14674 (N_14674,N_14475,N_14559);
nor U14675 (N_14675,N_14511,N_14479);
xnor U14676 (N_14676,N_14546,N_14447);
and U14677 (N_14677,N_14468,N_14534);
xnor U14678 (N_14678,N_14524,N_14506);
or U14679 (N_14679,N_14489,N_14400);
nor U14680 (N_14680,N_14582,N_14544);
or U14681 (N_14681,N_14578,N_14587);
nor U14682 (N_14682,N_14442,N_14522);
nand U14683 (N_14683,N_14460,N_14499);
xor U14684 (N_14684,N_14492,N_14472);
or U14685 (N_14685,N_14430,N_14542);
and U14686 (N_14686,N_14548,N_14416);
or U14687 (N_14687,N_14592,N_14463);
nor U14688 (N_14688,N_14466,N_14418);
nor U14689 (N_14689,N_14572,N_14517);
and U14690 (N_14690,N_14527,N_14457);
nand U14691 (N_14691,N_14490,N_14547);
nor U14692 (N_14692,N_14533,N_14464);
and U14693 (N_14693,N_14415,N_14555);
or U14694 (N_14694,N_14483,N_14586);
nor U14695 (N_14695,N_14526,N_14467);
nor U14696 (N_14696,N_14498,N_14557);
nor U14697 (N_14697,N_14417,N_14451);
nor U14698 (N_14698,N_14477,N_14576);
nand U14699 (N_14699,N_14532,N_14562);
or U14700 (N_14700,N_14585,N_14589);
and U14701 (N_14701,N_14467,N_14584);
and U14702 (N_14702,N_14543,N_14512);
nand U14703 (N_14703,N_14412,N_14544);
nand U14704 (N_14704,N_14474,N_14548);
xnor U14705 (N_14705,N_14527,N_14413);
and U14706 (N_14706,N_14534,N_14449);
or U14707 (N_14707,N_14468,N_14568);
and U14708 (N_14708,N_14411,N_14597);
nand U14709 (N_14709,N_14582,N_14508);
nand U14710 (N_14710,N_14517,N_14516);
xnor U14711 (N_14711,N_14575,N_14569);
or U14712 (N_14712,N_14402,N_14530);
or U14713 (N_14713,N_14404,N_14495);
and U14714 (N_14714,N_14541,N_14464);
nand U14715 (N_14715,N_14477,N_14570);
and U14716 (N_14716,N_14408,N_14427);
nor U14717 (N_14717,N_14457,N_14558);
or U14718 (N_14718,N_14482,N_14597);
or U14719 (N_14719,N_14501,N_14496);
xor U14720 (N_14720,N_14585,N_14591);
or U14721 (N_14721,N_14426,N_14500);
xnor U14722 (N_14722,N_14492,N_14480);
nor U14723 (N_14723,N_14445,N_14497);
nand U14724 (N_14724,N_14500,N_14436);
xnor U14725 (N_14725,N_14597,N_14451);
nor U14726 (N_14726,N_14429,N_14470);
nor U14727 (N_14727,N_14422,N_14501);
nor U14728 (N_14728,N_14439,N_14491);
nor U14729 (N_14729,N_14584,N_14523);
or U14730 (N_14730,N_14508,N_14478);
nor U14731 (N_14731,N_14545,N_14476);
or U14732 (N_14732,N_14501,N_14463);
or U14733 (N_14733,N_14596,N_14545);
or U14734 (N_14734,N_14547,N_14458);
and U14735 (N_14735,N_14442,N_14429);
and U14736 (N_14736,N_14570,N_14544);
and U14737 (N_14737,N_14527,N_14468);
xnor U14738 (N_14738,N_14518,N_14470);
nand U14739 (N_14739,N_14566,N_14428);
nor U14740 (N_14740,N_14400,N_14485);
nand U14741 (N_14741,N_14550,N_14408);
or U14742 (N_14742,N_14528,N_14401);
xnor U14743 (N_14743,N_14579,N_14547);
and U14744 (N_14744,N_14436,N_14513);
nand U14745 (N_14745,N_14544,N_14523);
nand U14746 (N_14746,N_14466,N_14520);
or U14747 (N_14747,N_14565,N_14590);
nor U14748 (N_14748,N_14474,N_14428);
nor U14749 (N_14749,N_14565,N_14533);
nand U14750 (N_14750,N_14478,N_14481);
and U14751 (N_14751,N_14412,N_14425);
or U14752 (N_14752,N_14480,N_14417);
nor U14753 (N_14753,N_14574,N_14473);
nor U14754 (N_14754,N_14466,N_14437);
xnor U14755 (N_14755,N_14513,N_14408);
nor U14756 (N_14756,N_14540,N_14544);
and U14757 (N_14757,N_14407,N_14534);
nand U14758 (N_14758,N_14418,N_14490);
nand U14759 (N_14759,N_14597,N_14518);
nand U14760 (N_14760,N_14505,N_14499);
and U14761 (N_14761,N_14463,N_14568);
nand U14762 (N_14762,N_14562,N_14538);
nor U14763 (N_14763,N_14493,N_14509);
and U14764 (N_14764,N_14578,N_14413);
or U14765 (N_14765,N_14500,N_14558);
or U14766 (N_14766,N_14510,N_14466);
nor U14767 (N_14767,N_14469,N_14512);
nor U14768 (N_14768,N_14417,N_14529);
nand U14769 (N_14769,N_14582,N_14463);
and U14770 (N_14770,N_14466,N_14557);
or U14771 (N_14771,N_14436,N_14507);
or U14772 (N_14772,N_14502,N_14494);
or U14773 (N_14773,N_14504,N_14502);
and U14774 (N_14774,N_14449,N_14518);
or U14775 (N_14775,N_14503,N_14484);
nand U14776 (N_14776,N_14514,N_14404);
and U14777 (N_14777,N_14447,N_14470);
and U14778 (N_14778,N_14488,N_14585);
or U14779 (N_14779,N_14400,N_14578);
and U14780 (N_14780,N_14495,N_14460);
or U14781 (N_14781,N_14481,N_14504);
or U14782 (N_14782,N_14496,N_14558);
or U14783 (N_14783,N_14501,N_14418);
nor U14784 (N_14784,N_14437,N_14413);
or U14785 (N_14785,N_14561,N_14477);
nor U14786 (N_14786,N_14469,N_14442);
and U14787 (N_14787,N_14576,N_14411);
and U14788 (N_14788,N_14438,N_14445);
nand U14789 (N_14789,N_14432,N_14423);
and U14790 (N_14790,N_14589,N_14571);
or U14791 (N_14791,N_14516,N_14460);
xor U14792 (N_14792,N_14485,N_14452);
and U14793 (N_14793,N_14408,N_14570);
and U14794 (N_14794,N_14543,N_14553);
xor U14795 (N_14795,N_14586,N_14548);
nand U14796 (N_14796,N_14480,N_14487);
or U14797 (N_14797,N_14544,N_14478);
nor U14798 (N_14798,N_14528,N_14542);
nor U14799 (N_14799,N_14552,N_14410);
or U14800 (N_14800,N_14691,N_14653);
xnor U14801 (N_14801,N_14700,N_14695);
nor U14802 (N_14802,N_14636,N_14613);
or U14803 (N_14803,N_14660,N_14739);
nor U14804 (N_14804,N_14777,N_14756);
nand U14805 (N_14805,N_14799,N_14774);
xor U14806 (N_14806,N_14627,N_14626);
and U14807 (N_14807,N_14712,N_14758);
nor U14808 (N_14808,N_14654,N_14642);
or U14809 (N_14809,N_14658,N_14771);
and U14810 (N_14810,N_14787,N_14731);
or U14811 (N_14811,N_14671,N_14718);
nand U14812 (N_14812,N_14728,N_14606);
nand U14813 (N_14813,N_14666,N_14741);
xor U14814 (N_14814,N_14701,N_14619);
and U14815 (N_14815,N_14721,N_14692);
nor U14816 (N_14816,N_14738,N_14724);
xnor U14817 (N_14817,N_14750,N_14765);
nand U14818 (N_14818,N_14649,N_14664);
nand U14819 (N_14819,N_14639,N_14600);
nand U14820 (N_14820,N_14678,N_14707);
or U14821 (N_14821,N_14632,N_14672);
and U14822 (N_14822,N_14734,N_14633);
nor U14823 (N_14823,N_14785,N_14635);
nor U14824 (N_14824,N_14770,N_14608);
nand U14825 (N_14825,N_14711,N_14648);
nor U14826 (N_14826,N_14674,N_14745);
nand U14827 (N_14827,N_14623,N_14614);
and U14828 (N_14828,N_14719,N_14652);
nand U14829 (N_14829,N_14759,N_14729);
or U14830 (N_14830,N_14610,N_14735);
or U14831 (N_14831,N_14783,N_14789);
and U14832 (N_14832,N_14616,N_14710);
xnor U14833 (N_14833,N_14618,N_14763);
and U14834 (N_14834,N_14643,N_14647);
nor U14835 (N_14835,N_14629,N_14628);
nor U14836 (N_14836,N_14732,N_14780);
and U14837 (N_14837,N_14687,N_14762);
and U14838 (N_14838,N_14798,N_14661);
nor U14839 (N_14839,N_14768,N_14645);
and U14840 (N_14840,N_14650,N_14673);
and U14841 (N_14841,N_14611,N_14630);
nand U14842 (N_14842,N_14743,N_14605);
or U14843 (N_14843,N_14602,N_14754);
or U14844 (N_14844,N_14740,N_14681);
or U14845 (N_14845,N_14742,N_14684);
xnor U14846 (N_14846,N_14634,N_14625);
xor U14847 (N_14847,N_14790,N_14655);
nor U14848 (N_14848,N_14683,N_14705);
nand U14849 (N_14849,N_14656,N_14663);
and U14850 (N_14850,N_14795,N_14607);
and U14851 (N_14851,N_14644,N_14796);
nor U14852 (N_14852,N_14669,N_14709);
nor U14853 (N_14853,N_14752,N_14677);
and U14854 (N_14854,N_14675,N_14764);
or U14855 (N_14855,N_14665,N_14631);
and U14856 (N_14856,N_14638,N_14690);
or U14857 (N_14857,N_14730,N_14708);
xnor U14858 (N_14858,N_14791,N_14640);
and U14859 (N_14859,N_14714,N_14615);
nand U14860 (N_14860,N_14679,N_14723);
nor U14861 (N_14861,N_14736,N_14609);
nor U14862 (N_14862,N_14689,N_14668);
nand U14863 (N_14863,N_14746,N_14755);
nor U14864 (N_14864,N_14688,N_14757);
or U14865 (N_14865,N_14775,N_14797);
nand U14866 (N_14866,N_14792,N_14766);
nand U14867 (N_14867,N_14779,N_14703);
nor U14868 (N_14868,N_14637,N_14760);
and U14869 (N_14869,N_14697,N_14667);
nor U14870 (N_14870,N_14737,N_14720);
or U14871 (N_14871,N_14733,N_14601);
and U14872 (N_14872,N_14651,N_14686);
or U14873 (N_14873,N_14704,N_14682);
or U14874 (N_14874,N_14622,N_14751);
nand U14875 (N_14875,N_14753,N_14717);
or U14876 (N_14876,N_14715,N_14769);
nand U14877 (N_14877,N_14776,N_14670);
xnor U14878 (N_14878,N_14722,N_14676);
or U14879 (N_14879,N_14726,N_14727);
xnor U14880 (N_14880,N_14646,N_14782);
and U14881 (N_14881,N_14778,N_14603);
and U14882 (N_14882,N_14749,N_14662);
xnor U14883 (N_14883,N_14699,N_14716);
nand U14884 (N_14884,N_14748,N_14784);
xor U14885 (N_14885,N_14773,N_14698);
or U14886 (N_14886,N_14781,N_14620);
and U14887 (N_14887,N_14696,N_14657);
and U14888 (N_14888,N_14744,N_14794);
or U14889 (N_14889,N_14761,N_14767);
or U14890 (N_14890,N_14706,N_14612);
nor U14891 (N_14891,N_14747,N_14786);
and U14892 (N_14892,N_14713,N_14793);
nand U14893 (N_14893,N_14680,N_14641);
or U14894 (N_14894,N_14702,N_14617);
nand U14895 (N_14895,N_14772,N_14694);
or U14896 (N_14896,N_14621,N_14685);
nand U14897 (N_14897,N_14659,N_14788);
nand U14898 (N_14898,N_14693,N_14725);
nor U14899 (N_14899,N_14624,N_14604);
xnor U14900 (N_14900,N_14657,N_14772);
nor U14901 (N_14901,N_14772,N_14692);
nand U14902 (N_14902,N_14708,N_14741);
nor U14903 (N_14903,N_14651,N_14744);
xor U14904 (N_14904,N_14763,N_14778);
nand U14905 (N_14905,N_14713,N_14703);
nand U14906 (N_14906,N_14607,N_14770);
nand U14907 (N_14907,N_14649,N_14737);
or U14908 (N_14908,N_14663,N_14702);
and U14909 (N_14909,N_14780,N_14605);
and U14910 (N_14910,N_14723,N_14656);
nor U14911 (N_14911,N_14682,N_14715);
nand U14912 (N_14912,N_14709,N_14673);
nand U14913 (N_14913,N_14749,N_14646);
and U14914 (N_14914,N_14609,N_14615);
or U14915 (N_14915,N_14687,N_14737);
nand U14916 (N_14916,N_14625,N_14783);
nand U14917 (N_14917,N_14776,N_14797);
nor U14918 (N_14918,N_14662,N_14623);
or U14919 (N_14919,N_14671,N_14687);
or U14920 (N_14920,N_14615,N_14795);
nand U14921 (N_14921,N_14794,N_14658);
and U14922 (N_14922,N_14758,N_14789);
nor U14923 (N_14923,N_14675,N_14749);
or U14924 (N_14924,N_14625,N_14744);
and U14925 (N_14925,N_14642,N_14664);
nand U14926 (N_14926,N_14746,N_14794);
nor U14927 (N_14927,N_14652,N_14646);
nor U14928 (N_14928,N_14753,N_14688);
nor U14929 (N_14929,N_14727,N_14616);
nor U14930 (N_14930,N_14735,N_14605);
nor U14931 (N_14931,N_14745,N_14655);
and U14932 (N_14932,N_14658,N_14705);
nor U14933 (N_14933,N_14786,N_14730);
nand U14934 (N_14934,N_14636,N_14638);
nand U14935 (N_14935,N_14725,N_14729);
nand U14936 (N_14936,N_14624,N_14756);
nor U14937 (N_14937,N_14744,N_14691);
or U14938 (N_14938,N_14605,N_14791);
nand U14939 (N_14939,N_14694,N_14622);
nand U14940 (N_14940,N_14787,N_14764);
nor U14941 (N_14941,N_14663,N_14729);
and U14942 (N_14942,N_14716,N_14652);
nor U14943 (N_14943,N_14650,N_14773);
nor U14944 (N_14944,N_14751,N_14697);
and U14945 (N_14945,N_14764,N_14659);
nor U14946 (N_14946,N_14603,N_14690);
nand U14947 (N_14947,N_14715,N_14675);
and U14948 (N_14948,N_14643,N_14655);
and U14949 (N_14949,N_14651,N_14662);
or U14950 (N_14950,N_14787,N_14720);
and U14951 (N_14951,N_14786,N_14688);
nand U14952 (N_14952,N_14762,N_14748);
nand U14953 (N_14953,N_14782,N_14628);
nand U14954 (N_14954,N_14719,N_14604);
nor U14955 (N_14955,N_14622,N_14604);
nand U14956 (N_14956,N_14696,N_14668);
nor U14957 (N_14957,N_14733,N_14761);
and U14958 (N_14958,N_14719,N_14684);
and U14959 (N_14959,N_14711,N_14636);
or U14960 (N_14960,N_14722,N_14723);
or U14961 (N_14961,N_14762,N_14658);
nor U14962 (N_14962,N_14686,N_14631);
nand U14963 (N_14963,N_14623,N_14762);
and U14964 (N_14964,N_14734,N_14625);
nor U14965 (N_14965,N_14653,N_14794);
xor U14966 (N_14966,N_14785,N_14790);
nor U14967 (N_14967,N_14774,N_14767);
or U14968 (N_14968,N_14619,N_14710);
nand U14969 (N_14969,N_14757,N_14676);
or U14970 (N_14970,N_14630,N_14703);
or U14971 (N_14971,N_14741,N_14686);
nor U14972 (N_14972,N_14629,N_14636);
nand U14973 (N_14973,N_14698,N_14735);
nor U14974 (N_14974,N_14657,N_14715);
nand U14975 (N_14975,N_14623,N_14733);
xor U14976 (N_14976,N_14632,N_14667);
and U14977 (N_14977,N_14771,N_14770);
nand U14978 (N_14978,N_14634,N_14759);
and U14979 (N_14979,N_14770,N_14795);
and U14980 (N_14980,N_14763,N_14672);
nand U14981 (N_14981,N_14658,N_14759);
nand U14982 (N_14982,N_14680,N_14710);
xor U14983 (N_14983,N_14613,N_14723);
or U14984 (N_14984,N_14675,N_14604);
nor U14985 (N_14985,N_14776,N_14772);
and U14986 (N_14986,N_14750,N_14662);
or U14987 (N_14987,N_14709,N_14702);
nand U14988 (N_14988,N_14694,N_14605);
nor U14989 (N_14989,N_14797,N_14743);
nand U14990 (N_14990,N_14792,N_14639);
nor U14991 (N_14991,N_14718,N_14605);
nand U14992 (N_14992,N_14710,N_14781);
nand U14993 (N_14993,N_14694,N_14660);
nor U14994 (N_14994,N_14694,N_14610);
xnor U14995 (N_14995,N_14603,N_14641);
nand U14996 (N_14996,N_14755,N_14792);
and U14997 (N_14997,N_14615,N_14793);
xor U14998 (N_14998,N_14746,N_14629);
nor U14999 (N_14999,N_14721,N_14771);
nand UO_0 (O_0,N_14978,N_14840);
and UO_1 (O_1,N_14819,N_14944);
xnor UO_2 (O_2,N_14852,N_14821);
nor UO_3 (O_3,N_14930,N_14846);
xor UO_4 (O_4,N_14904,N_14807);
nand UO_5 (O_5,N_14873,N_14876);
nor UO_6 (O_6,N_14857,N_14878);
and UO_7 (O_7,N_14896,N_14939);
nand UO_8 (O_8,N_14959,N_14877);
nor UO_9 (O_9,N_14940,N_14902);
nor UO_10 (O_10,N_14993,N_14991);
nand UO_11 (O_11,N_14874,N_14974);
xor UO_12 (O_12,N_14954,N_14864);
nor UO_13 (O_13,N_14910,N_14966);
nand UO_14 (O_14,N_14933,N_14950);
nor UO_15 (O_15,N_14975,N_14918);
and UO_16 (O_16,N_14947,N_14926);
nor UO_17 (O_17,N_14969,N_14943);
and UO_18 (O_18,N_14923,N_14838);
and UO_19 (O_19,N_14964,N_14855);
nor UO_20 (O_20,N_14880,N_14833);
or UO_21 (O_21,N_14800,N_14809);
nor UO_22 (O_22,N_14887,N_14998);
or UO_23 (O_23,N_14882,N_14837);
nor UO_24 (O_24,N_14937,N_14995);
or UO_25 (O_25,N_14850,N_14865);
or UO_26 (O_26,N_14936,N_14831);
and UO_27 (O_27,N_14823,N_14961);
and UO_28 (O_28,N_14989,N_14811);
or UO_29 (O_29,N_14982,N_14849);
and UO_30 (O_30,N_14919,N_14863);
and UO_31 (O_31,N_14962,N_14862);
nor UO_32 (O_32,N_14835,N_14928);
or UO_33 (O_33,N_14881,N_14883);
xor UO_34 (O_34,N_14909,N_14890);
nor UO_35 (O_35,N_14808,N_14911);
nand UO_36 (O_36,N_14951,N_14845);
nand UO_37 (O_37,N_14934,N_14903);
nor UO_38 (O_38,N_14888,N_14942);
nand UO_39 (O_39,N_14965,N_14972);
nor UO_40 (O_40,N_14822,N_14884);
xor UO_41 (O_41,N_14886,N_14971);
and UO_42 (O_42,N_14871,N_14957);
nor UO_43 (O_43,N_14851,N_14963);
nor UO_44 (O_44,N_14945,N_14858);
or UO_45 (O_45,N_14891,N_14805);
nand UO_46 (O_46,N_14872,N_14829);
nand UO_47 (O_47,N_14914,N_14815);
and UO_48 (O_48,N_14932,N_14906);
nor UO_49 (O_49,N_14924,N_14812);
nand UO_50 (O_50,N_14899,N_14856);
nor UO_51 (O_51,N_14960,N_14814);
nand UO_52 (O_52,N_14802,N_14996);
or UO_53 (O_53,N_14879,N_14860);
or UO_54 (O_54,N_14986,N_14810);
and UO_55 (O_55,N_14968,N_14967);
nor UO_56 (O_56,N_14981,N_14917);
and UO_57 (O_57,N_14867,N_14820);
or UO_58 (O_58,N_14915,N_14898);
and UO_59 (O_59,N_14894,N_14901);
and UO_60 (O_60,N_14987,N_14854);
or UO_61 (O_61,N_14817,N_14922);
and UO_62 (O_62,N_14893,N_14826);
or UO_63 (O_63,N_14853,N_14844);
nand UO_64 (O_64,N_14818,N_14828);
nor UO_65 (O_65,N_14806,N_14870);
and UO_66 (O_66,N_14920,N_14892);
nand UO_67 (O_67,N_14988,N_14834);
nand UO_68 (O_68,N_14983,N_14973);
or UO_69 (O_69,N_14946,N_14994);
or UO_70 (O_70,N_14953,N_14985);
and UO_71 (O_71,N_14916,N_14804);
xnor UO_72 (O_72,N_14992,N_14839);
or UO_73 (O_73,N_14825,N_14830);
nor UO_74 (O_74,N_14979,N_14908);
nand UO_75 (O_75,N_14866,N_14803);
xor UO_76 (O_76,N_14913,N_14827);
and UO_77 (O_77,N_14980,N_14999);
and UO_78 (O_78,N_14843,N_14927);
or UO_79 (O_79,N_14925,N_14958);
and UO_80 (O_80,N_14824,N_14970);
xor UO_81 (O_81,N_14931,N_14938);
xor UO_82 (O_82,N_14907,N_14897);
nand UO_83 (O_83,N_14935,N_14976);
nor UO_84 (O_84,N_14921,N_14868);
nor UO_85 (O_85,N_14941,N_14956);
or UO_86 (O_86,N_14861,N_14813);
nor UO_87 (O_87,N_14847,N_14859);
nand UO_88 (O_88,N_14885,N_14842);
nor UO_89 (O_89,N_14905,N_14900);
nand UO_90 (O_90,N_14948,N_14955);
and UO_91 (O_91,N_14889,N_14848);
or UO_92 (O_92,N_14895,N_14832);
or UO_93 (O_93,N_14990,N_14929);
nand UO_94 (O_94,N_14836,N_14997);
nor UO_95 (O_95,N_14912,N_14952);
and UO_96 (O_96,N_14949,N_14875);
or UO_97 (O_97,N_14801,N_14816);
or UO_98 (O_98,N_14841,N_14984);
nand UO_99 (O_99,N_14869,N_14977);
nand UO_100 (O_100,N_14880,N_14809);
nor UO_101 (O_101,N_14956,N_14889);
nand UO_102 (O_102,N_14927,N_14894);
nor UO_103 (O_103,N_14961,N_14970);
or UO_104 (O_104,N_14934,N_14913);
nor UO_105 (O_105,N_14995,N_14987);
and UO_106 (O_106,N_14968,N_14915);
or UO_107 (O_107,N_14891,N_14888);
xnor UO_108 (O_108,N_14897,N_14959);
or UO_109 (O_109,N_14938,N_14980);
or UO_110 (O_110,N_14957,N_14938);
xor UO_111 (O_111,N_14918,N_14907);
or UO_112 (O_112,N_14830,N_14872);
nor UO_113 (O_113,N_14992,N_14837);
xnor UO_114 (O_114,N_14859,N_14856);
nor UO_115 (O_115,N_14806,N_14888);
or UO_116 (O_116,N_14995,N_14931);
and UO_117 (O_117,N_14915,N_14923);
and UO_118 (O_118,N_14904,N_14845);
nand UO_119 (O_119,N_14801,N_14895);
or UO_120 (O_120,N_14910,N_14877);
or UO_121 (O_121,N_14847,N_14933);
and UO_122 (O_122,N_14877,N_14827);
or UO_123 (O_123,N_14838,N_14925);
nand UO_124 (O_124,N_14917,N_14864);
and UO_125 (O_125,N_14841,N_14952);
nand UO_126 (O_126,N_14850,N_14848);
xor UO_127 (O_127,N_14803,N_14825);
nand UO_128 (O_128,N_14804,N_14892);
nand UO_129 (O_129,N_14831,N_14917);
and UO_130 (O_130,N_14834,N_14998);
and UO_131 (O_131,N_14918,N_14833);
nor UO_132 (O_132,N_14921,N_14922);
or UO_133 (O_133,N_14973,N_14815);
and UO_134 (O_134,N_14912,N_14807);
or UO_135 (O_135,N_14991,N_14858);
and UO_136 (O_136,N_14946,N_14812);
xnor UO_137 (O_137,N_14919,N_14850);
xor UO_138 (O_138,N_14870,N_14987);
or UO_139 (O_139,N_14926,N_14909);
nor UO_140 (O_140,N_14818,N_14845);
nor UO_141 (O_141,N_14899,N_14839);
and UO_142 (O_142,N_14933,N_14877);
xnor UO_143 (O_143,N_14811,N_14837);
xnor UO_144 (O_144,N_14805,N_14811);
and UO_145 (O_145,N_14918,N_14861);
or UO_146 (O_146,N_14942,N_14914);
nor UO_147 (O_147,N_14933,N_14999);
or UO_148 (O_148,N_14920,N_14833);
nand UO_149 (O_149,N_14943,N_14870);
and UO_150 (O_150,N_14966,N_14890);
nand UO_151 (O_151,N_14969,N_14997);
nor UO_152 (O_152,N_14828,N_14824);
and UO_153 (O_153,N_14854,N_14840);
and UO_154 (O_154,N_14868,N_14940);
nor UO_155 (O_155,N_14958,N_14870);
nor UO_156 (O_156,N_14942,N_14921);
and UO_157 (O_157,N_14886,N_14904);
nor UO_158 (O_158,N_14828,N_14960);
nor UO_159 (O_159,N_14920,N_14829);
or UO_160 (O_160,N_14828,N_14939);
nand UO_161 (O_161,N_14919,N_14899);
or UO_162 (O_162,N_14816,N_14908);
and UO_163 (O_163,N_14920,N_14809);
nor UO_164 (O_164,N_14860,N_14817);
nor UO_165 (O_165,N_14876,N_14879);
and UO_166 (O_166,N_14927,N_14803);
or UO_167 (O_167,N_14854,N_14887);
nand UO_168 (O_168,N_14896,N_14815);
and UO_169 (O_169,N_14871,N_14948);
and UO_170 (O_170,N_14848,N_14819);
nand UO_171 (O_171,N_14851,N_14863);
nor UO_172 (O_172,N_14807,N_14810);
or UO_173 (O_173,N_14889,N_14976);
or UO_174 (O_174,N_14801,N_14868);
nor UO_175 (O_175,N_14878,N_14940);
or UO_176 (O_176,N_14876,N_14929);
nor UO_177 (O_177,N_14855,N_14810);
or UO_178 (O_178,N_14818,N_14928);
or UO_179 (O_179,N_14963,N_14956);
and UO_180 (O_180,N_14918,N_14887);
and UO_181 (O_181,N_14957,N_14828);
nor UO_182 (O_182,N_14838,N_14921);
nor UO_183 (O_183,N_14866,N_14842);
nand UO_184 (O_184,N_14920,N_14816);
nand UO_185 (O_185,N_14980,N_14939);
nand UO_186 (O_186,N_14929,N_14884);
xor UO_187 (O_187,N_14883,N_14863);
and UO_188 (O_188,N_14900,N_14894);
nand UO_189 (O_189,N_14893,N_14837);
nand UO_190 (O_190,N_14963,N_14910);
and UO_191 (O_191,N_14877,N_14980);
xnor UO_192 (O_192,N_14945,N_14881);
nor UO_193 (O_193,N_14854,N_14941);
and UO_194 (O_194,N_14962,N_14811);
xor UO_195 (O_195,N_14828,N_14833);
and UO_196 (O_196,N_14999,N_14902);
xor UO_197 (O_197,N_14978,N_14988);
nor UO_198 (O_198,N_14961,N_14814);
and UO_199 (O_199,N_14885,N_14880);
or UO_200 (O_200,N_14958,N_14993);
xor UO_201 (O_201,N_14906,N_14821);
or UO_202 (O_202,N_14847,N_14823);
nand UO_203 (O_203,N_14894,N_14973);
or UO_204 (O_204,N_14887,N_14838);
and UO_205 (O_205,N_14869,N_14850);
and UO_206 (O_206,N_14858,N_14817);
and UO_207 (O_207,N_14995,N_14884);
nand UO_208 (O_208,N_14954,N_14903);
nand UO_209 (O_209,N_14985,N_14832);
or UO_210 (O_210,N_14910,N_14946);
nor UO_211 (O_211,N_14981,N_14924);
and UO_212 (O_212,N_14856,N_14874);
nor UO_213 (O_213,N_14807,N_14981);
xor UO_214 (O_214,N_14809,N_14892);
or UO_215 (O_215,N_14972,N_14800);
nand UO_216 (O_216,N_14821,N_14897);
and UO_217 (O_217,N_14982,N_14987);
or UO_218 (O_218,N_14979,N_14946);
nor UO_219 (O_219,N_14848,N_14989);
or UO_220 (O_220,N_14951,N_14950);
nor UO_221 (O_221,N_14918,N_14999);
nor UO_222 (O_222,N_14917,N_14960);
nand UO_223 (O_223,N_14843,N_14929);
or UO_224 (O_224,N_14877,N_14884);
or UO_225 (O_225,N_14962,N_14991);
or UO_226 (O_226,N_14901,N_14882);
and UO_227 (O_227,N_14883,N_14888);
or UO_228 (O_228,N_14870,N_14873);
or UO_229 (O_229,N_14933,N_14864);
nor UO_230 (O_230,N_14824,N_14871);
and UO_231 (O_231,N_14935,N_14938);
nand UO_232 (O_232,N_14989,N_14934);
and UO_233 (O_233,N_14901,N_14989);
nor UO_234 (O_234,N_14933,N_14980);
or UO_235 (O_235,N_14865,N_14925);
and UO_236 (O_236,N_14835,N_14887);
nand UO_237 (O_237,N_14985,N_14973);
nand UO_238 (O_238,N_14935,N_14912);
and UO_239 (O_239,N_14801,N_14858);
and UO_240 (O_240,N_14981,N_14829);
or UO_241 (O_241,N_14988,N_14945);
nand UO_242 (O_242,N_14912,N_14993);
nand UO_243 (O_243,N_14920,N_14840);
and UO_244 (O_244,N_14810,N_14989);
or UO_245 (O_245,N_14809,N_14870);
xor UO_246 (O_246,N_14905,N_14975);
nand UO_247 (O_247,N_14947,N_14984);
nand UO_248 (O_248,N_14940,N_14829);
nand UO_249 (O_249,N_14968,N_14817);
nor UO_250 (O_250,N_14966,N_14924);
or UO_251 (O_251,N_14970,N_14984);
nand UO_252 (O_252,N_14951,N_14931);
or UO_253 (O_253,N_14923,N_14866);
nand UO_254 (O_254,N_14990,N_14827);
nor UO_255 (O_255,N_14951,N_14809);
xnor UO_256 (O_256,N_14844,N_14868);
xnor UO_257 (O_257,N_14926,N_14883);
and UO_258 (O_258,N_14986,N_14862);
nor UO_259 (O_259,N_14849,N_14834);
xnor UO_260 (O_260,N_14944,N_14902);
or UO_261 (O_261,N_14806,N_14974);
or UO_262 (O_262,N_14954,N_14995);
nor UO_263 (O_263,N_14857,N_14999);
nor UO_264 (O_264,N_14979,N_14977);
or UO_265 (O_265,N_14936,N_14893);
and UO_266 (O_266,N_14956,N_14873);
nand UO_267 (O_267,N_14999,N_14855);
and UO_268 (O_268,N_14845,N_14930);
and UO_269 (O_269,N_14829,N_14864);
nor UO_270 (O_270,N_14892,N_14973);
nand UO_271 (O_271,N_14969,N_14876);
nor UO_272 (O_272,N_14830,N_14928);
or UO_273 (O_273,N_14845,N_14996);
or UO_274 (O_274,N_14996,N_14976);
xnor UO_275 (O_275,N_14904,N_14958);
nand UO_276 (O_276,N_14976,N_14886);
or UO_277 (O_277,N_14954,N_14866);
and UO_278 (O_278,N_14874,N_14830);
nor UO_279 (O_279,N_14801,N_14813);
nand UO_280 (O_280,N_14973,N_14809);
or UO_281 (O_281,N_14971,N_14912);
nand UO_282 (O_282,N_14927,N_14889);
nand UO_283 (O_283,N_14889,N_14985);
nor UO_284 (O_284,N_14897,N_14923);
xnor UO_285 (O_285,N_14937,N_14898);
or UO_286 (O_286,N_14872,N_14902);
nor UO_287 (O_287,N_14997,N_14890);
and UO_288 (O_288,N_14903,N_14899);
nand UO_289 (O_289,N_14942,N_14852);
xnor UO_290 (O_290,N_14803,N_14923);
or UO_291 (O_291,N_14869,N_14928);
and UO_292 (O_292,N_14941,N_14825);
nand UO_293 (O_293,N_14951,N_14818);
or UO_294 (O_294,N_14959,N_14938);
and UO_295 (O_295,N_14902,N_14841);
and UO_296 (O_296,N_14891,N_14942);
nand UO_297 (O_297,N_14843,N_14809);
or UO_298 (O_298,N_14865,N_14837);
nand UO_299 (O_299,N_14919,N_14975);
and UO_300 (O_300,N_14998,N_14929);
and UO_301 (O_301,N_14858,N_14907);
or UO_302 (O_302,N_14854,N_14845);
nor UO_303 (O_303,N_14999,N_14976);
and UO_304 (O_304,N_14964,N_14925);
nand UO_305 (O_305,N_14965,N_14999);
xor UO_306 (O_306,N_14805,N_14858);
xor UO_307 (O_307,N_14897,N_14960);
and UO_308 (O_308,N_14884,N_14925);
and UO_309 (O_309,N_14801,N_14817);
nor UO_310 (O_310,N_14968,N_14883);
xnor UO_311 (O_311,N_14985,N_14932);
xor UO_312 (O_312,N_14987,N_14850);
nor UO_313 (O_313,N_14984,N_14848);
nor UO_314 (O_314,N_14964,N_14836);
xnor UO_315 (O_315,N_14898,N_14922);
nand UO_316 (O_316,N_14981,N_14994);
or UO_317 (O_317,N_14929,N_14919);
nor UO_318 (O_318,N_14940,N_14913);
or UO_319 (O_319,N_14919,N_14819);
nand UO_320 (O_320,N_14878,N_14957);
and UO_321 (O_321,N_14914,N_14939);
nand UO_322 (O_322,N_14891,N_14820);
nand UO_323 (O_323,N_14997,N_14991);
or UO_324 (O_324,N_14981,N_14869);
nand UO_325 (O_325,N_14856,N_14915);
nor UO_326 (O_326,N_14829,N_14939);
nor UO_327 (O_327,N_14821,N_14904);
nor UO_328 (O_328,N_14921,N_14952);
nor UO_329 (O_329,N_14851,N_14976);
or UO_330 (O_330,N_14992,N_14813);
and UO_331 (O_331,N_14976,N_14896);
and UO_332 (O_332,N_14933,N_14853);
xor UO_333 (O_333,N_14860,N_14814);
or UO_334 (O_334,N_14955,N_14954);
xnor UO_335 (O_335,N_14951,N_14963);
or UO_336 (O_336,N_14928,N_14959);
or UO_337 (O_337,N_14881,N_14826);
nor UO_338 (O_338,N_14864,N_14827);
xor UO_339 (O_339,N_14823,N_14955);
nand UO_340 (O_340,N_14839,N_14855);
nand UO_341 (O_341,N_14831,N_14942);
nor UO_342 (O_342,N_14839,N_14927);
and UO_343 (O_343,N_14869,N_14857);
and UO_344 (O_344,N_14857,N_14922);
nor UO_345 (O_345,N_14921,N_14991);
and UO_346 (O_346,N_14863,N_14977);
nand UO_347 (O_347,N_14982,N_14980);
nor UO_348 (O_348,N_14993,N_14923);
nand UO_349 (O_349,N_14873,N_14860);
nor UO_350 (O_350,N_14801,N_14979);
or UO_351 (O_351,N_14987,N_14808);
or UO_352 (O_352,N_14939,N_14867);
nor UO_353 (O_353,N_14916,N_14907);
nand UO_354 (O_354,N_14980,N_14803);
nor UO_355 (O_355,N_14806,N_14869);
nand UO_356 (O_356,N_14887,N_14970);
nand UO_357 (O_357,N_14887,N_14874);
and UO_358 (O_358,N_14968,N_14985);
nand UO_359 (O_359,N_14860,N_14913);
nand UO_360 (O_360,N_14855,N_14956);
and UO_361 (O_361,N_14967,N_14999);
nand UO_362 (O_362,N_14813,N_14949);
or UO_363 (O_363,N_14890,N_14926);
nor UO_364 (O_364,N_14999,N_14856);
or UO_365 (O_365,N_14884,N_14801);
or UO_366 (O_366,N_14845,N_14897);
nor UO_367 (O_367,N_14815,N_14818);
or UO_368 (O_368,N_14845,N_14862);
nand UO_369 (O_369,N_14853,N_14831);
nor UO_370 (O_370,N_14953,N_14865);
and UO_371 (O_371,N_14885,N_14808);
and UO_372 (O_372,N_14918,N_14862);
or UO_373 (O_373,N_14804,N_14802);
nor UO_374 (O_374,N_14820,N_14887);
nand UO_375 (O_375,N_14845,N_14988);
or UO_376 (O_376,N_14865,N_14948);
and UO_377 (O_377,N_14925,N_14955);
nand UO_378 (O_378,N_14865,N_14981);
nor UO_379 (O_379,N_14803,N_14845);
nand UO_380 (O_380,N_14859,N_14889);
nand UO_381 (O_381,N_14890,N_14936);
and UO_382 (O_382,N_14837,N_14862);
nand UO_383 (O_383,N_14819,N_14957);
and UO_384 (O_384,N_14965,N_14860);
xnor UO_385 (O_385,N_14818,N_14822);
or UO_386 (O_386,N_14917,N_14806);
nand UO_387 (O_387,N_14903,N_14868);
and UO_388 (O_388,N_14843,N_14946);
or UO_389 (O_389,N_14891,N_14926);
and UO_390 (O_390,N_14943,N_14871);
or UO_391 (O_391,N_14844,N_14927);
nor UO_392 (O_392,N_14808,N_14927);
nor UO_393 (O_393,N_14830,N_14982);
nor UO_394 (O_394,N_14941,N_14837);
or UO_395 (O_395,N_14914,N_14950);
nand UO_396 (O_396,N_14835,N_14969);
nand UO_397 (O_397,N_14839,N_14904);
or UO_398 (O_398,N_14932,N_14845);
xor UO_399 (O_399,N_14997,N_14910);
nor UO_400 (O_400,N_14807,N_14867);
nand UO_401 (O_401,N_14947,N_14950);
or UO_402 (O_402,N_14909,N_14918);
nor UO_403 (O_403,N_14827,N_14956);
and UO_404 (O_404,N_14809,N_14826);
nand UO_405 (O_405,N_14945,N_14896);
nor UO_406 (O_406,N_14834,N_14987);
nand UO_407 (O_407,N_14883,N_14879);
nand UO_408 (O_408,N_14840,N_14977);
or UO_409 (O_409,N_14932,N_14875);
or UO_410 (O_410,N_14911,N_14878);
and UO_411 (O_411,N_14946,N_14927);
or UO_412 (O_412,N_14926,N_14921);
xor UO_413 (O_413,N_14802,N_14914);
xor UO_414 (O_414,N_14846,N_14982);
xor UO_415 (O_415,N_14852,N_14929);
nand UO_416 (O_416,N_14861,N_14962);
nand UO_417 (O_417,N_14861,N_14926);
or UO_418 (O_418,N_14972,N_14903);
nor UO_419 (O_419,N_14810,N_14978);
nor UO_420 (O_420,N_14985,N_14807);
or UO_421 (O_421,N_14812,N_14935);
nand UO_422 (O_422,N_14937,N_14949);
nand UO_423 (O_423,N_14844,N_14956);
nand UO_424 (O_424,N_14821,N_14925);
xor UO_425 (O_425,N_14978,N_14965);
or UO_426 (O_426,N_14974,N_14805);
or UO_427 (O_427,N_14856,N_14900);
or UO_428 (O_428,N_14958,N_14913);
and UO_429 (O_429,N_14811,N_14931);
and UO_430 (O_430,N_14857,N_14949);
xor UO_431 (O_431,N_14848,N_14815);
nand UO_432 (O_432,N_14904,N_14859);
or UO_433 (O_433,N_14856,N_14847);
nor UO_434 (O_434,N_14952,N_14978);
and UO_435 (O_435,N_14881,N_14909);
nor UO_436 (O_436,N_14817,N_14800);
nand UO_437 (O_437,N_14812,N_14873);
nor UO_438 (O_438,N_14957,N_14846);
nor UO_439 (O_439,N_14894,N_14985);
nand UO_440 (O_440,N_14854,N_14997);
xor UO_441 (O_441,N_14992,N_14878);
or UO_442 (O_442,N_14904,N_14952);
or UO_443 (O_443,N_14997,N_14840);
nor UO_444 (O_444,N_14937,N_14974);
nand UO_445 (O_445,N_14856,N_14977);
xor UO_446 (O_446,N_14871,N_14817);
and UO_447 (O_447,N_14800,N_14815);
nand UO_448 (O_448,N_14810,N_14850);
nand UO_449 (O_449,N_14854,N_14994);
or UO_450 (O_450,N_14957,N_14857);
nand UO_451 (O_451,N_14833,N_14989);
and UO_452 (O_452,N_14809,N_14933);
nand UO_453 (O_453,N_14888,N_14851);
nor UO_454 (O_454,N_14890,N_14934);
and UO_455 (O_455,N_14900,N_14878);
and UO_456 (O_456,N_14863,N_14821);
nor UO_457 (O_457,N_14849,N_14959);
nor UO_458 (O_458,N_14920,N_14962);
and UO_459 (O_459,N_14873,N_14924);
and UO_460 (O_460,N_14836,N_14842);
or UO_461 (O_461,N_14801,N_14970);
nor UO_462 (O_462,N_14816,N_14806);
xor UO_463 (O_463,N_14904,N_14921);
nor UO_464 (O_464,N_14903,N_14982);
nand UO_465 (O_465,N_14800,N_14910);
nor UO_466 (O_466,N_14822,N_14819);
xor UO_467 (O_467,N_14950,N_14930);
nor UO_468 (O_468,N_14823,N_14886);
or UO_469 (O_469,N_14980,N_14932);
nor UO_470 (O_470,N_14905,N_14963);
and UO_471 (O_471,N_14946,N_14894);
or UO_472 (O_472,N_14816,N_14935);
or UO_473 (O_473,N_14898,N_14891);
and UO_474 (O_474,N_14887,N_14808);
and UO_475 (O_475,N_14999,N_14826);
or UO_476 (O_476,N_14986,N_14918);
nor UO_477 (O_477,N_14801,N_14909);
nor UO_478 (O_478,N_14895,N_14887);
and UO_479 (O_479,N_14811,N_14817);
and UO_480 (O_480,N_14857,N_14889);
or UO_481 (O_481,N_14939,N_14898);
xnor UO_482 (O_482,N_14840,N_14875);
or UO_483 (O_483,N_14933,N_14837);
nand UO_484 (O_484,N_14883,N_14855);
nand UO_485 (O_485,N_14956,N_14886);
and UO_486 (O_486,N_14937,N_14828);
nand UO_487 (O_487,N_14850,N_14858);
or UO_488 (O_488,N_14855,N_14985);
nor UO_489 (O_489,N_14818,N_14821);
or UO_490 (O_490,N_14965,N_14888);
xnor UO_491 (O_491,N_14883,N_14940);
and UO_492 (O_492,N_14905,N_14981);
nor UO_493 (O_493,N_14850,N_14974);
nand UO_494 (O_494,N_14975,N_14842);
and UO_495 (O_495,N_14833,N_14995);
nand UO_496 (O_496,N_14931,N_14841);
or UO_497 (O_497,N_14833,N_14980);
nand UO_498 (O_498,N_14909,N_14921);
nand UO_499 (O_499,N_14878,N_14959);
and UO_500 (O_500,N_14934,N_14809);
nor UO_501 (O_501,N_14812,N_14864);
and UO_502 (O_502,N_14998,N_14939);
or UO_503 (O_503,N_14889,N_14968);
xor UO_504 (O_504,N_14807,N_14908);
nand UO_505 (O_505,N_14998,N_14856);
nand UO_506 (O_506,N_14994,N_14836);
or UO_507 (O_507,N_14998,N_14846);
or UO_508 (O_508,N_14940,N_14867);
and UO_509 (O_509,N_14818,N_14990);
and UO_510 (O_510,N_14844,N_14835);
nor UO_511 (O_511,N_14837,N_14895);
xor UO_512 (O_512,N_14810,N_14995);
nor UO_513 (O_513,N_14980,N_14974);
nand UO_514 (O_514,N_14942,N_14885);
nor UO_515 (O_515,N_14810,N_14875);
and UO_516 (O_516,N_14867,N_14925);
or UO_517 (O_517,N_14855,N_14951);
nand UO_518 (O_518,N_14836,N_14919);
and UO_519 (O_519,N_14841,N_14911);
or UO_520 (O_520,N_14851,N_14994);
nand UO_521 (O_521,N_14957,N_14923);
nor UO_522 (O_522,N_14927,N_14962);
xnor UO_523 (O_523,N_14839,N_14907);
and UO_524 (O_524,N_14992,N_14838);
nand UO_525 (O_525,N_14877,N_14882);
xor UO_526 (O_526,N_14931,N_14918);
and UO_527 (O_527,N_14946,N_14905);
or UO_528 (O_528,N_14949,N_14996);
and UO_529 (O_529,N_14902,N_14855);
and UO_530 (O_530,N_14937,N_14926);
or UO_531 (O_531,N_14835,N_14831);
and UO_532 (O_532,N_14909,N_14968);
xor UO_533 (O_533,N_14939,N_14955);
or UO_534 (O_534,N_14901,N_14866);
xnor UO_535 (O_535,N_14877,N_14978);
nor UO_536 (O_536,N_14830,N_14916);
and UO_537 (O_537,N_14907,N_14968);
or UO_538 (O_538,N_14863,N_14861);
nand UO_539 (O_539,N_14821,N_14879);
nor UO_540 (O_540,N_14947,N_14967);
and UO_541 (O_541,N_14988,N_14822);
or UO_542 (O_542,N_14925,N_14965);
nand UO_543 (O_543,N_14828,N_14815);
nand UO_544 (O_544,N_14911,N_14915);
or UO_545 (O_545,N_14805,N_14832);
and UO_546 (O_546,N_14888,N_14902);
and UO_547 (O_547,N_14835,N_14919);
or UO_548 (O_548,N_14920,N_14874);
nand UO_549 (O_549,N_14977,N_14892);
and UO_550 (O_550,N_14986,N_14838);
nor UO_551 (O_551,N_14819,N_14812);
and UO_552 (O_552,N_14880,N_14989);
nor UO_553 (O_553,N_14809,N_14878);
nor UO_554 (O_554,N_14870,N_14949);
or UO_555 (O_555,N_14917,N_14897);
nand UO_556 (O_556,N_14972,N_14971);
or UO_557 (O_557,N_14996,N_14915);
nand UO_558 (O_558,N_14929,N_14959);
nor UO_559 (O_559,N_14882,N_14921);
nor UO_560 (O_560,N_14821,N_14956);
or UO_561 (O_561,N_14903,N_14866);
nor UO_562 (O_562,N_14856,N_14834);
nor UO_563 (O_563,N_14955,N_14914);
nor UO_564 (O_564,N_14945,N_14808);
nand UO_565 (O_565,N_14812,N_14823);
or UO_566 (O_566,N_14831,N_14802);
nand UO_567 (O_567,N_14846,N_14841);
nand UO_568 (O_568,N_14946,N_14924);
and UO_569 (O_569,N_14953,N_14902);
xnor UO_570 (O_570,N_14867,N_14992);
and UO_571 (O_571,N_14988,N_14993);
or UO_572 (O_572,N_14882,N_14967);
nand UO_573 (O_573,N_14909,N_14862);
and UO_574 (O_574,N_14993,N_14810);
and UO_575 (O_575,N_14805,N_14844);
nand UO_576 (O_576,N_14936,N_14851);
nand UO_577 (O_577,N_14843,N_14949);
nor UO_578 (O_578,N_14919,N_14942);
nor UO_579 (O_579,N_14866,N_14925);
and UO_580 (O_580,N_14841,N_14847);
nor UO_581 (O_581,N_14983,N_14817);
nor UO_582 (O_582,N_14882,N_14929);
xor UO_583 (O_583,N_14987,N_14894);
nor UO_584 (O_584,N_14882,N_14926);
or UO_585 (O_585,N_14945,N_14900);
and UO_586 (O_586,N_14805,N_14920);
nor UO_587 (O_587,N_14987,N_14981);
nand UO_588 (O_588,N_14820,N_14827);
nor UO_589 (O_589,N_14857,N_14986);
xor UO_590 (O_590,N_14861,N_14800);
and UO_591 (O_591,N_14981,N_14948);
and UO_592 (O_592,N_14922,N_14809);
nand UO_593 (O_593,N_14807,N_14895);
xor UO_594 (O_594,N_14895,N_14843);
and UO_595 (O_595,N_14944,N_14947);
nor UO_596 (O_596,N_14836,N_14983);
or UO_597 (O_597,N_14952,N_14977);
nand UO_598 (O_598,N_14808,N_14878);
nand UO_599 (O_599,N_14935,N_14879);
nand UO_600 (O_600,N_14930,N_14925);
or UO_601 (O_601,N_14904,N_14846);
nand UO_602 (O_602,N_14961,N_14853);
or UO_603 (O_603,N_14880,N_14808);
or UO_604 (O_604,N_14935,N_14929);
or UO_605 (O_605,N_14840,N_14973);
nor UO_606 (O_606,N_14822,N_14862);
and UO_607 (O_607,N_14962,N_14845);
and UO_608 (O_608,N_14951,N_14991);
xnor UO_609 (O_609,N_14902,N_14998);
nor UO_610 (O_610,N_14890,N_14801);
or UO_611 (O_611,N_14811,N_14859);
nand UO_612 (O_612,N_14909,N_14943);
or UO_613 (O_613,N_14862,N_14846);
nand UO_614 (O_614,N_14926,N_14929);
nand UO_615 (O_615,N_14872,N_14839);
or UO_616 (O_616,N_14847,N_14807);
and UO_617 (O_617,N_14910,N_14932);
and UO_618 (O_618,N_14954,N_14912);
and UO_619 (O_619,N_14902,N_14828);
nand UO_620 (O_620,N_14883,N_14891);
xnor UO_621 (O_621,N_14861,N_14940);
nor UO_622 (O_622,N_14928,N_14936);
xnor UO_623 (O_623,N_14846,N_14806);
nand UO_624 (O_624,N_14814,N_14827);
and UO_625 (O_625,N_14903,N_14824);
xnor UO_626 (O_626,N_14992,N_14810);
nor UO_627 (O_627,N_14827,N_14972);
or UO_628 (O_628,N_14991,N_14837);
xnor UO_629 (O_629,N_14949,N_14800);
nand UO_630 (O_630,N_14867,N_14846);
and UO_631 (O_631,N_14928,N_14942);
nand UO_632 (O_632,N_14848,N_14852);
and UO_633 (O_633,N_14856,N_14805);
or UO_634 (O_634,N_14896,N_14981);
and UO_635 (O_635,N_14940,N_14979);
and UO_636 (O_636,N_14901,N_14823);
and UO_637 (O_637,N_14875,N_14805);
or UO_638 (O_638,N_14802,N_14937);
nor UO_639 (O_639,N_14865,N_14964);
and UO_640 (O_640,N_14950,N_14991);
or UO_641 (O_641,N_14889,N_14896);
or UO_642 (O_642,N_14916,N_14993);
and UO_643 (O_643,N_14998,N_14961);
nor UO_644 (O_644,N_14955,N_14887);
and UO_645 (O_645,N_14948,N_14954);
or UO_646 (O_646,N_14867,N_14835);
and UO_647 (O_647,N_14998,N_14866);
or UO_648 (O_648,N_14997,N_14967);
nand UO_649 (O_649,N_14909,N_14979);
and UO_650 (O_650,N_14878,N_14926);
and UO_651 (O_651,N_14808,N_14957);
nand UO_652 (O_652,N_14969,N_14911);
or UO_653 (O_653,N_14806,N_14938);
or UO_654 (O_654,N_14874,N_14867);
nor UO_655 (O_655,N_14966,N_14982);
xor UO_656 (O_656,N_14860,N_14935);
or UO_657 (O_657,N_14913,N_14968);
nand UO_658 (O_658,N_14953,N_14822);
nand UO_659 (O_659,N_14936,N_14995);
nor UO_660 (O_660,N_14921,N_14821);
or UO_661 (O_661,N_14880,N_14814);
or UO_662 (O_662,N_14996,N_14807);
nor UO_663 (O_663,N_14876,N_14821);
or UO_664 (O_664,N_14950,N_14833);
or UO_665 (O_665,N_14876,N_14933);
nor UO_666 (O_666,N_14902,N_14832);
nand UO_667 (O_667,N_14899,N_14909);
nor UO_668 (O_668,N_14833,N_14917);
xor UO_669 (O_669,N_14960,N_14831);
nand UO_670 (O_670,N_14913,N_14912);
and UO_671 (O_671,N_14832,N_14845);
nor UO_672 (O_672,N_14806,N_14800);
and UO_673 (O_673,N_14889,N_14996);
and UO_674 (O_674,N_14885,N_14857);
nand UO_675 (O_675,N_14855,N_14807);
nor UO_676 (O_676,N_14802,N_14930);
nand UO_677 (O_677,N_14877,N_14975);
nand UO_678 (O_678,N_14833,N_14893);
or UO_679 (O_679,N_14910,N_14905);
nor UO_680 (O_680,N_14865,N_14895);
and UO_681 (O_681,N_14945,N_14957);
or UO_682 (O_682,N_14839,N_14838);
or UO_683 (O_683,N_14900,N_14844);
nor UO_684 (O_684,N_14987,N_14966);
nand UO_685 (O_685,N_14886,N_14948);
nor UO_686 (O_686,N_14947,N_14959);
and UO_687 (O_687,N_14895,N_14846);
nor UO_688 (O_688,N_14817,N_14942);
nor UO_689 (O_689,N_14810,N_14931);
and UO_690 (O_690,N_14932,N_14827);
nor UO_691 (O_691,N_14933,N_14932);
and UO_692 (O_692,N_14849,N_14833);
or UO_693 (O_693,N_14855,N_14880);
and UO_694 (O_694,N_14906,N_14975);
xnor UO_695 (O_695,N_14806,N_14972);
or UO_696 (O_696,N_14872,N_14961);
and UO_697 (O_697,N_14949,N_14824);
nand UO_698 (O_698,N_14839,N_14813);
xor UO_699 (O_699,N_14965,N_14889);
and UO_700 (O_700,N_14850,N_14851);
nand UO_701 (O_701,N_14862,N_14891);
nand UO_702 (O_702,N_14913,N_14804);
nand UO_703 (O_703,N_14921,N_14806);
and UO_704 (O_704,N_14992,N_14982);
or UO_705 (O_705,N_14980,N_14834);
or UO_706 (O_706,N_14948,N_14877);
xor UO_707 (O_707,N_14818,N_14980);
nand UO_708 (O_708,N_14937,N_14845);
xor UO_709 (O_709,N_14898,N_14907);
and UO_710 (O_710,N_14987,N_14943);
or UO_711 (O_711,N_14879,N_14885);
nand UO_712 (O_712,N_14926,N_14886);
nor UO_713 (O_713,N_14805,N_14979);
nor UO_714 (O_714,N_14808,N_14841);
and UO_715 (O_715,N_14850,N_14932);
nor UO_716 (O_716,N_14824,N_14986);
or UO_717 (O_717,N_14832,N_14962);
xor UO_718 (O_718,N_14923,N_14906);
xor UO_719 (O_719,N_14857,N_14840);
or UO_720 (O_720,N_14822,N_14816);
nand UO_721 (O_721,N_14876,N_14944);
or UO_722 (O_722,N_14875,N_14967);
nor UO_723 (O_723,N_14897,N_14982);
or UO_724 (O_724,N_14973,N_14854);
nor UO_725 (O_725,N_14994,N_14925);
and UO_726 (O_726,N_14815,N_14860);
nand UO_727 (O_727,N_14919,N_14968);
xor UO_728 (O_728,N_14973,N_14936);
and UO_729 (O_729,N_14846,N_14905);
or UO_730 (O_730,N_14844,N_14810);
nor UO_731 (O_731,N_14808,N_14883);
nand UO_732 (O_732,N_14946,N_14933);
nand UO_733 (O_733,N_14800,N_14987);
or UO_734 (O_734,N_14986,N_14964);
nand UO_735 (O_735,N_14894,N_14960);
and UO_736 (O_736,N_14855,N_14882);
nor UO_737 (O_737,N_14961,N_14836);
nor UO_738 (O_738,N_14815,N_14866);
and UO_739 (O_739,N_14927,N_14878);
or UO_740 (O_740,N_14831,N_14981);
and UO_741 (O_741,N_14982,N_14831);
or UO_742 (O_742,N_14954,N_14911);
nand UO_743 (O_743,N_14911,N_14887);
or UO_744 (O_744,N_14811,N_14823);
and UO_745 (O_745,N_14935,N_14825);
nand UO_746 (O_746,N_14807,N_14891);
nor UO_747 (O_747,N_14986,N_14944);
and UO_748 (O_748,N_14876,N_14982);
nand UO_749 (O_749,N_14910,N_14836);
or UO_750 (O_750,N_14887,N_14872);
and UO_751 (O_751,N_14884,N_14874);
or UO_752 (O_752,N_14891,N_14980);
and UO_753 (O_753,N_14969,N_14959);
nor UO_754 (O_754,N_14911,N_14811);
xor UO_755 (O_755,N_14811,N_14922);
nand UO_756 (O_756,N_14990,N_14831);
and UO_757 (O_757,N_14919,N_14932);
nor UO_758 (O_758,N_14942,N_14876);
nor UO_759 (O_759,N_14869,N_14812);
or UO_760 (O_760,N_14879,N_14905);
and UO_761 (O_761,N_14865,N_14804);
and UO_762 (O_762,N_14960,N_14861);
and UO_763 (O_763,N_14848,N_14866);
and UO_764 (O_764,N_14817,N_14946);
nand UO_765 (O_765,N_14942,N_14900);
nor UO_766 (O_766,N_14806,N_14805);
nand UO_767 (O_767,N_14982,N_14856);
nor UO_768 (O_768,N_14948,N_14900);
nor UO_769 (O_769,N_14880,N_14866);
and UO_770 (O_770,N_14873,N_14880);
xor UO_771 (O_771,N_14907,N_14868);
nand UO_772 (O_772,N_14945,N_14829);
and UO_773 (O_773,N_14943,N_14818);
xnor UO_774 (O_774,N_14807,N_14889);
or UO_775 (O_775,N_14945,N_14932);
nor UO_776 (O_776,N_14959,N_14867);
and UO_777 (O_777,N_14830,N_14993);
nor UO_778 (O_778,N_14938,N_14842);
nand UO_779 (O_779,N_14953,N_14952);
and UO_780 (O_780,N_14861,N_14906);
xnor UO_781 (O_781,N_14909,N_14805);
or UO_782 (O_782,N_14950,N_14925);
or UO_783 (O_783,N_14998,N_14994);
xnor UO_784 (O_784,N_14922,N_14935);
or UO_785 (O_785,N_14999,N_14890);
nand UO_786 (O_786,N_14923,N_14891);
and UO_787 (O_787,N_14835,N_14955);
xnor UO_788 (O_788,N_14979,N_14864);
xor UO_789 (O_789,N_14879,N_14803);
or UO_790 (O_790,N_14835,N_14957);
or UO_791 (O_791,N_14812,N_14862);
nand UO_792 (O_792,N_14853,N_14912);
nor UO_793 (O_793,N_14979,N_14957);
nand UO_794 (O_794,N_14879,N_14853);
nand UO_795 (O_795,N_14970,N_14865);
nor UO_796 (O_796,N_14882,N_14951);
nor UO_797 (O_797,N_14801,N_14904);
or UO_798 (O_798,N_14951,N_14914);
nor UO_799 (O_799,N_14962,N_14851);
nand UO_800 (O_800,N_14908,N_14800);
and UO_801 (O_801,N_14982,N_14916);
and UO_802 (O_802,N_14839,N_14994);
nor UO_803 (O_803,N_14809,N_14955);
xor UO_804 (O_804,N_14922,N_14911);
nor UO_805 (O_805,N_14952,N_14837);
xnor UO_806 (O_806,N_14919,N_14833);
nor UO_807 (O_807,N_14929,N_14955);
nor UO_808 (O_808,N_14893,N_14928);
nand UO_809 (O_809,N_14934,N_14988);
xor UO_810 (O_810,N_14850,N_14982);
xnor UO_811 (O_811,N_14812,N_14996);
and UO_812 (O_812,N_14839,N_14965);
or UO_813 (O_813,N_14831,N_14888);
xnor UO_814 (O_814,N_14828,N_14925);
or UO_815 (O_815,N_14915,N_14813);
nor UO_816 (O_816,N_14828,N_14944);
xnor UO_817 (O_817,N_14956,N_14945);
nand UO_818 (O_818,N_14806,N_14892);
nand UO_819 (O_819,N_14824,N_14923);
or UO_820 (O_820,N_14860,N_14943);
nor UO_821 (O_821,N_14951,N_14968);
nand UO_822 (O_822,N_14831,N_14970);
nand UO_823 (O_823,N_14938,N_14966);
nand UO_824 (O_824,N_14979,N_14989);
nand UO_825 (O_825,N_14856,N_14916);
and UO_826 (O_826,N_14946,N_14995);
nor UO_827 (O_827,N_14856,N_14948);
nand UO_828 (O_828,N_14977,N_14873);
and UO_829 (O_829,N_14815,N_14833);
nor UO_830 (O_830,N_14816,N_14857);
or UO_831 (O_831,N_14888,N_14916);
or UO_832 (O_832,N_14993,N_14945);
and UO_833 (O_833,N_14933,N_14940);
and UO_834 (O_834,N_14949,N_14979);
or UO_835 (O_835,N_14933,N_14834);
nand UO_836 (O_836,N_14801,N_14812);
nor UO_837 (O_837,N_14983,N_14841);
or UO_838 (O_838,N_14985,N_14954);
nor UO_839 (O_839,N_14985,N_14802);
xnor UO_840 (O_840,N_14889,N_14800);
or UO_841 (O_841,N_14948,N_14951);
nand UO_842 (O_842,N_14869,N_14890);
nand UO_843 (O_843,N_14944,N_14981);
xor UO_844 (O_844,N_14899,N_14938);
nand UO_845 (O_845,N_14932,N_14822);
nor UO_846 (O_846,N_14950,N_14826);
nand UO_847 (O_847,N_14895,N_14855);
nor UO_848 (O_848,N_14943,N_14983);
nor UO_849 (O_849,N_14917,N_14998);
nand UO_850 (O_850,N_14997,N_14865);
and UO_851 (O_851,N_14949,N_14989);
and UO_852 (O_852,N_14833,N_14826);
and UO_853 (O_853,N_14878,N_14840);
nand UO_854 (O_854,N_14815,N_14942);
and UO_855 (O_855,N_14966,N_14810);
xnor UO_856 (O_856,N_14990,N_14840);
and UO_857 (O_857,N_14971,N_14964);
nand UO_858 (O_858,N_14975,N_14917);
and UO_859 (O_859,N_14942,N_14911);
xnor UO_860 (O_860,N_14908,N_14919);
nand UO_861 (O_861,N_14827,N_14897);
or UO_862 (O_862,N_14927,N_14818);
or UO_863 (O_863,N_14882,N_14994);
xor UO_864 (O_864,N_14970,N_14858);
nor UO_865 (O_865,N_14926,N_14823);
or UO_866 (O_866,N_14811,N_14853);
and UO_867 (O_867,N_14877,N_14898);
and UO_868 (O_868,N_14899,N_14885);
nor UO_869 (O_869,N_14879,N_14925);
nor UO_870 (O_870,N_14915,N_14918);
nor UO_871 (O_871,N_14952,N_14930);
xor UO_872 (O_872,N_14835,N_14828);
nand UO_873 (O_873,N_14960,N_14835);
nand UO_874 (O_874,N_14821,N_14934);
and UO_875 (O_875,N_14848,N_14807);
nor UO_876 (O_876,N_14813,N_14969);
and UO_877 (O_877,N_14837,N_14956);
or UO_878 (O_878,N_14907,N_14810);
xnor UO_879 (O_879,N_14886,N_14855);
or UO_880 (O_880,N_14973,N_14842);
or UO_881 (O_881,N_14859,N_14956);
and UO_882 (O_882,N_14823,N_14803);
and UO_883 (O_883,N_14931,N_14993);
or UO_884 (O_884,N_14840,N_14992);
nand UO_885 (O_885,N_14968,N_14922);
and UO_886 (O_886,N_14880,N_14810);
and UO_887 (O_887,N_14974,N_14994);
xnor UO_888 (O_888,N_14890,N_14805);
and UO_889 (O_889,N_14975,N_14960);
nor UO_890 (O_890,N_14810,N_14936);
nand UO_891 (O_891,N_14927,N_14831);
nand UO_892 (O_892,N_14950,N_14824);
and UO_893 (O_893,N_14920,N_14953);
nor UO_894 (O_894,N_14924,N_14938);
nand UO_895 (O_895,N_14948,N_14878);
nand UO_896 (O_896,N_14838,N_14966);
or UO_897 (O_897,N_14860,N_14914);
or UO_898 (O_898,N_14857,N_14865);
nand UO_899 (O_899,N_14868,N_14894);
or UO_900 (O_900,N_14926,N_14904);
xnor UO_901 (O_901,N_14897,N_14849);
or UO_902 (O_902,N_14910,N_14968);
nor UO_903 (O_903,N_14931,N_14942);
nor UO_904 (O_904,N_14901,N_14821);
and UO_905 (O_905,N_14930,N_14955);
nor UO_906 (O_906,N_14963,N_14993);
and UO_907 (O_907,N_14869,N_14839);
nand UO_908 (O_908,N_14871,N_14899);
nor UO_909 (O_909,N_14932,N_14847);
nand UO_910 (O_910,N_14925,N_14927);
nor UO_911 (O_911,N_14997,N_14987);
and UO_912 (O_912,N_14889,N_14887);
xor UO_913 (O_913,N_14997,N_14800);
or UO_914 (O_914,N_14845,N_14809);
and UO_915 (O_915,N_14820,N_14888);
nor UO_916 (O_916,N_14835,N_14892);
and UO_917 (O_917,N_14933,N_14881);
nor UO_918 (O_918,N_14858,N_14946);
and UO_919 (O_919,N_14900,N_14936);
nand UO_920 (O_920,N_14861,N_14888);
and UO_921 (O_921,N_14818,N_14846);
nand UO_922 (O_922,N_14982,N_14880);
and UO_923 (O_923,N_14918,N_14903);
and UO_924 (O_924,N_14910,N_14825);
nand UO_925 (O_925,N_14965,N_14896);
and UO_926 (O_926,N_14813,N_14847);
nand UO_927 (O_927,N_14983,N_14979);
nand UO_928 (O_928,N_14855,N_14946);
and UO_929 (O_929,N_14878,N_14811);
or UO_930 (O_930,N_14923,N_14946);
or UO_931 (O_931,N_14818,N_14853);
nor UO_932 (O_932,N_14916,N_14800);
or UO_933 (O_933,N_14860,N_14911);
nand UO_934 (O_934,N_14967,N_14889);
and UO_935 (O_935,N_14990,N_14955);
nand UO_936 (O_936,N_14831,N_14874);
xor UO_937 (O_937,N_14834,N_14938);
and UO_938 (O_938,N_14884,N_14811);
nand UO_939 (O_939,N_14882,N_14819);
and UO_940 (O_940,N_14903,N_14818);
xor UO_941 (O_941,N_14951,N_14957);
or UO_942 (O_942,N_14862,N_14902);
or UO_943 (O_943,N_14930,N_14966);
nor UO_944 (O_944,N_14887,N_14825);
xnor UO_945 (O_945,N_14964,N_14830);
nor UO_946 (O_946,N_14815,N_14851);
and UO_947 (O_947,N_14861,N_14829);
xnor UO_948 (O_948,N_14901,N_14910);
nor UO_949 (O_949,N_14813,N_14973);
and UO_950 (O_950,N_14820,N_14814);
or UO_951 (O_951,N_14999,N_14877);
and UO_952 (O_952,N_14962,N_14989);
nor UO_953 (O_953,N_14887,N_14806);
nor UO_954 (O_954,N_14859,N_14936);
or UO_955 (O_955,N_14855,N_14856);
or UO_956 (O_956,N_14928,N_14819);
nand UO_957 (O_957,N_14856,N_14833);
xnor UO_958 (O_958,N_14815,N_14936);
nand UO_959 (O_959,N_14813,N_14911);
xor UO_960 (O_960,N_14891,N_14878);
xor UO_961 (O_961,N_14948,N_14987);
and UO_962 (O_962,N_14847,N_14960);
xnor UO_963 (O_963,N_14870,N_14922);
and UO_964 (O_964,N_14897,N_14944);
and UO_965 (O_965,N_14823,N_14975);
or UO_966 (O_966,N_14944,N_14811);
nand UO_967 (O_967,N_14890,N_14881);
and UO_968 (O_968,N_14940,N_14866);
and UO_969 (O_969,N_14859,N_14877);
nand UO_970 (O_970,N_14976,N_14802);
nand UO_971 (O_971,N_14964,N_14938);
xor UO_972 (O_972,N_14822,N_14881);
and UO_973 (O_973,N_14885,N_14969);
nand UO_974 (O_974,N_14870,N_14997);
nor UO_975 (O_975,N_14851,N_14895);
nor UO_976 (O_976,N_14885,N_14987);
and UO_977 (O_977,N_14925,N_14800);
or UO_978 (O_978,N_14998,N_14868);
nand UO_979 (O_979,N_14846,N_14871);
and UO_980 (O_980,N_14897,N_14814);
and UO_981 (O_981,N_14995,N_14842);
xnor UO_982 (O_982,N_14863,N_14850);
xor UO_983 (O_983,N_14913,N_14809);
nand UO_984 (O_984,N_14930,N_14885);
xor UO_985 (O_985,N_14942,N_14906);
xor UO_986 (O_986,N_14859,N_14967);
xor UO_987 (O_987,N_14948,N_14889);
or UO_988 (O_988,N_14943,N_14924);
nand UO_989 (O_989,N_14823,N_14862);
and UO_990 (O_990,N_14985,N_14996);
or UO_991 (O_991,N_14919,N_14937);
or UO_992 (O_992,N_14804,N_14995);
nor UO_993 (O_993,N_14872,N_14907);
and UO_994 (O_994,N_14845,N_14933);
or UO_995 (O_995,N_14993,N_14811);
nand UO_996 (O_996,N_14920,N_14836);
or UO_997 (O_997,N_14892,N_14881);
nor UO_998 (O_998,N_14840,N_14807);
and UO_999 (O_999,N_14870,N_14970);
nand UO_1000 (O_1000,N_14874,N_14897);
or UO_1001 (O_1001,N_14860,N_14991);
and UO_1002 (O_1002,N_14956,N_14959);
nor UO_1003 (O_1003,N_14839,N_14818);
and UO_1004 (O_1004,N_14982,N_14853);
or UO_1005 (O_1005,N_14934,N_14904);
nand UO_1006 (O_1006,N_14969,N_14956);
nor UO_1007 (O_1007,N_14830,N_14883);
nand UO_1008 (O_1008,N_14935,N_14866);
nand UO_1009 (O_1009,N_14880,N_14979);
xor UO_1010 (O_1010,N_14835,N_14971);
or UO_1011 (O_1011,N_14898,N_14863);
nor UO_1012 (O_1012,N_14987,N_14918);
xnor UO_1013 (O_1013,N_14972,N_14975);
nor UO_1014 (O_1014,N_14931,N_14955);
nand UO_1015 (O_1015,N_14982,N_14821);
nor UO_1016 (O_1016,N_14904,N_14950);
nor UO_1017 (O_1017,N_14813,N_14951);
nor UO_1018 (O_1018,N_14973,N_14947);
or UO_1019 (O_1019,N_14924,N_14916);
or UO_1020 (O_1020,N_14962,N_14990);
and UO_1021 (O_1021,N_14832,N_14884);
or UO_1022 (O_1022,N_14973,N_14929);
nor UO_1023 (O_1023,N_14947,N_14834);
nand UO_1024 (O_1024,N_14858,N_14967);
nand UO_1025 (O_1025,N_14984,N_14843);
and UO_1026 (O_1026,N_14990,N_14961);
or UO_1027 (O_1027,N_14912,N_14940);
or UO_1028 (O_1028,N_14939,N_14996);
nand UO_1029 (O_1029,N_14976,N_14906);
nor UO_1030 (O_1030,N_14867,N_14853);
or UO_1031 (O_1031,N_14852,N_14800);
or UO_1032 (O_1032,N_14935,N_14995);
nor UO_1033 (O_1033,N_14967,N_14872);
xor UO_1034 (O_1034,N_14871,N_14984);
nand UO_1035 (O_1035,N_14965,N_14800);
and UO_1036 (O_1036,N_14881,N_14946);
xor UO_1037 (O_1037,N_14830,N_14929);
or UO_1038 (O_1038,N_14843,N_14834);
nand UO_1039 (O_1039,N_14922,N_14993);
or UO_1040 (O_1040,N_14914,N_14861);
nand UO_1041 (O_1041,N_14857,N_14892);
and UO_1042 (O_1042,N_14985,N_14982);
and UO_1043 (O_1043,N_14859,N_14810);
or UO_1044 (O_1044,N_14932,N_14884);
nor UO_1045 (O_1045,N_14832,N_14955);
nand UO_1046 (O_1046,N_14932,N_14937);
or UO_1047 (O_1047,N_14896,N_14809);
or UO_1048 (O_1048,N_14893,N_14937);
nor UO_1049 (O_1049,N_14978,N_14928);
or UO_1050 (O_1050,N_14814,N_14937);
or UO_1051 (O_1051,N_14820,N_14935);
or UO_1052 (O_1052,N_14998,N_14967);
nor UO_1053 (O_1053,N_14951,N_14986);
or UO_1054 (O_1054,N_14925,N_14877);
and UO_1055 (O_1055,N_14950,N_14988);
nor UO_1056 (O_1056,N_14806,N_14943);
nand UO_1057 (O_1057,N_14862,N_14811);
or UO_1058 (O_1058,N_14957,N_14856);
and UO_1059 (O_1059,N_14977,N_14817);
nand UO_1060 (O_1060,N_14821,N_14944);
nor UO_1061 (O_1061,N_14877,N_14987);
and UO_1062 (O_1062,N_14962,N_14965);
nand UO_1063 (O_1063,N_14874,N_14956);
nor UO_1064 (O_1064,N_14861,N_14987);
nand UO_1065 (O_1065,N_14926,N_14966);
nand UO_1066 (O_1066,N_14890,N_14921);
nor UO_1067 (O_1067,N_14936,N_14933);
and UO_1068 (O_1068,N_14823,N_14897);
xnor UO_1069 (O_1069,N_14917,N_14944);
nor UO_1070 (O_1070,N_14832,N_14828);
nor UO_1071 (O_1071,N_14878,N_14826);
nor UO_1072 (O_1072,N_14968,N_14997);
or UO_1073 (O_1073,N_14829,N_14862);
nand UO_1074 (O_1074,N_14958,N_14886);
nand UO_1075 (O_1075,N_14857,N_14960);
and UO_1076 (O_1076,N_14919,N_14807);
nand UO_1077 (O_1077,N_14973,N_14956);
or UO_1078 (O_1078,N_14941,N_14858);
nand UO_1079 (O_1079,N_14946,N_14916);
and UO_1080 (O_1080,N_14958,N_14901);
nor UO_1081 (O_1081,N_14923,N_14830);
xnor UO_1082 (O_1082,N_14883,N_14807);
nor UO_1083 (O_1083,N_14972,N_14835);
and UO_1084 (O_1084,N_14853,N_14876);
or UO_1085 (O_1085,N_14857,N_14876);
nand UO_1086 (O_1086,N_14818,N_14850);
and UO_1087 (O_1087,N_14854,N_14934);
nor UO_1088 (O_1088,N_14854,N_14968);
and UO_1089 (O_1089,N_14896,N_14836);
and UO_1090 (O_1090,N_14982,N_14872);
nand UO_1091 (O_1091,N_14912,N_14885);
or UO_1092 (O_1092,N_14890,N_14927);
or UO_1093 (O_1093,N_14807,N_14821);
nand UO_1094 (O_1094,N_14933,N_14948);
or UO_1095 (O_1095,N_14928,N_14938);
nand UO_1096 (O_1096,N_14862,N_14954);
or UO_1097 (O_1097,N_14852,N_14822);
or UO_1098 (O_1098,N_14841,N_14856);
nor UO_1099 (O_1099,N_14863,N_14876);
xor UO_1100 (O_1100,N_14841,N_14850);
nor UO_1101 (O_1101,N_14903,N_14829);
and UO_1102 (O_1102,N_14886,N_14842);
or UO_1103 (O_1103,N_14882,N_14808);
xor UO_1104 (O_1104,N_14868,N_14886);
xor UO_1105 (O_1105,N_14830,N_14846);
nor UO_1106 (O_1106,N_14918,N_14838);
nand UO_1107 (O_1107,N_14983,N_14842);
and UO_1108 (O_1108,N_14849,N_14953);
and UO_1109 (O_1109,N_14931,N_14971);
or UO_1110 (O_1110,N_14956,N_14802);
xnor UO_1111 (O_1111,N_14809,N_14815);
xor UO_1112 (O_1112,N_14975,N_14929);
nor UO_1113 (O_1113,N_14847,N_14801);
or UO_1114 (O_1114,N_14879,N_14916);
or UO_1115 (O_1115,N_14822,N_14805);
or UO_1116 (O_1116,N_14873,N_14813);
or UO_1117 (O_1117,N_14847,N_14902);
or UO_1118 (O_1118,N_14843,N_14865);
nor UO_1119 (O_1119,N_14959,N_14955);
or UO_1120 (O_1120,N_14883,N_14970);
and UO_1121 (O_1121,N_14909,N_14931);
or UO_1122 (O_1122,N_14951,N_14852);
nand UO_1123 (O_1123,N_14963,N_14929);
and UO_1124 (O_1124,N_14860,N_14902);
xnor UO_1125 (O_1125,N_14936,N_14802);
xor UO_1126 (O_1126,N_14834,N_14976);
or UO_1127 (O_1127,N_14938,N_14920);
and UO_1128 (O_1128,N_14866,N_14983);
nand UO_1129 (O_1129,N_14948,N_14805);
nor UO_1130 (O_1130,N_14873,N_14962);
nor UO_1131 (O_1131,N_14936,N_14839);
and UO_1132 (O_1132,N_14931,N_14826);
xor UO_1133 (O_1133,N_14988,N_14821);
nand UO_1134 (O_1134,N_14878,N_14952);
and UO_1135 (O_1135,N_14898,N_14967);
nand UO_1136 (O_1136,N_14942,N_14865);
and UO_1137 (O_1137,N_14896,N_14866);
xnor UO_1138 (O_1138,N_14823,N_14877);
or UO_1139 (O_1139,N_14830,N_14991);
or UO_1140 (O_1140,N_14819,N_14937);
or UO_1141 (O_1141,N_14898,N_14903);
and UO_1142 (O_1142,N_14904,N_14837);
nor UO_1143 (O_1143,N_14983,N_14886);
and UO_1144 (O_1144,N_14802,N_14864);
or UO_1145 (O_1145,N_14940,N_14948);
nor UO_1146 (O_1146,N_14820,N_14862);
xor UO_1147 (O_1147,N_14966,N_14848);
or UO_1148 (O_1148,N_14972,N_14973);
and UO_1149 (O_1149,N_14989,N_14919);
and UO_1150 (O_1150,N_14921,N_14938);
nor UO_1151 (O_1151,N_14805,N_14842);
and UO_1152 (O_1152,N_14939,N_14935);
nand UO_1153 (O_1153,N_14983,N_14883);
nand UO_1154 (O_1154,N_14897,N_14945);
nand UO_1155 (O_1155,N_14935,N_14920);
nor UO_1156 (O_1156,N_14944,N_14952);
nand UO_1157 (O_1157,N_14840,N_14909);
nand UO_1158 (O_1158,N_14846,N_14874);
nor UO_1159 (O_1159,N_14974,N_14831);
nand UO_1160 (O_1160,N_14884,N_14842);
and UO_1161 (O_1161,N_14933,N_14880);
nand UO_1162 (O_1162,N_14877,N_14879);
nand UO_1163 (O_1163,N_14933,N_14956);
nor UO_1164 (O_1164,N_14828,N_14949);
nand UO_1165 (O_1165,N_14980,N_14804);
and UO_1166 (O_1166,N_14873,N_14832);
nand UO_1167 (O_1167,N_14879,N_14858);
and UO_1168 (O_1168,N_14973,N_14849);
and UO_1169 (O_1169,N_14826,N_14942);
and UO_1170 (O_1170,N_14834,N_14877);
and UO_1171 (O_1171,N_14991,N_14983);
nor UO_1172 (O_1172,N_14882,N_14801);
nand UO_1173 (O_1173,N_14820,N_14948);
and UO_1174 (O_1174,N_14922,N_14856);
or UO_1175 (O_1175,N_14831,N_14908);
and UO_1176 (O_1176,N_14996,N_14815);
xor UO_1177 (O_1177,N_14905,N_14930);
or UO_1178 (O_1178,N_14814,N_14885);
and UO_1179 (O_1179,N_14925,N_14863);
nand UO_1180 (O_1180,N_14968,N_14939);
and UO_1181 (O_1181,N_14836,N_14907);
xnor UO_1182 (O_1182,N_14849,N_14907);
or UO_1183 (O_1183,N_14817,N_14816);
or UO_1184 (O_1184,N_14921,N_14809);
and UO_1185 (O_1185,N_14944,N_14822);
xor UO_1186 (O_1186,N_14933,N_14959);
nand UO_1187 (O_1187,N_14979,N_14945);
or UO_1188 (O_1188,N_14903,N_14906);
nor UO_1189 (O_1189,N_14927,N_14851);
xnor UO_1190 (O_1190,N_14957,N_14985);
xnor UO_1191 (O_1191,N_14836,N_14946);
and UO_1192 (O_1192,N_14823,N_14831);
and UO_1193 (O_1193,N_14978,N_14898);
nand UO_1194 (O_1194,N_14821,N_14907);
nand UO_1195 (O_1195,N_14915,N_14802);
and UO_1196 (O_1196,N_14856,N_14923);
and UO_1197 (O_1197,N_14884,N_14946);
and UO_1198 (O_1198,N_14966,N_14843);
nand UO_1199 (O_1199,N_14967,N_14963);
nor UO_1200 (O_1200,N_14947,N_14925);
nand UO_1201 (O_1201,N_14996,N_14831);
and UO_1202 (O_1202,N_14999,N_14975);
and UO_1203 (O_1203,N_14815,N_14948);
nor UO_1204 (O_1204,N_14890,N_14914);
or UO_1205 (O_1205,N_14959,N_14859);
nand UO_1206 (O_1206,N_14985,N_14876);
nor UO_1207 (O_1207,N_14969,N_14828);
or UO_1208 (O_1208,N_14985,N_14884);
nor UO_1209 (O_1209,N_14849,N_14823);
or UO_1210 (O_1210,N_14947,N_14825);
and UO_1211 (O_1211,N_14934,N_14944);
or UO_1212 (O_1212,N_14928,N_14891);
nand UO_1213 (O_1213,N_14953,N_14861);
xnor UO_1214 (O_1214,N_14955,N_14899);
nand UO_1215 (O_1215,N_14915,N_14965);
nor UO_1216 (O_1216,N_14855,N_14871);
and UO_1217 (O_1217,N_14939,N_14936);
nand UO_1218 (O_1218,N_14963,N_14802);
nor UO_1219 (O_1219,N_14827,N_14873);
or UO_1220 (O_1220,N_14926,N_14946);
or UO_1221 (O_1221,N_14825,N_14950);
nor UO_1222 (O_1222,N_14985,N_14821);
nand UO_1223 (O_1223,N_14849,N_14963);
nand UO_1224 (O_1224,N_14975,N_14987);
nand UO_1225 (O_1225,N_14963,N_14809);
or UO_1226 (O_1226,N_14903,N_14822);
nand UO_1227 (O_1227,N_14986,N_14938);
or UO_1228 (O_1228,N_14982,N_14923);
nor UO_1229 (O_1229,N_14980,N_14883);
and UO_1230 (O_1230,N_14954,N_14801);
xnor UO_1231 (O_1231,N_14896,N_14900);
and UO_1232 (O_1232,N_14915,N_14844);
nor UO_1233 (O_1233,N_14959,N_14953);
xor UO_1234 (O_1234,N_14823,N_14971);
and UO_1235 (O_1235,N_14892,N_14971);
xnor UO_1236 (O_1236,N_14943,N_14848);
nand UO_1237 (O_1237,N_14824,N_14884);
or UO_1238 (O_1238,N_14824,N_14825);
nand UO_1239 (O_1239,N_14862,N_14824);
and UO_1240 (O_1240,N_14983,N_14829);
nor UO_1241 (O_1241,N_14897,N_14824);
nor UO_1242 (O_1242,N_14844,N_14960);
nand UO_1243 (O_1243,N_14945,N_14893);
nand UO_1244 (O_1244,N_14983,N_14914);
xnor UO_1245 (O_1245,N_14818,N_14875);
or UO_1246 (O_1246,N_14898,N_14803);
nand UO_1247 (O_1247,N_14829,N_14941);
and UO_1248 (O_1248,N_14939,N_14907);
nor UO_1249 (O_1249,N_14981,N_14912);
or UO_1250 (O_1250,N_14996,N_14859);
or UO_1251 (O_1251,N_14925,N_14810);
nor UO_1252 (O_1252,N_14869,N_14963);
or UO_1253 (O_1253,N_14960,N_14882);
or UO_1254 (O_1254,N_14938,N_14805);
nand UO_1255 (O_1255,N_14802,N_14953);
nand UO_1256 (O_1256,N_14819,N_14994);
nor UO_1257 (O_1257,N_14893,N_14854);
or UO_1258 (O_1258,N_14919,N_14867);
nor UO_1259 (O_1259,N_14828,N_14929);
nand UO_1260 (O_1260,N_14863,N_14967);
or UO_1261 (O_1261,N_14911,N_14950);
and UO_1262 (O_1262,N_14850,N_14922);
nand UO_1263 (O_1263,N_14988,N_14972);
nor UO_1264 (O_1264,N_14917,N_14964);
nor UO_1265 (O_1265,N_14985,N_14896);
and UO_1266 (O_1266,N_14940,N_14843);
nand UO_1267 (O_1267,N_14807,N_14974);
or UO_1268 (O_1268,N_14815,N_14924);
or UO_1269 (O_1269,N_14806,N_14875);
and UO_1270 (O_1270,N_14881,N_14922);
nand UO_1271 (O_1271,N_14919,N_14880);
or UO_1272 (O_1272,N_14835,N_14995);
xor UO_1273 (O_1273,N_14800,N_14901);
xnor UO_1274 (O_1274,N_14817,N_14970);
and UO_1275 (O_1275,N_14841,N_14996);
and UO_1276 (O_1276,N_14843,N_14901);
and UO_1277 (O_1277,N_14919,N_14862);
and UO_1278 (O_1278,N_14822,N_14952);
and UO_1279 (O_1279,N_14816,N_14805);
nand UO_1280 (O_1280,N_14951,N_14864);
nor UO_1281 (O_1281,N_14857,N_14998);
and UO_1282 (O_1282,N_14814,N_14840);
xnor UO_1283 (O_1283,N_14887,N_14930);
and UO_1284 (O_1284,N_14995,N_14986);
nor UO_1285 (O_1285,N_14914,N_14814);
and UO_1286 (O_1286,N_14831,N_14930);
and UO_1287 (O_1287,N_14929,N_14887);
nand UO_1288 (O_1288,N_14815,N_14972);
or UO_1289 (O_1289,N_14866,N_14877);
and UO_1290 (O_1290,N_14912,N_14959);
xnor UO_1291 (O_1291,N_14952,N_14976);
and UO_1292 (O_1292,N_14815,N_14964);
nand UO_1293 (O_1293,N_14969,N_14880);
and UO_1294 (O_1294,N_14873,N_14944);
and UO_1295 (O_1295,N_14862,N_14851);
nand UO_1296 (O_1296,N_14991,N_14972);
nor UO_1297 (O_1297,N_14919,N_14938);
nor UO_1298 (O_1298,N_14805,N_14927);
nor UO_1299 (O_1299,N_14948,N_14946);
nor UO_1300 (O_1300,N_14952,N_14826);
xnor UO_1301 (O_1301,N_14839,N_14953);
and UO_1302 (O_1302,N_14810,N_14981);
xor UO_1303 (O_1303,N_14931,N_14969);
or UO_1304 (O_1304,N_14811,N_14860);
nand UO_1305 (O_1305,N_14912,N_14927);
nand UO_1306 (O_1306,N_14951,N_14808);
or UO_1307 (O_1307,N_14806,N_14933);
nor UO_1308 (O_1308,N_14972,N_14829);
nor UO_1309 (O_1309,N_14844,N_14907);
or UO_1310 (O_1310,N_14894,N_14817);
and UO_1311 (O_1311,N_14890,N_14823);
or UO_1312 (O_1312,N_14835,N_14877);
or UO_1313 (O_1313,N_14850,N_14816);
or UO_1314 (O_1314,N_14920,N_14869);
nand UO_1315 (O_1315,N_14841,N_14883);
nand UO_1316 (O_1316,N_14925,N_14966);
nand UO_1317 (O_1317,N_14932,N_14921);
and UO_1318 (O_1318,N_14927,N_14884);
nor UO_1319 (O_1319,N_14973,N_14960);
nand UO_1320 (O_1320,N_14997,N_14883);
and UO_1321 (O_1321,N_14857,N_14993);
nor UO_1322 (O_1322,N_14949,N_14994);
or UO_1323 (O_1323,N_14925,N_14908);
nand UO_1324 (O_1324,N_14857,N_14836);
nand UO_1325 (O_1325,N_14840,N_14907);
nor UO_1326 (O_1326,N_14840,N_14805);
nor UO_1327 (O_1327,N_14969,N_14954);
xor UO_1328 (O_1328,N_14924,N_14933);
or UO_1329 (O_1329,N_14962,N_14988);
nand UO_1330 (O_1330,N_14860,N_14957);
nand UO_1331 (O_1331,N_14828,N_14874);
or UO_1332 (O_1332,N_14944,N_14861);
or UO_1333 (O_1333,N_14989,N_14978);
nor UO_1334 (O_1334,N_14869,N_14893);
nor UO_1335 (O_1335,N_14866,N_14886);
or UO_1336 (O_1336,N_14972,N_14873);
xnor UO_1337 (O_1337,N_14802,N_14944);
nor UO_1338 (O_1338,N_14869,N_14814);
or UO_1339 (O_1339,N_14885,N_14887);
or UO_1340 (O_1340,N_14870,N_14994);
or UO_1341 (O_1341,N_14947,N_14949);
nor UO_1342 (O_1342,N_14858,N_14819);
or UO_1343 (O_1343,N_14897,N_14891);
and UO_1344 (O_1344,N_14995,N_14875);
nand UO_1345 (O_1345,N_14960,N_14863);
nand UO_1346 (O_1346,N_14979,N_14916);
or UO_1347 (O_1347,N_14857,N_14971);
nand UO_1348 (O_1348,N_14948,N_14922);
or UO_1349 (O_1349,N_14857,N_14901);
nor UO_1350 (O_1350,N_14855,N_14861);
and UO_1351 (O_1351,N_14906,N_14842);
nor UO_1352 (O_1352,N_14930,N_14894);
and UO_1353 (O_1353,N_14897,N_14832);
nor UO_1354 (O_1354,N_14802,N_14862);
or UO_1355 (O_1355,N_14854,N_14848);
nor UO_1356 (O_1356,N_14969,N_14806);
xnor UO_1357 (O_1357,N_14978,N_14844);
nand UO_1358 (O_1358,N_14951,N_14829);
and UO_1359 (O_1359,N_14910,N_14876);
or UO_1360 (O_1360,N_14890,N_14967);
nand UO_1361 (O_1361,N_14900,N_14840);
nand UO_1362 (O_1362,N_14830,N_14943);
nor UO_1363 (O_1363,N_14999,N_14875);
and UO_1364 (O_1364,N_14819,N_14856);
nand UO_1365 (O_1365,N_14935,N_14954);
and UO_1366 (O_1366,N_14945,N_14959);
nor UO_1367 (O_1367,N_14898,N_14836);
and UO_1368 (O_1368,N_14845,N_14863);
nand UO_1369 (O_1369,N_14839,N_14977);
or UO_1370 (O_1370,N_14859,N_14865);
and UO_1371 (O_1371,N_14829,N_14814);
nand UO_1372 (O_1372,N_14809,N_14944);
nor UO_1373 (O_1373,N_14961,N_14903);
or UO_1374 (O_1374,N_14972,N_14872);
nor UO_1375 (O_1375,N_14899,N_14800);
and UO_1376 (O_1376,N_14864,N_14910);
nor UO_1377 (O_1377,N_14963,N_14887);
nor UO_1378 (O_1378,N_14812,N_14895);
nand UO_1379 (O_1379,N_14869,N_14841);
and UO_1380 (O_1380,N_14888,N_14949);
and UO_1381 (O_1381,N_14904,N_14847);
nand UO_1382 (O_1382,N_14886,N_14895);
or UO_1383 (O_1383,N_14812,N_14926);
nor UO_1384 (O_1384,N_14995,N_14920);
or UO_1385 (O_1385,N_14853,N_14805);
or UO_1386 (O_1386,N_14944,N_14915);
and UO_1387 (O_1387,N_14927,N_14901);
or UO_1388 (O_1388,N_14953,N_14847);
nand UO_1389 (O_1389,N_14989,N_14967);
or UO_1390 (O_1390,N_14907,N_14975);
and UO_1391 (O_1391,N_14886,N_14986);
xnor UO_1392 (O_1392,N_14961,N_14953);
nor UO_1393 (O_1393,N_14977,N_14851);
nor UO_1394 (O_1394,N_14865,N_14914);
nor UO_1395 (O_1395,N_14894,N_14836);
xor UO_1396 (O_1396,N_14811,N_14808);
nand UO_1397 (O_1397,N_14897,N_14997);
or UO_1398 (O_1398,N_14803,N_14914);
nand UO_1399 (O_1399,N_14873,N_14920);
nand UO_1400 (O_1400,N_14961,N_14992);
xnor UO_1401 (O_1401,N_14923,N_14869);
nand UO_1402 (O_1402,N_14921,N_14906);
and UO_1403 (O_1403,N_14971,N_14986);
nand UO_1404 (O_1404,N_14803,N_14990);
or UO_1405 (O_1405,N_14932,N_14944);
nand UO_1406 (O_1406,N_14970,N_14908);
nor UO_1407 (O_1407,N_14982,N_14943);
or UO_1408 (O_1408,N_14929,N_14981);
nor UO_1409 (O_1409,N_14818,N_14885);
xnor UO_1410 (O_1410,N_14846,N_14977);
or UO_1411 (O_1411,N_14823,N_14824);
nor UO_1412 (O_1412,N_14861,N_14895);
or UO_1413 (O_1413,N_14990,N_14852);
nor UO_1414 (O_1414,N_14993,N_14924);
xnor UO_1415 (O_1415,N_14839,N_14898);
or UO_1416 (O_1416,N_14892,N_14900);
nand UO_1417 (O_1417,N_14889,N_14951);
nand UO_1418 (O_1418,N_14929,N_14976);
nor UO_1419 (O_1419,N_14876,N_14973);
nand UO_1420 (O_1420,N_14907,N_14861);
nand UO_1421 (O_1421,N_14883,N_14843);
nor UO_1422 (O_1422,N_14999,N_14960);
or UO_1423 (O_1423,N_14923,N_14823);
nor UO_1424 (O_1424,N_14852,N_14870);
and UO_1425 (O_1425,N_14896,N_14975);
or UO_1426 (O_1426,N_14900,N_14998);
nor UO_1427 (O_1427,N_14961,N_14958);
or UO_1428 (O_1428,N_14828,N_14923);
or UO_1429 (O_1429,N_14880,N_14920);
nand UO_1430 (O_1430,N_14888,N_14857);
and UO_1431 (O_1431,N_14974,N_14934);
nor UO_1432 (O_1432,N_14816,N_14818);
or UO_1433 (O_1433,N_14935,N_14968);
nor UO_1434 (O_1434,N_14960,N_14801);
nand UO_1435 (O_1435,N_14964,N_14890);
nand UO_1436 (O_1436,N_14902,N_14997);
nor UO_1437 (O_1437,N_14971,N_14918);
and UO_1438 (O_1438,N_14962,N_14976);
or UO_1439 (O_1439,N_14867,N_14811);
nand UO_1440 (O_1440,N_14826,N_14913);
xor UO_1441 (O_1441,N_14811,N_14983);
xnor UO_1442 (O_1442,N_14810,N_14854);
nand UO_1443 (O_1443,N_14984,N_14850);
nor UO_1444 (O_1444,N_14812,N_14920);
nor UO_1445 (O_1445,N_14971,N_14987);
or UO_1446 (O_1446,N_14872,N_14860);
nor UO_1447 (O_1447,N_14880,N_14972);
nor UO_1448 (O_1448,N_14822,N_14973);
nand UO_1449 (O_1449,N_14991,N_14884);
and UO_1450 (O_1450,N_14884,N_14953);
or UO_1451 (O_1451,N_14974,N_14858);
xnor UO_1452 (O_1452,N_14862,N_14904);
nand UO_1453 (O_1453,N_14967,N_14920);
nor UO_1454 (O_1454,N_14927,N_14990);
nand UO_1455 (O_1455,N_14833,N_14939);
nor UO_1456 (O_1456,N_14871,N_14974);
nor UO_1457 (O_1457,N_14957,N_14972);
and UO_1458 (O_1458,N_14987,N_14924);
nand UO_1459 (O_1459,N_14853,N_14929);
nand UO_1460 (O_1460,N_14969,N_14991);
nor UO_1461 (O_1461,N_14947,N_14810);
nor UO_1462 (O_1462,N_14850,N_14912);
nor UO_1463 (O_1463,N_14868,N_14943);
nand UO_1464 (O_1464,N_14857,N_14833);
nor UO_1465 (O_1465,N_14964,N_14880);
and UO_1466 (O_1466,N_14854,N_14864);
xor UO_1467 (O_1467,N_14902,N_14851);
nand UO_1468 (O_1468,N_14939,N_14810);
xnor UO_1469 (O_1469,N_14868,N_14897);
or UO_1470 (O_1470,N_14940,N_14975);
nand UO_1471 (O_1471,N_14873,N_14939);
nand UO_1472 (O_1472,N_14878,N_14898);
and UO_1473 (O_1473,N_14858,N_14984);
xnor UO_1474 (O_1474,N_14878,N_14931);
and UO_1475 (O_1475,N_14945,N_14954);
and UO_1476 (O_1476,N_14848,N_14853);
nand UO_1477 (O_1477,N_14939,N_14858);
or UO_1478 (O_1478,N_14939,N_14866);
and UO_1479 (O_1479,N_14885,N_14914);
nand UO_1480 (O_1480,N_14870,N_14921);
xor UO_1481 (O_1481,N_14868,N_14804);
nand UO_1482 (O_1482,N_14892,N_14944);
xnor UO_1483 (O_1483,N_14851,N_14842);
nand UO_1484 (O_1484,N_14858,N_14842);
nand UO_1485 (O_1485,N_14956,N_14993);
and UO_1486 (O_1486,N_14954,N_14919);
nor UO_1487 (O_1487,N_14807,N_14977);
nor UO_1488 (O_1488,N_14983,N_14820);
nand UO_1489 (O_1489,N_14912,N_14820);
and UO_1490 (O_1490,N_14930,N_14889);
and UO_1491 (O_1491,N_14948,N_14962);
or UO_1492 (O_1492,N_14836,N_14805);
nor UO_1493 (O_1493,N_14809,N_14871);
or UO_1494 (O_1494,N_14883,N_14924);
xnor UO_1495 (O_1495,N_14899,N_14814);
nand UO_1496 (O_1496,N_14882,N_14920);
nor UO_1497 (O_1497,N_14995,N_14984);
and UO_1498 (O_1498,N_14926,N_14820);
nand UO_1499 (O_1499,N_14895,N_14972);
xor UO_1500 (O_1500,N_14808,N_14995);
or UO_1501 (O_1501,N_14987,N_14947);
or UO_1502 (O_1502,N_14866,N_14869);
or UO_1503 (O_1503,N_14926,N_14834);
nor UO_1504 (O_1504,N_14818,N_14958);
nor UO_1505 (O_1505,N_14911,N_14986);
nor UO_1506 (O_1506,N_14891,N_14906);
and UO_1507 (O_1507,N_14984,N_14986);
or UO_1508 (O_1508,N_14826,N_14864);
and UO_1509 (O_1509,N_14824,N_14956);
xnor UO_1510 (O_1510,N_14988,N_14838);
nand UO_1511 (O_1511,N_14917,N_14900);
and UO_1512 (O_1512,N_14901,N_14871);
nor UO_1513 (O_1513,N_14892,N_14946);
nand UO_1514 (O_1514,N_14873,N_14858);
xor UO_1515 (O_1515,N_14918,N_14801);
and UO_1516 (O_1516,N_14801,N_14809);
or UO_1517 (O_1517,N_14896,N_14811);
nor UO_1518 (O_1518,N_14907,N_14977);
nor UO_1519 (O_1519,N_14836,N_14941);
xnor UO_1520 (O_1520,N_14930,N_14810);
or UO_1521 (O_1521,N_14891,N_14822);
xnor UO_1522 (O_1522,N_14855,N_14816);
or UO_1523 (O_1523,N_14872,N_14962);
nor UO_1524 (O_1524,N_14915,N_14830);
and UO_1525 (O_1525,N_14816,N_14892);
xor UO_1526 (O_1526,N_14968,N_14998);
or UO_1527 (O_1527,N_14895,N_14990);
nor UO_1528 (O_1528,N_14898,N_14862);
or UO_1529 (O_1529,N_14955,N_14811);
nand UO_1530 (O_1530,N_14834,N_14944);
or UO_1531 (O_1531,N_14908,N_14896);
nand UO_1532 (O_1532,N_14847,N_14924);
and UO_1533 (O_1533,N_14980,N_14898);
nor UO_1534 (O_1534,N_14920,N_14803);
nand UO_1535 (O_1535,N_14908,N_14900);
nor UO_1536 (O_1536,N_14915,N_14933);
and UO_1537 (O_1537,N_14873,N_14845);
and UO_1538 (O_1538,N_14936,N_14976);
or UO_1539 (O_1539,N_14843,N_14939);
xor UO_1540 (O_1540,N_14988,N_14853);
and UO_1541 (O_1541,N_14973,N_14820);
and UO_1542 (O_1542,N_14941,N_14827);
and UO_1543 (O_1543,N_14812,N_14870);
nand UO_1544 (O_1544,N_14871,N_14950);
nand UO_1545 (O_1545,N_14960,N_14864);
or UO_1546 (O_1546,N_14871,N_14854);
xnor UO_1547 (O_1547,N_14951,N_14913);
nor UO_1548 (O_1548,N_14990,N_14887);
or UO_1549 (O_1549,N_14983,N_14939);
nor UO_1550 (O_1550,N_14883,N_14941);
nor UO_1551 (O_1551,N_14894,N_14880);
or UO_1552 (O_1552,N_14932,N_14943);
nor UO_1553 (O_1553,N_14927,N_14974);
and UO_1554 (O_1554,N_14839,N_14997);
or UO_1555 (O_1555,N_14859,N_14834);
xnor UO_1556 (O_1556,N_14866,N_14820);
or UO_1557 (O_1557,N_14810,N_14885);
and UO_1558 (O_1558,N_14926,N_14830);
nor UO_1559 (O_1559,N_14932,N_14830);
or UO_1560 (O_1560,N_14820,N_14976);
and UO_1561 (O_1561,N_14825,N_14902);
nand UO_1562 (O_1562,N_14933,N_14919);
nand UO_1563 (O_1563,N_14929,N_14934);
and UO_1564 (O_1564,N_14811,N_14941);
nor UO_1565 (O_1565,N_14809,N_14872);
nand UO_1566 (O_1566,N_14866,N_14816);
nor UO_1567 (O_1567,N_14991,N_14846);
and UO_1568 (O_1568,N_14801,N_14881);
and UO_1569 (O_1569,N_14839,N_14937);
nor UO_1570 (O_1570,N_14848,N_14824);
or UO_1571 (O_1571,N_14831,N_14882);
or UO_1572 (O_1572,N_14829,N_14853);
and UO_1573 (O_1573,N_14895,N_14983);
nor UO_1574 (O_1574,N_14891,N_14802);
nor UO_1575 (O_1575,N_14882,N_14864);
and UO_1576 (O_1576,N_14945,N_14928);
nor UO_1577 (O_1577,N_14911,N_14989);
nand UO_1578 (O_1578,N_14947,N_14997);
nand UO_1579 (O_1579,N_14978,N_14804);
nor UO_1580 (O_1580,N_14974,N_14902);
nor UO_1581 (O_1581,N_14982,N_14895);
or UO_1582 (O_1582,N_14881,N_14856);
or UO_1583 (O_1583,N_14836,N_14979);
xor UO_1584 (O_1584,N_14952,N_14802);
or UO_1585 (O_1585,N_14887,N_14880);
or UO_1586 (O_1586,N_14805,N_14879);
nand UO_1587 (O_1587,N_14823,N_14984);
nor UO_1588 (O_1588,N_14824,N_14892);
nor UO_1589 (O_1589,N_14835,N_14975);
nand UO_1590 (O_1590,N_14885,N_14963);
or UO_1591 (O_1591,N_14863,N_14893);
and UO_1592 (O_1592,N_14898,N_14968);
and UO_1593 (O_1593,N_14860,N_14918);
nor UO_1594 (O_1594,N_14944,N_14942);
nor UO_1595 (O_1595,N_14930,N_14809);
nor UO_1596 (O_1596,N_14995,N_14907);
nor UO_1597 (O_1597,N_14933,N_14906);
xnor UO_1598 (O_1598,N_14922,N_14969);
or UO_1599 (O_1599,N_14981,N_14956);
or UO_1600 (O_1600,N_14940,N_14892);
nand UO_1601 (O_1601,N_14915,N_14973);
and UO_1602 (O_1602,N_14926,N_14898);
or UO_1603 (O_1603,N_14928,N_14851);
nor UO_1604 (O_1604,N_14839,N_14847);
nor UO_1605 (O_1605,N_14832,N_14938);
nor UO_1606 (O_1606,N_14928,N_14875);
xor UO_1607 (O_1607,N_14915,N_14959);
and UO_1608 (O_1608,N_14873,N_14957);
nor UO_1609 (O_1609,N_14911,N_14867);
and UO_1610 (O_1610,N_14882,N_14979);
nand UO_1611 (O_1611,N_14852,N_14937);
nand UO_1612 (O_1612,N_14912,N_14907);
nand UO_1613 (O_1613,N_14933,N_14891);
and UO_1614 (O_1614,N_14934,N_14922);
xor UO_1615 (O_1615,N_14889,N_14963);
nand UO_1616 (O_1616,N_14874,N_14882);
or UO_1617 (O_1617,N_14947,N_14822);
xor UO_1618 (O_1618,N_14821,N_14977);
nand UO_1619 (O_1619,N_14955,N_14980);
and UO_1620 (O_1620,N_14987,N_14804);
nand UO_1621 (O_1621,N_14870,N_14950);
nor UO_1622 (O_1622,N_14995,N_14989);
or UO_1623 (O_1623,N_14900,N_14946);
nand UO_1624 (O_1624,N_14913,N_14901);
and UO_1625 (O_1625,N_14898,N_14813);
or UO_1626 (O_1626,N_14830,N_14821);
or UO_1627 (O_1627,N_14956,N_14971);
nor UO_1628 (O_1628,N_14905,N_14945);
nand UO_1629 (O_1629,N_14871,N_14972);
and UO_1630 (O_1630,N_14974,N_14992);
nor UO_1631 (O_1631,N_14847,N_14909);
xor UO_1632 (O_1632,N_14868,N_14957);
or UO_1633 (O_1633,N_14888,N_14863);
and UO_1634 (O_1634,N_14908,N_14864);
or UO_1635 (O_1635,N_14903,N_14932);
and UO_1636 (O_1636,N_14942,N_14864);
and UO_1637 (O_1637,N_14830,N_14997);
or UO_1638 (O_1638,N_14812,N_14977);
or UO_1639 (O_1639,N_14871,N_14983);
nor UO_1640 (O_1640,N_14993,N_14941);
nand UO_1641 (O_1641,N_14828,N_14970);
and UO_1642 (O_1642,N_14923,N_14950);
and UO_1643 (O_1643,N_14803,N_14861);
or UO_1644 (O_1644,N_14961,N_14806);
or UO_1645 (O_1645,N_14850,N_14998);
and UO_1646 (O_1646,N_14831,N_14820);
or UO_1647 (O_1647,N_14990,N_14935);
and UO_1648 (O_1648,N_14840,N_14958);
and UO_1649 (O_1649,N_14871,N_14804);
nand UO_1650 (O_1650,N_14934,N_14946);
nor UO_1651 (O_1651,N_14919,N_14972);
and UO_1652 (O_1652,N_14818,N_14992);
and UO_1653 (O_1653,N_14975,N_14995);
nand UO_1654 (O_1654,N_14885,N_14892);
nor UO_1655 (O_1655,N_14897,N_14885);
xor UO_1656 (O_1656,N_14867,N_14897);
nand UO_1657 (O_1657,N_14926,N_14810);
nor UO_1658 (O_1658,N_14881,N_14852);
nor UO_1659 (O_1659,N_14982,N_14968);
and UO_1660 (O_1660,N_14813,N_14891);
and UO_1661 (O_1661,N_14894,N_14891);
xor UO_1662 (O_1662,N_14886,N_14953);
or UO_1663 (O_1663,N_14830,N_14867);
or UO_1664 (O_1664,N_14875,N_14824);
xnor UO_1665 (O_1665,N_14828,N_14846);
xnor UO_1666 (O_1666,N_14803,N_14945);
nor UO_1667 (O_1667,N_14829,N_14838);
nor UO_1668 (O_1668,N_14819,N_14988);
nand UO_1669 (O_1669,N_14998,N_14892);
or UO_1670 (O_1670,N_14923,N_14994);
or UO_1671 (O_1671,N_14949,N_14948);
or UO_1672 (O_1672,N_14913,N_14992);
or UO_1673 (O_1673,N_14860,N_14997);
and UO_1674 (O_1674,N_14909,N_14885);
nand UO_1675 (O_1675,N_14913,N_14885);
xnor UO_1676 (O_1676,N_14910,N_14974);
nor UO_1677 (O_1677,N_14847,N_14850);
xor UO_1678 (O_1678,N_14829,N_14952);
nor UO_1679 (O_1679,N_14844,N_14970);
nor UO_1680 (O_1680,N_14925,N_14960);
nand UO_1681 (O_1681,N_14970,N_14973);
or UO_1682 (O_1682,N_14816,N_14845);
nand UO_1683 (O_1683,N_14970,N_14841);
or UO_1684 (O_1684,N_14905,N_14857);
and UO_1685 (O_1685,N_14984,N_14907);
nand UO_1686 (O_1686,N_14833,N_14927);
nor UO_1687 (O_1687,N_14994,N_14999);
and UO_1688 (O_1688,N_14924,N_14868);
and UO_1689 (O_1689,N_14950,N_14961);
nor UO_1690 (O_1690,N_14807,N_14957);
nor UO_1691 (O_1691,N_14936,N_14914);
and UO_1692 (O_1692,N_14956,N_14905);
or UO_1693 (O_1693,N_14807,N_14903);
nand UO_1694 (O_1694,N_14887,N_14924);
nor UO_1695 (O_1695,N_14993,N_14992);
nor UO_1696 (O_1696,N_14906,N_14847);
or UO_1697 (O_1697,N_14854,N_14850);
nor UO_1698 (O_1698,N_14862,N_14970);
or UO_1699 (O_1699,N_14965,N_14963);
nand UO_1700 (O_1700,N_14850,N_14825);
xnor UO_1701 (O_1701,N_14842,N_14992);
nor UO_1702 (O_1702,N_14881,N_14972);
and UO_1703 (O_1703,N_14990,N_14936);
and UO_1704 (O_1704,N_14825,N_14852);
or UO_1705 (O_1705,N_14846,N_14902);
and UO_1706 (O_1706,N_14879,N_14888);
nand UO_1707 (O_1707,N_14800,N_14887);
or UO_1708 (O_1708,N_14859,N_14914);
and UO_1709 (O_1709,N_14834,N_14863);
nand UO_1710 (O_1710,N_14952,N_14915);
and UO_1711 (O_1711,N_14834,N_14870);
nand UO_1712 (O_1712,N_14953,N_14974);
and UO_1713 (O_1713,N_14998,N_14813);
or UO_1714 (O_1714,N_14880,N_14844);
nand UO_1715 (O_1715,N_14821,N_14803);
or UO_1716 (O_1716,N_14998,N_14997);
and UO_1717 (O_1717,N_14964,N_14844);
and UO_1718 (O_1718,N_14885,N_14878);
and UO_1719 (O_1719,N_14961,N_14973);
nor UO_1720 (O_1720,N_14922,N_14865);
nand UO_1721 (O_1721,N_14944,N_14804);
nand UO_1722 (O_1722,N_14967,N_14931);
and UO_1723 (O_1723,N_14836,N_14915);
or UO_1724 (O_1724,N_14854,N_14822);
or UO_1725 (O_1725,N_14958,N_14809);
or UO_1726 (O_1726,N_14874,N_14817);
or UO_1727 (O_1727,N_14887,N_14939);
xnor UO_1728 (O_1728,N_14848,N_14977);
or UO_1729 (O_1729,N_14809,N_14806);
or UO_1730 (O_1730,N_14965,N_14858);
nor UO_1731 (O_1731,N_14972,N_14801);
nor UO_1732 (O_1732,N_14868,N_14893);
nor UO_1733 (O_1733,N_14802,N_14853);
or UO_1734 (O_1734,N_14957,N_14839);
and UO_1735 (O_1735,N_14933,N_14894);
nor UO_1736 (O_1736,N_14863,N_14832);
nand UO_1737 (O_1737,N_14811,N_14954);
and UO_1738 (O_1738,N_14840,N_14954);
nor UO_1739 (O_1739,N_14966,N_14913);
nand UO_1740 (O_1740,N_14898,N_14938);
nor UO_1741 (O_1741,N_14845,N_14828);
or UO_1742 (O_1742,N_14962,N_14806);
and UO_1743 (O_1743,N_14873,N_14917);
nand UO_1744 (O_1744,N_14897,N_14855);
and UO_1745 (O_1745,N_14936,N_14981);
nand UO_1746 (O_1746,N_14900,N_14914);
and UO_1747 (O_1747,N_14905,N_14898);
and UO_1748 (O_1748,N_14879,N_14868);
and UO_1749 (O_1749,N_14904,N_14894);
or UO_1750 (O_1750,N_14832,N_14961);
nand UO_1751 (O_1751,N_14963,N_14999);
and UO_1752 (O_1752,N_14875,N_14834);
and UO_1753 (O_1753,N_14945,N_14953);
nand UO_1754 (O_1754,N_14979,N_14856);
nand UO_1755 (O_1755,N_14844,N_14903);
or UO_1756 (O_1756,N_14922,N_14888);
and UO_1757 (O_1757,N_14954,N_14879);
or UO_1758 (O_1758,N_14900,N_14886);
nor UO_1759 (O_1759,N_14956,N_14863);
nand UO_1760 (O_1760,N_14820,N_14965);
and UO_1761 (O_1761,N_14815,N_14962);
or UO_1762 (O_1762,N_14985,N_14816);
nand UO_1763 (O_1763,N_14902,N_14958);
and UO_1764 (O_1764,N_14811,N_14987);
and UO_1765 (O_1765,N_14837,N_14962);
nand UO_1766 (O_1766,N_14919,N_14966);
or UO_1767 (O_1767,N_14816,N_14912);
or UO_1768 (O_1768,N_14952,N_14849);
or UO_1769 (O_1769,N_14907,N_14877);
nor UO_1770 (O_1770,N_14970,N_14815);
and UO_1771 (O_1771,N_14824,N_14954);
nand UO_1772 (O_1772,N_14893,N_14873);
and UO_1773 (O_1773,N_14920,N_14999);
nor UO_1774 (O_1774,N_14998,N_14977);
xnor UO_1775 (O_1775,N_14879,N_14943);
or UO_1776 (O_1776,N_14912,N_14906);
and UO_1777 (O_1777,N_14993,N_14936);
nand UO_1778 (O_1778,N_14964,N_14966);
nor UO_1779 (O_1779,N_14949,N_14809);
nor UO_1780 (O_1780,N_14939,N_14946);
nand UO_1781 (O_1781,N_14877,N_14998);
nor UO_1782 (O_1782,N_14975,N_14847);
and UO_1783 (O_1783,N_14901,N_14846);
xnor UO_1784 (O_1784,N_14800,N_14944);
nor UO_1785 (O_1785,N_14880,N_14805);
nand UO_1786 (O_1786,N_14806,N_14973);
nor UO_1787 (O_1787,N_14931,N_14914);
nand UO_1788 (O_1788,N_14804,N_14933);
xor UO_1789 (O_1789,N_14931,N_14948);
nand UO_1790 (O_1790,N_14858,N_14999);
xor UO_1791 (O_1791,N_14977,N_14860);
nor UO_1792 (O_1792,N_14971,N_14820);
xnor UO_1793 (O_1793,N_14899,N_14952);
and UO_1794 (O_1794,N_14943,N_14959);
or UO_1795 (O_1795,N_14975,N_14812);
nor UO_1796 (O_1796,N_14812,N_14963);
nor UO_1797 (O_1797,N_14910,N_14896);
and UO_1798 (O_1798,N_14978,N_14827);
and UO_1799 (O_1799,N_14950,N_14835);
or UO_1800 (O_1800,N_14982,N_14973);
nor UO_1801 (O_1801,N_14838,N_14821);
and UO_1802 (O_1802,N_14916,N_14808);
xnor UO_1803 (O_1803,N_14826,N_14982);
or UO_1804 (O_1804,N_14820,N_14886);
nand UO_1805 (O_1805,N_14960,N_14892);
or UO_1806 (O_1806,N_14825,N_14991);
or UO_1807 (O_1807,N_14968,N_14948);
nor UO_1808 (O_1808,N_14950,N_14861);
xnor UO_1809 (O_1809,N_14843,N_14896);
nor UO_1810 (O_1810,N_14906,N_14974);
nand UO_1811 (O_1811,N_14963,N_14888);
or UO_1812 (O_1812,N_14913,N_14833);
and UO_1813 (O_1813,N_14828,N_14850);
and UO_1814 (O_1814,N_14954,N_14883);
nand UO_1815 (O_1815,N_14859,N_14805);
xor UO_1816 (O_1816,N_14986,N_14806);
nor UO_1817 (O_1817,N_14809,N_14867);
nor UO_1818 (O_1818,N_14810,N_14858);
nand UO_1819 (O_1819,N_14966,N_14978);
nand UO_1820 (O_1820,N_14994,N_14935);
nand UO_1821 (O_1821,N_14980,N_14839);
or UO_1822 (O_1822,N_14898,N_14827);
nor UO_1823 (O_1823,N_14924,N_14929);
xor UO_1824 (O_1824,N_14828,N_14936);
xnor UO_1825 (O_1825,N_14937,N_14817);
xnor UO_1826 (O_1826,N_14936,N_14901);
and UO_1827 (O_1827,N_14988,N_14951);
nor UO_1828 (O_1828,N_14998,N_14882);
and UO_1829 (O_1829,N_14803,N_14974);
and UO_1830 (O_1830,N_14899,N_14947);
nand UO_1831 (O_1831,N_14839,N_14862);
nor UO_1832 (O_1832,N_14978,N_14942);
nor UO_1833 (O_1833,N_14801,N_14811);
xnor UO_1834 (O_1834,N_14800,N_14940);
and UO_1835 (O_1835,N_14842,N_14875);
nand UO_1836 (O_1836,N_14869,N_14959);
and UO_1837 (O_1837,N_14869,N_14933);
nor UO_1838 (O_1838,N_14870,N_14902);
nor UO_1839 (O_1839,N_14855,N_14977);
xnor UO_1840 (O_1840,N_14973,N_14962);
or UO_1841 (O_1841,N_14871,N_14814);
and UO_1842 (O_1842,N_14997,N_14821);
nand UO_1843 (O_1843,N_14804,N_14879);
nor UO_1844 (O_1844,N_14800,N_14984);
nand UO_1845 (O_1845,N_14834,N_14882);
and UO_1846 (O_1846,N_14834,N_14899);
and UO_1847 (O_1847,N_14934,N_14887);
and UO_1848 (O_1848,N_14902,N_14814);
nor UO_1849 (O_1849,N_14956,N_14812);
nand UO_1850 (O_1850,N_14963,N_14971);
nor UO_1851 (O_1851,N_14809,N_14986);
nand UO_1852 (O_1852,N_14977,N_14995);
or UO_1853 (O_1853,N_14824,N_14973);
and UO_1854 (O_1854,N_14878,N_14942);
or UO_1855 (O_1855,N_14941,N_14841);
xor UO_1856 (O_1856,N_14835,N_14843);
nand UO_1857 (O_1857,N_14835,N_14999);
nand UO_1858 (O_1858,N_14922,N_14849);
nor UO_1859 (O_1859,N_14897,N_14980);
or UO_1860 (O_1860,N_14826,N_14804);
and UO_1861 (O_1861,N_14823,N_14874);
xnor UO_1862 (O_1862,N_14883,N_14857);
nand UO_1863 (O_1863,N_14884,N_14899);
nor UO_1864 (O_1864,N_14840,N_14965);
nor UO_1865 (O_1865,N_14841,N_14912);
or UO_1866 (O_1866,N_14808,N_14802);
nor UO_1867 (O_1867,N_14837,N_14987);
or UO_1868 (O_1868,N_14921,N_14919);
nand UO_1869 (O_1869,N_14841,N_14998);
and UO_1870 (O_1870,N_14913,N_14967);
nand UO_1871 (O_1871,N_14987,N_14898);
xnor UO_1872 (O_1872,N_14876,N_14822);
or UO_1873 (O_1873,N_14898,N_14841);
nor UO_1874 (O_1874,N_14807,N_14836);
xnor UO_1875 (O_1875,N_14967,N_14975);
and UO_1876 (O_1876,N_14883,N_14831);
and UO_1877 (O_1877,N_14981,N_14952);
nand UO_1878 (O_1878,N_14908,N_14858);
nor UO_1879 (O_1879,N_14996,N_14938);
nor UO_1880 (O_1880,N_14905,N_14834);
xor UO_1881 (O_1881,N_14822,N_14861);
nor UO_1882 (O_1882,N_14983,N_14827);
or UO_1883 (O_1883,N_14917,N_14978);
or UO_1884 (O_1884,N_14956,N_14997);
or UO_1885 (O_1885,N_14838,N_14888);
nor UO_1886 (O_1886,N_14868,N_14823);
or UO_1887 (O_1887,N_14958,N_14924);
or UO_1888 (O_1888,N_14828,N_14981);
or UO_1889 (O_1889,N_14868,N_14802);
nand UO_1890 (O_1890,N_14885,N_14838);
and UO_1891 (O_1891,N_14916,N_14817);
or UO_1892 (O_1892,N_14908,N_14884);
or UO_1893 (O_1893,N_14872,N_14954);
and UO_1894 (O_1894,N_14907,N_14946);
nor UO_1895 (O_1895,N_14912,N_14976);
nor UO_1896 (O_1896,N_14820,N_14896);
or UO_1897 (O_1897,N_14810,N_14900);
or UO_1898 (O_1898,N_14992,N_14890);
nor UO_1899 (O_1899,N_14894,N_14819);
nand UO_1900 (O_1900,N_14838,N_14847);
nand UO_1901 (O_1901,N_14904,N_14842);
and UO_1902 (O_1902,N_14860,N_14830);
and UO_1903 (O_1903,N_14862,N_14863);
xor UO_1904 (O_1904,N_14841,N_14810);
and UO_1905 (O_1905,N_14976,N_14811);
nor UO_1906 (O_1906,N_14989,N_14819);
and UO_1907 (O_1907,N_14903,N_14975);
nand UO_1908 (O_1908,N_14958,N_14839);
nand UO_1909 (O_1909,N_14961,N_14869);
nor UO_1910 (O_1910,N_14917,N_14829);
or UO_1911 (O_1911,N_14833,N_14966);
nor UO_1912 (O_1912,N_14898,N_14824);
nor UO_1913 (O_1913,N_14992,N_14987);
or UO_1914 (O_1914,N_14803,N_14901);
and UO_1915 (O_1915,N_14801,N_14916);
nand UO_1916 (O_1916,N_14982,N_14862);
and UO_1917 (O_1917,N_14992,N_14865);
or UO_1918 (O_1918,N_14983,N_14865);
nand UO_1919 (O_1919,N_14977,N_14923);
or UO_1920 (O_1920,N_14954,N_14959);
nor UO_1921 (O_1921,N_14922,N_14823);
or UO_1922 (O_1922,N_14972,N_14924);
nor UO_1923 (O_1923,N_14894,N_14992);
or UO_1924 (O_1924,N_14841,N_14876);
xnor UO_1925 (O_1925,N_14996,N_14905);
or UO_1926 (O_1926,N_14849,N_14813);
nor UO_1927 (O_1927,N_14939,N_14956);
nor UO_1928 (O_1928,N_14999,N_14977);
nand UO_1929 (O_1929,N_14971,N_14813);
or UO_1930 (O_1930,N_14912,N_14992);
nand UO_1931 (O_1931,N_14877,N_14927);
nor UO_1932 (O_1932,N_14949,N_14969);
nand UO_1933 (O_1933,N_14842,N_14830);
nor UO_1934 (O_1934,N_14901,N_14865);
nor UO_1935 (O_1935,N_14851,N_14855);
and UO_1936 (O_1936,N_14956,N_14946);
xor UO_1937 (O_1937,N_14956,N_14887);
nor UO_1938 (O_1938,N_14975,N_14898);
nand UO_1939 (O_1939,N_14949,N_14897);
nor UO_1940 (O_1940,N_14969,N_14862);
and UO_1941 (O_1941,N_14981,N_14939);
or UO_1942 (O_1942,N_14980,N_14920);
xor UO_1943 (O_1943,N_14823,N_14980);
nor UO_1944 (O_1944,N_14897,N_14955);
and UO_1945 (O_1945,N_14934,N_14850);
nor UO_1946 (O_1946,N_14829,N_14836);
or UO_1947 (O_1947,N_14827,N_14830);
nand UO_1948 (O_1948,N_14912,N_14811);
and UO_1949 (O_1949,N_14985,N_14847);
xnor UO_1950 (O_1950,N_14936,N_14909);
nand UO_1951 (O_1951,N_14831,N_14865);
or UO_1952 (O_1952,N_14837,N_14986);
and UO_1953 (O_1953,N_14994,N_14931);
nand UO_1954 (O_1954,N_14851,N_14958);
xnor UO_1955 (O_1955,N_14983,N_14980);
nand UO_1956 (O_1956,N_14911,N_14803);
or UO_1957 (O_1957,N_14896,N_14952);
or UO_1958 (O_1958,N_14876,N_14839);
and UO_1959 (O_1959,N_14800,N_14880);
and UO_1960 (O_1960,N_14803,N_14955);
nor UO_1961 (O_1961,N_14974,N_14997);
and UO_1962 (O_1962,N_14966,N_14800);
and UO_1963 (O_1963,N_14926,N_14928);
nor UO_1964 (O_1964,N_14963,N_14858);
nor UO_1965 (O_1965,N_14917,N_14853);
or UO_1966 (O_1966,N_14981,N_14973);
xor UO_1967 (O_1967,N_14890,N_14878);
and UO_1968 (O_1968,N_14828,N_14977);
nand UO_1969 (O_1969,N_14879,N_14830);
xor UO_1970 (O_1970,N_14943,N_14958);
nand UO_1971 (O_1971,N_14840,N_14859);
or UO_1972 (O_1972,N_14821,N_14943);
nand UO_1973 (O_1973,N_14918,N_14885);
nand UO_1974 (O_1974,N_14900,N_14818);
nand UO_1975 (O_1975,N_14924,N_14856);
and UO_1976 (O_1976,N_14872,N_14856);
or UO_1977 (O_1977,N_14941,N_14918);
nor UO_1978 (O_1978,N_14933,N_14858);
or UO_1979 (O_1979,N_14962,N_14813);
nand UO_1980 (O_1980,N_14828,N_14932);
xor UO_1981 (O_1981,N_14863,N_14988);
nand UO_1982 (O_1982,N_14982,N_14808);
and UO_1983 (O_1983,N_14817,N_14849);
nor UO_1984 (O_1984,N_14805,N_14818);
nor UO_1985 (O_1985,N_14840,N_14828);
or UO_1986 (O_1986,N_14822,N_14955);
and UO_1987 (O_1987,N_14866,N_14864);
and UO_1988 (O_1988,N_14940,N_14931);
and UO_1989 (O_1989,N_14865,N_14834);
nor UO_1990 (O_1990,N_14845,N_14989);
and UO_1991 (O_1991,N_14901,N_14829);
and UO_1992 (O_1992,N_14882,N_14818);
nand UO_1993 (O_1993,N_14811,N_14803);
or UO_1994 (O_1994,N_14920,N_14922);
nand UO_1995 (O_1995,N_14923,N_14848);
nand UO_1996 (O_1996,N_14970,N_14837);
nor UO_1997 (O_1997,N_14831,N_14950);
and UO_1998 (O_1998,N_14842,N_14811);
nor UO_1999 (O_1999,N_14844,N_14984);
endmodule