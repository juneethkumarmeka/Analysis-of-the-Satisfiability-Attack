module basic_2500_25000_3000_5_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
and U0 (N_0,In_304,In_642);
nor U1 (N_1,In_1333,In_1325);
nor U2 (N_2,In_2412,In_2485);
nand U3 (N_3,In_2456,In_981);
or U4 (N_4,In_1535,In_1244);
xor U5 (N_5,In_1030,In_375);
and U6 (N_6,In_708,In_91);
nor U7 (N_7,In_436,In_1875);
nor U8 (N_8,In_136,In_747);
or U9 (N_9,In_2365,In_1582);
nor U10 (N_10,In_330,In_1874);
and U11 (N_11,In_1612,In_2154);
xor U12 (N_12,In_955,In_982);
nand U13 (N_13,In_201,In_346);
and U14 (N_14,In_1881,In_1024);
nor U15 (N_15,In_1630,In_2116);
nand U16 (N_16,In_1093,In_348);
or U17 (N_17,In_352,In_783);
xor U18 (N_18,In_1563,In_2137);
or U19 (N_19,In_1588,In_1367);
and U20 (N_20,In_2413,In_2119);
nand U21 (N_21,In_1692,In_1757);
xnor U22 (N_22,In_385,In_1720);
nor U23 (N_23,In_2249,In_1061);
xnor U24 (N_24,In_714,In_2173);
or U25 (N_25,In_769,In_261);
nor U26 (N_26,In_2449,In_415);
or U27 (N_27,In_478,In_1899);
or U28 (N_28,In_958,In_1355);
xor U29 (N_29,In_210,In_414);
or U30 (N_30,In_2262,In_442);
xnor U31 (N_31,In_876,In_485);
nand U32 (N_32,In_860,In_1837);
or U33 (N_33,In_1507,In_2024);
and U34 (N_34,In_251,In_1082);
nor U35 (N_35,In_1859,In_932);
and U36 (N_36,In_1790,In_1877);
and U37 (N_37,In_1980,In_426);
or U38 (N_38,In_2201,In_1112);
or U39 (N_39,In_417,In_2041);
and U40 (N_40,In_320,In_2356);
nand U41 (N_41,In_46,In_1710);
or U42 (N_42,In_897,In_649);
and U43 (N_43,In_337,In_1649);
and U44 (N_44,In_1767,In_940);
nor U45 (N_45,In_64,In_12);
nand U46 (N_46,In_2327,In_738);
nor U47 (N_47,In_779,In_1696);
nand U48 (N_48,In_1388,In_1516);
nor U49 (N_49,In_490,In_1044);
nor U50 (N_50,In_573,In_373);
xnor U51 (N_51,In_2372,In_281);
and U52 (N_52,In_2126,In_1258);
xnor U53 (N_53,In_845,In_915);
nor U54 (N_54,In_1756,In_1362);
nor U55 (N_55,In_1293,In_2232);
nor U56 (N_56,In_1597,In_120);
nor U57 (N_57,In_1286,In_2400);
nand U58 (N_58,In_1403,In_1533);
or U59 (N_59,In_889,In_1762);
xor U60 (N_60,In_2259,In_1032);
and U61 (N_61,In_1556,In_2434);
xnor U62 (N_62,In_2139,In_1285);
nor U63 (N_63,In_122,In_1482);
or U64 (N_64,In_628,In_1595);
nand U65 (N_65,In_2210,In_474);
and U66 (N_66,In_1050,In_2273);
nand U67 (N_67,In_2033,In_1348);
nor U68 (N_68,In_140,In_1891);
and U69 (N_69,In_661,In_991);
and U70 (N_70,In_569,In_662);
nand U71 (N_71,In_728,In_2427);
or U72 (N_72,In_2007,In_2329);
nor U73 (N_73,In_70,In_2280);
or U74 (N_74,In_1856,In_2282);
nor U75 (N_75,In_2158,In_419);
xor U76 (N_76,In_2492,In_1919);
or U77 (N_77,In_1042,In_2392);
nor U78 (N_78,In_984,In_2157);
nand U79 (N_79,In_302,In_1198);
or U80 (N_80,In_2398,In_928);
or U81 (N_81,In_1989,In_163);
or U82 (N_82,In_503,In_1070);
xor U83 (N_83,In_960,In_542);
and U84 (N_84,In_879,In_1177);
nand U85 (N_85,In_1107,In_189);
xnor U86 (N_86,In_1067,In_2040);
nor U87 (N_87,In_2230,In_872);
nand U88 (N_88,In_1769,In_1094);
nand U89 (N_89,In_2130,In_630);
and U90 (N_90,In_1438,In_276);
or U91 (N_91,In_129,In_1211);
nor U92 (N_92,In_396,In_2393);
xor U93 (N_93,In_1755,In_30);
and U94 (N_94,In_395,In_102);
or U95 (N_95,In_2240,In_2145);
nor U96 (N_96,In_786,In_2405);
or U97 (N_97,In_1263,In_366);
or U98 (N_98,In_1686,In_2233);
and U99 (N_99,In_1677,In_386);
or U100 (N_100,In_1065,In_155);
and U101 (N_101,In_772,In_1134);
or U102 (N_102,In_933,In_2307);
nor U103 (N_103,In_220,In_697);
or U104 (N_104,In_498,In_1206);
xnor U105 (N_105,In_596,In_139);
nor U106 (N_106,In_574,In_2483);
nand U107 (N_107,In_421,In_1749);
xnor U108 (N_108,In_1129,In_1529);
and U109 (N_109,In_654,In_2475);
and U110 (N_110,In_1862,In_1074);
nand U111 (N_111,In_531,In_1879);
and U112 (N_112,In_58,In_215);
nand U113 (N_113,In_1713,In_2431);
xor U114 (N_114,In_2346,In_1930);
or U115 (N_115,In_506,In_1666);
and U116 (N_116,In_935,In_602);
nor U117 (N_117,In_1709,In_878);
nor U118 (N_118,In_1814,In_1851);
nand U119 (N_119,In_1075,In_1440);
nor U120 (N_120,In_1733,In_944);
xnor U121 (N_121,In_1858,In_724);
or U122 (N_122,In_2344,In_619);
xnor U123 (N_123,In_918,In_432);
nor U124 (N_124,In_2010,In_2044);
or U125 (N_125,In_159,In_1151);
xnor U126 (N_126,In_970,In_2097);
xnor U127 (N_127,In_411,In_26);
xor U128 (N_128,In_2121,In_2343);
and U129 (N_129,In_880,In_35);
xor U130 (N_130,In_121,In_1185);
nor U131 (N_131,In_1542,In_1261);
nor U132 (N_132,In_1646,In_2422);
and U133 (N_133,In_2000,In_28);
xnor U134 (N_134,In_1832,In_1275);
or U135 (N_135,In_1117,In_1548);
or U136 (N_136,In_951,In_443);
nand U137 (N_137,In_992,In_393);
and U138 (N_138,In_1267,In_1602);
xor U139 (N_139,In_264,In_1958);
xor U140 (N_140,In_465,In_1173);
nand U141 (N_141,In_2229,In_966);
or U142 (N_142,In_92,In_644);
nand U143 (N_143,In_2275,In_2094);
nand U144 (N_144,In_855,In_1265);
xor U145 (N_145,In_59,In_481);
or U146 (N_146,In_200,In_1239);
nor U147 (N_147,In_2191,In_51);
xor U148 (N_148,In_1627,In_1121);
or U149 (N_149,In_1271,In_2270);
or U150 (N_150,In_227,In_1090);
nor U151 (N_151,In_1658,In_864);
and U152 (N_152,In_528,In_978);
nor U153 (N_153,In_1169,In_2016);
nor U154 (N_154,In_93,In_2134);
and U155 (N_155,In_1489,In_871);
nor U156 (N_156,In_1260,In_2378);
nand U157 (N_157,In_2179,In_948);
nand U158 (N_158,In_126,In_2418);
xor U159 (N_159,In_424,In_1160);
or U160 (N_160,In_1819,In_370);
or U161 (N_161,In_1472,In_1182);
and U162 (N_162,In_910,In_1812);
and U163 (N_163,In_987,In_775);
or U164 (N_164,In_1601,In_909);
nand U165 (N_165,In_1576,In_1643);
nand U166 (N_166,In_1158,In_2051);
xnor U167 (N_167,In_2142,In_234);
nor U168 (N_168,In_1096,In_1526);
and U169 (N_169,In_240,In_1017);
xnor U170 (N_170,In_2314,In_2034);
and U171 (N_171,In_1184,In_577);
and U172 (N_172,In_275,In_2473);
xnor U173 (N_173,In_547,In_2242);
nor U174 (N_174,In_1353,In_176);
nor U175 (N_175,In_2212,In_735);
or U176 (N_176,In_530,In_2339);
xor U177 (N_177,In_1560,In_983);
nand U178 (N_178,In_98,In_488);
xnor U179 (N_179,In_1728,In_678);
nand U180 (N_180,In_1194,In_326);
nand U181 (N_181,In_343,In_974);
xor U182 (N_182,In_2257,In_1327);
nor U183 (N_183,In_952,In_911);
or U184 (N_184,In_1101,In_19);
nor U185 (N_185,In_824,In_342);
nand U186 (N_186,In_1113,In_821);
xnor U187 (N_187,In_44,In_535);
xnor U188 (N_188,In_1705,In_1857);
and U189 (N_189,In_1305,In_119);
nand U190 (N_190,In_1810,In_2155);
or U191 (N_191,In_1869,In_1673);
nand U192 (N_192,In_514,In_1543);
and U193 (N_193,In_1479,In_1785);
nand U194 (N_194,In_621,In_1599);
xor U195 (N_195,In_891,In_2127);
nand U196 (N_196,In_1906,In_104);
xnor U197 (N_197,In_1896,In_2370);
nor U198 (N_198,In_1849,In_1702);
nand U199 (N_199,In_144,In_936);
or U200 (N_200,In_1176,In_610);
or U201 (N_201,In_1414,In_2053);
and U202 (N_202,In_1469,In_269);
nand U203 (N_203,In_731,In_209);
nor U204 (N_204,In_1833,In_1624);
and U205 (N_205,In_2361,In_2439);
or U206 (N_206,In_1283,In_1782);
or U207 (N_207,In_8,In_2246);
and U208 (N_208,In_2383,In_2099);
nor U209 (N_209,In_655,In_1621);
nand U210 (N_210,In_777,In_1852);
xor U211 (N_211,In_67,In_1156);
nor U212 (N_212,In_1947,In_1780);
xnor U213 (N_213,In_1080,In_2075);
nand U214 (N_214,In_22,In_1339);
xor U215 (N_215,In_172,In_1886);
nor U216 (N_216,In_2103,In_68);
nand U217 (N_217,In_1365,In_1667);
nand U218 (N_218,In_539,In_545);
nand U219 (N_219,In_903,In_441);
or U220 (N_220,In_1034,In_1056);
or U221 (N_221,In_907,In_392);
nor U222 (N_222,In_1337,In_527);
or U223 (N_223,In_757,In_1828);
or U224 (N_224,In_1086,In_288);
nand U225 (N_225,In_1227,In_435);
nor U226 (N_226,In_515,In_241);
nor U227 (N_227,In_2237,In_739);
or U228 (N_228,In_842,In_685);
xor U229 (N_229,In_2018,In_2328);
xnor U230 (N_230,In_762,In_1064);
xor U231 (N_231,In_1207,In_1104);
xnor U232 (N_232,In_2029,In_2480);
xor U233 (N_233,In_305,In_2079);
nand U234 (N_234,In_1689,In_2188);
or U235 (N_235,In_1213,In_1736);
and U236 (N_236,In_1111,In_712);
and U237 (N_237,In_1025,In_11);
nor U238 (N_238,In_1000,In_460);
xor U239 (N_239,In_1091,In_1256);
nand U240 (N_240,In_565,In_1396);
nand U241 (N_241,In_1591,In_1638);
nor U242 (N_242,In_612,In_1737);
nor U243 (N_243,In_764,In_298);
xnor U244 (N_244,In_459,In_862);
xnor U245 (N_245,In_1486,In_1954);
nand U246 (N_246,In_1953,In_2493);
xnor U247 (N_247,In_1701,In_648);
nor U248 (N_248,In_1521,In_2243);
xor U249 (N_249,In_469,In_1888);
and U250 (N_250,In_895,In_1610);
xor U251 (N_251,In_2274,In_806);
or U252 (N_252,In_483,In_1029);
or U253 (N_253,In_2388,In_1924);
xor U254 (N_254,In_1490,In_318);
nor U255 (N_255,In_585,In_2235);
xor U256 (N_256,In_2202,In_1149);
nor U257 (N_257,In_639,In_1987);
nor U258 (N_258,In_1309,In_282);
and U259 (N_259,In_1495,In_826);
and U260 (N_260,In_1600,In_869);
nor U261 (N_261,In_892,In_546);
or U262 (N_262,In_1625,In_2069);
xor U263 (N_263,In_2047,In_1043);
nor U264 (N_264,In_1335,In_1800);
nor U265 (N_265,In_80,In_1512);
nor U266 (N_266,In_1188,In_601);
and U267 (N_267,In_1497,In_849);
nand U268 (N_268,In_124,In_445);
or U269 (N_269,In_1456,In_2156);
or U270 (N_270,In_152,In_2283);
nor U271 (N_271,In_1341,In_303);
nand U272 (N_272,In_193,In_2305);
nor U273 (N_273,In_919,In_2009);
nand U274 (N_274,In_1680,In_1741);
nor U275 (N_275,In_2481,In_2023);
nor U276 (N_276,In_2124,In_709);
or U277 (N_277,In_33,In_2181);
nand U278 (N_278,In_1272,In_570);
or U279 (N_279,In_778,In_239);
nor U280 (N_280,In_169,In_618);
nand U281 (N_281,In_2447,In_2495);
or U282 (N_282,In_2064,In_150);
nor U283 (N_283,In_812,In_1864);
nand U284 (N_284,In_489,In_881);
or U285 (N_285,In_859,In_312);
or U286 (N_286,In_1855,In_2381);
xor U287 (N_287,In_1975,In_2036);
nand U288 (N_288,In_1170,In_180);
nand U289 (N_289,In_2006,In_187);
and U290 (N_290,In_624,In_549);
xnor U291 (N_291,In_1407,In_805);
nand U292 (N_292,In_633,In_428);
nor U293 (N_293,In_2291,In_249);
nand U294 (N_294,In_1369,In_765);
and U295 (N_295,In_389,In_339);
and U296 (N_296,In_1083,In_1389);
or U297 (N_297,In_203,In_2465);
nand U298 (N_298,In_1829,In_1312);
nor U299 (N_299,In_1161,In_259);
or U300 (N_300,In_930,In_744);
xnor U301 (N_301,In_1427,In_1307);
or U302 (N_302,In_2138,In_2399);
and U303 (N_303,In_1932,In_1847);
xnor U304 (N_304,In_153,In_663);
nor U305 (N_305,In_74,In_1536);
and U306 (N_306,In_293,In_2019);
and U307 (N_307,In_253,In_1606);
nand U308 (N_308,In_1985,In_1742);
nor U309 (N_309,In_1817,In_2433);
nand U310 (N_310,In_1834,In_283);
nand U311 (N_311,In_1352,In_1253);
nand U312 (N_312,In_1897,In_716);
nor U313 (N_313,In_519,In_835);
nor U314 (N_314,In_785,In_1779);
nand U315 (N_315,In_946,In_2027);
nor U316 (N_316,In_922,In_1063);
and U317 (N_317,In_2227,In_1128);
or U318 (N_318,In_416,In_1498);
xor U319 (N_319,In_484,In_611);
and U320 (N_320,In_736,In_776);
xnor U321 (N_321,In_1060,In_1290);
and U322 (N_322,In_2248,In_1138);
or U323 (N_323,In_1870,In_1910);
or U324 (N_324,In_784,In_1171);
xnor U325 (N_325,In_2135,In_2382);
nor U326 (N_326,In_164,In_555);
nor U327 (N_327,In_837,In_2411);
xnor U328 (N_328,In_453,In_1269);
or U329 (N_329,In_1722,In_492);
and U330 (N_330,In_1445,In_995);
xnor U331 (N_331,In_1216,In_1528);
xor U332 (N_332,In_1883,In_605);
xnor U333 (N_333,In_1802,In_1463);
and U334 (N_334,In_1381,In_248);
xor U335 (N_335,In_2466,In_541);
nor U336 (N_336,In_2470,In_2334);
xnor U337 (N_337,In_230,In_62);
nand U338 (N_338,In_1907,In_1088);
xor U339 (N_339,In_2204,In_2389);
nand U340 (N_340,In_130,In_2070);
nor U341 (N_341,In_734,In_560);
nor U342 (N_342,In_1687,In_963);
xnor U343 (N_343,In_1633,In_16);
xnor U344 (N_344,In_1822,In_477);
and U345 (N_345,In_562,In_1843);
nor U346 (N_346,In_1187,In_2083);
nand U347 (N_347,In_1840,In_1531);
xor U348 (N_348,In_2195,In_1904);
nor U349 (N_349,In_1478,In_359);
nand U350 (N_350,In_2115,In_2368);
xnor U351 (N_351,In_1977,In_1152);
xor U352 (N_352,In_289,In_2357);
and U353 (N_353,In_2395,In_2113);
nand U354 (N_354,In_1991,In_76);
nor U355 (N_355,In_2436,In_1234);
xnor U356 (N_356,In_224,In_2298);
nand U357 (N_357,In_37,In_2359);
nand U358 (N_358,In_692,In_252);
or U359 (N_359,In_1842,In_1517);
and U360 (N_360,In_2182,In_1719);
nor U361 (N_361,In_1890,In_486);
xnor U362 (N_362,In_479,In_927);
or U363 (N_363,In_24,In_133);
nand U364 (N_364,In_2123,In_1202);
nor U365 (N_365,In_1506,In_1386);
nand U366 (N_366,In_1552,In_1683);
and U367 (N_367,In_976,In_1297);
nand U368 (N_368,In_43,In_174);
or U369 (N_369,In_1662,In_563);
nand U370 (N_370,In_1608,In_2310);
nor U371 (N_371,In_473,In_1248);
and U372 (N_372,In_1228,In_524);
xor U373 (N_373,In_2120,In_313);
or U374 (N_374,In_1220,In_627);
xnor U375 (N_375,In_1519,In_998);
nor U376 (N_376,In_1190,In_1108);
and U377 (N_377,In_613,In_740);
and U378 (N_378,In_1679,In_1371);
xor U379 (N_379,In_158,In_719);
or U380 (N_380,In_1532,In_667);
and U381 (N_381,In_1006,In_843);
xor U382 (N_382,In_2011,In_2286);
and U383 (N_383,In_1745,In_1962);
or U384 (N_384,In_658,In_1923);
nand U385 (N_385,In_1321,In_2108);
or U386 (N_386,In_760,In_183);
and U387 (N_387,In_1073,In_360);
or U388 (N_388,In_1446,In_1825);
nor U389 (N_389,In_1058,In_1768);
and U390 (N_390,In_1114,In_962);
and U391 (N_391,In_1148,In_2444);
and U392 (N_392,In_2407,In_1580);
or U393 (N_393,In_1081,In_310);
nor U394 (N_394,In_1944,In_1648);
nor U395 (N_395,In_1671,In_247);
or U396 (N_396,In_1708,In_2349);
nand U397 (N_397,In_1483,In_766);
xor U398 (N_398,In_873,In_1603);
and U399 (N_399,In_270,In_699);
xor U400 (N_400,In_2301,In_2272);
nand U401 (N_401,In_1415,In_1379);
xnor U402 (N_402,In_271,In_1640);
or U403 (N_403,In_1392,In_1420);
nand U404 (N_404,In_2043,In_73);
nand U405 (N_405,In_78,In_1417);
nor U406 (N_406,In_1476,In_727);
xor U407 (N_407,In_2429,In_664);
and U408 (N_408,In_1848,In_2039);
and U409 (N_409,In_846,In_1986);
nand U410 (N_410,In_1147,In_1178);
or U411 (N_411,In_1133,In_1541);
nor U412 (N_412,In_1295,In_943);
nand U413 (N_413,In_88,In_1098);
and U414 (N_414,In_711,In_1019);
or U415 (N_415,In_1399,In_1815);
xor U416 (N_416,In_1300,In_69);
nor U417 (N_417,In_1022,In_1957);
and U418 (N_418,In_1008,In_300);
nor U419 (N_419,In_818,In_448);
or U420 (N_420,In_1794,In_2164);
xor U421 (N_421,In_368,In_1278);
or U422 (N_422,In_2147,In_502);
nand U423 (N_423,In_875,In_2213);
and U424 (N_424,In_1903,In_1209);
or U425 (N_425,In_1480,In_1565);
nand U426 (N_426,In_1926,In_1137);
xor U427 (N_427,In_1558,In_2266);
xnor U428 (N_428,In_191,In_795);
nand U429 (N_429,In_2153,In_1193);
xnor U430 (N_430,In_333,In_1912);
or U431 (N_431,In_1411,In_2199);
xor U432 (N_432,In_2284,In_2425);
or U433 (N_433,In_1659,In_1831);
and U434 (N_434,In_1895,In_487);
and U435 (N_435,In_412,In_1804);
nand U436 (N_436,In_1505,In_1394);
nand U437 (N_437,In_245,In_1681);
and U438 (N_438,In_780,In_1240);
or U439 (N_439,In_2261,In_1009);
or U440 (N_440,In_10,In_1015);
nor U441 (N_441,In_212,In_1795);
nand U442 (N_442,In_2498,In_2348);
nor U443 (N_443,In_2256,In_2253);
and U444 (N_444,In_851,In_1798);
and U445 (N_445,In_2453,In_1873);
xnor U446 (N_446,In_2358,In_60);
or U447 (N_447,In_1577,In_2110);
xnor U448 (N_448,In_801,In_482);
nand U449 (N_449,In_316,In_827);
or U450 (N_450,In_1118,In_1301);
and U451 (N_451,In_1229,In_1661);
xnor U452 (N_452,In_1324,In_2285);
nand U453 (N_453,In_108,In_1007);
or U454 (N_454,In_1868,In_1845);
nand U455 (N_455,In_750,In_1437);
or U456 (N_456,In_2168,In_290);
and U457 (N_457,In_2002,In_50);
xnor U458 (N_458,In_1846,In_2289);
and U459 (N_459,In_1436,In_1502);
and U460 (N_460,In_1511,In_507);
nand U461 (N_461,In_829,In_847);
nand U462 (N_462,In_1314,In_1778);
nor U463 (N_463,In_349,In_1751);
nand U464 (N_464,In_2351,In_763);
or U465 (N_465,In_1066,In_1346);
xnor U466 (N_466,In_1761,In_457);
or U467 (N_467,In_1690,In_2028);
or U468 (N_468,In_743,In_1328);
nand U469 (N_469,In_1494,In_580);
and U470 (N_470,In_1893,In_1550);
and U471 (N_471,In_2129,In_1753);
and U472 (N_472,In_647,In_746);
or U473 (N_473,In_1911,In_2445);
or U474 (N_474,In_1377,In_1046);
and U475 (N_475,In_625,In_410);
xor U476 (N_476,In_540,In_905);
nor U477 (N_477,In_2420,In_1639);
and U478 (N_478,In_1718,In_1827);
nor U479 (N_479,In_1288,In_2321);
nand U480 (N_480,In_931,In_950);
and U481 (N_481,In_14,In_2068);
nor U482 (N_482,In_1759,In_2165);
or U483 (N_483,In_631,In_61);
nor U484 (N_484,In_645,In_1928);
and U485 (N_485,In_2193,In_2017);
xnor U486 (N_486,In_1995,In_345);
and U487 (N_487,In_518,In_401);
and U488 (N_488,In_2278,In_31);
and U489 (N_489,In_2189,In_1306);
xnor U490 (N_490,In_2058,In_942);
nand U491 (N_491,In_1725,In_1100);
and U492 (N_492,In_2364,In_2476);
xnor U493 (N_493,In_49,In_285);
nand U494 (N_494,In_323,In_1882);
or U495 (N_495,In_2323,In_199);
nand U496 (N_496,In_1583,In_2457);
and U497 (N_497,In_1540,In_1450);
xnor U498 (N_498,In_2062,In_551);
xnor U499 (N_499,In_1808,In_674);
nand U500 (N_500,In_1539,In_1553);
nand U501 (N_501,In_472,In_954);
nand U502 (N_502,In_42,In_2149);
nand U503 (N_503,In_986,In_405);
and U504 (N_504,In_23,In_823);
xor U505 (N_505,In_431,In_670);
and U506 (N_506,In_1653,In_749);
nor U507 (N_507,In_2384,In_1222);
and U508 (N_508,In_358,In_1370);
xnor U509 (N_509,In_2360,In_1525);
or U510 (N_510,In_2146,In_2144);
nor U511 (N_511,In_165,In_1537);
nor U512 (N_512,In_2437,In_21);
xor U513 (N_513,In_904,In_299);
or U514 (N_514,In_1033,In_1455);
nor U515 (N_515,In_117,In_1452);
nand U516 (N_516,In_188,In_1935);
nor U517 (N_517,In_1534,In_1145);
or U518 (N_518,In_1071,In_195);
xnor U519 (N_519,In_1281,In_1783);
nor U520 (N_520,In_620,In_787);
nand U521 (N_521,In_1250,In_1703);
nor U522 (N_522,In_1706,In_336);
or U523 (N_523,In_1201,In_2484);
nand U524 (N_524,In_242,In_1549);
nand U525 (N_525,In_1865,In_36);
xor U526 (N_526,In_1245,In_1574);
or U527 (N_527,In_2464,In_2373);
nor U528 (N_528,In_953,In_816);
and U529 (N_529,In_870,In_362);
and U530 (N_530,In_2221,In_646);
nand U531 (N_531,In_1223,In_687);
or U532 (N_532,In_286,In_1791);
nor U533 (N_533,In_1045,In_1270);
or U534 (N_534,In_1296,In_1254);
xnor U535 (N_535,In_1039,In_185);
and U536 (N_536,In_1500,In_1226);
nand U537 (N_537,In_2319,In_184);
nor U538 (N_538,In_1885,In_1084);
or U539 (N_539,In_1927,In_1950);
nor U540 (N_540,In_1077,In_1429);
and U541 (N_541,In_588,In_1503);
nor U542 (N_542,In_1393,In_236);
or U543 (N_543,In_1976,In_1023);
nand U544 (N_544,In_79,In_2271);
or U545 (N_545,In_913,In_1788);
or U546 (N_546,In_2125,In_1587);
or U547 (N_547,In_1674,In_2394);
nor U548 (N_548,In_1038,In_2200);
and U549 (N_549,In_1465,In_1789);
nor U550 (N_550,In_1315,In_404);
and U551 (N_551,In_109,In_1329);
nor U552 (N_552,In_964,In_1747);
xnor U553 (N_553,In_399,In_497);
xor U554 (N_554,In_2320,In_961);
or U555 (N_555,In_2008,In_197);
and U556 (N_556,In_1347,In_1447);
or U557 (N_557,In_1485,In_854);
nand U558 (N_558,In_141,In_2208);
or U559 (N_559,In_840,In_255);
xor U560 (N_560,In_1375,In_990);
xor U561 (N_561,In_694,In_1937);
nand U562 (N_562,In_883,In_717);
nor U563 (N_563,In_454,In_1515);
nor U564 (N_564,In_499,In_2454);
nand U565 (N_565,In_2299,In_1634);
nand U566 (N_566,In_2251,In_756);
nor U567 (N_567,In_1492,In_1338);
nor U568 (N_568,In_1996,In_1821);
or U569 (N_569,In_2219,In_2086);
xnor U570 (N_570,In_113,In_194);
or U571 (N_571,In_1434,In_56);
nor U572 (N_572,In_1391,In_464);
nor U573 (N_573,In_564,In_607);
xor U574 (N_574,In_1344,In_2183);
or U575 (N_575,In_205,In_2265);
nor U576 (N_576,In_1125,In_82);
or U577 (N_577,In_2055,In_2112);
or U578 (N_578,In_244,In_494);
and U579 (N_579,In_2366,In_2176);
or U580 (N_580,In_383,In_1754);
xor U581 (N_581,In_1654,In_836);
xnor U582 (N_582,In_956,In_1569);
or U583 (N_583,In_2020,In_382);
nor U584 (N_584,In_2192,In_1772);
nor U585 (N_585,In_1357,In_123);
or U586 (N_586,In_2052,In_2311);
nand U587 (N_587,In_1838,In_2258);
nor U588 (N_588,In_2045,In_1345);
nand U589 (N_589,In_2102,In_2306);
xor U590 (N_590,In_4,In_1830);
xnor U591 (N_591,In_1488,In_53);
and U592 (N_592,In_1428,In_2117);
or U593 (N_593,In_886,In_2424);
xor U594 (N_594,In_2175,In_2264);
nor U595 (N_595,In_972,In_589);
xnor U596 (N_596,In_1711,In_491);
xnor U597 (N_597,In_1656,In_1934);
or U598 (N_598,In_190,In_1243);
nor U599 (N_599,In_231,In_614);
xor U600 (N_600,In_277,In_1605);
xor U601 (N_601,In_2267,In_675);
nor U602 (N_602,In_20,In_1774);
and U603 (N_603,In_2252,In_27);
nor U604 (N_604,In_221,In_598);
or U605 (N_605,In_550,In_45);
nand U606 (N_606,In_1509,In_2312);
and U607 (N_607,In_1908,In_2005);
or U608 (N_608,In_1586,In_2255);
and U609 (N_609,In_1963,In_914);
nor U610 (N_610,In_1433,In_311);
nand U611 (N_611,In_512,In_774);
nor U612 (N_612,In_1004,In_1183);
nand U613 (N_613,In_103,In_101);
or U614 (N_614,In_1217,In_1473);
xnor U615 (N_615,In_1116,In_1663);
nor U616 (N_616,In_1252,In_1124);
xor U617 (N_617,In_1806,In_771);
nor U618 (N_618,In_1920,In_480);
and U619 (N_619,In_1451,In_798);
nand U620 (N_620,In_996,In_830);
or U621 (N_621,In_650,In_1308);
nor U622 (N_622,In_444,In_1796);
or U623 (N_623,In_55,In_1763);
xnor U624 (N_624,In_637,In_1637);
nor U625 (N_625,In_582,In_1439);
or U626 (N_626,In_1670,In_81);
nand U627 (N_627,In_1655,In_237);
or U628 (N_628,In_423,In_1435);
and U629 (N_629,In_1418,In_1887);
or U630 (N_630,In_2474,In_476);
nor U631 (N_631,In_781,In_1518);
xor U632 (N_632,In_2281,In_1641);
or U633 (N_633,In_1900,In_2460);
nor U634 (N_634,In_773,In_2244);
and U635 (N_635,In_705,In_523);
and U636 (N_636,In_344,In_1913);
nor U637 (N_637,In_817,In_1232);
nand U638 (N_638,In_1162,In_1432);
nor U639 (N_639,In_2448,In_1021);
nand U640 (N_640,In_422,In_1037);
xnor U641 (N_641,In_38,In_1257);
or U642 (N_642,In_1562,In_2304);
or U643 (N_643,In_924,In_916);
or U644 (N_644,In_1334,In_2297);
and U645 (N_645,In_1598,In_1316);
and U646 (N_646,In_2078,In_160);
xor U647 (N_647,In_2118,In_604);
nand U648 (N_648,In_1336,In_2087);
xnor U649 (N_649,In_814,In_179);
nand U650 (N_650,In_451,In_17);
or U651 (N_651,In_1750,In_354);
or U652 (N_652,In_808,In_114);
nand U653 (N_653,In_355,In_2057);
nand U654 (N_654,In_1400,In_1457);
and U655 (N_655,In_1404,In_623);
and U656 (N_656,In_2211,In_1318);
xnor U657 (N_657,In_1547,In_7);
nand U658 (N_658,In_1551,In_1310);
and U659 (N_659,In_2417,In_25);
xor U660 (N_660,In_2186,In_387);
nor U661 (N_661,In_2421,In_2414);
and U662 (N_662,In_659,In_2468);
nand U663 (N_663,In_1915,In_1983);
or U664 (N_664,In_1921,In_722);
or U665 (N_665,In_543,In_1323);
or U666 (N_666,In_700,In_463);
nand U667 (N_667,In_1105,In_1035);
xnor U668 (N_668,In_989,In_1233);
nand U669 (N_669,In_1501,In_732);
xnor U670 (N_670,In_520,In_1467);
nor U671 (N_671,In_1055,In_1803);
nand U672 (N_672,In_2,In_985);
and U673 (N_673,In_1970,In_584);
nor U674 (N_674,In_307,In_198);
and U675 (N_675,In_890,In_1444);
and U676 (N_676,In_553,In_206);
nor U677 (N_677,In_2239,In_606);
nor U678 (N_678,In_599,In_1642);
xnor U679 (N_679,In_1441,In_347);
xnor U680 (N_680,In_1203,In_1878);
xnor U681 (N_681,In_1048,In_720);
nand U682 (N_682,In_1902,In_768);
or U683 (N_683,In_1165,In_1062);
xnor U684 (N_684,In_1664,In_325);
xor U685 (N_685,In_1,In_938);
nand U686 (N_686,In_1844,In_1880);
nor U687 (N_687,In_1106,In_1766);
or U688 (N_688,In_467,In_1771);
xor U689 (N_689,In_751,In_522);
nor U690 (N_690,In_1123,In_29);
xor U691 (N_691,In_272,In_2486);
nor U692 (N_692,In_632,In_2003);
and U693 (N_693,In_748,In_1011);
nand U694 (N_694,In_175,In_1564);
nand U695 (N_695,In_2106,In_437);
or U696 (N_696,In_887,In_666);
or U697 (N_697,In_427,In_306);
or U698 (N_698,In_468,In_268);
or U699 (N_699,In_1298,In_1652);
nor U700 (N_700,In_1368,In_1669);
and U701 (N_701,In_1787,In_761);
xnor U702 (N_702,In_1972,In_1945);
nand U703 (N_703,In_2214,In_47);
and U704 (N_704,In_689,In_576);
or U705 (N_705,In_820,In_334);
nand U706 (N_706,In_2472,In_2317);
nand U707 (N_707,In_2025,In_2315);
nand U708 (N_708,In_1554,In_72);
or U709 (N_709,In_1898,In_1949);
nand U710 (N_710,In_204,In_2236);
and U711 (N_711,In_364,In_1131);
or U712 (N_712,In_733,In_1740);
or U713 (N_713,In_15,In_2385);
xnor U714 (N_714,In_1099,In_1320);
nand U715 (N_715,In_1775,In_1726);
xnor U716 (N_716,In_844,In_1317);
or U717 (N_717,In_857,In_18);
nor U718 (N_718,In_1734,In_810);
nor U719 (N_719,In_2065,In_63);
nor U720 (N_720,In_1573,In_138);
nand U721 (N_721,In_2050,In_537);
nor U722 (N_722,In_696,In_446);
xnor U723 (N_723,In_425,In_752);
nor U724 (N_724,In_1287,In_1130);
and U725 (N_725,In_568,In_1835);
or U726 (N_726,In_2338,In_1933);
nand U727 (N_727,In_1423,In_2461);
or U728 (N_728,In_745,In_1914);
and U729 (N_729,In_1631,In_1623);
xnor U730 (N_730,In_1967,In_1186);
nor U731 (N_731,In_2111,In_1527);
nor U732 (N_732,In_2038,In_1195);
nand U733 (N_733,In_1443,In_83);
or U734 (N_734,In_1072,In_1508);
or U735 (N_735,In_1292,In_2178);
and U736 (N_736,In_1714,In_403);
and U737 (N_737,In_89,In_85);
nor U738 (N_738,In_173,In_1102);
xnor U739 (N_739,In_1697,In_363);
nand U740 (N_740,In_2180,In_71);
xnor U741 (N_741,In_2030,In_438);
xnor U742 (N_742,In_2463,In_2067);
nand U743 (N_743,In_1236,In_327);
xor U744 (N_744,In_1020,In_2222);
and U745 (N_745,In_1241,In_48);
nand U746 (N_746,In_2172,In_1922);
xor U747 (N_747,In_521,In_1629);
xnor U748 (N_748,In_447,In_538);
or U749 (N_749,In_192,In_341);
nand U750 (N_750,In_1361,In_110);
nand U751 (N_751,In_2060,In_683);
xor U752 (N_752,In_1461,In_1235);
nor U753 (N_753,In_1383,In_2330);
nor U754 (N_754,In_1068,In_819);
xnor U755 (N_755,In_2318,In_1717);
or U756 (N_756,In_1012,In_471);
or U757 (N_757,In_1694,In_533);
and U758 (N_758,In_2263,In_314);
nor U759 (N_759,In_1496,In_1390);
nand U760 (N_760,In_1951,In_1425);
and U761 (N_761,In_86,In_603);
and U762 (N_762,In_1952,In_1054);
or U763 (N_763,In_380,In_291);
and U764 (N_764,In_939,In_2293);
nand U765 (N_765,In_2162,In_1238);
nand U766 (N_766,In_378,In_1331);
or U767 (N_767,In_317,In_332);
and U768 (N_768,In_1163,In_1729);
nor U769 (N_769,In_759,In_1466);
and U770 (N_770,In_2071,In_848);
and U771 (N_771,In_2374,In_2026);
nand U772 (N_772,In_284,In_1559);
xor U773 (N_773,In_2441,In_2035);
nor U774 (N_774,In_1251,In_1579);
or U775 (N_775,In_1892,In_581);
xor U776 (N_776,In_2059,In_1140);
nand U777 (N_777,In_2093,In_1929);
xnor U778 (N_778,In_796,In_229);
xnor U779 (N_779,In_1424,In_1999);
or U780 (N_780,In_171,In_295);
nand U781 (N_781,In_1731,In_1946);
and U782 (N_782,In_877,In_99);
and U783 (N_783,In_797,In_1960);
and U784 (N_784,In_2101,In_208);
or U785 (N_785,In_1053,In_1426);
xor U786 (N_786,In_1136,In_1453);
xnor U787 (N_787,In_2455,In_2497);
nand U788 (N_788,In_372,In_1635);
and U789 (N_789,In_1412,In_475);
nand U790 (N_790,In_1909,In_2488);
nand U791 (N_791,In_1342,In_1982);
nor U792 (N_792,In_1311,In_2198);
xor U793 (N_793,In_1861,In_1948);
and U794 (N_794,In_2088,In_2001);
xnor U795 (N_795,In_1675,In_858);
or U796 (N_796,In_2491,In_2241);
nor U797 (N_797,In_508,In_643);
xor U798 (N_798,In_2196,In_1570);
nand U799 (N_799,In_1695,In_1820);
xor U800 (N_800,In_2496,In_900);
or U801 (N_801,In_178,In_406);
and U802 (N_802,In_794,In_90);
and U803 (N_803,In_297,In_1470);
nor U804 (N_804,In_2063,In_1363);
xnor U805 (N_805,In_578,In_1567);
and U806 (N_806,In_1401,In_331);
nor U807 (N_807,In_52,In_1115);
and U808 (N_808,In_1351,In_1786);
nand U809 (N_809,In_1979,In_1384);
and U810 (N_810,In_1961,In_941);
or U811 (N_811,In_496,In_1454);
nor U812 (N_812,In_1752,In_2250);
and U813 (N_813,In_947,In_9);
or U814 (N_814,In_2287,In_2390);
nand U815 (N_815,In_1973,In_753);
xor U816 (N_816,In_526,In_676);
nand U817 (N_817,In_671,In_1262);
nor U818 (N_818,In_95,In_1459);
nand U819 (N_819,In_1504,In_2049);
nand U820 (N_820,In_510,In_1572);
xor U821 (N_821,In_407,In_1993);
xor U822 (N_822,In_207,In_591);
and U823 (N_823,In_1997,In_713);
nor U824 (N_824,In_1049,In_118);
xor U825 (N_825,In_1224,In_1616);
or U826 (N_826,In_1302,In_1644);
and U827 (N_827,In_1744,In_1359);
nand U828 (N_828,In_525,In_673);
xor U829 (N_829,In_2013,In_287);
xor U830 (N_830,In_850,In_267);
or U831 (N_831,In_351,In_2479);
nand U832 (N_832,In_1167,In_1585);
nand U833 (N_833,In_397,In_87);
xnor U834 (N_834,In_1571,In_994);
xnor U835 (N_835,In_2409,In_2467);
and U836 (N_836,In_1524,In_1340);
xnor U837 (N_837,In_1615,In_1095);
xnor U838 (N_838,In_2369,In_594);
or U839 (N_839,In_2122,In_2452);
nor U840 (N_840,In_371,In_2353);
or U841 (N_841,In_949,In_1279);
nand U842 (N_842,In_1707,In_1264);
or U843 (N_843,In_2316,In_698);
nor U844 (N_844,In_2428,In_1699);
or U845 (N_845,In_154,In_1069);
nand U846 (N_846,In_1322,In_1448);
nor U847 (N_847,In_799,In_1818);
and U848 (N_848,In_2313,In_2406);
or U849 (N_849,In_1589,In_434);
and U850 (N_850,In_1974,In_754);
xnor U851 (N_851,In_1406,In_1356);
or U852 (N_852,In_0,In_1611);
xnor U853 (N_853,In_1594,In_2203);
or U854 (N_854,In_2169,In_321);
xor U855 (N_855,In_1650,In_1319);
nor U856 (N_856,In_2426,In_1764);
xor U857 (N_857,In_959,In_196);
xor U858 (N_858,In_1372,In_1360);
nand U859 (N_859,In_1618,In_157);
or U860 (N_860,In_926,In_934);
nor U861 (N_861,In_902,In_2326);
xnor U862 (N_862,In_1575,In_148);
and U863 (N_863,In_418,In_2469);
or U864 (N_864,In_2218,In_2081);
xnor U865 (N_865,In_105,In_888);
nand U866 (N_866,In_629,In_1231);
xor U867 (N_867,In_1159,In_718);
nand U868 (N_868,In_75,In_1555);
xnor U869 (N_869,In_408,In_2054);
nor U870 (N_870,In_1918,In_1700);
nand U871 (N_871,In_2231,In_1174);
nor U872 (N_872,In_1041,In_1513);
or U873 (N_873,In_2295,In_1510);
or U874 (N_874,In_1809,In_1590);
or U875 (N_875,In_706,In_2014);
xor U876 (N_876,In_617,In_2435);
and U877 (N_877,In_260,In_1487);
and U878 (N_878,In_867,In_292);
and U879 (N_879,In_1358,In_1366);
xor U880 (N_880,In_703,In_161);
xor U881 (N_881,In_2234,In_1792);
and U882 (N_882,In_232,In_149);
or U883 (N_883,In_1028,In_2152);
nand U884 (N_884,In_684,In_1956);
or U885 (N_885,In_1884,In_1632);
nand U886 (N_886,In_1561,In_2276);
nor U887 (N_887,In_758,In_1966);
nand U888 (N_888,In_2074,In_2098);
nand U889 (N_889,In_1402,In_957);
and U890 (N_890,In_2022,In_1617);
or U891 (N_891,In_2224,In_1823);
or U892 (N_892,In_39,In_634);
nand U893 (N_893,In_2170,In_898);
nand U894 (N_894,In_653,In_1164);
xnor U895 (N_895,In_213,In_896);
and U896 (N_896,In_968,In_322);
or U897 (N_897,In_1204,In_2177);
nor U898 (N_898,In_162,In_2084);
or U899 (N_899,In_1421,In_1805);
nor U900 (N_900,In_2095,In_908);
nand U901 (N_901,In_1917,In_1010);
xnor U902 (N_902,In_1596,In_2408);
and U903 (N_903,In_638,In_1964);
nor U904 (N_904,In_566,In_1781);
nor U905 (N_905,In_2300,In_1978);
xor U906 (N_906,In_1614,In_832);
or U907 (N_907,In_2223,In_1197);
nor U908 (N_908,In_906,In_1628);
nand U909 (N_909,In_501,In_1304);
and U910 (N_910,In_504,In_1994);
nor U911 (N_911,In_1943,In_1657);
nand U912 (N_912,In_54,In_841);
or U913 (N_913,In_2215,In_2220);
nor U914 (N_914,In_534,In_2396);
nand U915 (N_915,In_587,In_1350);
and U916 (N_916,In_2438,In_353);
or U917 (N_917,In_455,In_626);
and U918 (N_918,In_863,In_789);
nand U919 (N_919,In_2362,In_107);
or U920 (N_920,In_1931,In_2048);
nor U921 (N_921,In_665,In_202);
xor U922 (N_922,In_1132,In_1196);
or U923 (N_923,In_971,In_579);
nand U924 (N_924,In_2415,In_513);
xor U925 (N_925,In_1225,In_2254);
nor U926 (N_926,In_1191,In_885);
nor U927 (N_927,In_1397,In_1807);
or U928 (N_928,In_1839,In_458);
or U929 (N_929,In_294,In_263);
or U930 (N_930,In_361,In_800);
nor U931 (N_931,In_381,In_1349);
or U932 (N_932,In_1210,In_567);
nand U933 (N_933,In_2294,In_2303);
and U934 (N_934,In_1684,In_2459);
and U935 (N_935,In_544,In_5);
nor U936 (N_936,In_517,In_2072);
xnor U937 (N_937,In_917,In_1691);
xor U938 (N_938,In_1604,In_379);
nor U939 (N_939,In_557,In_1374);
and U940 (N_940,In_384,In_1557);
nor U941 (N_941,In_257,In_1801);
nor U942 (N_942,In_1221,In_767);
and U943 (N_943,In_1636,In_1493);
xor U944 (N_944,In_688,In_1430);
xnor U945 (N_945,In_1863,In_116);
or U946 (N_946,In_2277,In_2073);
nor U947 (N_947,In_181,In_672);
or U948 (N_948,In_1698,In_1255);
and U949 (N_949,In_1076,In_340);
nor U950 (N_950,In_975,In_500);
xnor U951 (N_951,In_1724,In_1715);
and U952 (N_952,In_1793,In_2159);
and U953 (N_953,In_1016,In_2021);
nand U954 (N_954,In_301,In_2238);
xnor U955 (N_955,In_1938,In_1354);
xor U956 (N_956,In_1925,In_145);
and U957 (N_957,In_388,In_1431);
nand U958 (N_958,In_1704,In_2471);
nor U959 (N_959,In_1155,In_1141);
and U960 (N_960,In_2379,In_1992);
nand U961 (N_961,In_803,In_2296);
or U962 (N_962,In_106,In_1854);
or U963 (N_963,In_1089,In_2410);
xnor U964 (N_964,In_308,In_365);
or U965 (N_965,In_583,In_1758);
and U966 (N_966,In_1530,In_1916);
or U967 (N_967,In_258,In_1268);
nor U968 (N_968,In_636,In_1871);
and U969 (N_969,In_1523,In_2499);
nand U970 (N_970,In_1475,In_2228);
or U971 (N_971,In_1274,In_1079);
or U972 (N_972,In_1647,In_2292);
nand U973 (N_973,In_128,In_1464);
or U974 (N_974,In_616,In_640);
and U975 (N_975,In_838,In_211);
nand U976 (N_976,In_1014,In_593);
or U977 (N_977,In_2324,In_1409);
or U978 (N_978,In_2226,In_2322);
nor U979 (N_979,In_2217,In_2185);
and U980 (N_980,In_532,In_882);
nand U981 (N_981,In_223,In_1219);
nor U982 (N_982,In_2066,In_2302);
xor U983 (N_983,In_1449,In_695);
xnor U984 (N_984,In_2080,In_1273);
xnor U985 (N_985,In_1143,In_374);
or U986 (N_986,In_2160,In_1395);
nand U987 (N_987,In_1735,In_1622);
or U988 (N_988,In_1481,In_2404);
nor U989 (N_989,In_1799,In_1180);
nor U990 (N_990,In_420,In_2352);
or U991 (N_991,In_2089,In_2477);
and U992 (N_992,In_1144,In_723);
nand U993 (N_993,In_228,In_41);
nand U994 (N_994,In_143,In_2288);
xnor U995 (N_995,In_1959,In_329);
or U996 (N_996,In_182,In_2443);
nand U997 (N_997,In_597,In_466);
and U998 (N_998,In_218,In_1811);
nand U999 (N_999,In_1860,In_2131);
xor U1000 (N_1000,In_668,In_1040);
nand U1001 (N_1001,In_977,In_726);
xnor U1002 (N_1002,In_315,In_1119);
and U1003 (N_1003,In_937,In_1013);
xnor U1004 (N_1004,In_2190,In_1276);
and U1005 (N_1005,In_884,In_741);
nand U1006 (N_1006,In_2076,In_704);
nor U1007 (N_1007,In_1965,In_505);
or U1008 (N_1008,In_2197,In_2042);
or U1009 (N_1009,In_2309,In_3);
xor U1010 (N_1010,In_693,In_2489);
nor U1011 (N_1011,In_1092,In_1001);
and U1012 (N_1012,In_127,In_656);
and U1013 (N_1013,In_265,In_651);
or U1014 (N_1014,In_710,In_1784);
nand U1015 (N_1015,In_973,In_1036);
xnor U1016 (N_1016,In_1154,In_1739);
and U1017 (N_1017,In_132,In_1867);
nand U1018 (N_1018,In_1721,In_2430);
nor U1019 (N_1019,In_622,In_2105);
nand U1020 (N_1020,In_1199,In_1816);
and U1021 (N_1021,In_226,In_168);
nor U1022 (N_1022,In_1103,In_1078);
xor U1023 (N_1023,In_2478,In_214);
or U1024 (N_1024,In_1520,In_409);
nor U1025 (N_1025,In_2225,In_1477);
or U1026 (N_1026,In_865,In_2100);
xnor U1027 (N_1027,In_1514,In_2342);
and U1028 (N_1028,In_969,In_2148);
nor U1029 (N_1029,In_235,In_1376);
and U1030 (N_1030,In_1192,In_1474);
nand U1031 (N_1031,In_151,In_721);
or U1032 (N_1032,In_1955,In_1969);
nand U1033 (N_1033,In_1110,In_635);
and U1034 (N_1034,In_852,In_225);
nor U1035 (N_1035,In_1166,In_2163);
nor U1036 (N_1036,In_1332,In_1208);
nand U1037 (N_1037,In_1546,In_679);
or U1038 (N_1038,In_1181,In_2335);
nor U1039 (N_1039,In_1836,In_1894);
or U1040 (N_1040,In_1538,In_2114);
and U1041 (N_1041,In_2268,In_1127);
or U1042 (N_1042,In_2350,In_1280);
or U1043 (N_1043,In_413,In_2096);
nand U1044 (N_1044,In_2403,In_811);
or U1045 (N_1045,In_219,In_2216);
nor U1046 (N_1046,In_1051,In_2377);
nand U1047 (N_1047,In_657,In_1578);
nand U1048 (N_1048,In_2206,In_682);
xnor U1049 (N_1049,In_755,In_1584);
nor U1050 (N_1050,In_1770,In_1364);
nor U1051 (N_1051,In_2082,In_686);
nand U1052 (N_1052,In_1712,In_1566);
or U1053 (N_1053,In_357,In_1303);
xor U1054 (N_1054,In_1087,In_1027);
nand U1055 (N_1055,In_2247,In_1135);
nand U1056 (N_1056,In_1971,In_1826);
and U1057 (N_1057,In_1246,In_669);
nand U1058 (N_1058,In_2194,In_254);
xnor U1059 (N_1059,In_243,In_2401);
nor U1060 (N_1060,In_246,In_742);
or U1061 (N_1061,In_2091,In_2490);
and U1062 (N_1062,In_572,In_135);
or U1063 (N_1063,In_554,In_2107);
and U1064 (N_1064,In_833,In_217);
xnor U1065 (N_1065,In_1291,In_391);
nand U1066 (N_1066,In_791,In_1230);
or U1067 (N_1067,In_1047,In_147);
xor U1068 (N_1068,In_1097,In_2279);
nor U1069 (N_1069,In_1545,In_828);
and U1070 (N_1070,In_1205,In_2487);
or U1071 (N_1071,In_456,In_1727);
and U1072 (N_1072,In_262,In_170);
nor U1073 (N_1073,In_398,In_788);
or U1074 (N_1074,In_2077,In_2442);
nand U1075 (N_1075,In_461,In_1746);
nand U1076 (N_1076,In_1398,In_1581);
or U1077 (N_1077,In_238,In_1085);
or U1078 (N_1078,In_925,In_980);
xor U1079 (N_1079,In_273,In_115);
or U1080 (N_1080,In_2260,In_400);
or U1081 (N_1081,In_1380,In_793);
nand U1082 (N_1082,In_1688,In_556);
xnor U1083 (N_1083,In_1544,In_2446);
nand U1084 (N_1084,In_279,In_2090);
nand U1085 (N_1085,In_34,In_2141);
and U1086 (N_1086,In_861,In_1408);
nor U1087 (N_1087,In_2037,In_1026);
or U1088 (N_1088,In_100,In_377);
or U1089 (N_1089,In_1990,In_921);
or U1090 (N_1090,In_177,In_2331);
and U1091 (N_1091,In_112,In_1005);
nand U1092 (N_1092,In_338,In_2355);
nor U1093 (N_1093,In_2166,In_595);
xnor U1094 (N_1094,In_142,In_1284);
and U1095 (N_1095,In_552,In_2494);
nor U1096 (N_1096,In_1748,In_1378);
xor U1097 (N_1097,In_2423,In_1939);
xor U1098 (N_1098,In_1672,In_1330);
and U1099 (N_1099,In_536,In_1716);
or U1100 (N_1100,In_470,In_1277);
and U1101 (N_1101,In_770,In_600);
or U1102 (N_1102,In_1249,In_1872);
nor U1103 (N_1103,In_2341,In_2387);
nor U1104 (N_1104,In_608,In_2371);
and U1105 (N_1105,In_2375,In_1343);
xor U1106 (N_1106,In_965,In_2336);
and U1107 (N_1107,In_1981,In_701);
nand U1108 (N_1108,In_923,In_233);
xnor U1109 (N_1109,In_2151,In_390);
or U1110 (N_1110,In_1693,In_1179);
or U1111 (N_1111,In_256,In_509);
and U1112 (N_1112,In_2092,In_2136);
and U1113 (N_1113,In_2308,In_2132);
nand U1114 (N_1114,In_2345,In_999);
nand U1115 (N_1115,In_660,In_997);
or U1116 (N_1116,In_1057,In_6);
xor U1117 (N_1117,In_1120,In_1522);
nand U1118 (N_1118,In_65,In_1373);
and U1119 (N_1119,In_2347,In_1218);
or U1120 (N_1120,In_1189,In_1968);
nor U1121 (N_1121,In_1212,In_2046);
xor U1122 (N_1122,In_2419,In_1942);
nand U1123 (N_1123,In_825,In_216);
nor U1124 (N_1124,In_1462,In_40);
xnor U1125 (N_1125,In_2450,In_988);
or U1126 (N_1126,In_1732,In_309);
xor U1127 (N_1127,In_1743,In_1471);
nor U1128 (N_1128,In_1214,In_324);
or U1129 (N_1129,In_894,In_1660);
xnor U1130 (N_1130,In_440,In_462);
or U1131 (N_1131,In_2290,In_1175);
or U1132 (N_1132,In_1592,In_1813);
nand U1133 (N_1133,In_156,In_402);
xor U1134 (N_1134,In_993,In_1266);
and U1135 (N_1135,In_1410,In_1685);
xor U1136 (N_1136,In_912,In_2061);
nand U1137 (N_1137,In_920,In_813);
and U1138 (N_1138,In_369,In_1242);
nand U1139 (N_1139,In_2174,In_807);
nor U1140 (N_1140,In_1153,In_111);
and U1141 (N_1141,In_1200,In_802);
or U1142 (N_1142,In_1853,In_2397);
xor U1143 (N_1143,In_166,In_1850);
and U1144 (N_1144,In_2402,In_2161);
or U1145 (N_1145,In_1002,In_274);
xnor U1146 (N_1146,In_2325,In_1405);
xnor U1147 (N_1147,In_1387,In_609);
nand U1148 (N_1148,In_2458,In_167);
or U1149 (N_1149,In_2269,In_1299);
nor U1150 (N_1150,In_2391,In_1776);
nor U1151 (N_1151,In_715,In_2332);
nor U1152 (N_1152,In_1442,In_559);
and U1153 (N_1153,In_250,In_2012);
nand U1154 (N_1154,In_1460,In_1866);
xnor U1155 (N_1155,In_1122,In_1259);
nor U1156 (N_1156,In_2333,In_350);
or U1157 (N_1157,In_77,In_1419);
xor U1158 (N_1158,In_1619,In_809);
xnor U1159 (N_1159,In_278,In_586);
and U1160 (N_1160,In_853,In_356);
xnor U1161 (N_1161,In_2140,In_1665);
and U1162 (N_1162,In_571,In_1941);
and U1163 (N_1163,In_874,In_2482);
nand U1164 (N_1164,In_495,In_2363);
or U1165 (N_1165,In_2209,In_1682);
and U1166 (N_1166,In_834,In_2462);
or U1167 (N_1167,In_280,In_707);
xor U1168 (N_1168,In_725,In_782);
xor U1169 (N_1169,In_450,In_2171);
or U1170 (N_1170,In_328,In_2109);
or U1171 (N_1171,In_2143,In_1668);
or U1172 (N_1172,In_792,In_2184);
xor U1173 (N_1173,In_1901,In_1988);
xor U1174 (N_1174,In_899,In_1723);
or U1175 (N_1175,In_2376,In_831);
and U1176 (N_1176,In_1215,In_222);
or U1177 (N_1177,In_2207,In_1282);
nand U1178 (N_1178,In_737,In_2367);
xnor U1179 (N_1179,In_1626,In_1936);
or U1180 (N_1180,In_1765,In_2056);
nand U1181 (N_1181,In_1157,In_516);
or U1182 (N_1182,In_1313,In_430);
nor U1183 (N_1183,In_2150,In_367);
nand U1184 (N_1184,In_1126,In_1593);
nand U1185 (N_1185,In_97,In_1422);
or U1186 (N_1186,In_1676,In_266);
nand U1187 (N_1187,In_558,In_1651);
nand U1188 (N_1188,In_1146,In_1247);
nand U1189 (N_1189,In_839,In_1609);
and U1190 (N_1190,In_2133,In_1237);
xnor U1191 (N_1191,In_2386,In_822);
xor U1192 (N_1192,In_2128,In_66);
nor U1193 (N_1193,In_511,In_146);
xnor U1194 (N_1194,In_439,In_94);
nand U1195 (N_1195,In_1458,In_1150);
and U1196 (N_1196,In_945,In_652);
or U1197 (N_1197,In_529,In_131);
or U1198 (N_1198,In_2432,In_137);
and U1199 (N_1199,In_493,In_1326);
nand U1200 (N_1200,In_2245,In_641);
nor U1201 (N_1201,In_815,In_2031);
nor U1202 (N_1202,In_2340,In_2032);
xnor U1203 (N_1203,In_1059,In_2451);
xnor U1204 (N_1204,In_2380,In_1738);
nand U1205 (N_1205,In_1645,In_590);
nor U1206 (N_1206,In_929,In_702);
xor U1207 (N_1207,In_866,In_2354);
or U1208 (N_1208,In_125,In_615);
xnor U1209 (N_1209,In_2440,In_1416);
or U1210 (N_1210,In_1289,In_790);
xor U1211 (N_1211,In_1294,In_452);
xnor U1212 (N_1212,In_2104,In_1841);
nand U1213 (N_1213,In_1168,In_186);
or U1214 (N_1214,In_1984,In_1382);
and U1215 (N_1215,In_1613,In_967);
or U1216 (N_1216,In_296,In_429);
or U1217 (N_1217,In_1678,In_1385);
nor U1218 (N_1218,In_57,In_2167);
nand U1219 (N_1219,In_13,In_1607);
xnor U1220 (N_1220,In_433,In_1142);
nor U1221 (N_1221,In_84,In_2416);
nor U1222 (N_1222,In_561,In_681);
nor U1223 (N_1223,In_1109,In_376);
nor U1224 (N_1224,In_868,In_319);
or U1225 (N_1225,In_690,In_680);
and U1226 (N_1226,In_1620,In_1468);
or U1227 (N_1227,In_1491,In_1031);
or U1228 (N_1228,In_691,In_1773);
xor U1229 (N_1229,In_1730,In_394);
nor U1230 (N_1230,In_2187,In_1568);
xnor U1231 (N_1231,In_1777,In_901);
nor U1232 (N_1232,In_1824,In_677);
nand U1233 (N_1233,In_1413,In_2015);
and U1234 (N_1234,In_729,In_1499);
or U1235 (N_1235,In_1940,In_1889);
or U1236 (N_1236,In_1998,In_730);
and U1237 (N_1237,In_134,In_449);
and U1238 (N_1238,In_32,In_2004);
or U1239 (N_1239,In_1172,In_1905);
xor U1240 (N_1240,In_856,In_335);
and U1241 (N_1241,In_804,In_1876);
or U1242 (N_1242,In_979,In_548);
nor U1243 (N_1243,In_592,In_2337);
or U1244 (N_1244,In_1484,In_575);
xnor U1245 (N_1245,In_1018,In_1797);
or U1246 (N_1246,In_1003,In_2205);
nand U1247 (N_1247,In_1139,In_2085);
and U1248 (N_1248,In_96,In_1760);
xor U1249 (N_1249,In_893,In_1052);
and U1250 (N_1250,In_2448,In_459);
xor U1251 (N_1251,In_135,In_498);
nand U1252 (N_1252,In_179,In_128);
nor U1253 (N_1253,In_134,In_372);
xor U1254 (N_1254,In_1651,In_556);
nor U1255 (N_1255,In_214,In_1619);
xnor U1256 (N_1256,In_1177,In_123);
xnor U1257 (N_1257,In_1502,In_105);
or U1258 (N_1258,In_1447,In_105);
and U1259 (N_1259,In_1368,In_1601);
or U1260 (N_1260,In_2271,In_2449);
nor U1261 (N_1261,In_1467,In_2195);
xor U1262 (N_1262,In_2102,In_1106);
nand U1263 (N_1263,In_1042,In_876);
and U1264 (N_1264,In_25,In_2165);
nor U1265 (N_1265,In_2083,In_553);
xnor U1266 (N_1266,In_2407,In_1914);
or U1267 (N_1267,In_812,In_59);
nand U1268 (N_1268,In_176,In_195);
and U1269 (N_1269,In_1696,In_31);
nand U1270 (N_1270,In_1988,In_261);
or U1271 (N_1271,In_261,In_2198);
or U1272 (N_1272,In_685,In_1958);
nor U1273 (N_1273,In_2018,In_2093);
nor U1274 (N_1274,In_295,In_2299);
or U1275 (N_1275,In_606,In_2367);
or U1276 (N_1276,In_1699,In_2462);
or U1277 (N_1277,In_1138,In_1811);
and U1278 (N_1278,In_1020,In_1547);
xnor U1279 (N_1279,In_482,In_92);
nor U1280 (N_1280,In_1156,In_2297);
xnor U1281 (N_1281,In_2430,In_2261);
nand U1282 (N_1282,In_990,In_684);
or U1283 (N_1283,In_1476,In_654);
xnor U1284 (N_1284,In_734,In_1669);
or U1285 (N_1285,In_61,In_1959);
xnor U1286 (N_1286,In_36,In_217);
or U1287 (N_1287,In_2208,In_1137);
and U1288 (N_1288,In_1180,In_1731);
nand U1289 (N_1289,In_2068,In_1096);
xnor U1290 (N_1290,In_1883,In_236);
and U1291 (N_1291,In_1963,In_752);
and U1292 (N_1292,In_548,In_579);
xnor U1293 (N_1293,In_2439,In_1902);
nor U1294 (N_1294,In_780,In_1117);
and U1295 (N_1295,In_1110,In_190);
nand U1296 (N_1296,In_906,In_2184);
xor U1297 (N_1297,In_527,In_1391);
or U1298 (N_1298,In_1460,In_946);
or U1299 (N_1299,In_717,In_2158);
nand U1300 (N_1300,In_1936,In_588);
nand U1301 (N_1301,In_1117,In_2266);
xnor U1302 (N_1302,In_2309,In_916);
or U1303 (N_1303,In_1532,In_2216);
nor U1304 (N_1304,In_1610,In_1362);
nand U1305 (N_1305,In_432,In_1951);
xor U1306 (N_1306,In_1672,In_1592);
xor U1307 (N_1307,In_2244,In_145);
xnor U1308 (N_1308,In_376,In_855);
or U1309 (N_1309,In_912,In_216);
nor U1310 (N_1310,In_1402,In_2281);
nor U1311 (N_1311,In_717,In_754);
xnor U1312 (N_1312,In_773,In_29);
or U1313 (N_1313,In_1396,In_1154);
or U1314 (N_1314,In_641,In_2073);
nand U1315 (N_1315,In_459,In_1947);
nor U1316 (N_1316,In_648,In_1385);
nand U1317 (N_1317,In_1567,In_2469);
or U1318 (N_1318,In_2386,In_313);
nand U1319 (N_1319,In_387,In_2420);
and U1320 (N_1320,In_1041,In_1119);
nand U1321 (N_1321,In_162,In_1613);
or U1322 (N_1322,In_926,In_1942);
and U1323 (N_1323,In_221,In_1166);
nor U1324 (N_1324,In_2310,In_1455);
nor U1325 (N_1325,In_2301,In_899);
nor U1326 (N_1326,In_1593,In_63);
nand U1327 (N_1327,In_1629,In_2374);
or U1328 (N_1328,In_159,In_1347);
or U1329 (N_1329,In_440,In_121);
nor U1330 (N_1330,In_793,In_2202);
nor U1331 (N_1331,In_1103,In_683);
xnor U1332 (N_1332,In_2255,In_1030);
or U1333 (N_1333,In_861,In_1366);
and U1334 (N_1334,In_1712,In_1124);
xor U1335 (N_1335,In_210,In_769);
nor U1336 (N_1336,In_357,In_1016);
nor U1337 (N_1337,In_806,In_1111);
xor U1338 (N_1338,In_2494,In_1772);
xor U1339 (N_1339,In_1087,In_530);
nor U1340 (N_1340,In_2091,In_393);
and U1341 (N_1341,In_33,In_1945);
or U1342 (N_1342,In_1469,In_2362);
or U1343 (N_1343,In_2212,In_28);
xor U1344 (N_1344,In_1555,In_1176);
nor U1345 (N_1345,In_1223,In_1052);
or U1346 (N_1346,In_1607,In_145);
and U1347 (N_1347,In_455,In_2203);
nor U1348 (N_1348,In_595,In_343);
xnor U1349 (N_1349,In_1854,In_2058);
nor U1350 (N_1350,In_1630,In_1049);
nor U1351 (N_1351,In_2076,In_1830);
or U1352 (N_1352,In_549,In_1796);
and U1353 (N_1353,In_2442,In_2071);
nor U1354 (N_1354,In_1794,In_2193);
and U1355 (N_1355,In_866,In_1813);
or U1356 (N_1356,In_2173,In_252);
nand U1357 (N_1357,In_1304,In_1777);
nand U1358 (N_1358,In_1974,In_2356);
and U1359 (N_1359,In_2253,In_1207);
nand U1360 (N_1360,In_1467,In_1406);
and U1361 (N_1361,In_2197,In_2214);
and U1362 (N_1362,In_1035,In_1155);
nor U1363 (N_1363,In_1064,In_714);
and U1364 (N_1364,In_775,In_2390);
and U1365 (N_1365,In_1238,In_1641);
and U1366 (N_1366,In_64,In_320);
xnor U1367 (N_1367,In_61,In_2462);
xor U1368 (N_1368,In_2422,In_690);
nor U1369 (N_1369,In_2186,In_1625);
and U1370 (N_1370,In_1369,In_607);
nand U1371 (N_1371,In_1782,In_2040);
nand U1372 (N_1372,In_1241,In_1415);
or U1373 (N_1373,In_2316,In_612);
or U1374 (N_1374,In_1279,In_2329);
nand U1375 (N_1375,In_2054,In_1740);
and U1376 (N_1376,In_1369,In_1136);
nand U1377 (N_1377,In_1868,In_355);
nor U1378 (N_1378,In_978,In_1715);
xor U1379 (N_1379,In_1052,In_59);
nor U1380 (N_1380,In_1198,In_2269);
nor U1381 (N_1381,In_152,In_1936);
nor U1382 (N_1382,In_470,In_2484);
xnor U1383 (N_1383,In_908,In_2183);
and U1384 (N_1384,In_1755,In_1636);
nor U1385 (N_1385,In_923,In_254);
nand U1386 (N_1386,In_2329,In_1385);
or U1387 (N_1387,In_2358,In_2109);
xor U1388 (N_1388,In_24,In_2011);
and U1389 (N_1389,In_584,In_623);
nand U1390 (N_1390,In_487,In_2415);
and U1391 (N_1391,In_685,In_784);
xor U1392 (N_1392,In_1603,In_693);
nor U1393 (N_1393,In_257,In_740);
nand U1394 (N_1394,In_1824,In_1810);
xnor U1395 (N_1395,In_2366,In_1319);
or U1396 (N_1396,In_1361,In_2360);
nor U1397 (N_1397,In_2300,In_725);
nor U1398 (N_1398,In_631,In_157);
nor U1399 (N_1399,In_713,In_2059);
or U1400 (N_1400,In_2428,In_1550);
nor U1401 (N_1401,In_1276,In_224);
nor U1402 (N_1402,In_1154,In_1409);
and U1403 (N_1403,In_852,In_1149);
xor U1404 (N_1404,In_1590,In_2252);
or U1405 (N_1405,In_1149,In_600);
nand U1406 (N_1406,In_2377,In_121);
or U1407 (N_1407,In_819,In_2348);
xnor U1408 (N_1408,In_1856,In_675);
nor U1409 (N_1409,In_1203,In_96);
and U1410 (N_1410,In_1523,In_462);
nor U1411 (N_1411,In_1579,In_808);
xor U1412 (N_1412,In_832,In_1340);
nor U1413 (N_1413,In_1994,In_116);
or U1414 (N_1414,In_327,In_2282);
and U1415 (N_1415,In_369,In_177);
or U1416 (N_1416,In_2452,In_474);
xnor U1417 (N_1417,In_732,In_1174);
and U1418 (N_1418,In_842,In_1800);
nand U1419 (N_1419,In_2359,In_1247);
or U1420 (N_1420,In_1512,In_1375);
and U1421 (N_1421,In_651,In_2248);
nand U1422 (N_1422,In_2318,In_787);
or U1423 (N_1423,In_1023,In_1582);
xnor U1424 (N_1424,In_1602,In_307);
or U1425 (N_1425,In_1719,In_1713);
nor U1426 (N_1426,In_1786,In_545);
xnor U1427 (N_1427,In_1867,In_315);
xor U1428 (N_1428,In_2069,In_2233);
nor U1429 (N_1429,In_1940,In_1898);
or U1430 (N_1430,In_2363,In_850);
and U1431 (N_1431,In_153,In_725);
and U1432 (N_1432,In_628,In_383);
xor U1433 (N_1433,In_314,In_2217);
nor U1434 (N_1434,In_480,In_1763);
nand U1435 (N_1435,In_1061,In_904);
and U1436 (N_1436,In_1118,In_1659);
and U1437 (N_1437,In_2218,In_2027);
and U1438 (N_1438,In_1147,In_333);
or U1439 (N_1439,In_1524,In_1337);
nor U1440 (N_1440,In_522,In_1826);
or U1441 (N_1441,In_1164,In_282);
and U1442 (N_1442,In_1736,In_1686);
nor U1443 (N_1443,In_1402,In_1753);
xnor U1444 (N_1444,In_842,In_185);
nor U1445 (N_1445,In_2094,In_1666);
and U1446 (N_1446,In_384,In_1586);
and U1447 (N_1447,In_1147,In_285);
xnor U1448 (N_1448,In_1612,In_1337);
and U1449 (N_1449,In_243,In_29);
nor U1450 (N_1450,In_1613,In_1852);
xnor U1451 (N_1451,In_2129,In_439);
nand U1452 (N_1452,In_875,In_1183);
nor U1453 (N_1453,In_495,In_2420);
nand U1454 (N_1454,In_1885,In_272);
nor U1455 (N_1455,In_1019,In_324);
and U1456 (N_1456,In_1823,In_1952);
nand U1457 (N_1457,In_546,In_1499);
and U1458 (N_1458,In_1774,In_1167);
nor U1459 (N_1459,In_972,In_533);
or U1460 (N_1460,In_1485,In_771);
nand U1461 (N_1461,In_51,In_2092);
or U1462 (N_1462,In_408,In_460);
xor U1463 (N_1463,In_1205,In_212);
nand U1464 (N_1464,In_1610,In_1910);
or U1465 (N_1465,In_297,In_278);
and U1466 (N_1466,In_1116,In_2232);
nand U1467 (N_1467,In_616,In_2386);
or U1468 (N_1468,In_2365,In_1448);
or U1469 (N_1469,In_1520,In_582);
or U1470 (N_1470,In_669,In_1933);
xnor U1471 (N_1471,In_367,In_1900);
nand U1472 (N_1472,In_1935,In_1097);
nor U1473 (N_1473,In_1539,In_411);
nor U1474 (N_1474,In_569,In_1226);
and U1475 (N_1475,In_1980,In_2199);
nor U1476 (N_1476,In_1842,In_2242);
nand U1477 (N_1477,In_2322,In_689);
and U1478 (N_1478,In_590,In_1990);
nor U1479 (N_1479,In_1400,In_1197);
xor U1480 (N_1480,In_2336,In_2382);
nor U1481 (N_1481,In_827,In_2257);
nor U1482 (N_1482,In_928,In_2123);
and U1483 (N_1483,In_1693,In_2407);
nor U1484 (N_1484,In_1031,In_1133);
nand U1485 (N_1485,In_2190,In_806);
and U1486 (N_1486,In_775,In_261);
or U1487 (N_1487,In_921,In_1658);
or U1488 (N_1488,In_2381,In_2400);
and U1489 (N_1489,In_2127,In_1081);
and U1490 (N_1490,In_1,In_2439);
nor U1491 (N_1491,In_42,In_745);
nor U1492 (N_1492,In_815,In_65);
nor U1493 (N_1493,In_2347,In_2091);
nor U1494 (N_1494,In_853,In_1161);
xnor U1495 (N_1495,In_414,In_2245);
and U1496 (N_1496,In_1635,In_1398);
nor U1497 (N_1497,In_2338,In_841);
xor U1498 (N_1498,In_2386,In_1904);
or U1499 (N_1499,In_1081,In_1306);
and U1500 (N_1500,In_237,In_215);
and U1501 (N_1501,In_2152,In_1472);
and U1502 (N_1502,In_48,In_848);
and U1503 (N_1503,In_2189,In_2196);
xor U1504 (N_1504,In_2152,In_1494);
nor U1505 (N_1505,In_924,In_313);
or U1506 (N_1506,In_410,In_668);
or U1507 (N_1507,In_990,In_776);
or U1508 (N_1508,In_2347,In_763);
or U1509 (N_1509,In_186,In_1949);
nand U1510 (N_1510,In_2483,In_2333);
nor U1511 (N_1511,In_1439,In_2270);
and U1512 (N_1512,In_543,In_2239);
xor U1513 (N_1513,In_2363,In_769);
and U1514 (N_1514,In_1804,In_1587);
xnor U1515 (N_1515,In_1585,In_1154);
nor U1516 (N_1516,In_1362,In_2452);
xnor U1517 (N_1517,In_1544,In_521);
nand U1518 (N_1518,In_2054,In_2496);
and U1519 (N_1519,In_2375,In_1244);
xnor U1520 (N_1520,In_213,In_2194);
and U1521 (N_1521,In_1336,In_1297);
nand U1522 (N_1522,In_576,In_1085);
and U1523 (N_1523,In_1153,In_1320);
xnor U1524 (N_1524,In_1673,In_788);
and U1525 (N_1525,In_256,In_737);
nor U1526 (N_1526,In_1443,In_2265);
or U1527 (N_1527,In_391,In_1576);
and U1528 (N_1528,In_1021,In_1739);
nand U1529 (N_1529,In_1682,In_879);
or U1530 (N_1530,In_1129,In_2348);
nor U1531 (N_1531,In_1125,In_1630);
nor U1532 (N_1532,In_908,In_2174);
nor U1533 (N_1533,In_1727,In_114);
and U1534 (N_1534,In_2469,In_1729);
nand U1535 (N_1535,In_1084,In_45);
and U1536 (N_1536,In_1728,In_2217);
nand U1537 (N_1537,In_550,In_359);
or U1538 (N_1538,In_1412,In_2034);
and U1539 (N_1539,In_798,In_432);
nand U1540 (N_1540,In_1228,In_703);
xnor U1541 (N_1541,In_122,In_1120);
xnor U1542 (N_1542,In_2145,In_826);
xor U1543 (N_1543,In_994,In_1489);
xnor U1544 (N_1544,In_2348,In_2236);
and U1545 (N_1545,In_1781,In_1712);
and U1546 (N_1546,In_410,In_291);
nand U1547 (N_1547,In_1675,In_1097);
nor U1548 (N_1548,In_77,In_1863);
and U1549 (N_1549,In_1542,In_309);
nor U1550 (N_1550,In_590,In_2281);
nand U1551 (N_1551,In_2496,In_343);
nand U1552 (N_1552,In_546,In_368);
or U1553 (N_1553,In_1245,In_1766);
and U1554 (N_1554,In_1860,In_1769);
xor U1555 (N_1555,In_1327,In_45);
nor U1556 (N_1556,In_1421,In_204);
nor U1557 (N_1557,In_864,In_2168);
nand U1558 (N_1558,In_1822,In_486);
nand U1559 (N_1559,In_377,In_1681);
xor U1560 (N_1560,In_2017,In_1992);
nor U1561 (N_1561,In_310,In_1429);
nor U1562 (N_1562,In_1873,In_6);
nor U1563 (N_1563,In_1428,In_420);
or U1564 (N_1564,In_172,In_647);
nand U1565 (N_1565,In_1978,In_2183);
or U1566 (N_1566,In_587,In_643);
or U1567 (N_1567,In_174,In_1235);
or U1568 (N_1568,In_814,In_189);
nor U1569 (N_1569,In_847,In_274);
xor U1570 (N_1570,In_1662,In_1429);
and U1571 (N_1571,In_250,In_1092);
and U1572 (N_1572,In_527,In_140);
and U1573 (N_1573,In_1141,In_1361);
or U1574 (N_1574,In_979,In_98);
nor U1575 (N_1575,In_1298,In_352);
nor U1576 (N_1576,In_2437,In_336);
or U1577 (N_1577,In_957,In_778);
and U1578 (N_1578,In_2283,In_1472);
xnor U1579 (N_1579,In_249,In_192);
xnor U1580 (N_1580,In_290,In_1356);
or U1581 (N_1581,In_1565,In_1721);
or U1582 (N_1582,In_2071,In_2298);
or U1583 (N_1583,In_2031,In_958);
and U1584 (N_1584,In_2185,In_1215);
nand U1585 (N_1585,In_2326,In_2392);
xnor U1586 (N_1586,In_2270,In_1404);
nand U1587 (N_1587,In_443,In_831);
and U1588 (N_1588,In_1197,In_661);
nand U1589 (N_1589,In_211,In_1941);
or U1590 (N_1590,In_95,In_1594);
nor U1591 (N_1591,In_1061,In_1663);
xnor U1592 (N_1592,In_2418,In_829);
xor U1593 (N_1593,In_1351,In_137);
xnor U1594 (N_1594,In_2493,In_742);
nand U1595 (N_1595,In_867,In_1612);
nor U1596 (N_1596,In_1322,In_824);
nor U1597 (N_1597,In_830,In_1134);
or U1598 (N_1598,In_1904,In_1963);
nand U1599 (N_1599,In_250,In_1856);
nand U1600 (N_1600,In_1835,In_237);
or U1601 (N_1601,In_2304,In_1546);
xor U1602 (N_1602,In_1151,In_1821);
or U1603 (N_1603,In_1248,In_850);
nor U1604 (N_1604,In_1980,In_2397);
nor U1605 (N_1605,In_2007,In_993);
xor U1606 (N_1606,In_778,In_1945);
and U1607 (N_1607,In_714,In_2364);
or U1608 (N_1608,In_1894,In_594);
xor U1609 (N_1609,In_981,In_1008);
and U1610 (N_1610,In_1584,In_2374);
or U1611 (N_1611,In_265,In_2434);
and U1612 (N_1612,In_62,In_180);
nor U1613 (N_1613,In_1009,In_909);
nand U1614 (N_1614,In_1042,In_2344);
or U1615 (N_1615,In_442,In_1011);
or U1616 (N_1616,In_1240,In_2129);
xnor U1617 (N_1617,In_585,In_916);
xnor U1618 (N_1618,In_1234,In_107);
and U1619 (N_1619,In_2379,In_1787);
xor U1620 (N_1620,In_873,In_1102);
and U1621 (N_1621,In_454,In_1263);
xor U1622 (N_1622,In_615,In_92);
xnor U1623 (N_1623,In_589,In_610);
xor U1624 (N_1624,In_1003,In_998);
nor U1625 (N_1625,In_1246,In_1454);
xor U1626 (N_1626,In_2055,In_2206);
nor U1627 (N_1627,In_1936,In_634);
nor U1628 (N_1628,In_732,In_446);
or U1629 (N_1629,In_294,In_564);
and U1630 (N_1630,In_41,In_848);
nand U1631 (N_1631,In_747,In_727);
and U1632 (N_1632,In_1409,In_1310);
or U1633 (N_1633,In_306,In_475);
xor U1634 (N_1634,In_1909,In_446);
and U1635 (N_1635,In_1104,In_440);
xnor U1636 (N_1636,In_606,In_2005);
nand U1637 (N_1637,In_718,In_307);
nor U1638 (N_1638,In_850,In_1229);
nor U1639 (N_1639,In_624,In_1365);
or U1640 (N_1640,In_826,In_347);
nand U1641 (N_1641,In_774,In_1924);
nor U1642 (N_1642,In_1865,In_268);
xnor U1643 (N_1643,In_663,In_418);
nand U1644 (N_1644,In_414,In_1927);
xnor U1645 (N_1645,In_40,In_1844);
xnor U1646 (N_1646,In_1355,In_1017);
or U1647 (N_1647,In_1624,In_944);
nor U1648 (N_1648,In_2408,In_1086);
xnor U1649 (N_1649,In_1635,In_1263);
nand U1650 (N_1650,In_1285,In_928);
and U1651 (N_1651,In_869,In_2408);
nand U1652 (N_1652,In_2350,In_317);
or U1653 (N_1653,In_900,In_768);
or U1654 (N_1654,In_2185,In_863);
nand U1655 (N_1655,In_2009,In_179);
nand U1656 (N_1656,In_2388,In_1201);
nand U1657 (N_1657,In_1943,In_1557);
nand U1658 (N_1658,In_2382,In_205);
nor U1659 (N_1659,In_186,In_425);
nand U1660 (N_1660,In_2130,In_485);
and U1661 (N_1661,In_1476,In_190);
or U1662 (N_1662,In_1701,In_1721);
nand U1663 (N_1663,In_1764,In_2082);
or U1664 (N_1664,In_2292,In_2496);
or U1665 (N_1665,In_523,In_1874);
xnor U1666 (N_1666,In_2277,In_1111);
xnor U1667 (N_1667,In_2081,In_2389);
nor U1668 (N_1668,In_2461,In_878);
xnor U1669 (N_1669,In_1294,In_1113);
nor U1670 (N_1670,In_1895,In_2492);
nand U1671 (N_1671,In_263,In_1873);
or U1672 (N_1672,In_180,In_373);
xor U1673 (N_1673,In_1330,In_936);
nand U1674 (N_1674,In_1983,In_2296);
nand U1675 (N_1675,In_1583,In_1375);
nand U1676 (N_1676,In_999,In_1022);
or U1677 (N_1677,In_739,In_720);
nor U1678 (N_1678,In_382,In_54);
nor U1679 (N_1679,In_1987,In_1111);
nand U1680 (N_1680,In_1032,In_708);
nand U1681 (N_1681,In_479,In_25);
nor U1682 (N_1682,In_1608,In_1400);
nor U1683 (N_1683,In_1950,In_61);
xor U1684 (N_1684,In_1878,In_1250);
nor U1685 (N_1685,In_2272,In_1756);
and U1686 (N_1686,In_2380,In_1281);
nor U1687 (N_1687,In_1980,In_362);
nand U1688 (N_1688,In_1186,In_360);
nor U1689 (N_1689,In_709,In_1997);
or U1690 (N_1690,In_2109,In_2020);
and U1691 (N_1691,In_1181,In_2084);
nand U1692 (N_1692,In_1149,In_570);
xor U1693 (N_1693,In_1617,In_236);
xnor U1694 (N_1694,In_821,In_534);
xor U1695 (N_1695,In_104,In_418);
nor U1696 (N_1696,In_291,In_1764);
nand U1697 (N_1697,In_783,In_20);
and U1698 (N_1698,In_1491,In_2414);
xnor U1699 (N_1699,In_1590,In_1902);
nor U1700 (N_1700,In_2259,In_1786);
nor U1701 (N_1701,In_745,In_2447);
nor U1702 (N_1702,In_209,In_2070);
and U1703 (N_1703,In_816,In_833);
or U1704 (N_1704,In_1611,In_1657);
and U1705 (N_1705,In_2472,In_1469);
xor U1706 (N_1706,In_2470,In_424);
or U1707 (N_1707,In_205,In_627);
xnor U1708 (N_1708,In_1006,In_74);
xor U1709 (N_1709,In_586,In_1510);
xnor U1710 (N_1710,In_2311,In_535);
nand U1711 (N_1711,In_2492,In_1826);
nor U1712 (N_1712,In_464,In_1845);
nand U1713 (N_1713,In_1198,In_2221);
xor U1714 (N_1714,In_1233,In_18);
xnor U1715 (N_1715,In_2026,In_501);
or U1716 (N_1716,In_1566,In_1411);
nor U1717 (N_1717,In_239,In_531);
nor U1718 (N_1718,In_2064,In_1657);
and U1719 (N_1719,In_551,In_942);
nor U1720 (N_1720,In_2168,In_2492);
nand U1721 (N_1721,In_116,In_2034);
nand U1722 (N_1722,In_1297,In_1875);
xnor U1723 (N_1723,In_1595,In_936);
nor U1724 (N_1724,In_1185,In_2117);
and U1725 (N_1725,In_1307,In_105);
xor U1726 (N_1726,In_947,In_1499);
nand U1727 (N_1727,In_1782,In_1618);
nand U1728 (N_1728,In_537,In_1570);
or U1729 (N_1729,In_1207,In_983);
nand U1730 (N_1730,In_369,In_2359);
or U1731 (N_1731,In_1889,In_50);
or U1732 (N_1732,In_270,In_2185);
nand U1733 (N_1733,In_1414,In_2191);
or U1734 (N_1734,In_1262,In_767);
or U1735 (N_1735,In_898,In_895);
xor U1736 (N_1736,In_2353,In_1769);
or U1737 (N_1737,In_1963,In_1987);
nor U1738 (N_1738,In_1933,In_678);
xor U1739 (N_1739,In_1435,In_2315);
or U1740 (N_1740,In_330,In_263);
nand U1741 (N_1741,In_1775,In_2421);
nand U1742 (N_1742,In_2093,In_1388);
and U1743 (N_1743,In_354,In_1838);
or U1744 (N_1744,In_522,In_613);
nor U1745 (N_1745,In_73,In_1424);
or U1746 (N_1746,In_2068,In_1772);
nand U1747 (N_1747,In_141,In_1429);
nor U1748 (N_1748,In_126,In_473);
nand U1749 (N_1749,In_833,In_94);
and U1750 (N_1750,In_1502,In_1625);
nor U1751 (N_1751,In_350,In_459);
or U1752 (N_1752,In_541,In_1072);
and U1753 (N_1753,In_1789,In_615);
xnor U1754 (N_1754,In_595,In_2330);
xnor U1755 (N_1755,In_929,In_935);
and U1756 (N_1756,In_2334,In_1950);
nand U1757 (N_1757,In_1544,In_1453);
and U1758 (N_1758,In_1327,In_1827);
or U1759 (N_1759,In_2136,In_2362);
nor U1760 (N_1760,In_434,In_1271);
and U1761 (N_1761,In_485,In_2010);
and U1762 (N_1762,In_2204,In_1601);
or U1763 (N_1763,In_1958,In_2267);
or U1764 (N_1764,In_977,In_2069);
nor U1765 (N_1765,In_1747,In_2387);
or U1766 (N_1766,In_736,In_290);
or U1767 (N_1767,In_1365,In_498);
and U1768 (N_1768,In_2223,In_1669);
xor U1769 (N_1769,In_698,In_1197);
nor U1770 (N_1770,In_80,In_1509);
and U1771 (N_1771,In_1998,In_1364);
nand U1772 (N_1772,In_1521,In_723);
xor U1773 (N_1773,In_877,In_1342);
xor U1774 (N_1774,In_565,In_171);
and U1775 (N_1775,In_1082,In_104);
nor U1776 (N_1776,In_455,In_2289);
xor U1777 (N_1777,In_347,In_654);
xor U1778 (N_1778,In_527,In_1977);
nand U1779 (N_1779,In_1617,In_1403);
or U1780 (N_1780,In_1651,In_2282);
nor U1781 (N_1781,In_1796,In_1217);
nand U1782 (N_1782,In_1691,In_607);
or U1783 (N_1783,In_1547,In_538);
and U1784 (N_1784,In_1637,In_1742);
xnor U1785 (N_1785,In_1216,In_1091);
and U1786 (N_1786,In_2492,In_1621);
and U1787 (N_1787,In_2182,In_231);
nand U1788 (N_1788,In_1211,In_86);
or U1789 (N_1789,In_97,In_394);
xor U1790 (N_1790,In_1519,In_887);
nor U1791 (N_1791,In_1994,In_2183);
and U1792 (N_1792,In_1319,In_467);
and U1793 (N_1793,In_999,In_1336);
nor U1794 (N_1794,In_2433,In_1980);
nand U1795 (N_1795,In_825,In_1274);
nor U1796 (N_1796,In_851,In_72);
nand U1797 (N_1797,In_208,In_1195);
xor U1798 (N_1798,In_1479,In_1672);
and U1799 (N_1799,In_1726,In_1264);
xor U1800 (N_1800,In_2319,In_858);
nand U1801 (N_1801,In_1641,In_816);
xnor U1802 (N_1802,In_937,In_1582);
nand U1803 (N_1803,In_1650,In_2292);
nor U1804 (N_1804,In_465,In_1929);
or U1805 (N_1805,In_1857,In_540);
nand U1806 (N_1806,In_426,In_1374);
or U1807 (N_1807,In_937,In_1938);
xor U1808 (N_1808,In_177,In_1037);
xnor U1809 (N_1809,In_1566,In_1898);
nand U1810 (N_1810,In_514,In_46);
nand U1811 (N_1811,In_2445,In_1182);
and U1812 (N_1812,In_2301,In_626);
nand U1813 (N_1813,In_2190,In_187);
xnor U1814 (N_1814,In_928,In_1836);
nand U1815 (N_1815,In_2138,In_1731);
and U1816 (N_1816,In_309,In_1790);
nor U1817 (N_1817,In_2304,In_1005);
and U1818 (N_1818,In_2341,In_339);
or U1819 (N_1819,In_360,In_1958);
xnor U1820 (N_1820,In_2233,In_1421);
or U1821 (N_1821,In_2106,In_1887);
xnor U1822 (N_1822,In_733,In_1974);
xnor U1823 (N_1823,In_655,In_2335);
nor U1824 (N_1824,In_983,In_1579);
nor U1825 (N_1825,In_202,In_2175);
or U1826 (N_1826,In_1186,In_19);
or U1827 (N_1827,In_1067,In_576);
nor U1828 (N_1828,In_1092,In_1336);
or U1829 (N_1829,In_2413,In_1789);
nor U1830 (N_1830,In_2272,In_475);
and U1831 (N_1831,In_1222,In_1800);
xnor U1832 (N_1832,In_1504,In_2407);
nor U1833 (N_1833,In_617,In_926);
xnor U1834 (N_1834,In_2035,In_98);
or U1835 (N_1835,In_1730,In_1922);
nand U1836 (N_1836,In_394,In_1605);
and U1837 (N_1837,In_1937,In_2303);
nor U1838 (N_1838,In_1620,In_2150);
and U1839 (N_1839,In_212,In_1395);
nand U1840 (N_1840,In_233,In_382);
xor U1841 (N_1841,In_497,In_1777);
xor U1842 (N_1842,In_1,In_1673);
or U1843 (N_1843,In_182,In_311);
and U1844 (N_1844,In_2349,In_1339);
nand U1845 (N_1845,In_444,In_996);
xnor U1846 (N_1846,In_1943,In_1424);
xnor U1847 (N_1847,In_976,In_2347);
and U1848 (N_1848,In_2430,In_847);
or U1849 (N_1849,In_1829,In_1463);
or U1850 (N_1850,In_1950,In_424);
and U1851 (N_1851,In_1799,In_850);
xor U1852 (N_1852,In_1879,In_1349);
or U1853 (N_1853,In_410,In_1138);
or U1854 (N_1854,In_229,In_2013);
and U1855 (N_1855,In_1063,In_1671);
nand U1856 (N_1856,In_1347,In_2440);
and U1857 (N_1857,In_1534,In_958);
nand U1858 (N_1858,In_206,In_862);
nor U1859 (N_1859,In_2220,In_2393);
xor U1860 (N_1860,In_1973,In_2429);
xor U1861 (N_1861,In_775,In_712);
and U1862 (N_1862,In_1923,In_1029);
nand U1863 (N_1863,In_1315,In_981);
xnor U1864 (N_1864,In_885,In_1214);
nand U1865 (N_1865,In_519,In_1335);
or U1866 (N_1866,In_1601,In_1615);
nand U1867 (N_1867,In_2144,In_1487);
nor U1868 (N_1868,In_824,In_1251);
nand U1869 (N_1869,In_2444,In_1507);
nand U1870 (N_1870,In_2319,In_166);
or U1871 (N_1871,In_436,In_503);
xor U1872 (N_1872,In_1915,In_2473);
nor U1873 (N_1873,In_2164,In_323);
and U1874 (N_1874,In_421,In_910);
nand U1875 (N_1875,In_2417,In_958);
nor U1876 (N_1876,In_1829,In_1177);
nor U1877 (N_1877,In_83,In_1840);
nor U1878 (N_1878,In_1739,In_2290);
xor U1879 (N_1879,In_1627,In_401);
xnor U1880 (N_1880,In_1328,In_181);
nor U1881 (N_1881,In_1082,In_379);
or U1882 (N_1882,In_1149,In_1139);
nor U1883 (N_1883,In_383,In_1636);
and U1884 (N_1884,In_614,In_1154);
xnor U1885 (N_1885,In_2153,In_2420);
nand U1886 (N_1886,In_1545,In_1435);
and U1887 (N_1887,In_378,In_202);
or U1888 (N_1888,In_1744,In_2275);
xnor U1889 (N_1889,In_2396,In_1770);
xor U1890 (N_1890,In_1517,In_1494);
nor U1891 (N_1891,In_260,In_376);
nand U1892 (N_1892,In_2484,In_666);
or U1893 (N_1893,In_2201,In_1598);
or U1894 (N_1894,In_2257,In_1361);
nor U1895 (N_1895,In_1562,In_227);
nor U1896 (N_1896,In_102,In_2151);
xnor U1897 (N_1897,In_1908,In_2181);
xor U1898 (N_1898,In_863,In_1106);
nor U1899 (N_1899,In_2062,In_529);
or U1900 (N_1900,In_386,In_897);
nand U1901 (N_1901,In_1707,In_503);
nor U1902 (N_1902,In_796,In_66);
nor U1903 (N_1903,In_1909,In_629);
nand U1904 (N_1904,In_679,In_581);
and U1905 (N_1905,In_1175,In_22);
and U1906 (N_1906,In_1244,In_1657);
or U1907 (N_1907,In_2205,In_496);
xor U1908 (N_1908,In_2166,In_632);
and U1909 (N_1909,In_1377,In_1830);
and U1910 (N_1910,In_63,In_1979);
xnor U1911 (N_1911,In_1833,In_207);
nand U1912 (N_1912,In_897,In_1899);
nor U1913 (N_1913,In_123,In_2005);
nand U1914 (N_1914,In_1783,In_2310);
or U1915 (N_1915,In_721,In_1682);
nor U1916 (N_1916,In_319,In_745);
and U1917 (N_1917,In_1617,In_932);
nand U1918 (N_1918,In_1257,In_1501);
and U1919 (N_1919,In_727,In_370);
nand U1920 (N_1920,In_517,In_1901);
xor U1921 (N_1921,In_2024,In_1547);
or U1922 (N_1922,In_1597,In_1639);
or U1923 (N_1923,In_36,In_229);
nand U1924 (N_1924,In_538,In_613);
xnor U1925 (N_1925,In_1909,In_657);
xor U1926 (N_1926,In_2135,In_84);
and U1927 (N_1927,In_1358,In_300);
nor U1928 (N_1928,In_1624,In_937);
nand U1929 (N_1929,In_263,In_2193);
and U1930 (N_1930,In_210,In_1091);
or U1931 (N_1931,In_351,In_1401);
nand U1932 (N_1932,In_2308,In_1945);
or U1933 (N_1933,In_887,In_1852);
and U1934 (N_1934,In_1544,In_1777);
and U1935 (N_1935,In_64,In_1676);
xnor U1936 (N_1936,In_822,In_703);
and U1937 (N_1937,In_2222,In_1046);
nor U1938 (N_1938,In_1206,In_273);
xor U1939 (N_1939,In_1079,In_1530);
xnor U1940 (N_1940,In_598,In_1017);
xor U1941 (N_1941,In_1018,In_508);
nor U1942 (N_1942,In_2345,In_1951);
nand U1943 (N_1943,In_272,In_2101);
nand U1944 (N_1944,In_2271,In_2169);
xnor U1945 (N_1945,In_1329,In_1160);
nand U1946 (N_1946,In_1505,In_608);
nor U1947 (N_1947,In_615,In_879);
or U1948 (N_1948,In_1028,In_2168);
xor U1949 (N_1949,In_221,In_1461);
xor U1950 (N_1950,In_2005,In_1436);
and U1951 (N_1951,In_558,In_1054);
xor U1952 (N_1952,In_1976,In_853);
xnor U1953 (N_1953,In_951,In_370);
nor U1954 (N_1954,In_1898,In_1622);
xor U1955 (N_1955,In_54,In_1101);
xor U1956 (N_1956,In_160,In_1029);
nor U1957 (N_1957,In_1160,In_1419);
xnor U1958 (N_1958,In_1021,In_559);
or U1959 (N_1959,In_686,In_1036);
and U1960 (N_1960,In_1729,In_460);
nand U1961 (N_1961,In_238,In_559);
and U1962 (N_1962,In_1235,In_2181);
nand U1963 (N_1963,In_1635,In_24);
nand U1964 (N_1964,In_142,In_294);
and U1965 (N_1965,In_321,In_259);
or U1966 (N_1966,In_1638,In_2198);
nor U1967 (N_1967,In_83,In_2064);
nand U1968 (N_1968,In_2050,In_916);
xnor U1969 (N_1969,In_2366,In_1618);
nand U1970 (N_1970,In_1830,In_1891);
or U1971 (N_1971,In_587,In_1974);
nor U1972 (N_1972,In_1544,In_985);
and U1973 (N_1973,In_593,In_588);
and U1974 (N_1974,In_2441,In_1269);
and U1975 (N_1975,In_1284,In_1263);
nand U1976 (N_1976,In_904,In_2188);
or U1977 (N_1977,In_1572,In_1904);
and U1978 (N_1978,In_1989,In_1004);
nor U1979 (N_1979,In_459,In_1258);
nor U1980 (N_1980,In_1504,In_988);
nor U1981 (N_1981,In_1843,In_894);
nor U1982 (N_1982,In_2295,In_2045);
nand U1983 (N_1983,In_1184,In_184);
or U1984 (N_1984,In_587,In_1057);
or U1985 (N_1985,In_790,In_1670);
or U1986 (N_1986,In_945,In_2499);
nor U1987 (N_1987,In_1903,In_1750);
and U1988 (N_1988,In_2027,In_1563);
and U1989 (N_1989,In_15,In_1139);
xnor U1990 (N_1990,In_1820,In_2302);
xnor U1991 (N_1991,In_825,In_244);
and U1992 (N_1992,In_1099,In_1542);
xor U1993 (N_1993,In_141,In_2432);
and U1994 (N_1994,In_1025,In_1881);
xnor U1995 (N_1995,In_2364,In_797);
nand U1996 (N_1996,In_2460,In_2114);
or U1997 (N_1997,In_207,In_1781);
xor U1998 (N_1998,In_1540,In_2348);
nand U1999 (N_1999,In_1600,In_2347);
and U2000 (N_2000,In_1251,In_1073);
or U2001 (N_2001,In_4,In_227);
or U2002 (N_2002,In_36,In_2093);
nand U2003 (N_2003,In_1722,In_827);
xnor U2004 (N_2004,In_774,In_200);
and U2005 (N_2005,In_1805,In_968);
nor U2006 (N_2006,In_4,In_2358);
nand U2007 (N_2007,In_1402,In_371);
nand U2008 (N_2008,In_860,In_513);
nand U2009 (N_2009,In_1684,In_197);
nor U2010 (N_2010,In_825,In_1317);
nand U2011 (N_2011,In_612,In_1613);
or U2012 (N_2012,In_28,In_1830);
xor U2013 (N_2013,In_2291,In_61);
nor U2014 (N_2014,In_1497,In_201);
nor U2015 (N_2015,In_2296,In_4);
nand U2016 (N_2016,In_116,In_81);
xnor U2017 (N_2017,In_1274,In_1648);
or U2018 (N_2018,In_970,In_1441);
or U2019 (N_2019,In_2466,In_1595);
nor U2020 (N_2020,In_43,In_646);
nor U2021 (N_2021,In_136,In_1456);
nand U2022 (N_2022,In_1518,In_2227);
nand U2023 (N_2023,In_1126,In_1251);
nand U2024 (N_2024,In_2410,In_1602);
nor U2025 (N_2025,In_576,In_914);
and U2026 (N_2026,In_836,In_1765);
xor U2027 (N_2027,In_1673,In_1916);
nor U2028 (N_2028,In_1852,In_2070);
nor U2029 (N_2029,In_1654,In_978);
nand U2030 (N_2030,In_457,In_393);
or U2031 (N_2031,In_370,In_290);
xnor U2032 (N_2032,In_788,In_905);
xor U2033 (N_2033,In_1440,In_750);
or U2034 (N_2034,In_1991,In_1589);
nor U2035 (N_2035,In_1235,In_2017);
or U2036 (N_2036,In_2033,In_1607);
and U2037 (N_2037,In_1266,In_2010);
or U2038 (N_2038,In_1750,In_1410);
nor U2039 (N_2039,In_870,In_1648);
or U2040 (N_2040,In_2027,In_1202);
nor U2041 (N_2041,In_471,In_528);
nor U2042 (N_2042,In_331,In_1875);
xnor U2043 (N_2043,In_2263,In_819);
and U2044 (N_2044,In_1456,In_1146);
nand U2045 (N_2045,In_1549,In_2046);
nand U2046 (N_2046,In_432,In_606);
nor U2047 (N_2047,In_1396,In_458);
xor U2048 (N_2048,In_2067,In_928);
nor U2049 (N_2049,In_1015,In_2072);
xor U2050 (N_2050,In_1991,In_1231);
xor U2051 (N_2051,In_2247,In_446);
or U2052 (N_2052,In_469,In_1297);
nand U2053 (N_2053,In_124,In_1090);
or U2054 (N_2054,In_787,In_1990);
or U2055 (N_2055,In_1350,In_1227);
nor U2056 (N_2056,In_113,In_1113);
and U2057 (N_2057,In_324,In_1817);
nor U2058 (N_2058,In_914,In_567);
or U2059 (N_2059,In_950,In_2352);
xnor U2060 (N_2060,In_1037,In_2359);
xnor U2061 (N_2061,In_2336,In_137);
nand U2062 (N_2062,In_52,In_1898);
or U2063 (N_2063,In_2237,In_1136);
or U2064 (N_2064,In_913,In_72);
nand U2065 (N_2065,In_1157,In_1335);
and U2066 (N_2066,In_873,In_2136);
nor U2067 (N_2067,In_1979,In_929);
nor U2068 (N_2068,In_957,In_810);
or U2069 (N_2069,In_2337,In_2468);
nand U2070 (N_2070,In_2062,In_901);
nor U2071 (N_2071,In_1159,In_897);
nor U2072 (N_2072,In_211,In_2099);
xor U2073 (N_2073,In_761,In_2455);
nand U2074 (N_2074,In_2287,In_2035);
nand U2075 (N_2075,In_248,In_722);
xnor U2076 (N_2076,In_1407,In_514);
xor U2077 (N_2077,In_375,In_2248);
and U2078 (N_2078,In_400,In_2012);
nor U2079 (N_2079,In_607,In_1636);
nand U2080 (N_2080,In_649,In_163);
xnor U2081 (N_2081,In_2144,In_137);
and U2082 (N_2082,In_664,In_886);
xnor U2083 (N_2083,In_1651,In_1018);
or U2084 (N_2084,In_9,In_1686);
nor U2085 (N_2085,In_617,In_246);
xnor U2086 (N_2086,In_1395,In_1301);
nor U2087 (N_2087,In_1985,In_2355);
or U2088 (N_2088,In_1813,In_1896);
and U2089 (N_2089,In_1878,In_1484);
nor U2090 (N_2090,In_487,In_1932);
or U2091 (N_2091,In_1308,In_2269);
nand U2092 (N_2092,In_2074,In_1900);
nor U2093 (N_2093,In_397,In_1464);
and U2094 (N_2094,In_1562,In_1303);
and U2095 (N_2095,In_1816,In_1128);
nand U2096 (N_2096,In_2448,In_702);
nor U2097 (N_2097,In_1614,In_1361);
and U2098 (N_2098,In_2255,In_1071);
nand U2099 (N_2099,In_1959,In_1006);
or U2100 (N_2100,In_102,In_691);
and U2101 (N_2101,In_26,In_1781);
and U2102 (N_2102,In_1579,In_2429);
and U2103 (N_2103,In_1980,In_2493);
or U2104 (N_2104,In_925,In_189);
nor U2105 (N_2105,In_139,In_1187);
or U2106 (N_2106,In_1238,In_1294);
nand U2107 (N_2107,In_683,In_2087);
xor U2108 (N_2108,In_782,In_2172);
or U2109 (N_2109,In_2159,In_193);
nand U2110 (N_2110,In_1754,In_1336);
nor U2111 (N_2111,In_2290,In_303);
nor U2112 (N_2112,In_1147,In_687);
xnor U2113 (N_2113,In_469,In_2038);
xor U2114 (N_2114,In_583,In_1533);
nand U2115 (N_2115,In_2445,In_1214);
or U2116 (N_2116,In_1872,In_767);
nand U2117 (N_2117,In_315,In_1200);
or U2118 (N_2118,In_2098,In_1872);
nand U2119 (N_2119,In_89,In_1218);
nor U2120 (N_2120,In_2453,In_1504);
and U2121 (N_2121,In_1954,In_2158);
xnor U2122 (N_2122,In_879,In_821);
and U2123 (N_2123,In_254,In_1143);
and U2124 (N_2124,In_1727,In_1696);
and U2125 (N_2125,In_2418,In_1275);
or U2126 (N_2126,In_1977,In_1729);
nand U2127 (N_2127,In_1617,In_2415);
xnor U2128 (N_2128,In_1283,In_2277);
or U2129 (N_2129,In_2411,In_1665);
xor U2130 (N_2130,In_1218,In_1074);
xor U2131 (N_2131,In_44,In_1041);
and U2132 (N_2132,In_2381,In_2149);
xor U2133 (N_2133,In_2325,In_2040);
xnor U2134 (N_2134,In_699,In_1667);
or U2135 (N_2135,In_289,In_137);
nand U2136 (N_2136,In_2395,In_2388);
nand U2137 (N_2137,In_225,In_329);
nand U2138 (N_2138,In_2458,In_1992);
nor U2139 (N_2139,In_97,In_1265);
nor U2140 (N_2140,In_812,In_397);
and U2141 (N_2141,In_8,In_1654);
xor U2142 (N_2142,In_1178,In_272);
nor U2143 (N_2143,In_1698,In_484);
nand U2144 (N_2144,In_1118,In_400);
xor U2145 (N_2145,In_1723,In_1475);
nor U2146 (N_2146,In_1793,In_149);
and U2147 (N_2147,In_1850,In_630);
nand U2148 (N_2148,In_644,In_954);
or U2149 (N_2149,In_1308,In_631);
nor U2150 (N_2150,In_1240,In_137);
nand U2151 (N_2151,In_487,In_1109);
xnor U2152 (N_2152,In_866,In_1459);
nor U2153 (N_2153,In_613,In_1159);
or U2154 (N_2154,In_213,In_1817);
nand U2155 (N_2155,In_2018,In_329);
and U2156 (N_2156,In_1832,In_1294);
nor U2157 (N_2157,In_1335,In_314);
xnor U2158 (N_2158,In_1685,In_1326);
or U2159 (N_2159,In_2301,In_2282);
nand U2160 (N_2160,In_2120,In_1580);
xnor U2161 (N_2161,In_2462,In_811);
and U2162 (N_2162,In_1209,In_1500);
or U2163 (N_2163,In_1177,In_1002);
nor U2164 (N_2164,In_1546,In_1308);
or U2165 (N_2165,In_2239,In_1970);
xor U2166 (N_2166,In_442,In_897);
xnor U2167 (N_2167,In_100,In_27);
nor U2168 (N_2168,In_1666,In_467);
nand U2169 (N_2169,In_2425,In_2451);
or U2170 (N_2170,In_1679,In_445);
xor U2171 (N_2171,In_462,In_918);
nor U2172 (N_2172,In_63,In_565);
or U2173 (N_2173,In_460,In_802);
nor U2174 (N_2174,In_435,In_2347);
nor U2175 (N_2175,In_1061,In_686);
nor U2176 (N_2176,In_278,In_349);
nand U2177 (N_2177,In_1916,In_710);
nor U2178 (N_2178,In_1409,In_821);
xor U2179 (N_2179,In_1781,In_1490);
xor U2180 (N_2180,In_1549,In_2364);
and U2181 (N_2181,In_32,In_1238);
nor U2182 (N_2182,In_1721,In_1435);
nand U2183 (N_2183,In_2061,In_2243);
xor U2184 (N_2184,In_402,In_978);
nand U2185 (N_2185,In_50,In_708);
nor U2186 (N_2186,In_2406,In_2156);
and U2187 (N_2187,In_155,In_1061);
or U2188 (N_2188,In_220,In_2177);
and U2189 (N_2189,In_1375,In_1883);
or U2190 (N_2190,In_601,In_756);
and U2191 (N_2191,In_1796,In_1375);
nor U2192 (N_2192,In_1641,In_1480);
or U2193 (N_2193,In_2489,In_701);
xor U2194 (N_2194,In_316,In_1349);
nand U2195 (N_2195,In_635,In_550);
or U2196 (N_2196,In_1614,In_1779);
nand U2197 (N_2197,In_155,In_271);
xor U2198 (N_2198,In_280,In_970);
xor U2199 (N_2199,In_1890,In_1684);
nand U2200 (N_2200,In_401,In_1173);
nor U2201 (N_2201,In_2030,In_522);
or U2202 (N_2202,In_616,In_1035);
nand U2203 (N_2203,In_2,In_2352);
xnor U2204 (N_2204,In_570,In_1713);
or U2205 (N_2205,In_1641,In_1613);
nand U2206 (N_2206,In_729,In_1418);
nor U2207 (N_2207,In_299,In_1637);
xor U2208 (N_2208,In_2490,In_1745);
and U2209 (N_2209,In_2178,In_1766);
or U2210 (N_2210,In_2247,In_583);
or U2211 (N_2211,In_1781,In_2384);
nor U2212 (N_2212,In_2248,In_1271);
xor U2213 (N_2213,In_591,In_2464);
and U2214 (N_2214,In_1347,In_1770);
or U2215 (N_2215,In_317,In_739);
xor U2216 (N_2216,In_802,In_1030);
or U2217 (N_2217,In_362,In_1591);
nand U2218 (N_2218,In_432,In_2209);
and U2219 (N_2219,In_586,In_1634);
xor U2220 (N_2220,In_2116,In_1711);
nor U2221 (N_2221,In_426,In_119);
xnor U2222 (N_2222,In_1892,In_718);
or U2223 (N_2223,In_245,In_495);
or U2224 (N_2224,In_144,In_1448);
nand U2225 (N_2225,In_2462,In_427);
nor U2226 (N_2226,In_1325,In_1657);
and U2227 (N_2227,In_2286,In_290);
xnor U2228 (N_2228,In_1708,In_1502);
nand U2229 (N_2229,In_1090,In_2085);
or U2230 (N_2230,In_849,In_1465);
nand U2231 (N_2231,In_725,In_1581);
nor U2232 (N_2232,In_1903,In_444);
or U2233 (N_2233,In_2261,In_1186);
and U2234 (N_2234,In_751,In_1412);
nand U2235 (N_2235,In_2234,In_981);
or U2236 (N_2236,In_2090,In_1241);
nor U2237 (N_2237,In_646,In_522);
nor U2238 (N_2238,In_2373,In_1116);
nand U2239 (N_2239,In_2402,In_1962);
nor U2240 (N_2240,In_1846,In_1470);
and U2241 (N_2241,In_413,In_63);
xor U2242 (N_2242,In_665,In_676);
xor U2243 (N_2243,In_1224,In_495);
xnor U2244 (N_2244,In_1917,In_914);
nand U2245 (N_2245,In_227,In_316);
nor U2246 (N_2246,In_877,In_1410);
nand U2247 (N_2247,In_1778,In_1580);
or U2248 (N_2248,In_30,In_1671);
xnor U2249 (N_2249,In_1753,In_2346);
and U2250 (N_2250,In_1216,In_824);
or U2251 (N_2251,In_2294,In_1642);
nor U2252 (N_2252,In_1036,In_2496);
or U2253 (N_2253,In_84,In_1158);
and U2254 (N_2254,In_521,In_91);
nor U2255 (N_2255,In_473,In_35);
nand U2256 (N_2256,In_945,In_1324);
or U2257 (N_2257,In_855,In_1338);
xnor U2258 (N_2258,In_1460,In_354);
nor U2259 (N_2259,In_1195,In_922);
nand U2260 (N_2260,In_964,In_1485);
nand U2261 (N_2261,In_43,In_70);
nand U2262 (N_2262,In_748,In_1604);
and U2263 (N_2263,In_635,In_2162);
nand U2264 (N_2264,In_1331,In_218);
xnor U2265 (N_2265,In_2008,In_886);
and U2266 (N_2266,In_2207,In_1402);
and U2267 (N_2267,In_826,In_439);
and U2268 (N_2268,In_1464,In_2149);
nor U2269 (N_2269,In_1852,In_295);
xnor U2270 (N_2270,In_2170,In_1801);
or U2271 (N_2271,In_820,In_402);
xnor U2272 (N_2272,In_2247,In_1086);
nor U2273 (N_2273,In_1587,In_2181);
and U2274 (N_2274,In_684,In_2141);
and U2275 (N_2275,In_1019,In_655);
or U2276 (N_2276,In_1960,In_1991);
xor U2277 (N_2277,In_511,In_1828);
and U2278 (N_2278,In_763,In_812);
xor U2279 (N_2279,In_641,In_1224);
or U2280 (N_2280,In_7,In_2461);
and U2281 (N_2281,In_876,In_1628);
or U2282 (N_2282,In_1451,In_731);
and U2283 (N_2283,In_268,In_685);
and U2284 (N_2284,In_36,In_622);
xnor U2285 (N_2285,In_1765,In_115);
nand U2286 (N_2286,In_800,In_353);
nor U2287 (N_2287,In_522,In_1754);
and U2288 (N_2288,In_1917,In_913);
or U2289 (N_2289,In_471,In_925);
nand U2290 (N_2290,In_1564,In_1294);
nor U2291 (N_2291,In_1302,In_1896);
nand U2292 (N_2292,In_1342,In_2415);
nand U2293 (N_2293,In_2303,In_382);
nor U2294 (N_2294,In_1239,In_406);
xor U2295 (N_2295,In_1528,In_2223);
nand U2296 (N_2296,In_1724,In_62);
xor U2297 (N_2297,In_1862,In_708);
nor U2298 (N_2298,In_933,In_1885);
xnor U2299 (N_2299,In_1500,In_788);
nor U2300 (N_2300,In_2469,In_77);
nor U2301 (N_2301,In_676,In_2025);
nand U2302 (N_2302,In_812,In_483);
or U2303 (N_2303,In_134,In_359);
nor U2304 (N_2304,In_2010,In_2149);
nand U2305 (N_2305,In_1877,In_274);
and U2306 (N_2306,In_2346,In_1675);
nand U2307 (N_2307,In_389,In_7);
or U2308 (N_2308,In_927,In_345);
and U2309 (N_2309,In_99,In_1621);
nand U2310 (N_2310,In_876,In_1313);
nand U2311 (N_2311,In_912,In_1545);
or U2312 (N_2312,In_2370,In_1431);
and U2313 (N_2313,In_421,In_306);
nor U2314 (N_2314,In_2108,In_1423);
or U2315 (N_2315,In_212,In_458);
nor U2316 (N_2316,In_1749,In_1853);
nor U2317 (N_2317,In_1063,In_1191);
nand U2318 (N_2318,In_1827,In_2071);
nor U2319 (N_2319,In_2269,In_1182);
and U2320 (N_2320,In_1074,In_681);
xnor U2321 (N_2321,In_1716,In_204);
or U2322 (N_2322,In_1950,In_31);
or U2323 (N_2323,In_50,In_2153);
xnor U2324 (N_2324,In_941,In_264);
nor U2325 (N_2325,In_299,In_85);
xnor U2326 (N_2326,In_120,In_1465);
or U2327 (N_2327,In_556,In_872);
nand U2328 (N_2328,In_1993,In_782);
xor U2329 (N_2329,In_2404,In_883);
xor U2330 (N_2330,In_2053,In_295);
xnor U2331 (N_2331,In_2423,In_2104);
or U2332 (N_2332,In_1757,In_682);
and U2333 (N_2333,In_1883,In_109);
nand U2334 (N_2334,In_330,In_148);
nand U2335 (N_2335,In_309,In_2143);
nor U2336 (N_2336,In_2454,In_2413);
nand U2337 (N_2337,In_1802,In_1925);
nor U2338 (N_2338,In_1738,In_1619);
and U2339 (N_2339,In_217,In_1208);
and U2340 (N_2340,In_590,In_1711);
and U2341 (N_2341,In_1606,In_1801);
nor U2342 (N_2342,In_2489,In_2133);
or U2343 (N_2343,In_59,In_1521);
or U2344 (N_2344,In_416,In_737);
and U2345 (N_2345,In_951,In_1420);
nor U2346 (N_2346,In_1811,In_481);
xor U2347 (N_2347,In_272,In_541);
nand U2348 (N_2348,In_345,In_2195);
or U2349 (N_2349,In_1581,In_1845);
or U2350 (N_2350,In_1961,In_950);
and U2351 (N_2351,In_627,In_1341);
or U2352 (N_2352,In_1163,In_236);
nand U2353 (N_2353,In_767,In_2158);
or U2354 (N_2354,In_2281,In_928);
or U2355 (N_2355,In_962,In_1740);
nor U2356 (N_2356,In_127,In_1005);
nor U2357 (N_2357,In_1313,In_305);
nor U2358 (N_2358,In_97,In_741);
and U2359 (N_2359,In_616,In_1902);
and U2360 (N_2360,In_2049,In_2209);
or U2361 (N_2361,In_794,In_22);
nand U2362 (N_2362,In_498,In_1686);
or U2363 (N_2363,In_908,In_384);
nand U2364 (N_2364,In_170,In_944);
and U2365 (N_2365,In_143,In_2446);
nand U2366 (N_2366,In_114,In_1101);
nand U2367 (N_2367,In_1856,In_2196);
xnor U2368 (N_2368,In_2077,In_1321);
nand U2369 (N_2369,In_740,In_347);
nand U2370 (N_2370,In_2178,In_889);
and U2371 (N_2371,In_1820,In_2479);
or U2372 (N_2372,In_1207,In_2065);
and U2373 (N_2373,In_1865,In_1214);
nand U2374 (N_2374,In_670,In_2332);
nand U2375 (N_2375,In_2317,In_554);
xor U2376 (N_2376,In_2248,In_449);
nor U2377 (N_2377,In_1912,In_665);
nor U2378 (N_2378,In_2353,In_1162);
nor U2379 (N_2379,In_2332,In_367);
nand U2380 (N_2380,In_722,In_1078);
nor U2381 (N_2381,In_1147,In_473);
or U2382 (N_2382,In_1233,In_384);
nand U2383 (N_2383,In_712,In_875);
and U2384 (N_2384,In_714,In_1946);
xor U2385 (N_2385,In_1626,In_2269);
nand U2386 (N_2386,In_1333,In_43);
or U2387 (N_2387,In_781,In_1039);
and U2388 (N_2388,In_286,In_1345);
nand U2389 (N_2389,In_1409,In_695);
and U2390 (N_2390,In_501,In_2161);
or U2391 (N_2391,In_1336,In_434);
xor U2392 (N_2392,In_521,In_1293);
or U2393 (N_2393,In_1149,In_1938);
and U2394 (N_2394,In_349,In_727);
or U2395 (N_2395,In_2412,In_1822);
and U2396 (N_2396,In_2418,In_365);
nor U2397 (N_2397,In_2153,In_1861);
nor U2398 (N_2398,In_1291,In_450);
xor U2399 (N_2399,In_1404,In_384);
or U2400 (N_2400,In_180,In_1488);
xnor U2401 (N_2401,In_2128,In_1549);
xnor U2402 (N_2402,In_2231,In_29);
xor U2403 (N_2403,In_391,In_2414);
or U2404 (N_2404,In_2165,In_604);
or U2405 (N_2405,In_724,In_1801);
nand U2406 (N_2406,In_713,In_162);
or U2407 (N_2407,In_3,In_1321);
nor U2408 (N_2408,In_1092,In_86);
nand U2409 (N_2409,In_1424,In_1529);
nor U2410 (N_2410,In_1798,In_134);
xnor U2411 (N_2411,In_402,In_1909);
nand U2412 (N_2412,In_1733,In_589);
xnor U2413 (N_2413,In_2074,In_1007);
or U2414 (N_2414,In_470,In_36);
or U2415 (N_2415,In_1203,In_726);
and U2416 (N_2416,In_850,In_1409);
nor U2417 (N_2417,In_2117,In_103);
and U2418 (N_2418,In_1475,In_735);
and U2419 (N_2419,In_2258,In_511);
nand U2420 (N_2420,In_2056,In_1335);
and U2421 (N_2421,In_1757,In_1339);
nand U2422 (N_2422,In_73,In_1405);
or U2423 (N_2423,In_423,In_2379);
nand U2424 (N_2424,In_1837,In_1736);
nand U2425 (N_2425,In_788,In_239);
or U2426 (N_2426,In_361,In_920);
nand U2427 (N_2427,In_1587,In_1303);
nor U2428 (N_2428,In_574,In_919);
xnor U2429 (N_2429,In_210,In_149);
nand U2430 (N_2430,In_1759,In_705);
and U2431 (N_2431,In_337,In_458);
xnor U2432 (N_2432,In_1950,In_371);
nand U2433 (N_2433,In_1050,In_691);
and U2434 (N_2434,In_1440,In_2233);
xnor U2435 (N_2435,In_120,In_997);
or U2436 (N_2436,In_846,In_297);
and U2437 (N_2437,In_374,In_512);
nand U2438 (N_2438,In_1375,In_497);
nor U2439 (N_2439,In_859,In_1784);
nor U2440 (N_2440,In_1341,In_610);
nor U2441 (N_2441,In_2265,In_111);
and U2442 (N_2442,In_957,In_1102);
or U2443 (N_2443,In_837,In_1882);
xnor U2444 (N_2444,In_1771,In_1576);
nand U2445 (N_2445,In_864,In_1401);
xor U2446 (N_2446,In_6,In_1802);
and U2447 (N_2447,In_1590,In_869);
and U2448 (N_2448,In_842,In_1834);
nand U2449 (N_2449,In_1124,In_1973);
and U2450 (N_2450,In_193,In_1340);
nand U2451 (N_2451,In_1335,In_2183);
nor U2452 (N_2452,In_2345,In_306);
nand U2453 (N_2453,In_741,In_945);
or U2454 (N_2454,In_1862,In_1356);
and U2455 (N_2455,In_79,In_2425);
xnor U2456 (N_2456,In_2187,In_1913);
and U2457 (N_2457,In_511,In_563);
and U2458 (N_2458,In_326,In_1908);
and U2459 (N_2459,In_889,In_1851);
nor U2460 (N_2460,In_1032,In_2127);
or U2461 (N_2461,In_130,In_1928);
and U2462 (N_2462,In_1080,In_284);
xor U2463 (N_2463,In_2181,In_2174);
or U2464 (N_2464,In_2234,In_1954);
nand U2465 (N_2465,In_943,In_1765);
nor U2466 (N_2466,In_1435,In_1197);
xnor U2467 (N_2467,In_2226,In_2233);
xor U2468 (N_2468,In_207,In_1600);
and U2469 (N_2469,In_2320,In_949);
nand U2470 (N_2470,In_1219,In_103);
and U2471 (N_2471,In_1022,In_2395);
or U2472 (N_2472,In_1957,In_2230);
or U2473 (N_2473,In_1530,In_1160);
xor U2474 (N_2474,In_1697,In_1065);
xor U2475 (N_2475,In_982,In_2121);
xnor U2476 (N_2476,In_1988,In_252);
and U2477 (N_2477,In_106,In_571);
nor U2478 (N_2478,In_1378,In_1690);
nor U2479 (N_2479,In_553,In_2366);
xnor U2480 (N_2480,In_1311,In_104);
and U2481 (N_2481,In_1831,In_2295);
nor U2482 (N_2482,In_898,In_1488);
or U2483 (N_2483,In_2354,In_1621);
or U2484 (N_2484,In_1467,In_750);
nor U2485 (N_2485,In_309,In_219);
and U2486 (N_2486,In_2271,In_11);
xnor U2487 (N_2487,In_738,In_1922);
xnor U2488 (N_2488,In_2498,In_2306);
xnor U2489 (N_2489,In_707,In_1674);
nor U2490 (N_2490,In_2278,In_861);
nor U2491 (N_2491,In_1745,In_2090);
xor U2492 (N_2492,In_2241,In_1387);
nand U2493 (N_2493,In_481,In_1725);
and U2494 (N_2494,In_170,In_367);
nor U2495 (N_2495,In_406,In_577);
nor U2496 (N_2496,In_1014,In_2451);
and U2497 (N_2497,In_1901,In_1976);
or U2498 (N_2498,In_496,In_2074);
xnor U2499 (N_2499,In_787,In_1405);
nand U2500 (N_2500,In_1108,In_203);
xnor U2501 (N_2501,In_628,In_26);
and U2502 (N_2502,In_2025,In_1365);
xnor U2503 (N_2503,In_2281,In_1600);
nand U2504 (N_2504,In_2426,In_1608);
and U2505 (N_2505,In_46,In_495);
or U2506 (N_2506,In_1526,In_363);
xor U2507 (N_2507,In_1983,In_23);
xor U2508 (N_2508,In_2439,In_1051);
or U2509 (N_2509,In_1863,In_1150);
or U2510 (N_2510,In_2053,In_448);
xnor U2511 (N_2511,In_1389,In_1707);
xnor U2512 (N_2512,In_2413,In_2022);
nand U2513 (N_2513,In_1999,In_1601);
nand U2514 (N_2514,In_566,In_1864);
and U2515 (N_2515,In_2257,In_42);
or U2516 (N_2516,In_503,In_1163);
nor U2517 (N_2517,In_2248,In_1190);
nor U2518 (N_2518,In_692,In_1999);
or U2519 (N_2519,In_111,In_1920);
or U2520 (N_2520,In_2067,In_1460);
or U2521 (N_2521,In_2104,In_844);
xnor U2522 (N_2522,In_220,In_2209);
and U2523 (N_2523,In_1642,In_1153);
and U2524 (N_2524,In_1605,In_2275);
nor U2525 (N_2525,In_948,In_246);
xnor U2526 (N_2526,In_616,In_808);
nor U2527 (N_2527,In_1969,In_677);
nand U2528 (N_2528,In_302,In_1199);
and U2529 (N_2529,In_493,In_243);
or U2530 (N_2530,In_2194,In_1589);
nand U2531 (N_2531,In_444,In_1971);
nor U2532 (N_2532,In_418,In_2136);
nand U2533 (N_2533,In_1507,In_791);
nand U2534 (N_2534,In_437,In_1617);
and U2535 (N_2535,In_1714,In_1815);
nor U2536 (N_2536,In_20,In_1841);
xnor U2537 (N_2537,In_777,In_313);
or U2538 (N_2538,In_1910,In_1097);
and U2539 (N_2539,In_265,In_1434);
nor U2540 (N_2540,In_976,In_876);
and U2541 (N_2541,In_2229,In_1967);
or U2542 (N_2542,In_759,In_1974);
xnor U2543 (N_2543,In_2209,In_2461);
xor U2544 (N_2544,In_326,In_1256);
and U2545 (N_2545,In_145,In_937);
or U2546 (N_2546,In_2459,In_2270);
nand U2547 (N_2547,In_609,In_2115);
and U2548 (N_2548,In_436,In_2028);
and U2549 (N_2549,In_2478,In_1898);
nand U2550 (N_2550,In_663,In_1707);
xor U2551 (N_2551,In_797,In_247);
nor U2552 (N_2552,In_2023,In_2229);
xor U2553 (N_2553,In_1738,In_2103);
nand U2554 (N_2554,In_556,In_475);
xnor U2555 (N_2555,In_473,In_1813);
nand U2556 (N_2556,In_1490,In_1330);
or U2557 (N_2557,In_1567,In_1654);
nand U2558 (N_2558,In_330,In_680);
xnor U2559 (N_2559,In_2195,In_1121);
xor U2560 (N_2560,In_1924,In_1588);
nand U2561 (N_2561,In_1775,In_1077);
or U2562 (N_2562,In_2164,In_48);
or U2563 (N_2563,In_1355,In_137);
or U2564 (N_2564,In_1543,In_288);
or U2565 (N_2565,In_1505,In_1661);
nor U2566 (N_2566,In_434,In_360);
nand U2567 (N_2567,In_2069,In_2067);
xnor U2568 (N_2568,In_1260,In_1611);
or U2569 (N_2569,In_2324,In_197);
and U2570 (N_2570,In_743,In_2480);
nor U2571 (N_2571,In_2448,In_1906);
or U2572 (N_2572,In_1976,In_1593);
nor U2573 (N_2573,In_674,In_2165);
or U2574 (N_2574,In_1130,In_351);
or U2575 (N_2575,In_1404,In_1694);
nand U2576 (N_2576,In_2206,In_1852);
or U2577 (N_2577,In_632,In_2054);
nand U2578 (N_2578,In_1055,In_1169);
nor U2579 (N_2579,In_510,In_1440);
or U2580 (N_2580,In_626,In_730);
or U2581 (N_2581,In_1492,In_1913);
and U2582 (N_2582,In_327,In_998);
xor U2583 (N_2583,In_852,In_689);
nor U2584 (N_2584,In_1775,In_2390);
and U2585 (N_2585,In_316,In_875);
and U2586 (N_2586,In_1294,In_1807);
nand U2587 (N_2587,In_512,In_545);
or U2588 (N_2588,In_2082,In_2410);
nand U2589 (N_2589,In_1478,In_33);
or U2590 (N_2590,In_2012,In_1618);
or U2591 (N_2591,In_20,In_1563);
and U2592 (N_2592,In_355,In_2422);
nand U2593 (N_2593,In_460,In_1601);
xor U2594 (N_2594,In_2316,In_133);
and U2595 (N_2595,In_2287,In_2367);
xnor U2596 (N_2596,In_1832,In_2234);
and U2597 (N_2597,In_1319,In_2075);
or U2598 (N_2598,In_1379,In_2488);
nand U2599 (N_2599,In_363,In_2420);
or U2600 (N_2600,In_1379,In_2152);
and U2601 (N_2601,In_2093,In_1674);
xnor U2602 (N_2602,In_1338,In_1487);
xnor U2603 (N_2603,In_282,In_1747);
xnor U2604 (N_2604,In_2072,In_1957);
and U2605 (N_2605,In_1154,In_516);
xor U2606 (N_2606,In_1710,In_773);
nor U2607 (N_2607,In_1172,In_1502);
nor U2608 (N_2608,In_2467,In_1863);
xor U2609 (N_2609,In_1140,In_2075);
nand U2610 (N_2610,In_711,In_478);
nand U2611 (N_2611,In_1123,In_65);
xnor U2612 (N_2612,In_836,In_968);
nor U2613 (N_2613,In_939,In_1001);
nand U2614 (N_2614,In_1763,In_2490);
xnor U2615 (N_2615,In_927,In_2324);
nor U2616 (N_2616,In_964,In_1831);
nand U2617 (N_2617,In_1391,In_1456);
nand U2618 (N_2618,In_1537,In_353);
and U2619 (N_2619,In_1910,In_568);
nor U2620 (N_2620,In_437,In_1456);
nor U2621 (N_2621,In_1803,In_2293);
xor U2622 (N_2622,In_1866,In_253);
or U2623 (N_2623,In_510,In_2311);
xor U2624 (N_2624,In_2007,In_1976);
xor U2625 (N_2625,In_1307,In_548);
nand U2626 (N_2626,In_1846,In_851);
nand U2627 (N_2627,In_617,In_291);
nand U2628 (N_2628,In_1078,In_63);
or U2629 (N_2629,In_1018,In_1653);
nor U2630 (N_2630,In_1745,In_1709);
and U2631 (N_2631,In_1284,In_2242);
xor U2632 (N_2632,In_1517,In_2105);
nand U2633 (N_2633,In_2087,In_1829);
nor U2634 (N_2634,In_272,In_1555);
nand U2635 (N_2635,In_960,In_91);
and U2636 (N_2636,In_1304,In_2450);
or U2637 (N_2637,In_540,In_921);
and U2638 (N_2638,In_1733,In_1319);
or U2639 (N_2639,In_1055,In_2386);
and U2640 (N_2640,In_2165,In_1087);
nand U2641 (N_2641,In_710,In_2198);
nand U2642 (N_2642,In_1993,In_1047);
and U2643 (N_2643,In_1786,In_2406);
xnor U2644 (N_2644,In_1354,In_1741);
xor U2645 (N_2645,In_2324,In_1786);
nor U2646 (N_2646,In_1205,In_2253);
nor U2647 (N_2647,In_756,In_2330);
nand U2648 (N_2648,In_1681,In_113);
nor U2649 (N_2649,In_1634,In_1714);
nand U2650 (N_2650,In_834,In_572);
nor U2651 (N_2651,In_759,In_372);
and U2652 (N_2652,In_1149,In_631);
or U2653 (N_2653,In_967,In_1671);
nor U2654 (N_2654,In_2045,In_260);
nand U2655 (N_2655,In_601,In_1242);
nand U2656 (N_2656,In_2096,In_1448);
nand U2657 (N_2657,In_1916,In_452);
or U2658 (N_2658,In_210,In_938);
xnor U2659 (N_2659,In_1280,In_221);
or U2660 (N_2660,In_1939,In_221);
nand U2661 (N_2661,In_984,In_931);
nor U2662 (N_2662,In_694,In_693);
and U2663 (N_2663,In_1262,In_321);
nor U2664 (N_2664,In_2338,In_616);
and U2665 (N_2665,In_25,In_196);
nor U2666 (N_2666,In_1763,In_1548);
nor U2667 (N_2667,In_1247,In_1047);
nor U2668 (N_2668,In_2265,In_1182);
nand U2669 (N_2669,In_18,In_2185);
or U2670 (N_2670,In_1398,In_413);
nor U2671 (N_2671,In_355,In_1230);
nand U2672 (N_2672,In_299,In_2234);
nor U2673 (N_2673,In_1821,In_667);
nor U2674 (N_2674,In_1463,In_1420);
nor U2675 (N_2675,In_1343,In_1878);
nand U2676 (N_2676,In_2435,In_1604);
or U2677 (N_2677,In_2121,In_1657);
nand U2678 (N_2678,In_713,In_392);
nand U2679 (N_2679,In_1263,In_1644);
or U2680 (N_2680,In_582,In_1672);
nor U2681 (N_2681,In_2430,In_799);
and U2682 (N_2682,In_1883,In_1121);
and U2683 (N_2683,In_350,In_895);
or U2684 (N_2684,In_1450,In_1115);
and U2685 (N_2685,In_1909,In_546);
and U2686 (N_2686,In_1245,In_1355);
or U2687 (N_2687,In_1808,In_1373);
or U2688 (N_2688,In_522,In_1901);
xnor U2689 (N_2689,In_1015,In_232);
nor U2690 (N_2690,In_2315,In_942);
or U2691 (N_2691,In_2121,In_2352);
xor U2692 (N_2692,In_557,In_11);
and U2693 (N_2693,In_2242,In_983);
or U2694 (N_2694,In_1800,In_311);
xor U2695 (N_2695,In_1809,In_940);
nor U2696 (N_2696,In_2086,In_1292);
or U2697 (N_2697,In_1949,In_822);
or U2698 (N_2698,In_1318,In_2369);
or U2699 (N_2699,In_87,In_940);
xnor U2700 (N_2700,In_932,In_1488);
nor U2701 (N_2701,In_2215,In_2255);
and U2702 (N_2702,In_2207,In_403);
or U2703 (N_2703,In_1681,In_1693);
nor U2704 (N_2704,In_1324,In_2468);
nand U2705 (N_2705,In_1015,In_1741);
and U2706 (N_2706,In_2043,In_943);
nand U2707 (N_2707,In_527,In_965);
and U2708 (N_2708,In_157,In_2275);
xnor U2709 (N_2709,In_1032,In_1716);
xnor U2710 (N_2710,In_179,In_1509);
and U2711 (N_2711,In_1117,In_382);
nor U2712 (N_2712,In_914,In_660);
nand U2713 (N_2713,In_1148,In_2099);
nand U2714 (N_2714,In_2197,In_523);
or U2715 (N_2715,In_388,In_2062);
and U2716 (N_2716,In_1204,In_634);
xnor U2717 (N_2717,In_309,In_2484);
or U2718 (N_2718,In_13,In_1909);
or U2719 (N_2719,In_526,In_2203);
or U2720 (N_2720,In_686,In_1306);
nor U2721 (N_2721,In_1458,In_1354);
and U2722 (N_2722,In_1993,In_460);
xnor U2723 (N_2723,In_1900,In_2377);
xnor U2724 (N_2724,In_629,In_4);
nor U2725 (N_2725,In_1127,In_271);
nand U2726 (N_2726,In_1883,In_168);
and U2727 (N_2727,In_837,In_1165);
and U2728 (N_2728,In_242,In_889);
nand U2729 (N_2729,In_1163,In_1933);
xor U2730 (N_2730,In_1694,In_1024);
nand U2731 (N_2731,In_1226,In_1859);
nor U2732 (N_2732,In_2024,In_571);
xnor U2733 (N_2733,In_1080,In_1019);
xnor U2734 (N_2734,In_1223,In_903);
nor U2735 (N_2735,In_1628,In_451);
nand U2736 (N_2736,In_361,In_174);
and U2737 (N_2737,In_389,In_58);
and U2738 (N_2738,In_1408,In_2171);
nor U2739 (N_2739,In_625,In_2457);
nand U2740 (N_2740,In_530,In_2335);
nor U2741 (N_2741,In_44,In_724);
nand U2742 (N_2742,In_2128,In_1462);
and U2743 (N_2743,In_2345,In_837);
xor U2744 (N_2744,In_2352,In_1508);
and U2745 (N_2745,In_1333,In_965);
or U2746 (N_2746,In_301,In_2277);
or U2747 (N_2747,In_282,In_1533);
or U2748 (N_2748,In_1706,In_1572);
nor U2749 (N_2749,In_1818,In_1881);
and U2750 (N_2750,In_2112,In_817);
nand U2751 (N_2751,In_2333,In_988);
and U2752 (N_2752,In_377,In_1902);
nand U2753 (N_2753,In_2061,In_2458);
or U2754 (N_2754,In_1411,In_1481);
xnor U2755 (N_2755,In_1099,In_1047);
or U2756 (N_2756,In_2475,In_428);
and U2757 (N_2757,In_2208,In_2000);
nand U2758 (N_2758,In_1447,In_996);
nor U2759 (N_2759,In_122,In_81);
nor U2760 (N_2760,In_1218,In_1627);
or U2761 (N_2761,In_690,In_572);
or U2762 (N_2762,In_1044,In_432);
xnor U2763 (N_2763,In_2322,In_1511);
nand U2764 (N_2764,In_1108,In_263);
nand U2765 (N_2765,In_1454,In_272);
nand U2766 (N_2766,In_1410,In_2035);
nor U2767 (N_2767,In_2065,In_152);
or U2768 (N_2768,In_1912,In_430);
nor U2769 (N_2769,In_1372,In_455);
nor U2770 (N_2770,In_2207,In_183);
or U2771 (N_2771,In_1672,In_716);
xnor U2772 (N_2772,In_1218,In_453);
and U2773 (N_2773,In_1632,In_469);
and U2774 (N_2774,In_2381,In_1448);
nand U2775 (N_2775,In_2017,In_403);
or U2776 (N_2776,In_357,In_912);
nor U2777 (N_2777,In_2193,In_1298);
xor U2778 (N_2778,In_2441,In_1273);
nor U2779 (N_2779,In_1447,In_490);
xor U2780 (N_2780,In_1564,In_536);
xor U2781 (N_2781,In_818,In_1039);
or U2782 (N_2782,In_222,In_1911);
or U2783 (N_2783,In_301,In_1866);
nand U2784 (N_2784,In_2062,In_944);
nor U2785 (N_2785,In_1507,In_2314);
or U2786 (N_2786,In_1845,In_933);
xor U2787 (N_2787,In_2316,In_1395);
nand U2788 (N_2788,In_1932,In_2362);
nor U2789 (N_2789,In_896,In_2336);
or U2790 (N_2790,In_2493,In_183);
xor U2791 (N_2791,In_1841,In_488);
or U2792 (N_2792,In_2125,In_1104);
nand U2793 (N_2793,In_495,In_1631);
nor U2794 (N_2794,In_2026,In_2145);
or U2795 (N_2795,In_453,In_2392);
xor U2796 (N_2796,In_2420,In_2055);
xor U2797 (N_2797,In_1446,In_344);
and U2798 (N_2798,In_383,In_1574);
nand U2799 (N_2799,In_315,In_2009);
nor U2800 (N_2800,In_1316,In_2075);
nor U2801 (N_2801,In_368,In_2343);
and U2802 (N_2802,In_1715,In_531);
or U2803 (N_2803,In_2022,In_1171);
nand U2804 (N_2804,In_1302,In_1539);
xnor U2805 (N_2805,In_806,In_1474);
nor U2806 (N_2806,In_1961,In_731);
or U2807 (N_2807,In_1747,In_204);
xor U2808 (N_2808,In_2348,In_625);
nand U2809 (N_2809,In_1061,In_1234);
or U2810 (N_2810,In_1926,In_1454);
xnor U2811 (N_2811,In_997,In_462);
and U2812 (N_2812,In_1245,In_2225);
or U2813 (N_2813,In_25,In_1064);
and U2814 (N_2814,In_365,In_1955);
and U2815 (N_2815,In_2240,In_1882);
or U2816 (N_2816,In_931,In_85);
and U2817 (N_2817,In_2054,In_1898);
and U2818 (N_2818,In_408,In_2309);
nor U2819 (N_2819,In_107,In_2038);
nand U2820 (N_2820,In_1056,In_2005);
or U2821 (N_2821,In_1934,In_687);
xnor U2822 (N_2822,In_1441,In_951);
or U2823 (N_2823,In_2156,In_627);
nor U2824 (N_2824,In_2433,In_1063);
or U2825 (N_2825,In_1598,In_1306);
xor U2826 (N_2826,In_1098,In_1573);
xnor U2827 (N_2827,In_37,In_114);
xor U2828 (N_2828,In_2029,In_632);
xor U2829 (N_2829,In_290,In_782);
and U2830 (N_2830,In_1141,In_2092);
xor U2831 (N_2831,In_1417,In_1936);
xnor U2832 (N_2832,In_2264,In_388);
nand U2833 (N_2833,In_990,In_877);
and U2834 (N_2834,In_1043,In_296);
nand U2835 (N_2835,In_782,In_765);
or U2836 (N_2836,In_1170,In_1792);
or U2837 (N_2837,In_450,In_1135);
nand U2838 (N_2838,In_1339,In_729);
or U2839 (N_2839,In_1006,In_1423);
nand U2840 (N_2840,In_457,In_1299);
nor U2841 (N_2841,In_1255,In_1543);
or U2842 (N_2842,In_1188,In_2474);
nand U2843 (N_2843,In_153,In_2159);
xor U2844 (N_2844,In_182,In_1059);
nand U2845 (N_2845,In_1858,In_1306);
nor U2846 (N_2846,In_2262,In_708);
nand U2847 (N_2847,In_2146,In_948);
xnor U2848 (N_2848,In_1192,In_2098);
nor U2849 (N_2849,In_1275,In_1479);
or U2850 (N_2850,In_1740,In_201);
nor U2851 (N_2851,In_827,In_611);
and U2852 (N_2852,In_428,In_1197);
xor U2853 (N_2853,In_1354,In_751);
and U2854 (N_2854,In_869,In_1776);
nand U2855 (N_2855,In_1660,In_1442);
nand U2856 (N_2856,In_853,In_220);
nand U2857 (N_2857,In_1278,In_277);
or U2858 (N_2858,In_1696,In_122);
xnor U2859 (N_2859,In_808,In_695);
nor U2860 (N_2860,In_2324,In_60);
and U2861 (N_2861,In_256,In_1543);
or U2862 (N_2862,In_1584,In_1575);
or U2863 (N_2863,In_93,In_1161);
nand U2864 (N_2864,In_634,In_1027);
or U2865 (N_2865,In_1865,In_690);
nor U2866 (N_2866,In_115,In_244);
nand U2867 (N_2867,In_2330,In_2248);
xor U2868 (N_2868,In_1506,In_2366);
nand U2869 (N_2869,In_2342,In_908);
or U2870 (N_2870,In_2148,In_1708);
nor U2871 (N_2871,In_1756,In_64);
and U2872 (N_2872,In_1430,In_1844);
nand U2873 (N_2873,In_2007,In_2380);
xnor U2874 (N_2874,In_2169,In_48);
nor U2875 (N_2875,In_4,In_1187);
nand U2876 (N_2876,In_2226,In_2386);
nor U2877 (N_2877,In_1767,In_965);
and U2878 (N_2878,In_1249,In_1889);
xnor U2879 (N_2879,In_2409,In_1186);
nand U2880 (N_2880,In_1776,In_1133);
nor U2881 (N_2881,In_956,In_2092);
or U2882 (N_2882,In_27,In_1303);
nand U2883 (N_2883,In_1225,In_1705);
nor U2884 (N_2884,In_1516,In_1618);
xor U2885 (N_2885,In_510,In_1910);
xnor U2886 (N_2886,In_709,In_50);
xor U2887 (N_2887,In_1612,In_2173);
nand U2888 (N_2888,In_252,In_2224);
nand U2889 (N_2889,In_2052,In_2340);
or U2890 (N_2890,In_472,In_1414);
and U2891 (N_2891,In_2417,In_1302);
or U2892 (N_2892,In_1792,In_230);
and U2893 (N_2893,In_719,In_2375);
nor U2894 (N_2894,In_1762,In_2461);
nand U2895 (N_2895,In_1092,In_2475);
xnor U2896 (N_2896,In_459,In_1966);
nand U2897 (N_2897,In_2047,In_726);
nor U2898 (N_2898,In_1206,In_767);
nor U2899 (N_2899,In_2028,In_293);
and U2900 (N_2900,In_1795,In_1206);
nand U2901 (N_2901,In_387,In_935);
nand U2902 (N_2902,In_490,In_1122);
xor U2903 (N_2903,In_726,In_1447);
nand U2904 (N_2904,In_2423,In_1464);
nor U2905 (N_2905,In_2126,In_2158);
and U2906 (N_2906,In_254,In_2453);
or U2907 (N_2907,In_871,In_1455);
xnor U2908 (N_2908,In_1984,In_1324);
and U2909 (N_2909,In_1837,In_766);
or U2910 (N_2910,In_460,In_273);
nand U2911 (N_2911,In_2238,In_286);
nor U2912 (N_2912,In_1890,In_533);
and U2913 (N_2913,In_2499,In_1860);
nand U2914 (N_2914,In_127,In_769);
or U2915 (N_2915,In_1750,In_271);
or U2916 (N_2916,In_1230,In_943);
or U2917 (N_2917,In_2037,In_50);
nand U2918 (N_2918,In_19,In_510);
nand U2919 (N_2919,In_1945,In_1440);
or U2920 (N_2920,In_2008,In_1255);
or U2921 (N_2921,In_2407,In_2035);
xor U2922 (N_2922,In_893,In_1289);
nor U2923 (N_2923,In_2406,In_538);
nand U2924 (N_2924,In_131,In_1183);
nand U2925 (N_2925,In_366,In_1136);
nand U2926 (N_2926,In_812,In_191);
nor U2927 (N_2927,In_1230,In_919);
xnor U2928 (N_2928,In_1923,In_1455);
or U2929 (N_2929,In_2382,In_1265);
nor U2930 (N_2930,In_1648,In_2014);
and U2931 (N_2931,In_191,In_1702);
or U2932 (N_2932,In_1090,In_1421);
nand U2933 (N_2933,In_2049,In_645);
and U2934 (N_2934,In_389,In_1560);
nand U2935 (N_2935,In_844,In_1657);
and U2936 (N_2936,In_2470,In_239);
xnor U2937 (N_2937,In_215,In_208);
nor U2938 (N_2938,In_1948,In_882);
xor U2939 (N_2939,In_758,In_2198);
xor U2940 (N_2940,In_1794,In_1081);
xnor U2941 (N_2941,In_2055,In_306);
xnor U2942 (N_2942,In_637,In_883);
and U2943 (N_2943,In_145,In_1288);
and U2944 (N_2944,In_2146,In_1729);
nor U2945 (N_2945,In_1601,In_1230);
nor U2946 (N_2946,In_1929,In_1340);
and U2947 (N_2947,In_1003,In_2197);
or U2948 (N_2948,In_1312,In_1551);
nor U2949 (N_2949,In_86,In_403);
nor U2950 (N_2950,In_2292,In_1494);
nand U2951 (N_2951,In_353,In_2179);
or U2952 (N_2952,In_2169,In_339);
xnor U2953 (N_2953,In_2485,In_1573);
nor U2954 (N_2954,In_1273,In_205);
xnor U2955 (N_2955,In_2455,In_1415);
nand U2956 (N_2956,In_1242,In_918);
nor U2957 (N_2957,In_2204,In_1358);
and U2958 (N_2958,In_559,In_1883);
xnor U2959 (N_2959,In_521,In_1104);
nor U2960 (N_2960,In_1424,In_1687);
xor U2961 (N_2961,In_1560,In_1963);
xor U2962 (N_2962,In_1080,In_10);
xor U2963 (N_2963,In_2313,In_1558);
nor U2964 (N_2964,In_1193,In_993);
nor U2965 (N_2965,In_1654,In_614);
nor U2966 (N_2966,In_83,In_1918);
xnor U2967 (N_2967,In_2055,In_751);
and U2968 (N_2968,In_1318,In_699);
and U2969 (N_2969,In_1263,In_442);
nor U2970 (N_2970,In_1633,In_705);
xnor U2971 (N_2971,In_2375,In_913);
nor U2972 (N_2972,In_2343,In_120);
and U2973 (N_2973,In_455,In_788);
and U2974 (N_2974,In_2368,In_2162);
nor U2975 (N_2975,In_1536,In_2098);
xnor U2976 (N_2976,In_444,In_2193);
nor U2977 (N_2977,In_121,In_468);
nand U2978 (N_2978,In_1455,In_1880);
nor U2979 (N_2979,In_1149,In_890);
nand U2980 (N_2980,In_382,In_1709);
nor U2981 (N_2981,In_302,In_1172);
nor U2982 (N_2982,In_1646,In_1492);
nand U2983 (N_2983,In_752,In_1183);
nor U2984 (N_2984,In_1449,In_1901);
nand U2985 (N_2985,In_342,In_1491);
and U2986 (N_2986,In_609,In_514);
and U2987 (N_2987,In_2129,In_2357);
nand U2988 (N_2988,In_867,In_374);
nand U2989 (N_2989,In_575,In_2059);
nor U2990 (N_2990,In_1037,In_765);
nor U2991 (N_2991,In_904,In_2451);
or U2992 (N_2992,In_1079,In_1216);
nor U2993 (N_2993,In_2340,In_1323);
or U2994 (N_2994,In_773,In_621);
or U2995 (N_2995,In_1429,In_1209);
xnor U2996 (N_2996,In_1642,In_124);
and U2997 (N_2997,In_830,In_1668);
and U2998 (N_2998,In_1228,In_2197);
nand U2999 (N_2999,In_395,In_1130);
nand U3000 (N_3000,In_2090,In_1920);
or U3001 (N_3001,In_1869,In_461);
nand U3002 (N_3002,In_127,In_907);
and U3003 (N_3003,In_2164,In_842);
xnor U3004 (N_3004,In_1913,In_335);
and U3005 (N_3005,In_1172,In_750);
nor U3006 (N_3006,In_1660,In_1798);
nor U3007 (N_3007,In_586,In_318);
or U3008 (N_3008,In_12,In_1381);
xnor U3009 (N_3009,In_784,In_842);
nand U3010 (N_3010,In_2154,In_2468);
or U3011 (N_3011,In_1550,In_2424);
xor U3012 (N_3012,In_301,In_323);
and U3013 (N_3013,In_1691,In_1317);
xor U3014 (N_3014,In_1119,In_1520);
nand U3015 (N_3015,In_518,In_751);
nor U3016 (N_3016,In_1139,In_1186);
nand U3017 (N_3017,In_1822,In_528);
and U3018 (N_3018,In_1114,In_1501);
nor U3019 (N_3019,In_1418,In_2023);
xor U3020 (N_3020,In_2199,In_2366);
or U3021 (N_3021,In_1538,In_2205);
nor U3022 (N_3022,In_2120,In_642);
nor U3023 (N_3023,In_1479,In_522);
xor U3024 (N_3024,In_1285,In_2470);
nor U3025 (N_3025,In_1311,In_50);
and U3026 (N_3026,In_2257,In_73);
and U3027 (N_3027,In_1971,In_2178);
xor U3028 (N_3028,In_2449,In_642);
nand U3029 (N_3029,In_17,In_989);
and U3030 (N_3030,In_1990,In_2246);
or U3031 (N_3031,In_288,In_329);
or U3032 (N_3032,In_231,In_1073);
nand U3033 (N_3033,In_892,In_2462);
nor U3034 (N_3034,In_848,In_215);
and U3035 (N_3035,In_2016,In_1191);
nand U3036 (N_3036,In_2087,In_2234);
nor U3037 (N_3037,In_236,In_430);
nor U3038 (N_3038,In_953,In_1398);
nor U3039 (N_3039,In_1597,In_1623);
xor U3040 (N_3040,In_1661,In_889);
or U3041 (N_3041,In_948,In_1382);
and U3042 (N_3042,In_462,In_143);
and U3043 (N_3043,In_2240,In_849);
nor U3044 (N_3044,In_1483,In_261);
and U3045 (N_3045,In_2479,In_1076);
nor U3046 (N_3046,In_71,In_47);
xnor U3047 (N_3047,In_1559,In_1178);
xor U3048 (N_3048,In_111,In_272);
nor U3049 (N_3049,In_1313,In_162);
nor U3050 (N_3050,In_1279,In_707);
or U3051 (N_3051,In_695,In_2457);
xnor U3052 (N_3052,In_754,In_2022);
nor U3053 (N_3053,In_2030,In_1456);
nand U3054 (N_3054,In_1591,In_571);
xor U3055 (N_3055,In_1491,In_2038);
and U3056 (N_3056,In_413,In_313);
xor U3057 (N_3057,In_1880,In_1820);
nor U3058 (N_3058,In_279,In_624);
nor U3059 (N_3059,In_1109,In_872);
xor U3060 (N_3060,In_2445,In_2204);
and U3061 (N_3061,In_1912,In_1436);
xor U3062 (N_3062,In_1462,In_1549);
nand U3063 (N_3063,In_95,In_1660);
and U3064 (N_3064,In_1056,In_1913);
xnor U3065 (N_3065,In_958,In_660);
and U3066 (N_3066,In_2177,In_1439);
and U3067 (N_3067,In_1919,In_1082);
nor U3068 (N_3068,In_2315,In_172);
and U3069 (N_3069,In_526,In_474);
xnor U3070 (N_3070,In_1807,In_1598);
and U3071 (N_3071,In_1181,In_226);
xnor U3072 (N_3072,In_1215,In_125);
xnor U3073 (N_3073,In_1453,In_1421);
or U3074 (N_3074,In_777,In_1377);
and U3075 (N_3075,In_67,In_1268);
nand U3076 (N_3076,In_275,In_740);
nand U3077 (N_3077,In_963,In_2336);
and U3078 (N_3078,In_1602,In_1517);
nand U3079 (N_3079,In_9,In_660);
or U3080 (N_3080,In_1331,In_1275);
xnor U3081 (N_3081,In_1705,In_592);
or U3082 (N_3082,In_315,In_1604);
and U3083 (N_3083,In_1964,In_1541);
xnor U3084 (N_3084,In_1838,In_1551);
nand U3085 (N_3085,In_1495,In_1584);
nand U3086 (N_3086,In_485,In_1900);
and U3087 (N_3087,In_872,In_2491);
nor U3088 (N_3088,In_1918,In_251);
nand U3089 (N_3089,In_1278,In_2084);
nor U3090 (N_3090,In_137,In_758);
xor U3091 (N_3091,In_884,In_1831);
and U3092 (N_3092,In_395,In_233);
or U3093 (N_3093,In_605,In_140);
nor U3094 (N_3094,In_1316,In_494);
nand U3095 (N_3095,In_1083,In_448);
or U3096 (N_3096,In_2453,In_1959);
nand U3097 (N_3097,In_209,In_2389);
xor U3098 (N_3098,In_679,In_1171);
or U3099 (N_3099,In_476,In_1371);
and U3100 (N_3100,In_1806,In_939);
nor U3101 (N_3101,In_2069,In_2112);
xor U3102 (N_3102,In_368,In_1026);
and U3103 (N_3103,In_1852,In_277);
or U3104 (N_3104,In_261,In_1040);
and U3105 (N_3105,In_2107,In_1802);
nor U3106 (N_3106,In_325,In_616);
or U3107 (N_3107,In_252,In_1749);
or U3108 (N_3108,In_2366,In_524);
nor U3109 (N_3109,In_2139,In_1266);
and U3110 (N_3110,In_2251,In_361);
xnor U3111 (N_3111,In_2314,In_362);
xnor U3112 (N_3112,In_183,In_2246);
nor U3113 (N_3113,In_1782,In_526);
or U3114 (N_3114,In_2180,In_2036);
xnor U3115 (N_3115,In_577,In_2010);
xor U3116 (N_3116,In_420,In_0);
and U3117 (N_3117,In_599,In_44);
xor U3118 (N_3118,In_657,In_2442);
nand U3119 (N_3119,In_1866,In_1552);
and U3120 (N_3120,In_179,In_2456);
xnor U3121 (N_3121,In_733,In_1800);
xor U3122 (N_3122,In_767,In_1263);
nand U3123 (N_3123,In_675,In_1938);
xnor U3124 (N_3124,In_1799,In_140);
nand U3125 (N_3125,In_1532,In_794);
and U3126 (N_3126,In_1223,In_458);
nand U3127 (N_3127,In_1483,In_1100);
and U3128 (N_3128,In_308,In_2302);
nor U3129 (N_3129,In_2388,In_2205);
nor U3130 (N_3130,In_245,In_2409);
nand U3131 (N_3131,In_1521,In_780);
and U3132 (N_3132,In_1632,In_1481);
nor U3133 (N_3133,In_329,In_2216);
or U3134 (N_3134,In_864,In_1314);
nand U3135 (N_3135,In_2326,In_2426);
and U3136 (N_3136,In_439,In_393);
nor U3137 (N_3137,In_1612,In_1318);
or U3138 (N_3138,In_1427,In_734);
and U3139 (N_3139,In_1585,In_1678);
and U3140 (N_3140,In_845,In_2099);
or U3141 (N_3141,In_1202,In_132);
and U3142 (N_3142,In_1102,In_1425);
or U3143 (N_3143,In_791,In_1030);
and U3144 (N_3144,In_1966,In_926);
nor U3145 (N_3145,In_471,In_305);
or U3146 (N_3146,In_256,In_1615);
nand U3147 (N_3147,In_371,In_1891);
and U3148 (N_3148,In_877,In_712);
nand U3149 (N_3149,In_809,In_239);
xor U3150 (N_3150,In_2073,In_2158);
or U3151 (N_3151,In_2065,In_2195);
nand U3152 (N_3152,In_559,In_613);
nor U3153 (N_3153,In_899,In_2445);
or U3154 (N_3154,In_1174,In_1484);
and U3155 (N_3155,In_816,In_144);
nor U3156 (N_3156,In_761,In_1227);
nor U3157 (N_3157,In_493,In_716);
nand U3158 (N_3158,In_2190,In_1921);
nor U3159 (N_3159,In_2065,In_2360);
nor U3160 (N_3160,In_447,In_2202);
or U3161 (N_3161,In_1964,In_205);
and U3162 (N_3162,In_1805,In_1456);
or U3163 (N_3163,In_1477,In_1422);
nor U3164 (N_3164,In_1079,In_226);
nor U3165 (N_3165,In_1439,In_1046);
or U3166 (N_3166,In_1842,In_2411);
nand U3167 (N_3167,In_2316,In_516);
nor U3168 (N_3168,In_1135,In_325);
and U3169 (N_3169,In_1540,In_878);
or U3170 (N_3170,In_1615,In_1443);
and U3171 (N_3171,In_2025,In_207);
or U3172 (N_3172,In_404,In_2209);
nor U3173 (N_3173,In_231,In_1715);
xnor U3174 (N_3174,In_628,In_2150);
nor U3175 (N_3175,In_1284,In_716);
nor U3176 (N_3176,In_1171,In_2362);
xor U3177 (N_3177,In_463,In_2425);
nand U3178 (N_3178,In_241,In_2242);
and U3179 (N_3179,In_1314,In_210);
or U3180 (N_3180,In_821,In_539);
and U3181 (N_3181,In_1044,In_1737);
nor U3182 (N_3182,In_2017,In_453);
and U3183 (N_3183,In_2392,In_1302);
and U3184 (N_3184,In_570,In_2329);
nand U3185 (N_3185,In_1208,In_287);
nor U3186 (N_3186,In_570,In_300);
or U3187 (N_3187,In_1220,In_110);
xor U3188 (N_3188,In_829,In_535);
and U3189 (N_3189,In_1864,In_1745);
nor U3190 (N_3190,In_2123,In_1216);
and U3191 (N_3191,In_1494,In_534);
xor U3192 (N_3192,In_2318,In_309);
and U3193 (N_3193,In_2438,In_971);
nand U3194 (N_3194,In_1749,In_572);
xor U3195 (N_3195,In_1482,In_1114);
and U3196 (N_3196,In_174,In_1417);
xnor U3197 (N_3197,In_378,In_1688);
nor U3198 (N_3198,In_1440,In_1678);
and U3199 (N_3199,In_2331,In_1589);
nor U3200 (N_3200,In_1859,In_868);
and U3201 (N_3201,In_1040,In_649);
nor U3202 (N_3202,In_1715,In_1774);
and U3203 (N_3203,In_2163,In_2326);
nor U3204 (N_3204,In_1049,In_1753);
and U3205 (N_3205,In_506,In_2495);
and U3206 (N_3206,In_301,In_599);
and U3207 (N_3207,In_1415,In_1934);
xor U3208 (N_3208,In_1220,In_2455);
nand U3209 (N_3209,In_2285,In_1872);
or U3210 (N_3210,In_968,In_305);
nand U3211 (N_3211,In_377,In_1016);
and U3212 (N_3212,In_260,In_1423);
and U3213 (N_3213,In_659,In_2473);
or U3214 (N_3214,In_967,In_2220);
and U3215 (N_3215,In_110,In_1018);
or U3216 (N_3216,In_1871,In_1985);
xor U3217 (N_3217,In_675,In_655);
xor U3218 (N_3218,In_1886,In_1908);
nand U3219 (N_3219,In_1745,In_1850);
xor U3220 (N_3220,In_689,In_208);
xor U3221 (N_3221,In_1262,In_1506);
nand U3222 (N_3222,In_1628,In_378);
xnor U3223 (N_3223,In_2236,In_509);
nor U3224 (N_3224,In_357,In_2057);
nand U3225 (N_3225,In_990,In_2113);
nor U3226 (N_3226,In_624,In_446);
nand U3227 (N_3227,In_751,In_1563);
and U3228 (N_3228,In_698,In_2085);
nor U3229 (N_3229,In_403,In_51);
nand U3230 (N_3230,In_1849,In_1261);
or U3231 (N_3231,In_1237,In_1791);
or U3232 (N_3232,In_2342,In_1198);
xor U3233 (N_3233,In_1200,In_1199);
xnor U3234 (N_3234,In_2030,In_1552);
or U3235 (N_3235,In_2045,In_1626);
nand U3236 (N_3236,In_1287,In_1884);
or U3237 (N_3237,In_2304,In_1872);
nand U3238 (N_3238,In_1875,In_1054);
or U3239 (N_3239,In_91,In_1743);
xnor U3240 (N_3240,In_1715,In_800);
and U3241 (N_3241,In_1742,In_765);
and U3242 (N_3242,In_667,In_2337);
and U3243 (N_3243,In_1015,In_2357);
xor U3244 (N_3244,In_836,In_296);
and U3245 (N_3245,In_1720,In_379);
or U3246 (N_3246,In_893,In_827);
and U3247 (N_3247,In_593,In_1398);
and U3248 (N_3248,In_503,In_1783);
or U3249 (N_3249,In_2389,In_1641);
nand U3250 (N_3250,In_1055,In_2007);
or U3251 (N_3251,In_1573,In_1775);
nand U3252 (N_3252,In_296,In_1343);
nand U3253 (N_3253,In_1347,In_1152);
nand U3254 (N_3254,In_1791,In_2308);
and U3255 (N_3255,In_584,In_1198);
nor U3256 (N_3256,In_2215,In_2445);
nand U3257 (N_3257,In_783,In_967);
and U3258 (N_3258,In_1090,In_159);
and U3259 (N_3259,In_1081,In_1710);
or U3260 (N_3260,In_2421,In_2069);
xor U3261 (N_3261,In_1173,In_1764);
and U3262 (N_3262,In_2312,In_288);
nand U3263 (N_3263,In_508,In_1610);
nand U3264 (N_3264,In_2255,In_231);
xnor U3265 (N_3265,In_2487,In_1038);
nand U3266 (N_3266,In_1452,In_951);
and U3267 (N_3267,In_2488,In_68);
nor U3268 (N_3268,In_1593,In_2177);
nor U3269 (N_3269,In_1433,In_605);
nand U3270 (N_3270,In_1647,In_2017);
or U3271 (N_3271,In_1094,In_2400);
and U3272 (N_3272,In_311,In_1278);
and U3273 (N_3273,In_1519,In_1820);
or U3274 (N_3274,In_942,In_187);
nor U3275 (N_3275,In_1485,In_895);
nor U3276 (N_3276,In_17,In_777);
or U3277 (N_3277,In_1121,In_2150);
xnor U3278 (N_3278,In_141,In_955);
and U3279 (N_3279,In_1297,In_2444);
xnor U3280 (N_3280,In_1383,In_1247);
xor U3281 (N_3281,In_1474,In_116);
xor U3282 (N_3282,In_694,In_1823);
nor U3283 (N_3283,In_2309,In_1753);
or U3284 (N_3284,In_2163,In_2454);
nand U3285 (N_3285,In_333,In_1975);
and U3286 (N_3286,In_1818,In_1510);
nor U3287 (N_3287,In_300,In_1030);
nor U3288 (N_3288,In_573,In_1235);
xnor U3289 (N_3289,In_2275,In_1036);
or U3290 (N_3290,In_221,In_1566);
nor U3291 (N_3291,In_1177,In_1384);
nand U3292 (N_3292,In_942,In_1436);
xnor U3293 (N_3293,In_2210,In_1664);
nand U3294 (N_3294,In_1262,In_793);
xnor U3295 (N_3295,In_1514,In_810);
nor U3296 (N_3296,In_480,In_1835);
nand U3297 (N_3297,In_1045,In_2490);
xor U3298 (N_3298,In_634,In_2007);
nor U3299 (N_3299,In_701,In_1350);
xor U3300 (N_3300,In_832,In_291);
nand U3301 (N_3301,In_754,In_471);
xnor U3302 (N_3302,In_951,In_1150);
nand U3303 (N_3303,In_1072,In_568);
and U3304 (N_3304,In_307,In_1285);
and U3305 (N_3305,In_811,In_1389);
and U3306 (N_3306,In_257,In_351);
or U3307 (N_3307,In_684,In_1532);
or U3308 (N_3308,In_2340,In_472);
xor U3309 (N_3309,In_867,In_888);
nand U3310 (N_3310,In_1886,In_1810);
and U3311 (N_3311,In_1946,In_1198);
nand U3312 (N_3312,In_1536,In_327);
nor U3313 (N_3313,In_352,In_1103);
nand U3314 (N_3314,In_100,In_859);
xor U3315 (N_3315,In_711,In_2499);
nand U3316 (N_3316,In_2397,In_225);
nor U3317 (N_3317,In_1094,In_1708);
nor U3318 (N_3318,In_1199,In_24);
or U3319 (N_3319,In_101,In_45);
xnor U3320 (N_3320,In_1375,In_498);
or U3321 (N_3321,In_909,In_222);
nand U3322 (N_3322,In_1693,In_1773);
and U3323 (N_3323,In_1513,In_1468);
nand U3324 (N_3324,In_2270,In_118);
xnor U3325 (N_3325,In_2083,In_1495);
xnor U3326 (N_3326,In_513,In_566);
or U3327 (N_3327,In_1152,In_1204);
nand U3328 (N_3328,In_1301,In_315);
nor U3329 (N_3329,In_1268,In_1040);
or U3330 (N_3330,In_420,In_1561);
and U3331 (N_3331,In_464,In_2409);
or U3332 (N_3332,In_1242,In_1997);
and U3333 (N_3333,In_349,In_758);
or U3334 (N_3334,In_1382,In_1987);
or U3335 (N_3335,In_1966,In_64);
nand U3336 (N_3336,In_669,In_1982);
xnor U3337 (N_3337,In_2342,In_137);
nor U3338 (N_3338,In_141,In_286);
or U3339 (N_3339,In_88,In_1039);
nor U3340 (N_3340,In_2215,In_2279);
or U3341 (N_3341,In_817,In_1330);
xor U3342 (N_3342,In_2328,In_2453);
and U3343 (N_3343,In_422,In_286);
and U3344 (N_3344,In_962,In_1535);
nor U3345 (N_3345,In_2127,In_425);
or U3346 (N_3346,In_724,In_1012);
xnor U3347 (N_3347,In_1074,In_767);
nand U3348 (N_3348,In_2052,In_702);
nor U3349 (N_3349,In_1791,In_2078);
and U3350 (N_3350,In_1168,In_1870);
nor U3351 (N_3351,In_1993,In_1996);
and U3352 (N_3352,In_814,In_610);
xor U3353 (N_3353,In_1438,In_1906);
nor U3354 (N_3354,In_862,In_1985);
nand U3355 (N_3355,In_597,In_821);
nor U3356 (N_3356,In_1521,In_1818);
or U3357 (N_3357,In_228,In_1259);
and U3358 (N_3358,In_2001,In_1406);
nand U3359 (N_3359,In_1456,In_1986);
and U3360 (N_3360,In_758,In_1650);
and U3361 (N_3361,In_1989,In_2466);
nor U3362 (N_3362,In_2252,In_2072);
nand U3363 (N_3363,In_1573,In_629);
nor U3364 (N_3364,In_1710,In_764);
and U3365 (N_3365,In_1807,In_1677);
nor U3366 (N_3366,In_2126,In_121);
nand U3367 (N_3367,In_458,In_2147);
nand U3368 (N_3368,In_1580,In_1065);
nor U3369 (N_3369,In_1042,In_813);
and U3370 (N_3370,In_603,In_2262);
or U3371 (N_3371,In_370,In_1441);
xor U3372 (N_3372,In_1907,In_595);
nor U3373 (N_3373,In_1544,In_709);
nor U3374 (N_3374,In_2000,In_101);
xnor U3375 (N_3375,In_1075,In_320);
nand U3376 (N_3376,In_891,In_977);
and U3377 (N_3377,In_1529,In_1761);
or U3378 (N_3378,In_1522,In_1574);
nor U3379 (N_3379,In_973,In_787);
nand U3380 (N_3380,In_1249,In_1471);
and U3381 (N_3381,In_680,In_1726);
and U3382 (N_3382,In_2351,In_684);
and U3383 (N_3383,In_2177,In_2331);
or U3384 (N_3384,In_706,In_1761);
nand U3385 (N_3385,In_2335,In_496);
nand U3386 (N_3386,In_700,In_1205);
and U3387 (N_3387,In_265,In_1784);
nand U3388 (N_3388,In_2127,In_842);
nand U3389 (N_3389,In_705,In_2371);
nor U3390 (N_3390,In_2223,In_352);
xnor U3391 (N_3391,In_542,In_1400);
nand U3392 (N_3392,In_1391,In_1782);
xor U3393 (N_3393,In_2232,In_668);
nand U3394 (N_3394,In_2288,In_1154);
and U3395 (N_3395,In_560,In_2181);
nand U3396 (N_3396,In_1007,In_944);
nand U3397 (N_3397,In_542,In_1722);
xor U3398 (N_3398,In_1761,In_2122);
or U3399 (N_3399,In_1040,In_1785);
and U3400 (N_3400,In_1721,In_972);
xnor U3401 (N_3401,In_1408,In_641);
nand U3402 (N_3402,In_1726,In_331);
and U3403 (N_3403,In_2232,In_2298);
nand U3404 (N_3404,In_2046,In_1162);
nand U3405 (N_3405,In_1100,In_1582);
xor U3406 (N_3406,In_1747,In_893);
nor U3407 (N_3407,In_2337,In_1199);
nor U3408 (N_3408,In_481,In_964);
xnor U3409 (N_3409,In_2283,In_1208);
xor U3410 (N_3410,In_244,In_452);
xor U3411 (N_3411,In_2403,In_1226);
or U3412 (N_3412,In_1945,In_849);
and U3413 (N_3413,In_256,In_121);
or U3414 (N_3414,In_1196,In_1493);
nand U3415 (N_3415,In_39,In_643);
nor U3416 (N_3416,In_613,In_1462);
and U3417 (N_3417,In_923,In_140);
xnor U3418 (N_3418,In_724,In_1788);
nor U3419 (N_3419,In_1383,In_699);
or U3420 (N_3420,In_2425,In_925);
xnor U3421 (N_3421,In_1052,In_1656);
nand U3422 (N_3422,In_1951,In_951);
and U3423 (N_3423,In_2033,In_2115);
and U3424 (N_3424,In_531,In_1190);
xor U3425 (N_3425,In_1779,In_1935);
nor U3426 (N_3426,In_1190,In_568);
xor U3427 (N_3427,In_1120,In_2177);
or U3428 (N_3428,In_432,In_1393);
nor U3429 (N_3429,In_455,In_2023);
nand U3430 (N_3430,In_2235,In_1231);
nor U3431 (N_3431,In_2491,In_39);
nand U3432 (N_3432,In_1790,In_2361);
or U3433 (N_3433,In_401,In_531);
or U3434 (N_3434,In_2219,In_289);
xor U3435 (N_3435,In_2190,In_978);
nor U3436 (N_3436,In_2489,In_1972);
or U3437 (N_3437,In_1778,In_1691);
nor U3438 (N_3438,In_894,In_147);
nand U3439 (N_3439,In_863,In_748);
nor U3440 (N_3440,In_2364,In_1602);
nor U3441 (N_3441,In_1405,In_1134);
and U3442 (N_3442,In_1184,In_1340);
nand U3443 (N_3443,In_1421,In_1473);
nor U3444 (N_3444,In_224,In_1354);
nand U3445 (N_3445,In_1122,In_329);
nor U3446 (N_3446,In_1040,In_617);
nand U3447 (N_3447,In_1147,In_1704);
nor U3448 (N_3448,In_658,In_2084);
nand U3449 (N_3449,In_1096,In_1278);
xnor U3450 (N_3450,In_1991,In_670);
and U3451 (N_3451,In_254,In_2181);
nand U3452 (N_3452,In_277,In_1325);
nor U3453 (N_3453,In_1613,In_2453);
nor U3454 (N_3454,In_2322,In_2202);
or U3455 (N_3455,In_326,In_605);
xnor U3456 (N_3456,In_1810,In_163);
and U3457 (N_3457,In_2378,In_1506);
nand U3458 (N_3458,In_1202,In_2255);
xnor U3459 (N_3459,In_260,In_1034);
nand U3460 (N_3460,In_63,In_2413);
xnor U3461 (N_3461,In_1855,In_758);
xor U3462 (N_3462,In_2072,In_1843);
or U3463 (N_3463,In_450,In_2065);
xor U3464 (N_3464,In_2310,In_1369);
or U3465 (N_3465,In_2106,In_792);
or U3466 (N_3466,In_411,In_1001);
xnor U3467 (N_3467,In_2475,In_1305);
nor U3468 (N_3468,In_1464,In_89);
and U3469 (N_3469,In_1524,In_684);
and U3470 (N_3470,In_643,In_190);
xor U3471 (N_3471,In_1242,In_351);
or U3472 (N_3472,In_1251,In_121);
or U3473 (N_3473,In_620,In_1947);
and U3474 (N_3474,In_2293,In_656);
nand U3475 (N_3475,In_1037,In_116);
nor U3476 (N_3476,In_2076,In_870);
and U3477 (N_3477,In_654,In_277);
and U3478 (N_3478,In_2335,In_933);
nand U3479 (N_3479,In_2307,In_157);
nor U3480 (N_3480,In_897,In_1016);
xor U3481 (N_3481,In_572,In_1549);
nor U3482 (N_3482,In_402,In_954);
or U3483 (N_3483,In_2373,In_299);
and U3484 (N_3484,In_1671,In_1265);
xor U3485 (N_3485,In_579,In_138);
nor U3486 (N_3486,In_1681,In_2297);
nor U3487 (N_3487,In_1192,In_1057);
or U3488 (N_3488,In_1448,In_594);
and U3489 (N_3489,In_47,In_644);
and U3490 (N_3490,In_1330,In_1835);
nand U3491 (N_3491,In_1473,In_703);
nor U3492 (N_3492,In_2360,In_2044);
nand U3493 (N_3493,In_1112,In_2394);
nand U3494 (N_3494,In_513,In_743);
xor U3495 (N_3495,In_1589,In_1145);
xnor U3496 (N_3496,In_1608,In_820);
xnor U3497 (N_3497,In_2263,In_451);
nor U3498 (N_3498,In_1697,In_41);
nand U3499 (N_3499,In_156,In_1837);
nand U3500 (N_3500,In_2255,In_410);
or U3501 (N_3501,In_1515,In_1949);
nand U3502 (N_3502,In_993,In_19);
nand U3503 (N_3503,In_2087,In_1742);
nor U3504 (N_3504,In_941,In_1883);
nand U3505 (N_3505,In_2124,In_1275);
xnor U3506 (N_3506,In_335,In_904);
or U3507 (N_3507,In_1873,In_119);
nand U3508 (N_3508,In_1077,In_2075);
xnor U3509 (N_3509,In_2045,In_97);
nor U3510 (N_3510,In_2240,In_1250);
nand U3511 (N_3511,In_384,In_1669);
nand U3512 (N_3512,In_499,In_2043);
nor U3513 (N_3513,In_2066,In_954);
nand U3514 (N_3514,In_2221,In_874);
nor U3515 (N_3515,In_1333,In_76);
xnor U3516 (N_3516,In_669,In_1259);
xnor U3517 (N_3517,In_1801,In_1985);
and U3518 (N_3518,In_1903,In_1312);
nor U3519 (N_3519,In_40,In_1357);
nor U3520 (N_3520,In_2153,In_579);
or U3521 (N_3521,In_1416,In_596);
and U3522 (N_3522,In_1588,In_951);
or U3523 (N_3523,In_1611,In_1567);
and U3524 (N_3524,In_261,In_1853);
and U3525 (N_3525,In_781,In_1268);
nor U3526 (N_3526,In_91,In_579);
xnor U3527 (N_3527,In_2231,In_1912);
nor U3528 (N_3528,In_1550,In_663);
nand U3529 (N_3529,In_347,In_2120);
nand U3530 (N_3530,In_1583,In_864);
xor U3531 (N_3531,In_2091,In_2353);
nor U3532 (N_3532,In_2232,In_1306);
nand U3533 (N_3533,In_950,In_2314);
and U3534 (N_3534,In_2370,In_121);
xor U3535 (N_3535,In_2136,In_525);
xnor U3536 (N_3536,In_1048,In_1440);
xnor U3537 (N_3537,In_1921,In_2418);
nor U3538 (N_3538,In_1163,In_109);
or U3539 (N_3539,In_1090,In_1069);
nor U3540 (N_3540,In_1973,In_1254);
and U3541 (N_3541,In_2196,In_424);
nor U3542 (N_3542,In_388,In_1967);
or U3543 (N_3543,In_2276,In_873);
and U3544 (N_3544,In_1027,In_615);
nor U3545 (N_3545,In_1392,In_2291);
nor U3546 (N_3546,In_2414,In_1176);
nor U3547 (N_3547,In_498,In_404);
nor U3548 (N_3548,In_1214,In_1333);
xnor U3549 (N_3549,In_2488,In_313);
nor U3550 (N_3550,In_2137,In_1551);
nand U3551 (N_3551,In_1957,In_357);
nand U3552 (N_3552,In_2211,In_2075);
and U3553 (N_3553,In_691,In_718);
or U3554 (N_3554,In_917,In_1457);
xor U3555 (N_3555,In_2230,In_1531);
nand U3556 (N_3556,In_2230,In_2236);
nand U3557 (N_3557,In_2316,In_1263);
nand U3558 (N_3558,In_702,In_2151);
nand U3559 (N_3559,In_205,In_1695);
nor U3560 (N_3560,In_2437,In_1115);
xor U3561 (N_3561,In_1839,In_1382);
nand U3562 (N_3562,In_11,In_2440);
nor U3563 (N_3563,In_798,In_661);
and U3564 (N_3564,In_502,In_1322);
xor U3565 (N_3565,In_1266,In_470);
xor U3566 (N_3566,In_558,In_210);
or U3567 (N_3567,In_1823,In_1608);
nand U3568 (N_3568,In_246,In_1687);
nand U3569 (N_3569,In_1481,In_1170);
nor U3570 (N_3570,In_241,In_1360);
nor U3571 (N_3571,In_1533,In_1510);
or U3572 (N_3572,In_1335,In_368);
nor U3573 (N_3573,In_1708,In_881);
or U3574 (N_3574,In_418,In_664);
xnor U3575 (N_3575,In_670,In_199);
and U3576 (N_3576,In_1565,In_1059);
or U3577 (N_3577,In_1676,In_2087);
nor U3578 (N_3578,In_1206,In_206);
xnor U3579 (N_3579,In_1764,In_254);
and U3580 (N_3580,In_2450,In_2436);
or U3581 (N_3581,In_657,In_2208);
or U3582 (N_3582,In_2060,In_1130);
xor U3583 (N_3583,In_171,In_425);
nand U3584 (N_3584,In_1960,In_1699);
xnor U3585 (N_3585,In_1517,In_1450);
nand U3586 (N_3586,In_2486,In_1560);
and U3587 (N_3587,In_1315,In_1411);
nand U3588 (N_3588,In_1979,In_2321);
nand U3589 (N_3589,In_1942,In_1927);
and U3590 (N_3590,In_2092,In_354);
or U3591 (N_3591,In_1993,In_284);
nand U3592 (N_3592,In_277,In_2347);
or U3593 (N_3593,In_2086,In_1325);
nand U3594 (N_3594,In_1805,In_1698);
nor U3595 (N_3595,In_1705,In_1169);
and U3596 (N_3596,In_2006,In_2368);
nor U3597 (N_3597,In_357,In_2373);
nand U3598 (N_3598,In_2460,In_953);
xnor U3599 (N_3599,In_297,In_1768);
nor U3600 (N_3600,In_1783,In_389);
or U3601 (N_3601,In_171,In_26);
and U3602 (N_3602,In_1410,In_1245);
and U3603 (N_3603,In_1898,In_277);
and U3604 (N_3604,In_1482,In_352);
nand U3605 (N_3605,In_345,In_1136);
nor U3606 (N_3606,In_656,In_502);
or U3607 (N_3607,In_1549,In_1725);
nand U3608 (N_3608,In_705,In_750);
and U3609 (N_3609,In_1914,In_451);
xor U3610 (N_3610,In_1512,In_989);
and U3611 (N_3611,In_2384,In_1139);
nand U3612 (N_3612,In_1013,In_1863);
or U3613 (N_3613,In_2216,In_659);
xnor U3614 (N_3614,In_175,In_200);
nor U3615 (N_3615,In_1007,In_290);
and U3616 (N_3616,In_160,In_1278);
xor U3617 (N_3617,In_1035,In_1628);
nor U3618 (N_3618,In_1424,In_1932);
nor U3619 (N_3619,In_1416,In_1082);
nand U3620 (N_3620,In_2440,In_1407);
nand U3621 (N_3621,In_2116,In_1673);
or U3622 (N_3622,In_18,In_313);
and U3623 (N_3623,In_1065,In_877);
xnor U3624 (N_3624,In_1511,In_190);
nand U3625 (N_3625,In_614,In_1139);
nand U3626 (N_3626,In_619,In_379);
and U3627 (N_3627,In_97,In_2288);
xnor U3628 (N_3628,In_1908,In_366);
nand U3629 (N_3629,In_915,In_518);
nor U3630 (N_3630,In_2116,In_233);
or U3631 (N_3631,In_1303,In_2067);
nand U3632 (N_3632,In_2026,In_226);
nor U3633 (N_3633,In_2251,In_1591);
xnor U3634 (N_3634,In_449,In_10);
or U3635 (N_3635,In_2038,In_1367);
xor U3636 (N_3636,In_752,In_1749);
nand U3637 (N_3637,In_2490,In_380);
and U3638 (N_3638,In_1093,In_2438);
and U3639 (N_3639,In_895,In_2061);
xnor U3640 (N_3640,In_536,In_1392);
nor U3641 (N_3641,In_1034,In_709);
and U3642 (N_3642,In_2375,In_2279);
xnor U3643 (N_3643,In_1888,In_967);
xnor U3644 (N_3644,In_1716,In_765);
nor U3645 (N_3645,In_1713,In_1948);
and U3646 (N_3646,In_2136,In_1542);
or U3647 (N_3647,In_1314,In_660);
xnor U3648 (N_3648,In_2429,In_624);
and U3649 (N_3649,In_141,In_354);
xnor U3650 (N_3650,In_2185,In_295);
xnor U3651 (N_3651,In_45,In_1411);
and U3652 (N_3652,In_351,In_1868);
xnor U3653 (N_3653,In_153,In_72);
or U3654 (N_3654,In_1431,In_311);
nor U3655 (N_3655,In_1995,In_2467);
nor U3656 (N_3656,In_139,In_219);
and U3657 (N_3657,In_450,In_2351);
or U3658 (N_3658,In_647,In_1383);
xor U3659 (N_3659,In_1726,In_2077);
and U3660 (N_3660,In_1652,In_2462);
nor U3661 (N_3661,In_57,In_601);
xnor U3662 (N_3662,In_384,In_1122);
and U3663 (N_3663,In_348,In_1730);
nor U3664 (N_3664,In_1676,In_972);
nand U3665 (N_3665,In_1159,In_236);
nor U3666 (N_3666,In_644,In_335);
xor U3667 (N_3667,In_721,In_2109);
xor U3668 (N_3668,In_1522,In_735);
and U3669 (N_3669,In_1212,In_1838);
nor U3670 (N_3670,In_2202,In_76);
and U3671 (N_3671,In_2279,In_1111);
nor U3672 (N_3672,In_184,In_681);
or U3673 (N_3673,In_2042,In_1868);
and U3674 (N_3674,In_1974,In_949);
xnor U3675 (N_3675,In_2254,In_688);
xor U3676 (N_3676,In_1626,In_508);
and U3677 (N_3677,In_492,In_769);
or U3678 (N_3678,In_57,In_202);
and U3679 (N_3679,In_907,In_654);
and U3680 (N_3680,In_2199,In_1611);
and U3681 (N_3681,In_530,In_141);
xor U3682 (N_3682,In_400,In_2429);
or U3683 (N_3683,In_647,In_1105);
nand U3684 (N_3684,In_417,In_2431);
nor U3685 (N_3685,In_528,In_1421);
nand U3686 (N_3686,In_143,In_558);
and U3687 (N_3687,In_1600,In_1666);
and U3688 (N_3688,In_973,In_1550);
nor U3689 (N_3689,In_1340,In_1457);
nor U3690 (N_3690,In_864,In_2460);
nand U3691 (N_3691,In_1632,In_1262);
xnor U3692 (N_3692,In_155,In_1393);
nor U3693 (N_3693,In_2060,In_1516);
nand U3694 (N_3694,In_942,In_1615);
and U3695 (N_3695,In_2161,In_1858);
xor U3696 (N_3696,In_1769,In_687);
nor U3697 (N_3697,In_2008,In_331);
and U3698 (N_3698,In_2300,In_1779);
or U3699 (N_3699,In_1899,In_1900);
nand U3700 (N_3700,In_429,In_1809);
and U3701 (N_3701,In_88,In_1539);
and U3702 (N_3702,In_1182,In_1394);
nor U3703 (N_3703,In_1704,In_2157);
or U3704 (N_3704,In_1703,In_1941);
and U3705 (N_3705,In_2266,In_2458);
nand U3706 (N_3706,In_2313,In_2022);
nor U3707 (N_3707,In_2326,In_1400);
and U3708 (N_3708,In_1227,In_1919);
nor U3709 (N_3709,In_517,In_2346);
or U3710 (N_3710,In_1112,In_2185);
xor U3711 (N_3711,In_469,In_1074);
xor U3712 (N_3712,In_1163,In_2421);
nor U3713 (N_3713,In_1085,In_1266);
nand U3714 (N_3714,In_547,In_1128);
xor U3715 (N_3715,In_1267,In_1994);
or U3716 (N_3716,In_1389,In_509);
nor U3717 (N_3717,In_2206,In_31);
and U3718 (N_3718,In_322,In_2391);
nand U3719 (N_3719,In_1591,In_1351);
xnor U3720 (N_3720,In_2209,In_827);
nand U3721 (N_3721,In_769,In_1518);
or U3722 (N_3722,In_2327,In_1038);
xor U3723 (N_3723,In_399,In_1252);
or U3724 (N_3724,In_873,In_1917);
and U3725 (N_3725,In_70,In_289);
xor U3726 (N_3726,In_1564,In_1860);
xor U3727 (N_3727,In_1310,In_1047);
nand U3728 (N_3728,In_1969,In_180);
and U3729 (N_3729,In_2306,In_416);
xor U3730 (N_3730,In_1700,In_967);
or U3731 (N_3731,In_1273,In_925);
or U3732 (N_3732,In_2039,In_279);
nand U3733 (N_3733,In_697,In_2050);
xnor U3734 (N_3734,In_589,In_463);
nor U3735 (N_3735,In_112,In_614);
xor U3736 (N_3736,In_417,In_986);
xnor U3737 (N_3737,In_534,In_1448);
xnor U3738 (N_3738,In_1575,In_347);
nor U3739 (N_3739,In_721,In_45);
and U3740 (N_3740,In_2475,In_1259);
or U3741 (N_3741,In_2261,In_1982);
xnor U3742 (N_3742,In_674,In_1689);
nor U3743 (N_3743,In_1060,In_2151);
xor U3744 (N_3744,In_2212,In_1933);
xor U3745 (N_3745,In_1652,In_200);
or U3746 (N_3746,In_839,In_2268);
or U3747 (N_3747,In_1128,In_1690);
xor U3748 (N_3748,In_2335,In_103);
nand U3749 (N_3749,In_911,In_1584);
and U3750 (N_3750,In_1687,In_503);
nand U3751 (N_3751,In_272,In_23);
or U3752 (N_3752,In_155,In_1143);
and U3753 (N_3753,In_1946,In_2263);
nor U3754 (N_3754,In_666,In_1189);
nor U3755 (N_3755,In_1476,In_221);
nand U3756 (N_3756,In_1892,In_1322);
nor U3757 (N_3757,In_1130,In_1958);
xnor U3758 (N_3758,In_1751,In_1446);
and U3759 (N_3759,In_747,In_475);
or U3760 (N_3760,In_1557,In_161);
nor U3761 (N_3761,In_1968,In_1230);
or U3762 (N_3762,In_98,In_883);
nand U3763 (N_3763,In_2124,In_105);
or U3764 (N_3764,In_260,In_1902);
and U3765 (N_3765,In_1109,In_1998);
and U3766 (N_3766,In_2185,In_1642);
nand U3767 (N_3767,In_556,In_87);
nor U3768 (N_3768,In_1118,In_2369);
and U3769 (N_3769,In_1543,In_1715);
xor U3770 (N_3770,In_2402,In_1996);
or U3771 (N_3771,In_1466,In_1027);
nor U3772 (N_3772,In_1529,In_972);
xnor U3773 (N_3773,In_2014,In_2409);
nor U3774 (N_3774,In_443,In_561);
and U3775 (N_3775,In_371,In_1306);
xnor U3776 (N_3776,In_442,In_62);
xor U3777 (N_3777,In_973,In_47);
and U3778 (N_3778,In_1733,In_2445);
and U3779 (N_3779,In_1343,In_1512);
or U3780 (N_3780,In_1742,In_2012);
nand U3781 (N_3781,In_540,In_878);
xnor U3782 (N_3782,In_1775,In_1402);
xor U3783 (N_3783,In_676,In_606);
or U3784 (N_3784,In_610,In_2301);
and U3785 (N_3785,In_1606,In_1068);
and U3786 (N_3786,In_811,In_2221);
or U3787 (N_3787,In_1101,In_2121);
or U3788 (N_3788,In_2330,In_663);
xor U3789 (N_3789,In_800,In_751);
nor U3790 (N_3790,In_1268,In_2138);
or U3791 (N_3791,In_1426,In_1422);
or U3792 (N_3792,In_87,In_261);
or U3793 (N_3793,In_325,In_67);
nor U3794 (N_3794,In_558,In_683);
nand U3795 (N_3795,In_1117,In_1345);
nand U3796 (N_3796,In_2166,In_2433);
nand U3797 (N_3797,In_686,In_809);
xnor U3798 (N_3798,In_1457,In_1522);
xnor U3799 (N_3799,In_1970,In_2036);
and U3800 (N_3800,In_1217,In_2144);
xnor U3801 (N_3801,In_1348,In_1412);
nor U3802 (N_3802,In_927,In_1647);
or U3803 (N_3803,In_1944,In_218);
and U3804 (N_3804,In_343,In_2359);
nor U3805 (N_3805,In_77,In_1336);
nor U3806 (N_3806,In_450,In_2399);
and U3807 (N_3807,In_2083,In_333);
nand U3808 (N_3808,In_158,In_553);
nand U3809 (N_3809,In_1640,In_2085);
nand U3810 (N_3810,In_602,In_959);
nand U3811 (N_3811,In_899,In_204);
nand U3812 (N_3812,In_1088,In_2169);
xor U3813 (N_3813,In_1918,In_444);
or U3814 (N_3814,In_542,In_1072);
or U3815 (N_3815,In_1723,In_1453);
nand U3816 (N_3816,In_2193,In_68);
nand U3817 (N_3817,In_575,In_2056);
nor U3818 (N_3818,In_2380,In_2427);
xnor U3819 (N_3819,In_955,In_1654);
nor U3820 (N_3820,In_625,In_306);
nor U3821 (N_3821,In_941,In_1630);
nand U3822 (N_3822,In_1276,In_126);
nor U3823 (N_3823,In_691,In_209);
and U3824 (N_3824,In_907,In_265);
nand U3825 (N_3825,In_1362,In_901);
or U3826 (N_3826,In_859,In_2492);
nor U3827 (N_3827,In_1071,In_915);
or U3828 (N_3828,In_699,In_2174);
nand U3829 (N_3829,In_691,In_82);
xor U3830 (N_3830,In_843,In_926);
and U3831 (N_3831,In_1848,In_1681);
and U3832 (N_3832,In_1769,In_2273);
xor U3833 (N_3833,In_783,In_950);
nand U3834 (N_3834,In_699,In_1158);
nand U3835 (N_3835,In_778,In_2001);
or U3836 (N_3836,In_1408,In_404);
nor U3837 (N_3837,In_1936,In_290);
xor U3838 (N_3838,In_647,In_934);
xor U3839 (N_3839,In_1352,In_875);
xor U3840 (N_3840,In_897,In_208);
and U3841 (N_3841,In_588,In_30);
or U3842 (N_3842,In_213,In_835);
nor U3843 (N_3843,In_201,In_116);
and U3844 (N_3844,In_261,In_35);
nand U3845 (N_3845,In_2289,In_1214);
xor U3846 (N_3846,In_2304,In_466);
nor U3847 (N_3847,In_225,In_547);
and U3848 (N_3848,In_1489,In_1209);
nand U3849 (N_3849,In_706,In_243);
nor U3850 (N_3850,In_2384,In_1743);
or U3851 (N_3851,In_934,In_2098);
and U3852 (N_3852,In_802,In_890);
and U3853 (N_3853,In_1237,In_2206);
nand U3854 (N_3854,In_1729,In_544);
nor U3855 (N_3855,In_1576,In_2252);
and U3856 (N_3856,In_352,In_36);
nand U3857 (N_3857,In_2309,In_2280);
nand U3858 (N_3858,In_420,In_1498);
and U3859 (N_3859,In_392,In_1528);
and U3860 (N_3860,In_1737,In_292);
or U3861 (N_3861,In_487,In_690);
and U3862 (N_3862,In_2256,In_309);
and U3863 (N_3863,In_1374,In_942);
or U3864 (N_3864,In_2486,In_2066);
xnor U3865 (N_3865,In_2051,In_188);
and U3866 (N_3866,In_2123,In_2113);
xnor U3867 (N_3867,In_468,In_1366);
xnor U3868 (N_3868,In_709,In_2148);
nand U3869 (N_3869,In_1635,In_1671);
or U3870 (N_3870,In_396,In_1760);
and U3871 (N_3871,In_1748,In_2209);
or U3872 (N_3872,In_1127,In_1899);
or U3873 (N_3873,In_1087,In_1366);
xor U3874 (N_3874,In_392,In_1411);
and U3875 (N_3875,In_854,In_1723);
nor U3876 (N_3876,In_2044,In_279);
or U3877 (N_3877,In_1671,In_1372);
or U3878 (N_3878,In_1431,In_597);
nand U3879 (N_3879,In_2070,In_2204);
nand U3880 (N_3880,In_403,In_1314);
or U3881 (N_3881,In_1024,In_2007);
nor U3882 (N_3882,In_181,In_1525);
or U3883 (N_3883,In_1881,In_312);
nor U3884 (N_3884,In_888,In_1666);
and U3885 (N_3885,In_1560,In_523);
xnor U3886 (N_3886,In_387,In_899);
xnor U3887 (N_3887,In_1267,In_464);
xor U3888 (N_3888,In_588,In_1841);
or U3889 (N_3889,In_1455,In_1238);
and U3890 (N_3890,In_1828,In_806);
nand U3891 (N_3891,In_2186,In_716);
or U3892 (N_3892,In_2208,In_2252);
nor U3893 (N_3893,In_364,In_2239);
and U3894 (N_3894,In_74,In_698);
xnor U3895 (N_3895,In_878,In_2341);
nand U3896 (N_3896,In_1713,In_253);
or U3897 (N_3897,In_1946,In_410);
nand U3898 (N_3898,In_1410,In_1352);
nor U3899 (N_3899,In_216,In_1433);
nand U3900 (N_3900,In_137,In_1418);
nor U3901 (N_3901,In_1736,In_2042);
nor U3902 (N_3902,In_407,In_2035);
nand U3903 (N_3903,In_2477,In_997);
and U3904 (N_3904,In_1108,In_1085);
or U3905 (N_3905,In_2283,In_2173);
and U3906 (N_3906,In_400,In_1298);
or U3907 (N_3907,In_1943,In_2313);
nand U3908 (N_3908,In_949,In_891);
nor U3909 (N_3909,In_14,In_1310);
or U3910 (N_3910,In_2264,In_1700);
nor U3911 (N_3911,In_349,In_2199);
and U3912 (N_3912,In_2447,In_360);
xnor U3913 (N_3913,In_6,In_1125);
xnor U3914 (N_3914,In_84,In_146);
and U3915 (N_3915,In_228,In_823);
xnor U3916 (N_3916,In_1717,In_1561);
and U3917 (N_3917,In_2413,In_1448);
and U3918 (N_3918,In_1782,In_2114);
xnor U3919 (N_3919,In_2042,In_1867);
xor U3920 (N_3920,In_1294,In_2485);
or U3921 (N_3921,In_152,In_987);
nand U3922 (N_3922,In_773,In_417);
nand U3923 (N_3923,In_1894,In_1681);
nor U3924 (N_3924,In_2317,In_1104);
xor U3925 (N_3925,In_167,In_1785);
nor U3926 (N_3926,In_1998,In_2340);
and U3927 (N_3927,In_264,In_2207);
nor U3928 (N_3928,In_311,In_708);
nand U3929 (N_3929,In_638,In_1178);
xor U3930 (N_3930,In_1925,In_2104);
and U3931 (N_3931,In_613,In_1583);
xor U3932 (N_3932,In_406,In_834);
or U3933 (N_3933,In_217,In_530);
xor U3934 (N_3934,In_723,In_1303);
nand U3935 (N_3935,In_1094,In_1858);
nor U3936 (N_3936,In_2293,In_1089);
nor U3937 (N_3937,In_2379,In_1263);
nand U3938 (N_3938,In_2103,In_1590);
or U3939 (N_3939,In_1164,In_793);
or U3940 (N_3940,In_1410,In_460);
or U3941 (N_3941,In_2481,In_1936);
and U3942 (N_3942,In_1276,In_967);
xor U3943 (N_3943,In_1384,In_2180);
and U3944 (N_3944,In_1755,In_115);
nor U3945 (N_3945,In_158,In_585);
and U3946 (N_3946,In_2433,In_751);
nand U3947 (N_3947,In_1622,In_2158);
nand U3948 (N_3948,In_1942,In_2128);
nand U3949 (N_3949,In_1330,In_314);
and U3950 (N_3950,In_1687,In_536);
nand U3951 (N_3951,In_521,In_1699);
or U3952 (N_3952,In_846,In_484);
or U3953 (N_3953,In_939,In_167);
nor U3954 (N_3954,In_543,In_1996);
xor U3955 (N_3955,In_1063,In_2213);
nand U3956 (N_3956,In_1465,In_2269);
xor U3957 (N_3957,In_1614,In_589);
or U3958 (N_3958,In_1167,In_1345);
xnor U3959 (N_3959,In_341,In_1172);
and U3960 (N_3960,In_669,In_1180);
nor U3961 (N_3961,In_2422,In_1170);
xor U3962 (N_3962,In_1525,In_1937);
nor U3963 (N_3963,In_193,In_1200);
xnor U3964 (N_3964,In_773,In_1113);
nor U3965 (N_3965,In_807,In_785);
xor U3966 (N_3966,In_66,In_256);
nor U3967 (N_3967,In_925,In_1576);
nand U3968 (N_3968,In_1004,In_1149);
xor U3969 (N_3969,In_554,In_1883);
or U3970 (N_3970,In_157,In_2350);
or U3971 (N_3971,In_395,In_2345);
and U3972 (N_3972,In_500,In_285);
nand U3973 (N_3973,In_641,In_1665);
xnor U3974 (N_3974,In_1861,In_2396);
nand U3975 (N_3975,In_158,In_957);
nor U3976 (N_3976,In_1036,In_2418);
nor U3977 (N_3977,In_1016,In_677);
or U3978 (N_3978,In_2350,In_245);
nor U3979 (N_3979,In_1793,In_645);
nand U3980 (N_3980,In_2082,In_1740);
or U3981 (N_3981,In_1245,In_1825);
nor U3982 (N_3982,In_675,In_1567);
or U3983 (N_3983,In_2051,In_1636);
nor U3984 (N_3984,In_605,In_405);
xnor U3985 (N_3985,In_1786,In_1813);
nand U3986 (N_3986,In_604,In_799);
or U3987 (N_3987,In_1371,In_1398);
nand U3988 (N_3988,In_516,In_913);
nor U3989 (N_3989,In_2366,In_1472);
nor U3990 (N_3990,In_1511,In_343);
and U3991 (N_3991,In_1824,In_1076);
nand U3992 (N_3992,In_512,In_1123);
nor U3993 (N_3993,In_1221,In_562);
nand U3994 (N_3994,In_612,In_471);
and U3995 (N_3995,In_1341,In_1709);
xnor U3996 (N_3996,In_1323,In_865);
and U3997 (N_3997,In_923,In_317);
xnor U3998 (N_3998,In_2378,In_817);
and U3999 (N_3999,In_638,In_1288);
xor U4000 (N_4000,In_1848,In_33);
and U4001 (N_4001,In_111,In_1428);
and U4002 (N_4002,In_1429,In_402);
nand U4003 (N_4003,In_471,In_289);
or U4004 (N_4004,In_2149,In_958);
nand U4005 (N_4005,In_2009,In_1119);
and U4006 (N_4006,In_2166,In_1553);
or U4007 (N_4007,In_779,In_121);
and U4008 (N_4008,In_589,In_253);
nand U4009 (N_4009,In_2084,In_2188);
and U4010 (N_4010,In_1076,In_2208);
nor U4011 (N_4011,In_128,In_1455);
nor U4012 (N_4012,In_697,In_278);
and U4013 (N_4013,In_2397,In_204);
nand U4014 (N_4014,In_2328,In_819);
nor U4015 (N_4015,In_1175,In_153);
or U4016 (N_4016,In_907,In_194);
and U4017 (N_4017,In_407,In_8);
xnor U4018 (N_4018,In_1880,In_1265);
xnor U4019 (N_4019,In_29,In_1086);
or U4020 (N_4020,In_528,In_178);
and U4021 (N_4021,In_2070,In_360);
and U4022 (N_4022,In_125,In_1323);
nand U4023 (N_4023,In_622,In_677);
nor U4024 (N_4024,In_420,In_332);
nor U4025 (N_4025,In_623,In_1990);
nor U4026 (N_4026,In_131,In_1341);
and U4027 (N_4027,In_2437,In_2261);
or U4028 (N_4028,In_1037,In_1234);
nor U4029 (N_4029,In_900,In_128);
xnor U4030 (N_4030,In_1812,In_91);
nand U4031 (N_4031,In_1525,In_1513);
and U4032 (N_4032,In_565,In_564);
nor U4033 (N_4033,In_681,In_1879);
and U4034 (N_4034,In_104,In_1831);
nand U4035 (N_4035,In_652,In_587);
and U4036 (N_4036,In_1094,In_81);
xnor U4037 (N_4037,In_1460,In_2164);
or U4038 (N_4038,In_192,In_1694);
nand U4039 (N_4039,In_574,In_768);
nand U4040 (N_4040,In_1842,In_2484);
nand U4041 (N_4041,In_2158,In_2174);
xor U4042 (N_4042,In_2072,In_1146);
nor U4043 (N_4043,In_1507,In_1240);
nor U4044 (N_4044,In_612,In_1012);
nor U4045 (N_4045,In_1799,In_235);
and U4046 (N_4046,In_1806,In_2450);
or U4047 (N_4047,In_132,In_413);
and U4048 (N_4048,In_2101,In_155);
xnor U4049 (N_4049,In_496,In_362);
nor U4050 (N_4050,In_1665,In_248);
nor U4051 (N_4051,In_149,In_992);
nor U4052 (N_4052,In_2426,In_2211);
nand U4053 (N_4053,In_1089,In_608);
and U4054 (N_4054,In_2477,In_566);
nor U4055 (N_4055,In_1132,In_684);
nand U4056 (N_4056,In_2027,In_1510);
xnor U4057 (N_4057,In_775,In_792);
and U4058 (N_4058,In_1618,In_306);
nor U4059 (N_4059,In_139,In_626);
and U4060 (N_4060,In_410,In_527);
or U4061 (N_4061,In_2264,In_1224);
or U4062 (N_4062,In_927,In_2465);
or U4063 (N_4063,In_442,In_1443);
nand U4064 (N_4064,In_2046,In_1932);
nand U4065 (N_4065,In_980,In_1081);
or U4066 (N_4066,In_2167,In_2317);
or U4067 (N_4067,In_822,In_2145);
or U4068 (N_4068,In_133,In_2049);
nand U4069 (N_4069,In_1387,In_1151);
or U4070 (N_4070,In_82,In_2299);
nor U4071 (N_4071,In_2448,In_949);
nand U4072 (N_4072,In_1524,In_539);
or U4073 (N_4073,In_285,In_1461);
and U4074 (N_4074,In_1272,In_1655);
xor U4075 (N_4075,In_887,In_2156);
nor U4076 (N_4076,In_445,In_2452);
and U4077 (N_4077,In_1228,In_987);
xnor U4078 (N_4078,In_2044,In_1678);
nand U4079 (N_4079,In_57,In_2184);
xnor U4080 (N_4080,In_759,In_301);
or U4081 (N_4081,In_1161,In_170);
xnor U4082 (N_4082,In_1114,In_608);
or U4083 (N_4083,In_2288,In_1109);
nand U4084 (N_4084,In_1050,In_143);
xnor U4085 (N_4085,In_2430,In_720);
nand U4086 (N_4086,In_1751,In_1950);
nand U4087 (N_4087,In_334,In_2334);
or U4088 (N_4088,In_1043,In_2339);
nor U4089 (N_4089,In_938,In_1320);
nand U4090 (N_4090,In_434,In_1172);
and U4091 (N_4091,In_1470,In_364);
or U4092 (N_4092,In_533,In_823);
and U4093 (N_4093,In_705,In_1449);
nor U4094 (N_4094,In_172,In_2341);
or U4095 (N_4095,In_425,In_2237);
or U4096 (N_4096,In_136,In_468);
and U4097 (N_4097,In_2363,In_74);
xor U4098 (N_4098,In_61,In_138);
or U4099 (N_4099,In_336,In_904);
nand U4100 (N_4100,In_1099,In_1996);
nor U4101 (N_4101,In_334,In_1067);
xnor U4102 (N_4102,In_1244,In_298);
or U4103 (N_4103,In_2120,In_1143);
xor U4104 (N_4104,In_2277,In_811);
or U4105 (N_4105,In_654,In_358);
or U4106 (N_4106,In_810,In_972);
xor U4107 (N_4107,In_62,In_342);
xnor U4108 (N_4108,In_444,In_1515);
nand U4109 (N_4109,In_683,In_1661);
and U4110 (N_4110,In_1354,In_1472);
xnor U4111 (N_4111,In_1541,In_599);
nand U4112 (N_4112,In_1773,In_1875);
xnor U4113 (N_4113,In_765,In_2347);
or U4114 (N_4114,In_800,In_632);
and U4115 (N_4115,In_1493,In_332);
or U4116 (N_4116,In_405,In_358);
or U4117 (N_4117,In_2200,In_1933);
and U4118 (N_4118,In_149,In_421);
and U4119 (N_4119,In_1511,In_2136);
xor U4120 (N_4120,In_1717,In_1062);
nor U4121 (N_4121,In_125,In_2098);
nor U4122 (N_4122,In_844,In_2289);
nand U4123 (N_4123,In_2000,In_2497);
and U4124 (N_4124,In_2473,In_1977);
and U4125 (N_4125,In_1114,In_323);
nor U4126 (N_4126,In_1577,In_1325);
xnor U4127 (N_4127,In_1931,In_1245);
nor U4128 (N_4128,In_384,In_1331);
nor U4129 (N_4129,In_1116,In_827);
or U4130 (N_4130,In_842,In_280);
nand U4131 (N_4131,In_2291,In_1218);
xor U4132 (N_4132,In_1436,In_1860);
nand U4133 (N_4133,In_1856,In_1230);
or U4134 (N_4134,In_63,In_1707);
nand U4135 (N_4135,In_1314,In_353);
and U4136 (N_4136,In_166,In_362);
and U4137 (N_4137,In_420,In_2285);
nand U4138 (N_4138,In_2247,In_1073);
xnor U4139 (N_4139,In_1643,In_600);
or U4140 (N_4140,In_624,In_2105);
xnor U4141 (N_4141,In_1933,In_2151);
xnor U4142 (N_4142,In_1911,In_1463);
xnor U4143 (N_4143,In_409,In_598);
nor U4144 (N_4144,In_1347,In_411);
or U4145 (N_4145,In_628,In_420);
or U4146 (N_4146,In_848,In_2297);
or U4147 (N_4147,In_1232,In_1767);
nor U4148 (N_4148,In_1770,In_1616);
nor U4149 (N_4149,In_1430,In_2246);
and U4150 (N_4150,In_3,In_2481);
and U4151 (N_4151,In_1500,In_59);
or U4152 (N_4152,In_1261,In_378);
and U4153 (N_4153,In_1476,In_1281);
xor U4154 (N_4154,In_1338,In_2364);
nor U4155 (N_4155,In_1630,In_1635);
and U4156 (N_4156,In_779,In_1187);
or U4157 (N_4157,In_2297,In_2349);
xnor U4158 (N_4158,In_262,In_2170);
and U4159 (N_4159,In_610,In_2177);
nand U4160 (N_4160,In_1830,In_2452);
xor U4161 (N_4161,In_626,In_1208);
nand U4162 (N_4162,In_1325,In_574);
nor U4163 (N_4163,In_822,In_2122);
xor U4164 (N_4164,In_2467,In_387);
and U4165 (N_4165,In_896,In_1648);
or U4166 (N_4166,In_1408,In_2184);
nor U4167 (N_4167,In_499,In_2375);
and U4168 (N_4168,In_1881,In_1033);
and U4169 (N_4169,In_1775,In_1025);
nand U4170 (N_4170,In_972,In_326);
or U4171 (N_4171,In_464,In_1604);
nor U4172 (N_4172,In_369,In_825);
and U4173 (N_4173,In_2416,In_2243);
and U4174 (N_4174,In_642,In_1704);
or U4175 (N_4175,In_1017,In_280);
xnor U4176 (N_4176,In_61,In_1381);
nand U4177 (N_4177,In_682,In_862);
and U4178 (N_4178,In_1323,In_373);
nand U4179 (N_4179,In_832,In_325);
nand U4180 (N_4180,In_1605,In_588);
xor U4181 (N_4181,In_2092,In_355);
nand U4182 (N_4182,In_1553,In_1442);
xor U4183 (N_4183,In_1136,In_1247);
xnor U4184 (N_4184,In_1465,In_964);
or U4185 (N_4185,In_1381,In_1152);
nand U4186 (N_4186,In_1919,In_407);
and U4187 (N_4187,In_789,In_1962);
and U4188 (N_4188,In_1792,In_16);
or U4189 (N_4189,In_1245,In_108);
nor U4190 (N_4190,In_324,In_2335);
and U4191 (N_4191,In_1428,In_459);
nand U4192 (N_4192,In_848,In_150);
nor U4193 (N_4193,In_642,In_848);
nor U4194 (N_4194,In_357,In_1931);
nor U4195 (N_4195,In_942,In_1624);
nand U4196 (N_4196,In_1535,In_794);
or U4197 (N_4197,In_1122,In_2010);
nand U4198 (N_4198,In_1170,In_1647);
and U4199 (N_4199,In_2149,In_1471);
xnor U4200 (N_4200,In_356,In_503);
nand U4201 (N_4201,In_2281,In_571);
nand U4202 (N_4202,In_1447,In_361);
nor U4203 (N_4203,In_1509,In_1553);
and U4204 (N_4204,In_923,In_715);
and U4205 (N_4205,In_357,In_644);
and U4206 (N_4206,In_886,In_1589);
nor U4207 (N_4207,In_1388,In_1821);
and U4208 (N_4208,In_339,In_2167);
nand U4209 (N_4209,In_1706,In_1878);
and U4210 (N_4210,In_2443,In_143);
nor U4211 (N_4211,In_1350,In_469);
or U4212 (N_4212,In_490,In_1539);
and U4213 (N_4213,In_762,In_604);
xnor U4214 (N_4214,In_666,In_741);
nor U4215 (N_4215,In_2130,In_651);
nor U4216 (N_4216,In_1698,In_53);
xor U4217 (N_4217,In_1300,In_1966);
or U4218 (N_4218,In_445,In_1393);
xnor U4219 (N_4219,In_409,In_836);
xnor U4220 (N_4220,In_302,In_1973);
and U4221 (N_4221,In_444,In_1712);
and U4222 (N_4222,In_2330,In_307);
nor U4223 (N_4223,In_2146,In_1672);
nand U4224 (N_4224,In_1090,In_1808);
and U4225 (N_4225,In_1912,In_1400);
xor U4226 (N_4226,In_436,In_899);
nand U4227 (N_4227,In_1117,In_584);
and U4228 (N_4228,In_1197,In_449);
and U4229 (N_4229,In_2189,In_2231);
or U4230 (N_4230,In_517,In_2067);
xor U4231 (N_4231,In_1472,In_2025);
xnor U4232 (N_4232,In_1866,In_1913);
xnor U4233 (N_4233,In_1490,In_1950);
and U4234 (N_4234,In_1232,In_1625);
and U4235 (N_4235,In_101,In_985);
xnor U4236 (N_4236,In_465,In_1914);
nand U4237 (N_4237,In_2245,In_350);
nor U4238 (N_4238,In_1765,In_1045);
nand U4239 (N_4239,In_1200,In_2472);
nor U4240 (N_4240,In_1091,In_1230);
or U4241 (N_4241,In_1972,In_2295);
nand U4242 (N_4242,In_1786,In_1776);
xor U4243 (N_4243,In_449,In_865);
nand U4244 (N_4244,In_2088,In_2228);
xor U4245 (N_4245,In_1254,In_1782);
or U4246 (N_4246,In_1476,In_2115);
or U4247 (N_4247,In_2488,In_1739);
xnor U4248 (N_4248,In_1408,In_207);
or U4249 (N_4249,In_1948,In_247);
nand U4250 (N_4250,In_878,In_587);
nand U4251 (N_4251,In_1226,In_2279);
nand U4252 (N_4252,In_1444,In_2284);
nor U4253 (N_4253,In_789,In_750);
nand U4254 (N_4254,In_2216,In_1450);
or U4255 (N_4255,In_369,In_2061);
or U4256 (N_4256,In_3,In_582);
or U4257 (N_4257,In_2287,In_2051);
and U4258 (N_4258,In_1224,In_1403);
or U4259 (N_4259,In_185,In_596);
nor U4260 (N_4260,In_2212,In_1342);
xnor U4261 (N_4261,In_1473,In_2173);
nor U4262 (N_4262,In_413,In_316);
or U4263 (N_4263,In_244,In_1606);
and U4264 (N_4264,In_2048,In_1089);
and U4265 (N_4265,In_2314,In_788);
or U4266 (N_4266,In_646,In_1036);
nor U4267 (N_4267,In_976,In_1423);
or U4268 (N_4268,In_1681,In_1565);
xor U4269 (N_4269,In_1796,In_816);
nand U4270 (N_4270,In_723,In_57);
nor U4271 (N_4271,In_631,In_109);
nand U4272 (N_4272,In_1027,In_676);
nand U4273 (N_4273,In_2180,In_2108);
nor U4274 (N_4274,In_1885,In_663);
nand U4275 (N_4275,In_2069,In_1633);
nand U4276 (N_4276,In_1610,In_1855);
and U4277 (N_4277,In_2004,In_54);
xnor U4278 (N_4278,In_849,In_380);
nor U4279 (N_4279,In_122,In_565);
nor U4280 (N_4280,In_1047,In_503);
xor U4281 (N_4281,In_1482,In_1136);
and U4282 (N_4282,In_72,In_670);
nand U4283 (N_4283,In_1409,In_1755);
nand U4284 (N_4284,In_437,In_1910);
xnor U4285 (N_4285,In_90,In_371);
xnor U4286 (N_4286,In_2148,In_1061);
nor U4287 (N_4287,In_1245,In_301);
nand U4288 (N_4288,In_2357,In_299);
nor U4289 (N_4289,In_952,In_915);
nand U4290 (N_4290,In_244,In_17);
xor U4291 (N_4291,In_584,In_1031);
nor U4292 (N_4292,In_1512,In_2068);
or U4293 (N_4293,In_559,In_656);
or U4294 (N_4294,In_1376,In_2068);
nor U4295 (N_4295,In_1086,In_2023);
nand U4296 (N_4296,In_2144,In_1671);
or U4297 (N_4297,In_392,In_571);
nand U4298 (N_4298,In_2426,In_1082);
or U4299 (N_4299,In_2402,In_1869);
and U4300 (N_4300,In_537,In_1651);
xnor U4301 (N_4301,In_355,In_1723);
nand U4302 (N_4302,In_1247,In_1786);
or U4303 (N_4303,In_345,In_683);
nor U4304 (N_4304,In_1632,In_822);
or U4305 (N_4305,In_736,In_2428);
or U4306 (N_4306,In_489,In_1073);
xor U4307 (N_4307,In_2069,In_239);
or U4308 (N_4308,In_573,In_1494);
or U4309 (N_4309,In_1356,In_515);
nor U4310 (N_4310,In_821,In_1531);
xnor U4311 (N_4311,In_872,In_1512);
nor U4312 (N_4312,In_1290,In_1156);
xnor U4313 (N_4313,In_350,In_615);
xor U4314 (N_4314,In_1222,In_843);
and U4315 (N_4315,In_2047,In_852);
or U4316 (N_4316,In_2210,In_1757);
nand U4317 (N_4317,In_1842,In_1729);
xnor U4318 (N_4318,In_1828,In_861);
xor U4319 (N_4319,In_307,In_1775);
and U4320 (N_4320,In_650,In_864);
and U4321 (N_4321,In_1934,In_2355);
or U4322 (N_4322,In_2161,In_1237);
nor U4323 (N_4323,In_780,In_1435);
xnor U4324 (N_4324,In_2264,In_1800);
or U4325 (N_4325,In_452,In_1704);
xnor U4326 (N_4326,In_506,In_1735);
and U4327 (N_4327,In_2499,In_1066);
xor U4328 (N_4328,In_770,In_890);
and U4329 (N_4329,In_1636,In_303);
and U4330 (N_4330,In_666,In_910);
or U4331 (N_4331,In_2170,In_121);
nand U4332 (N_4332,In_2427,In_641);
and U4333 (N_4333,In_484,In_2145);
xor U4334 (N_4334,In_1808,In_543);
nor U4335 (N_4335,In_897,In_261);
xnor U4336 (N_4336,In_1913,In_642);
or U4337 (N_4337,In_1994,In_2025);
nor U4338 (N_4338,In_1684,In_1003);
nor U4339 (N_4339,In_585,In_1923);
nor U4340 (N_4340,In_274,In_1901);
or U4341 (N_4341,In_258,In_1604);
xor U4342 (N_4342,In_1390,In_1286);
nand U4343 (N_4343,In_1545,In_903);
xnor U4344 (N_4344,In_1209,In_498);
and U4345 (N_4345,In_1791,In_297);
or U4346 (N_4346,In_1006,In_2422);
xor U4347 (N_4347,In_210,In_1841);
nor U4348 (N_4348,In_184,In_452);
nor U4349 (N_4349,In_2204,In_588);
nand U4350 (N_4350,In_838,In_1832);
nand U4351 (N_4351,In_350,In_1386);
nor U4352 (N_4352,In_1571,In_438);
or U4353 (N_4353,In_1340,In_2422);
and U4354 (N_4354,In_2304,In_12);
xnor U4355 (N_4355,In_1647,In_1413);
xor U4356 (N_4356,In_1017,In_1471);
or U4357 (N_4357,In_1800,In_2184);
and U4358 (N_4358,In_843,In_2404);
or U4359 (N_4359,In_1086,In_1259);
nand U4360 (N_4360,In_500,In_2224);
and U4361 (N_4361,In_1364,In_1490);
nor U4362 (N_4362,In_1203,In_603);
and U4363 (N_4363,In_1126,In_1492);
nand U4364 (N_4364,In_730,In_1132);
and U4365 (N_4365,In_260,In_1654);
nand U4366 (N_4366,In_1664,In_610);
or U4367 (N_4367,In_360,In_2251);
nand U4368 (N_4368,In_725,In_1163);
or U4369 (N_4369,In_1964,In_2434);
nor U4370 (N_4370,In_328,In_2152);
xor U4371 (N_4371,In_1452,In_1999);
xor U4372 (N_4372,In_2165,In_1968);
xnor U4373 (N_4373,In_1041,In_1653);
nand U4374 (N_4374,In_363,In_694);
nand U4375 (N_4375,In_1030,In_1043);
and U4376 (N_4376,In_2246,In_526);
and U4377 (N_4377,In_635,In_1197);
or U4378 (N_4378,In_1577,In_1428);
nand U4379 (N_4379,In_21,In_710);
or U4380 (N_4380,In_544,In_1883);
nor U4381 (N_4381,In_695,In_519);
and U4382 (N_4382,In_58,In_1688);
xnor U4383 (N_4383,In_2258,In_587);
nor U4384 (N_4384,In_1248,In_1596);
nor U4385 (N_4385,In_284,In_519);
xnor U4386 (N_4386,In_1046,In_1457);
xnor U4387 (N_4387,In_240,In_1896);
or U4388 (N_4388,In_1159,In_619);
or U4389 (N_4389,In_230,In_1013);
xor U4390 (N_4390,In_581,In_1724);
nor U4391 (N_4391,In_2082,In_864);
xor U4392 (N_4392,In_989,In_2386);
nand U4393 (N_4393,In_223,In_1448);
nand U4394 (N_4394,In_207,In_820);
or U4395 (N_4395,In_2380,In_1558);
nor U4396 (N_4396,In_1513,In_2255);
and U4397 (N_4397,In_708,In_959);
nand U4398 (N_4398,In_409,In_1467);
and U4399 (N_4399,In_985,In_1939);
or U4400 (N_4400,In_2233,In_723);
and U4401 (N_4401,In_1111,In_1915);
xor U4402 (N_4402,In_472,In_1155);
or U4403 (N_4403,In_1303,In_720);
and U4404 (N_4404,In_1156,In_255);
nand U4405 (N_4405,In_1914,In_182);
nand U4406 (N_4406,In_1221,In_2053);
nand U4407 (N_4407,In_1664,In_50);
nor U4408 (N_4408,In_1050,In_6);
xnor U4409 (N_4409,In_675,In_263);
or U4410 (N_4410,In_1305,In_1682);
nor U4411 (N_4411,In_2406,In_73);
nand U4412 (N_4412,In_1580,In_803);
or U4413 (N_4413,In_1783,In_1882);
or U4414 (N_4414,In_57,In_1305);
or U4415 (N_4415,In_2361,In_646);
or U4416 (N_4416,In_843,In_849);
or U4417 (N_4417,In_1248,In_2415);
and U4418 (N_4418,In_1871,In_469);
nor U4419 (N_4419,In_2057,In_1950);
or U4420 (N_4420,In_2256,In_910);
nand U4421 (N_4421,In_1349,In_2497);
and U4422 (N_4422,In_1523,In_1557);
nor U4423 (N_4423,In_1807,In_2006);
xnor U4424 (N_4424,In_1174,In_246);
and U4425 (N_4425,In_2413,In_2385);
xnor U4426 (N_4426,In_1464,In_2103);
nor U4427 (N_4427,In_87,In_2452);
nand U4428 (N_4428,In_1699,In_2156);
nand U4429 (N_4429,In_988,In_252);
nor U4430 (N_4430,In_189,In_2437);
nor U4431 (N_4431,In_551,In_329);
nor U4432 (N_4432,In_1150,In_1982);
and U4433 (N_4433,In_2189,In_1829);
xor U4434 (N_4434,In_198,In_137);
nor U4435 (N_4435,In_1221,In_2003);
nand U4436 (N_4436,In_1528,In_24);
or U4437 (N_4437,In_2497,In_2261);
and U4438 (N_4438,In_1744,In_1567);
and U4439 (N_4439,In_632,In_667);
xor U4440 (N_4440,In_2256,In_1662);
or U4441 (N_4441,In_870,In_542);
nand U4442 (N_4442,In_100,In_2227);
xnor U4443 (N_4443,In_1353,In_1003);
nand U4444 (N_4444,In_870,In_1558);
nand U4445 (N_4445,In_2102,In_1997);
nand U4446 (N_4446,In_82,In_898);
nor U4447 (N_4447,In_1657,In_1168);
xor U4448 (N_4448,In_2204,In_410);
xor U4449 (N_4449,In_1846,In_1648);
nor U4450 (N_4450,In_498,In_2444);
or U4451 (N_4451,In_863,In_339);
and U4452 (N_4452,In_2340,In_1347);
nor U4453 (N_4453,In_1369,In_2004);
and U4454 (N_4454,In_618,In_969);
nand U4455 (N_4455,In_1340,In_702);
nand U4456 (N_4456,In_1326,In_1078);
nor U4457 (N_4457,In_1843,In_494);
and U4458 (N_4458,In_39,In_1712);
nor U4459 (N_4459,In_186,In_882);
and U4460 (N_4460,In_1372,In_1317);
xor U4461 (N_4461,In_1291,In_1627);
nor U4462 (N_4462,In_2324,In_1800);
nand U4463 (N_4463,In_1319,In_52);
nor U4464 (N_4464,In_724,In_24);
or U4465 (N_4465,In_517,In_320);
or U4466 (N_4466,In_345,In_395);
xnor U4467 (N_4467,In_24,In_549);
nand U4468 (N_4468,In_2149,In_379);
and U4469 (N_4469,In_1856,In_1366);
xor U4470 (N_4470,In_320,In_1920);
xor U4471 (N_4471,In_1611,In_2357);
or U4472 (N_4472,In_1527,In_2010);
xnor U4473 (N_4473,In_148,In_503);
nand U4474 (N_4474,In_1433,In_2191);
nand U4475 (N_4475,In_938,In_1149);
or U4476 (N_4476,In_1745,In_323);
nor U4477 (N_4477,In_1979,In_1256);
xor U4478 (N_4478,In_644,In_2180);
nor U4479 (N_4479,In_2305,In_2459);
xor U4480 (N_4480,In_562,In_1974);
xnor U4481 (N_4481,In_1516,In_281);
or U4482 (N_4482,In_394,In_1665);
or U4483 (N_4483,In_765,In_2039);
or U4484 (N_4484,In_358,In_1918);
xor U4485 (N_4485,In_944,In_600);
xnor U4486 (N_4486,In_538,In_957);
or U4487 (N_4487,In_1850,In_1101);
nor U4488 (N_4488,In_2189,In_905);
nor U4489 (N_4489,In_2231,In_113);
xor U4490 (N_4490,In_2312,In_2263);
nor U4491 (N_4491,In_2006,In_1209);
and U4492 (N_4492,In_794,In_595);
xnor U4493 (N_4493,In_352,In_892);
nand U4494 (N_4494,In_2326,In_1354);
or U4495 (N_4495,In_1731,In_1968);
nand U4496 (N_4496,In_1214,In_454);
nand U4497 (N_4497,In_328,In_1484);
and U4498 (N_4498,In_1168,In_2169);
or U4499 (N_4499,In_907,In_1234);
nand U4500 (N_4500,In_1355,In_171);
nand U4501 (N_4501,In_786,In_854);
xor U4502 (N_4502,In_1657,In_1561);
and U4503 (N_4503,In_2233,In_1171);
xnor U4504 (N_4504,In_133,In_2300);
and U4505 (N_4505,In_1768,In_1586);
or U4506 (N_4506,In_1300,In_784);
xor U4507 (N_4507,In_1613,In_1397);
or U4508 (N_4508,In_1873,In_894);
and U4509 (N_4509,In_693,In_234);
or U4510 (N_4510,In_2015,In_23);
and U4511 (N_4511,In_874,In_1380);
nand U4512 (N_4512,In_1618,In_824);
and U4513 (N_4513,In_981,In_488);
nor U4514 (N_4514,In_1874,In_130);
xor U4515 (N_4515,In_1353,In_2206);
or U4516 (N_4516,In_93,In_2486);
or U4517 (N_4517,In_931,In_945);
nor U4518 (N_4518,In_35,In_1826);
nor U4519 (N_4519,In_2168,In_1897);
nand U4520 (N_4520,In_343,In_2192);
or U4521 (N_4521,In_1418,In_508);
nor U4522 (N_4522,In_2297,In_1474);
and U4523 (N_4523,In_822,In_74);
xnor U4524 (N_4524,In_1271,In_1657);
nor U4525 (N_4525,In_1484,In_605);
xnor U4526 (N_4526,In_2177,In_926);
nor U4527 (N_4527,In_5,In_1692);
nand U4528 (N_4528,In_39,In_2485);
or U4529 (N_4529,In_701,In_730);
or U4530 (N_4530,In_2077,In_1811);
or U4531 (N_4531,In_2155,In_2116);
or U4532 (N_4532,In_1042,In_61);
or U4533 (N_4533,In_189,In_2074);
and U4534 (N_4534,In_58,In_101);
and U4535 (N_4535,In_1823,In_1464);
or U4536 (N_4536,In_1739,In_1816);
nand U4537 (N_4537,In_1548,In_2424);
nand U4538 (N_4538,In_493,In_601);
and U4539 (N_4539,In_1993,In_1555);
nor U4540 (N_4540,In_688,In_831);
xor U4541 (N_4541,In_2441,In_966);
or U4542 (N_4542,In_2063,In_1522);
nand U4543 (N_4543,In_64,In_905);
and U4544 (N_4544,In_1108,In_2100);
xor U4545 (N_4545,In_1358,In_1107);
and U4546 (N_4546,In_1867,In_1717);
xnor U4547 (N_4547,In_2062,In_806);
nor U4548 (N_4548,In_1909,In_159);
and U4549 (N_4549,In_2325,In_1772);
and U4550 (N_4550,In_1424,In_2278);
or U4551 (N_4551,In_1676,In_659);
and U4552 (N_4552,In_725,In_929);
nand U4553 (N_4553,In_854,In_1184);
or U4554 (N_4554,In_1060,In_1687);
nor U4555 (N_4555,In_2225,In_2135);
or U4556 (N_4556,In_857,In_1949);
xor U4557 (N_4557,In_2497,In_2375);
nand U4558 (N_4558,In_1790,In_2107);
nand U4559 (N_4559,In_489,In_1077);
nand U4560 (N_4560,In_333,In_1976);
nand U4561 (N_4561,In_114,In_1110);
nor U4562 (N_4562,In_388,In_1699);
nor U4563 (N_4563,In_1320,In_2469);
nor U4564 (N_4564,In_1063,In_1579);
xor U4565 (N_4565,In_1221,In_898);
nand U4566 (N_4566,In_1194,In_249);
or U4567 (N_4567,In_1202,In_548);
and U4568 (N_4568,In_2445,In_2107);
or U4569 (N_4569,In_1253,In_2287);
or U4570 (N_4570,In_1277,In_2225);
xor U4571 (N_4571,In_1374,In_3);
xor U4572 (N_4572,In_1302,In_1975);
nand U4573 (N_4573,In_619,In_178);
xnor U4574 (N_4574,In_959,In_1804);
and U4575 (N_4575,In_1713,In_1280);
nand U4576 (N_4576,In_691,In_2000);
or U4577 (N_4577,In_1123,In_1030);
or U4578 (N_4578,In_2353,In_1458);
and U4579 (N_4579,In_1019,In_455);
nand U4580 (N_4580,In_1312,In_922);
nand U4581 (N_4581,In_703,In_1536);
nor U4582 (N_4582,In_2208,In_211);
nor U4583 (N_4583,In_713,In_1433);
and U4584 (N_4584,In_124,In_1806);
or U4585 (N_4585,In_1641,In_1789);
and U4586 (N_4586,In_1381,In_1655);
and U4587 (N_4587,In_157,In_681);
and U4588 (N_4588,In_107,In_1940);
and U4589 (N_4589,In_1431,In_2133);
xnor U4590 (N_4590,In_976,In_971);
or U4591 (N_4591,In_1487,In_1057);
xor U4592 (N_4592,In_1263,In_1760);
nor U4593 (N_4593,In_2495,In_1444);
nand U4594 (N_4594,In_2096,In_1967);
nor U4595 (N_4595,In_1287,In_429);
nand U4596 (N_4596,In_939,In_62);
xnor U4597 (N_4597,In_1345,In_312);
or U4598 (N_4598,In_230,In_1129);
nand U4599 (N_4599,In_455,In_1694);
nor U4600 (N_4600,In_790,In_311);
nor U4601 (N_4601,In_1594,In_2106);
nor U4602 (N_4602,In_427,In_568);
and U4603 (N_4603,In_896,In_2211);
and U4604 (N_4604,In_757,In_138);
nand U4605 (N_4605,In_943,In_225);
xor U4606 (N_4606,In_2248,In_767);
or U4607 (N_4607,In_2246,In_2339);
and U4608 (N_4608,In_1712,In_352);
nand U4609 (N_4609,In_1398,In_1933);
or U4610 (N_4610,In_1713,In_2335);
or U4611 (N_4611,In_1028,In_2249);
and U4612 (N_4612,In_1417,In_1500);
and U4613 (N_4613,In_1693,In_1867);
nand U4614 (N_4614,In_1,In_2266);
nor U4615 (N_4615,In_673,In_743);
and U4616 (N_4616,In_2086,In_377);
xnor U4617 (N_4617,In_2356,In_194);
and U4618 (N_4618,In_962,In_1932);
and U4619 (N_4619,In_1489,In_1);
or U4620 (N_4620,In_430,In_1683);
or U4621 (N_4621,In_494,In_2036);
or U4622 (N_4622,In_756,In_1496);
nor U4623 (N_4623,In_2443,In_361);
nand U4624 (N_4624,In_1367,In_2469);
or U4625 (N_4625,In_1540,In_2369);
and U4626 (N_4626,In_2143,In_741);
and U4627 (N_4627,In_618,In_1619);
nor U4628 (N_4628,In_1687,In_917);
or U4629 (N_4629,In_1029,In_801);
nand U4630 (N_4630,In_1829,In_1758);
xor U4631 (N_4631,In_2107,In_151);
nand U4632 (N_4632,In_997,In_424);
xor U4633 (N_4633,In_2431,In_943);
nor U4634 (N_4634,In_1900,In_155);
nor U4635 (N_4635,In_2190,In_1640);
xor U4636 (N_4636,In_1318,In_1904);
nor U4637 (N_4637,In_1089,In_761);
nand U4638 (N_4638,In_1078,In_2496);
nor U4639 (N_4639,In_1634,In_525);
or U4640 (N_4640,In_60,In_1755);
nor U4641 (N_4641,In_1493,In_277);
or U4642 (N_4642,In_2327,In_138);
nand U4643 (N_4643,In_1881,In_216);
or U4644 (N_4644,In_1997,In_2430);
xnor U4645 (N_4645,In_1643,In_16);
xnor U4646 (N_4646,In_2356,In_638);
and U4647 (N_4647,In_1341,In_2371);
or U4648 (N_4648,In_2176,In_1955);
or U4649 (N_4649,In_1900,In_738);
or U4650 (N_4650,In_783,In_1005);
or U4651 (N_4651,In_682,In_1727);
xnor U4652 (N_4652,In_1063,In_499);
nand U4653 (N_4653,In_1709,In_2166);
nand U4654 (N_4654,In_346,In_205);
and U4655 (N_4655,In_467,In_415);
or U4656 (N_4656,In_2239,In_266);
nor U4657 (N_4657,In_1954,In_45);
or U4658 (N_4658,In_321,In_2370);
and U4659 (N_4659,In_27,In_2001);
and U4660 (N_4660,In_280,In_1352);
and U4661 (N_4661,In_749,In_301);
and U4662 (N_4662,In_1399,In_548);
xor U4663 (N_4663,In_1854,In_100);
and U4664 (N_4664,In_875,In_789);
nor U4665 (N_4665,In_2251,In_42);
and U4666 (N_4666,In_1202,In_637);
or U4667 (N_4667,In_1183,In_102);
nand U4668 (N_4668,In_289,In_890);
nand U4669 (N_4669,In_1906,In_594);
nand U4670 (N_4670,In_559,In_1953);
nor U4671 (N_4671,In_2216,In_2120);
nor U4672 (N_4672,In_1338,In_1218);
or U4673 (N_4673,In_2079,In_63);
or U4674 (N_4674,In_1051,In_1044);
and U4675 (N_4675,In_1642,In_1797);
or U4676 (N_4676,In_487,In_1935);
nor U4677 (N_4677,In_1522,In_2364);
nor U4678 (N_4678,In_266,In_760);
and U4679 (N_4679,In_1508,In_482);
and U4680 (N_4680,In_444,In_2268);
and U4681 (N_4681,In_2437,In_404);
nand U4682 (N_4682,In_2080,In_672);
xor U4683 (N_4683,In_1235,In_778);
nand U4684 (N_4684,In_264,In_1093);
nor U4685 (N_4685,In_636,In_2139);
nand U4686 (N_4686,In_1698,In_840);
and U4687 (N_4687,In_219,In_1736);
and U4688 (N_4688,In_2004,In_2326);
xor U4689 (N_4689,In_168,In_857);
or U4690 (N_4690,In_830,In_2398);
xor U4691 (N_4691,In_1449,In_2466);
nand U4692 (N_4692,In_1490,In_1602);
and U4693 (N_4693,In_2230,In_2142);
xor U4694 (N_4694,In_2399,In_1093);
xor U4695 (N_4695,In_625,In_828);
or U4696 (N_4696,In_1482,In_1981);
nand U4697 (N_4697,In_247,In_269);
nor U4698 (N_4698,In_1874,In_924);
nor U4699 (N_4699,In_1072,In_1309);
nor U4700 (N_4700,In_303,In_1499);
nor U4701 (N_4701,In_1241,In_1250);
nand U4702 (N_4702,In_1771,In_974);
and U4703 (N_4703,In_1229,In_7);
and U4704 (N_4704,In_1125,In_2397);
nor U4705 (N_4705,In_1891,In_697);
xor U4706 (N_4706,In_1723,In_250);
xnor U4707 (N_4707,In_1494,In_692);
nand U4708 (N_4708,In_2223,In_2314);
or U4709 (N_4709,In_1341,In_1807);
nand U4710 (N_4710,In_1339,In_1733);
xor U4711 (N_4711,In_189,In_486);
nand U4712 (N_4712,In_139,In_2187);
xnor U4713 (N_4713,In_564,In_1682);
xor U4714 (N_4714,In_2101,In_1132);
and U4715 (N_4715,In_2326,In_1248);
and U4716 (N_4716,In_2454,In_1896);
or U4717 (N_4717,In_1481,In_2411);
xnor U4718 (N_4718,In_960,In_361);
nor U4719 (N_4719,In_1976,In_516);
or U4720 (N_4720,In_1813,In_2488);
nor U4721 (N_4721,In_1295,In_2270);
and U4722 (N_4722,In_1482,In_780);
or U4723 (N_4723,In_2282,In_1330);
nor U4724 (N_4724,In_1023,In_2359);
or U4725 (N_4725,In_1039,In_1528);
or U4726 (N_4726,In_1505,In_1225);
nand U4727 (N_4727,In_2327,In_328);
or U4728 (N_4728,In_1072,In_326);
xnor U4729 (N_4729,In_1347,In_1558);
nor U4730 (N_4730,In_1952,In_832);
xnor U4731 (N_4731,In_2133,In_394);
or U4732 (N_4732,In_569,In_2401);
nand U4733 (N_4733,In_1634,In_693);
xor U4734 (N_4734,In_1931,In_1521);
nor U4735 (N_4735,In_2466,In_1534);
xor U4736 (N_4736,In_767,In_883);
or U4737 (N_4737,In_1215,In_1811);
or U4738 (N_4738,In_1411,In_1936);
xnor U4739 (N_4739,In_2204,In_1946);
nor U4740 (N_4740,In_2349,In_1086);
nand U4741 (N_4741,In_2241,In_933);
and U4742 (N_4742,In_1352,In_1856);
and U4743 (N_4743,In_2448,In_2240);
and U4744 (N_4744,In_643,In_1339);
xnor U4745 (N_4745,In_883,In_572);
or U4746 (N_4746,In_305,In_2296);
or U4747 (N_4747,In_18,In_2177);
and U4748 (N_4748,In_1373,In_1169);
nand U4749 (N_4749,In_1696,In_445);
nor U4750 (N_4750,In_350,In_1542);
xnor U4751 (N_4751,In_1928,In_65);
or U4752 (N_4752,In_2283,In_1621);
and U4753 (N_4753,In_1555,In_2318);
nand U4754 (N_4754,In_1996,In_542);
nor U4755 (N_4755,In_2398,In_591);
nand U4756 (N_4756,In_1167,In_1344);
or U4757 (N_4757,In_2424,In_2038);
nor U4758 (N_4758,In_2217,In_201);
nor U4759 (N_4759,In_1215,In_610);
or U4760 (N_4760,In_701,In_1493);
xnor U4761 (N_4761,In_1095,In_2030);
nand U4762 (N_4762,In_2099,In_437);
nor U4763 (N_4763,In_683,In_2006);
xnor U4764 (N_4764,In_2420,In_859);
and U4765 (N_4765,In_86,In_435);
nand U4766 (N_4766,In_2326,In_319);
nand U4767 (N_4767,In_486,In_1761);
nor U4768 (N_4768,In_724,In_1914);
and U4769 (N_4769,In_2075,In_679);
and U4770 (N_4770,In_1639,In_750);
nand U4771 (N_4771,In_2491,In_500);
or U4772 (N_4772,In_737,In_2430);
xnor U4773 (N_4773,In_330,In_2098);
or U4774 (N_4774,In_1992,In_824);
xnor U4775 (N_4775,In_326,In_435);
and U4776 (N_4776,In_133,In_210);
nor U4777 (N_4777,In_2494,In_536);
and U4778 (N_4778,In_1016,In_1472);
and U4779 (N_4779,In_570,In_2137);
xor U4780 (N_4780,In_1504,In_1723);
and U4781 (N_4781,In_1444,In_1961);
xor U4782 (N_4782,In_1112,In_757);
or U4783 (N_4783,In_415,In_2262);
nor U4784 (N_4784,In_1626,In_432);
nand U4785 (N_4785,In_1491,In_59);
and U4786 (N_4786,In_2184,In_1926);
and U4787 (N_4787,In_1405,In_814);
xor U4788 (N_4788,In_1298,In_1574);
nor U4789 (N_4789,In_628,In_1443);
nand U4790 (N_4790,In_43,In_1815);
nand U4791 (N_4791,In_1527,In_1207);
and U4792 (N_4792,In_125,In_99);
xor U4793 (N_4793,In_2059,In_1051);
xor U4794 (N_4794,In_1788,In_1282);
nor U4795 (N_4795,In_190,In_2476);
and U4796 (N_4796,In_552,In_1693);
nand U4797 (N_4797,In_244,In_564);
nor U4798 (N_4798,In_731,In_868);
nor U4799 (N_4799,In_1280,In_341);
nor U4800 (N_4800,In_1668,In_912);
nand U4801 (N_4801,In_1183,In_308);
nor U4802 (N_4802,In_978,In_1817);
nand U4803 (N_4803,In_1741,In_2429);
xnor U4804 (N_4804,In_288,In_858);
or U4805 (N_4805,In_2362,In_1340);
nand U4806 (N_4806,In_1218,In_1730);
xor U4807 (N_4807,In_1606,In_2431);
xnor U4808 (N_4808,In_235,In_1717);
and U4809 (N_4809,In_510,In_2266);
nor U4810 (N_4810,In_628,In_524);
nand U4811 (N_4811,In_610,In_654);
nor U4812 (N_4812,In_1204,In_7);
nand U4813 (N_4813,In_1199,In_1646);
nand U4814 (N_4814,In_1359,In_976);
nor U4815 (N_4815,In_697,In_2192);
xor U4816 (N_4816,In_764,In_352);
nand U4817 (N_4817,In_1996,In_822);
nand U4818 (N_4818,In_974,In_1898);
nor U4819 (N_4819,In_332,In_1069);
nor U4820 (N_4820,In_1189,In_1460);
nand U4821 (N_4821,In_1497,In_1278);
nand U4822 (N_4822,In_1070,In_1967);
xor U4823 (N_4823,In_1318,In_2348);
xor U4824 (N_4824,In_1645,In_1602);
nor U4825 (N_4825,In_1170,In_2136);
nand U4826 (N_4826,In_2453,In_893);
xor U4827 (N_4827,In_2306,In_1541);
xor U4828 (N_4828,In_2350,In_1919);
nand U4829 (N_4829,In_129,In_1070);
nor U4830 (N_4830,In_1661,In_2128);
nand U4831 (N_4831,In_963,In_1432);
nand U4832 (N_4832,In_1672,In_2186);
nor U4833 (N_4833,In_1518,In_1432);
xor U4834 (N_4834,In_858,In_323);
or U4835 (N_4835,In_1799,In_1806);
nor U4836 (N_4836,In_936,In_691);
nor U4837 (N_4837,In_2442,In_1067);
xnor U4838 (N_4838,In_2021,In_1037);
nand U4839 (N_4839,In_180,In_2478);
or U4840 (N_4840,In_1122,In_133);
xnor U4841 (N_4841,In_387,In_1688);
xnor U4842 (N_4842,In_1754,In_1606);
nor U4843 (N_4843,In_952,In_235);
and U4844 (N_4844,In_175,In_718);
nand U4845 (N_4845,In_1188,In_2098);
and U4846 (N_4846,In_1307,In_1703);
xor U4847 (N_4847,In_1367,In_1755);
xor U4848 (N_4848,In_590,In_1676);
nor U4849 (N_4849,In_2300,In_1421);
and U4850 (N_4850,In_288,In_2034);
and U4851 (N_4851,In_416,In_799);
or U4852 (N_4852,In_1578,In_186);
and U4853 (N_4853,In_2103,In_985);
nor U4854 (N_4854,In_1948,In_1553);
nand U4855 (N_4855,In_938,In_2372);
and U4856 (N_4856,In_958,In_826);
and U4857 (N_4857,In_49,In_1701);
xor U4858 (N_4858,In_997,In_1168);
and U4859 (N_4859,In_1095,In_1523);
xor U4860 (N_4860,In_84,In_633);
and U4861 (N_4861,In_2022,In_404);
nor U4862 (N_4862,In_1587,In_2133);
or U4863 (N_4863,In_1400,In_1270);
xnor U4864 (N_4864,In_1008,In_1281);
nand U4865 (N_4865,In_2049,In_1315);
or U4866 (N_4866,In_1872,In_844);
nand U4867 (N_4867,In_2088,In_1738);
xor U4868 (N_4868,In_435,In_300);
nor U4869 (N_4869,In_1480,In_2064);
xnor U4870 (N_4870,In_221,In_1153);
xnor U4871 (N_4871,In_1710,In_1329);
nor U4872 (N_4872,In_1851,In_1284);
and U4873 (N_4873,In_1429,In_273);
or U4874 (N_4874,In_606,In_484);
xnor U4875 (N_4875,In_1630,In_2257);
nor U4876 (N_4876,In_181,In_235);
and U4877 (N_4877,In_254,In_2210);
and U4878 (N_4878,In_2363,In_351);
and U4879 (N_4879,In_2020,In_916);
nor U4880 (N_4880,In_339,In_733);
xnor U4881 (N_4881,In_1358,In_1483);
and U4882 (N_4882,In_1960,In_348);
nand U4883 (N_4883,In_232,In_1007);
and U4884 (N_4884,In_945,In_1848);
nor U4885 (N_4885,In_1451,In_594);
and U4886 (N_4886,In_876,In_1894);
or U4887 (N_4887,In_1913,In_2368);
xor U4888 (N_4888,In_2063,In_1473);
nand U4889 (N_4889,In_1170,In_660);
and U4890 (N_4890,In_841,In_2336);
nand U4891 (N_4891,In_2026,In_1300);
or U4892 (N_4892,In_1757,In_2370);
nor U4893 (N_4893,In_1957,In_22);
xnor U4894 (N_4894,In_2274,In_2313);
and U4895 (N_4895,In_963,In_927);
or U4896 (N_4896,In_2493,In_1138);
xor U4897 (N_4897,In_1200,In_1566);
and U4898 (N_4898,In_215,In_3);
nor U4899 (N_4899,In_1713,In_2125);
nor U4900 (N_4900,In_2270,In_824);
or U4901 (N_4901,In_867,In_578);
nor U4902 (N_4902,In_45,In_1227);
xnor U4903 (N_4903,In_1560,In_741);
nor U4904 (N_4904,In_282,In_1354);
xor U4905 (N_4905,In_385,In_2434);
nor U4906 (N_4906,In_2208,In_156);
xnor U4907 (N_4907,In_334,In_412);
xnor U4908 (N_4908,In_2140,In_369);
or U4909 (N_4909,In_1953,In_705);
and U4910 (N_4910,In_1863,In_816);
xnor U4911 (N_4911,In_1156,In_1353);
or U4912 (N_4912,In_477,In_2431);
or U4913 (N_4913,In_243,In_424);
xnor U4914 (N_4914,In_655,In_1805);
nand U4915 (N_4915,In_1591,In_2436);
xor U4916 (N_4916,In_2218,In_1876);
or U4917 (N_4917,In_2311,In_858);
and U4918 (N_4918,In_735,In_1501);
nand U4919 (N_4919,In_182,In_1420);
xor U4920 (N_4920,In_2272,In_2107);
or U4921 (N_4921,In_1261,In_1588);
xnor U4922 (N_4922,In_1404,In_34);
xnor U4923 (N_4923,In_65,In_105);
xnor U4924 (N_4924,In_1206,In_2049);
nor U4925 (N_4925,In_85,In_1128);
nor U4926 (N_4926,In_1815,In_701);
or U4927 (N_4927,In_1236,In_478);
nand U4928 (N_4928,In_1803,In_1673);
and U4929 (N_4929,In_1770,In_2274);
and U4930 (N_4930,In_1732,In_1455);
xnor U4931 (N_4931,In_150,In_2304);
nand U4932 (N_4932,In_152,In_1163);
or U4933 (N_4933,In_571,In_1911);
xor U4934 (N_4934,In_978,In_631);
and U4935 (N_4935,In_1459,In_461);
nand U4936 (N_4936,In_2367,In_1597);
or U4937 (N_4937,In_1536,In_557);
nand U4938 (N_4938,In_2470,In_1018);
nor U4939 (N_4939,In_2148,In_450);
and U4940 (N_4940,In_1882,In_1127);
nand U4941 (N_4941,In_664,In_1400);
or U4942 (N_4942,In_2199,In_1893);
nand U4943 (N_4943,In_2472,In_639);
nand U4944 (N_4944,In_561,In_128);
xnor U4945 (N_4945,In_1264,In_733);
nand U4946 (N_4946,In_1071,In_1899);
or U4947 (N_4947,In_1877,In_1430);
or U4948 (N_4948,In_1838,In_2088);
xnor U4949 (N_4949,In_808,In_1570);
nor U4950 (N_4950,In_69,In_1940);
nor U4951 (N_4951,In_661,In_1105);
and U4952 (N_4952,In_1121,In_747);
nor U4953 (N_4953,In_1500,In_2453);
or U4954 (N_4954,In_744,In_1855);
nand U4955 (N_4955,In_246,In_1345);
or U4956 (N_4956,In_290,In_815);
nand U4957 (N_4957,In_654,In_1473);
nor U4958 (N_4958,In_225,In_391);
or U4959 (N_4959,In_2360,In_2191);
nand U4960 (N_4960,In_1317,In_552);
nand U4961 (N_4961,In_1226,In_2296);
or U4962 (N_4962,In_43,In_335);
nor U4963 (N_4963,In_333,In_468);
and U4964 (N_4964,In_415,In_1058);
xnor U4965 (N_4965,In_1691,In_1677);
or U4966 (N_4966,In_1024,In_1099);
and U4967 (N_4967,In_1092,In_524);
nand U4968 (N_4968,In_122,In_512);
nand U4969 (N_4969,In_162,In_742);
xor U4970 (N_4970,In_450,In_1900);
or U4971 (N_4971,In_2347,In_2187);
or U4972 (N_4972,In_2148,In_941);
nand U4973 (N_4973,In_2451,In_1074);
and U4974 (N_4974,In_2416,In_1036);
or U4975 (N_4975,In_1078,In_1453);
or U4976 (N_4976,In_1527,In_93);
nor U4977 (N_4977,In_2003,In_1817);
and U4978 (N_4978,In_371,In_2274);
nor U4979 (N_4979,In_416,In_311);
xnor U4980 (N_4980,In_2437,In_294);
nand U4981 (N_4981,In_1407,In_108);
nor U4982 (N_4982,In_2318,In_1938);
and U4983 (N_4983,In_880,In_360);
xnor U4984 (N_4984,In_2306,In_946);
nor U4985 (N_4985,In_717,In_306);
and U4986 (N_4986,In_923,In_1429);
nor U4987 (N_4987,In_2073,In_1551);
nor U4988 (N_4988,In_2148,In_397);
xnor U4989 (N_4989,In_2046,In_1779);
xor U4990 (N_4990,In_818,In_1207);
nor U4991 (N_4991,In_2144,In_2098);
nor U4992 (N_4992,In_1229,In_1709);
or U4993 (N_4993,In_1068,In_799);
xnor U4994 (N_4994,In_1804,In_677);
nand U4995 (N_4995,In_429,In_278);
nor U4996 (N_4996,In_1238,In_528);
nor U4997 (N_4997,In_1177,In_247);
or U4998 (N_4998,In_1715,In_1802);
and U4999 (N_4999,In_2414,In_2366);
nor U5000 (N_5000,N_2311,N_4374);
or U5001 (N_5001,N_1849,N_2383);
nand U5002 (N_5002,N_4684,N_4344);
or U5003 (N_5003,N_2784,N_47);
nand U5004 (N_5004,N_2359,N_4595);
or U5005 (N_5005,N_4362,N_3734);
or U5006 (N_5006,N_2476,N_2105);
nand U5007 (N_5007,N_2143,N_3079);
nor U5008 (N_5008,N_3839,N_3856);
nand U5009 (N_5009,N_2252,N_1461);
or U5010 (N_5010,N_4430,N_898);
and U5011 (N_5011,N_2696,N_3254);
nor U5012 (N_5012,N_567,N_114);
nor U5013 (N_5013,N_2795,N_4337);
xor U5014 (N_5014,N_1886,N_2415);
nand U5015 (N_5015,N_1848,N_3260);
nand U5016 (N_5016,N_4030,N_4327);
or U5017 (N_5017,N_1941,N_216);
and U5018 (N_5018,N_857,N_714);
nand U5019 (N_5019,N_2655,N_4198);
or U5020 (N_5020,N_2894,N_853);
xnor U5021 (N_5021,N_3950,N_326);
or U5022 (N_5022,N_1925,N_2686);
nor U5023 (N_5023,N_4321,N_4774);
nor U5024 (N_5024,N_4864,N_4531);
or U5025 (N_5025,N_1757,N_1193);
nor U5026 (N_5026,N_3933,N_1123);
or U5027 (N_5027,N_2702,N_2590);
or U5028 (N_5028,N_4706,N_2613);
xor U5029 (N_5029,N_4471,N_921);
xor U5030 (N_5030,N_1746,N_58);
xnor U5031 (N_5031,N_8,N_1896);
xnor U5032 (N_5032,N_3269,N_1114);
xor U5033 (N_5033,N_1228,N_2422);
and U5034 (N_5034,N_2244,N_4691);
or U5035 (N_5035,N_673,N_4793);
and U5036 (N_5036,N_4074,N_2392);
or U5037 (N_5037,N_2744,N_4623);
nand U5038 (N_5038,N_4933,N_2358);
nor U5039 (N_5039,N_1620,N_4723);
or U5040 (N_5040,N_4508,N_4218);
and U5041 (N_5041,N_2088,N_153);
and U5042 (N_5042,N_1401,N_2939);
nor U5043 (N_5043,N_629,N_4491);
or U5044 (N_5044,N_3581,N_1706);
nand U5045 (N_5045,N_4289,N_4903);
or U5046 (N_5046,N_240,N_3018);
nand U5047 (N_5047,N_2432,N_1214);
nand U5048 (N_5048,N_467,N_977);
or U5049 (N_5049,N_4283,N_3215);
or U5050 (N_5050,N_2023,N_3812);
nor U5051 (N_5051,N_3411,N_3611);
xnor U5052 (N_5052,N_1898,N_1614);
xor U5053 (N_5053,N_980,N_4310);
xnor U5054 (N_5054,N_777,N_760);
nor U5055 (N_5055,N_273,N_3625);
xnor U5056 (N_5056,N_930,N_4637);
xor U5057 (N_5057,N_3474,N_143);
nor U5058 (N_5058,N_1168,N_2460);
and U5059 (N_5059,N_2994,N_3831);
nand U5060 (N_5060,N_185,N_2247);
and U5061 (N_5061,N_141,N_4584);
xnor U5062 (N_5062,N_4827,N_3298);
and U5063 (N_5063,N_3374,N_1295);
and U5064 (N_5064,N_3761,N_1264);
xnor U5065 (N_5065,N_3597,N_3988);
or U5066 (N_5066,N_4567,N_3067);
nand U5067 (N_5067,N_2434,N_2548);
nor U5068 (N_5068,N_4400,N_3667);
nand U5069 (N_5069,N_4000,N_4718);
nand U5070 (N_5070,N_1185,N_171);
or U5071 (N_5071,N_3525,N_4475);
xnor U5072 (N_5072,N_927,N_1675);
nor U5073 (N_5073,N_229,N_965);
nand U5074 (N_5074,N_4085,N_2341);
xor U5075 (N_5075,N_2141,N_1732);
and U5076 (N_5076,N_4216,N_4200);
nor U5077 (N_5077,N_3589,N_1521);
or U5078 (N_5078,N_2833,N_1987);
xnor U5079 (N_5079,N_4311,N_3267);
nand U5080 (N_5080,N_532,N_2623);
nand U5081 (N_5081,N_3913,N_496);
nor U5082 (N_5082,N_4186,N_831);
or U5083 (N_5083,N_3743,N_3570);
xnor U5084 (N_5084,N_1233,N_4973);
nor U5085 (N_5085,N_2324,N_3698);
nor U5086 (N_5086,N_908,N_1206);
and U5087 (N_5087,N_3307,N_786);
or U5088 (N_5088,N_4168,N_2391);
xnor U5089 (N_5089,N_2123,N_1854);
and U5090 (N_5090,N_843,N_1215);
or U5091 (N_5091,N_2877,N_4188);
or U5092 (N_5092,N_1238,N_1314);
and U5093 (N_5093,N_4641,N_4309);
and U5094 (N_5094,N_1218,N_2114);
nand U5095 (N_5095,N_366,N_1667);
nand U5096 (N_5096,N_1663,N_3894);
xor U5097 (N_5097,N_487,N_2474);
or U5098 (N_5098,N_2618,N_3863);
and U5099 (N_5099,N_353,N_307);
xnor U5100 (N_5100,N_2307,N_660);
and U5101 (N_5101,N_2614,N_4214);
and U5102 (N_5102,N_2317,N_133);
nand U5103 (N_5103,N_995,N_4631);
nor U5104 (N_5104,N_1357,N_2718);
or U5105 (N_5105,N_36,N_2478);
and U5106 (N_5106,N_3828,N_489);
and U5107 (N_5107,N_3763,N_4087);
or U5108 (N_5108,N_3131,N_2039);
nand U5109 (N_5109,N_3476,N_2799);
xnor U5110 (N_5110,N_4660,N_1492);
nor U5111 (N_5111,N_493,N_4834);
xor U5112 (N_5112,N_1042,N_3336);
xor U5113 (N_5113,N_4683,N_3769);
or U5114 (N_5114,N_4833,N_3931);
xnor U5115 (N_5115,N_4288,N_4889);
nor U5116 (N_5116,N_4078,N_1782);
or U5117 (N_5117,N_4876,N_984);
nor U5118 (N_5118,N_4225,N_2954);
and U5119 (N_5119,N_4746,N_124);
or U5120 (N_5120,N_2189,N_4043);
xnor U5121 (N_5121,N_1138,N_2427);
or U5122 (N_5122,N_3437,N_2900);
xor U5123 (N_5123,N_2679,N_2031);
xor U5124 (N_5124,N_4788,N_211);
nand U5125 (N_5125,N_4279,N_4921);
xnor U5126 (N_5126,N_2825,N_563);
nor U5127 (N_5127,N_3665,N_25);
and U5128 (N_5128,N_832,N_359);
xor U5129 (N_5129,N_4205,N_4487);
xnor U5130 (N_5130,N_26,N_1255);
nor U5131 (N_5131,N_3952,N_2394);
nand U5132 (N_5132,N_4373,N_3320);
and U5133 (N_5133,N_2801,N_2891);
nand U5134 (N_5134,N_3469,N_1626);
or U5135 (N_5135,N_936,N_4448);
nor U5136 (N_5136,N_2804,N_2689);
nor U5137 (N_5137,N_3429,N_4952);
nand U5138 (N_5138,N_3259,N_2664);
nor U5139 (N_5139,N_361,N_4850);
and U5140 (N_5140,N_2085,N_906);
or U5141 (N_5141,N_687,N_1668);
xnor U5142 (N_5142,N_797,N_3517);
and U5143 (N_5143,N_3112,N_872);
nand U5144 (N_5144,N_4737,N_157);
xnor U5145 (N_5145,N_1093,N_497);
xnor U5146 (N_5146,N_1921,N_4017);
and U5147 (N_5147,N_1810,N_3020);
nor U5148 (N_5148,N_976,N_2274);
nand U5149 (N_5149,N_1652,N_4433);
nor U5150 (N_5150,N_722,N_1120);
and U5151 (N_5151,N_4519,N_2227);
nand U5152 (N_5152,N_4483,N_3833);
and U5153 (N_5153,N_3006,N_1894);
xnor U5154 (N_5154,N_3540,N_3277);
and U5155 (N_5155,N_1633,N_4208);
nor U5156 (N_5156,N_795,N_1355);
nand U5157 (N_5157,N_705,N_3739);
nand U5158 (N_5158,N_1587,N_2916);
xor U5159 (N_5159,N_1767,N_3696);
nor U5160 (N_5160,N_4629,N_2362);
xor U5161 (N_5161,N_880,N_1376);
nand U5162 (N_5162,N_84,N_3163);
or U5163 (N_5163,N_1117,N_2593);
or U5164 (N_5164,N_4410,N_627);
and U5165 (N_5165,N_473,N_2334);
or U5166 (N_5166,N_3998,N_4156);
xor U5167 (N_5167,N_4944,N_1005);
or U5168 (N_5168,N_3255,N_3342);
or U5169 (N_5169,N_4968,N_2643);
nor U5170 (N_5170,N_1707,N_3485);
nand U5171 (N_5171,N_2826,N_1385);
and U5172 (N_5172,N_680,N_4735);
and U5173 (N_5173,N_1531,N_2923);
nand U5174 (N_5174,N_3648,N_1125);
or U5175 (N_5175,N_1473,N_1934);
nor U5176 (N_5176,N_4338,N_2232);
nand U5177 (N_5177,N_769,N_3184);
nand U5178 (N_5178,N_710,N_1323);
nor U5179 (N_5179,N_1060,N_2456);
nand U5180 (N_5180,N_796,N_1805);
and U5181 (N_5181,N_4831,N_4807);
xnor U5182 (N_5182,N_510,N_1300);
xor U5183 (N_5183,N_1992,N_2626);
xnor U5184 (N_5184,N_1680,N_83);
or U5185 (N_5185,N_2024,N_2823);
nor U5186 (N_5186,N_2037,N_1332);
nor U5187 (N_5187,N_807,N_3407);
nand U5188 (N_5188,N_3680,N_1616);
xor U5189 (N_5189,N_778,N_1037);
and U5190 (N_5190,N_1286,N_1544);
nand U5191 (N_5191,N_1474,N_973);
and U5192 (N_5192,N_4932,N_3183);
or U5193 (N_5193,N_3993,N_698);
or U5194 (N_5194,N_2264,N_754);
and U5195 (N_5195,N_674,N_517);
xor U5196 (N_5196,N_882,N_606);
and U5197 (N_5197,N_4233,N_623);
or U5198 (N_5198,N_1421,N_1855);
xnor U5199 (N_5199,N_4565,N_1351);
nand U5200 (N_5200,N_3808,N_334);
and U5201 (N_5201,N_1610,N_416);
nand U5202 (N_5202,N_4387,N_4756);
or U5203 (N_5203,N_2172,N_155);
xnor U5204 (N_5204,N_1662,N_2756);
nand U5205 (N_5205,N_937,N_998);
xnor U5206 (N_5206,N_2015,N_4758);
and U5207 (N_5207,N_3512,N_2814);
nor U5208 (N_5208,N_4420,N_528);
and U5209 (N_5209,N_2872,N_2812);
or U5210 (N_5210,N_4866,N_1009);
nand U5211 (N_5211,N_772,N_1811);
xnor U5212 (N_5212,N_223,N_767);
and U5213 (N_5213,N_2707,N_3296);
xor U5214 (N_5214,N_1289,N_3519);
nor U5215 (N_5215,N_2206,N_2908);
xnor U5216 (N_5216,N_1584,N_1577);
and U5217 (N_5217,N_4947,N_2737);
nand U5218 (N_5218,N_1210,N_3503);
nand U5219 (N_5219,N_2638,N_2766);
xor U5220 (N_5220,N_1787,N_4800);
nor U5221 (N_5221,N_1635,N_2910);
or U5222 (N_5222,N_4426,N_1743);
nand U5223 (N_5223,N_2300,N_397);
or U5224 (N_5224,N_92,N_4719);
nor U5225 (N_5225,N_2061,N_1397);
xnor U5226 (N_5226,N_3608,N_3271);
or U5227 (N_5227,N_1498,N_1151);
nor U5228 (N_5228,N_3225,N_3669);
and U5229 (N_5229,N_2204,N_258);
nand U5230 (N_5230,N_536,N_3069);
or U5231 (N_5231,N_1651,N_524);
nor U5232 (N_5232,N_218,N_4069);
nand U5233 (N_5233,N_782,N_4496);
and U5234 (N_5234,N_2694,N_2741);
or U5235 (N_5235,N_2156,N_4014);
nand U5236 (N_5236,N_390,N_2387);
xnor U5237 (N_5237,N_2722,N_780);
or U5238 (N_5238,N_1755,N_4934);
nor U5239 (N_5239,N_2289,N_3791);
nand U5240 (N_5240,N_3126,N_1001);
or U5241 (N_5241,N_2670,N_2742);
or U5242 (N_5242,N_4731,N_4408);
and U5243 (N_5243,N_3257,N_446);
and U5244 (N_5244,N_2134,N_4114);
nor U5245 (N_5245,N_1362,N_4878);
xnor U5246 (N_5246,N_426,N_958);
xnor U5247 (N_5247,N_2064,N_1287);
and U5248 (N_5248,N_929,N_2082);
nor U5249 (N_5249,N_4484,N_3068);
nand U5250 (N_5250,N_1022,N_424);
nor U5251 (N_5251,N_3562,N_4906);
nand U5252 (N_5252,N_963,N_806);
nand U5253 (N_5253,N_3528,N_3409);
and U5254 (N_5254,N_564,N_2537);
nor U5255 (N_5255,N_1209,N_4058);
xnor U5256 (N_5256,N_1561,N_3160);
xnor U5257 (N_5257,N_1298,N_2897);
and U5258 (N_5258,N_3132,N_2229);
and U5259 (N_5259,N_2688,N_2177);
xnor U5260 (N_5260,N_4281,N_4521);
xnor U5261 (N_5261,N_2410,N_4514);
xor U5262 (N_5262,N_3527,N_3331);
nor U5263 (N_5263,N_2265,N_1163);
and U5264 (N_5264,N_1491,N_2016);
nor U5265 (N_5265,N_3820,N_4231);
and U5266 (N_5266,N_2103,N_2067);
or U5267 (N_5267,N_3287,N_2892);
or U5268 (N_5268,N_942,N_2859);
nand U5269 (N_5269,N_4237,N_3016);
nand U5270 (N_5270,N_715,N_88);
or U5271 (N_5271,N_1660,N_2561);
or U5272 (N_5272,N_4974,N_1970);
and U5273 (N_5273,N_4507,N_2190);
and U5274 (N_5274,N_3561,N_1236);
nand U5275 (N_5275,N_636,N_521);
xnor U5276 (N_5276,N_1570,N_2927);
or U5277 (N_5277,N_2257,N_1137);
nand U5278 (N_5278,N_1033,N_2087);
xnor U5279 (N_5279,N_2312,N_2122);
and U5280 (N_5280,N_1156,N_3560);
nand U5281 (N_5281,N_4398,N_3177);
xor U5282 (N_5282,N_2116,N_2763);
xnor U5283 (N_5283,N_4382,N_2370);
nand U5284 (N_5284,N_2426,N_186);
nor U5285 (N_5285,N_2789,N_3379);
nand U5286 (N_5286,N_1200,N_3951);
nor U5287 (N_5287,N_4460,N_11);
nor U5288 (N_5288,N_3710,N_1337);
and U5289 (N_5289,N_3550,N_1982);
or U5290 (N_5290,N_2651,N_1831);
or U5291 (N_5291,N_725,N_3154);
and U5292 (N_5292,N_2622,N_3681);
xnor U5293 (N_5293,N_1601,N_4154);
nand U5294 (N_5294,N_1965,N_324);
nand U5295 (N_5295,N_896,N_3724);
or U5296 (N_5296,N_888,N_1496);
or U5297 (N_5297,N_1103,N_222);
nand U5298 (N_5298,N_175,N_4312);
nor U5299 (N_5299,N_276,N_672);
nand U5300 (N_5300,N_2621,N_2045);
xor U5301 (N_5301,N_619,N_1960);
or U5302 (N_5302,N_311,N_1179);
nand U5303 (N_5303,N_1551,N_3347);
or U5304 (N_5304,N_1150,N_2231);
xnor U5305 (N_5305,N_4054,N_2302);
nand U5306 (N_5306,N_2647,N_1230);
nor U5307 (N_5307,N_2915,N_638);
and U5308 (N_5308,N_1268,N_1352);
nand U5309 (N_5309,N_3182,N_4005);
nor U5310 (N_5310,N_2163,N_4953);
xor U5311 (N_5311,N_520,N_1371);
xnor U5312 (N_5312,N_4776,N_3719);
and U5313 (N_5313,N_213,N_2092);
xor U5314 (N_5314,N_731,N_4192);
or U5315 (N_5315,N_2620,N_631);
nand U5316 (N_5316,N_4012,N_1052);
or U5317 (N_5317,N_3157,N_2184);
or U5318 (N_5318,N_523,N_3393);
or U5319 (N_5319,N_996,N_1423);
and U5320 (N_5320,N_4651,N_4928);
and U5321 (N_5321,N_21,N_800);
nor U5322 (N_5322,N_2882,N_52);
or U5323 (N_5323,N_3577,N_4948);
and U5324 (N_5324,N_848,N_884);
nor U5325 (N_5325,N_2008,N_4345);
nand U5326 (N_5326,N_957,N_1276);
or U5327 (N_5327,N_3616,N_4326);
nor U5328 (N_5328,N_4232,N_3613);
nand U5329 (N_5329,N_2389,N_4703);
nor U5330 (N_5330,N_3420,N_286);
or U5331 (N_5331,N_2608,N_1526);
and U5332 (N_5332,N_1350,N_3678);
nand U5333 (N_5333,N_4416,N_4379);
or U5334 (N_5334,N_539,N_3238);
nor U5335 (N_5335,N_2076,N_4634);
nor U5336 (N_5336,N_3108,N_3633);
nor U5337 (N_5337,N_4848,N_4429);
nor U5338 (N_5338,N_2893,N_3246);
xor U5339 (N_5339,N_220,N_1629);
or U5340 (N_5340,N_3451,N_3524);
and U5341 (N_5341,N_2830,N_4183);
or U5342 (N_5342,N_4590,N_2332);
xor U5343 (N_5343,N_3899,N_2152);
nand U5344 (N_5344,N_3210,N_1847);
xor U5345 (N_5345,N_4422,N_4015);
nand U5346 (N_5346,N_3859,N_4529);
nor U5347 (N_5347,N_1784,N_50);
nor U5348 (N_5348,N_1760,N_2529);
nand U5349 (N_5349,N_821,N_176);
or U5350 (N_5350,N_4388,N_4882);
xor U5351 (N_5351,N_3504,N_1962);
and U5352 (N_5352,N_126,N_2711);
nand U5353 (N_5353,N_2513,N_2490);
nor U5354 (N_5354,N_379,N_2695);
xnor U5355 (N_5355,N_1866,N_641);
nor U5356 (N_5356,N_1013,N_4658);
xor U5357 (N_5357,N_4927,N_4667);
or U5358 (N_5358,N_2497,N_91);
and U5359 (N_5359,N_3384,N_3941);
nand U5360 (N_5360,N_3236,N_2933);
or U5361 (N_5361,N_3602,N_3072);
or U5362 (N_5362,N_2261,N_1541);
nand U5363 (N_5363,N_3663,N_3115);
and U5364 (N_5364,N_3333,N_1140);
or U5365 (N_5365,N_1945,N_2841);
xnor U5366 (N_5366,N_1862,N_4438);
nor U5367 (N_5367,N_764,N_835);
nand U5368 (N_5368,N_130,N_1549);
xor U5369 (N_5369,N_1924,N_4481);
xnor U5370 (N_5370,N_3980,N_3073);
nor U5371 (N_5371,N_1155,N_1441);
or U5372 (N_5372,N_4956,N_4239);
or U5373 (N_5373,N_465,N_1900);
and U5374 (N_5374,N_3426,N_891);
or U5375 (N_5375,N_3280,N_1598);
or U5376 (N_5376,N_4393,N_4212);
nor U5377 (N_5377,N_112,N_2902);
xor U5378 (N_5378,N_3448,N_62);
nor U5379 (N_5379,N_1061,N_3679);
nand U5380 (N_5380,N_3551,N_3180);
or U5381 (N_5381,N_10,N_3930);
nor U5382 (N_5382,N_3354,N_165);
nand U5383 (N_5383,N_1416,N_2221);
and U5384 (N_5384,N_4525,N_4712);
nor U5385 (N_5385,N_3552,N_3397);
nand U5386 (N_5386,N_4072,N_4645);
nor U5387 (N_5387,N_3310,N_2671);
nor U5388 (N_5388,N_879,N_642);
or U5389 (N_5389,N_2486,N_3684);
nor U5390 (N_5390,N_3687,N_345);
and U5391 (N_5391,N_504,N_2106);
nand U5392 (N_5392,N_3169,N_3065);
and U5393 (N_5393,N_3650,N_4193);
nand U5394 (N_5394,N_4613,N_1603);
xor U5395 (N_5395,N_4897,N_4228);
xor U5396 (N_5396,N_2691,N_4818);
xnor U5397 (N_5397,N_989,N_3646);
and U5398 (N_5398,N_1475,N_1187);
nand U5399 (N_5399,N_1260,N_3450);
nand U5400 (N_5400,N_2027,N_4315);
nor U5401 (N_5401,N_1546,N_2381);
nand U5402 (N_5402,N_2878,N_138);
nor U5403 (N_5403,N_471,N_2555);
nor U5404 (N_5404,N_380,N_2747);
or U5405 (N_5405,N_4185,N_2165);
nor U5406 (N_5406,N_322,N_4498);
or U5407 (N_5407,N_1841,N_615);
xnor U5408 (N_5408,N_3243,N_1888);
and U5409 (N_5409,N_3850,N_2175);
xor U5410 (N_5410,N_242,N_4767);
nand U5411 (N_5411,N_1803,N_1783);
and U5412 (N_5412,N_584,N_3500);
nor U5413 (N_5413,N_1222,N_971);
xor U5414 (N_5414,N_4971,N_4126);
nand U5415 (N_5415,N_1636,N_1208);
or U5416 (N_5416,N_1876,N_4568);
nand U5417 (N_5417,N_555,N_2730);
or U5418 (N_5418,N_1297,N_1948);
nor U5419 (N_5419,N_3111,N_704);
xnor U5420 (N_5420,N_146,N_3113);
nor U5421 (N_5421,N_4517,N_1356);
nor U5422 (N_5422,N_2198,N_3738);
xor U5423 (N_5423,N_2019,N_1802);
nor U5424 (N_5424,N_164,N_414);
or U5425 (N_5425,N_3092,N_1535);
or U5426 (N_5426,N_3935,N_2192);
and U5427 (N_5427,N_1372,N_1065);
nor U5428 (N_5428,N_877,N_855);
and U5429 (N_5429,N_2303,N_779);
and U5430 (N_5430,N_3702,N_2491);
and U5431 (N_5431,N_3505,N_4273);
and U5432 (N_5432,N_1143,N_2790);
or U5433 (N_5433,N_2652,N_907);
nand U5434 (N_5434,N_4226,N_2544);
xnor U5435 (N_5435,N_2319,N_1464);
and U5436 (N_5436,N_3846,N_3226);
or U5437 (N_5437,N_4450,N_3019);
or U5438 (N_5438,N_2805,N_3219);
and U5439 (N_5439,N_1607,N_19);
and U5440 (N_5440,N_3779,N_4655);
xnor U5441 (N_5441,N_708,N_4358);
xnor U5442 (N_5442,N_2551,N_3050);
xnor U5443 (N_5443,N_2329,N_3645);
nand U5444 (N_5444,N_931,N_1861);
or U5445 (N_5445,N_3604,N_2011);
nor U5446 (N_5446,N_3371,N_851);
nor U5447 (N_5447,N_508,N_1688);
nor U5448 (N_5448,N_1919,N_320);
nor U5449 (N_5449,N_1807,N_4992);
nand U5450 (N_5450,N_4900,N_2495);
and U5451 (N_5451,N_2993,N_3799);
nor U5452 (N_5452,N_2769,N_2148);
or U5453 (N_5453,N_607,N_596);
xor U5454 (N_5454,N_509,N_3447);
xor U5455 (N_5455,N_1035,N_2835);
or U5456 (N_5456,N_2179,N_1578);
xor U5457 (N_5457,N_4136,N_1380);
and U5458 (N_5458,N_2539,N_3892);
nor U5459 (N_5459,N_4249,N_4474);
nor U5460 (N_5460,N_2428,N_4802);
nor U5461 (N_5461,N_2568,N_1937);
nor U5462 (N_5462,N_3704,N_2477);
nor U5463 (N_5463,N_2922,N_1413);
and U5464 (N_5464,N_4275,N_1012);
xor U5465 (N_5465,N_4,N_1056);
xnor U5466 (N_5466,N_347,N_1183);
or U5467 (N_5467,N_4624,N_1341);
xnor U5468 (N_5468,N_4190,N_1290);
nor U5469 (N_5469,N_576,N_411);
nor U5470 (N_5470,N_2453,N_4270);
nand U5471 (N_5471,N_2018,N_3502);
nor U5472 (N_5472,N_2225,N_251);
and U5473 (N_5473,N_4144,N_1216);
nand U5474 (N_5474,N_4899,N_1558);
and U5475 (N_5475,N_336,N_3143);
and U5476 (N_5476,N_4317,N_3804);
and U5477 (N_5477,N_4284,N_1487);
nand U5478 (N_5478,N_2339,N_2454);
nand U5479 (N_5479,N_2502,N_2278);
xor U5480 (N_5480,N_2489,N_48);
and U5481 (N_5481,N_2964,N_3634);
and U5482 (N_5482,N_1701,N_4694);
xnor U5483 (N_5483,N_2071,N_4930);
or U5484 (N_5484,N_3355,N_2338);
or U5485 (N_5485,N_4415,N_3725);
xor U5486 (N_5486,N_1991,N_3281);
xor U5487 (N_5487,N_1511,N_3127);
or U5488 (N_5488,N_2136,N_1147);
and U5489 (N_5489,N_1481,N_2880);
xnor U5490 (N_5490,N_1345,N_3455);
nand U5491 (N_5491,N_4151,N_1870);
nor U5492 (N_5492,N_3035,N_3161);
nor U5493 (N_5493,N_2459,N_4621);
nor U5494 (N_5494,N_2547,N_423);
and U5495 (N_5495,N_2108,N_2386);
and U5496 (N_5496,N_2211,N_621);
nor U5497 (N_5497,N_1204,N_4469);
xor U5498 (N_5498,N_2824,N_1983);
nor U5499 (N_5499,N_613,N_970);
nand U5500 (N_5500,N_3489,N_1829);
xor U5501 (N_5501,N_1101,N_3723);
xnor U5502 (N_5502,N_28,N_1665);
xnor U5503 (N_5503,N_71,N_648);
nor U5504 (N_5504,N_3549,N_3882);
nand U5505 (N_5505,N_4561,N_1608);
or U5506 (N_5506,N_2785,N_2308);
and U5507 (N_5507,N_3901,N_2776);
or U5508 (N_5508,N_1694,N_2467);
nor U5509 (N_5509,N_2021,N_4242);
or U5510 (N_5510,N_1926,N_1837);
nor U5511 (N_5511,N_4985,N_2848);
nand U5512 (N_5512,N_3153,N_2736);
or U5513 (N_5513,N_3900,N_40);
nor U5514 (N_5514,N_4763,N_1661);
nand U5515 (N_5515,N_1265,N_1243);
or U5516 (N_5516,N_3903,N_1692);
nand U5517 (N_5517,N_2273,N_1106);
nand U5518 (N_5518,N_2820,N_3);
and U5519 (N_5519,N_4206,N_1762);
nand U5520 (N_5520,N_3506,N_4159);
nand U5521 (N_5521,N_3599,N_3387);
and U5522 (N_5522,N_587,N_4711);
and U5523 (N_5523,N_3797,N_2582);
or U5524 (N_5524,N_140,N_966);
and U5525 (N_5525,N_4562,N_2395);
or U5526 (N_5526,N_2093,N_1806);
or U5527 (N_5527,N_1754,N_1529);
nand U5528 (N_5528,N_4065,N_2077);
xnor U5529 (N_5529,N_3554,N_2838);
and U5530 (N_5530,N_20,N_1878);
xnor U5531 (N_5531,N_3830,N_3647);
xor U5532 (N_5532,N_2619,N_3975);
xor U5533 (N_5533,N_3526,N_2684);
xor U5534 (N_5534,N_243,N_4534);
xor U5535 (N_5535,N_1508,N_4642);
nor U5536 (N_5536,N_1099,N_4830);
nand U5537 (N_5537,N_788,N_2693);
or U5538 (N_5538,N_4923,N_2592);
and U5539 (N_5539,N_2533,N_3746);
xnor U5540 (N_5540,N_4530,N_1655);
nor U5541 (N_5541,N_2762,N_4445);
xor U5542 (N_5542,N_1044,N_734);
nor U5543 (N_5543,N_2276,N_1358);
and U5544 (N_5544,N_3224,N_2286);
or U5545 (N_5545,N_3173,N_2726);
or U5546 (N_5546,N_2199,N_601);
nand U5547 (N_5547,N_659,N_2151);
xor U5548 (N_5548,N_1109,N_4399);
nand U5549 (N_5549,N_585,N_4856);
nor U5550 (N_5550,N_1972,N_4073);
or U5551 (N_5551,N_3195,N_4022);
or U5552 (N_5552,N_2078,N_1440);
and U5553 (N_5553,N_102,N_3178);
or U5554 (N_5554,N_382,N_1766);
and U5555 (N_5555,N_230,N_2305);
nor U5556 (N_5556,N_1325,N_4180);
or U5557 (N_5557,N_476,N_1504);
and U5558 (N_5558,N_4195,N_291);
or U5559 (N_5559,N_4427,N_4598);
nor U5560 (N_5560,N_3410,N_1917);
nor U5561 (N_5561,N_2487,N_878);
or U5562 (N_5562,N_4449,N_2831);
and U5563 (N_5563,N_4732,N_1733);
or U5564 (N_5564,N_2944,N_3413);
and U5565 (N_5565,N_2752,N_3241);
xor U5566 (N_5566,N_4323,N_4976);
and U5567 (N_5567,N_2042,N_3919);
nor U5568 (N_5568,N_282,N_430);
xor U5569 (N_5569,N_4207,N_538);
nor U5570 (N_5570,N_2234,N_2809);
xor U5571 (N_5571,N_3285,N_2003);
and U5572 (N_5572,N_2860,N_4236);
xor U5573 (N_5573,N_4025,N_210);
nand U5574 (N_5574,N_1146,N_1073);
or U5575 (N_5575,N_2480,N_4600);
xor U5576 (N_5576,N_1606,N_199);
nand U5577 (N_5577,N_3249,N_1500);
nor U5578 (N_5578,N_3459,N_679);
xor U5579 (N_5579,N_3836,N_1393);
or U5580 (N_5580,N_4113,N_3816);
nor U5581 (N_5581,N_1051,N_2032);
xor U5582 (N_5582,N_3605,N_3408);
and U5583 (N_5583,N_147,N_329);
xor U5584 (N_5584,N_2157,N_1205);
or U5585 (N_5585,N_3085,N_1769);
or U5586 (N_5586,N_2660,N_1048);
nand U5587 (N_5587,N_1846,N_2301);
or U5588 (N_5588,N_1815,N_979);
nor U5589 (N_5589,N_3340,N_4688);
nor U5590 (N_5590,N_1348,N_2417);
nor U5591 (N_5591,N_3498,N_1301);
xor U5592 (N_5592,N_1293,N_1063);
nor U5593 (N_5593,N_384,N_701);
nor U5594 (N_5594,N_739,N_3801);
and U5595 (N_5595,N_74,N_3025);
or U5596 (N_5596,N_2369,N_905);
and U5597 (N_5597,N_4939,N_3029);
xor U5598 (N_5598,N_4306,N_4581);
xnor U5599 (N_5599,N_3840,N_4537);
and U5600 (N_5600,N_265,N_2251);
nor U5601 (N_5601,N_3295,N_685);
or U5602 (N_5602,N_4988,N_41);
and U5603 (N_5603,N_4693,N_4049);
and U5604 (N_5604,N_2013,N_1986);
or U5605 (N_5605,N_2986,N_516);
nor U5606 (N_5606,N_4504,N_3187);
and U5607 (N_5607,N_2700,N_3706);
nor U5608 (N_5608,N_1826,N_4202);
nand U5609 (N_5609,N_3076,N_3610);
or U5610 (N_5610,N_1553,N_77);
or U5611 (N_5611,N_4247,N_2159);
nand U5612 (N_5612,N_4316,N_1130);
nand U5613 (N_5613,N_1538,N_4032);
or U5614 (N_5614,N_1710,N_3054);
nor U5615 (N_5615,N_2985,N_425);
and U5616 (N_5616,N_1014,N_30);
or U5617 (N_5617,N_1157,N_453);
xor U5618 (N_5618,N_3624,N_4617);
xnor U5619 (N_5619,N_3228,N_914);
nand U5620 (N_5620,N_3214,N_2559);
nand U5621 (N_5621,N_3428,N_304);
nand U5622 (N_5622,N_4341,N_3877);
or U5623 (N_5623,N_4486,N_2699);
and U5624 (N_5624,N_4840,N_4821);
nand U5625 (N_5625,N_2836,N_4219);
nor U5626 (N_5626,N_556,N_4630);
and U5627 (N_5627,N_3100,N_4385);
nor U5628 (N_5628,N_681,N_3538);
and U5629 (N_5629,N_4966,N_1302);
xor U5630 (N_5630,N_1716,N_183);
xnor U5631 (N_5631,N_3439,N_3027);
xnor U5632 (N_5632,N_1003,N_1654);
nor U5633 (N_5633,N_2585,N_4577);
nor U5634 (N_5634,N_4599,N_1429);
nor U5635 (N_5635,N_1158,N_4799);
xor U5636 (N_5636,N_2187,N_2236);
xnor U5637 (N_5637,N_3936,N_2522);
nor U5638 (N_5638,N_652,N_1000);
and U5639 (N_5639,N_2845,N_697);
and U5640 (N_5640,N_1055,N_4874);
nand U5641 (N_5641,N_750,N_558);
and U5642 (N_5642,N_2111,N_3268);
and U5643 (N_5643,N_4161,N_3628);
nand U5644 (N_5644,N_3477,N_870);
nor U5645 (N_5645,N_431,N_248);
nand U5646 (N_5646,N_3252,N_1477);
xnor U5647 (N_5647,N_4130,N_4084);
or U5648 (N_5648,N_2226,N_816);
or U5649 (N_5649,N_2095,N_2240);
nor U5650 (N_5650,N_1391,N_658);
nor U5651 (N_5651,N_4619,N_4877);
nand U5652 (N_5652,N_2966,N_274);
or U5653 (N_5653,N_3304,N_2365);
nor U5654 (N_5654,N_559,N_4860);
and U5655 (N_5655,N_2233,N_2052);
xor U5656 (N_5656,N_3015,N_459);
or U5657 (N_5657,N_2591,N_2917);
nor U5658 (N_5658,N_3405,N_3217);
or U5659 (N_5659,N_4582,N_4583);
nor U5660 (N_5660,N_974,N_4644);
nor U5661 (N_5661,N_4867,N_1340);
nand U5662 (N_5662,N_2352,N_2036);
nor U5663 (N_5663,N_314,N_4252);
nand U5664 (N_5664,N_1879,N_4227);
nor U5665 (N_5665,N_4516,N_2953);
nor U5666 (N_5666,N_4535,N_4785);
nand U5667 (N_5667,N_245,N_1547);
xor U5668 (N_5668,N_2949,N_1838);
or U5669 (N_5669,N_4419,N_1874);
and U5670 (N_5670,N_1560,N_4773);
nand U5671 (N_5671,N_644,N_1993);
nor U5672 (N_5672,N_4666,N_3629);
xor U5673 (N_5673,N_732,N_1374);
nand U5674 (N_5674,N_1967,N_2940);
nor U5675 (N_5675,N_605,N_172);
nand U5676 (N_5676,N_2887,N_849);
nand U5677 (N_5677,N_3683,N_1232);
or U5678 (N_5678,N_4943,N_802);
nor U5679 (N_5679,N_4407,N_1794);
xor U5680 (N_5680,N_4361,N_3579);
or U5681 (N_5681,N_1375,N_190);
and U5682 (N_5682,N_3999,N_3123);
and U5683 (N_5683,N_443,N_4700);
nand U5684 (N_5684,N_2874,N_4446);
nor U5685 (N_5685,N_2787,N_854);
nor U5686 (N_5686,N_2978,N_3400);
xor U5687 (N_5687,N_4772,N_3194);
or U5688 (N_5688,N_1312,N_1657);
or U5689 (N_5689,N_2816,N_66);
nor U5690 (N_5690,N_1964,N_3878);
or U5691 (N_5691,N_2594,N_2363);
xnor U5692 (N_5692,N_460,N_1226);
xnor U5693 (N_5693,N_492,N_3148);
or U5694 (N_5694,N_433,N_4518);
nor U5695 (N_5695,N_773,N_2050);
nand U5696 (N_5696,N_3635,N_1775);
xnor U5697 (N_5697,N_2038,N_4499);
and U5698 (N_5698,N_69,N_2437);
nand U5699 (N_5699,N_4554,N_2068);
and U5700 (N_5700,N_1534,N_2135);
and U5701 (N_5701,N_250,N_1316);
nor U5702 (N_5702,N_2727,N_2249);
xnor U5703 (N_5703,N_2657,N_4266);
xor U5704 (N_5704,N_3446,N_2001);
nor U5705 (N_5705,N_4938,N_2402);
xor U5706 (N_5706,N_4217,N_723);
or U5707 (N_5707,N_2739,N_2617);
nand U5708 (N_5708,N_1167,N_362);
xor U5709 (N_5709,N_4412,N_3651);
and U5710 (N_5710,N_1556,N_2574);
nor U5711 (N_5711,N_4099,N_4477);
or U5712 (N_5712,N_4836,N_1039);
xor U5713 (N_5713,N_4768,N_2757);
nor U5714 (N_5714,N_33,N_12);
xnor U5715 (N_5715,N_972,N_177);
nor U5716 (N_5716,N_1075,N_1944);
or U5717 (N_5717,N_742,N_4787);
and U5718 (N_5718,N_2119,N_3957);
nand U5719 (N_5719,N_3416,N_2290);
xor U5720 (N_5720,N_1721,N_4670);
and U5721 (N_5721,N_2403,N_2270);
nand U5722 (N_5722,N_654,N_4124);
or U5723 (N_5723,N_4575,N_3375);
nor U5724 (N_5724,N_4425,N_499);
and U5725 (N_5725,N_139,N_4298);
and U5726 (N_5726,N_1468,N_389);
nor U5727 (N_5727,N_4869,N_239);
xor U5728 (N_5728,N_1478,N_4910);
and U5729 (N_5729,N_1306,N_1785);
nand U5730 (N_5730,N_1364,N_3244);
nor U5731 (N_5731,N_3879,N_75);
xor U5732 (N_5732,N_3264,N_2633);
xnor U5733 (N_5733,N_3688,N_915);
nand U5734 (N_5734,N_4633,N_3099);
nand U5735 (N_5735,N_3927,N_3363);
and U5736 (N_5736,N_2368,N_2778);
or U5737 (N_5737,N_2147,N_4302);
or U5738 (N_5738,N_932,N_890);
nand U5739 (N_5739,N_4238,N_573);
or U5740 (N_5740,N_346,N_4829);
and U5741 (N_5741,N_4485,N_290);
or U5742 (N_5742,N_3475,N_755);
nand U5743 (N_5743,N_2697,N_4360);
nor U5744 (N_5744,N_18,N_427);
or U5745 (N_5745,N_2484,N_1624);
nor U5746 (N_5746,N_4333,N_2458);
nor U5747 (N_5747,N_275,N_2216);
xor U5748 (N_5748,N_3851,N_811);
and U5749 (N_5749,N_315,N_1928);
or U5750 (N_5750,N_4489,N_610);
nor U5751 (N_5751,N_3961,N_2348);
nand U5752 (N_5752,N_3134,N_3530);
or U5753 (N_5753,N_1905,N_3832);
nand U5754 (N_5754,N_3120,N_2853);
nand U5755 (N_5755,N_2269,N_4784);
or U5756 (N_5756,N_4888,N_814);
nor U5757 (N_5757,N_4588,N_4241);
or U5758 (N_5758,N_1679,N_3104);
or U5759 (N_5759,N_1088,N_2506);
xor U5760 (N_5760,N_4771,N_2755);
xor U5761 (N_5761,N_3837,N_1020);
xnor U5762 (N_5762,N_57,N_4319);
nor U5763 (N_5763,N_859,N_377);
xor U5764 (N_5764,N_1909,N_1324);
xor U5765 (N_5765,N_2945,N_3038);
xnor U5766 (N_5766,N_1175,N_643);
nor U5767 (N_5767,N_4117,N_1571);
nor U5768 (N_5768,N_3796,N_45);
and U5769 (N_5769,N_993,N_668);
nor U5770 (N_5770,N_3086,N_356);
or U5771 (N_5771,N_3391,N_2310);
nor U5772 (N_5772,N_4569,N_2132);
nand U5773 (N_5773,N_3162,N_340);
xnor U5774 (N_5774,N_3205,N_1913);
nor U5775 (N_5775,N_2174,N_97);
nand U5776 (N_5776,N_1822,N_4954);
nand U5777 (N_5777,N_3891,N_2337);
xor U5778 (N_5778,N_2550,N_3574);
nor U5779 (N_5779,N_3897,N_4134);
nor U5780 (N_5780,N_3314,N_2705);
nor U5781 (N_5781,N_3692,N_2740);
or U5782 (N_5782,N_4175,N_2677);
xnor U5783 (N_5783,N_2443,N_1720);
nand U5784 (N_5784,N_2999,N_2377);
or U5785 (N_5785,N_3491,N_3572);
nand U5786 (N_5786,N_1734,N_2656);
nand U5787 (N_5787,N_1197,N_1465);
nand U5788 (N_5788,N_292,N_535);
xnor U5789 (N_5789,N_2208,N_4296);
nand U5790 (N_5790,N_3081,N_4411);
xnor U5791 (N_5791,N_4221,N_2479);
nand U5792 (N_5792,N_4993,N_4563);
nand U5793 (N_5793,N_3872,N_159);
or U5794 (N_5794,N_4152,N_1951);
nor U5795 (N_5795,N_2873,N_3609);
nor U5796 (N_5796,N_264,N_4880);
nand U5797 (N_5797,N_224,N_568);
nor U5798 (N_5798,N_1486,N_938);
nor U5799 (N_5799,N_2262,N_3768);
and U5800 (N_5800,N_2393,N_1084);
or U5801 (N_5801,N_4322,N_4754);
and U5802 (N_5802,N_3920,N_4133);
nand U5803 (N_5803,N_865,N_967);
nor U5804 (N_5804,N_2971,N_1751);
nand U5805 (N_5805,N_2420,N_682);
and U5806 (N_5806,N_4792,N_3303);
and U5807 (N_5807,N_3780,N_2672);
nand U5808 (N_5808,N_491,N_2188);
and U5809 (N_5809,N_4959,N_4984);
nand U5810 (N_5810,N_726,N_3559);
or U5811 (N_5811,N_2983,N_4203);
or U5812 (N_5812,N_2161,N_4359);
nand U5813 (N_5813,N_3094,N_561);
nand U5814 (N_5814,N_1684,N_246);
xnor U5815 (N_5815,N_1390,N_2056);
nand U5816 (N_5816,N_4853,N_4278);
nor U5817 (N_5817,N_418,N_1502);
nand U5818 (N_5818,N_1269,N_3864);
xor U5819 (N_5819,N_2904,N_4402);
or U5820 (N_5820,N_1892,N_3818);
and U5821 (N_5821,N_3757,N_3926);
nor U5822 (N_5822,N_2745,N_2280);
xor U5823 (N_5823,N_299,N_4146);
nor U5824 (N_5824,N_2714,N_3353);
or U5825 (N_5825,N_774,N_4352);
or U5826 (N_5826,N_2284,N_1650);
nand U5827 (N_5827,N_4791,N_3586);
and U5828 (N_5828,N_323,N_272);
xnor U5829 (N_5829,N_3227,N_827);
nand U5830 (N_5830,N_4465,N_1067);
nand U5831 (N_5831,N_707,N_99);
xor U5832 (N_5832,N_1844,N_232);
xor U5833 (N_5833,N_1425,N_1176);
nand U5834 (N_5834,N_4077,N_2586);
nand U5835 (N_5835,N_4002,N_983);
xnor U5836 (N_5836,N_3300,N_2948);
and U5837 (N_5837,N_2010,N_3346);
and U5838 (N_5838,N_4081,N_3248);
and U5839 (N_5839,N_3778,N_934);
nor U5840 (N_5840,N_4304,N_1501);
nor U5841 (N_5841,N_1952,N_4949);
nor U5842 (N_5842,N_635,N_1245);
and U5843 (N_5843,N_4372,N_4805);
and U5844 (N_5844,N_4034,N_4295);
and U5845 (N_5845,N_2988,N_1586);
nand U5846 (N_5846,N_1823,N_3232);
nand U5847 (N_5847,N_4778,N_3440);
or U5848 (N_5848,N_3676,N_1181);
and U5849 (N_5849,N_4125,N_2524);
and U5850 (N_5850,N_2025,N_1462);
nand U5851 (N_5851,N_2463,N_271);
and U5852 (N_5852,N_4677,N_396);
xor U5853 (N_5853,N_3932,N_4704);
nand U5854 (N_5854,N_4162,N_1619);
xnor U5855 (N_5855,N_398,N_4495);
or U5856 (N_5856,N_3388,N_4194);
and U5857 (N_5857,N_137,N_1749);
nor U5858 (N_5858,N_871,N_3731);
nand U5859 (N_5859,N_388,N_3753);
nor U5860 (N_5860,N_1516,N_1873);
nand U5861 (N_5861,N_413,N_4696);
or U5862 (N_5862,N_3003,N_3368);
and U5863 (N_5863,N_4604,N_4614);
or U5864 (N_5864,N_4743,N_4246);
xor U5865 (N_5865,N_1131,N_4605);
nor U5866 (N_5866,N_579,N_3198);
nand U5867 (N_5867,N_226,N_1400);
nor U5868 (N_5868,N_3457,N_4292);
or U5869 (N_5869,N_3861,N_590);
nand U5870 (N_5870,N_2847,N_595);
and U5871 (N_5871,N_3078,N_301);
nand U5872 (N_5872,N_4559,N_3305);
nor U5873 (N_5873,N_696,N_3773);
nand U5874 (N_5874,N_992,N_4040);
or U5875 (N_5875,N_2912,N_784);
xnor U5876 (N_5876,N_458,N_501);
xnor U5877 (N_5877,N_3898,N_2683);
nor U5878 (N_5878,N_3766,N_2867);
xor U5879 (N_5879,N_4436,N_3534);
and U5880 (N_5880,N_1431,N_3977);
xor U5881 (N_5881,N_1115,N_2323);
and U5882 (N_5882,N_3656,N_59);
xnor U5883 (N_5883,N_3486,N_2720);
or U5884 (N_5884,N_1778,N_2104);
nor U5885 (N_5885,N_4849,N_378);
xor U5886 (N_5886,N_4455,N_252);
nand U5887 (N_5887,N_828,N_3666);
xnor U5888 (N_5888,N_1081,N_4894);
nand U5889 (N_5889,N_131,N_1284);
xor U5890 (N_5890,N_1770,N_2576);
or U5891 (N_5891,N_449,N_1852);
nand U5892 (N_5892,N_3370,N_3747);
and U5893 (N_5893,N_287,N_4845);
nand U5894 (N_5894,N_3617,N_2968);
nor U5895 (N_5895,N_3179,N_1235);
xnor U5896 (N_5896,N_881,N_3953);
or U5897 (N_5897,N_2666,N_574);
nand U5898 (N_5898,N_3484,N_60);
or U5899 (N_5899,N_2054,N_1882);
or U5900 (N_5900,N_3720,N_1148);
or U5901 (N_5901,N_4458,N_3063);
nand U5902 (N_5902,N_1484,N_3438);
xor U5903 (N_5903,N_197,N_61);
xnor U5904 (N_5904,N_3427,N_1028);
and U5905 (N_5905,N_161,N_3390);
xnor U5906 (N_5906,N_279,N_3121);
or U5907 (N_5907,N_3944,N_4201);
xor U5908 (N_5908,N_1761,N_2782);
or U5909 (N_5909,N_2120,N_1932);
nand U5910 (N_5910,N_3415,N_2074);
or U5911 (N_5911,N_2865,N_3508);
nor U5912 (N_5912,N_3037,N_3070);
or U5913 (N_5913,N_4452,N_3402);
nor U5914 (N_5914,N_3261,N_3575);
nor U5915 (N_5915,N_1221,N_3740);
or U5916 (N_5916,N_4434,N_4142);
or U5917 (N_5917,N_14,N_4511);
or U5918 (N_5918,N_889,N_4290);
and U5919 (N_5919,N_4008,N_876);
xnor U5920 (N_5920,N_468,N_2531);
nand U5921 (N_5921,N_946,N_2517);
nor U5922 (N_5922,N_4364,N_2941);
or U5923 (N_5923,N_4401,N_3467);
and U5924 (N_5924,N_1463,N_86);
nor U5925 (N_5925,N_333,N_2743);
or U5926 (N_5926,N_1327,N_4942);
nand U5927 (N_5927,N_2538,N_3661);
or U5928 (N_5928,N_4441,N_3708);
xnor U5929 (N_5929,N_2209,N_1880);
nor U5930 (N_5930,N_2072,N_939);
or U5931 (N_5931,N_3658,N_2807);
xor U5932 (N_5932,N_4390,N_4522);
and U5933 (N_5933,N_4902,N_1250);
xor U5934 (N_5934,N_3318,N_3514);
and U5935 (N_5935,N_548,N_1645);
xnor U5936 (N_5936,N_3767,N_1621);
xnor U5937 (N_5937,N_4710,N_3406);
and U5938 (N_5938,N_1656,N_3022);
nand U5939 (N_5939,N_3095,N_4618);
nor U5940 (N_5940,N_2218,N_405);
nor U5941 (N_5941,N_1195,N_3585);
or U5942 (N_5942,N_118,N_2012);
xor U5943 (N_5943,N_1773,N_2382);
or U5944 (N_5944,N_2399,N_1647);
or U5945 (N_5945,N_4095,N_3434);
nor U5946 (N_5946,N_1672,N_3293);
nor U5947 (N_5947,N_663,N_1912);
xnor U5948 (N_5948,N_2808,N_766);
or U5949 (N_5949,N_4736,N_2212);
nor U5950 (N_5950,N_3535,N_4549);
and U5951 (N_5951,N_2678,N_3852);
nor U5952 (N_5952,N_1687,N_920);
and U5953 (N_5953,N_744,N_1703);
or U5954 (N_5954,N_4505,N_589);
nand U5955 (N_5955,N_2889,N_363);
nand U5956 (N_5956,N_4782,N_4417);
and U5957 (N_5957,N_3712,N_89);
or U5958 (N_5958,N_2967,N_1470);
xor U5959 (N_5959,N_3311,N_2802);
and U5960 (N_5960,N_2952,N_1054);
and U5961 (N_5961,N_1087,N_2167);
or U5962 (N_5962,N_3752,N_393);
and U5963 (N_5963,N_3986,N_3984);
xnor U5964 (N_5964,N_1377,N_163);
or U5965 (N_5965,N_4272,N_1234);
nor U5966 (N_5966,N_4409,N_2504);
nor U5967 (N_5967,N_1827,N_1683);
and U5968 (N_5968,N_2662,N_3974);
nor U5969 (N_5969,N_2850,N_1779);
nand U5970 (N_5970,N_2572,N_2430);
and U5971 (N_5971,N_634,N_4539);
nor U5972 (N_5972,N_3316,N_2055);
nand U5973 (N_5973,N_594,N_3216);
xnor U5974 (N_5974,N_794,N_3848);
or U5975 (N_5975,N_761,N_3654);
nor U5976 (N_5976,N_5,N_4267);
xor U5977 (N_5977,N_4813,N_65);
or U5978 (N_5978,N_2842,N_4363);
nor U5979 (N_5979,N_1008,N_3381);
xor U5980 (N_5980,N_1097,N_3359);
nor U5981 (N_5981,N_3135,N_2294);
xnor U5982 (N_5982,N_4503,N_4480);
and U5983 (N_5983,N_3857,N_4354);
nand U5984 (N_5984,N_2612,N_1902);
or U5985 (N_5985,N_1713,N_2183);
xnor U5986 (N_5986,N_1172,N_2788);
and U5987 (N_5987,N_3620,N_944);
and U5988 (N_5988,N_1396,N_3805);
xor U5989 (N_5989,N_3265,N_4204);
and U5990 (N_5990,N_3181,N_991);
and U5991 (N_5991,N_3795,N_1446);
nor U5992 (N_5992,N_950,N_2905);
and U5993 (N_5993,N_4795,N_810);
nand U5994 (N_5994,N_4775,N_2026);
xor U5995 (N_5995,N_196,N_2629);
xnor U5996 (N_5996,N_1360,N_4357);
nor U5997 (N_5997,N_893,N_2315);
and U5998 (N_5998,N_1189,N_100);
or U5999 (N_5999,N_2815,N_2140);
xor U6000 (N_6000,N_2768,N_82);
nor U6001 (N_6001,N_620,N_2729);
xor U6002 (N_6002,N_1171,N_2710);
nand U6003 (N_6003,N_2791,N_1510);
nor U6004 (N_6004,N_1002,N_3051);
nand U6005 (N_6005,N_534,N_3925);
nor U6006 (N_6006,N_789,N_2552);
and U6007 (N_6007,N_1096,N_1567);
and U6008 (N_6008,N_1190,N_2932);
xor U6009 (N_6009,N_3989,N_1808);
nand U6010 (N_6010,N_1279,N_550);
or U6011 (N_6011,N_609,N_3947);
nand U6012 (N_6012,N_1532,N_3614);
and U6013 (N_6013,N_3668,N_758);
xnor U6014 (N_6014,N_81,N_4846);
xnor U6015 (N_6015,N_3497,N_207);
and U6016 (N_6016,N_2911,N_2125);
nor U6017 (N_6017,N_4041,N_2595);
or U6018 (N_6018,N_3571,N_2864);
xor U6019 (N_6019,N_798,N_4962);
or U6020 (N_6020,N_1399,N_2759);
nor U6021 (N_6021,N_770,N_4256);
nand U6022 (N_6022,N_2663,N_2584);
nor U6023 (N_6023,N_688,N_4989);
or U6024 (N_6024,N_1904,N_1664);
nand U6025 (N_6025,N_799,N_2566);
nor U6026 (N_6026,N_2758,N_4697);
or U6027 (N_6027,N_1191,N_4324);
nor U6028 (N_6028,N_1071,N_3921);
nor U6029 (N_6029,N_4570,N_2275);
and U6030 (N_6030,N_474,N_4919);
and U6031 (N_6031,N_1135,N_926);
or U6032 (N_6032,N_3495,N_4890);
nand U6033 (N_6033,N_1648,N_1528);
nor U6034 (N_6034,N_3621,N_4812);
and U6035 (N_6035,N_412,N_597);
nand U6036 (N_6036,N_4680,N_1877);
and U6037 (N_6037,N_1082,N_1127);
nand U6038 (N_6038,N_1819,N_885);
nor U6039 (N_6039,N_2468,N_2347);
xnor U6040 (N_6040,N_3144,N_1451);
nand U6041 (N_6041,N_4612,N_68);
or U6042 (N_6042,N_4018,N_1433);
nor U6043 (N_6043,N_225,N_3880);
xor U6044 (N_6044,N_1469,N_2464);
nand U6045 (N_6045,N_1918,N_572);
nor U6046 (N_6046,N_4961,N_1046);
or U6047 (N_6047,N_3518,N_2378);
nor U6048 (N_6048,N_2094,N_3590);
xor U6049 (N_6049,N_3556,N_4076);
and U6050 (N_6050,N_1700,N_2154);
or U6051 (N_6051,N_3636,N_1644);
nand U6052 (N_6052,N_711,N_3618);
or U6053 (N_6053,N_1995,N_456);
nor U6054 (N_6054,N_1637,N_1110);
or U6055 (N_6055,N_3971,N_4262);
or U6056 (N_6056,N_3566,N_1062);
or U6057 (N_6057,N_2407,N_1581);
nand U6058 (N_6058,N_2081,N_3443);
nor U6059 (N_6059,N_591,N_1812);
nand U6060 (N_6060,N_2020,N_3223);
nor U6061 (N_6061,N_1557,N_4153);
and U6062 (N_6062,N_1402,N_503);
or U6063 (N_6063,N_2146,N_392);
nor U6064 (N_6064,N_3673,N_3785);
nor U6065 (N_6065,N_1029,N_3292);
xor U6066 (N_6066,N_2098,N_4515);
or U6067 (N_6067,N_270,N_4277);
xor U6068 (N_6068,N_1126,N_2771);
or U6069 (N_6069,N_765,N_2903);
and U6070 (N_6070,N_895,N_2318);
nor U6071 (N_6071,N_3970,N_181);
xnor U6072 (N_6072,N_1957,N_1241);
xnor U6073 (N_6073,N_1443,N_3270);
nor U6074 (N_6074,N_4922,N_4047);
xor U6075 (N_6075,N_1404,N_3166);
nand U6076 (N_6076,N_830,N_3150);
xnor U6077 (N_6077,N_3367,N_3881);
and U6078 (N_6078,N_3315,N_3356);
and U6079 (N_6079,N_4166,N_4303);
or U6080 (N_6080,N_2350,N_3943);
xor U6081 (N_6081,N_1045,N_244);
nand U6082 (N_6082,N_3229,N_3907);
nand U6083 (N_6083,N_4726,N_2268);
or U6084 (N_6084,N_2195,N_3671);
nor U6085 (N_6085,N_2316,N_4794);
xor U6086 (N_6086,N_2035,N_331);
or U6087 (N_6087,N_4285,N_956);
and U6088 (N_6088,N_2577,N_1789);
or U6089 (N_6089,N_986,N_2376);
nor U6090 (N_6090,N_4972,N_2505);
nor U6091 (N_6091,N_2283,N_3396);
nand U6092 (N_6092,N_2637,N_3471);
nand U6093 (N_6093,N_1875,N_4646);
nor U6094 (N_6094,N_759,N_3959);
or U6095 (N_6095,N_990,N_1833);
nor U6096 (N_6096,N_2980,N_187);
nand U6097 (N_6097,N_4083,N_267);
and U6098 (N_6098,N_577,N_4187);
nand U6099 (N_6099,N_54,N_4964);
nand U6100 (N_6100,N_228,N_3973);
and U6101 (N_6101,N_4115,N_1455);
or U6102 (N_6102,N_3028,N_4991);
nand U6103 (N_6103,N_2235,N_3060);
nand U6104 (N_6104,N_2746,N_1843);
nor U6105 (N_6105,N_3532,N_4730);
and U6106 (N_6106,N_2043,N_1165);
and U6107 (N_6107,N_3212,N_671);
or U6108 (N_6108,N_2404,N_3902);
or U6109 (N_6109,N_612,N_2063);
xnor U6110 (N_6110,N_1712,N_3090);
nor U6111 (N_6111,N_3843,N_289);
nor U6112 (N_6112,N_1786,N_4139);
or U6113 (N_6113,N_3004,N_1344);
and U6114 (N_6114,N_2009,N_4862);
or U6115 (N_6115,N_1708,N_2005);
or U6116 (N_6116,N_3717,N_3317);
and U6117 (N_6117,N_2224,N_3197);
or U6118 (N_6118,N_1973,N_4107);
nand U6119 (N_6119,N_2961,N_4639);
nor U6120 (N_6120,N_2934,N_2396);
xor U6121 (N_6121,N_4090,N_863);
and U6122 (N_6122,N_2772,N_278);
nand U6123 (N_6123,N_150,N_280);
nand U6124 (N_6124,N_2452,N_1220);
and U6125 (N_6125,N_3329,N_49);
xnor U6126 (N_6126,N_4591,N_649);
nand U6127 (N_6127,N_4061,N_1627);
or U6128 (N_6128,N_2906,N_2130);
nor U6129 (N_6129,N_3911,N_781);
xnor U6130 (N_6130,N_4523,N_2034);
nand U6131 (N_6131,N_4546,N_867);
and U6132 (N_6132,N_419,N_3644);
or U6133 (N_6133,N_3274,N_308);
or U6134 (N_6134,N_402,N_1955);
or U6135 (N_6135,N_3705,N_4325);
nand U6136 (N_6136,N_4643,N_4350);
xnor U6137 (N_6137,N_3091,N_4681);
or U6138 (N_6138,N_3266,N_438);
and U6139 (N_6139,N_3458,N_3501);
xnor U6140 (N_6140,N_3023,N_2271);
or U6141 (N_6141,N_360,N_4493);
or U6142 (N_6142,N_3573,N_4199);
nor U6143 (N_6143,N_4891,N_4585);
nand U6144 (N_6144,N_3075,N_954);
nor U6145 (N_6145,N_639,N_645);
nor U6146 (N_6146,N_1588,N_3118);
nand U6147 (N_6147,N_1998,N_4958);
nor U6148 (N_6148,N_1615,N_4293);
nand U6149 (N_6149,N_1954,N_1457);
nand U6150 (N_6150,N_3968,N_1006);
nand U6151 (N_6151,N_145,N_2075);
nand U6152 (N_6152,N_134,N_27);
nor U6153 (N_6153,N_1697,N_3672);
or U6154 (N_6154,N_4924,N_2914);
and U6155 (N_6155,N_338,N_2253);
xnor U6156 (N_6156,N_4640,N_4045);
xnor U6157 (N_6157,N_3987,N_3385);
nor U6158 (N_6158,N_2041,N_4823);
xor U6159 (N_6159,N_236,N_4979);
and U6160 (N_6160,N_2571,N_4606);
or U6161 (N_6161,N_3730,N_1122);
or U6162 (N_6162,N_4803,N_3382);
or U6163 (N_6163,N_1958,N_624);
or U6164 (N_6164,N_1975,N_2196);
xor U6165 (N_6165,N_3815,N_1548);
xnor U6166 (N_6166,N_4396,N_188);
xnor U6167 (N_6167,N_1476,N_3364);
or U6168 (N_6168,N_1728,N_4728);
nor U6169 (N_6169,N_2958,N_3639);
xnor U6170 (N_6170,N_4179,N_1311);
xnor U6171 (N_6171,N_1,N_743);
or U6172 (N_6172,N_2228,N_1225);
or U6173 (N_6173,N_128,N_2266);
xnor U6174 (N_6174,N_1309,N_3962);
xor U6175 (N_6175,N_3643,N_2107);
and U6176 (N_6176,N_3008,N_3357);
xnor U6177 (N_6177,N_3496,N_1426);
and U6178 (N_6178,N_4094,N_868);
xor U6179 (N_6179,N_4001,N_483);
nand U6180 (N_6180,N_3594,N_234);
and U6181 (N_6181,N_1507,N_381);
nor U6182 (N_6182,N_2543,N_1930);
nand U6183 (N_6183,N_4406,N_1288);
nor U6184 (N_6184,N_4589,N_2436);
nand U6185 (N_6185,N_1435,N_3956);
nor U6186 (N_6186,N_442,N_2079);
and U6187 (N_6187,N_4761,N_2440);
and U6188 (N_6188,N_4263,N_4118);
and U6189 (N_6189,N_2811,N_98);
and U6190 (N_6190,N_4510,N_1069);
or U6191 (N_6191,N_0,N_588);
xnor U6192 (N_6192,N_3955,N_1759);
nand U6193 (N_6193,N_2515,N_650);
nand U6194 (N_6194,N_4053,N_2222);
nor U6195 (N_6195,N_646,N_2998);
xor U6196 (N_6196,N_3313,N_3110);
nand U6197 (N_6197,N_864,N_4798);
or U6198 (N_6198,N_4287,N_3677);
and U6199 (N_6199,N_1495,N_103);
nand U6200 (N_6200,N_9,N_1820);
or U6201 (N_6201,N_120,N_409);
or U6202 (N_6202,N_4229,N_842);
and U6203 (N_6203,N_1261,N_2388);
nand U6204 (N_6204,N_3630,N_2818);
or U6205 (N_6205,N_4137,N_350);
and U6206 (N_6206,N_4339,N_3449);
nor U6207 (N_6207,N_1388,N_825);
nor U6208 (N_6208,N_2855,N_494);
nor U6209 (N_6209,N_2866,N_3741);
nor U6210 (N_6210,N_923,N_4854);
nand U6211 (N_6211,N_195,N_2200);
and U6212 (N_6212,N_3640,N_391);
or U6213 (N_6213,N_3047,N_4442);
or U6214 (N_6214,N_2821,N_2441);
xor U6215 (N_6215,N_3584,N_4026);
or U6216 (N_6216,N_1795,N_3714);
nor U6217 (N_6217,N_2128,N_151);
or U6218 (N_6218,N_4941,N_1144);
and U6219 (N_6219,N_3905,N_951);
nand U6220 (N_6220,N_4838,N_1299);
or U6221 (N_6221,N_2503,N_4080);
xor U6222 (N_6222,N_2084,N_737);
and U6223 (N_6223,N_586,N_1518);
or U6224 (N_6224,N_4123,N_1382);
or U6225 (N_6225,N_4855,N_1800);
nor U6226 (N_6226,N_4527,N_1213);
nand U6227 (N_6227,N_4010,N_410);
nand U6228 (N_6228,N_2685,N_1550);
nand U6229 (N_6229,N_4883,N_997);
or U6230 (N_6230,N_2343,N_571);
nand U6231 (N_6231,N_2322,N_2137);
nand U6232 (N_6232,N_2260,N_3191);
nor U6233 (N_6233,N_2527,N_2786);
or U6234 (N_6234,N_2965,N_4873);
nand U6235 (N_6235,N_4259,N_3803);
xor U6236 (N_6236,N_4729,N_4628);
nand U6237 (N_6237,N_4885,N_4108);
and U6238 (N_6238,N_4828,N_2645);
or U6239 (N_6239,N_1899,N_4822);
nor U6240 (N_6240,N_321,N_3130);
or U6241 (N_6241,N_3158,N_4329);
or U6242 (N_6242,N_281,N_4037);
and U6243 (N_6243,N_1793,N_3507);
and U6244 (N_6244,N_1201,N_4764);
and U6245 (N_6245,N_399,N_3203);
nor U6246 (N_6246,N_2950,N_4024);
or U6247 (N_6247,N_3171,N_4698);
and U6248 (N_6248,N_1253,N_505);
nand U6249 (N_6249,N_3151,N_4987);
nand U6250 (N_6250,N_1936,N_1690);
or U6251 (N_6251,N_1034,N_3889);
and U6252 (N_6252,N_2287,N_2238);
xnor U6253 (N_6253,N_1906,N_383);
nand U6254 (N_6254,N_4926,N_1911);
and U6255 (N_6255,N_2242,N_3233);
nor U6256 (N_6256,N_2895,N_952);
and U6257 (N_6257,N_2682,N_3481);
and U6258 (N_6258,N_2150,N_1968);
nor U6259 (N_6259,N_2258,N_3297);
nand U6260 (N_6260,N_1454,N_179);
and U6261 (N_6261,N_569,N_618);
and U6262 (N_6262,N_1319,N_1649);
nor U6263 (N_6263,N_3299,N_1895);
nor U6264 (N_6264,N_3478,N_3456);
xnor U6265 (N_6265,N_1040,N_3749);
nand U6266 (N_6266,N_2803,N_4067);
nand U6267 (N_6267,N_490,N_2390);
nor U6268 (N_6268,N_4870,N_2044);
nand U6269 (N_6269,N_3083,N_3289);
or U6270 (N_6270,N_526,N_3199);
xor U6271 (N_6271,N_4673,N_2255);
or U6272 (N_6272,N_4692,N_3854);
nand U6273 (N_6273,N_4770,N_3211);
nor U6274 (N_6274,N_4121,N_746);
or U6275 (N_6275,N_4593,N_2138);
nor U6276 (N_6276,N_506,N_4392);
and U6277 (N_6277,N_3032,N_2419);
nand U6278 (N_6278,N_3258,N_713);
nand U6279 (N_6279,N_3771,N_3939);
and U6280 (N_6280,N_677,N_2588);
xor U6281 (N_6281,N_2797,N_4742);
nand U6282 (N_6282,N_4075,N_1494);
and U6283 (N_6283,N_132,N_237);
nor U6284 (N_6284,N_1308,N_3155);
or U6285 (N_6285,N_3234,N_479);
xor U6286 (N_6286,N_4375,N_1519);
and U6287 (N_6287,N_2979,N_4781);
or U6288 (N_6288,N_2931,N_691);
or U6289 (N_6289,N_3546,N_2509);
nand U6290 (N_6290,N_87,N_4951);
xnor U6291 (N_6291,N_2049,N_2272);
xnor U6292 (N_6292,N_1752,N_184);
xor U6293 (N_6293,N_4555,N_2549);
xnor U6294 (N_6294,N_2017,N_2060);
xnor U6295 (N_6295,N_2599,N_2277);
nor U6296 (N_6296,N_1835,N_962);
and U6297 (N_6297,N_4940,N_4169);
nand U6298 (N_6298,N_2627,N_4608);
and U6299 (N_6299,N_1428,N_3824);
and U6300 (N_6300,N_2411,N_4428);
nand U6301 (N_6301,N_4020,N_1244);
or U6302 (N_6302,N_3093,N_2553);
or U6303 (N_6303,N_1851,N_502);
and U6304 (N_6304,N_332,N_1333);
or U6305 (N_6305,N_1996,N_1666);
xor U6306 (N_6306,N_4044,N_4576);
xor U6307 (N_6307,N_1517,N_2913);
xnor U6308 (N_6308,N_2051,N_3096);
and U6309 (N_6309,N_507,N_1194);
nand U6310 (N_6310,N_4421,N_3533);
xnor U6311 (N_6311,N_604,N_1594);
or U6312 (N_6312,N_4636,N_3945);
or U6313 (N_6313,N_415,N_4257);
or U6314 (N_6314,N_3755,N_4300);
and U6315 (N_6315,N_440,N_374);
nand U6316 (N_6316,N_3001,N_4937);
nand U6317 (N_6317,N_530,N_1489);
xnor U6318 (N_6318,N_2047,N_2121);
or U6319 (N_6319,N_4033,N_1537);
xor U6320 (N_6320,N_537,N_3494);
nand U6321 (N_6321,N_2924,N_2540);
nand U6322 (N_6322,N_3479,N_4431);
nor U6323 (N_6323,N_3923,N_3691);
xor U6324 (N_6324,N_198,N_664);
or U6325 (N_6325,N_3810,N_4986);
nor U6326 (N_6326,N_3792,N_4547);
nand U6327 (N_6327,N_4865,N_2615);
or U6328 (N_6328,N_1296,N_3652);
xor U6329 (N_6329,N_4592,N_1791);
nor U6330 (N_6330,N_4007,N_2062);
and U6331 (N_6331,N_2542,N_2640);
or U6332 (N_6332,N_3383,N_3052);
xor U6333 (N_6333,N_3464,N_614);
xnor U6334 (N_6334,N_4622,N_4690);
or U6335 (N_6335,N_1180,N_2798);
and U6336 (N_6336,N_1107,N_238);
or U6337 (N_6337,N_1980,N_1479);
xnor U6338 (N_6338,N_3967,N_2641);
nand U6339 (N_6339,N_2256,N_3694);
xor U6340 (N_6340,N_525,N_1410);
nor U6341 (N_6341,N_1134,N_4171);
nor U6342 (N_6342,N_3569,N_349);
nor U6343 (N_6343,N_625,N_1612);
nand U6344 (N_6344,N_3139,N_1080);
or U6345 (N_6345,N_1686,N_3940);
nor U6346 (N_6346,N_4995,N_1719);
nor U6347 (N_6347,N_6,N_3414);
xor U6348 (N_6348,N_2709,N_253);
and U6349 (N_6349,N_2472,N_4935);
nor U6350 (N_6350,N_4815,N_975);
xor U6351 (N_6351,N_1611,N_3098);
and U6352 (N_6352,N_2754,N_3064);
or U6353 (N_6353,N_2501,N_1430);
xnor U6354 (N_6354,N_495,N_3213);
nand U6355 (N_6355,N_1015,N_3376);
xnor U6356 (N_6356,N_3841,N_1872);
and U6357 (N_6357,N_1622,N_981);
nor U6358 (N_6358,N_709,N_182);
xor U6359 (N_6359,N_3809,N_1074);
nor U6360 (N_6360,N_551,N_3909);
nor U6361 (N_6361,N_3784,N_3176);
xnor U6362 (N_6362,N_2033,N_1922);
and U6363 (N_6363,N_543,N_1963);
xnor U6364 (N_6364,N_892,N_4950);
nand U6365 (N_6365,N_3733,N_2281);
xnor U6366 (N_6366,N_3659,N_1025);
xor U6367 (N_6367,N_1320,N_3709);
xnor U6368 (N_6368,N_435,N_3136);
xnor U6369 (N_6369,N_2733,N_2385);
or U6370 (N_6370,N_4674,N_4757);
xor U6371 (N_6371,N_174,N_4777);
or U6372 (N_6372,N_4100,N_4196);
nand U6373 (N_6373,N_1623,N_3145);
nand U6374 (N_6374,N_17,N_3567);
nand U6375 (N_6375,N_4189,N_3034);
xnor U6376 (N_6376,N_562,N_3606);
nor U6377 (N_6377,N_1321,N_2854);
nand U6378 (N_6378,N_123,N_1513);
and U6379 (N_6379,N_2676,N_3576);
or U6380 (N_6380,N_3838,N_1671);
xnor U6381 (N_6381,N_1251,N_3306);
nand U6382 (N_6382,N_189,N_1969);
nand U6383 (N_6383,N_4335,N_1953);
nor U6384 (N_6384,N_692,N_1098);
or U6385 (N_6385,N_4716,N_1058);
and U6386 (N_6386,N_2560,N_4820);
or U6387 (N_6387,N_498,N_2987);
or U6388 (N_6388,N_2920,N_4104);
nor U6389 (N_6389,N_2673,N_452);
nand U6390 (N_6390,N_4064,N_860);
nand U6391 (N_6391,N_1329,N_1166);
or U6392 (N_6392,N_2990,N_1595);
or U6393 (N_6393,N_1405,N_4245);
nand U6394 (N_6394,N_720,N_325);
nand U6395 (N_6395,N_804,N_78);
and U6396 (N_6396,N_847,N_1506);
and U6397 (N_6397,N_4616,N_4093);
or U6398 (N_6398,N_833,N_2485);
or U6399 (N_6399,N_3220,N_2708);
and U6400 (N_6400,N_4843,N_2288);
xor U6401 (N_6401,N_1303,N_51);
nor U6402 (N_6402,N_3338,N_2962);
or U6403 (N_6403,N_4454,N_1085);
nand U6404 (N_6404,N_1335,N_3462);
and U6405 (N_6405,N_3380,N_22);
and U6406 (N_6406,N_1493,N_763);
and U6407 (N_6407,N_570,N_4762);
xor U6408 (N_6408,N_1047,N_1722);
nand U6409 (N_6409,N_4824,N_4620);
xor U6410 (N_6410,N_4378,N_3595);
xor U6411 (N_6411,N_3934,N_2351);
xor U6412 (N_6412,N_2837,N_1499);
nor U6413 (N_6413,N_4440,N_4671);
nand U6414 (N_6414,N_1745,N_875);
nor U6415 (N_6415,N_312,N_3273);
xnor U6416 (N_6416,N_3545,N_1642);
xor U6417 (N_6417,N_1349,N_1839);
xor U6418 (N_6418,N_1154,N_700);
and U6419 (N_6419,N_1153,N_655);
xnor U6420 (N_6420,N_2494,N_4557);
nand U6421 (N_6421,N_3906,N_1273);
xor U6422 (N_6422,N_4209,N_4573);
nor U6423 (N_6423,N_4369,N_2601);
nor U6424 (N_6424,N_935,N_3834);
xor U6425 (N_6425,N_358,N_4297);
xor U6426 (N_6426,N_1338,N_1609);
nor U6427 (N_6427,N_4603,N_2510);
nand U6428 (N_6428,N_3783,N_4258);
and U6429 (N_6429,N_2400,N_23);
nand U6430 (N_6430,N_2587,N_2153);
and U6431 (N_6431,N_1094,N_1102);
or U6432 (N_6432,N_933,N_53);
and U6433 (N_6433,N_3759,N_1903);
nand U6434 (N_6434,N_1108,N_1883);
and U6435 (N_6435,N_3432,N_46);
nor U6436 (N_6436,N_2610,N_1389);
nand U6437 (N_6437,N_2483,N_3835);
and U6438 (N_6438,N_818,N_1272);
nor U6439 (N_6439,N_1453,N_3386);
and U6440 (N_6440,N_1639,N_4170);
nand U6441 (N_6441,N_3728,N_298);
nand U6442 (N_6442,N_3924,N_4230);
xnor U6443 (N_6443,N_2360,N_2665);
and U6444 (N_6444,N_354,N_3140);
or U6445 (N_6445,N_4432,N_4235);
nand U6446 (N_6446,N_531,N_4857);
or U6447 (N_6447,N_4244,N_2002);
and U6448 (N_6448,N_2648,N_96);
and U6449 (N_6449,N_961,N_3056);
or U6450 (N_6450,N_3874,N_1813);
nand U6451 (N_6451,N_719,N_721);
or U6452 (N_6452,N_4804,N_2888);
nor U6453 (N_6453,N_1142,N_3002);
and U6454 (N_6454,N_4602,N_2567);
nand U6455 (N_6455,N_1407,N_2004);
and U6456 (N_6456,N_3327,N_628);
and U6457 (N_6457,N_204,N_4211);
or U6458 (N_6458,N_518,N_3722);
and U6459 (N_6459,N_729,N_2445);
or U6460 (N_6460,N_2578,N_167);
xor U6461 (N_6461,N_343,N_1116);
and U6462 (N_6462,N_2876,N_1893);
xnor U6463 (N_6463,N_1160,N_1522);
and U6464 (N_6464,N_3463,N_3726);
nor U6465 (N_6465,N_169,N_4308);
and U6466 (N_6466,N_1274,N_1990);
xor U6467 (N_6467,N_599,N_4872);
or U6468 (N_6468,N_1774,N_3963);
nor U6469 (N_6469,N_1979,N_3916);
and U6470 (N_6470,N_469,N_4351);
or U6471 (N_6471,N_1041,N_3829);
nand U6472 (N_6472,N_2997,N_3873);
nor U6473 (N_6473,N_2525,N_4042);
and U6474 (N_6474,N_1442,N_4750);
nor U6475 (N_6475,N_3915,N_1427);
xnor U6476 (N_6476,N_1676,N_4395);
and U6477 (N_6477,N_4467,N_2447);
and U6478 (N_6478,N_3742,N_3811);
nand U6479 (N_6479,N_4753,N_1593);
and U6480 (N_6480,N_2201,N_2712);
or U6481 (N_6481,N_4003,N_3750);
and U6482 (N_6482,N_1505,N_866);
xnor U6483 (N_6483,N_2444,N_2030);
xor U6484 (N_6484,N_3789,N_3543);
nand U6485 (N_6485,N_3071,N_2058);
or U6486 (N_6486,N_910,N_4502);
nor U6487 (N_6487,N_2439,N_3565);
nand U6488 (N_6488,N_3122,N_3884);
nor U6489 (N_6489,N_695,N_4470);
nor U6490 (N_6490,N_1989,N_1186);
nand U6491 (N_6491,N_1277,N_519);
xor U6492 (N_6492,N_1378,N_2493);
or U6493 (N_6493,N_4320,N_3867);
and U6494 (N_6494,N_3084,N_4663);
nor U6495 (N_6495,N_3592,N_1574);
nand U6496 (N_6496,N_1702,N_1693);
nor U6497 (N_6497,N_3777,N_3030);
xnor U6498 (N_6498,N_3328,N_3200);
or U6499 (N_6499,N_39,N_2995);
nor U6500 (N_6500,N_1092,N_4101);
or U6501 (N_6501,N_3209,N_2898);
nor U6502 (N_6502,N_3221,N_2083);
xnor U6503 (N_6503,N_1539,N_370);
xnor U6504 (N_6504,N_3716,N_2295);
or U6505 (N_6505,N_1869,N_106);
xor U6506 (N_6506,N_3583,N_3129);
or U6507 (N_6507,N_4881,N_35);
or U6508 (N_6508,N_554,N_4473);
xor U6509 (N_6509,N_2886,N_919);
nand U6510 (N_6510,N_2602,N_4911);
nand U6511 (N_6511,N_63,N_689);
nor U6512 (N_6512,N_4384,N_2096);
and U6513 (N_6513,N_4975,N_792);
and U6514 (N_6514,N_4488,N_4574);
or U6515 (N_6515,N_1417,N_3515);
and U6516 (N_6516,N_2069,N_1907);
xor U6517 (N_6517,N_3675,N_4466);
and U6518 (N_6518,N_2717,N_2581);
xor U6519 (N_6519,N_2455,N_1867);
or U6520 (N_6520,N_3822,N_745);
nor U6521 (N_6521,N_2649,N_4028);
xor U6522 (N_6522,N_296,N_1592);
and U6523 (N_6523,N_4334,N_4587);
or U6524 (N_6524,N_4965,N_2164);
xor U6525 (N_6525,N_1436,N_1007);
nand U6526 (N_6526,N_4625,N_3403);
or U6527 (N_6527,N_342,N_1076);
xor U6528 (N_6528,N_3937,N_2977);
nor U6529 (N_6529,N_1381,N_3849);
xor U6530 (N_6530,N_834,N_170);
and U6531 (N_6531,N_261,N_1533);
xnor U6532 (N_6532,N_42,N_1890);
or U6533 (N_6533,N_1342,N_2241);
nor U6534 (N_6534,N_2658,N_1940);
nor U6535 (N_6535,N_3764,N_740);
nand U6536 (N_6536,N_3703,N_4999);
xnor U6537 (N_6537,N_1370,N_1354);
nand U6538 (N_6538,N_540,N_3701);
nand U6539 (N_6539,N_2749,N_1845);
nand U6540 (N_6540,N_1780,N_762);
nor U6541 (N_6541,N_337,N_3326);
or U6542 (N_6542,N_3756,N_4886);
or U6543 (N_6543,N_447,N_2416);
xnor U6544 (N_6544,N_2203,N_233);
and U6545 (N_6545,N_1977,N_4301);
and U6546 (N_6546,N_2796,N_2519);
nand U6547 (N_6547,N_4342,N_1555);
and U6548 (N_6548,N_2406,N_1790);
and U6549 (N_6549,N_4901,N_464);
nor U6550 (N_6550,N_1409,N_3417);
xnor U6551 (N_6551,N_2178,N_3010);
or U6552 (N_6552,N_904,N_3107);
nor U6553 (N_6553,N_511,N_4250);
or U6554 (N_6554,N_2180,N_3017);
nor U6555 (N_6555,N_1192,N_406);
nor U6556 (N_6556,N_3876,N_2523);
xor U6557 (N_6557,N_4983,N_217);
xnor U6558 (N_6558,N_4745,N_4268);
xnor U6559 (N_6559,N_3480,N_4394);
nor U6560 (N_6560,N_1857,N_2073);
or U6561 (N_6561,N_4665,N_3910);
and U6562 (N_6562,N_1458,N_2057);
nor U6563 (N_6563,N_1580,N_4540);
xnor U6564 (N_6564,N_3425,N_1856);
and U6565 (N_6565,N_4528,N_3352);
and U6566 (N_6566,N_1090,N_1439);
nor U6567 (N_6567,N_2938,N_1961);
nand U6568 (N_6568,N_987,N_616);
or U6569 (N_6569,N_717,N_454);
or U6570 (N_6570,N_3553,N_1248);
xor U6571 (N_6571,N_2644,N_1520);
or U6572 (N_6572,N_3745,N_4861);
or U6573 (N_6573,N_4164,N_344);
nand U6574 (N_6574,N_3853,N_461);
and U6575 (N_6575,N_3012,N_4553);
nand U6576 (N_6576,N_4414,N_4669);
or U6577 (N_6577,N_372,N_2100);
and U6578 (N_6578,N_4063,N_1366);
and U6579 (N_6579,N_4814,N_3192);
and U6580 (N_6580,N_656,N_1935);
xnor U6581 (N_6581,N_247,N_3235);
xor U6582 (N_6582,N_2628,N_757);
xnor U6583 (N_6583,N_1334,N_4255);
nand U6584 (N_6584,N_219,N_1043);
nand U6585 (N_6585,N_2423,N_3825);
and U6586 (N_6586,N_4490,N_2);
or U6587 (N_6587,N_1792,N_2059);
nor U6588 (N_6588,N_2115,N_4128);
nor U6589 (N_6589,N_2007,N_1984);
or U6590 (N_6590,N_3057,N_330);
or U6591 (N_6591,N_1978,N_110);
nor U6592 (N_6592,N_776,N_4520);
nor U6593 (N_6593,N_2214,N_3398);
xnor U6594 (N_6594,N_1368,N_1411);
or U6595 (N_6595,N_420,N_2751);
and U6596 (N_6596,N_4029,N_1384);
nor U6597 (N_6597,N_4062,N_4340);
or U6598 (N_6598,N_3541,N_3168);
xnor U6599 (N_6599,N_4538,N_3788);
and U6600 (N_6600,N_4844,N_2346);
nor U6601 (N_6601,N_209,N_1735);
nand U6602 (N_6602,N_4163,N_3389);
and U6603 (N_6603,N_4721,N_4722);
and U6604 (N_6604,N_2182,N_1017);
nor U6605 (N_6605,N_3682,N_1403);
or U6606 (N_6606,N_3954,N_3994);
or U6607 (N_6607,N_3964,N_2397);
xnor U6608 (N_6608,N_2863,N_2777);
nor U6609 (N_6609,N_73,N_712);
nor U6610 (N_6610,N_2960,N_4808);
and U6611 (N_6611,N_72,N_1678);
or U6612 (N_6612,N_617,N_1240);
nand U6613 (N_6613,N_4148,N_2006);
nand U6614 (N_6614,N_208,N_1386);
or U6615 (N_6615,N_513,N_2972);
nand U6616 (N_6616,N_1136,N_2438);
and U6617 (N_6617,N_1641,N_3424);
nor U6618 (N_6618,N_2674,N_3309);
nor U6619 (N_6619,N_2207,N_2331);
nand U6620 (N_6620,N_294,N_1605);
nor U6621 (N_6621,N_1572,N_1118);
xor U6622 (N_6622,N_899,N_2937);
nand U6623 (N_6623,N_2817,N_4524);
nand U6624 (N_6624,N_3372,N_3591);
or U6625 (N_6625,N_4269,N_2521);
nor U6626 (N_6626,N_2557,N_109);
xor U6627 (N_6627,N_4858,N_191);
and U6628 (N_6628,N_2706,N_3547);
xor U6629 (N_6629,N_4271,N_3460);
and U6630 (N_6630,N_1853,N_375);
or U6631 (N_6631,N_3435,N_4668);
or U6632 (N_6632,N_4918,N_4705);
nor U6633 (N_6633,N_4817,N_3729);
or U6634 (N_6634,N_4036,N_335);
nor U6635 (N_6635,N_1658,N_2661);
nand U6636 (N_6636,N_4155,N_1415);
and U6637 (N_6637,N_2435,N_4752);
or U6638 (N_6638,N_4119,N_3563);
and U6639 (N_6639,N_310,N_1741);
and U6640 (N_6640,N_592,N_1322);
nor U6641 (N_6641,N_4089,N_4996);
or U6642 (N_6642,N_817,N_791);
xor U6643 (N_6643,N_3253,N_2409);
nand U6644 (N_6644,N_837,N_328);
nor U6645 (N_6645,N_480,N_2750);
nand U6646 (N_6646,N_2947,N_2133);
xor U6647 (N_6647,N_1801,N_1164);
and U6648 (N_6648,N_1885,N_1596);
xor U6649 (N_6649,N_2605,N_2230);
nand U6650 (N_6650,N_1939,N_1599);
xor U6651 (N_6651,N_1207,N_2296);
or U6652 (N_6652,N_913,N_2461);
nand U6653 (N_6653,N_3330,N_4896);
or U6654 (N_6654,N_3021,N_1089);
and U6655 (N_6655,N_844,N_214);
or U6656 (N_6656,N_4556,N_2800);
nor U6657 (N_6657,N_1689,N_3529);
nand U6658 (N_6658,N_4079,N_348);
nor U6659 (N_6659,N_4916,N_1174);
or U6660 (N_6660,N_1582,N_235);
nand U6661 (N_6661,N_647,N_3807);
xnor U6662 (N_6662,N_3344,N_1078);
or U6663 (N_6663,N_3695,N_4343);
nor U6664 (N_6664,N_667,N_3845);
and U6665 (N_6665,N_4887,N_736);
and U6666 (N_6666,N_3077,N_2545);
nor U6667 (N_6667,N_4141,N_1602);
nor U6668 (N_6668,N_545,N_3088);
nand U6669 (N_6669,N_4609,N_1949);
nand U6670 (N_6670,N_3377,N_1211);
or U6671 (N_6671,N_3433,N_2091);
nand U6672 (N_6672,N_3146,N_1483);
nor U6673 (N_6673,N_533,N_1938);
and U6674 (N_6674,N_262,N_1777);
and U6675 (N_6675,N_3523,N_3102);
and U6676 (N_6676,N_4879,N_4251);
or U6677 (N_6677,N_3242,N_1395);
or U6678 (N_6678,N_3031,N_1564);
nand U6679 (N_6679,N_2374,N_4157);
nor U6680 (N_6680,N_3046,N_4727);
nor U6681 (N_6681,N_3821,N_3369);
xor U6682 (N_6682,N_2046,N_1943);
and U6683 (N_6683,N_1696,N_1600);
nand U6684 (N_6684,N_2704,N_3557);
nor U6685 (N_6685,N_3548,N_1729);
or U6686 (N_6686,N_142,N_2775);
nor U6687 (N_6687,N_3638,N_4371);
and U6688 (N_6688,N_249,N_2896);
and U6689 (N_6689,N_3978,N_3655);
nor U6690 (N_6690,N_2963,N_2239);
nand U6691 (N_6691,N_787,N_3990);
nand U6692 (N_6692,N_4512,N_4165);
or U6693 (N_6693,N_2534,N_462);
xnor U6694 (N_6694,N_3868,N_4868);
or U6695 (N_6695,N_1536,N_1889);
nand U6696 (N_6696,N_168,N_3786);
nor U6697 (N_6697,N_2541,N_4702);
nand U6698 (N_6698,N_115,N_3172);
and U6699 (N_6699,N_395,N_3442);
nand U6700 (N_6700,N_206,N_2327);
xnor U6701 (N_6701,N_4478,N_3751);
nor U6702 (N_6702,N_1618,N_1257);
nor U6703 (N_6703,N_3862,N_1188);
and U6704 (N_6704,N_3700,N_675);
xor U6705 (N_6705,N_4066,N_355);
or U6706 (N_6706,N_4656,N_1748);
or U6707 (N_6707,N_897,N_1929);
and U6708 (N_6708,N_448,N_4626);
nand U6709 (N_6709,N_661,N_3674);
or U6710 (N_6710,N_809,N_3817);
and U6711 (N_6711,N_2398,N_2942);
or U6712 (N_6712,N_3908,N_3544);
and U6713 (N_6713,N_2171,N_2884);
and U6714 (N_6714,N_2418,N_3802);
and U6715 (N_6715,N_2220,N_44);
nor U6716 (N_6716,N_1514,N_4661);
or U6717 (N_6717,N_1715,N_1653);
nor U6718 (N_6718,N_2881,N_162);
nand U6719 (N_6719,N_4895,N_2469);
nor U6720 (N_6720,N_3542,N_640);
or U6721 (N_6721,N_4331,N_3013);
or U6722 (N_6722,N_2883,N_522);
nor U6723 (N_6723,N_3521,N_775);
nand U6724 (N_6724,N_70,N_2951);
or U6725 (N_6725,N_1064,N_3653);
nor U6726 (N_6726,N_385,N_2792);
nor U6727 (N_6727,N_4627,N_4149);
nor U6728 (N_6728,N_1383,N_4960);
xor U6729 (N_6729,N_2223,N_1018);
xor U6730 (N_6730,N_4435,N_466);
and U6731 (N_6731,N_999,N_2372);
xnor U6732 (N_6732,N_180,N_1418);
or U6733 (N_6733,N_598,N_1049);
nand U6734 (N_6734,N_2110,N_4013);
or U6735 (N_6735,N_2996,N_2526);
and U6736 (N_6736,N_3847,N_3765);
or U6737 (N_6737,N_4459,N_144);
xor U6738 (N_6738,N_135,N_1414);
or U6739 (N_6739,N_436,N_1315);
nand U6740 (N_6740,N_978,N_753);
nor U6741 (N_6741,N_1966,N_1740);
xnor U6742 (N_6742,N_2481,N_3421);
nand U6743 (N_6743,N_4367,N_3164);
nand U6744 (N_6744,N_4070,N_1231);
nand U6745 (N_6745,N_417,N_3490);
nor U6746 (N_6746,N_2819,N_2611);
and U6747 (N_6747,N_4182,N_2099);
and U6748 (N_6748,N_3312,N_3218);
and U6749 (N_6749,N_3465,N_305);
and U6750 (N_6750,N_4526,N_1613);
nand U6751 (N_6751,N_2144,N_125);
and U6752 (N_6752,N_127,N_4875);
xnor U6753 (N_6753,N_4955,N_2909);
nor U6754 (N_6754,N_2668,N_2616);
nand U6755 (N_6755,N_894,N_2291);
or U6756 (N_6756,N_3972,N_2982);
or U6757 (N_6757,N_3580,N_3904);
or U6758 (N_6758,N_2162,N_3601);
nor U6759 (N_6759,N_3826,N_2899);
xor U6760 (N_6760,N_2943,N_1927);
xnor U6761 (N_6761,N_3080,N_3942);
or U6762 (N_6762,N_3142,N_922);
nor U6763 (N_6763,N_2806,N_3637);
nand U6764 (N_6764,N_2344,N_4116);
nand U6765 (N_6765,N_3323,N_3009);
nand U6766 (N_6766,N_2380,N_2753);
or U6767 (N_6767,N_783,N_2959);
nor U6768 (N_6768,N_2259,N_2687);
and U6769 (N_6769,N_4914,N_3794);
nand U6770 (N_6770,N_3319,N_4649);
and U6771 (N_6771,N_4769,N_2408);
and U6772 (N_6772,N_948,N_4541);
and U6773 (N_6773,N_1997,N_3736);
or U6774 (N_6774,N_4749,N_1347);
or U6775 (N_6775,N_2890,N_4365);
and U6776 (N_6776,N_3045,N_4977);
nand U6777 (N_6777,N_4280,N_829);
nor U6778 (N_6778,N_2129,N_2554);
xnor U6779 (N_6779,N_2810,N_212);
nor U6780 (N_6780,N_4110,N_4741);
or U6781 (N_6781,N_2794,N_2158);
xor U6782 (N_6782,N_4027,N_4492);
nor U6783 (N_6783,N_2530,N_1394);
nand U6784 (N_6784,N_2029,N_4479);
nand U6785 (N_6785,N_2117,N_2304);
nand U6786 (N_6786,N_203,N_2498);
nand U6787 (N_6787,N_1617,N_2834);
and U6788 (N_6788,N_4779,N_3564);
xnor U6789 (N_6789,N_300,N_2869);
and U6790 (N_6790,N_3156,N_1447);
or U6791 (N_6791,N_3014,N_3082);
nand U6792 (N_6792,N_421,N_2449);
or U6793 (N_6793,N_2690,N_1219);
nand U6794 (N_6794,N_1543,N_148);
xor U6795 (N_6795,N_858,N_1674);
nand U6796 (N_6796,N_3256,N_1908);
or U6797 (N_6797,N_1552,N_1031);
nor U6798 (N_6798,N_2328,N_3483);
and U6799 (N_6799,N_3324,N_2429);
and U6800 (N_6800,N_4353,N_1834);
or U6801 (N_6801,N_34,N_549);
nand U6802 (N_6802,N_2361,N_158);
or U6803 (N_6803,N_4990,N_803);
nor U6804 (N_6804,N_1242,N_1950);
nor U6805 (N_6805,N_4635,N_2669);
and U6806 (N_6806,N_2843,N_3250);
xor U6807 (N_6807,N_3201,N_874);
nand U6808 (N_6808,N_4724,N_1685);
and U6809 (N_6809,N_3555,N_4676);
and U6810 (N_6810,N_2109,N_2774);
or U6811 (N_6811,N_1971,N_4558);
and U6812 (N_6812,N_2748,N_1026);
or U6813 (N_6813,N_1121,N_2101);
nor U6814 (N_6814,N_3718,N_512);
xnor U6815 (N_6815,N_1527,N_2237);
xor U6816 (N_6816,N_3061,N_4098);
nor U6817 (N_6817,N_2355,N_1068);
and U6818 (N_6818,N_4500,N_1563);
xnor U6819 (N_6819,N_925,N_4234);
nor U6820 (N_6820,N_4091,N_4650);
xor U6821 (N_6821,N_3401,N_3174);
or U6822 (N_6822,N_1758,N_1750);
nand U6823 (N_6823,N_2492,N_2827);
or U6824 (N_6824,N_4689,N_1224);
and U6825 (N_6825,N_3631,N_1814);
nand U6826 (N_6826,N_3412,N_1038);
and U6827 (N_6827,N_4816,N_93);
or U6828 (N_6828,N_4835,N_1480);
or U6829 (N_6829,N_3011,N_3049);
xor U6830 (N_6830,N_457,N_4023);
and U6831 (N_6831,N_2250,N_1119);
or U6832 (N_6832,N_2760,N_3468);
and U6833 (N_6833,N_2470,N_2875);
or U6834 (N_6834,N_263,N_4679);
or U6835 (N_6835,N_4313,N_368);
nand U6836 (N_6836,N_2532,N_676);
nand U6837 (N_6837,N_121,N_277);
nand U6838 (N_6838,N_2624,N_3627);
and U6839 (N_6839,N_173,N_2511);
nand U6840 (N_6840,N_3290,N_2731);
xnor U6841 (N_6841,N_2767,N_4884);
or U6842 (N_6842,N_903,N_1711);
xnor U6843 (N_6843,N_1999,N_4224);
nand U6844 (N_6844,N_2773,N_3286);
nor U6845 (N_6845,N_4052,N_4863);
xnor U6846 (N_6846,N_839,N_4243);
xnor U6847 (N_6847,N_901,N_2353);
and U6848 (N_6848,N_2457,N_2066);
or U6849 (N_6849,N_3715,N_4536);
or U6850 (N_6850,N_3568,N_2320);
and U6851 (N_6851,N_1981,N_1246);
xor U6852 (N_6852,N_4905,N_1840);
xor U6853 (N_6853,N_1259,N_1488);
nor U6854 (N_6854,N_529,N_1763);
or U6855 (N_6855,N_1162,N_3251);
xor U6856 (N_6856,N_3536,N_2462);
nor U6857 (N_6857,N_4057,N_3727);
nor U6858 (N_6858,N_1202,N_3883);
nor U6859 (N_6859,N_1974,N_2650);
nor U6860 (N_6860,N_2698,N_1361);
or U6861 (N_6861,N_1104,N_3053);
and U6862 (N_6862,N_4912,N_4509);
xnor U6863 (N_6863,N_4982,N_154);
xor U6864 (N_6864,N_2142,N_969);
xnor U6865 (N_6865,N_3444,N_3662);
nor U6866 (N_6866,N_3033,N_3995);
xnor U6867 (N_6867,N_2597,N_2974);
nand U6868 (N_6868,N_741,N_3612);
xnor U6869 (N_6869,N_4105,N_1437);
xnor U6870 (N_6870,N_2070,N_1699);
or U6871 (N_6871,N_4709,N_749);
nand U6872 (N_6872,N_3997,N_3685);
xnor U6873 (N_6873,N_1788,N_85);
nand U6874 (N_6874,N_317,N_2342);
or U6875 (N_6875,N_3294,N_2634);
and U6876 (N_6876,N_582,N_3819);
nor U6877 (N_6877,N_2413,N_3928);
xor U6878 (N_6878,N_3949,N_4648);
nand U6879 (N_6879,N_4424,N_400);
or U6880 (N_6880,N_1145,N_404);
nor U6881 (N_6881,N_16,N_2871);
nor U6882 (N_6882,N_2340,N_4578);
nor U6883 (N_6883,N_4264,N_1212);
nand U6884 (N_6884,N_4127,N_152);
nand U6885 (N_6885,N_428,N_3870);
and U6886 (N_6886,N_2975,N_309);
or U6887 (N_6887,N_3175,N_1363);
nand U6888 (N_6888,N_3946,N_4580);
xnor U6889 (N_6889,N_4810,N_4173);
xor U6890 (N_6890,N_1897,N_3737);
nor U6891 (N_6891,N_2844,N_2401);
nor U6892 (N_6892,N_4610,N_651);
and U6893 (N_6893,N_4444,N_1432);
and U6894 (N_6894,N_1634,N_771);
and U6895 (N_6895,N_3886,N_2448);
nand U6896 (N_6896,N_2170,N_339);
and U6897 (N_6897,N_578,N_3349);
and U6898 (N_6898,N_2761,N_4806);
nor U6899 (N_6899,N_1196,N_3660);
and U6900 (N_6900,N_3159,N_575);
or U6901 (N_6901,N_3760,N_302);
nand U6902 (N_6902,N_838,N_836);
nor U6903 (N_6903,N_727,N_24);
and U6904 (N_6904,N_2518,N_2112);
and U6905 (N_6905,N_2723,N_1283);
or U6906 (N_6906,N_4738,N_3048);
and U6907 (N_6907,N_1111,N_2089);
nand U6908 (N_6908,N_637,N_3152);
or U6909 (N_6909,N_4031,N_1771);
and U6910 (N_6910,N_805,N_1583);
xor U6911 (N_6911,N_3598,N_4859);
nand U6912 (N_6912,N_3275,N_1237);
xor U6913 (N_6913,N_947,N_4751);
or U6914 (N_6914,N_3141,N_3103);
or U6915 (N_6915,N_2813,N_2936);
or U6916 (N_6916,N_486,N_3026);
nand U6917 (N_6917,N_3188,N_2832);
and U6918 (N_6918,N_900,N_924);
and U6919 (N_6919,N_3325,N_4223);
or U6920 (N_6920,N_751,N_4909);
nor U6921 (N_6921,N_3697,N_2569);
xor U6922 (N_6922,N_1291,N_429);
xnor U6923 (N_6923,N_2989,N_4571);
nor U6924 (N_6924,N_4786,N_2185);
and U6925 (N_6925,N_3522,N_2014);
and U6926 (N_6926,N_4898,N_3454);
xor U6927 (N_6927,N_1159,N_515);
and U6928 (N_6928,N_2681,N_2976);
nor U6929 (N_6929,N_4917,N_3492);
nand U6930 (N_6930,N_4544,N_2925);
nand U6931 (N_6931,N_3231,N_4055);
nand U6932 (N_6932,N_2169,N_202);
nand U6933 (N_6933,N_2563,N_3758);
and U6934 (N_6934,N_4131,N_2197);
or U6935 (N_6935,N_119,N_683);
nor U6936 (N_6936,N_841,N_1482);
nor U6937 (N_6937,N_4140,N_4945);
xor U6938 (N_6938,N_632,N_90);
nor U6939 (N_6939,N_3039,N_3689);
nor U6940 (N_6940,N_231,N_822);
or U6941 (N_6941,N_1445,N_960);
nor U6942 (N_6942,N_2326,N_3466);
xnor U6943 (N_6943,N_2131,N_748);
xnor U6944 (N_6944,N_2292,N_3282);
and U6945 (N_6945,N_2625,N_488);
nand U6946 (N_6946,N_2636,N_1821);
or U6947 (N_6947,N_3230,N_2446);
nor U6948 (N_6948,N_1369,N_37);
nand U6949 (N_6949,N_2570,N_4579);
or U6950 (N_6950,N_4046,N_2336);
xnor U6951 (N_6951,N_3748,N_1281);
or U6952 (N_6952,N_1444,N_2546);
xor U6953 (N_6953,N_4004,N_4908);
nand U6954 (N_6954,N_790,N_3283);
nand U6955 (N_6955,N_1004,N_387);
nand U6956 (N_6956,N_1459,N_1817);
and U6957 (N_6957,N_2245,N_2512);
xor U6958 (N_6958,N_1066,N_2849);
and U6959 (N_6959,N_1270,N_3041);
xnor U6960 (N_6960,N_4550,N_205);
nor U6961 (N_6961,N_4739,N_1247);
nor U6962 (N_6962,N_254,N_968);
or U6963 (N_6963,N_3844,N_953);
or U6964 (N_6964,N_369,N_1139);
xor U6965 (N_6965,N_1254,N_3147);
nand U6966 (N_6966,N_2654,N_4780);
and U6967 (N_6967,N_4158,N_3321);
xnor U6968 (N_6968,N_728,N_2127);
nor U6969 (N_6969,N_192,N_1576);
or U6970 (N_6970,N_450,N_4403);
and U6971 (N_6971,N_2992,N_4109);
and U6972 (N_6972,N_2839,N_1313);
and U6973 (N_6973,N_3461,N_3341);
nand U6974 (N_6974,N_3790,N_3059);
and U6975 (N_6975,N_2321,N_1565);
nand U6976 (N_6976,N_285,N_3711);
xnor U6977 (N_6977,N_3473,N_1070);
nand U6978 (N_6978,N_662,N_434);
and U6979 (N_6979,N_2166,N_4019);
xnor U6980 (N_6980,N_684,N_3520);
or U6981 (N_6981,N_1695,N_3917);
nor U6982 (N_6982,N_3493,N_4260);
nor U6983 (N_6983,N_940,N_3074);
nand U6984 (N_6984,N_678,N_1133);
nor U6985 (N_6985,N_1317,N_2053);
xor U6986 (N_6986,N_2499,N_3969);
nor U6987 (N_6987,N_3394,N_1199);
nand U6988 (N_6988,N_1956,N_1659);
xnor U6989 (N_6989,N_1178,N_3431);
xnor U6990 (N_6990,N_4181,N_2298);
nor U6991 (N_6991,N_1994,N_1346);
xnor U6992 (N_6992,N_2639,N_2632);
xor U6993 (N_6993,N_160,N_3912);
nor U6994 (N_6994,N_1509,N_1579);
nand U6995 (N_6995,N_2248,N_1832);
nand U6996 (N_6996,N_4892,N_4240);
nand U6997 (N_6997,N_1628,N_463);
or U6998 (N_6998,N_4586,N_4068);
and U6999 (N_6999,N_4717,N_2719);
nor U7000 (N_7000,N_484,N_4366);
nor U7001 (N_7001,N_527,N_4734);
nor U7002 (N_7002,N_2732,N_845);
xnor U7003 (N_7003,N_622,N_3302);
and U7004 (N_7004,N_303,N_166);
xor U7005 (N_7005,N_2919,N_3263);
nand U7006 (N_7006,N_1339,N_3657);
and U7007 (N_7007,N_3170,N_580);
nor U7008 (N_7008,N_4566,N_4851);
or U7009 (N_7009,N_1670,N_4543);
nor U7010 (N_7010,N_3596,N_7);
and U7011 (N_7011,N_2635,N_313);
xnor U7012 (N_7012,N_2217,N_2728);
or U7013 (N_7013,N_1472,N_4381);
xor U7014 (N_7014,N_560,N_3348);
nor U7015 (N_7015,N_1942,N_1336);
and U7016 (N_7016,N_3482,N_1490);
nor U7017 (N_7017,N_477,N_1530);
xor U7018 (N_7018,N_1630,N_2379);
nor U7019 (N_7019,N_4981,N_2779);
or U7020 (N_7020,N_3781,N_437);
and U7021 (N_7021,N_3922,N_432);
nor U7022 (N_7022,N_1095,N_2535);
or U7023 (N_7023,N_455,N_341);
nand U7024 (N_7024,N_4532,N_1797);
nand U7025 (N_7025,N_2558,N_4759);
nand U7026 (N_7026,N_3875,N_1079);
and U7027 (N_7027,N_2868,N_3770);
nand U7028 (N_7028,N_4050,N_3649);
xnor U7029 (N_7029,N_3288,N_918);
xor U7030 (N_7030,N_32,N_136);
nand U7031 (N_7031,N_3334,N_1730);
nor U7032 (N_7032,N_3365,N_2118);
and U7033 (N_7033,N_111,N_79);
xor U7034 (N_7034,N_2375,N_4178);
nor U7035 (N_7035,N_2609,N_241);
nand U7036 (N_7036,N_852,N_1677);
nor U7037 (N_7037,N_4191,N_67);
or U7038 (N_7038,N_3670,N_600);
nor U7039 (N_7039,N_820,N_4552);
nor U7040 (N_7040,N_257,N_3806);
xor U7041 (N_7041,N_1915,N_1566);
or U7042 (N_7042,N_4464,N_13);
nand U7043 (N_7043,N_56,N_4714);
nor U7044 (N_7044,N_255,N_3418);
xnor U7045 (N_7045,N_2102,N_909);
nand U7046 (N_7046,N_2764,N_4016);
xor U7047 (N_7047,N_4056,N_3488);
nor U7048 (N_7048,N_3866,N_1169);
nor U7049 (N_7049,N_1714,N_1698);
and U7050 (N_7050,N_3895,N_2279);
nand U7051 (N_7051,N_1523,N_3332);
or U7052 (N_7052,N_4513,N_4494);
and U7053 (N_7053,N_2243,N_1285);
and U7054 (N_7054,N_1132,N_3239);
nor U7055 (N_7055,N_3472,N_3422);
nor U7056 (N_7056,N_4497,N_1258);
or U7057 (N_7057,N_4819,N_2356);
or U7058 (N_7058,N_3366,N_1830);
or U7059 (N_7059,N_1010,N_3058);
nor U7060 (N_7060,N_2357,N_3929);
or U7061 (N_7061,N_3860,N_2425);
nor U7062 (N_7062,N_3707,N_1161);
and U7063 (N_7063,N_451,N_2956);
and U7064 (N_7064,N_1731,N_4248);
nor U7065 (N_7065,N_318,N_1438);
and U7066 (N_7066,N_2921,N_4708);
and U7067 (N_7067,N_1083,N_3938);
and U7068 (N_7068,N_4437,N_4744);
nor U7069 (N_7069,N_4695,N_3042);
nor U7070 (N_7070,N_4801,N_3603);
nand U7071 (N_7071,N_1353,N_982);
or U7072 (N_7072,N_1318,N_3509);
and U7073 (N_7073,N_3222,N_542);
nor U7074 (N_7074,N_284,N_4597);
nor U7075 (N_7075,N_2065,N_2822);
nor U7076 (N_7076,N_2299,N_1568);
and U7077 (N_7077,N_117,N_1030);
and U7078 (N_7078,N_3276,N_3106);
nor U7079 (N_7079,N_4482,N_3607);
and U7080 (N_7080,N_43,N_2282);
nor U7081 (N_7081,N_2564,N_4913);
nand U7082 (N_7082,N_3055,N_3000);
xor U7083 (N_7083,N_200,N_1448);
xnor U7084 (N_7084,N_4707,N_2667);
or U7085 (N_7085,N_80,N_1901);
nor U7086 (N_7086,N_793,N_4097);
or U7087 (N_7087,N_2465,N_916);
and U7088 (N_7088,N_2579,N_2969);
and U7089 (N_7089,N_4551,N_3452);
nor U7090 (N_7090,N_1515,N_1072);
nor U7091 (N_7091,N_422,N_2565);
nor U7092 (N_7092,N_3531,N_1266);
xor U7093 (N_7093,N_4994,N_2928);
or U7094 (N_7094,N_227,N_2364);
xor U7095 (N_7095,N_2926,N_371);
xnor U7096 (N_7096,N_1456,N_94);
nand U7097 (N_7097,N_1524,N_4122);
or U7098 (N_7098,N_4006,N_1239);
or U7099 (N_7099,N_4184,N_2366);
or U7100 (N_7100,N_1818,N_4647);
xnor U7101 (N_7101,N_3985,N_3793);
or U7102 (N_7102,N_2191,N_1781);
and U7103 (N_7103,N_3754,N_2556);
and U7104 (N_7104,N_1359,N_887);
or U7105 (N_7105,N_3186,N_2781);
and U7106 (N_7106,N_1591,N_4389);
nand U7107 (N_7107,N_3958,N_38);
or U7108 (N_7108,N_1643,N_3204);
or U7109 (N_7109,N_2313,N_4715);
or U7110 (N_7110,N_3782,N_1764);
nor U7111 (N_7111,N_4443,N_104);
nor U7112 (N_7112,N_1640,N_1256);
xor U7113 (N_7113,N_1328,N_2500);
nor U7114 (N_7114,N_2829,N_4796);
and U7115 (N_7115,N_2514,N_105);
or U7116 (N_7116,N_2335,N_514);
nand U7117 (N_7117,N_2642,N_2405);
or U7118 (N_7118,N_3138,N_481);
nand U7119 (N_7119,N_4453,N_3888);
xnor U7120 (N_7120,N_3322,N_4129);
nor U7121 (N_7121,N_2145,N_4701);
or U7122 (N_7122,N_4789,N_1294);
nor U7123 (N_7123,N_4294,N_3842);
and U7124 (N_7124,N_1471,N_259);
or U7125 (N_7125,N_4451,N_4839);
or U7126 (N_7126,N_1850,N_1406);
nor U7127 (N_7127,N_2724,N_4051);
nand U7128 (N_7128,N_1747,N_4220);
nor U7129 (N_7129,N_1776,N_3623);
xor U7130 (N_7130,N_3133,N_4048);
nor U7131 (N_7131,N_2149,N_4418);
xnor U7132 (N_7132,N_1023,N_1753);
nor U7133 (N_7133,N_3732,N_3419);
nor U7134 (N_7134,N_4970,N_4967);
nor U7135 (N_7135,N_4462,N_4760);
and U7136 (N_7136,N_4009,N_3362);
xnor U7137 (N_7137,N_4662,N_1059);
nand U7138 (N_7138,N_4907,N_4213);
nor U7139 (N_7139,N_699,N_4336);
nand U7140 (N_7140,N_1021,N_4011);
nor U7141 (N_7141,N_4765,N_724);
or U7142 (N_7142,N_3776,N_3981);
nand U7143 (N_7143,N_1589,N_394);
or U7144 (N_7144,N_3499,N_1704);
nor U7145 (N_7145,N_552,N_475);
and U7146 (N_7146,N_819,N_3337);
nor U7147 (N_7147,N_1307,N_1545);
nand U7148 (N_7148,N_3430,N_4447);
nor U7149 (N_7149,N_2596,N_3358);
or U7150 (N_7150,N_4615,N_2856);
nand U7151 (N_7151,N_3813,N_4611);
nor U7152 (N_7152,N_3622,N_1343);
or U7153 (N_7153,N_3699,N_2048);
and U7154 (N_7154,N_4725,N_2168);
and U7155 (N_7155,N_3240,N_4713);
xnor U7156 (N_7156,N_1933,N_928);
xnor U7157 (N_7157,N_3693,N_1016);
xor U7158 (N_7158,N_2246,N_2090);
xor U7159 (N_7159,N_840,N_1871);
nand U7160 (N_7160,N_3167,N_541);
nor U7161 (N_7161,N_1910,N_2205);
nand U7162 (N_7162,N_3823,N_1946);
xnor U7163 (N_7163,N_949,N_3996);
or U7164 (N_7164,N_76,N_3966);
nand U7165 (N_7165,N_4825,N_3869);
nand U7166 (N_7166,N_1724,N_4172);
or U7167 (N_7167,N_1310,N_4135);
nor U7168 (N_7168,N_2589,N_1113);
and U7169 (N_7169,N_470,N_2367);
and U7170 (N_7170,N_2984,N_4305);
xor U7171 (N_7171,N_1100,N_2496);
or U7172 (N_7172,N_4472,N_288);
nor U7173 (N_7173,N_1227,N_1742);
nor U7174 (N_7174,N_113,N_439);
nor U7175 (N_7175,N_2520,N_2861);
nand U7176 (N_7176,N_985,N_1863);
and U7177 (N_7177,N_4678,N_4657);
and U7178 (N_7178,N_1091,N_327);
nor U7179 (N_7179,N_2600,N_1466);
and U7180 (N_7180,N_1717,N_4747);
and U7181 (N_7181,N_1057,N_2575);
nor U7182 (N_7182,N_653,N_716);
and U7183 (N_7183,N_1809,N_2333);
and U7184 (N_7184,N_3245,N_1646);
or U7185 (N_7185,N_221,N_3960);
nor U7186 (N_7186,N_2254,N_4978);
xnor U7187 (N_7187,N_553,N_4355);
nor U7188 (N_7188,N_2267,N_3885);
and U7189 (N_7189,N_2973,N_3343);
and U7190 (N_7190,N_2210,N_665);
xnor U7191 (N_7191,N_4456,N_2734);
xor U7192 (N_7192,N_1223,N_2675);
and U7193 (N_7193,N_4039,N_4330);
or U7194 (N_7194,N_1262,N_2451);
or U7195 (N_7195,N_3117,N_2735);
xnor U7196 (N_7196,N_116,N_4946);
nor U7197 (N_7197,N_4654,N_2885);
xor U7198 (N_7198,N_3339,N_4370);
nor U7199 (N_7199,N_4210,N_1422);
and U7200 (N_7200,N_2901,N_2851);
nand U7201 (N_7201,N_4035,N_4904);
nand U7202 (N_7202,N_747,N_2701);
or U7203 (N_7203,N_1450,N_883);
and U7204 (N_7204,N_3858,N_3089);
nor U7205 (N_7205,N_2935,N_3787);
or U7206 (N_7206,N_2703,N_4842);
nand U7207 (N_7207,N_295,N_4461);
xor U7208 (N_7208,N_1590,N_4720);
or U7209 (N_7209,N_2580,N_1691);
xnor U7210 (N_7210,N_2692,N_547);
nor U7211 (N_7211,N_3798,N_1916);
nand U7212 (N_7212,N_500,N_4925);
xnor U7213 (N_7213,N_1112,N_2160);
nor U7214 (N_7214,N_4463,N_4652);
or U7215 (N_7215,N_812,N_4685);
xor U7216 (N_7216,N_1705,N_1141);
xnor U7217 (N_7217,N_266,N_1379);
xnor U7218 (N_7218,N_603,N_1988);
xnor U7219 (N_7219,N_2086,N_2630);
nor U7220 (N_7220,N_669,N_367);
xnor U7221 (N_7221,N_3202,N_768);
nand U7222 (N_7222,N_4545,N_3278);
nand U7223 (N_7223,N_3247,N_1292);
nand U7224 (N_7224,N_3510,N_3642);
nor U7225 (N_7225,N_703,N_4145);
nand U7226 (N_7226,N_407,N_4174);
nand U7227 (N_7227,N_2607,N_693);
nand U7228 (N_7228,N_1931,N_3558);
nor U7229 (N_7229,N_4060,N_608);
xnor U7230 (N_7230,N_1554,N_201);
nor U7231 (N_7231,N_4542,N_4998);
nor U7232 (N_7232,N_1129,N_4607);
and U7233 (N_7233,N_785,N_4915);
or U7234 (N_7234,N_4963,N_3423);
nand U7235 (N_7235,N_4687,N_3105);
and U7236 (N_7236,N_824,N_2293);
nand U7237 (N_7237,N_912,N_633);
or U7238 (N_7238,N_3378,N_1331);
nand U7239 (N_7239,N_4038,N_869);
nand U7240 (N_7240,N_2879,N_352);
and U7241 (N_7241,N_4147,N_3137);
nor U7242 (N_7242,N_2155,N_215);
and U7243 (N_7243,N_2857,N_4222);
nor U7244 (N_7244,N_4291,N_945);
nor U7245 (N_7245,N_3291,N_3664);
xor U7246 (N_7246,N_1542,N_862);
nor U7247 (N_7247,N_4143,N_3578);
and U7248 (N_7248,N_2475,N_4797);
and U7249 (N_7249,N_4177,N_4318);
nor U7250 (N_7250,N_122,N_4120);
nor U7251 (N_7251,N_1424,N_3626);
and U7252 (N_7252,N_3721,N_2970);
or U7253 (N_7253,N_3097,N_1267);
or U7254 (N_7254,N_815,N_702);
and U7255 (N_7255,N_4533,N_364);
and U7256 (N_7256,N_31,N_3114);
or U7257 (N_7257,N_2840,N_4893);
and U7258 (N_7258,N_3992,N_1177);
xnor U7259 (N_7259,N_4150,N_2562);
or U7260 (N_7260,N_478,N_2215);
or U7261 (N_7261,N_1053,N_886);
nor U7262 (N_7262,N_1249,N_3036);
and U7263 (N_7263,N_4682,N_3101);
nand U7264 (N_7264,N_813,N_3890);
and U7265 (N_7265,N_3887,N_2713);
nand U7266 (N_7266,N_306,N_4286);
nor U7267 (N_7267,N_269,N_193);
or U7268 (N_7268,N_3044,N_4871);
xnor U7269 (N_7269,N_3279,N_3979);
and U7270 (N_7270,N_2097,N_1709);
nand U7271 (N_7271,N_4086,N_3615);
nand U7272 (N_7272,N_2309,N_1798);
and U7273 (N_7273,N_2285,N_3062);
and U7274 (N_7274,N_1859,N_4811);
nor U7275 (N_7275,N_2738,N_626);
or U7276 (N_7276,N_4111,N_2507);
nor U7277 (N_7277,N_4160,N_1923);
or U7278 (N_7278,N_2573,N_3335);
nor U7279 (N_7279,N_4594,N_1304);
nand U7280 (N_7280,N_4790,N_149);
nor U7281 (N_7281,N_2471,N_2022);
xor U7282 (N_7282,N_107,N_2981);
xor U7283 (N_7283,N_4847,N_3116);
nor U7284 (N_7284,N_3470,N_1739);
and U7285 (N_7285,N_4276,N_1198);
nor U7286 (N_7286,N_565,N_4476);
and U7287 (N_7287,N_1559,N_1865);
nand U7288 (N_7288,N_1842,N_3991);
nand U7289 (N_7289,N_1275,N_718);
xor U7290 (N_7290,N_4596,N_2955);
nand U7291 (N_7291,N_1744,N_1914);
or U7292 (N_7292,N_2193,N_3109);
nor U7293 (N_7293,N_730,N_1420);
nand U7294 (N_7294,N_3284,N_1229);
nand U7295 (N_7295,N_1868,N_706);
nand U7296 (N_7296,N_3373,N_3124);
xnor U7297 (N_7297,N_4852,N_2646);
xor U7298 (N_7298,N_873,N_3308);
and U7299 (N_7299,N_3262,N_955);
xor U7300 (N_7300,N_3360,N_403);
xor U7301 (N_7301,N_4307,N_4274);
nand U7302 (N_7302,N_2725,N_4653);
xor U7303 (N_7303,N_3208,N_1625);
nand U7304 (N_7304,N_1631,N_3914);
nor U7305 (N_7305,N_4837,N_4997);
or U7306 (N_7306,N_3005,N_2870);
nor U7307 (N_7307,N_1825,N_3865);
nand U7308 (N_7308,N_1467,N_3600);
or U7309 (N_7309,N_3713,N_856);
and U7310 (N_7310,N_826,N_4920);
nand U7311 (N_7311,N_1392,N_3588);
or U7312 (N_7312,N_1387,N_686);
and U7313 (N_7313,N_2603,N_1681);
nor U7314 (N_7314,N_1497,N_1884);
and U7315 (N_7315,N_1149,N_3965);
nand U7316 (N_7316,N_4254,N_4957);
nand U7317 (N_7317,N_2680,N_95);
xor U7318 (N_7318,N_3237,N_2488);
nand U7319 (N_7319,N_2846,N_2176);
or U7320 (N_7320,N_1799,N_1398);
nand U7321 (N_7321,N_2858,N_4423);
nor U7322 (N_7322,N_1836,N_2862);
or U7323 (N_7323,N_657,N_3066);
or U7324 (N_7324,N_911,N_2202);
nand U7325 (N_7325,N_1562,N_1173);
and U7326 (N_7326,N_1449,N_4082);
or U7327 (N_7327,N_3774,N_4103);
xnor U7328 (N_7328,N_4377,N_4936);
nor U7329 (N_7329,N_2000,N_3827);
and U7330 (N_7330,N_3772,N_2028);
and U7331 (N_7331,N_3686,N_1796);
xor U7332 (N_7332,N_256,N_1673);
or U7333 (N_7333,N_3487,N_2918);
nor U7334 (N_7334,N_1280,N_2384);
and U7335 (N_7335,N_2991,N_2929);
nand U7336 (N_7336,N_441,N_3537);
or U7337 (N_7337,N_1756,N_1726);
or U7338 (N_7338,N_4071,N_129);
or U7339 (N_7339,N_3593,N_4261);
and U7340 (N_7340,N_2124,N_260);
or U7341 (N_7341,N_4740,N_1263);
nand U7342 (N_7342,N_752,N_3441);
and U7343 (N_7343,N_3345,N_1011);
xor U7344 (N_7344,N_3149,N_2770);
or U7345 (N_7345,N_2186,N_3404);
and U7346 (N_7346,N_376,N_4176);
xor U7347 (N_7347,N_1540,N_4929);
nand U7348 (N_7348,N_1460,N_316);
and U7349 (N_7349,N_4832,N_4349);
and U7350 (N_7350,N_3893,N_3128);
and U7351 (N_7351,N_566,N_2173);
nand U7352 (N_7352,N_3775,N_3814);
and U7353 (N_7353,N_4548,N_3871);
and U7354 (N_7354,N_1170,N_1947);
xnor U7355 (N_7355,N_2373,N_386);
nand U7356 (N_7356,N_482,N_1452);
xnor U7357 (N_7357,N_3024,N_2194);
nor U7358 (N_7358,N_293,N_4167);
and U7359 (N_7359,N_4969,N_351);
xnor U7360 (N_7360,N_3351,N_1828);
or U7361 (N_7361,N_4809,N_2306);
and U7362 (N_7362,N_690,N_544);
nand U7363 (N_7363,N_3185,N_4560);
nand U7364 (N_7364,N_2907,N_3582);
nor U7365 (N_7365,N_1725,N_2414);
and U7366 (N_7366,N_1182,N_3043);
nand U7367 (N_7367,N_4391,N_1976);
nand U7368 (N_7368,N_1050,N_4380);
nor U7369 (N_7369,N_4980,N_1027);
xnor U7370 (N_7370,N_1278,N_3119);
nand U7371 (N_7371,N_694,N_808);
or U7372 (N_7372,N_3190,N_756);
and U7373 (N_7373,N_1881,N_297);
nor U7374 (N_7374,N_2721,N_1569);
nor U7375 (N_7375,N_3436,N_2297);
or U7376 (N_7376,N_29,N_1128);
or U7377 (N_7377,N_15,N_2431);
and U7378 (N_7378,N_2765,N_1736);
xor U7379 (N_7379,N_1184,N_4564);
xor U7380 (N_7380,N_4638,N_4346);
nand U7381 (N_7381,N_3516,N_1412);
nand U7382 (N_7382,N_602,N_3301);
and U7383 (N_7383,N_4282,N_319);
and U7384 (N_7384,N_2946,N_1305);
or U7385 (N_7385,N_4672,N_670);
xor U7386 (N_7386,N_4197,N_2263);
or U7387 (N_7387,N_1765,N_1525);
and U7388 (N_7388,N_3007,N_2466);
nor U7389 (N_7389,N_557,N_4439);
and U7390 (N_7390,N_988,N_4931);
and U7391 (N_7391,N_2213,N_2659);
nor U7392 (N_7392,N_4699,N_445);
nor U7393 (N_7393,N_1086,N_2631);
or U7394 (N_7394,N_964,N_108);
nor U7395 (N_7395,N_2412,N_1036);
or U7396 (N_7396,N_2345,N_1408);
or U7397 (N_7397,N_4766,N_3165);
and U7398 (N_7398,N_55,N_1718);
xnor U7399 (N_7399,N_1738,N_2113);
xnor U7400 (N_7400,N_3125,N_3976);
or U7401 (N_7401,N_1860,N_801);
nor U7402 (N_7402,N_1891,N_4733);
xor U7403 (N_7403,N_3983,N_1503);
or U7404 (N_7404,N_1024,N_1573);
or U7405 (N_7405,N_4397,N_2126);
nor U7406 (N_7406,N_3587,N_2139);
and U7407 (N_7407,N_4457,N_2040);
and U7408 (N_7408,N_4506,N_2508);
nand U7409 (N_7409,N_4299,N_1597);
nor U7410 (N_7410,N_4405,N_2583);
nor U7411 (N_7411,N_1604,N_4686);
xor U7412 (N_7412,N_1434,N_850);
and U7413 (N_7413,N_735,N_4748);
nor U7414 (N_7414,N_4841,N_4413);
or U7415 (N_7415,N_902,N_2783);
xor U7416 (N_7416,N_2424,N_3392);
xnor U7417 (N_7417,N_4265,N_2930);
nand U7418 (N_7418,N_268,N_3399);
nand U7419 (N_7419,N_1419,N_941);
nand U7420 (N_7420,N_3855,N_1217);
or U7421 (N_7421,N_581,N_373);
or U7422 (N_7422,N_2482,N_1632);
xor U7423 (N_7423,N_3800,N_472);
xor U7424 (N_7424,N_823,N_583);
nand U7425 (N_7425,N_2780,N_4328);
nand U7426 (N_7426,N_666,N_4332);
and U7427 (N_7427,N_2349,N_2852);
and U7428 (N_7428,N_3982,N_3641);
nor U7429 (N_7429,N_2080,N_917);
nor U7430 (N_7430,N_2181,N_2957);
or U7431 (N_7431,N_4021,N_2528);
nor U7432 (N_7432,N_4468,N_401);
nand U7433 (N_7433,N_3193,N_2330);
nand U7434 (N_7434,N_1326,N_1252);
or U7435 (N_7435,N_1638,N_3896);
or U7436 (N_7436,N_1772,N_1804);
or U7437 (N_7437,N_4059,N_4138);
nor U7438 (N_7438,N_3619,N_3948);
xor U7439 (N_7439,N_2828,N_4755);
xor U7440 (N_7440,N_4348,N_4632);
nor U7441 (N_7441,N_2715,N_4368);
or U7442 (N_7442,N_3395,N_1152);
and U7443 (N_7443,N_4376,N_4664);
xor U7444 (N_7444,N_4572,N_593);
xnor U7445 (N_7445,N_1858,N_3272);
nor U7446 (N_7446,N_1105,N_1682);
and U7447 (N_7447,N_2604,N_3361);
and U7448 (N_7448,N_3189,N_2450);
nand U7449 (N_7449,N_4092,N_3206);
and U7450 (N_7450,N_3762,N_4783);
nand U7451 (N_7451,N_444,N_4659);
nor U7452 (N_7452,N_2536,N_4253);
xor U7453 (N_7453,N_283,N_4314);
and U7454 (N_7454,N_4404,N_3513);
nor U7455 (N_7455,N_2421,N_101);
and U7456 (N_7456,N_1985,N_1282);
nor U7457 (N_7457,N_3453,N_4501);
xor U7458 (N_7458,N_178,N_611);
and U7459 (N_7459,N_1737,N_2325);
and U7460 (N_7460,N_2516,N_1669);
and U7461 (N_7461,N_2606,N_1824);
xnor U7462 (N_7462,N_4826,N_4356);
nand U7463 (N_7463,N_2314,N_1019);
and U7464 (N_7464,N_156,N_3087);
nand U7465 (N_7465,N_1959,N_2473);
and U7466 (N_7466,N_733,N_1585);
nor U7467 (N_7467,N_4096,N_1920);
and U7468 (N_7468,N_3207,N_1864);
xnor U7469 (N_7469,N_408,N_4383);
or U7470 (N_7470,N_4102,N_4088);
or U7471 (N_7471,N_4112,N_846);
xor U7472 (N_7472,N_4347,N_1575);
nor U7473 (N_7473,N_3350,N_1271);
nand U7474 (N_7474,N_3735,N_2433);
or U7475 (N_7475,N_3040,N_4215);
xor U7476 (N_7476,N_485,N_2653);
nand U7477 (N_7477,N_1512,N_2598);
nand U7478 (N_7478,N_1887,N_2793);
nor U7479 (N_7479,N_2716,N_4386);
nand U7480 (N_7480,N_994,N_357);
nor U7481 (N_7481,N_4601,N_861);
xnor U7482 (N_7482,N_546,N_2219);
nor U7483 (N_7483,N_738,N_1485);
and U7484 (N_7484,N_1373,N_2442);
nor U7485 (N_7485,N_959,N_2371);
nor U7486 (N_7486,N_943,N_64);
nand U7487 (N_7487,N_3918,N_1723);
nor U7488 (N_7488,N_2354,N_1124);
nand U7489 (N_7489,N_1816,N_1365);
nor U7490 (N_7490,N_1367,N_3445);
nand U7491 (N_7491,N_3744,N_365);
and U7492 (N_7492,N_1330,N_3511);
nor U7493 (N_7493,N_1768,N_3632);
nand U7494 (N_7494,N_3690,N_4675);
or U7495 (N_7495,N_4106,N_630);
and U7496 (N_7496,N_4132,N_1727);
nand U7497 (N_7497,N_1032,N_1077);
nor U7498 (N_7498,N_1203,N_3539);
xor U7499 (N_7499,N_194,N_3196);
nor U7500 (N_7500,N_4064,N_692);
nand U7501 (N_7501,N_121,N_2294);
and U7502 (N_7502,N_1704,N_1906);
xor U7503 (N_7503,N_2454,N_3325);
nor U7504 (N_7504,N_3785,N_943);
and U7505 (N_7505,N_4923,N_4339);
or U7506 (N_7506,N_1067,N_3873);
and U7507 (N_7507,N_97,N_4338);
or U7508 (N_7508,N_2615,N_2481);
nand U7509 (N_7509,N_428,N_2747);
nor U7510 (N_7510,N_2992,N_4360);
or U7511 (N_7511,N_3945,N_3144);
and U7512 (N_7512,N_4198,N_3413);
or U7513 (N_7513,N_2514,N_4206);
nor U7514 (N_7514,N_3534,N_3731);
and U7515 (N_7515,N_4905,N_2218);
nand U7516 (N_7516,N_2200,N_2574);
nor U7517 (N_7517,N_850,N_513);
xnor U7518 (N_7518,N_887,N_4134);
nor U7519 (N_7519,N_3778,N_1151);
and U7520 (N_7520,N_2241,N_2420);
xnor U7521 (N_7521,N_20,N_2315);
xor U7522 (N_7522,N_215,N_1643);
or U7523 (N_7523,N_34,N_2395);
xor U7524 (N_7524,N_1977,N_2092);
and U7525 (N_7525,N_598,N_2343);
nand U7526 (N_7526,N_3302,N_2151);
or U7527 (N_7527,N_4710,N_1763);
and U7528 (N_7528,N_3683,N_398);
xnor U7529 (N_7529,N_777,N_535);
and U7530 (N_7530,N_1697,N_3723);
xor U7531 (N_7531,N_1729,N_301);
and U7532 (N_7532,N_2070,N_4453);
and U7533 (N_7533,N_3829,N_4967);
nand U7534 (N_7534,N_873,N_1876);
xnor U7535 (N_7535,N_1734,N_2039);
and U7536 (N_7536,N_3673,N_100);
xor U7537 (N_7537,N_489,N_1076);
and U7538 (N_7538,N_1833,N_3218);
nor U7539 (N_7539,N_1363,N_904);
and U7540 (N_7540,N_3345,N_1182);
nor U7541 (N_7541,N_1965,N_212);
and U7542 (N_7542,N_1538,N_3763);
xor U7543 (N_7543,N_3003,N_3619);
and U7544 (N_7544,N_4939,N_2605);
xnor U7545 (N_7545,N_2365,N_385);
xnor U7546 (N_7546,N_1059,N_2904);
xor U7547 (N_7547,N_1242,N_2443);
or U7548 (N_7548,N_4015,N_4121);
or U7549 (N_7549,N_262,N_1793);
xnor U7550 (N_7550,N_4835,N_3751);
xnor U7551 (N_7551,N_947,N_438);
nand U7552 (N_7552,N_1878,N_3735);
nor U7553 (N_7553,N_147,N_2032);
nand U7554 (N_7554,N_3082,N_759);
and U7555 (N_7555,N_1724,N_1841);
xnor U7556 (N_7556,N_3808,N_3555);
nor U7557 (N_7557,N_783,N_4184);
and U7558 (N_7558,N_3118,N_2315);
xnor U7559 (N_7559,N_248,N_1502);
nor U7560 (N_7560,N_2304,N_2354);
nor U7561 (N_7561,N_1396,N_4468);
xnor U7562 (N_7562,N_223,N_1692);
and U7563 (N_7563,N_3406,N_2554);
xor U7564 (N_7564,N_3688,N_2507);
xor U7565 (N_7565,N_3368,N_1154);
xor U7566 (N_7566,N_4694,N_2290);
nor U7567 (N_7567,N_1067,N_1573);
and U7568 (N_7568,N_418,N_277);
and U7569 (N_7569,N_3184,N_3988);
or U7570 (N_7570,N_3171,N_3473);
or U7571 (N_7571,N_1422,N_2135);
and U7572 (N_7572,N_2416,N_1936);
nor U7573 (N_7573,N_800,N_3321);
xor U7574 (N_7574,N_3701,N_3988);
nor U7575 (N_7575,N_4317,N_2699);
and U7576 (N_7576,N_4767,N_1044);
or U7577 (N_7577,N_2755,N_1367);
and U7578 (N_7578,N_4887,N_51);
xnor U7579 (N_7579,N_661,N_3759);
and U7580 (N_7580,N_2100,N_1287);
nor U7581 (N_7581,N_4799,N_146);
nand U7582 (N_7582,N_3526,N_4426);
nor U7583 (N_7583,N_3305,N_3215);
and U7584 (N_7584,N_2603,N_2550);
or U7585 (N_7585,N_3598,N_1191);
and U7586 (N_7586,N_2882,N_2734);
or U7587 (N_7587,N_4240,N_1184);
or U7588 (N_7588,N_2716,N_4356);
or U7589 (N_7589,N_10,N_4999);
nand U7590 (N_7590,N_650,N_2094);
or U7591 (N_7591,N_2822,N_1021);
or U7592 (N_7592,N_2101,N_344);
nand U7593 (N_7593,N_3855,N_506);
or U7594 (N_7594,N_4108,N_2128);
nor U7595 (N_7595,N_3860,N_4306);
nor U7596 (N_7596,N_1102,N_4391);
xnor U7597 (N_7597,N_1813,N_1691);
or U7598 (N_7598,N_3561,N_907);
nor U7599 (N_7599,N_1775,N_3384);
nand U7600 (N_7600,N_244,N_2928);
and U7601 (N_7601,N_3238,N_2230);
and U7602 (N_7602,N_3321,N_3677);
or U7603 (N_7603,N_100,N_2439);
xor U7604 (N_7604,N_4455,N_2125);
or U7605 (N_7605,N_2967,N_193);
and U7606 (N_7606,N_4650,N_3315);
nand U7607 (N_7607,N_878,N_1750);
nand U7608 (N_7608,N_1900,N_1553);
and U7609 (N_7609,N_183,N_2591);
nand U7610 (N_7610,N_3072,N_3488);
nand U7611 (N_7611,N_1543,N_1857);
xnor U7612 (N_7612,N_3353,N_2575);
or U7613 (N_7613,N_1720,N_2572);
or U7614 (N_7614,N_1888,N_4210);
nor U7615 (N_7615,N_1187,N_618);
nand U7616 (N_7616,N_1727,N_4734);
nor U7617 (N_7617,N_1867,N_2845);
nor U7618 (N_7618,N_4164,N_3993);
or U7619 (N_7619,N_320,N_2980);
and U7620 (N_7620,N_4777,N_1680);
nand U7621 (N_7621,N_696,N_1597);
or U7622 (N_7622,N_4579,N_943);
or U7623 (N_7623,N_1719,N_530);
and U7624 (N_7624,N_2932,N_1362);
and U7625 (N_7625,N_3109,N_688);
or U7626 (N_7626,N_4417,N_3649);
or U7627 (N_7627,N_4785,N_2112);
or U7628 (N_7628,N_192,N_4985);
and U7629 (N_7629,N_118,N_1426);
xor U7630 (N_7630,N_3163,N_2017);
nor U7631 (N_7631,N_3569,N_926);
xor U7632 (N_7632,N_2879,N_2133);
nor U7633 (N_7633,N_3062,N_4047);
nor U7634 (N_7634,N_3682,N_64);
and U7635 (N_7635,N_4550,N_1680);
nor U7636 (N_7636,N_3682,N_102);
nand U7637 (N_7637,N_625,N_3673);
nor U7638 (N_7638,N_3775,N_1117);
xor U7639 (N_7639,N_426,N_3513);
nand U7640 (N_7640,N_3081,N_878);
nand U7641 (N_7641,N_3613,N_717);
xnor U7642 (N_7642,N_1336,N_3926);
and U7643 (N_7643,N_1279,N_1162);
or U7644 (N_7644,N_390,N_1200);
or U7645 (N_7645,N_2798,N_4683);
and U7646 (N_7646,N_3994,N_1984);
nand U7647 (N_7647,N_3802,N_1844);
and U7648 (N_7648,N_1839,N_4923);
xnor U7649 (N_7649,N_1157,N_1330);
or U7650 (N_7650,N_1315,N_2282);
nor U7651 (N_7651,N_843,N_3518);
or U7652 (N_7652,N_2028,N_4155);
xnor U7653 (N_7653,N_4348,N_1979);
xor U7654 (N_7654,N_2721,N_2773);
nand U7655 (N_7655,N_1904,N_1880);
and U7656 (N_7656,N_3524,N_1481);
xor U7657 (N_7657,N_4654,N_3872);
xnor U7658 (N_7658,N_1932,N_1564);
and U7659 (N_7659,N_1919,N_2266);
nor U7660 (N_7660,N_1178,N_1858);
and U7661 (N_7661,N_1530,N_2443);
xor U7662 (N_7662,N_396,N_55);
or U7663 (N_7663,N_990,N_1515);
xnor U7664 (N_7664,N_3971,N_2249);
and U7665 (N_7665,N_3797,N_3857);
xor U7666 (N_7666,N_1794,N_3710);
nand U7667 (N_7667,N_1008,N_508);
nor U7668 (N_7668,N_3236,N_3091);
nand U7669 (N_7669,N_4204,N_369);
nor U7670 (N_7670,N_2797,N_4025);
nand U7671 (N_7671,N_1285,N_306);
nand U7672 (N_7672,N_4995,N_970);
xor U7673 (N_7673,N_1399,N_4052);
nor U7674 (N_7674,N_1224,N_3994);
and U7675 (N_7675,N_1427,N_1850);
nor U7676 (N_7676,N_4206,N_1689);
nand U7677 (N_7677,N_1908,N_1236);
xor U7678 (N_7678,N_1282,N_3361);
nand U7679 (N_7679,N_4302,N_2666);
xnor U7680 (N_7680,N_1809,N_647);
or U7681 (N_7681,N_1253,N_2906);
xor U7682 (N_7682,N_4466,N_1780);
nor U7683 (N_7683,N_3902,N_3611);
nor U7684 (N_7684,N_3095,N_1546);
nor U7685 (N_7685,N_4457,N_4916);
or U7686 (N_7686,N_3345,N_527);
nand U7687 (N_7687,N_3381,N_766);
nand U7688 (N_7688,N_1268,N_3589);
nor U7689 (N_7689,N_2487,N_3230);
nand U7690 (N_7690,N_1728,N_558);
nand U7691 (N_7691,N_3675,N_2598);
nand U7692 (N_7692,N_4084,N_3710);
nand U7693 (N_7693,N_2753,N_1261);
nor U7694 (N_7694,N_4364,N_3127);
nand U7695 (N_7695,N_4197,N_1541);
nand U7696 (N_7696,N_3794,N_3427);
nor U7697 (N_7697,N_228,N_1460);
nor U7698 (N_7698,N_4184,N_1919);
and U7699 (N_7699,N_4918,N_3401);
nand U7700 (N_7700,N_4102,N_935);
nor U7701 (N_7701,N_2553,N_2247);
xor U7702 (N_7702,N_2421,N_3923);
xnor U7703 (N_7703,N_4851,N_2375);
or U7704 (N_7704,N_3950,N_1090);
or U7705 (N_7705,N_3111,N_2442);
or U7706 (N_7706,N_4031,N_1608);
nor U7707 (N_7707,N_4812,N_2862);
xor U7708 (N_7708,N_4853,N_1374);
xor U7709 (N_7709,N_3031,N_53);
or U7710 (N_7710,N_4044,N_392);
nand U7711 (N_7711,N_4650,N_4615);
and U7712 (N_7712,N_4851,N_1471);
nand U7713 (N_7713,N_1782,N_138);
xor U7714 (N_7714,N_4136,N_3121);
xnor U7715 (N_7715,N_3587,N_1389);
xor U7716 (N_7716,N_1027,N_3224);
or U7717 (N_7717,N_2703,N_2013);
nor U7718 (N_7718,N_4740,N_1628);
nand U7719 (N_7719,N_3730,N_3988);
and U7720 (N_7720,N_1967,N_160);
nor U7721 (N_7721,N_1023,N_4428);
nand U7722 (N_7722,N_1406,N_4139);
xor U7723 (N_7723,N_2653,N_4699);
and U7724 (N_7724,N_3406,N_23);
xor U7725 (N_7725,N_2379,N_4676);
and U7726 (N_7726,N_3672,N_1223);
and U7727 (N_7727,N_3529,N_2548);
nor U7728 (N_7728,N_923,N_2204);
nand U7729 (N_7729,N_1716,N_1025);
and U7730 (N_7730,N_4383,N_3765);
and U7731 (N_7731,N_2507,N_120);
or U7732 (N_7732,N_4012,N_4688);
or U7733 (N_7733,N_4127,N_3038);
and U7734 (N_7734,N_2626,N_3213);
nand U7735 (N_7735,N_4592,N_722);
and U7736 (N_7736,N_4804,N_1133);
xor U7737 (N_7737,N_2677,N_1669);
xnor U7738 (N_7738,N_4670,N_817);
xor U7739 (N_7739,N_969,N_4857);
and U7740 (N_7740,N_1099,N_1182);
or U7741 (N_7741,N_4320,N_4905);
nor U7742 (N_7742,N_274,N_331);
and U7743 (N_7743,N_4705,N_433);
and U7744 (N_7744,N_3313,N_4076);
and U7745 (N_7745,N_3948,N_3649);
or U7746 (N_7746,N_4807,N_2705);
nor U7747 (N_7747,N_4192,N_2738);
or U7748 (N_7748,N_1546,N_2453);
nand U7749 (N_7749,N_193,N_4049);
or U7750 (N_7750,N_560,N_2921);
xnor U7751 (N_7751,N_2047,N_255);
nand U7752 (N_7752,N_2768,N_4585);
nor U7753 (N_7753,N_1967,N_2042);
nand U7754 (N_7754,N_1977,N_381);
and U7755 (N_7755,N_3714,N_835);
or U7756 (N_7756,N_2595,N_4517);
and U7757 (N_7757,N_2399,N_1956);
nor U7758 (N_7758,N_4576,N_4387);
nor U7759 (N_7759,N_1880,N_3705);
nand U7760 (N_7760,N_1940,N_4620);
nor U7761 (N_7761,N_1155,N_1222);
nand U7762 (N_7762,N_4948,N_3823);
nand U7763 (N_7763,N_82,N_444);
xor U7764 (N_7764,N_2624,N_4849);
nor U7765 (N_7765,N_4959,N_1785);
xnor U7766 (N_7766,N_495,N_332);
and U7767 (N_7767,N_811,N_599);
xnor U7768 (N_7768,N_3627,N_748);
nand U7769 (N_7769,N_1404,N_1530);
and U7770 (N_7770,N_2217,N_1883);
or U7771 (N_7771,N_512,N_4597);
nor U7772 (N_7772,N_2895,N_3914);
and U7773 (N_7773,N_1485,N_2793);
nor U7774 (N_7774,N_4479,N_5);
or U7775 (N_7775,N_2261,N_2231);
xnor U7776 (N_7776,N_4453,N_3869);
xor U7777 (N_7777,N_1563,N_4222);
nand U7778 (N_7778,N_448,N_4214);
and U7779 (N_7779,N_3980,N_4152);
nor U7780 (N_7780,N_1867,N_4698);
or U7781 (N_7781,N_3008,N_3800);
nor U7782 (N_7782,N_3794,N_28);
and U7783 (N_7783,N_3255,N_1265);
and U7784 (N_7784,N_1298,N_632);
or U7785 (N_7785,N_121,N_1354);
xnor U7786 (N_7786,N_885,N_1642);
nor U7787 (N_7787,N_4137,N_981);
xnor U7788 (N_7788,N_2146,N_4305);
nand U7789 (N_7789,N_4124,N_107);
xor U7790 (N_7790,N_2786,N_4695);
nand U7791 (N_7791,N_2078,N_230);
or U7792 (N_7792,N_985,N_4263);
and U7793 (N_7793,N_418,N_1915);
nand U7794 (N_7794,N_1145,N_2341);
nor U7795 (N_7795,N_1259,N_2081);
and U7796 (N_7796,N_2727,N_4673);
nor U7797 (N_7797,N_4634,N_3519);
xnor U7798 (N_7798,N_2078,N_522);
nand U7799 (N_7799,N_3206,N_1943);
xnor U7800 (N_7800,N_1286,N_430);
and U7801 (N_7801,N_284,N_2970);
nor U7802 (N_7802,N_4909,N_3287);
xnor U7803 (N_7803,N_1012,N_4788);
nor U7804 (N_7804,N_1401,N_2141);
nor U7805 (N_7805,N_432,N_4277);
nor U7806 (N_7806,N_950,N_4965);
nand U7807 (N_7807,N_4117,N_691);
xnor U7808 (N_7808,N_632,N_4599);
or U7809 (N_7809,N_2957,N_1432);
nor U7810 (N_7810,N_1281,N_108);
or U7811 (N_7811,N_1504,N_3572);
xnor U7812 (N_7812,N_4333,N_1946);
xor U7813 (N_7813,N_1210,N_1087);
or U7814 (N_7814,N_1077,N_3846);
nand U7815 (N_7815,N_3179,N_583);
and U7816 (N_7816,N_2687,N_3112);
or U7817 (N_7817,N_741,N_4339);
nand U7818 (N_7818,N_3052,N_751);
nand U7819 (N_7819,N_3709,N_11);
xnor U7820 (N_7820,N_3709,N_3554);
nand U7821 (N_7821,N_2892,N_4398);
and U7822 (N_7822,N_496,N_396);
or U7823 (N_7823,N_4286,N_709);
nand U7824 (N_7824,N_3868,N_4529);
xnor U7825 (N_7825,N_4728,N_3187);
nor U7826 (N_7826,N_860,N_2384);
or U7827 (N_7827,N_531,N_2666);
xnor U7828 (N_7828,N_4947,N_3606);
xnor U7829 (N_7829,N_3705,N_805);
nor U7830 (N_7830,N_2225,N_1514);
or U7831 (N_7831,N_1124,N_440);
xor U7832 (N_7832,N_4295,N_3431);
nor U7833 (N_7833,N_4988,N_1035);
nor U7834 (N_7834,N_4599,N_3925);
xor U7835 (N_7835,N_4663,N_3764);
nor U7836 (N_7836,N_3143,N_4221);
nor U7837 (N_7837,N_4304,N_4340);
nor U7838 (N_7838,N_4720,N_2778);
or U7839 (N_7839,N_3373,N_2815);
nor U7840 (N_7840,N_2708,N_103);
nand U7841 (N_7841,N_4379,N_3088);
xnor U7842 (N_7842,N_3152,N_2137);
and U7843 (N_7843,N_3135,N_2167);
xnor U7844 (N_7844,N_3444,N_3958);
xnor U7845 (N_7845,N_4007,N_80);
nor U7846 (N_7846,N_3780,N_4879);
nor U7847 (N_7847,N_4671,N_149);
or U7848 (N_7848,N_137,N_3805);
and U7849 (N_7849,N_3920,N_4147);
and U7850 (N_7850,N_112,N_3353);
and U7851 (N_7851,N_2188,N_3779);
or U7852 (N_7852,N_4055,N_2805);
or U7853 (N_7853,N_625,N_1767);
xor U7854 (N_7854,N_970,N_4400);
xnor U7855 (N_7855,N_4429,N_4786);
and U7856 (N_7856,N_1809,N_756);
and U7857 (N_7857,N_4463,N_4810);
or U7858 (N_7858,N_4275,N_3250);
and U7859 (N_7859,N_4713,N_808);
xnor U7860 (N_7860,N_636,N_2350);
nand U7861 (N_7861,N_1523,N_2671);
and U7862 (N_7862,N_3464,N_3797);
nor U7863 (N_7863,N_2852,N_1754);
nand U7864 (N_7864,N_4733,N_42);
nand U7865 (N_7865,N_4932,N_3878);
nand U7866 (N_7866,N_1358,N_3999);
or U7867 (N_7867,N_3867,N_3696);
or U7868 (N_7868,N_4929,N_4748);
nand U7869 (N_7869,N_2592,N_1522);
or U7870 (N_7870,N_4247,N_2065);
xor U7871 (N_7871,N_480,N_3070);
or U7872 (N_7872,N_4521,N_3701);
xnor U7873 (N_7873,N_4031,N_1036);
or U7874 (N_7874,N_1301,N_3482);
nor U7875 (N_7875,N_4397,N_1047);
nand U7876 (N_7876,N_4078,N_3759);
nor U7877 (N_7877,N_2575,N_3133);
and U7878 (N_7878,N_1205,N_3891);
or U7879 (N_7879,N_3260,N_1155);
and U7880 (N_7880,N_2819,N_2824);
nand U7881 (N_7881,N_1983,N_1110);
nor U7882 (N_7882,N_595,N_937);
nand U7883 (N_7883,N_1949,N_2095);
nand U7884 (N_7884,N_771,N_2503);
or U7885 (N_7885,N_3742,N_1162);
xor U7886 (N_7886,N_990,N_2867);
nand U7887 (N_7887,N_35,N_3048);
xor U7888 (N_7888,N_30,N_1849);
or U7889 (N_7889,N_4006,N_1709);
nor U7890 (N_7890,N_2931,N_1969);
nor U7891 (N_7891,N_1538,N_1185);
or U7892 (N_7892,N_1144,N_1789);
or U7893 (N_7893,N_4575,N_365);
xnor U7894 (N_7894,N_3212,N_4070);
nor U7895 (N_7895,N_2069,N_3046);
and U7896 (N_7896,N_3373,N_1289);
nor U7897 (N_7897,N_4716,N_3297);
nand U7898 (N_7898,N_4833,N_3926);
xor U7899 (N_7899,N_737,N_3262);
and U7900 (N_7900,N_481,N_63);
nand U7901 (N_7901,N_762,N_4853);
and U7902 (N_7902,N_2623,N_3836);
and U7903 (N_7903,N_4523,N_4749);
and U7904 (N_7904,N_1796,N_176);
and U7905 (N_7905,N_3344,N_4215);
xor U7906 (N_7906,N_3203,N_800);
or U7907 (N_7907,N_1694,N_3944);
xnor U7908 (N_7908,N_4415,N_4968);
and U7909 (N_7909,N_3502,N_1869);
nor U7910 (N_7910,N_2890,N_494);
nand U7911 (N_7911,N_3333,N_2189);
or U7912 (N_7912,N_4680,N_1901);
nor U7913 (N_7913,N_3340,N_2838);
nand U7914 (N_7914,N_1160,N_432);
nand U7915 (N_7915,N_542,N_2836);
or U7916 (N_7916,N_3795,N_2383);
and U7917 (N_7917,N_4094,N_70);
nand U7918 (N_7918,N_1544,N_4984);
xnor U7919 (N_7919,N_4833,N_4718);
nand U7920 (N_7920,N_832,N_3441);
or U7921 (N_7921,N_1102,N_1991);
nand U7922 (N_7922,N_2813,N_262);
xor U7923 (N_7923,N_3983,N_205);
or U7924 (N_7924,N_3397,N_2447);
and U7925 (N_7925,N_1439,N_2632);
nand U7926 (N_7926,N_4168,N_3918);
or U7927 (N_7927,N_3072,N_4213);
nor U7928 (N_7928,N_353,N_1503);
nor U7929 (N_7929,N_1644,N_2009);
nand U7930 (N_7930,N_4876,N_3792);
nand U7931 (N_7931,N_1444,N_895);
xor U7932 (N_7932,N_1152,N_4214);
or U7933 (N_7933,N_2486,N_849);
or U7934 (N_7934,N_3815,N_3421);
xnor U7935 (N_7935,N_833,N_2847);
nor U7936 (N_7936,N_4695,N_4647);
and U7937 (N_7937,N_1445,N_3411);
xnor U7938 (N_7938,N_2944,N_4119);
xnor U7939 (N_7939,N_816,N_723);
xnor U7940 (N_7940,N_4317,N_4281);
nor U7941 (N_7941,N_2909,N_3243);
xnor U7942 (N_7942,N_4100,N_4377);
and U7943 (N_7943,N_1896,N_1094);
xnor U7944 (N_7944,N_3506,N_1070);
nand U7945 (N_7945,N_568,N_1206);
nand U7946 (N_7946,N_59,N_4237);
or U7947 (N_7947,N_4268,N_446);
xnor U7948 (N_7948,N_1994,N_1634);
nor U7949 (N_7949,N_2166,N_3574);
xnor U7950 (N_7950,N_4894,N_4327);
and U7951 (N_7951,N_3071,N_1059);
xor U7952 (N_7952,N_2985,N_1986);
nand U7953 (N_7953,N_67,N_461);
and U7954 (N_7954,N_2639,N_1443);
xor U7955 (N_7955,N_68,N_3818);
nor U7956 (N_7956,N_3530,N_459);
nor U7957 (N_7957,N_9,N_322);
and U7958 (N_7958,N_1562,N_1056);
nand U7959 (N_7959,N_2346,N_638);
nor U7960 (N_7960,N_2868,N_2932);
nand U7961 (N_7961,N_3842,N_1628);
xor U7962 (N_7962,N_3724,N_4870);
xor U7963 (N_7963,N_693,N_295);
nand U7964 (N_7964,N_1948,N_2750);
xor U7965 (N_7965,N_596,N_665);
nor U7966 (N_7966,N_2946,N_3364);
and U7967 (N_7967,N_3361,N_3607);
or U7968 (N_7968,N_3634,N_4791);
and U7969 (N_7969,N_3323,N_4741);
nor U7970 (N_7970,N_898,N_4843);
or U7971 (N_7971,N_2594,N_3673);
and U7972 (N_7972,N_184,N_4659);
or U7973 (N_7973,N_797,N_2439);
and U7974 (N_7974,N_1033,N_3255);
or U7975 (N_7975,N_1967,N_2292);
and U7976 (N_7976,N_655,N_2348);
nand U7977 (N_7977,N_1564,N_1782);
nor U7978 (N_7978,N_2885,N_4225);
nor U7979 (N_7979,N_436,N_1093);
nand U7980 (N_7980,N_3473,N_2952);
or U7981 (N_7981,N_670,N_3190);
xor U7982 (N_7982,N_2093,N_3481);
nor U7983 (N_7983,N_478,N_2175);
or U7984 (N_7984,N_953,N_4402);
xnor U7985 (N_7985,N_1803,N_4682);
xnor U7986 (N_7986,N_4812,N_1778);
and U7987 (N_7987,N_333,N_4744);
nand U7988 (N_7988,N_3653,N_1187);
and U7989 (N_7989,N_3799,N_3401);
xor U7990 (N_7990,N_1691,N_891);
xnor U7991 (N_7991,N_1683,N_4151);
nand U7992 (N_7992,N_2860,N_3129);
nor U7993 (N_7993,N_2459,N_4533);
or U7994 (N_7994,N_2394,N_106);
or U7995 (N_7995,N_2714,N_3664);
nor U7996 (N_7996,N_2652,N_2706);
or U7997 (N_7997,N_1389,N_4695);
or U7998 (N_7998,N_4966,N_94);
and U7999 (N_7999,N_3879,N_1746);
xnor U8000 (N_8000,N_3375,N_730);
nand U8001 (N_8001,N_123,N_923);
or U8002 (N_8002,N_4655,N_1808);
and U8003 (N_8003,N_4192,N_3987);
xor U8004 (N_8004,N_144,N_1949);
nor U8005 (N_8005,N_4837,N_2919);
nor U8006 (N_8006,N_1893,N_99);
nand U8007 (N_8007,N_2403,N_4012);
xor U8008 (N_8008,N_939,N_1304);
nand U8009 (N_8009,N_4194,N_1864);
nor U8010 (N_8010,N_266,N_4224);
nand U8011 (N_8011,N_128,N_4511);
or U8012 (N_8012,N_2709,N_578);
nand U8013 (N_8013,N_3753,N_644);
xor U8014 (N_8014,N_3155,N_508);
nor U8015 (N_8015,N_775,N_3424);
nand U8016 (N_8016,N_2275,N_4786);
and U8017 (N_8017,N_3148,N_2709);
or U8018 (N_8018,N_4398,N_1803);
or U8019 (N_8019,N_2609,N_2861);
nand U8020 (N_8020,N_2649,N_2543);
or U8021 (N_8021,N_1110,N_341);
xor U8022 (N_8022,N_298,N_3507);
nand U8023 (N_8023,N_3459,N_1264);
nor U8024 (N_8024,N_4154,N_4135);
xor U8025 (N_8025,N_4663,N_2403);
nor U8026 (N_8026,N_930,N_4158);
and U8027 (N_8027,N_3719,N_3439);
or U8028 (N_8028,N_2555,N_4189);
nand U8029 (N_8029,N_1227,N_1345);
and U8030 (N_8030,N_2707,N_3689);
and U8031 (N_8031,N_76,N_3980);
or U8032 (N_8032,N_173,N_4119);
nand U8033 (N_8033,N_2369,N_12);
nor U8034 (N_8034,N_2952,N_952);
or U8035 (N_8035,N_1702,N_2344);
nand U8036 (N_8036,N_3882,N_2226);
or U8037 (N_8037,N_3055,N_4990);
and U8038 (N_8038,N_4404,N_670);
or U8039 (N_8039,N_3929,N_758);
and U8040 (N_8040,N_1643,N_1066);
and U8041 (N_8041,N_1671,N_4436);
and U8042 (N_8042,N_76,N_2740);
nor U8043 (N_8043,N_903,N_2006);
nand U8044 (N_8044,N_4907,N_22);
and U8045 (N_8045,N_86,N_4907);
nor U8046 (N_8046,N_4727,N_2883);
nand U8047 (N_8047,N_2695,N_2155);
xor U8048 (N_8048,N_1924,N_2172);
nand U8049 (N_8049,N_3213,N_675);
and U8050 (N_8050,N_956,N_652);
nand U8051 (N_8051,N_2964,N_4242);
and U8052 (N_8052,N_1952,N_3371);
nor U8053 (N_8053,N_3476,N_1596);
nor U8054 (N_8054,N_2713,N_1226);
and U8055 (N_8055,N_4595,N_246);
nor U8056 (N_8056,N_1411,N_3089);
xnor U8057 (N_8057,N_2804,N_3349);
or U8058 (N_8058,N_1317,N_2110);
xor U8059 (N_8059,N_3754,N_3423);
nand U8060 (N_8060,N_2870,N_1672);
xnor U8061 (N_8061,N_2705,N_4747);
or U8062 (N_8062,N_1636,N_3432);
xnor U8063 (N_8063,N_2357,N_3577);
or U8064 (N_8064,N_3460,N_2601);
nand U8065 (N_8065,N_4890,N_3056);
nand U8066 (N_8066,N_3640,N_1596);
nand U8067 (N_8067,N_2126,N_2324);
or U8068 (N_8068,N_3373,N_3837);
nand U8069 (N_8069,N_3698,N_4238);
xnor U8070 (N_8070,N_3120,N_4441);
nand U8071 (N_8071,N_2679,N_2962);
xnor U8072 (N_8072,N_3327,N_2777);
xor U8073 (N_8073,N_1481,N_775);
or U8074 (N_8074,N_743,N_2728);
or U8075 (N_8075,N_853,N_3678);
nor U8076 (N_8076,N_2064,N_1637);
or U8077 (N_8077,N_3325,N_3447);
nor U8078 (N_8078,N_3492,N_3736);
xnor U8079 (N_8079,N_993,N_1847);
xnor U8080 (N_8080,N_3731,N_228);
or U8081 (N_8081,N_3058,N_1710);
and U8082 (N_8082,N_4485,N_4149);
nor U8083 (N_8083,N_4476,N_3146);
and U8084 (N_8084,N_314,N_2203);
xor U8085 (N_8085,N_369,N_2785);
nand U8086 (N_8086,N_923,N_198);
or U8087 (N_8087,N_2842,N_586);
or U8088 (N_8088,N_2482,N_2013);
nand U8089 (N_8089,N_3189,N_3084);
or U8090 (N_8090,N_989,N_2160);
or U8091 (N_8091,N_1068,N_1566);
nand U8092 (N_8092,N_3921,N_2236);
nand U8093 (N_8093,N_2581,N_3172);
nand U8094 (N_8094,N_464,N_3600);
xor U8095 (N_8095,N_1659,N_2977);
or U8096 (N_8096,N_296,N_4387);
xor U8097 (N_8097,N_3926,N_929);
and U8098 (N_8098,N_2288,N_1225);
and U8099 (N_8099,N_1061,N_303);
and U8100 (N_8100,N_3111,N_617);
nand U8101 (N_8101,N_2061,N_4102);
or U8102 (N_8102,N_4817,N_941);
or U8103 (N_8103,N_3300,N_2241);
and U8104 (N_8104,N_1356,N_1869);
xnor U8105 (N_8105,N_2407,N_268);
or U8106 (N_8106,N_3124,N_1886);
or U8107 (N_8107,N_2499,N_229);
and U8108 (N_8108,N_2885,N_4069);
xnor U8109 (N_8109,N_2592,N_1728);
xnor U8110 (N_8110,N_2512,N_3049);
and U8111 (N_8111,N_2579,N_2790);
and U8112 (N_8112,N_2776,N_3355);
xnor U8113 (N_8113,N_353,N_4053);
nand U8114 (N_8114,N_1708,N_2787);
or U8115 (N_8115,N_214,N_54);
xor U8116 (N_8116,N_1564,N_3959);
and U8117 (N_8117,N_4064,N_2689);
nor U8118 (N_8118,N_1314,N_1439);
or U8119 (N_8119,N_1950,N_3112);
or U8120 (N_8120,N_1402,N_2051);
or U8121 (N_8121,N_3341,N_3795);
nor U8122 (N_8122,N_1258,N_2448);
nand U8123 (N_8123,N_1226,N_1558);
nor U8124 (N_8124,N_3276,N_4492);
or U8125 (N_8125,N_2163,N_3056);
or U8126 (N_8126,N_2900,N_502);
nor U8127 (N_8127,N_4825,N_1267);
nand U8128 (N_8128,N_3193,N_682);
or U8129 (N_8129,N_32,N_3189);
nor U8130 (N_8130,N_2839,N_4463);
and U8131 (N_8131,N_4129,N_3251);
nand U8132 (N_8132,N_4504,N_4203);
nor U8133 (N_8133,N_4896,N_2794);
nand U8134 (N_8134,N_801,N_3276);
nand U8135 (N_8135,N_1265,N_2666);
or U8136 (N_8136,N_4989,N_482);
nand U8137 (N_8137,N_4517,N_725);
and U8138 (N_8138,N_2498,N_1458);
or U8139 (N_8139,N_4905,N_698);
nor U8140 (N_8140,N_753,N_839);
or U8141 (N_8141,N_761,N_4012);
nor U8142 (N_8142,N_538,N_3973);
nand U8143 (N_8143,N_1131,N_1802);
or U8144 (N_8144,N_3090,N_4631);
or U8145 (N_8145,N_4390,N_3500);
nand U8146 (N_8146,N_952,N_4414);
or U8147 (N_8147,N_1594,N_4991);
xnor U8148 (N_8148,N_829,N_405);
xor U8149 (N_8149,N_1455,N_2303);
and U8150 (N_8150,N_2391,N_2250);
xnor U8151 (N_8151,N_4683,N_3437);
xnor U8152 (N_8152,N_4455,N_1546);
and U8153 (N_8153,N_968,N_1206);
or U8154 (N_8154,N_3429,N_4586);
xnor U8155 (N_8155,N_3139,N_4661);
nand U8156 (N_8156,N_1334,N_3496);
xnor U8157 (N_8157,N_4024,N_2792);
nor U8158 (N_8158,N_397,N_4290);
nor U8159 (N_8159,N_4530,N_3790);
or U8160 (N_8160,N_912,N_1405);
and U8161 (N_8161,N_905,N_1471);
and U8162 (N_8162,N_1197,N_4398);
or U8163 (N_8163,N_3129,N_2041);
or U8164 (N_8164,N_3540,N_1593);
nor U8165 (N_8165,N_2898,N_2273);
or U8166 (N_8166,N_3956,N_1017);
and U8167 (N_8167,N_745,N_2484);
nand U8168 (N_8168,N_3365,N_3582);
nor U8169 (N_8169,N_4015,N_791);
or U8170 (N_8170,N_64,N_3391);
nor U8171 (N_8171,N_1392,N_2100);
xnor U8172 (N_8172,N_3918,N_4744);
nor U8173 (N_8173,N_1521,N_1798);
xor U8174 (N_8174,N_2160,N_4324);
nand U8175 (N_8175,N_1776,N_3793);
xor U8176 (N_8176,N_944,N_3200);
nand U8177 (N_8177,N_2416,N_1139);
nor U8178 (N_8178,N_3165,N_1470);
and U8179 (N_8179,N_3710,N_1744);
or U8180 (N_8180,N_4058,N_1873);
nand U8181 (N_8181,N_3659,N_29);
or U8182 (N_8182,N_2019,N_997);
nand U8183 (N_8183,N_4064,N_427);
or U8184 (N_8184,N_1800,N_1697);
xnor U8185 (N_8185,N_3173,N_3842);
and U8186 (N_8186,N_1762,N_1919);
nor U8187 (N_8187,N_3842,N_2309);
xnor U8188 (N_8188,N_996,N_2554);
nand U8189 (N_8189,N_2105,N_933);
nor U8190 (N_8190,N_1012,N_3351);
or U8191 (N_8191,N_1601,N_2014);
xor U8192 (N_8192,N_815,N_4669);
nor U8193 (N_8193,N_1362,N_1338);
nor U8194 (N_8194,N_2610,N_4174);
xor U8195 (N_8195,N_3929,N_2183);
nand U8196 (N_8196,N_835,N_1874);
or U8197 (N_8197,N_3385,N_740);
nor U8198 (N_8198,N_4760,N_3213);
and U8199 (N_8199,N_2451,N_4754);
xor U8200 (N_8200,N_1118,N_1436);
nand U8201 (N_8201,N_4215,N_2980);
or U8202 (N_8202,N_4802,N_3693);
and U8203 (N_8203,N_3661,N_832);
and U8204 (N_8204,N_3173,N_3577);
and U8205 (N_8205,N_4786,N_2438);
or U8206 (N_8206,N_3202,N_3661);
or U8207 (N_8207,N_1052,N_538);
xnor U8208 (N_8208,N_192,N_926);
or U8209 (N_8209,N_699,N_651);
or U8210 (N_8210,N_3896,N_3187);
nor U8211 (N_8211,N_3265,N_2775);
nor U8212 (N_8212,N_4774,N_3484);
nand U8213 (N_8213,N_3775,N_973);
nand U8214 (N_8214,N_1090,N_634);
xnor U8215 (N_8215,N_2141,N_2714);
and U8216 (N_8216,N_2838,N_2978);
and U8217 (N_8217,N_317,N_3452);
or U8218 (N_8218,N_2391,N_4060);
and U8219 (N_8219,N_152,N_367);
or U8220 (N_8220,N_3649,N_1470);
xor U8221 (N_8221,N_2355,N_3238);
nand U8222 (N_8222,N_1521,N_3833);
nor U8223 (N_8223,N_994,N_3573);
and U8224 (N_8224,N_4342,N_2822);
xor U8225 (N_8225,N_4825,N_3341);
and U8226 (N_8226,N_3339,N_1269);
nand U8227 (N_8227,N_4683,N_4273);
xor U8228 (N_8228,N_4193,N_524);
or U8229 (N_8229,N_167,N_3844);
nand U8230 (N_8230,N_2940,N_3437);
nand U8231 (N_8231,N_3741,N_3204);
nand U8232 (N_8232,N_1285,N_427);
xnor U8233 (N_8233,N_3188,N_3140);
nand U8234 (N_8234,N_489,N_3550);
xnor U8235 (N_8235,N_305,N_3520);
xor U8236 (N_8236,N_4506,N_3325);
nor U8237 (N_8237,N_4609,N_4162);
or U8238 (N_8238,N_3808,N_2897);
or U8239 (N_8239,N_4306,N_3105);
nor U8240 (N_8240,N_3540,N_4715);
and U8241 (N_8241,N_4763,N_4082);
nor U8242 (N_8242,N_4655,N_4007);
or U8243 (N_8243,N_3452,N_2161);
and U8244 (N_8244,N_1981,N_1518);
and U8245 (N_8245,N_2686,N_2948);
xnor U8246 (N_8246,N_4148,N_1032);
and U8247 (N_8247,N_1611,N_105);
xor U8248 (N_8248,N_3514,N_3683);
xnor U8249 (N_8249,N_2334,N_3479);
or U8250 (N_8250,N_3574,N_2955);
or U8251 (N_8251,N_2205,N_4749);
and U8252 (N_8252,N_2178,N_1518);
xor U8253 (N_8253,N_4311,N_1603);
and U8254 (N_8254,N_3933,N_2657);
nand U8255 (N_8255,N_3217,N_2463);
nor U8256 (N_8256,N_327,N_3194);
and U8257 (N_8257,N_1660,N_4535);
xnor U8258 (N_8258,N_2297,N_2645);
xnor U8259 (N_8259,N_639,N_1923);
or U8260 (N_8260,N_1679,N_4888);
nor U8261 (N_8261,N_2117,N_3596);
and U8262 (N_8262,N_3034,N_3084);
nor U8263 (N_8263,N_4871,N_3728);
and U8264 (N_8264,N_2431,N_1584);
and U8265 (N_8265,N_57,N_55);
nand U8266 (N_8266,N_333,N_2703);
or U8267 (N_8267,N_1157,N_28);
xnor U8268 (N_8268,N_1112,N_3305);
nand U8269 (N_8269,N_4934,N_2851);
or U8270 (N_8270,N_72,N_198);
nor U8271 (N_8271,N_3888,N_2378);
and U8272 (N_8272,N_4592,N_2534);
nand U8273 (N_8273,N_629,N_671);
nand U8274 (N_8274,N_937,N_3025);
nand U8275 (N_8275,N_300,N_3819);
and U8276 (N_8276,N_4927,N_271);
nor U8277 (N_8277,N_2452,N_1350);
nor U8278 (N_8278,N_3414,N_1426);
nand U8279 (N_8279,N_279,N_4876);
nand U8280 (N_8280,N_2554,N_4592);
nand U8281 (N_8281,N_4843,N_2300);
nor U8282 (N_8282,N_1635,N_3193);
xnor U8283 (N_8283,N_2515,N_4569);
xor U8284 (N_8284,N_3782,N_2702);
or U8285 (N_8285,N_214,N_2775);
nand U8286 (N_8286,N_288,N_619);
nor U8287 (N_8287,N_557,N_4590);
nor U8288 (N_8288,N_2345,N_1828);
nor U8289 (N_8289,N_3746,N_4006);
nand U8290 (N_8290,N_2793,N_779);
nor U8291 (N_8291,N_4774,N_3876);
nor U8292 (N_8292,N_3042,N_1949);
and U8293 (N_8293,N_4565,N_3307);
or U8294 (N_8294,N_1065,N_4307);
nand U8295 (N_8295,N_285,N_4122);
or U8296 (N_8296,N_2827,N_2740);
and U8297 (N_8297,N_1734,N_3295);
nor U8298 (N_8298,N_3383,N_839);
and U8299 (N_8299,N_1492,N_3092);
nor U8300 (N_8300,N_2092,N_2156);
and U8301 (N_8301,N_3997,N_3489);
nand U8302 (N_8302,N_107,N_1618);
or U8303 (N_8303,N_1550,N_4081);
xnor U8304 (N_8304,N_2762,N_1892);
xor U8305 (N_8305,N_4351,N_4376);
nor U8306 (N_8306,N_2809,N_4541);
nand U8307 (N_8307,N_489,N_1450);
nand U8308 (N_8308,N_4522,N_850);
nand U8309 (N_8309,N_1294,N_181);
nor U8310 (N_8310,N_4874,N_4647);
xnor U8311 (N_8311,N_2975,N_2610);
nand U8312 (N_8312,N_174,N_3546);
xor U8313 (N_8313,N_4134,N_2297);
or U8314 (N_8314,N_895,N_4071);
nor U8315 (N_8315,N_4277,N_665);
and U8316 (N_8316,N_1268,N_1784);
or U8317 (N_8317,N_3468,N_4344);
or U8318 (N_8318,N_1876,N_1112);
nor U8319 (N_8319,N_2768,N_633);
xor U8320 (N_8320,N_2600,N_1461);
nand U8321 (N_8321,N_981,N_1926);
or U8322 (N_8322,N_2834,N_4186);
xor U8323 (N_8323,N_1623,N_1803);
and U8324 (N_8324,N_132,N_298);
nor U8325 (N_8325,N_1553,N_3451);
xnor U8326 (N_8326,N_3,N_4730);
nand U8327 (N_8327,N_3946,N_4349);
nor U8328 (N_8328,N_988,N_1308);
nor U8329 (N_8329,N_4267,N_1193);
and U8330 (N_8330,N_223,N_991);
nand U8331 (N_8331,N_2263,N_2676);
nor U8332 (N_8332,N_2441,N_910);
or U8333 (N_8333,N_3524,N_2539);
nand U8334 (N_8334,N_2077,N_1596);
or U8335 (N_8335,N_291,N_3195);
nor U8336 (N_8336,N_3186,N_211);
and U8337 (N_8337,N_1532,N_1487);
xor U8338 (N_8338,N_534,N_1329);
nor U8339 (N_8339,N_4903,N_1141);
and U8340 (N_8340,N_3185,N_4310);
nor U8341 (N_8341,N_4396,N_2508);
xnor U8342 (N_8342,N_1412,N_2927);
nor U8343 (N_8343,N_748,N_1204);
xnor U8344 (N_8344,N_4665,N_1165);
xor U8345 (N_8345,N_4491,N_2253);
nor U8346 (N_8346,N_4081,N_1233);
or U8347 (N_8347,N_839,N_2841);
or U8348 (N_8348,N_3943,N_542);
nor U8349 (N_8349,N_2557,N_2352);
and U8350 (N_8350,N_1638,N_116);
nand U8351 (N_8351,N_4062,N_4538);
xor U8352 (N_8352,N_2088,N_2824);
and U8353 (N_8353,N_598,N_1295);
or U8354 (N_8354,N_3614,N_3374);
xor U8355 (N_8355,N_4370,N_4016);
xor U8356 (N_8356,N_3549,N_2169);
and U8357 (N_8357,N_3808,N_2315);
and U8358 (N_8358,N_3888,N_43);
and U8359 (N_8359,N_2740,N_780);
xor U8360 (N_8360,N_3143,N_552);
nor U8361 (N_8361,N_1930,N_1468);
nand U8362 (N_8362,N_770,N_2268);
or U8363 (N_8363,N_812,N_4045);
and U8364 (N_8364,N_4649,N_479);
nor U8365 (N_8365,N_3934,N_3653);
xnor U8366 (N_8366,N_433,N_2588);
nor U8367 (N_8367,N_4275,N_3999);
or U8368 (N_8368,N_4681,N_1266);
nand U8369 (N_8369,N_2252,N_943);
xnor U8370 (N_8370,N_3923,N_2205);
xnor U8371 (N_8371,N_3648,N_1191);
xnor U8372 (N_8372,N_3182,N_557);
nor U8373 (N_8373,N_93,N_1245);
xnor U8374 (N_8374,N_1806,N_2407);
nand U8375 (N_8375,N_3865,N_794);
xor U8376 (N_8376,N_909,N_3310);
and U8377 (N_8377,N_1064,N_1669);
and U8378 (N_8378,N_1499,N_2983);
or U8379 (N_8379,N_571,N_4133);
nor U8380 (N_8380,N_1809,N_1510);
xor U8381 (N_8381,N_1581,N_1592);
or U8382 (N_8382,N_178,N_3127);
or U8383 (N_8383,N_1472,N_2130);
xnor U8384 (N_8384,N_4238,N_1961);
nor U8385 (N_8385,N_805,N_209);
nand U8386 (N_8386,N_1998,N_228);
and U8387 (N_8387,N_819,N_3685);
xnor U8388 (N_8388,N_152,N_3871);
or U8389 (N_8389,N_619,N_4192);
xnor U8390 (N_8390,N_1601,N_3963);
and U8391 (N_8391,N_4468,N_3610);
nand U8392 (N_8392,N_2015,N_1989);
or U8393 (N_8393,N_3171,N_2250);
nand U8394 (N_8394,N_2315,N_2990);
nor U8395 (N_8395,N_944,N_4297);
or U8396 (N_8396,N_2776,N_3361);
xor U8397 (N_8397,N_1498,N_1361);
or U8398 (N_8398,N_2523,N_4679);
xor U8399 (N_8399,N_4722,N_4631);
xnor U8400 (N_8400,N_234,N_2057);
and U8401 (N_8401,N_653,N_3084);
and U8402 (N_8402,N_119,N_2768);
or U8403 (N_8403,N_289,N_494);
or U8404 (N_8404,N_586,N_3478);
and U8405 (N_8405,N_2462,N_18);
or U8406 (N_8406,N_2605,N_3210);
xor U8407 (N_8407,N_2266,N_2188);
nor U8408 (N_8408,N_968,N_665);
nand U8409 (N_8409,N_2084,N_2582);
and U8410 (N_8410,N_4719,N_3255);
nand U8411 (N_8411,N_225,N_945);
nor U8412 (N_8412,N_4389,N_4062);
xor U8413 (N_8413,N_3058,N_4354);
xnor U8414 (N_8414,N_4355,N_4245);
xnor U8415 (N_8415,N_1746,N_2630);
nand U8416 (N_8416,N_155,N_3346);
nor U8417 (N_8417,N_1681,N_2112);
nor U8418 (N_8418,N_4927,N_1750);
and U8419 (N_8419,N_1703,N_2510);
or U8420 (N_8420,N_2219,N_1184);
nor U8421 (N_8421,N_4225,N_2683);
and U8422 (N_8422,N_1272,N_4911);
nor U8423 (N_8423,N_202,N_2060);
or U8424 (N_8424,N_176,N_258);
xnor U8425 (N_8425,N_3259,N_2393);
nor U8426 (N_8426,N_2165,N_3764);
nor U8427 (N_8427,N_4170,N_384);
nor U8428 (N_8428,N_528,N_1129);
or U8429 (N_8429,N_2126,N_4846);
or U8430 (N_8430,N_627,N_1156);
xor U8431 (N_8431,N_3194,N_3605);
and U8432 (N_8432,N_2912,N_4206);
and U8433 (N_8433,N_4560,N_4899);
or U8434 (N_8434,N_231,N_2639);
xnor U8435 (N_8435,N_4397,N_2196);
nor U8436 (N_8436,N_2949,N_1269);
and U8437 (N_8437,N_4477,N_3061);
or U8438 (N_8438,N_4401,N_2459);
nor U8439 (N_8439,N_1136,N_530);
nor U8440 (N_8440,N_4951,N_2002);
and U8441 (N_8441,N_629,N_2108);
or U8442 (N_8442,N_1284,N_2840);
or U8443 (N_8443,N_2476,N_82);
nand U8444 (N_8444,N_2472,N_1306);
or U8445 (N_8445,N_3759,N_3469);
nor U8446 (N_8446,N_12,N_1795);
nor U8447 (N_8447,N_4989,N_4831);
nand U8448 (N_8448,N_2793,N_1693);
or U8449 (N_8449,N_2372,N_2082);
or U8450 (N_8450,N_2232,N_252);
or U8451 (N_8451,N_2440,N_853);
nand U8452 (N_8452,N_3468,N_4281);
and U8453 (N_8453,N_3692,N_845);
and U8454 (N_8454,N_4989,N_3717);
or U8455 (N_8455,N_3374,N_1533);
nand U8456 (N_8456,N_1193,N_888);
and U8457 (N_8457,N_3213,N_2633);
nor U8458 (N_8458,N_4031,N_2277);
nor U8459 (N_8459,N_2782,N_3092);
and U8460 (N_8460,N_2678,N_1873);
or U8461 (N_8461,N_3562,N_4928);
and U8462 (N_8462,N_1585,N_1983);
xnor U8463 (N_8463,N_719,N_623);
and U8464 (N_8464,N_787,N_2238);
and U8465 (N_8465,N_1329,N_4887);
or U8466 (N_8466,N_4149,N_3116);
and U8467 (N_8467,N_823,N_3135);
nand U8468 (N_8468,N_3750,N_3175);
nor U8469 (N_8469,N_1676,N_868);
nor U8470 (N_8470,N_280,N_3962);
and U8471 (N_8471,N_1876,N_3201);
or U8472 (N_8472,N_2119,N_3660);
xor U8473 (N_8473,N_3948,N_4299);
or U8474 (N_8474,N_4724,N_4908);
or U8475 (N_8475,N_1359,N_2790);
nand U8476 (N_8476,N_3333,N_2270);
nor U8477 (N_8477,N_4325,N_1540);
and U8478 (N_8478,N_1627,N_1054);
nor U8479 (N_8479,N_516,N_4611);
or U8480 (N_8480,N_1310,N_2331);
or U8481 (N_8481,N_2975,N_2541);
nor U8482 (N_8482,N_1820,N_469);
xor U8483 (N_8483,N_218,N_3408);
nand U8484 (N_8484,N_2751,N_4050);
or U8485 (N_8485,N_2031,N_2478);
or U8486 (N_8486,N_1307,N_870);
xnor U8487 (N_8487,N_274,N_1981);
nand U8488 (N_8488,N_2567,N_694);
nor U8489 (N_8489,N_1813,N_1107);
nor U8490 (N_8490,N_4737,N_3891);
nor U8491 (N_8491,N_1571,N_334);
and U8492 (N_8492,N_734,N_4011);
nand U8493 (N_8493,N_2500,N_1202);
and U8494 (N_8494,N_1101,N_2708);
or U8495 (N_8495,N_4665,N_1622);
nand U8496 (N_8496,N_4033,N_4788);
xnor U8497 (N_8497,N_2159,N_2018);
xor U8498 (N_8498,N_3231,N_4963);
or U8499 (N_8499,N_198,N_2162);
or U8500 (N_8500,N_1880,N_213);
nand U8501 (N_8501,N_1614,N_2637);
and U8502 (N_8502,N_4237,N_2534);
and U8503 (N_8503,N_3687,N_4423);
or U8504 (N_8504,N_1161,N_1343);
xor U8505 (N_8505,N_3931,N_145);
and U8506 (N_8506,N_4329,N_2826);
nand U8507 (N_8507,N_1892,N_327);
nor U8508 (N_8508,N_748,N_1667);
and U8509 (N_8509,N_43,N_1791);
or U8510 (N_8510,N_523,N_1093);
and U8511 (N_8511,N_3117,N_2214);
nand U8512 (N_8512,N_3770,N_977);
or U8513 (N_8513,N_4964,N_2450);
nand U8514 (N_8514,N_4272,N_1340);
and U8515 (N_8515,N_3339,N_3245);
nand U8516 (N_8516,N_2661,N_2117);
nor U8517 (N_8517,N_955,N_3855);
nor U8518 (N_8518,N_563,N_353);
or U8519 (N_8519,N_3689,N_245);
nand U8520 (N_8520,N_1124,N_4072);
xor U8521 (N_8521,N_2145,N_2799);
xor U8522 (N_8522,N_4178,N_1381);
or U8523 (N_8523,N_1858,N_1560);
and U8524 (N_8524,N_611,N_3928);
and U8525 (N_8525,N_1499,N_2405);
nor U8526 (N_8526,N_2851,N_4280);
and U8527 (N_8527,N_4305,N_203);
nand U8528 (N_8528,N_157,N_3088);
nor U8529 (N_8529,N_2896,N_4374);
and U8530 (N_8530,N_3354,N_2907);
xnor U8531 (N_8531,N_755,N_1064);
and U8532 (N_8532,N_3348,N_2360);
nand U8533 (N_8533,N_3018,N_1441);
and U8534 (N_8534,N_1762,N_1428);
and U8535 (N_8535,N_4901,N_1258);
nand U8536 (N_8536,N_4003,N_3883);
nor U8537 (N_8537,N_3926,N_1796);
or U8538 (N_8538,N_3087,N_3383);
nand U8539 (N_8539,N_903,N_3791);
xor U8540 (N_8540,N_3613,N_1732);
and U8541 (N_8541,N_3068,N_1347);
or U8542 (N_8542,N_4698,N_455);
nor U8543 (N_8543,N_1971,N_2657);
or U8544 (N_8544,N_1462,N_3909);
nor U8545 (N_8545,N_2321,N_370);
nor U8546 (N_8546,N_1146,N_1995);
nor U8547 (N_8547,N_2059,N_2795);
nand U8548 (N_8548,N_956,N_4602);
nand U8549 (N_8549,N_3151,N_2130);
xnor U8550 (N_8550,N_1290,N_2312);
or U8551 (N_8551,N_2324,N_3966);
xor U8552 (N_8552,N_2323,N_2944);
nand U8553 (N_8553,N_1904,N_1111);
nor U8554 (N_8554,N_4475,N_2561);
or U8555 (N_8555,N_3251,N_4119);
nand U8556 (N_8556,N_2111,N_613);
nand U8557 (N_8557,N_4597,N_383);
nand U8558 (N_8558,N_2111,N_1031);
and U8559 (N_8559,N_2460,N_2318);
nand U8560 (N_8560,N_1867,N_2887);
and U8561 (N_8561,N_2197,N_4688);
and U8562 (N_8562,N_526,N_3209);
and U8563 (N_8563,N_4999,N_2534);
nand U8564 (N_8564,N_3556,N_272);
nand U8565 (N_8565,N_4438,N_2402);
or U8566 (N_8566,N_4822,N_486);
nor U8567 (N_8567,N_3592,N_304);
nand U8568 (N_8568,N_896,N_4278);
nor U8569 (N_8569,N_2009,N_1874);
nor U8570 (N_8570,N_4539,N_3997);
nor U8571 (N_8571,N_2663,N_4903);
or U8572 (N_8572,N_2855,N_3751);
nand U8573 (N_8573,N_1664,N_4851);
xor U8574 (N_8574,N_2478,N_4873);
or U8575 (N_8575,N_871,N_2354);
or U8576 (N_8576,N_3759,N_2636);
nand U8577 (N_8577,N_4103,N_4275);
nand U8578 (N_8578,N_2365,N_467);
nand U8579 (N_8579,N_4225,N_3042);
and U8580 (N_8580,N_2264,N_1336);
or U8581 (N_8581,N_4279,N_1374);
xor U8582 (N_8582,N_583,N_151);
or U8583 (N_8583,N_2180,N_1908);
nor U8584 (N_8584,N_2496,N_2598);
nor U8585 (N_8585,N_1214,N_2517);
xor U8586 (N_8586,N_1884,N_3853);
xor U8587 (N_8587,N_2471,N_781);
xnor U8588 (N_8588,N_1744,N_926);
and U8589 (N_8589,N_4904,N_4899);
xor U8590 (N_8590,N_1579,N_2037);
or U8591 (N_8591,N_508,N_2713);
and U8592 (N_8592,N_1960,N_4792);
xnor U8593 (N_8593,N_2709,N_301);
xnor U8594 (N_8594,N_2864,N_4899);
nor U8595 (N_8595,N_3585,N_4394);
xnor U8596 (N_8596,N_983,N_4890);
nor U8597 (N_8597,N_574,N_9);
or U8598 (N_8598,N_4348,N_4949);
and U8599 (N_8599,N_1755,N_3963);
and U8600 (N_8600,N_58,N_1673);
and U8601 (N_8601,N_4823,N_2581);
or U8602 (N_8602,N_4920,N_2000);
nand U8603 (N_8603,N_3587,N_2700);
nand U8604 (N_8604,N_3648,N_452);
xnor U8605 (N_8605,N_1045,N_4483);
xor U8606 (N_8606,N_4389,N_4574);
nor U8607 (N_8607,N_2246,N_968);
or U8608 (N_8608,N_2659,N_3245);
or U8609 (N_8609,N_1354,N_228);
xor U8610 (N_8610,N_2978,N_3463);
or U8611 (N_8611,N_739,N_33);
and U8612 (N_8612,N_3628,N_2897);
nand U8613 (N_8613,N_581,N_233);
and U8614 (N_8614,N_2378,N_2988);
or U8615 (N_8615,N_3749,N_327);
xnor U8616 (N_8616,N_3347,N_2126);
nand U8617 (N_8617,N_2325,N_826);
nand U8618 (N_8618,N_276,N_1412);
xor U8619 (N_8619,N_205,N_4677);
xor U8620 (N_8620,N_2630,N_1912);
nand U8621 (N_8621,N_2862,N_3170);
nor U8622 (N_8622,N_3064,N_2647);
or U8623 (N_8623,N_1883,N_4241);
nand U8624 (N_8624,N_4783,N_526);
xnor U8625 (N_8625,N_383,N_3246);
xnor U8626 (N_8626,N_1857,N_1207);
and U8627 (N_8627,N_217,N_2899);
xor U8628 (N_8628,N_3147,N_4718);
nand U8629 (N_8629,N_3676,N_2246);
or U8630 (N_8630,N_4560,N_662);
xnor U8631 (N_8631,N_431,N_1793);
nor U8632 (N_8632,N_1724,N_3947);
nand U8633 (N_8633,N_4093,N_1577);
and U8634 (N_8634,N_3985,N_1751);
xnor U8635 (N_8635,N_3123,N_2536);
nand U8636 (N_8636,N_296,N_3149);
xnor U8637 (N_8637,N_977,N_4323);
xnor U8638 (N_8638,N_2880,N_2520);
and U8639 (N_8639,N_2713,N_2800);
xnor U8640 (N_8640,N_1718,N_1203);
xor U8641 (N_8641,N_1452,N_1631);
nor U8642 (N_8642,N_4935,N_2680);
and U8643 (N_8643,N_2288,N_3216);
and U8644 (N_8644,N_2295,N_3600);
xnor U8645 (N_8645,N_3049,N_2432);
xnor U8646 (N_8646,N_3679,N_2117);
and U8647 (N_8647,N_3816,N_4898);
nand U8648 (N_8648,N_1538,N_3378);
nor U8649 (N_8649,N_2032,N_445);
nor U8650 (N_8650,N_264,N_3048);
xnor U8651 (N_8651,N_3829,N_4983);
nand U8652 (N_8652,N_4553,N_2556);
and U8653 (N_8653,N_889,N_1171);
and U8654 (N_8654,N_2360,N_3556);
and U8655 (N_8655,N_1382,N_2199);
or U8656 (N_8656,N_2608,N_3604);
and U8657 (N_8657,N_3476,N_4814);
xnor U8658 (N_8658,N_4412,N_4434);
and U8659 (N_8659,N_4730,N_4984);
xnor U8660 (N_8660,N_3417,N_196);
nor U8661 (N_8661,N_3110,N_1206);
and U8662 (N_8662,N_4056,N_2979);
xor U8663 (N_8663,N_596,N_1059);
nand U8664 (N_8664,N_2890,N_1081);
and U8665 (N_8665,N_3614,N_2965);
nor U8666 (N_8666,N_4009,N_1460);
xnor U8667 (N_8667,N_544,N_3604);
and U8668 (N_8668,N_3761,N_2054);
nor U8669 (N_8669,N_62,N_3946);
nand U8670 (N_8670,N_116,N_2958);
nand U8671 (N_8671,N_2028,N_746);
nand U8672 (N_8672,N_2237,N_1440);
nand U8673 (N_8673,N_2634,N_1339);
xnor U8674 (N_8674,N_3167,N_3960);
or U8675 (N_8675,N_4057,N_269);
nand U8676 (N_8676,N_1344,N_4315);
and U8677 (N_8677,N_623,N_2306);
or U8678 (N_8678,N_3525,N_1950);
nor U8679 (N_8679,N_2191,N_864);
xor U8680 (N_8680,N_1550,N_52);
and U8681 (N_8681,N_3106,N_3568);
and U8682 (N_8682,N_3915,N_79);
xnor U8683 (N_8683,N_3444,N_1111);
nand U8684 (N_8684,N_4830,N_3402);
nor U8685 (N_8685,N_3874,N_1014);
nand U8686 (N_8686,N_2507,N_796);
nand U8687 (N_8687,N_2237,N_2114);
and U8688 (N_8688,N_2413,N_3693);
or U8689 (N_8689,N_4890,N_821);
or U8690 (N_8690,N_4986,N_2567);
xnor U8691 (N_8691,N_796,N_4971);
nand U8692 (N_8692,N_4003,N_3298);
xnor U8693 (N_8693,N_2447,N_2170);
nor U8694 (N_8694,N_1593,N_4061);
or U8695 (N_8695,N_4140,N_3654);
or U8696 (N_8696,N_3211,N_785);
and U8697 (N_8697,N_3224,N_4138);
nor U8698 (N_8698,N_676,N_322);
or U8699 (N_8699,N_3217,N_1148);
nand U8700 (N_8700,N_280,N_4228);
nor U8701 (N_8701,N_2613,N_3426);
xnor U8702 (N_8702,N_3014,N_3505);
nand U8703 (N_8703,N_1255,N_3529);
nand U8704 (N_8704,N_1283,N_1784);
or U8705 (N_8705,N_4487,N_629);
nand U8706 (N_8706,N_4970,N_550);
nor U8707 (N_8707,N_4493,N_4958);
xor U8708 (N_8708,N_3028,N_1645);
and U8709 (N_8709,N_2862,N_1497);
or U8710 (N_8710,N_1365,N_2145);
and U8711 (N_8711,N_262,N_3871);
or U8712 (N_8712,N_1645,N_503);
xnor U8713 (N_8713,N_4002,N_4040);
and U8714 (N_8714,N_1441,N_904);
or U8715 (N_8715,N_71,N_1977);
nand U8716 (N_8716,N_4510,N_4140);
nor U8717 (N_8717,N_3945,N_3638);
nand U8718 (N_8718,N_2592,N_1507);
or U8719 (N_8719,N_639,N_4271);
or U8720 (N_8720,N_321,N_3339);
or U8721 (N_8721,N_1226,N_1131);
or U8722 (N_8722,N_2671,N_1667);
or U8723 (N_8723,N_4816,N_3914);
nand U8724 (N_8724,N_2673,N_4435);
nor U8725 (N_8725,N_3687,N_1743);
and U8726 (N_8726,N_2852,N_2364);
and U8727 (N_8727,N_3007,N_1698);
nand U8728 (N_8728,N_2254,N_268);
and U8729 (N_8729,N_1538,N_4785);
nor U8730 (N_8730,N_334,N_4311);
and U8731 (N_8731,N_1422,N_4822);
and U8732 (N_8732,N_2774,N_2986);
nand U8733 (N_8733,N_681,N_2840);
or U8734 (N_8734,N_153,N_1661);
nor U8735 (N_8735,N_730,N_2211);
xor U8736 (N_8736,N_4056,N_3444);
nand U8737 (N_8737,N_1430,N_2400);
or U8738 (N_8738,N_568,N_1388);
nor U8739 (N_8739,N_3318,N_3752);
nor U8740 (N_8740,N_3759,N_270);
xnor U8741 (N_8741,N_952,N_1966);
nand U8742 (N_8742,N_1623,N_1197);
and U8743 (N_8743,N_50,N_4387);
nand U8744 (N_8744,N_221,N_4192);
nand U8745 (N_8745,N_4625,N_488);
xnor U8746 (N_8746,N_1835,N_831);
nand U8747 (N_8747,N_2994,N_2781);
nand U8748 (N_8748,N_971,N_2371);
nand U8749 (N_8749,N_3497,N_4044);
or U8750 (N_8750,N_2938,N_978);
nand U8751 (N_8751,N_2356,N_4946);
nand U8752 (N_8752,N_3218,N_3654);
or U8753 (N_8753,N_2892,N_3315);
and U8754 (N_8754,N_4194,N_614);
nor U8755 (N_8755,N_408,N_2027);
and U8756 (N_8756,N_2780,N_2890);
nor U8757 (N_8757,N_2352,N_2207);
or U8758 (N_8758,N_1352,N_1186);
and U8759 (N_8759,N_3864,N_3090);
nand U8760 (N_8760,N_1920,N_533);
nor U8761 (N_8761,N_791,N_2835);
or U8762 (N_8762,N_3603,N_4319);
nand U8763 (N_8763,N_41,N_2585);
xnor U8764 (N_8764,N_52,N_2647);
or U8765 (N_8765,N_1127,N_3452);
or U8766 (N_8766,N_4317,N_567);
and U8767 (N_8767,N_4312,N_1770);
nand U8768 (N_8768,N_2210,N_2666);
nor U8769 (N_8769,N_2358,N_3675);
nand U8770 (N_8770,N_1806,N_2052);
xnor U8771 (N_8771,N_2074,N_1505);
nor U8772 (N_8772,N_1139,N_4090);
and U8773 (N_8773,N_3478,N_1084);
nand U8774 (N_8774,N_2280,N_1248);
and U8775 (N_8775,N_1935,N_2947);
nand U8776 (N_8776,N_1449,N_3588);
or U8777 (N_8777,N_1606,N_255);
nor U8778 (N_8778,N_120,N_2291);
nor U8779 (N_8779,N_525,N_2887);
and U8780 (N_8780,N_4432,N_2516);
nor U8781 (N_8781,N_3088,N_761);
nor U8782 (N_8782,N_3815,N_3370);
nand U8783 (N_8783,N_3049,N_4385);
and U8784 (N_8784,N_1171,N_2823);
nor U8785 (N_8785,N_1078,N_667);
or U8786 (N_8786,N_1005,N_594);
nand U8787 (N_8787,N_2090,N_603);
nand U8788 (N_8788,N_2701,N_4727);
and U8789 (N_8789,N_2649,N_424);
nor U8790 (N_8790,N_3374,N_4229);
or U8791 (N_8791,N_783,N_311);
or U8792 (N_8792,N_1042,N_949);
xor U8793 (N_8793,N_4784,N_749);
xor U8794 (N_8794,N_695,N_3180);
nor U8795 (N_8795,N_2047,N_2224);
nor U8796 (N_8796,N_1738,N_4242);
or U8797 (N_8797,N_2475,N_2309);
nor U8798 (N_8798,N_2201,N_4287);
nor U8799 (N_8799,N_9,N_2287);
and U8800 (N_8800,N_2844,N_26);
xor U8801 (N_8801,N_835,N_930);
xnor U8802 (N_8802,N_4827,N_4942);
or U8803 (N_8803,N_2490,N_1369);
xnor U8804 (N_8804,N_995,N_4481);
xor U8805 (N_8805,N_1091,N_3148);
xnor U8806 (N_8806,N_1949,N_3306);
or U8807 (N_8807,N_2020,N_1330);
nand U8808 (N_8808,N_1703,N_3276);
nor U8809 (N_8809,N_1249,N_2879);
xor U8810 (N_8810,N_72,N_4905);
nor U8811 (N_8811,N_3890,N_213);
nand U8812 (N_8812,N_3504,N_3344);
nand U8813 (N_8813,N_4169,N_1266);
xor U8814 (N_8814,N_2955,N_1633);
and U8815 (N_8815,N_3154,N_1480);
nand U8816 (N_8816,N_1705,N_2070);
and U8817 (N_8817,N_956,N_1315);
nand U8818 (N_8818,N_2093,N_4016);
and U8819 (N_8819,N_2922,N_4583);
xor U8820 (N_8820,N_362,N_3792);
or U8821 (N_8821,N_4308,N_1450);
and U8822 (N_8822,N_3109,N_989);
nor U8823 (N_8823,N_1279,N_445);
xor U8824 (N_8824,N_4748,N_3333);
or U8825 (N_8825,N_3826,N_4751);
nand U8826 (N_8826,N_1219,N_2885);
nand U8827 (N_8827,N_1617,N_3002);
nor U8828 (N_8828,N_3186,N_923);
xnor U8829 (N_8829,N_972,N_29);
and U8830 (N_8830,N_84,N_2962);
and U8831 (N_8831,N_1324,N_1236);
nor U8832 (N_8832,N_4212,N_1778);
or U8833 (N_8833,N_614,N_217);
xor U8834 (N_8834,N_3118,N_2626);
and U8835 (N_8835,N_3499,N_1529);
or U8836 (N_8836,N_1218,N_1910);
nand U8837 (N_8837,N_4012,N_2806);
or U8838 (N_8838,N_1558,N_1922);
or U8839 (N_8839,N_4213,N_3883);
or U8840 (N_8840,N_2727,N_4473);
nand U8841 (N_8841,N_3248,N_3622);
or U8842 (N_8842,N_1110,N_3804);
or U8843 (N_8843,N_507,N_2983);
nor U8844 (N_8844,N_4844,N_2507);
nand U8845 (N_8845,N_1032,N_2251);
xor U8846 (N_8846,N_341,N_2560);
xor U8847 (N_8847,N_4931,N_4880);
nor U8848 (N_8848,N_3206,N_895);
xnor U8849 (N_8849,N_4011,N_3974);
and U8850 (N_8850,N_745,N_2286);
and U8851 (N_8851,N_1060,N_4312);
nor U8852 (N_8852,N_758,N_4809);
xnor U8853 (N_8853,N_4216,N_4011);
nand U8854 (N_8854,N_1701,N_1668);
nor U8855 (N_8855,N_3309,N_4911);
and U8856 (N_8856,N_572,N_2908);
nor U8857 (N_8857,N_1990,N_3950);
nor U8858 (N_8858,N_4329,N_3862);
or U8859 (N_8859,N_1478,N_983);
xor U8860 (N_8860,N_2092,N_637);
nor U8861 (N_8861,N_1563,N_385);
nor U8862 (N_8862,N_1888,N_545);
or U8863 (N_8863,N_1508,N_4149);
or U8864 (N_8864,N_3387,N_3974);
and U8865 (N_8865,N_1999,N_4561);
nand U8866 (N_8866,N_2096,N_1927);
and U8867 (N_8867,N_161,N_2063);
xor U8868 (N_8868,N_3555,N_4798);
or U8869 (N_8869,N_737,N_1124);
nor U8870 (N_8870,N_966,N_2666);
xor U8871 (N_8871,N_223,N_3277);
nand U8872 (N_8872,N_3593,N_2456);
or U8873 (N_8873,N_1204,N_842);
and U8874 (N_8874,N_1263,N_2110);
nor U8875 (N_8875,N_3395,N_377);
and U8876 (N_8876,N_3126,N_3359);
or U8877 (N_8877,N_3604,N_547);
nand U8878 (N_8878,N_1058,N_789);
xor U8879 (N_8879,N_3179,N_757);
and U8880 (N_8880,N_2443,N_1816);
nor U8881 (N_8881,N_2193,N_2814);
nor U8882 (N_8882,N_3197,N_1441);
xor U8883 (N_8883,N_1438,N_943);
xnor U8884 (N_8884,N_1040,N_4650);
xnor U8885 (N_8885,N_4560,N_2674);
nand U8886 (N_8886,N_372,N_1025);
nor U8887 (N_8887,N_3642,N_4628);
nor U8888 (N_8888,N_734,N_4944);
xor U8889 (N_8889,N_2484,N_215);
xor U8890 (N_8890,N_564,N_4581);
xor U8891 (N_8891,N_1127,N_903);
xnor U8892 (N_8892,N_1674,N_3963);
nor U8893 (N_8893,N_4791,N_339);
nor U8894 (N_8894,N_1236,N_973);
xor U8895 (N_8895,N_2236,N_3941);
or U8896 (N_8896,N_367,N_3902);
xnor U8897 (N_8897,N_494,N_3677);
xor U8898 (N_8898,N_3640,N_2549);
nand U8899 (N_8899,N_4370,N_3862);
and U8900 (N_8900,N_4176,N_4412);
nor U8901 (N_8901,N_2530,N_3217);
xor U8902 (N_8902,N_4577,N_4836);
or U8903 (N_8903,N_2475,N_4946);
xnor U8904 (N_8904,N_548,N_328);
nand U8905 (N_8905,N_1020,N_2959);
nand U8906 (N_8906,N_1360,N_4374);
and U8907 (N_8907,N_1461,N_1622);
nand U8908 (N_8908,N_477,N_4390);
and U8909 (N_8909,N_3474,N_1359);
nand U8910 (N_8910,N_2422,N_600);
and U8911 (N_8911,N_4134,N_4019);
and U8912 (N_8912,N_159,N_4574);
and U8913 (N_8913,N_2158,N_4368);
xnor U8914 (N_8914,N_3977,N_526);
nand U8915 (N_8915,N_2700,N_3468);
xor U8916 (N_8916,N_4124,N_3784);
nand U8917 (N_8917,N_3272,N_3875);
xnor U8918 (N_8918,N_1203,N_1031);
nand U8919 (N_8919,N_1382,N_3852);
nand U8920 (N_8920,N_2263,N_535);
xor U8921 (N_8921,N_2383,N_1334);
nand U8922 (N_8922,N_489,N_3212);
nor U8923 (N_8923,N_4250,N_579);
nand U8924 (N_8924,N_2601,N_958);
nand U8925 (N_8925,N_4498,N_1937);
and U8926 (N_8926,N_2985,N_2856);
nor U8927 (N_8927,N_3977,N_3717);
nand U8928 (N_8928,N_2718,N_122);
xor U8929 (N_8929,N_169,N_4533);
and U8930 (N_8930,N_1821,N_2000);
or U8931 (N_8931,N_3407,N_3792);
or U8932 (N_8932,N_861,N_2897);
nand U8933 (N_8933,N_2930,N_4360);
nand U8934 (N_8934,N_4074,N_1008);
or U8935 (N_8935,N_4971,N_4191);
nor U8936 (N_8936,N_4514,N_1919);
nor U8937 (N_8937,N_3512,N_1917);
and U8938 (N_8938,N_919,N_3963);
and U8939 (N_8939,N_4315,N_3542);
xor U8940 (N_8940,N_893,N_3419);
nor U8941 (N_8941,N_397,N_3045);
nand U8942 (N_8942,N_3974,N_3729);
nand U8943 (N_8943,N_3199,N_1351);
nor U8944 (N_8944,N_4982,N_2703);
nand U8945 (N_8945,N_4915,N_3286);
and U8946 (N_8946,N_1667,N_3385);
nor U8947 (N_8947,N_2831,N_3682);
nand U8948 (N_8948,N_2970,N_2803);
nor U8949 (N_8949,N_2016,N_1170);
and U8950 (N_8950,N_1416,N_1148);
xor U8951 (N_8951,N_2355,N_821);
and U8952 (N_8952,N_2910,N_4205);
xnor U8953 (N_8953,N_168,N_2458);
nand U8954 (N_8954,N_3400,N_2125);
nor U8955 (N_8955,N_4868,N_4033);
and U8956 (N_8956,N_1051,N_3439);
nor U8957 (N_8957,N_1237,N_3417);
xor U8958 (N_8958,N_1792,N_1023);
xnor U8959 (N_8959,N_2565,N_1553);
xnor U8960 (N_8960,N_984,N_2016);
xnor U8961 (N_8961,N_79,N_2898);
xnor U8962 (N_8962,N_4573,N_146);
or U8963 (N_8963,N_2365,N_150);
and U8964 (N_8964,N_4721,N_902);
xnor U8965 (N_8965,N_2932,N_1449);
nor U8966 (N_8966,N_1589,N_3491);
xnor U8967 (N_8967,N_1675,N_3084);
nor U8968 (N_8968,N_4749,N_4318);
xnor U8969 (N_8969,N_3164,N_1317);
xnor U8970 (N_8970,N_4809,N_1956);
nand U8971 (N_8971,N_3286,N_4497);
or U8972 (N_8972,N_2547,N_2083);
and U8973 (N_8973,N_3024,N_4316);
and U8974 (N_8974,N_4419,N_2076);
nor U8975 (N_8975,N_1340,N_4508);
xnor U8976 (N_8976,N_3192,N_2907);
or U8977 (N_8977,N_1741,N_2020);
nor U8978 (N_8978,N_68,N_4258);
nor U8979 (N_8979,N_1857,N_3956);
nand U8980 (N_8980,N_3138,N_1734);
nand U8981 (N_8981,N_2419,N_600);
nor U8982 (N_8982,N_4336,N_2547);
and U8983 (N_8983,N_723,N_3453);
nand U8984 (N_8984,N_409,N_116);
nand U8985 (N_8985,N_4857,N_1970);
or U8986 (N_8986,N_4694,N_833);
and U8987 (N_8987,N_4873,N_2246);
or U8988 (N_8988,N_1845,N_280);
or U8989 (N_8989,N_1263,N_2149);
nand U8990 (N_8990,N_2786,N_3421);
or U8991 (N_8991,N_4652,N_2665);
xnor U8992 (N_8992,N_4957,N_4682);
nor U8993 (N_8993,N_1354,N_4462);
nand U8994 (N_8994,N_3248,N_3484);
nor U8995 (N_8995,N_3203,N_1062);
or U8996 (N_8996,N_3054,N_3752);
nand U8997 (N_8997,N_2156,N_2822);
xnor U8998 (N_8998,N_2225,N_2612);
xor U8999 (N_8999,N_1210,N_4034);
or U9000 (N_9000,N_3566,N_1300);
nand U9001 (N_9001,N_3783,N_1252);
nand U9002 (N_9002,N_1750,N_2175);
xor U9003 (N_9003,N_4946,N_2648);
nand U9004 (N_9004,N_1193,N_2553);
nand U9005 (N_9005,N_23,N_1772);
and U9006 (N_9006,N_3446,N_2801);
nand U9007 (N_9007,N_4243,N_522);
xor U9008 (N_9008,N_1358,N_4551);
or U9009 (N_9009,N_1589,N_884);
nor U9010 (N_9010,N_4449,N_331);
or U9011 (N_9011,N_3983,N_314);
and U9012 (N_9012,N_696,N_4208);
nand U9013 (N_9013,N_2638,N_4028);
nor U9014 (N_9014,N_4605,N_3009);
xor U9015 (N_9015,N_291,N_3402);
and U9016 (N_9016,N_1102,N_4909);
nand U9017 (N_9017,N_1535,N_4244);
nand U9018 (N_9018,N_4766,N_685);
and U9019 (N_9019,N_1162,N_3686);
nand U9020 (N_9020,N_3100,N_4712);
xnor U9021 (N_9021,N_2035,N_2187);
or U9022 (N_9022,N_4519,N_3259);
xnor U9023 (N_9023,N_1704,N_3798);
nand U9024 (N_9024,N_2125,N_1335);
nand U9025 (N_9025,N_3638,N_4348);
and U9026 (N_9026,N_4270,N_3213);
nand U9027 (N_9027,N_1437,N_1970);
or U9028 (N_9028,N_2692,N_4745);
xnor U9029 (N_9029,N_3823,N_3517);
xor U9030 (N_9030,N_2562,N_4960);
nor U9031 (N_9031,N_2527,N_1451);
xor U9032 (N_9032,N_4788,N_1164);
xnor U9033 (N_9033,N_3078,N_1979);
and U9034 (N_9034,N_4541,N_4955);
nand U9035 (N_9035,N_3463,N_136);
or U9036 (N_9036,N_4212,N_610);
nor U9037 (N_9037,N_1392,N_16);
or U9038 (N_9038,N_4711,N_1349);
xnor U9039 (N_9039,N_4568,N_4911);
nand U9040 (N_9040,N_3174,N_3709);
xor U9041 (N_9041,N_2577,N_3916);
xor U9042 (N_9042,N_2753,N_2266);
nand U9043 (N_9043,N_2628,N_3932);
xor U9044 (N_9044,N_830,N_3161);
nand U9045 (N_9045,N_4375,N_1230);
nor U9046 (N_9046,N_591,N_2148);
nor U9047 (N_9047,N_2677,N_4022);
nor U9048 (N_9048,N_4850,N_1153);
xor U9049 (N_9049,N_12,N_1525);
nand U9050 (N_9050,N_1454,N_3927);
or U9051 (N_9051,N_2989,N_1669);
nand U9052 (N_9052,N_3855,N_4046);
or U9053 (N_9053,N_4910,N_164);
nor U9054 (N_9054,N_3643,N_1860);
xnor U9055 (N_9055,N_4652,N_701);
nand U9056 (N_9056,N_211,N_4132);
nor U9057 (N_9057,N_2511,N_2686);
nand U9058 (N_9058,N_2237,N_4603);
and U9059 (N_9059,N_2757,N_368);
nor U9060 (N_9060,N_743,N_396);
nand U9061 (N_9061,N_3873,N_3041);
and U9062 (N_9062,N_4672,N_1285);
nor U9063 (N_9063,N_2347,N_3434);
nand U9064 (N_9064,N_772,N_3230);
nor U9065 (N_9065,N_2106,N_1907);
xor U9066 (N_9066,N_4179,N_3905);
nand U9067 (N_9067,N_1563,N_1542);
or U9068 (N_9068,N_1046,N_4092);
nor U9069 (N_9069,N_73,N_1558);
nor U9070 (N_9070,N_1911,N_2526);
xor U9071 (N_9071,N_3343,N_2552);
nor U9072 (N_9072,N_256,N_2689);
nand U9073 (N_9073,N_2708,N_1474);
xor U9074 (N_9074,N_610,N_1509);
xor U9075 (N_9075,N_3692,N_4529);
or U9076 (N_9076,N_1630,N_2765);
xor U9077 (N_9077,N_4344,N_3116);
nor U9078 (N_9078,N_4702,N_2911);
and U9079 (N_9079,N_1619,N_288);
nand U9080 (N_9080,N_1015,N_2821);
xor U9081 (N_9081,N_3037,N_2896);
and U9082 (N_9082,N_2843,N_597);
nor U9083 (N_9083,N_2251,N_2740);
or U9084 (N_9084,N_2149,N_70);
nor U9085 (N_9085,N_200,N_4833);
and U9086 (N_9086,N_1091,N_778);
nor U9087 (N_9087,N_3006,N_1968);
xor U9088 (N_9088,N_1804,N_4988);
and U9089 (N_9089,N_4377,N_462);
xor U9090 (N_9090,N_175,N_2211);
nand U9091 (N_9091,N_1308,N_2083);
nor U9092 (N_9092,N_363,N_934);
or U9093 (N_9093,N_2199,N_3064);
nor U9094 (N_9094,N_704,N_1922);
xnor U9095 (N_9095,N_672,N_604);
and U9096 (N_9096,N_464,N_902);
xor U9097 (N_9097,N_4337,N_34);
or U9098 (N_9098,N_3582,N_2798);
or U9099 (N_9099,N_3518,N_1839);
xor U9100 (N_9100,N_200,N_4651);
nor U9101 (N_9101,N_3332,N_4893);
xor U9102 (N_9102,N_4027,N_4733);
or U9103 (N_9103,N_177,N_3749);
or U9104 (N_9104,N_1529,N_2698);
nand U9105 (N_9105,N_451,N_1380);
or U9106 (N_9106,N_2199,N_2514);
and U9107 (N_9107,N_2540,N_2601);
and U9108 (N_9108,N_986,N_606);
or U9109 (N_9109,N_818,N_4178);
xor U9110 (N_9110,N_4998,N_4746);
xnor U9111 (N_9111,N_1363,N_2180);
nor U9112 (N_9112,N_3823,N_419);
and U9113 (N_9113,N_2540,N_4289);
and U9114 (N_9114,N_2855,N_541);
nor U9115 (N_9115,N_4834,N_3954);
nand U9116 (N_9116,N_4535,N_4433);
and U9117 (N_9117,N_2259,N_666);
and U9118 (N_9118,N_2290,N_4837);
or U9119 (N_9119,N_3796,N_4024);
and U9120 (N_9120,N_4225,N_2763);
or U9121 (N_9121,N_1442,N_3093);
or U9122 (N_9122,N_1384,N_1301);
nand U9123 (N_9123,N_4324,N_3756);
and U9124 (N_9124,N_1186,N_2760);
xor U9125 (N_9125,N_4271,N_2423);
xor U9126 (N_9126,N_3263,N_1343);
xor U9127 (N_9127,N_4712,N_463);
nor U9128 (N_9128,N_537,N_1612);
nand U9129 (N_9129,N_3900,N_2565);
and U9130 (N_9130,N_4618,N_3819);
and U9131 (N_9131,N_2775,N_551);
nor U9132 (N_9132,N_2255,N_1056);
xnor U9133 (N_9133,N_2531,N_650);
nand U9134 (N_9134,N_4573,N_4082);
xor U9135 (N_9135,N_4094,N_3673);
nand U9136 (N_9136,N_1996,N_1969);
nand U9137 (N_9137,N_3586,N_4561);
nand U9138 (N_9138,N_874,N_4630);
nand U9139 (N_9139,N_3006,N_3458);
or U9140 (N_9140,N_414,N_2904);
nor U9141 (N_9141,N_4082,N_4306);
nor U9142 (N_9142,N_1379,N_897);
xor U9143 (N_9143,N_4348,N_1036);
or U9144 (N_9144,N_437,N_1776);
xnor U9145 (N_9145,N_3647,N_3075);
and U9146 (N_9146,N_3987,N_3607);
or U9147 (N_9147,N_1292,N_3957);
or U9148 (N_9148,N_2437,N_4457);
nand U9149 (N_9149,N_161,N_265);
or U9150 (N_9150,N_4008,N_2690);
xor U9151 (N_9151,N_19,N_4122);
nand U9152 (N_9152,N_4768,N_3993);
and U9153 (N_9153,N_760,N_2398);
nand U9154 (N_9154,N_4825,N_3866);
or U9155 (N_9155,N_4157,N_1245);
or U9156 (N_9156,N_1143,N_2592);
xnor U9157 (N_9157,N_1642,N_4683);
nor U9158 (N_9158,N_4105,N_3539);
nor U9159 (N_9159,N_3905,N_1953);
and U9160 (N_9160,N_1285,N_4928);
xnor U9161 (N_9161,N_232,N_4039);
nand U9162 (N_9162,N_1892,N_4830);
nor U9163 (N_9163,N_1489,N_2313);
and U9164 (N_9164,N_2974,N_2031);
or U9165 (N_9165,N_1314,N_2120);
xnor U9166 (N_9166,N_2875,N_2472);
or U9167 (N_9167,N_446,N_2589);
or U9168 (N_9168,N_3594,N_3024);
and U9169 (N_9169,N_1370,N_475);
nand U9170 (N_9170,N_1310,N_2727);
nor U9171 (N_9171,N_717,N_3771);
xnor U9172 (N_9172,N_4376,N_3246);
xor U9173 (N_9173,N_854,N_3712);
nand U9174 (N_9174,N_3462,N_2197);
or U9175 (N_9175,N_1082,N_370);
nand U9176 (N_9176,N_4657,N_1063);
xor U9177 (N_9177,N_1386,N_4978);
nand U9178 (N_9178,N_2213,N_1838);
or U9179 (N_9179,N_4696,N_4065);
nand U9180 (N_9180,N_3820,N_3479);
or U9181 (N_9181,N_3839,N_4100);
or U9182 (N_9182,N_1136,N_4482);
nand U9183 (N_9183,N_270,N_156);
nor U9184 (N_9184,N_4330,N_697);
or U9185 (N_9185,N_650,N_873);
xnor U9186 (N_9186,N_564,N_4657);
nor U9187 (N_9187,N_4493,N_4751);
nand U9188 (N_9188,N_2507,N_495);
xnor U9189 (N_9189,N_2893,N_2442);
and U9190 (N_9190,N_4366,N_1935);
and U9191 (N_9191,N_4037,N_1999);
and U9192 (N_9192,N_3055,N_1172);
and U9193 (N_9193,N_2041,N_3638);
xor U9194 (N_9194,N_4508,N_368);
nor U9195 (N_9195,N_4026,N_1091);
or U9196 (N_9196,N_2122,N_4871);
xnor U9197 (N_9197,N_2283,N_4186);
nand U9198 (N_9198,N_2155,N_4674);
nor U9199 (N_9199,N_1434,N_3973);
nor U9200 (N_9200,N_1324,N_3332);
and U9201 (N_9201,N_2320,N_2769);
or U9202 (N_9202,N_4424,N_2103);
nor U9203 (N_9203,N_968,N_1965);
nor U9204 (N_9204,N_488,N_282);
xnor U9205 (N_9205,N_4503,N_1249);
nor U9206 (N_9206,N_4767,N_4315);
or U9207 (N_9207,N_3968,N_2283);
nand U9208 (N_9208,N_3542,N_4467);
and U9209 (N_9209,N_631,N_2116);
and U9210 (N_9210,N_4928,N_4217);
xor U9211 (N_9211,N_1164,N_52);
and U9212 (N_9212,N_2474,N_2895);
nor U9213 (N_9213,N_2601,N_985);
or U9214 (N_9214,N_2450,N_700);
or U9215 (N_9215,N_3917,N_4025);
and U9216 (N_9216,N_884,N_3234);
and U9217 (N_9217,N_3855,N_3098);
xor U9218 (N_9218,N_2816,N_2877);
or U9219 (N_9219,N_1335,N_2409);
and U9220 (N_9220,N_4280,N_1153);
and U9221 (N_9221,N_4715,N_724);
nor U9222 (N_9222,N_986,N_1448);
xnor U9223 (N_9223,N_3041,N_4487);
and U9224 (N_9224,N_1950,N_2869);
nor U9225 (N_9225,N_3815,N_2639);
nand U9226 (N_9226,N_4706,N_3621);
nor U9227 (N_9227,N_1408,N_1986);
and U9228 (N_9228,N_49,N_2417);
and U9229 (N_9229,N_3567,N_3103);
and U9230 (N_9230,N_172,N_3769);
xor U9231 (N_9231,N_2941,N_835);
or U9232 (N_9232,N_302,N_1948);
nand U9233 (N_9233,N_2955,N_492);
or U9234 (N_9234,N_739,N_1263);
nor U9235 (N_9235,N_1951,N_3238);
nand U9236 (N_9236,N_1560,N_2610);
or U9237 (N_9237,N_3622,N_3334);
and U9238 (N_9238,N_3477,N_3022);
or U9239 (N_9239,N_3189,N_1380);
xor U9240 (N_9240,N_2980,N_3275);
or U9241 (N_9241,N_4419,N_2521);
nor U9242 (N_9242,N_4527,N_998);
and U9243 (N_9243,N_3748,N_4708);
and U9244 (N_9244,N_3801,N_1697);
and U9245 (N_9245,N_2874,N_3593);
xnor U9246 (N_9246,N_4384,N_331);
nand U9247 (N_9247,N_940,N_3621);
nand U9248 (N_9248,N_1931,N_1051);
and U9249 (N_9249,N_3623,N_4626);
or U9250 (N_9250,N_3588,N_4770);
nand U9251 (N_9251,N_4822,N_3821);
and U9252 (N_9252,N_3690,N_3742);
xor U9253 (N_9253,N_1181,N_3840);
nand U9254 (N_9254,N_252,N_3281);
nand U9255 (N_9255,N_2320,N_1956);
or U9256 (N_9256,N_2869,N_3524);
nor U9257 (N_9257,N_1957,N_2113);
or U9258 (N_9258,N_310,N_1253);
and U9259 (N_9259,N_2926,N_1229);
or U9260 (N_9260,N_4188,N_2520);
and U9261 (N_9261,N_1952,N_2417);
xor U9262 (N_9262,N_4235,N_3671);
and U9263 (N_9263,N_4992,N_2247);
nor U9264 (N_9264,N_3109,N_915);
nand U9265 (N_9265,N_623,N_4275);
and U9266 (N_9266,N_2323,N_3257);
nand U9267 (N_9267,N_4595,N_3964);
or U9268 (N_9268,N_2171,N_71);
nor U9269 (N_9269,N_3223,N_4263);
xnor U9270 (N_9270,N_197,N_1256);
nand U9271 (N_9271,N_4976,N_4310);
nor U9272 (N_9272,N_1190,N_3813);
and U9273 (N_9273,N_2377,N_1716);
nand U9274 (N_9274,N_2064,N_2214);
xor U9275 (N_9275,N_2705,N_4231);
xnor U9276 (N_9276,N_812,N_3760);
xor U9277 (N_9277,N_4213,N_3544);
nand U9278 (N_9278,N_2539,N_1835);
nand U9279 (N_9279,N_415,N_2930);
nor U9280 (N_9280,N_3199,N_3205);
nor U9281 (N_9281,N_2798,N_2767);
and U9282 (N_9282,N_3307,N_1983);
nand U9283 (N_9283,N_4566,N_3812);
nand U9284 (N_9284,N_2558,N_2188);
and U9285 (N_9285,N_4663,N_562);
xnor U9286 (N_9286,N_373,N_4123);
nand U9287 (N_9287,N_1416,N_1935);
nor U9288 (N_9288,N_1264,N_4785);
xnor U9289 (N_9289,N_2568,N_2808);
or U9290 (N_9290,N_3564,N_4896);
nand U9291 (N_9291,N_4893,N_3685);
nor U9292 (N_9292,N_1237,N_4982);
nor U9293 (N_9293,N_4824,N_1227);
nor U9294 (N_9294,N_4550,N_960);
nor U9295 (N_9295,N_1832,N_2435);
nor U9296 (N_9296,N_4284,N_913);
or U9297 (N_9297,N_2596,N_1942);
xnor U9298 (N_9298,N_1294,N_1683);
nor U9299 (N_9299,N_4546,N_2958);
nor U9300 (N_9300,N_554,N_377);
xor U9301 (N_9301,N_2690,N_3799);
and U9302 (N_9302,N_3809,N_3883);
nand U9303 (N_9303,N_3577,N_1990);
or U9304 (N_9304,N_1467,N_3591);
xor U9305 (N_9305,N_4409,N_1838);
nand U9306 (N_9306,N_3358,N_3004);
or U9307 (N_9307,N_3131,N_4048);
nand U9308 (N_9308,N_888,N_3360);
xor U9309 (N_9309,N_3320,N_3010);
xor U9310 (N_9310,N_3344,N_3345);
nand U9311 (N_9311,N_2131,N_1053);
or U9312 (N_9312,N_3991,N_1439);
and U9313 (N_9313,N_1976,N_4653);
xor U9314 (N_9314,N_3200,N_3766);
xnor U9315 (N_9315,N_1598,N_4835);
nor U9316 (N_9316,N_1079,N_765);
nand U9317 (N_9317,N_3395,N_1047);
nand U9318 (N_9318,N_4877,N_2293);
nand U9319 (N_9319,N_1500,N_2865);
xnor U9320 (N_9320,N_1598,N_2735);
or U9321 (N_9321,N_2661,N_1948);
nand U9322 (N_9322,N_2346,N_443);
and U9323 (N_9323,N_4696,N_1516);
and U9324 (N_9324,N_4844,N_2701);
or U9325 (N_9325,N_1829,N_3787);
xor U9326 (N_9326,N_4307,N_4100);
nand U9327 (N_9327,N_452,N_4297);
or U9328 (N_9328,N_963,N_789);
xor U9329 (N_9329,N_0,N_1956);
xnor U9330 (N_9330,N_1289,N_786);
nand U9331 (N_9331,N_323,N_2960);
or U9332 (N_9332,N_4274,N_4804);
and U9333 (N_9333,N_1136,N_3779);
or U9334 (N_9334,N_3766,N_3195);
nor U9335 (N_9335,N_1059,N_3826);
or U9336 (N_9336,N_4174,N_1147);
or U9337 (N_9337,N_2354,N_528);
or U9338 (N_9338,N_918,N_702);
or U9339 (N_9339,N_28,N_2790);
xor U9340 (N_9340,N_2367,N_4218);
nor U9341 (N_9341,N_865,N_1524);
and U9342 (N_9342,N_177,N_4970);
nor U9343 (N_9343,N_439,N_2555);
nor U9344 (N_9344,N_1192,N_4341);
and U9345 (N_9345,N_2150,N_590);
or U9346 (N_9346,N_561,N_531);
nor U9347 (N_9347,N_2844,N_2900);
or U9348 (N_9348,N_3426,N_1725);
xor U9349 (N_9349,N_2207,N_2266);
nand U9350 (N_9350,N_117,N_2848);
nor U9351 (N_9351,N_2895,N_651);
or U9352 (N_9352,N_612,N_2083);
or U9353 (N_9353,N_3614,N_2334);
nor U9354 (N_9354,N_2810,N_3774);
or U9355 (N_9355,N_1346,N_63);
nand U9356 (N_9356,N_1928,N_4608);
nand U9357 (N_9357,N_1517,N_2781);
and U9358 (N_9358,N_1233,N_1072);
and U9359 (N_9359,N_884,N_2121);
nand U9360 (N_9360,N_1309,N_4862);
xnor U9361 (N_9361,N_1549,N_3330);
or U9362 (N_9362,N_2729,N_3204);
or U9363 (N_9363,N_3298,N_3065);
nor U9364 (N_9364,N_2799,N_2880);
xor U9365 (N_9365,N_999,N_1191);
nand U9366 (N_9366,N_951,N_4363);
or U9367 (N_9367,N_1657,N_2721);
nor U9368 (N_9368,N_2378,N_2839);
and U9369 (N_9369,N_3828,N_237);
nor U9370 (N_9370,N_1716,N_3965);
and U9371 (N_9371,N_2455,N_3356);
or U9372 (N_9372,N_3577,N_3155);
and U9373 (N_9373,N_2220,N_4484);
nand U9374 (N_9374,N_4826,N_2416);
or U9375 (N_9375,N_2012,N_4168);
xor U9376 (N_9376,N_707,N_4138);
nand U9377 (N_9377,N_4444,N_2229);
xnor U9378 (N_9378,N_3534,N_2250);
nand U9379 (N_9379,N_1815,N_3077);
xnor U9380 (N_9380,N_3857,N_3728);
or U9381 (N_9381,N_2457,N_1745);
or U9382 (N_9382,N_2820,N_1564);
nor U9383 (N_9383,N_3647,N_4373);
nor U9384 (N_9384,N_4887,N_4551);
or U9385 (N_9385,N_807,N_108);
nor U9386 (N_9386,N_3471,N_2013);
xor U9387 (N_9387,N_4173,N_619);
nand U9388 (N_9388,N_1971,N_2025);
nor U9389 (N_9389,N_3743,N_4910);
and U9390 (N_9390,N_3657,N_4410);
or U9391 (N_9391,N_3486,N_1513);
nor U9392 (N_9392,N_2475,N_4020);
or U9393 (N_9393,N_2979,N_1086);
nand U9394 (N_9394,N_3587,N_4870);
or U9395 (N_9395,N_614,N_2356);
nand U9396 (N_9396,N_33,N_4629);
and U9397 (N_9397,N_1857,N_2661);
or U9398 (N_9398,N_3498,N_2359);
nand U9399 (N_9399,N_2707,N_3346);
nor U9400 (N_9400,N_2314,N_411);
nand U9401 (N_9401,N_685,N_460);
or U9402 (N_9402,N_1841,N_2309);
nand U9403 (N_9403,N_4727,N_67);
nand U9404 (N_9404,N_2537,N_3143);
and U9405 (N_9405,N_213,N_722);
xnor U9406 (N_9406,N_3084,N_663);
nand U9407 (N_9407,N_3620,N_459);
or U9408 (N_9408,N_3425,N_1197);
nand U9409 (N_9409,N_3675,N_288);
nor U9410 (N_9410,N_3459,N_2846);
xor U9411 (N_9411,N_1279,N_317);
or U9412 (N_9412,N_1848,N_1594);
nor U9413 (N_9413,N_2207,N_3397);
or U9414 (N_9414,N_1242,N_2424);
nor U9415 (N_9415,N_1863,N_4826);
and U9416 (N_9416,N_2390,N_4374);
xor U9417 (N_9417,N_3110,N_3042);
nor U9418 (N_9418,N_4599,N_851);
and U9419 (N_9419,N_4151,N_3421);
nor U9420 (N_9420,N_1285,N_927);
or U9421 (N_9421,N_3630,N_4364);
or U9422 (N_9422,N_2139,N_1992);
or U9423 (N_9423,N_112,N_1758);
nand U9424 (N_9424,N_4023,N_2277);
or U9425 (N_9425,N_4992,N_2263);
nand U9426 (N_9426,N_4795,N_2334);
xor U9427 (N_9427,N_2670,N_2089);
and U9428 (N_9428,N_3835,N_519);
xor U9429 (N_9429,N_4911,N_1703);
nand U9430 (N_9430,N_3480,N_2231);
xnor U9431 (N_9431,N_747,N_2623);
nand U9432 (N_9432,N_2739,N_2709);
and U9433 (N_9433,N_2863,N_1679);
or U9434 (N_9434,N_2553,N_931);
nand U9435 (N_9435,N_3121,N_1270);
and U9436 (N_9436,N_2003,N_1091);
and U9437 (N_9437,N_3407,N_957);
and U9438 (N_9438,N_2767,N_1875);
nor U9439 (N_9439,N_3575,N_924);
or U9440 (N_9440,N_394,N_1241);
xnor U9441 (N_9441,N_904,N_2958);
and U9442 (N_9442,N_112,N_1843);
or U9443 (N_9443,N_1285,N_4905);
nand U9444 (N_9444,N_3855,N_2642);
nor U9445 (N_9445,N_475,N_1210);
xnor U9446 (N_9446,N_28,N_1146);
nand U9447 (N_9447,N_4142,N_2497);
nor U9448 (N_9448,N_1709,N_3288);
nor U9449 (N_9449,N_380,N_502);
xor U9450 (N_9450,N_3698,N_3228);
xnor U9451 (N_9451,N_1495,N_175);
nor U9452 (N_9452,N_4122,N_4958);
or U9453 (N_9453,N_1644,N_2786);
nand U9454 (N_9454,N_1798,N_1643);
xnor U9455 (N_9455,N_2285,N_4662);
or U9456 (N_9456,N_1808,N_1855);
xor U9457 (N_9457,N_876,N_1131);
nand U9458 (N_9458,N_4419,N_2730);
nand U9459 (N_9459,N_1867,N_4407);
xnor U9460 (N_9460,N_1022,N_4825);
and U9461 (N_9461,N_4924,N_75);
nor U9462 (N_9462,N_2000,N_1387);
or U9463 (N_9463,N_1568,N_928);
or U9464 (N_9464,N_2882,N_1706);
nand U9465 (N_9465,N_1924,N_1414);
xnor U9466 (N_9466,N_921,N_1743);
nand U9467 (N_9467,N_1386,N_2640);
or U9468 (N_9468,N_4923,N_4621);
and U9469 (N_9469,N_520,N_835);
xnor U9470 (N_9470,N_4728,N_2967);
nand U9471 (N_9471,N_3931,N_2905);
nor U9472 (N_9472,N_3859,N_2535);
nand U9473 (N_9473,N_4181,N_469);
nor U9474 (N_9474,N_1310,N_175);
and U9475 (N_9475,N_713,N_4184);
or U9476 (N_9476,N_1363,N_4143);
and U9477 (N_9477,N_3489,N_1468);
nand U9478 (N_9478,N_4891,N_3974);
nand U9479 (N_9479,N_1548,N_955);
nand U9480 (N_9480,N_2296,N_2756);
xor U9481 (N_9481,N_3976,N_4076);
or U9482 (N_9482,N_1412,N_1734);
and U9483 (N_9483,N_2415,N_4703);
or U9484 (N_9484,N_369,N_618);
or U9485 (N_9485,N_52,N_598);
nand U9486 (N_9486,N_1709,N_2993);
xnor U9487 (N_9487,N_644,N_1901);
xnor U9488 (N_9488,N_446,N_3297);
nor U9489 (N_9489,N_1874,N_1296);
or U9490 (N_9490,N_2337,N_3129);
nor U9491 (N_9491,N_3285,N_4968);
and U9492 (N_9492,N_769,N_1696);
xor U9493 (N_9493,N_4829,N_1668);
nand U9494 (N_9494,N_1570,N_4734);
and U9495 (N_9495,N_2761,N_1217);
xnor U9496 (N_9496,N_4703,N_4749);
xor U9497 (N_9497,N_1856,N_412);
nor U9498 (N_9498,N_2327,N_1947);
and U9499 (N_9499,N_4952,N_1751);
or U9500 (N_9500,N_1748,N_587);
and U9501 (N_9501,N_3473,N_3646);
and U9502 (N_9502,N_4748,N_1113);
nor U9503 (N_9503,N_1159,N_342);
nor U9504 (N_9504,N_2072,N_1587);
nor U9505 (N_9505,N_2480,N_1630);
nor U9506 (N_9506,N_3950,N_2544);
and U9507 (N_9507,N_4621,N_2783);
nand U9508 (N_9508,N_2589,N_4740);
nand U9509 (N_9509,N_1507,N_3438);
nor U9510 (N_9510,N_1011,N_1626);
and U9511 (N_9511,N_4435,N_4301);
xor U9512 (N_9512,N_2327,N_4106);
nand U9513 (N_9513,N_4576,N_3197);
and U9514 (N_9514,N_4194,N_1597);
nand U9515 (N_9515,N_3981,N_1644);
xnor U9516 (N_9516,N_4454,N_4872);
or U9517 (N_9517,N_3288,N_1245);
and U9518 (N_9518,N_4773,N_3915);
nor U9519 (N_9519,N_4197,N_2093);
nand U9520 (N_9520,N_937,N_2723);
nor U9521 (N_9521,N_3761,N_774);
or U9522 (N_9522,N_2651,N_4231);
or U9523 (N_9523,N_2083,N_4252);
and U9524 (N_9524,N_396,N_4060);
or U9525 (N_9525,N_2248,N_917);
nand U9526 (N_9526,N_1494,N_268);
and U9527 (N_9527,N_3409,N_2338);
xor U9528 (N_9528,N_2101,N_1949);
nor U9529 (N_9529,N_1434,N_4211);
or U9530 (N_9530,N_2828,N_2197);
and U9531 (N_9531,N_1587,N_616);
nand U9532 (N_9532,N_1690,N_4147);
and U9533 (N_9533,N_1878,N_3581);
nor U9534 (N_9534,N_3573,N_3706);
and U9535 (N_9535,N_4326,N_2546);
and U9536 (N_9536,N_248,N_2481);
xnor U9537 (N_9537,N_1876,N_825);
nand U9538 (N_9538,N_3179,N_2762);
and U9539 (N_9539,N_1586,N_4084);
xnor U9540 (N_9540,N_77,N_3604);
and U9541 (N_9541,N_3644,N_3331);
and U9542 (N_9542,N_2614,N_1105);
nor U9543 (N_9543,N_4579,N_1876);
nor U9544 (N_9544,N_3406,N_4841);
and U9545 (N_9545,N_859,N_1373);
and U9546 (N_9546,N_2957,N_3651);
or U9547 (N_9547,N_759,N_4319);
or U9548 (N_9548,N_2206,N_4400);
nand U9549 (N_9549,N_2267,N_2482);
nor U9550 (N_9550,N_2766,N_247);
or U9551 (N_9551,N_2649,N_3807);
and U9552 (N_9552,N_2836,N_1142);
xnor U9553 (N_9553,N_938,N_4959);
and U9554 (N_9554,N_520,N_3378);
or U9555 (N_9555,N_4384,N_3513);
or U9556 (N_9556,N_359,N_3116);
and U9557 (N_9557,N_4419,N_456);
nor U9558 (N_9558,N_3164,N_4869);
xnor U9559 (N_9559,N_2182,N_964);
nand U9560 (N_9560,N_604,N_592);
or U9561 (N_9561,N_2974,N_2969);
xnor U9562 (N_9562,N_3232,N_3515);
xnor U9563 (N_9563,N_330,N_719);
and U9564 (N_9564,N_936,N_1072);
nor U9565 (N_9565,N_2575,N_1843);
nor U9566 (N_9566,N_4118,N_177);
and U9567 (N_9567,N_3090,N_2130);
and U9568 (N_9568,N_1926,N_494);
or U9569 (N_9569,N_3958,N_2406);
nand U9570 (N_9570,N_4106,N_745);
nand U9571 (N_9571,N_654,N_1195);
xnor U9572 (N_9572,N_1336,N_3568);
nand U9573 (N_9573,N_2177,N_2382);
or U9574 (N_9574,N_923,N_912);
xor U9575 (N_9575,N_1439,N_425);
and U9576 (N_9576,N_2056,N_4749);
or U9577 (N_9577,N_3963,N_2644);
nor U9578 (N_9578,N_577,N_1349);
and U9579 (N_9579,N_4071,N_4512);
and U9580 (N_9580,N_2807,N_170);
xor U9581 (N_9581,N_866,N_2543);
and U9582 (N_9582,N_3623,N_4734);
or U9583 (N_9583,N_109,N_2381);
and U9584 (N_9584,N_4596,N_2889);
and U9585 (N_9585,N_3304,N_2593);
and U9586 (N_9586,N_103,N_1472);
nand U9587 (N_9587,N_4654,N_3244);
nor U9588 (N_9588,N_3266,N_2244);
and U9589 (N_9589,N_4555,N_647);
xor U9590 (N_9590,N_3654,N_284);
and U9591 (N_9591,N_4665,N_2148);
and U9592 (N_9592,N_4944,N_2531);
nor U9593 (N_9593,N_1079,N_3569);
nand U9594 (N_9594,N_567,N_1669);
nor U9595 (N_9595,N_1581,N_3377);
nand U9596 (N_9596,N_987,N_1311);
xnor U9597 (N_9597,N_678,N_4482);
and U9598 (N_9598,N_1598,N_1447);
or U9599 (N_9599,N_3112,N_4276);
or U9600 (N_9600,N_3132,N_838);
and U9601 (N_9601,N_373,N_4143);
or U9602 (N_9602,N_995,N_3839);
or U9603 (N_9603,N_1603,N_1290);
nand U9604 (N_9604,N_2711,N_3940);
and U9605 (N_9605,N_3757,N_594);
nand U9606 (N_9606,N_2878,N_4054);
or U9607 (N_9607,N_4616,N_488);
and U9608 (N_9608,N_3938,N_300);
or U9609 (N_9609,N_3738,N_2431);
xor U9610 (N_9610,N_2634,N_2809);
xor U9611 (N_9611,N_2420,N_332);
and U9612 (N_9612,N_1955,N_202);
nor U9613 (N_9613,N_3458,N_338);
nor U9614 (N_9614,N_2250,N_1417);
or U9615 (N_9615,N_2178,N_3394);
and U9616 (N_9616,N_1828,N_1426);
or U9617 (N_9617,N_1493,N_4842);
xor U9618 (N_9618,N_2762,N_4041);
nand U9619 (N_9619,N_2691,N_314);
nor U9620 (N_9620,N_4986,N_2835);
and U9621 (N_9621,N_3491,N_3990);
or U9622 (N_9622,N_265,N_4228);
or U9623 (N_9623,N_1558,N_2625);
nor U9624 (N_9624,N_3944,N_4987);
nand U9625 (N_9625,N_1074,N_4514);
xnor U9626 (N_9626,N_270,N_125);
nor U9627 (N_9627,N_989,N_617);
and U9628 (N_9628,N_4200,N_1261);
or U9629 (N_9629,N_1494,N_4203);
and U9630 (N_9630,N_663,N_2634);
and U9631 (N_9631,N_4863,N_66);
or U9632 (N_9632,N_2079,N_3645);
nand U9633 (N_9633,N_1487,N_3783);
xor U9634 (N_9634,N_1206,N_2956);
or U9635 (N_9635,N_3264,N_542);
nor U9636 (N_9636,N_2181,N_4425);
nor U9637 (N_9637,N_970,N_598);
and U9638 (N_9638,N_3039,N_4231);
and U9639 (N_9639,N_4901,N_4714);
xor U9640 (N_9640,N_4811,N_3790);
nand U9641 (N_9641,N_2028,N_718);
xor U9642 (N_9642,N_691,N_2881);
or U9643 (N_9643,N_1731,N_4647);
xnor U9644 (N_9644,N_4406,N_297);
and U9645 (N_9645,N_2657,N_1043);
nand U9646 (N_9646,N_4231,N_4654);
nand U9647 (N_9647,N_1041,N_3244);
nand U9648 (N_9648,N_625,N_2126);
and U9649 (N_9649,N_4143,N_4105);
and U9650 (N_9650,N_2249,N_1281);
and U9651 (N_9651,N_2928,N_1469);
or U9652 (N_9652,N_2764,N_2959);
xor U9653 (N_9653,N_958,N_1385);
or U9654 (N_9654,N_1389,N_2155);
xor U9655 (N_9655,N_4390,N_2119);
xor U9656 (N_9656,N_3752,N_4522);
or U9657 (N_9657,N_2072,N_4518);
xor U9658 (N_9658,N_4190,N_4216);
nand U9659 (N_9659,N_2286,N_3598);
or U9660 (N_9660,N_2797,N_486);
nand U9661 (N_9661,N_2082,N_3723);
xnor U9662 (N_9662,N_2662,N_2356);
and U9663 (N_9663,N_4196,N_4760);
xor U9664 (N_9664,N_858,N_2361);
nor U9665 (N_9665,N_4260,N_4935);
and U9666 (N_9666,N_2334,N_3853);
or U9667 (N_9667,N_3120,N_3589);
and U9668 (N_9668,N_2781,N_3511);
nor U9669 (N_9669,N_2930,N_306);
and U9670 (N_9670,N_1211,N_1821);
xnor U9671 (N_9671,N_1190,N_1065);
nor U9672 (N_9672,N_563,N_2890);
or U9673 (N_9673,N_1356,N_1615);
and U9674 (N_9674,N_200,N_3043);
or U9675 (N_9675,N_1834,N_3908);
nand U9676 (N_9676,N_1374,N_1905);
nor U9677 (N_9677,N_3250,N_1504);
nand U9678 (N_9678,N_2960,N_991);
xor U9679 (N_9679,N_3539,N_573);
and U9680 (N_9680,N_3189,N_4755);
or U9681 (N_9681,N_1771,N_552);
nor U9682 (N_9682,N_2116,N_3436);
nor U9683 (N_9683,N_879,N_4624);
xnor U9684 (N_9684,N_2234,N_1467);
or U9685 (N_9685,N_4031,N_4418);
and U9686 (N_9686,N_1301,N_549);
nor U9687 (N_9687,N_1718,N_1848);
nand U9688 (N_9688,N_4813,N_4025);
or U9689 (N_9689,N_4259,N_938);
or U9690 (N_9690,N_2129,N_1359);
nand U9691 (N_9691,N_3247,N_1334);
or U9692 (N_9692,N_322,N_4080);
and U9693 (N_9693,N_2319,N_249);
xnor U9694 (N_9694,N_2000,N_476);
and U9695 (N_9695,N_3450,N_1764);
nor U9696 (N_9696,N_968,N_2012);
xor U9697 (N_9697,N_4737,N_805);
xnor U9698 (N_9698,N_981,N_4925);
nor U9699 (N_9699,N_2852,N_2710);
xnor U9700 (N_9700,N_4402,N_4604);
nor U9701 (N_9701,N_4363,N_4689);
or U9702 (N_9702,N_549,N_242);
or U9703 (N_9703,N_51,N_3754);
nor U9704 (N_9704,N_1210,N_3255);
and U9705 (N_9705,N_1855,N_4876);
nor U9706 (N_9706,N_3885,N_49);
nor U9707 (N_9707,N_1214,N_1930);
or U9708 (N_9708,N_2726,N_988);
or U9709 (N_9709,N_3007,N_781);
nand U9710 (N_9710,N_1744,N_2798);
or U9711 (N_9711,N_4111,N_2012);
nand U9712 (N_9712,N_3728,N_3950);
xor U9713 (N_9713,N_1723,N_1773);
or U9714 (N_9714,N_595,N_3511);
nor U9715 (N_9715,N_3829,N_355);
or U9716 (N_9716,N_1572,N_920);
nor U9717 (N_9717,N_3966,N_2265);
nand U9718 (N_9718,N_686,N_1858);
nand U9719 (N_9719,N_542,N_2488);
xor U9720 (N_9720,N_1061,N_4031);
nand U9721 (N_9721,N_3173,N_2043);
xnor U9722 (N_9722,N_245,N_62);
or U9723 (N_9723,N_2907,N_395);
nor U9724 (N_9724,N_4003,N_4705);
nor U9725 (N_9725,N_3471,N_2277);
xor U9726 (N_9726,N_2575,N_1970);
and U9727 (N_9727,N_2363,N_3097);
or U9728 (N_9728,N_2584,N_3918);
nor U9729 (N_9729,N_180,N_1645);
or U9730 (N_9730,N_2338,N_4123);
nand U9731 (N_9731,N_3218,N_3152);
or U9732 (N_9732,N_2970,N_3193);
nand U9733 (N_9733,N_972,N_1711);
or U9734 (N_9734,N_1175,N_1949);
nand U9735 (N_9735,N_2042,N_1154);
and U9736 (N_9736,N_4929,N_4047);
or U9737 (N_9737,N_820,N_688);
xor U9738 (N_9738,N_1409,N_1957);
and U9739 (N_9739,N_989,N_2654);
and U9740 (N_9740,N_3327,N_1580);
or U9741 (N_9741,N_250,N_3427);
nor U9742 (N_9742,N_1537,N_2844);
or U9743 (N_9743,N_4018,N_786);
xor U9744 (N_9744,N_3690,N_2316);
xnor U9745 (N_9745,N_4869,N_3524);
and U9746 (N_9746,N_3103,N_726);
nand U9747 (N_9747,N_3091,N_2576);
and U9748 (N_9748,N_3868,N_3995);
nand U9749 (N_9749,N_1202,N_3485);
or U9750 (N_9750,N_2421,N_1721);
nor U9751 (N_9751,N_3457,N_4115);
and U9752 (N_9752,N_2792,N_167);
nor U9753 (N_9753,N_2354,N_4265);
and U9754 (N_9754,N_3538,N_1685);
and U9755 (N_9755,N_2781,N_1784);
nor U9756 (N_9756,N_4719,N_4484);
nor U9757 (N_9757,N_3165,N_4893);
xor U9758 (N_9758,N_482,N_2275);
and U9759 (N_9759,N_4524,N_3905);
or U9760 (N_9760,N_3838,N_1271);
and U9761 (N_9761,N_2036,N_1986);
or U9762 (N_9762,N_4073,N_4712);
or U9763 (N_9763,N_4368,N_4209);
nor U9764 (N_9764,N_2382,N_1687);
and U9765 (N_9765,N_4371,N_786);
nand U9766 (N_9766,N_1397,N_476);
nor U9767 (N_9767,N_1496,N_914);
or U9768 (N_9768,N_1328,N_4026);
or U9769 (N_9769,N_277,N_1015);
nand U9770 (N_9770,N_2751,N_922);
and U9771 (N_9771,N_3935,N_4018);
xnor U9772 (N_9772,N_2573,N_958);
or U9773 (N_9773,N_2537,N_3049);
xnor U9774 (N_9774,N_4856,N_4857);
and U9775 (N_9775,N_2701,N_1332);
xor U9776 (N_9776,N_4820,N_2818);
nand U9777 (N_9777,N_4268,N_874);
or U9778 (N_9778,N_333,N_1118);
nand U9779 (N_9779,N_887,N_3862);
nand U9780 (N_9780,N_1713,N_4833);
nor U9781 (N_9781,N_3609,N_4584);
or U9782 (N_9782,N_2593,N_327);
or U9783 (N_9783,N_1460,N_1497);
xnor U9784 (N_9784,N_3556,N_3117);
xor U9785 (N_9785,N_411,N_3924);
nand U9786 (N_9786,N_83,N_4006);
or U9787 (N_9787,N_446,N_3721);
or U9788 (N_9788,N_2568,N_3617);
nor U9789 (N_9789,N_4836,N_2749);
and U9790 (N_9790,N_3706,N_4313);
xnor U9791 (N_9791,N_1363,N_4181);
nor U9792 (N_9792,N_3912,N_930);
xnor U9793 (N_9793,N_4238,N_3693);
or U9794 (N_9794,N_2010,N_4528);
nand U9795 (N_9795,N_1922,N_4601);
nor U9796 (N_9796,N_2038,N_2521);
nor U9797 (N_9797,N_653,N_2920);
and U9798 (N_9798,N_4517,N_3974);
and U9799 (N_9799,N_2197,N_1420);
nor U9800 (N_9800,N_4981,N_3118);
nor U9801 (N_9801,N_1951,N_249);
nor U9802 (N_9802,N_835,N_3820);
xnor U9803 (N_9803,N_4661,N_3359);
or U9804 (N_9804,N_1775,N_446);
xor U9805 (N_9805,N_233,N_4445);
nor U9806 (N_9806,N_909,N_3928);
xor U9807 (N_9807,N_4165,N_4224);
or U9808 (N_9808,N_2302,N_2450);
nand U9809 (N_9809,N_1779,N_4061);
nor U9810 (N_9810,N_1268,N_1974);
or U9811 (N_9811,N_2911,N_50);
or U9812 (N_9812,N_4883,N_2621);
nor U9813 (N_9813,N_2639,N_3421);
and U9814 (N_9814,N_3328,N_1268);
or U9815 (N_9815,N_2783,N_633);
or U9816 (N_9816,N_3962,N_3623);
and U9817 (N_9817,N_4270,N_10);
nand U9818 (N_9818,N_1257,N_2218);
or U9819 (N_9819,N_1498,N_4310);
nand U9820 (N_9820,N_1096,N_4056);
xor U9821 (N_9821,N_2962,N_4403);
or U9822 (N_9822,N_2640,N_2591);
nand U9823 (N_9823,N_2095,N_4532);
xor U9824 (N_9824,N_493,N_1432);
nor U9825 (N_9825,N_1807,N_239);
or U9826 (N_9826,N_528,N_1476);
xnor U9827 (N_9827,N_4820,N_414);
nand U9828 (N_9828,N_1728,N_3868);
and U9829 (N_9829,N_137,N_1502);
nor U9830 (N_9830,N_1325,N_3405);
xor U9831 (N_9831,N_314,N_448);
xor U9832 (N_9832,N_150,N_615);
or U9833 (N_9833,N_2305,N_1036);
or U9834 (N_9834,N_875,N_1499);
and U9835 (N_9835,N_4919,N_3394);
or U9836 (N_9836,N_3190,N_1705);
nand U9837 (N_9837,N_4087,N_3528);
and U9838 (N_9838,N_2743,N_1028);
nand U9839 (N_9839,N_336,N_626);
nor U9840 (N_9840,N_3149,N_4212);
or U9841 (N_9841,N_912,N_2307);
and U9842 (N_9842,N_20,N_3479);
or U9843 (N_9843,N_3127,N_3424);
nor U9844 (N_9844,N_2458,N_2754);
or U9845 (N_9845,N_4538,N_151);
or U9846 (N_9846,N_3478,N_1176);
nand U9847 (N_9847,N_1817,N_1833);
nand U9848 (N_9848,N_559,N_4149);
and U9849 (N_9849,N_1182,N_1202);
or U9850 (N_9850,N_2797,N_4193);
or U9851 (N_9851,N_1332,N_3891);
and U9852 (N_9852,N_2241,N_338);
or U9853 (N_9853,N_2553,N_2576);
or U9854 (N_9854,N_2392,N_2335);
nor U9855 (N_9855,N_4675,N_2343);
or U9856 (N_9856,N_4996,N_4780);
xnor U9857 (N_9857,N_2602,N_313);
xnor U9858 (N_9858,N_1672,N_1013);
nor U9859 (N_9859,N_2514,N_2411);
xor U9860 (N_9860,N_1316,N_452);
or U9861 (N_9861,N_2231,N_639);
or U9862 (N_9862,N_3226,N_1484);
xnor U9863 (N_9863,N_985,N_4238);
and U9864 (N_9864,N_4153,N_1574);
nand U9865 (N_9865,N_2070,N_4601);
xor U9866 (N_9866,N_3852,N_4256);
xnor U9867 (N_9867,N_2646,N_4643);
xnor U9868 (N_9868,N_3262,N_3210);
nand U9869 (N_9869,N_2359,N_308);
nor U9870 (N_9870,N_2692,N_4845);
xor U9871 (N_9871,N_881,N_952);
or U9872 (N_9872,N_1754,N_3787);
nand U9873 (N_9873,N_3474,N_1684);
or U9874 (N_9874,N_2362,N_119);
nand U9875 (N_9875,N_255,N_3884);
xnor U9876 (N_9876,N_1804,N_2602);
and U9877 (N_9877,N_4380,N_4477);
or U9878 (N_9878,N_4604,N_690);
or U9879 (N_9879,N_4916,N_99);
or U9880 (N_9880,N_3883,N_3915);
xnor U9881 (N_9881,N_2370,N_239);
and U9882 (N_9882,N_921,N_3756);
xnor U9883 (N_9883,N_2257,N_549);
or U9884 (N_9884,N_767,N_1499);
nand U9885 (N_9885,N_2619,N_456);
and U9886 (N_9886,N_1115,N_1596);
xnor U9887 (N_9887,N_2567,N_1466);
and U9888 (N_9888,N_4063,N_3376);
or U9889 (N_9889,N_1004,N_318);
nor U9890 (N_9890,N_3474,N_25);
nor U9891 (N_9891,N_1570,N_3197);
and U9892 (N_9892,N_3982,N_4143);
nor U9893 (N_9893,N_3701,N_2182);
xnor U9894 (N_9894,N_4418,N_2567);
xor U9895 (N_9895,N_2963,N_2816);
or U9896 (N_9896,N_4085,N_2917);
nand U9897 (N_9897,N_4317,N_1717);
and U9898 (N_9898,N_2527,N_4743);
nand U9899 (N_9899,N_462,N_2201);
xor U9900 (N_9900,N_4182,N_4935);
nand U9901 (N_9901,N_1650,N_4486);
or U9902 (N_9902,N_2502,N_2994);
nand U9903 (N_9903,N_4787,N_1892);
and U9904 (N_9904,N_1086,N_3042);
and U9905 (N_9905,N_3112,N_1293);
nor U9906 (N_9906,N_2678,N_2077);
nor U9907 (N_9907,N_2737,N_3793);
xnor U9908 (N_9908,N_4102,N_1618);
xor U9909 (N_9909,N_1455,N_4960);
and U9910 (N_9910,N_1863,N_2080);
nor U9911 (N_9911,N_3897,N_2551);
nand U9912 (N_9912,N_4610,N_3230);
xor U9913 (N_9913,N_2517,N_3966);
xnor U9914 (N_9914,N_4253,N_357);
xnor U9915 (N_9915,N_11,N_1938);
nand U9916 (N_9916,N_2489,N_4718);
xor U9917 (N_9917,N_174,N_453);
nor U9918 (N_9918,N_2954,N_4090);
xor U9919 (N_9919,N_4272,N_2100);
xor U9920 (N_9920,N_2548,N_3306);
and U9921 (N_9921,N_1290,N_1214);
or U9922 (N_9922,N_119,N_4021);
nand U9923 (N_9923,N_1171,N_4112);
or U9924 (N_9924,N_898,N_3420);
nor U9925 (N_9925,N_747,N_2505);
xnor U9926 (N_9926,N_3737,N_663);
or U9927 (N_9927,N_747,N_600);
nor U9928 (N_9928,N_979,N_1777);
nor U9929 (N_9929,N_360,N_2939);
xor U9930 (N_9930,N_629,N_3682);
nand U9931 (N_9931,N_1135,N_717);
xor U9932 (N_9932,N_888,N_1696);
xnor U9933 (N_9933,N_4803,N_3628);
nand U9934 (N_9934,N_236,N_2622);
nand U9935 (N_9935,N_4238,N_3430);
or U9936 (N_9936,N_3794,N_2472);
nor U9937 (N_9937,N_65,N_2979);
nor U9938 (N_9938,N_4013,N_1917);
nand U9939 (N_9939,N_3344,N_4686);
nor U9940 (N_9940,N_3656,N_2718);
nand U9941 (N_9941,N_985,N_1135);
xor U9942 (N_9942,N_4668,N_3517);
xnor U9943 (N_9943,N_1138,N_1755);
xnor U9944 (N_9944,N_3444,N_3173);
or U9945 (N_9945,N_4969,N_1368);
or U9946 (N_9946,N_1872,N_2129);
nor U9947 (N_9947,N_4221,N_4404);
nand U9948 (N_9948,N_1100,N_2945);
and U9949 (N_9949,N_4408,N_508);
or U9950 (N_9950,N_4796,N_1866);
and U9951 (N_9951,N_4694,N_946);
xor U9952 (N_9952,N_4424,N_1599);
nor U9953 (N_9953,N_2352,N_2722);
or U9954 (N_9954,N_3083,N_199);
xor U9955 (N_9955,N_2466,N_60);
and U9956 (N_9956,N_625,N_768);
nand U9957 (N_9957,N_1905,N_1067);
or U9958 (N_9958,N_4625,N_4631);
nor U9959 (N_9959,N_2514,N_1917);
nand U9960 (N_9960,N_1507,N_2310);
nor U9961 (N_9961,N_2778,N_2673);
nand U9962 (N_9962,N_1284,N_153);
nor U9963 (N_9963,N_4557,N_2510);
xor U9964 (N_9964,N_3554,N_2347);
nor U9965 (N_9965,N_763,N_3132);
nand U9966 (N_9966,N_2723,N_4918);
nand U9967 (N_9967,N_3172,N_376);
nand U9968 (N_9968,N_619,N_4291);
nor U9969 (N_9969,N_4955,N_3450);
or U9970 (N_9970,N_4467,N_3553);
and U9971 (N_9971,N_4506,N_3252);
xor U9972 (N_9972,N_4228,N_269);
or U9973 (N_9973,N_2137,N_248);
or U9974 (N_9974,N_2108,N_1337);
nand U9975 (N_9975,N_684,N_792);
xnor U9976 (N_9976,N_2044,N_854);
xor U9977 (N_9977,N_2457,N_1124);
xor U9978 (N_9978,N_952,N_3329);
nor U9979 (N_9979,N_1503,N_2665);
nor U9980 (N_9980,N_2891,N_4766);
xnor U9981 (N_9981,N_4613,N_869);
and U9982 (N_9982,N_3462,N_973);
xor U9983 (N_9983,N_4800,N_1612);
nor U9984 (N_9984,N_3947,N_4119);
or U9985 (N_9985,N_3676,N_1263);
nor U9986 (N_9986,N_4185,N_711);
nand U9987 (N_9987,N_1893,N_4619);
and U9988 (N_9988,N_162,N_1027);
xnor U9989 (N_9989,N_3183,N_2885);
nor U9990 (N_9990,N_1040,N_4349);
xnor U9991 (N_9991,N_4384,N_4423);
nor U9992 (N_9992,N_2155,N_4845);
nand U9993 (N_9993,N_3027,N_332);
and U9994 (N_9994,N_818,N_1183);
nor U9995 (N_9995,N_3662,N_4910);
nand U9996 (N_9996,N_1046,N_1710);
or U9997 (N_9997,N_3499,N_2468);
nand U9998 (N_9998,N_4246,N_3455);
and U9999 (N_9999,N_1035,N_894);
or U10000 (N_10000,N_9631,N_7546);
or U10001 (N_10001,N_6897,N_6792);
and U10002 (N_10002,N_6547,N_9059);
or U10003 (N_10003,N_5666,N_8448);
nand U10004 (N_10004,N_8665,N_6657);
nand U10005 (N_10005,N_9434,N_8714);
and U10006 (N_10006,N_5465,N_5432);
or U10007 (N_10007,N_6829,N_9956);
and U10008 (N_10008,N_9755,N_8708);
or U10009 (N_10009,N_9689,N_8155);
nor U10010 (N_10010,N_5263,N_8329);
nand U10011 (N_10011,N_6425,N_6967);
xnor U10012 (N_10012,N_5604,N_6502);
and U10013 (N_10013,N_9833,N_7968);
nand U10014 (N_10014,N_8901,N_8897);
and U10015 (N_10015,N_5723,N_9342);
xnor U10016 (N_10016,N_9317,N_6024);
xnor U10017 (N_10017,N_5599,N_8760);
xor U10018 (N_10018,N_8612,N_7097);
xor U10019 (N_10019,N_6999,N_8356);
and U10020 (N_10020,N_8475,N_8138);
and U10021 (N_10021,N_5772,N_9111);
nor U10022 (N_10022,N_6621,N_7740);
nand U10023 (N_10023,N_8112,N_8094);
xor U10024 (N_10024,N_9516,N_9908);
or U10025 (N_10025,N_6428,N_7214);
nor U10026 (N_10026,N_9102,N_5467);
nand U10027 (N_10027,N_5710,N_7009);
xnor U10028 (N_10028,N_8966,N_7190);
xnor U10029 (N_10029,N_5522,N_5431);
or U10030 (N_10030,N_8316,N_8866);
or U10031 (N_10031,N_8693,N_9183);
nor U10032 (N_10032,N_7777,N_6185);
xnor U10033 (N_10033,N_6853,N_6316);
nand U10034 (N_10034,N_6697,N_7859);
nand U10035 (N_10035,N_5301,N_8028);
or U10036 (N_10036,N_7277,N_8829);
or U10037 (N_10037,N_8834,N_9145);
xor U10038 (N_10038,N_8869,N_6674);
nor U10039 (N_10039,N_5833,N_8682);
and U10040 (N_10040,N_9038,N_9246);
or U10041 (N_10041,N_9563,N_7269);
xor U10042 (N_10042,N_6130,N_5445);
xor U10043 (N_10043,N_9863,N_6911);
nand U10044 (N_10044,N_9674,N_7959);
or U10045 (N_10045,N_7231,N_8658);
nor U10046 (N_10046,N_8494,N_7579);
nand U10047 (N_10047,N_8501,N_5188);
or U10048 (N_10048,N_5125,N_5941);
or U10049 (N_10049,N_7517,N_5925);
nand U10050 (N_10050,N_5842,N_6073);
and U10051 (N_10051,N_8474,N_8018);
nand U10052 (N_10052,N_5179,N_8787);
nor U10053 (N_10053,N_8392,N_8046);
xnor U10054 (N_10054,N_7810,N_9235);
nor U10055 (N_10055,N_6904,N_8850);
or U10056 (N_10056,N_6727,N_7264);
xor U10057 (N_10057,N_7492,N_6492);
nand U10058 (N_10058,N_7100,N_8499);
or U10059 (N_10059,N_5657,N_5238);
nand U10060 (N_10060,N_7437,N_8201);
nand U10061 (N_10061,N_5759,N_6108);
or U10062 (N_10062,N_8275,N_6506);
and U10063 (N_10063,N_5998,N_8294);
and U10064 (N_10064,N_7762,N_5860);
nor U10065 (N_10065,N_7443,N_6921);
or U10066 (N_10066,N_9331,N_9813);
xor U10067 (N_10067,N_5069,N_8652);
nor U10068 (N_10068,N_9401,N_9670);
xor U10069 (N_10069,N_7922,N_6062);
xnor U10070 (N_10070,N_7849,N_5684);
nor U10071 (N_10071,N_6966,N_7656);
and U10072 (N_10072,N_6310,N_5953);
nand U10073 (N_10073,N_8958,N_9473);
nand U10074 (N_10074,N_7589,N_8740);
nand U10075 (N_10075,N_6679,N_9758);
xor U10076 (N_10076,N_6991,N_5575);
or U10077 (N_10077,N_9267,N_5758);
xnor U10078 (N_10078,N_8912,N_7911);
nor U10079 (N_10079,N_8167,N_9126);
or U10080 (N_10080,N_8991,N_9582);
nand U10081 (N_10081,N_6232,N_6040);
and U10082 (N_10082,N_7151,N_6916);
xnor U10083 (N_10083,N_5746,N_8809);
and U10084 (N_10084,N_8955,N_8166);
nand U10085 (N_10085,N_6034,N_6796);
or U10086 (N_10086,N_5903,N_5592);
xnor U10087 (N_10087,N_6417,N_5659);
nand U10088 (N_10088,N_9531,N_8491);
nand U10089 (N_10089,N_7555,N_9254);
and U10090 (N_10090,N_5270,N_6171);
xor U10091 (N_10091,N_9338,N_5668);
or U10092 (N_10092,N_9696,N_7882);
or U10093 (N_10093,N_5485,N_8468);
or U10094 (N_10094,N_8385,N_8214);
nand U10095 (N_10095,N_9451,N_6406);
nand U10096 (N_10096,N_6631,N_9536);
nor U10097 (N_10097,N_8697,N_5535);
nor U10098 (N_10098,N_6395,N_5434);
or U10099 (N_10099,N_9881,N_8456);
nor U10100 (N_10100,N_6128,N_8051);
or U10101 (N_10101,N_8997,N_8010);
nor U10102 (N_10102,N_9385,N_8146);
or U10103 (N_10103,N_8726,N_9284);
nand U10104 (N_10104,N_8815,N_8974);
or U10105 (N_10105,N_8030,N_7268);
nor U10106 (N_10106,N_7750,N_8766);
nor U10107 (N_10107,N_7928,N_7124);
xnor U10108 (N_10108,N_6685,N_8216);
xnor U10109 (N_10109,N_7748,N_6832);
or U10110 (N_10110,N_7973,N_6409);
nand U10111 (N_10111,N_5864,N_8916);
or U10112 (N_10112,N_8498,N_7789);
nand U10113 (N_10113,N_5131,N_5908);
nor U10114 (N_10114,N_9546,N_7294);
nand U10115 (N_10115,N_9868,N_7507);
and U10116 (N_10116,N_8909,N_9172);
xnor U10117 (N_10117,N_6422,N_9307);
xor U10118 (N_10118,N_5728,N_9879);
xnor U10119 (N_10119,N_9175,N_8221);
and U10120 (N_10120,N_7139,N_5168);
nand U10121 (N_10121,N_7909,N_9539);
nand U10122 (N_10122,N_8852,N_5486);
xnor U10123 (N_10123,N_9360,N_7431);
or U10124 (N_10124,N_8657,N_8281);
nand U10125 (N_10125,N_9333,N_7166);
nor U10126 (N_10126,N_5995,N_8607);
or U10127 (N_10127,N_8695,N_8126);
or U10128 (N_10128,N_5735,N_5001);
xnor U10129 (N_10129,N_7157,N_8649);
nor U10130 (N_10130,N_9819,N_5333);
or U10131 (N_10131,N_5816,N_7585);
xor U10132 (N_10132,N_9955,N_5958);
xnor U10133 (N_10133,N_9816,N_8836);
nand U10134 (N_10134,N_7705,N_6776);
or U10135 (N_10135,N_5137,N_9509);
or U10136 (N_10136,N_5399,N_6741);
and U10137 (N_10137,N_9469,N_9377);
or U10138 (N_10138,N_6733,N_5371);
and U10139 (N_10139,N_5021,N_7317);
and U10140 (N_10140,N_9047,N_6294);
nand U10141 (N_10141,N_6408,N_8034);
xor U10142 (N_10142,N_7474,N_7220);
or U10143 (N_10143,N_5652,N_7658);
xor U10144 (N_10144,N_5883,N_7417);
nand U10145 (N_10145,N_9514,N_5016);
nor U10146 (N_10146,N_5702,N_9060);
and U10147 (N_10147,N_7156,N_5039);
or U10148 (N_10148,N_5917,N_9089);
xnor U10149 (N_10149,N_6543,N_5002);
nand U10150 (N_10150,N_7797,N_6669);
nand U10151 (N_10151,N_6823,N_9297);
or U10152 (N_10152,N_7721,N_5897);
nor U10153 (N_10153,N_5950,N_6248);
and U10154 (N_10154,N_9131,N_9383);
and U10155 (N_10155,N_7240,N_9282);
or U10156 (N_10156,N_8659,N_9730);
or U10157 (N_10157,N_8336,N_8789);
or U10158 (N_10158,N_5916,N_7647);
nor U10159 (N_10159,N_5695,N_6524);
nor U10160 (N_10160,N_5305,N_7171);
nand U10161 (N_10161,N_9903,N_6244);
or U10162 (N_10162,N_6758,N_6884);
and U10163 (N_10163,N_7278,N_7618);
nand U10164 (N_10164,N_5559,N_8817);
nand U10165 (N_10165,N_8862,N_9084);
nand U10166 (N_10166,N_9015,N_5083);
or U10167 (N_10167,N_9750,N_6332);
nor U10168 (N_10168,N_9427,N_6311);
and U10169 (N_10169,N_5972,N_5286);
nor U10170 (N_10170,N_6893,N_6584);
nand U10171 (N_10171,N_7110,N_6362);
or U10172 (N_10172,N_9471,N_8195);
xnor U10173 (N_10173,N_6889,N_9814);
or U10174 (N_10174,N_8785,N_5080);
or U10175 (N_10175,N_6307,N_5082);
xnor U10176 (N_10176,N_6468,N_7062);
and U10177 (N_10177,N_6935,N_6116);
nor U10178 (N_10178,N_8502,N_5194);
and U10179 (N_10179,N_9849,N_6998);
and U10180 (N_10180,N_9654,N_5043);
nor U10181 (N_10181,N_7148,N_5888);
and U10182 (N_10182,N_8904,N_7074);
nand U10183 (N_10183,N_5169,N_8395);
nand U10184 (N_10184,N_6612,N_7219);
and U10185 (N_10185,N_7853,N_5354);
nor U10186 (N_10186,N_6512,N_7447);
and U10187 (N_10187,N_8527,N_8068);
or U10188 (N_10188,N_5598,N_8000);
or U10189 (N_10189,N_6732,N_5761);
nor U10190 (N_10190,N_8379,N_5546);
and U10191 (N_10191,N_9556,N_7629);
nor U10192 (N_10192,N_8405,N_6573);
and U10193 (N_10193,N_7847,N_7098);
or U10194 (N_10194,N_9732,N_5868);
xnor U10195 (N_10195,N_6634,N_5608);
xor U10196 (N_10196,N_9848,N_8238);
nor U10197 (N_10197,N_7760,N_8663);
and U10198 (N_10198,N_6483,N_6081);
nor U10199 (N_10199,N_8645,N_5412);
xor U10200 (N_10200,N_9238,N_7408);
xnor U10201 (N_10201,N_9652,N_6090);
or U10202 (N_10202,N_5554,N_8369);
nand U10203 (N_10203,N_9869,N_6389);
xnor U10204 (N_10204,N_7346,N_7085);
nand U10205 (N_10205,N_7920,N_6215);
nand U10206 (N_10206,N_8447,N_6557);
xor U10207 (N_10207,N_8193,N_9119);
xnor U10208 (N_10208,N_9229,N_7102);
or U10209 (N_10209,N_7374,N_5124);
and U10210 (N_10210,N_8187,N_5643);
or U10211 (N_10211,N_6943,N_5803);
nand U10212 (N_10212,N_5310,N_5247);
and U10213 (N_10213,N_9356,N_9421);
and U10214 (N_10214,N_6695,N_6815);
and U10215 (N_10215,N_9829,N_9265);
nand U10216 (N_10216,N_7837,N_5624);
and U10217 (N_10217,N_8826,N_8630);
or U10218 (N_10218,N_8360,N_7333);
or U10219 (N_10219,N_5831,N_5223);
and U10220 (N_10220,N_9523,N_9393);
nor U10221 (N_10221,N_7984,N_5519);
or U10222 (N_10222,N_8647,N_6193);
or U10223 (N_10223,N_8932,N_8305);
and U10224 (N_10224,N_9529,N_6055);
and U10225 (N_10225,N_7093,N_6811);
nor U10226 (N_10226,N_5778,N_8845);
nand U10227 (N_10227,N_5177,N_9057);
or U10228 (N_10228,N_8178,N_7203);
or U10229 (N_10229,N_7070,N_5924);
xor U10230 (N_10230,N_8581,N_7581);
and U10231 (N_10231,N_7173,N_6183);
nor U10232 (N_10232,N_9474,N_7245);
and U10233 (N_10233,N_9006,N_9880);
xor U10234 (N_10234,N_6749,N_8455);
nand U10235 (N_10235,N_7696,N_7530);
nand U10236 (N_10236,N_9715,N_8777);
nand U10237 (N_10237,N_5703,N_9362);
and U10238 (N_10238,N_5755,N_5515);
nor U10239 (N_10239,N_6374,N_8666);
xor U10240 (N_10240,N_8357,N_8733);
nor U10241 (N_10241,N_8765,N_5585);
nand U10242 (N_10242,N_7802,N_7573);
or U10243 (N_10243,N_9485,N_9032);
nor U10244 (N_10244,N_8082,N_6162);
nor U10245 (N_10245,N_8588,N_6706);
nand U10246 (N_10246,N_5322,N_7898);
xnor U10247 (N_10247,N_8044,N_5913);
or U10248 (N_10248,N_8457,N_8913);
nand U10249 (N_10249,N_9711,N_6281);
nor U10250 (N_10250,N_9208,N_8900);
and U10251 (N_10251,N_6987,N_8951);
and U10252 (N_10252,N_7636,N_5940);
nor U10253 (N_10253,N_6644,N_7778);
xor U10254 (N_10254,N_7635,N_9486);
nand U10255 (N_10255,N_6568,N_9454);
nor U10256 (N_10256,N_8846,N_6069);
and U10257 (N_10257,N_5784,N_9063);
and U10258 (N_10258,N_5549,N_8865);
nand U10259 (N_10259,N_5904,N_6887);
nor U10260 (N_10260,N_9649,N_9989);
or U10261 (N_10261,N_9919,N_7997);
xnor U10262 (N_10262,N_6835,N_5642);
xnor U10263 (N_10263,N_8495,N_6348);
and U10264 (N_10264,N_5662,N_7508);
nand U10265 (N_10265,N_8960,N_5437);
nand U10266 (N_10266,N_5867,N_7255);
xor U10267 (N_10267,N_7314,N_5335);
or U10268 (N_10268,N_9405,N_7529);
nor U10269 (N_10269,N_6646,N_7661);
nand U10270 (N_10270,N_8574,N_9325);
nand U10271 (N_10271,N_7996,N_6460);
and U10272 (N_10272,N_7838,N_9211);
nand U10273 (N_10273,N_7910,N_9097);
nand U10274 (N_10274,N_6444,N_5099);
or U10275 (N_10275,N_5203,N_5248);
and U10276 (N_10276,N_9044,N_5553);
or U10277 (N_10277,N_8505,N_6058);
xnor U10278 (N_10278,N_6005,N_9628);
nand U10279 (N_10279,N_6289,N_6440);
xor U10280 (N_10280,N_5729,N_9054);
nor U10281 (N_10281,N_6877,N_7514);
nand U10282 (N_10282,N_6447,N_8304);
xnor U10283 (N_10283,N_7484,N_5220);
nand U10284 (N_10284,N_5473,N_8349);
nand U10285 (N_10285,N_5423,N_8061);
nor U10286 (N_10286,N_8711,N_5356);
or U10287 (N_10287,N_7744,N_9984);
xor U10288 (N_10288,N_7205,N_9419);
nand U10289 (N_10289,N_8521,N_8081);
nand U10290 (N_10290,N_5147,N_9502);
or U10291 (N_10291,N_7160,N_5201);
nand U10292 (N_10292,N_8141,N_9672);
xnor U10293 (N_10293,N_6497,N_9422);
nor U10294 (N_10294,N_9125,N_9720);
nand U10295 (N_10295,N_5540,N_5312);
nand U10296 (N_10296,N_7518,N_8375);
and U10297 (N_10297,N_5954,N_9406);
nor U10298 (N_10298,N_7243,N_5128);
nor U10299 (N_10299,N_6910,N_7186);
and U10300 (N_10300,N_8319,N_8365);
nand U10301 (N_10301,N_8688,N_5190);
nor U10302 (N_10302,N_6230,N_7247);
nor U10303 (N_10303,N_9058,N_9043);
and U10304 (N_10304,N_5200,N_5199);
and U10305 (N_10305,N_8032,N_6586);
xnor U10306 (N_10306,N_6759,N_6849);
and U10307 (N_10307,N_9895,N_9252);
and U10308 (N_10308,N_7967,N_7500);
xnor U10309 (N_10309,N_8444,N_5284);
nand U10310 (N_10310,N_7653,N_8506);
or U10311 (N_10311,N_5006,N_6720);
xnor U10312 (N_10312,N_6735,N_9947);
and U10313 (N_10313,N_5550,N_5583);
or U10314 (N_10314,N_5104,N_5629);
nand U10315 (N_10315,N_8290,N_8824);
and U10316 (N_10316,N_8552,N_8282);
nor U10317 (N_10317,N_5588,N_9219);
or U10318 (N_10318,N_9533,N_9190);
nand U10319 (N_10319,N_6789,N_8935);
xor U10320 (N_10320,N_5479,N_7736);
nand U10321 (N_10321,N_6223,N_9936);
nand U10322 (N_10322,N_8377,N_9667);
and U10323 (N_10323,N_8429,N_6578);
nand U10324 (N_10324,N_5106,N_9453);
and U10325 (N_10325,N_8539,N_6773);
nand U10326 (N_10326,N_6595,N_9142);
or U10327 (N_10327,N_6534,N_5751);
xnor U10328 (N_10328,N_9818,N_8918);
nand U10329 (N_10329,N_7800,N_5173);
xor U10330 (N_10330,N_9821,N_7570);
or U10331 (N_10331,N_6477,N_8827);
xor U10332 (N_10332,N_9806,N_9226);
nand U10333 (N_10333,N_8397,N_5456);
xnor U10334 (N_10334,N_8119,N_5876);
xnor U10335 (N_10335,N_8313,N_9121);
nor U10336 (N_10336,N_8084,N_5385);
nand U10337 (N_10337,N_6737,N_7267);
and U10338 (N_10338,N_6400,N_5490);
xnor U10339 (N_10339,N_7767,N_8348);
nand U10340 (N_10340,N_7167,N_6672);
or U10341 (N_10341,N_7540,N_9718);
and U10342 (N_10342,N_6766,N_9756);
and U10343 (N_10343,N_9149,N_6583);
nor U10344 (N_10344,N_6820,N_6429);
or U10345 (N_10345,N_7120,N_8107);
xnor U10346 (N_10346,N_9040,N_6635);
and U10347 (N_10347,N_6828,N_5215);
or U10348 (N_10348,N_9929,N_7378);
or U10349 (N_10349,N_5225,N_6690);
and U10350 (N_10350,N_8315,N_6702);
nor U10351 (N_10351,N_6202,N_7329);
nand U10352 (N_10352,N_8611,N_5430);
nand U10353 (N_10353,N_9553,N_7979);
and U10354 (N_10354,N_7065,N_9329);
or U10355 (N_10355,N_6590,N_9200);
nand U10356 (N_10356,N_9852,N_7370);
or U10357 (N_10357,N_8863,N_8067);
nor U10358 (N_10358,N_9295,N_8985);
xor U10359 (N_10359,N_7908,N_5066);
nor U10360 (N_10360,N_9371,N_5073);
xor U10361 (N_10361,N_5115,N_8414);
nor U10362 (N_10362,N_5514,N_7929);
nor U10363 (N_10363,N_7526,N_6139);
or U10364 (N_10364,N_9260,N_9207);
xnor U10365 (N_10365,N_9538,N_6035);
or U10366 (N_10366,N_7196,N_7189);
nand U10367 (N_10367,N_6225,N_7468);
or U10368 (N_10368,N_9171,N_6436);
nor U10369 (N_10369,N_5476,N_7850);
or U10370 (N_10370,N_8871,N_8434);
xnor U10371 (N_10371,N_9289,N_7108);
nor U10372 (N_10372,N_9028,N_8684);
nor U10373 (N_10373,N_8860,N_9954);
nand U10374 (N_10374,N_9540,N_7622);
and U10375 (N_10375,N_7983,N_6495);
xnor U10376 (N_10376,N_5074,N_7538);
xor U10377 (N_10377,N_9633,N_9867);
and U10378 (N_10378,N_6950,N_6156);
nor U10379 (N_10379,N_8939,N_7690);
nand U10380 (N_10380,N_8259,N_6328);
xnor U10381 (N_10381,N_7819,N_6074);
or U10382 (N_10382,N_9993,N_5722);
xor U10383 (N_10383,N_9907,N_6504);
xnor U10384 (N_10384,N_6442,N_6196);
or U10385 (N_10385,N_7942,N_9447);
nor U10386 (N_10386,N_6656,N_5411);
and U10387 (N_10387,N_5108,N_8840);
and U10388 (N_10388,N_6216,N_6517);
nor U10389 (N_10389,N_5294,N_6698);
nand U10390 (N_10390,N_6012,N_7643);
nand U10391 (N_10391,N_8400,N_7498);
nor U10392 (N_10392,N_8274,N_5040);
or U10393 (N_10393,N_8022,N_5548);
nand U10394 (N_10394,N_7966,N_6859);
or U10395 (N_10395,N_8337,N_8592);
nand U10396 (N_10396,N_9702,N_8134);
nand U10397 (N_10397,N_5753,N_5407);
and U10398 (N_10398,N_5155,N_7044);
xnor U10399 (N_10399,N_6098,N_5697);
nand U10400 (N_10400,N_5576,N_8549);
nor U10401 (N_10401,N_5851,N_7752);
nand U10402 (N_10402,N_9855,N_8910);
nand U10403 (N_10403,N_7040,N_9775);
or U10404 (N_10404,N_9515,N_6218);
xor U10405 (N_10405,N_7300,N_5826);
and U10406 (N_10406,N_8393,N_8384);
xor U10407 (N_10407,N_5603,N_6742);
or U10408 (N_10408,N_8604,N_9290);
nand U10409 (N_10409,N_5366,N_7115);
nor U10410 (N_10410,N_9146,N_9668);
nor U10411 (N_10411,N_8739,N_8945);
nand U10412 (N_10412,N_7184,N_6404);
or U10413 (N_10413,N_8575,N_9986);
nand U10414 (N_10414,N_9739,N_6599);
nand U10415 (N_10415,N_5019,N_6153);
or U10416 (N_10416,N_8706,N_5853);
and U10417 (N_10417,N_6449,N_7473);
and U10418 (N_10418,N_6673,N_5834);
nor U10419 (N_10419,N_8266,N_8270);
and U10420 (N_10420,N_6653,N_5672);
nor U10421 (N_10421,N_6942,N_5180);
or U10422 (N_10422,N_6976,N_9999);
nor U10423 (N_10423,N_9657,N_6148);
nand U10424 (N_10424,N_6953,N_8524);
xor U10425 (N_10425,N_6858,N_8643);
nand U10426 (N_10426,N_8116,N_9321);
and U10427 (N_10427,N_9611,N_6700);
xnor U10428 (N_10428,N_6496,N_9817);
xnor U10429 (N_10429,N_7509,N_8778);
or U10430 (N_10430,N_8531,N_6151);
and U10431 (N_10431,N_6334,N_9217);
nor U10432 (N_10432,N_7117,N_6944);
nor U10433 (N_10433,N_8186,N_7860);
xor U10434 (N_10434,N_5339,N_7731);
or U10435 (N_10435,N_8048,N_6838);
or U10436 (N_10436,N_7071,N_9594);
nor U10437 (N_10437,N_6734,N_9547);
or U10438 (N_10438,N_9107,N_6474);
or U10439 (N_10439,N_7801,N_9607);
and U10440 (N_10440,N_5645,N_8914);
xor U10441 (N_10441,N_6813,N_5863);
xor U10442 (N_10442,N_7919,N_5494);
xnor U10443 (N_10443,N_8689,N_5796);
and U10444 (N_10444,N_7136,N_9932);
or U10445 (N_10445,N_9315,N_6561);
nand U10446 (N_10446,N_5785,N_8399);
xnor U10447 (N_10447,N_7449,N_7852);
or U10448 (N_10448,N_7805,N_8250);
or U10449 (N_10449,N_9724,N_6333);
nor U10450 (N_10450,N_5718,N_9931);
nand U10451 (N_10451,N_6964,N_6272);
or U10452 (N_10452,N_8308,N_7524);
or U10453 (N_10453,N_8424,N_6382);
nand U10454 (N_10454,N_5810,N_5397);
nand U10455 (N_10455,N_6782,N_5845);
nand U10456 (N_10456,N_8218,N_8302);
nor U10457 (N_10457,N_5383,N_7315);
and U10458 (N_10458,N_5633,N_6243);
xnor U10459 (N_10459,N_7497,N_8359);
and U10460 (N_10460,N_5480,N_9345);
xor U10461 (N_10461,N_5105,N_9964);
and U10462 (N_10462,N_5052,N_7487);
xnor U10463 (N_10463,N_8439,N_9928);
nand U10464 (N_10464,N_8234,N_8754);
nand U10465 (N_10465,N_6091,N_9468);
or U10466 (N_10466,N_5566,N_7980);
nor U10467 (N_10467,N_9640,N_9202);
and U10468 (N_10468,N_7265,N_7254);
or U10469 (N_10469,N_5113,N_5139);
xnor U10470 (N_10470,N_7904,N_8558);
nor U10471 (N_10471,N_8323,N_6668);
and U10472 (N_10472,N_5900,N_7651);
nor U10473 (N_10473,N_6963,N_5474);
or U10474 (N_10474,N_8350,N_9969);
and U10475 (N_10475,N_6433,N_8470);
xnor U10476 (N_10476,N_5240,N_9410);
or U10477 (N_10477,N_7357,N_8798);
nor U10478 (N_10478,N_8858,N_9568);
and U10479 (N_10479,N_5376,N_9379);
xor U10480 (N_10480,N_7554,N_6288);
nand U10481 (N_10481,N_8127,N_5462);
and U10482 (N_10482,N_9407,N_7745);
nor U10483 (N_10483,N_5902,N_5628);
nand U10484 (N_10484,N_5320,N_8841);
xnor U10485 (N_10485,N_5975,N_7703);
nand U10486 (N_10486,N_6762,N_9328);
or U10487 (N_10487,N_5616,N_7289);
or U10488 (N_10488,N_8398,N_6387);
and U10489 (N_10489,N_9092,N_6274);
nor U10490 (N_10490,N_9452,N_5438);
nand U10491 (N_10491,N_9206,N_6170);
nor U10492 (N_10492,N_5946,N_5389);
or U10493 (N_10493,N_7737,N_5939);
and U10494 (N_10494,N_8775,N_8964);
nand U10495 (N_10495,N_8299,N_6650);
and U10496 (N_10496,N_5891,N_9904);
or U10497 (N_10497,N_8838,N_5792);
and U10498 (N_10498,N_9095,N_7418);
nand U10499 (N_10499,N_6271,N_7272);
nand U10500 (N_10500,N_6095,N_7410);
nand U10501 (N_10501,N_6724,N_7769);
and U10502 (N_10502,N_9583,N_7930);
or U10503 (N_10503,N_5258,N_5675);
and U10504 (N_10504,N_6908,N_7130);
nor U10505 (N_10505,N_6349,N_7229);
nor U10506 (N_10506,N_9512,N_8861);
nor U10507 (N_10507,N_8412,N_9048);
or U10508 (N_10508,N_7562,N_9760);
xnor U10509 (N_10509,N_8569,N_8756);
xor U10510 (N_10510,N_9558,N_9710);
xnor U10511 (N_10511,N_6705,N_5622);
and U10512 (N_10512,N_9830,N_8965);
xor U10513 (N_10513,N_9236,N_9358);
nand U10514 (N_10514,N_9629,N_6262);
xnor U10515 (N_10515,N_6140,N_5373);
or U10516 (N_10516,N_8232,N_7328);
nor U10517 (N_10517,N_9638,N_6546);
nand U10518 (N_10518,N_6161,N_6390);
xor U10519 (N_10519,N_9279,N_7702);
or U10520 (N_10520,N_6801,N_7035);
and U10521 (N_10521,N_7181,N_8538);
or U10522 (N_10522,N_5517,N_5224);
xor U10523 (N_10523,N_9612,N_5931);
nand U10524 (N_10524,N_8477,N_9416);
nor U10525 (N_10525,N_7659,N_7131);
nor U10526 (N_10526,N_9905,N_8550);
and U10527 (N_10527,N_7488,N_9627);
nor U10528 (N_10528,N_9866,N_7271);
nand U10529 (N_10529,N_9354,N_5982);
and U10530 (N_10530,N_5817,N_7393);
nor U10531 (N_10531,N_6684,N_8883);
and U10532 (N_10532,N_8700,N_9094);
and U10533 (N_10533,N_5750,N_9293);
or U10534 (N_10534,N_5459,N_9274);
xnor U10535 (N_10535,N_5451,N_5823);
and U10536 (N_10536,N_5951,N_5731);
nor U10537 (N_10537,N_9162,N_6491);
or U10538 (N_10538,N_9165,N_9024);
nand U10539 (N_10539,N_8153,N_9648);
xnor U10540 (N_10540,N_9774,N_9554);
nand U10541 (N_10541,N_5318,N_9505);
nor U10542 (N_10542,N_5452,N_9692);
nand U10543 (N_10543,N_7896,N_6299);
or U10544 (N_10544,N_6461,N_5153);
xor U10545 (N_10545,N_8854,N_6445);
or U10546 (N_10546,N_9941,N_8980);
xnor U10547 (N_10547,N_9201,N_5390);
nor U10548 (N_10548,N_9911,N_8229);
nand U10549 (N_10549,N_6301,N_6687);
or U10550 (N_10550,N_7007,N_8781);
and U10551 (N_10551,N_9170,N_7052);
nand U10552 (N_10552,N_9676,N_5237);
nand U10553 (N_10553,N_5516,N_6637);
nand U10554 (N_10554,N_6509,N_5307);
nand U10555 (N_10555,N_5687,N_6628);
xor U10556 (N_10556,N_5667,N_6154);
nor U10557 (N_10557,N_9838,N_7954);
xnor U10558 (N_10558,N_7432,N_6804);
or U10559 (N_10559,N_5386,N_7577);
or U10560 (N_10560,N_8842,N_7757);
nor U10561 (N_10561,N_5890,N_9445);
or U10562 (N_10562,N_7844,N_7999);
nand U10563 (N_10563,N_9925,N_9924);
or U10564 (N_10564,N_8843,N_9917);
and U10565 (N_10565,N_9725,N_6806);
nor U10566 (N_10566,N_8047,N_6540);
xor U10567 (N_10567,N_6228,N_8536);
nor U10568 (N_10568,N_9576,N_9161);
nor U10569 (N_10569,N_7429,N_5369);
and U10570 (N_10570,N_7634,N_5055);
nand U10571 (N_10571,N_6971,N_8441);
and U10572 (N_10572,N_7121,N_7599);
or U10573 (N_10573,N_8076,N_6711);
and U10574 (N_10574,N_9087,N_8008);
nor U10575 (N_10575,N_9621,N_5911);
or U10576 (N_10576,N_5518,N_7187);
xor U10577 (N_10577,N_8496,N_7209);
nand U10578 (N_10578,N_6329,N_7695);
and U10579 (N_10579,N_6596,N_5738);
xnor U10580 (N_10580,N_6136,N_5565);
xor U10581 (N_10581,N_7128,N_7558);
nand U10582 (N_10582,N_7681,N_7461);
nand U10583 (N_10583,N_5988,N_8479);
or U10584 (N_10584,N_7854,N_6624);
nor U10585 (N_10585,N_5578,N_6753);
nand U10586 (N_10586,N_5461,N_5324);
and U10587 (N_10587,N_9898,N_7846);
or U10588 (N_10588,N_6948,N_8742);
nor U10589 (N_10589,N_8467,N_9042);
or U10590 (N_10590,N_8362,N_9365);
nor U10591 (N_10591,N_6376,N_8938);
nor U10592 (N_10592,N_8176,N_9687);
nand U10593 (N_10593,N_5906,N_8092);
or U10594 (N_10594,N_5768,N_6601);
nand U10595 (N_10595,N_8066,N_5062);
and U10596 (N_10596,N_9203,N_9461);
nor U10597 (N_10597,N_5351,N_7799);
nor U10598 (N_10598,N_6250,N_7666);
or U10599 (N_10599,N_8462,N_6319);
and U10600 (N_10600,N_9090,N_8318);
nor U10601 (N_10601,N_9458,N_5370);
and U10602 (N_10602,N_6723,N_8968);
and U10603 (N_10603,N_9831,N_9180);
nor U10604 (N_10604,N_9423,N_9415);
nor U10605 (N_10605,N_6844,N_5887);
nor U10606 (N_10606,N_6989,N_7215);
and U10607 (N_10607,N_9382,N_8300);
or U10608 (N_10608,N_8844,N_7101);
nor U10609 (N_10609,N_7824,N_9240);
xor U10610 (N_10610,N_7103,N_7192);
nand U10611 (N_10611,N_7326,N_9997);
nand U10612 (N_10612,N_8197,N_5261);
nor U10613 (N_10613,N_5713,N_6508);
or U10614 (N_10614,N_7786,N_5513);
or U10615 (N_10615,N_9220,N_5676);
or U10616 (N_10616,N_9264,N_9772);
xnor U10617 (N_10617,N_5274,N_5724);
or U10618 (N_10618,N_7361,N_9796);
nor U10619 (N_10619,N_6326,N_6107);
nand U10620 (N_10620,N_9744,N_8507);
nand U10621 (N_10621,N_7046,N_5292);
or U10622 (N_10622,N_9482,N_9645);
or U10623 (N_10623,N_8981,N_7282);
and U10624 (N_10624,N_5048,N_5646);
xor U10625 (N_10625,N_9521,N_5363);
or U10626 (N_10626,N_8483,N_9526);
nor U10627 (N_10627,N_9983,N_9595);
xnor U10628 (N_10628,N_5427,N_5495);
or U10629 (N_10629,N_5786,N_6938);
nand U10630 (N_10630,N_7918,N_7395);
xnor U10631 (N_10631,N_6515,N_9680);
xnor U10632 (N_10632,N_9444,N_6956);
or U10633 (N_10633,N_6752,N_6982);
or U10634 (N_10634,N_9950,N_9324);
or U10635 (N_10635,N_5135,N_9569);
xnor U10636 (N_10636,N_9266,N_6210);
xor U10637 (N_10637,N_6462,N_8156);
and U10638 (N_10638,N_5015,N_6039);
xnor U10639 (N_10639,N_5653,N_6774);
xor U10640 (N_10640,N_8303,N_7405);
or U10641 (N_10641,N_7932,N_8983);
or U10642 (N_10642,N_8425,N_6385);
nand U10643 (N_10643,N_8049,N_9386);
or U10644 (N_10644,N_7741,N_8628);
xnor U10645 (N_10645,N_9734,N_6235);
xor U10646 (N_10646,N_8731,N_7907);
or U10647 (N_10647,N_6048,N_6320);
nand U10648 (N_10648,N_5634,N_6338);
and U10649 (N_10649,N_9071,N_6527);
nor U10650 (N_10650,N_9476,N_5295);
nand U10651 (N_10651,N_5029,N_9204);
and U10652 (N_10652,N_5144,N_8389);
or U10653 (N_10653,N_7463,N_6659);
nor U10654 (N_10654,N_7667,N_6977);
xnor U10655 (N_10655,N_5647,N_7055);
and U10656 (N_10656,N_5571,N_6000);
and U10657 (N_10657,N_7234,N_8596);
or U10658 (N_10658,N_6855,N_5044);
nand U10659 (N_10659,N_6127,N_6498);
and U10660 (N_10660,N_5943,N_9943);
and U10661 (N_10661,N_7764,N_6101);
or U10662 (N_10662,N_8820,N_8407);
xnor U10663 (N_10663,N_6770,N_7153);
or U10664 (N_10664,N_9551,N_7336);
and U10665 (N_10665,N_6463,N_8987);
and U10666 (N_10666,N_8220,N_6340);
nor U10667 (N_10667,N_6063,N_8823);
xnor U10668 (N_10668,N_5671,N_6606);
and U10669 (N_10669,N_7041,N_6743);
nand U10670 (N_10670,N_7056,N_7457);
nor U10671 (N_10671,N_9270,N_7008);
nand U10672 (N_10672,N_8247,N_7733);
xor U10673 (N_10673,N_6488,N_8514);
xnor U10674 (N_10674,N_5770,N_7952);
nand U10675 (N_10675,N_9334,N_5299);
nor U10676 (N_10676,N_5036,N_9049);
and U10677 (N_10677,N_8252,N_6867);
nand U10678 (N_10678,N_8079,N_7568);
nor U10679 (N_10679,N_9854,N_7906);
and U10680 (N_10680,N_6526,N_5246);
xnor U10681 (N_10681,N_6709,N_8488);
nor U10682 (N_10682,N_5984,N_5410);
nor U10683 (N_10683,N_8940,N_6816);
xor U10684 (N_10684,N_5316,N_7149);
nor U10685 (N_10685,N_8872,N_9156);
nand U10686 (N_10686,N_9630,N_8183);
nand U10687 (N_10687,N_7665,N_5193);
xor U10688 (N_10688,N_9799,N_8922);
nor U10689 (N_10689,N_6375,N_7389);
nor U10690 (N_10690,N_6772,N_9343);
and U10691 (N_10691,N_7864,N_7360);
or U10692 (N_10692,N_6134,N_6995);
nor U10693 (N_10693,N_8644,N_7567);
nand U10694 (N_10694,N_9875,N_5726);
nand U10695 (N_10695,N_9948,N_9433);
nand U10696 (N_10696,N_5852,N_8915);
and U10697 (N_10697,N_5620,N_9101);
xor U10698 (N_10698,N_9185,N_7427);
or U10699 (N_10699,N_7931,N_9056);
xnor U10700 (N_10700,N_9311,N_9963);
nor U10701 (N_10701,N_8403,N_7195);
and U10702 (N_10702,N_8450,N_6514);
or U10703 (N_10703,N_5763,N_5297);
nor U10704 (N_10704,N_5268,N_6366);
or U10705 (N_10705,N_6181,N_7202);
and U10706 (N_10706,N_8096,N_8601);
nor U10707 (N_10707,N_6453,N_7869);
nor U10708 (N_10708,N_9103,N_5158);
and U10709 (N_10709,N_5568,N_9748);
xor U10710 (N_10710,N_8086,N_7645);
nor U10711 (N_10711,N_8625,N_8816);
or U10712 (N_10712,N_9273,N_6819);
nand U10713 (N_10713,N_7312,N_6380);
or U10714 (N_10714,N_7713,N_7366);
nor U10715 (N_10715,N_8203,N_5489);
nor U10716 (N_10716,N_5625,N_7230);
or U10717 (N_10717,N_5614,N_5789);
xnor U10718 (N_10718,N_9504,N_9800);
nor U10719 (N_10719,N_5425,N_5873);
xor U10720 (N_10720,N_8001,N_7286);
or U10721 (N_10721,N_5406,N_9389);
nand U10722 (N_10722,N_6109,N_6490);
nor U10723 (N_10723,N_9117,N_5504);
xnor U10724 (N_10724,N_7923,N_7226);
xnor U10725 (N_10725,N_6775,N_7944);
or U10726 (N_10726,N_7397,N_8572);
nor U10727 (N_10727,N_7670,N_8936);
nand U10728 (N_10728,N_6466,N_5313);
nand U10729 (N_10729,N_7521,N_7113);
nor U10730 (N_10730,N_5454,N_9641);
or U10731 (N_10731,N_8236,N_5872);
xor U10732 (N_10732,N_7594,N_5141);
nand U10733 (N_10733,N_9807,N_6336);
nand U10734 (N_10734,N_9637,N_8121);
nor U10735 (N_10735,N_6592,N_8005);
nand U10736 (N_10736,N_7018,N_5563);
xnor U10737 (N_10737,N_7902,N_9355);
nand U10738 (N_10738,N_5288,N_8279);
xnor U10739 (N_10739,N_9442,N_9198);
or U10740 (N_10740,N_8603,N_7325);
nand U10741 (N_10741,N_5737,N_5228);
nand U10742 (N_10742,N_7631,N_6010);
nand U10743 (N_10743,N_6293,N_8580);
xnor U10744 (N_10744,N_7158,N_8751);
xor U10745 (N_10745,N_8548,N_8573);
nor U10746 (N_10746,N_6682,N_8881);
and U10747 (N_10747,N_7894,N_9926);
nand U10748 (N_10748,N_8009,N_5387);
or U10749 (N_10749,N_8949,N_6620);
nand U10750 (N_10750,N_7597,N_8352);
nand U10751 (N_10751,N_5528,N_5715);
nor U10752 (N_10752,N_6939,N_8258);
nor U10753 (N_10753,N_7221,N_5742);
or U10754 (N_10754,N_5992,N_6285);
nand U10755 (N_10755,N_6664,N_8556);
xnor U10756 (N_10756,N_8800,N_7817);
and U10757 (N_10757,N_9008,N_7592);
nand U10758 (N_10758,N_9650,N_6710);
and U10759 (N_10759,N_8228,N_6686);
xnor U10760 (N_10760,N_8338,N_5532);
or U10761 (N_10761,N_6085,N_7058);
nor U10762 (N_10762,N_9605,N_5679);
xor U10763 (N_10763,N_7857,N_6997);
or U10764 (N_10764,N_6860,N_5812);
nand U10765 (N_10765,N_6845,N_9144);
nand U10766 (N_10766,N_9007,N_8864);
and U10767 (N_10767,N_9424,N_5837);
xor U10768 (N_10768,N_7316,N_5229);
nand U10769 (N_10769,N_6954,N_8262);
xor U10770 (N_10770,N_8181,N_5923);
nor U10771 (N_10771,N_8154,N_8118);
or U10772 (N_10772,N_6836,N_6187);
and U10773 (N_10773,N_9344,N_7717);
nor U10774 (N_10774,N_8255,N_5971);
or U10775 (N_10775,N_6298,N_6638);
or U10776 (N_10776,N_6393,N_5234);
nor U10777 (N_10777,N_6582,N_6739);
nand U10778 (N_10778,N_6826,N_7732);
xnor U10779 (N_10779,N_6625,N_9918);
and U10780 (N_10780,N_9834,N_5547);
xnor U10781 (N_10781,N_9952,N_7654);
nor U10782 (N_10782,N_7477,N_5025);
nor U10783 (N_10783,N_5483,N_6731);
nand U10784 (N_10784,N_8855,N_5067);
nor U10785 (N_10785,N_8265,N_7926);
nor U10786 (N_10786,N_8701,N_5391);
xor U10787 (N_10787,N_6747,N_6879);
xnor U10788 (N_10788,N_7588,N_7550);
and U10789 (N_10789,N_7632,N_5126);
and U10790 (N_10790,N_9972,N_7270);
or U10791 (N_10791,N_5615,N_9792);
or U10792 (N_10792,N_5457,N_8810);
nand U10793 (N_10793,N_5967,N_7304);
nand U10794 (N_10794,N_5804,N_7351);
and U10795 (N_10795,N_5520,N_8431);
nor U10796 (N_10796,N_6177,N_7891);
nand U10797 (N_10797,N_5944,N_5534);
nand U10798 (N_10798,N_8231,N_5418);
nand U10799 (N_10799,N_6356,N_7424);
and U10800 (N_10800,N_8977,N_5574);
nor U10801 (N_10801,N_9129,N_6236);
xnor U10802 (N_10802,N_9985,N_7352);
xnor U10803 (N_10803,N_5607,N_9751);
or U10804 (N_10804,N_9186,N_5334);
or U10805 (N_10805,N_8254,N_9392);
xor U10806 (N_10806,N_6450,N_6850);
or U10807 (N_10807,N_6864,N_7516);
or U10808 (N_10808,N_8857,N_7414);
and U10809 (N_10809,N_8595,N_5185);
xnor U10810 (N_10810,N_8559,N_6912);
or U10811 (N_10811,N_8687,N_7228);
and U10812 (N_10812,N_7122,N_9679);
or U10813 (N_10813,N_5420,N_6120);
nand U10814 (N_10814,N_8454,N_6302);
and U10815 (N_10815,N_9074,N_9046);
and U10816 (N_10816,N_6256,N_5774);
nand U10817 (N_10817,N_6266,N_6089);
and U10818 (N_10818,N_8664,N_9653);
nand U10819 (N_10819,N_6609,N_6655);
or U10820 (N_10820,N_5621,N_7216);
nand U10821 (N_10821,N_7332,N_5781);
or U10822 (N_10822,N_5754,N_5769);
nand U10823 (N_10823,N_9754,N_9599);
nor U10824 (N_10824,N_8029,N_9544);
or U10825 (N_10825,N_7435,N_6993);
xor U10826 (N_10826,N_7969,N_9864);
xnor U10827 (N_10827,N_5072,N_5858);
and U10828 (N_10828,N_6105,N_7616);
nor U10829 (N_10829,N_6651,N_8993);
nand U10830 (N_10830,N_9897,N_5290);
nor U10831 (N_10831,N_5444,N_7557);
or U10832 (N_10832,N_8077,N_5156);
nand U10833 (N_10833,N_7112,N_9798);
xor U10834 (N_10834,N_6785,N_6571);
xnor U10835 (N_10835,N_6072,N_9811);
nand U10836 (N_10836,N_9402,N_5303);
xor U10837 (N_10837,N_9408,N_8667);
and U10838 (N_10838,N_5719,N_6902);
and U10839 (N_10839,N_6464,N_8934);
nor U10840 (N_10840,N_6451,N_5112);
or U10841 (N_10841,N_9308,N_8248);
or U10842 (N_10842,N_9313,N_7503);
or U10843 (N_10843,N_8100,N_6042);
nand U10844 (N_10844,N_8136,N_9192);
or U10845 (N_10845,N_6576,N_7785);
and U10846 (N_10846,N_6671,N_9004);
xor U10847 (N_10847,N_7867,N_9076);
xnor U10848 (N_10848,N_7057,N_9414);
nor U10849 (N_10849,N_5918,N_7845);
xor U10850 (N_10850,N_5123,N_9322);
xor U10851 (N_10851,N_8790,N_5038);
nor U10852 (N_10852,N_6405,N_7460);
xor U10853 (N_10853,N_9050,N_9467);
and U10854 (N_10854,N_5880,N_5262);
nand U10855 (N_10855,N_9822,N_5449);
nand U10856 (N_10856,N_6009,N_6781);
nor U10857 (N_10857,N_5654,N_6234);
xor U10858 (N_10858,N_6952,N_9757);
or U10859 (N_10859,N_7440,N_6529);
or U10860 (N_10860,N_8091,N_7619);
and U10861 (N_10861,N_5569,N_6123);
and U10862 (N_10862,N_8602,N_6467);
or U10863 (N_10863,N_8788,N_6061);
nand U10864 (N_10864,N_5325,N_5696);
nor U10865 (N_10865,N_9900,N_6086);
xor U10866 (N_10866,N_7273,N_8818);
nor U10867 (N_10867,N_9671,N_8510);
xnor U10868 (N_10868,N_6036,N_7072);
and U10869 (N_10869,N_9882,N_5187);
or U10870 (N_10870,N_9193,N_8159);
nand U10871 (N_10871,N_5562,N_8374);
xor U10872 (N_10872,N_8103,N_7335);
xnor U10873 (N_10873,N_8438,N_5764);
and U10874 (N_10874,N_6407,N_5644);
nand U10875 (N_10875,N_6691,N_7506);
nor U10876 (N_10876,N_8492,N_8326);
nand U10877 (N_10877,N_9069,N_7812);
and U10878 (N_10878,N_9781,N_8710);
or U10879 (N_10879,N_9134,N_5976);
nand U10880 (N_10880,N_7610,N_5821);
nor U10881 (N_10881,N_9420,N_7830);
nor U10882 (N_10882,N_5338,N_9591);
and U10883 (N_10883,N_8376,N_6726);
or U10884 (N_10884,N_9228,N_5150);
and U10885 (N_10885,N_7861,N_7795);
or U10886 (N_10886,N_6501,N_9639);
and U10887 (N_10887,N_6714,N_5013);
nand U10888 (N_10888,N_9268,N_9797);
nand U10889 (N_10889,N_5878,N_7888);
xnor U10890 (N_10890,N_9256,N_5678);
xnor U10891 (N_10891,N_6986,N_8718);
nand U10892 (N_10892,N_8635,N_9285);
and U10893 (N_10893,N_9858,N_7020);
and U10894 (N_10894,N_9901,N_5464);
nand U10895 (N_10895,N_8998,N_7250);
and U10896 (N_10896,N_9588,N_9353);
or U10897 (N_10897,N_9197,N_5698);
nand U10898 (N_10898,N_7607,N_5708);
nor U10899 (N_10899,N_8608,N_5884);
xor U10900 (N_10900,N_9380,N_5707);
nand U10901 (N_10901,N_8656,N_7766);
or U10902 (N_10902,N_5093,N_6840);
or U10903 (N_10903,N_5100,N_9644);
and U10904 (N_10904,N_8345,N_7688);
or U10905 (N_10905,N_6277,N_9003);
xor U10906 (N_10906,N_9825,N_7527);
nand U10907 (N_10907,N_6615,N_6545);
nor U10908 (N_10908,N_8799,N_8727);
xor U10909 (N_10909,N_9340,N_6610);
xnor U10910 (N_10910,N_8241,N_9241);
or U10911 (N_10911,N_6352,N_9137);
nor U10912 (N_10912,N_9061,N_7412);
and U10913 (N_10913,N_6618,N_9384);
nor U10914 (N_10914,N_8674,N_9660);
nor U10915 (N_10915,N_7989,N_8433);
and U10916 (N_10916,N_5388,N_6861);
and U10917 (N_10917,N_9184,N_7476);
nor U10918 (N_10918,N_9278,N_7972);
or U10919 (N_10919,N_5865,N_5329);
nor U10920 (N_10920,N_8942,N_5589);
xnor U10921 (N_10921,N_9902,N_7483);
nand U10922 (N_10922,N_8380,N_7406);
xnor U10923 (N_10923,N_9013,N_7404);
or U10924 (N_10924,N_5460,N_7833);
nor U10925 (N_10925,N_7602,N_7840);
nor U10926 (N_10926,N_7925,N_7168);
or U10927 (N_10927,N_9615,N_6906);
nand U10928 (N_10928,N_6147,N_5683);
xnor U10929 (N_10929,N_7788,N_5930);
nor U10930 (N_10930,N_8738,N_5331);
and U10931 (N_10931,N_9021,N_6959);
nand U10932 (N_10932,N_6962,N_8283);
nor U10933 (N_10933,N_5612,N_6522);
xor U10934 (N_10934,N_6197,N_7279);
xnor U10935 (N_10935,N_7821,N_6818);
nand U10936 (N_10936,N_6029,N_5005);
or U10937 (N_10937,N_5208,N_7034);
or U10938 (N_10938,N_8472,N_8992);
nor U10939 (N_10939,N_7890,N_9542);
or U10940 (N_10940,N_9014,N_9977);
xnor U10941 (N_10941,N_5663,N_7499);
xor U10942 (N_10942,N_5086,N_8928);
nand U10943 (N_10943,N_6588,N_9376);
nor U10944 (N_10944,N_5251,N_9065);
and U10945 (N_10945,N_5980,N_7448);
or U10946 (N_10946,N_5912,N_9974);
xor U10947 (N_10947,N_5914,N_8073);
and U10948 (N_10948,N_5416,N_8055);
and U10949 (N_10949,N_6613,N_9979);
nor U10950 (N_10950,N_5506,N_5272);
nand U10951 (N_10951,N_8560,N_8387);
xor U10952 (N_10952,N_8173,N_9239);
or U10953 (N_10953,N_5143,N_7955);
or U10954 (N_10954,N_9697,N_6756);
or U10955 (N_10955,N_7396,N_5979);
and U10956 (N_10956,N_6345,N_6647);
or U10957 (N_10957,N_9723,N_5110);
xnor U10958 (N_10958,N_6064,N_8849);
or U10959 (N_10959,N_9098,N_5999);
or U10960 (N_10960,N_5289,N_5453);
nor U10961 (N_10961,N_7963,N_8463);
or U10962 (N_10962,N_6675,N_9112);
nor U10963 (N_10963,N_7515,N_6941);
nand U10964 (N_10964,N_5018,N_6304);
or U10965 (N_10965,N_8629,N_6699);
and U10966 (N_10966,N_6940,N_9403);
or U10967 (N_10967,N_9620,N_9052);
nand U10968 (N_10968,N_9114,N_9368);
xor U10969 (N_10969,N_8523,N_8052);
nand U10970 (N_10970,N_5997,N_8208);
xor U10971 (N_10971,N_9174,N_6337);
nand U10972 (N_10972,N_7095,N_9837);
nor U10973 (N_10973,N_5045,N_6158);
xnor U10974 (N_10974,N_5365,N_9862);
nand U10975 (N_10975,N_8671,N_7986);
nand U10976 (N_10976,N_7327,N_6562);
or U10977 (N_10977,N_5315,N_8070);
or U10978 (N_10978,N_7751,N_6198);
or U10979 (N_10979,N_8975,N_5448);
or U10980 (N_10980,N_5204,N_8984);
nand U10981 (N_10981,N_9669,N_9292);
and U10982 (N_10982,N_7479,N_9116);
xnor U10983 (N_10983,N_8924,N_8191);
and U10984 (N_10984,N_7587,N_5050);
and U10985 (N_10985,N_7604,N_9921);
or U10986 (N_10986,N_7652,N_8277);
and U10987 (N_10987,N_7340,N_5705);
nand U10988 (N_10988,N_8353,N_7401);
nor U10989 (N_10989,N_5957,N_7319);
nand U10990 (N_10990,N_6552,N_5650);
nor U10991 (N_10991,N_8114,N_5949);
xor U10992 (N_10992,N_5306,N_7032);
xor U10993 (N_10993,N_5157,N_5552);
xnor U10994 (N_10994,N_5843,N_8026);
or U10995 (N_10995,N_8544,N_9893);
nor U10996 (N_10996,N_7964,N_5840);
nand U10997 (N_10997,N_6359,N_8309);
nor U10998 (N_10998,N_9584,N_8217);
xnor U10999 (N_10999,N_6730,N_6361);
xor U11000 (N_11000,N_6814,N_9323);
or U11001 (N_11001,N_7212,N_7718);
nand U11002 (N_11002,N_8041,N_7719);
nor U11003 (N_11003,N_5236,N_9138);
nor U11004 (N_11004,N_9699,N_7003);
and U11005 (N_11005,N_8260,N_5529);
nor U11006 (N_11006,N_6060,N_6204);
or U11007 (N_11007,N_9559,N_9456);
xor U11008 (N_11008,N_8929,N_6186);
nand U11009 (N_11009,N_6633,N_9055);
nand U11010 (N_11010,N_6446,N_6563);
xnor U11011 (N_11011,N_7275,N_6037);
nor U11012 (N_11012,N_8020,N_6984);
nand U11013 (N_11013,N_8108,N_9369);
xor U11014 (N_11014,N_7863,N_8650);
nor U11015 (N_11015,N_8959,N_9913);
and U11016 (N_11016,N_5893,N_9143);
or U11017 (N_11017,N_6401,N_8819);
and U11018 (N_11018,N_7924,N_6799);
or U11019 (N_11019,N_8920,N_8833);
or U11020 (N_11020,N_7851,N_6059);
and U11021 (N_11021,N_7948,N_6876);
or U11022 (N_11022,N_9448,N_8194);
or U11023 (N_11023,N_6895,N_9878);
or U11024 (N_11024,N_6286,N_6926);
nand U11025 (N_11025,N_7341,N_7053);
xor U11026 (N_11026,N_6481,N_9223);
nand U11027 (N_11027,N_6099,N_5212);
nor U11028 (N_11028,N_7990,N_9537);
xor U11029 (N_11029,N_7338,N_7781);
nor U11030 (N_11030,N_6321,N_9844);
xnor U11031 (N_11031,N_7881,N_6871);
and U11032 (N_11032,N_9717,N_9332);
xor U11033 (N_11033,N_9351,N_7141);
and U11034 (N_11034,N_6505,N_8856);
nor U11035 (N_11035,N_9026,N_9216);
nor U11036 (N_11036,N_8140,N_7941);
nand U11037 (N_11037,N_7623,N_9743);
xor U11038 (N_11038,N_6001,N_8072);
or U11039 (N_11039,N_8889,N_8104);
nand U11040 (N_11040,N_5811,N_8415);
or U11041 (N_11041,N_8179,N_8967);
or U11042 (N_11042,N_9191,N_7297);
nor U11043 (N_11043,N_5171,N_7501);
xnor U11044 (N_11044,N_6883,N_7420);
nor U11045 (N_11045,N_5533,N_6652);
xnor U11046 (N_11046,N_7039,N_6260);
or U11047 (N_11047,N_5551,N_9975);
xor U11048 (N_11048,N_8449,N_8954);
xor U11049 (N_11049,N_5054,N_5347);
nand U11050 (N_11050,N_7433,N_7510);
xor U11051 (N_11051,N_7232,N_5771);
nand U11052 (N_11052,N_8828,N_5777);
nor U11053 (N_11053,N_9887,N_9336);
xor U11054 (N_11054,N_8805,N_5346);
nor U11055 (N_11055,N_8853,N_7376);
or U11056 (N_11056,N_5934,N_7641);
xor U11057 (N_11057,N_6873,N_8422);
or U11058 (N_11058,N_5443,N_5637);
or U11059 (N_11059,N_5794,N_8600);
nand U11060 (N_11060,N_7061,N_9659);
xnor U11061 (N_11061,N_8736,N_8175);
or U11062 (N_11062,N_8973,N_7385);
nor U11063 (N_11063,N_5531,N_7611);
xnor U11064 (N_11064,N_7892,N_6367);
nand U11065 (N_11065,N_6719,N_6831);
xor U11066 (N_11066,N_7029,N_9510);
and U11067 (N_11067,N_8225,N_7644);
nand U11068 (N_11068,N_8620,N_7525);
or U11069 (N_11069,N_5544,N_8594);
or U11070 (N_11070,N_7006,N_8157);
xnor U11071 (N_11071,N_8161,N_8568);
or U11072 (N_11072,N_5617,N_9269);
and U11073 (N_11073,N_6965,N_7027);
nor U11074 (N_11074,N_9976,N_8699);
or U11075 (N_11075,N_5627,N_7235);
or U11076 (N_11076,N_8420,N_7868);
nor U11077 (N_11077,N_9478,N_9437);
and U11078 (N_11078,N_7865,N_9673);
nor U11079 (N_11079,N_6566,N_7261);
or U11080 (N_11080,N_9643,N_7590);
or U11081 (N_11081,N_8648,N_9316);
nand U11082 (N_11082,N_7017,N_9337);
nand U11083 (N_11083,N_7807,N_9169);
nor U11084 (N_11084,N_8971,N_9487);
and U11085 (N_11085,N_6521,N_5673);
xor U11086 (N_11086,N_6335,N_8905);
xor U11087 (N_11087,N_5458,N_9372);
and U11088 (N_11088,N_8529,N_8837);
xnor U11089 (N_11089,N_9124,N_5409);
and U11090 (N_11090,N_9450,N_7490);
nor U11091 (N_11091,N_5162,N_5882);
nor U11092 (N_11092,N_5985,N_8423);
nor U11093 (N_11093,N_6049,N_5500);
nand U11094 (N_11094,N_8712,N_5343);
nand U11095 (N_11095,N_9596,N_5127);
nand U11096 (N_11096,N_6875,N_8050);
or U11097 (N_11097,N_8899,N_7455);
and U11098 (N_11098,N_5057,N_6688);
and U11099 (N_11099,N_6630,N_5658);
xnor U11100 (N_11100,N_9656,N_9397);
or U11101 (N_11101,N_9617,N_7045);
nand U11102 (N_11102,N_5595,N_9104);
nor U11103 (N_11103,N_6800,N_7321);
xnor U11104 (N_11104,N_8526,N_5560);
nor U11105 (N_11105,N_7126,N_7012);
or U11106 (N_11106,N_5990,N_8696);
nand U11107 (N_11107,N_6113,N_6642);
nor U11108 (N_11108,N_6915,N_6247);
nand U11109 (N_11109,N_6896,N_8370);
or U11110 (N_11110,N_7175,N_6600);
xnor U11111 (N_11111,N_7533,N_7411);
or U11112 (N_11112,N_6006,N_9874);
xnor U11113 (N_11113,N_9088,N_7444);
and U11114 (N_11114,N_6411,N_8485);
nor U11115 (N_11115,N_9783,N_5838);
xnor U11116 (N_11116,N_9080,N_8623);
xnor U11117 (N_11117,N_7913,N_8015);
xnor U11118 (N_11118,N_8297,N_8033);
nor U11119 (N_11119,N_5183,N_9574);
nand U11120 (N_11120,N_8520,N_8563);
or U11121 (N_11121,N_5854,N_6870);
nor U11122 (N_11122,N_8770,N_8848);
nand U11123 (N_11123,N_6159,N_9534);
and U11124 (N_11124,N_6209,N_6643);
nand U11125 (N_11125,N_6722,N_7109);
and U11126 (N_11126,N_7390,N_5802);
nor U11127 (N_11127,N_5825,N_9965);
nor U11128 (N_11128,N_8263,N_8642);
nand U11129 (N_11129,N_6283,N_7938);
and U11130 (N_11130,N_8487,N_9364);
nor U11131 (N_11131,N_7258,N_7064);
or U11132 (N_11132,N_5441,N_7459);
nand U11133 (N_11133,N_6725,N_5328);
nand U11134 (N_11134,N_7458,N_7409);
or U11135 (N_11135,N_8207,N_6351);
xor U11136 (N_11136,N_9301,N_7104);
nand U11137 (N_11137,N_9374,N_9404);
and U11138 (N_11138,N_9625,N_9843);
and U11139 (N_11139,N_6947,N_6882);
or U11140 (N_11140,N_6102,N_8634);
nor U11141 (N_11141,N_9141,N_7831);
and U11142 (N_11142,N_9847,N_5384);
xnor U11143 (N_11143,N_6539,N_5536);
xnor U11144 (N_11144,N_7609,N_8989);
nand U11145 (N_11145,N_8493,N_5920);
nor U11146 (N_11146,N_6420,N_9439);
or U11147 (N_11147,N_5291,N_7313);
nor U11148 (N_11148,N_7303,N_7689);
nand U11149 (N_11149,N_6949,N_5631);
and U11150 (N_11150,N_6097,N_7023);
xor U11151 (N_11151,N_9704,N_6043);
xor U11152 (N_11152,N_6729,N_7878);
or U11153 (N_11153,N_9319,N_5487);
xnor U11154 (N_11154,N_9396,N_7363);
or U11155 (N_11155,N_6032,N_7491);
nor U11156 (N_11156,N_6603,N_5053);
or U11157 (N_11157,N_9791,N_7475);
nor U11158 (N_11158,N_7993,N_7323);
xor U11159 (N_11159,N_9773,N_8812);
nor U11160 (N_11160,N_7816,N_9133);
and U11161 (N_11161,N_8367,N_9271);
nor U11162 (N_11162,N_5948,N_6025);
or U11163 (N_11163,N_8170,N_9642);
nor U11164 (N_11164,N_6717,N_5359);
nor U11165 (N_11165,N_6544,N_5577);
and U11166 (N_11166,N_6325,N_6008);
xnor U11167 (N_11167,N_7704,N_7161);
or U11168 (N_11168,N_6011,N_7302);
xor U11169 (N_11169,N_6254,N_8566);
and U11170 (N_11170,N_8877,N_6754);
xor U11171 (N_11171,N_9820,N_9571);
and U11172 (N_11172,N_7049,N_6144);
or U11173 (N_11173,N_9788,N_7825);
nor U11174 (N_11174,N_6200,N_8661);
nor U11175 (N_11175,N_6313,N_6054);
or U11176 (N_11176,N_9029,N_9978);
nor U11177 (N_11177,N_7422,N_9894);
xor U11178 (N_11178,N_6822,N_9616);
xor U11179 (N_11179,N_8090,N_5000);
xnor U11180 (N_11180,N_5264,N_5374);
nand U11181 (N_11181,N_5255,N_9600);
xor U11182 (N_11182,N_9840,N_8317);
nor U11183 (N_11183,N_8404,N_5721);
nand U11184 (N_11184,N_6150,N_5469);
nand U11185 (N_11185,N_5795,N_7756);
and U11186 (N_11186,N_9210,N_7305);
nand U11187 (N_11187,N_8898,N_8528);
xnor U11188 (N_11188,N_7353,N_6080);
and U11189 (N_11189,N_6594,N_5989);
nand U11190 (N_11190,N_9000,N_5145);
and U11191 (N_11191,N_9363,N_8322);
or U11192 (N_11192,N_6245,N_9933);
and U11193 (N_11193,N_8169,N_7249);
nor U11194 (N_11194,N_9922,N_9701);
nand U11195 (N_11195,N_7712,N_6833);
xor U11196 (N_11196,N_8062,N_7933);
nand U11197 (N_11197,N_5392,N_7154);
or U11198 (N_11198,N_5218,N_5132);
nand U11199 (N_11199,N_6689,N_8622);
or U11200 (N_11200,N_5507,N_7914);
or U11201 (N_11201,N_9610,N_9177);
nand U11202 (N_11202,N_9128,N_8382);
nand U11203 (N_11203,N_7545,N_7887);
xnor U11204 (N_11204,N_9934,N_8680);
nand U11205 (N_11205,N_6636,N_9655);
and U11206 (N_11206,N_5466,N_7077);
nor U11207 (N_11207,N_7107,N_7803);
nor U11208 (N_11208,N_6788,N_6485);
xnor U11209 (N_11209,N_7940,N_5857);
and U11210 (N_11210,N_8172,N_7083);
nand U11211 (N_11211,N_9237,N_7453);
and U11212 (N_11212,N_6106,N_5151);
or U11213 (N_11213,N_8578,N_7774);
and U11214 (N_11214,N_5609,N_7798);
nand U11215 (N_11215,N_7081,N_6598);
nor U11216 (N_11216,N_5780,N_7200);
and U11217 (N_11217,N_6662,N_9768);
or U11218 (N_11218,N_5163,N_5172);
or U11219 (N_11219,N_9647,N_6138);
xor U11220 (N_11220,N_5241,N_5776);
nand U11221 (N_11221,N_5730,N_7765);
or U11222 (N_11222,N_6798,N_5600);
and U11223 (N_11223,N_6480,N_8137);
xnor U11224 (N_11224,N_8147,N_6443);
or U11225 (N_11225,N_8184,N_8587);
xor U11226 (N_11226,N_7129,N_9779);
xnor U11227 (N_11227,N_5358,N_5889);
or U11228 (N_11228,N_7739,N_9009);
nand U11229 (N_11229,N_9598,N_8085);
and U11230 (N_11230,N_7330,N_7134);
and U11231 (N_11231,N_9891,N_5747);
or U11232 (N_11232,N_7900,N_5007);
and U11233 (N_11233,N_6981,N_9064);
nand U11234 (N_11234,N_8771,N_8083);
and U11235 (N_11235,N_5866,N_5964);
or U11236 (N_11236,N_5901,N_8088);
or U11237 (N_11237,N_7159,N_7388);
or U11238 (N_11238,N_6052,N_5686);
or U11239 (N_11239,N_5357,N_7382);
xor U11240 (N_11240,N_9249,N_5538);
nand U11241 (N_11241,N_8160,N_8589);
xnor U11242 (N_11242,N_5414,N_8410);
and U11243 (N_11243,N_7152,N_8814);
xor U11244 (N_11244,N_8115,N_9012);
or U11245 (N_11245,N_7520,N_6767);
nor U11246 (N_11246,N_8227,N_6415);
nand U11247 (N_11247,N_7253,N_7676);
xnor U11248 (N_11248,N_6378,N_8609);
nand U11249 (N_11249,N_9025,N_8192);
xnor U11250 (N_11250,N_7560,N_6067);
nor U11251 (N_11251,N_7091,N_6456);
and U11252 (N_11252,N_5829,N_5472);
xnor U11253 (N_11253,N_5511,N_6021);
nand U11254 (N_11254,N_7727,N_8240);
or U11255 (N_11255,N_5570,N_9346);
xor U11256 (N_11256,N_5210,N_6280);
nand U11257 (N_11257,N_7150,N_5497);
and U11258 (N_11258,N_9690,N_9314);
or U11259 (N_11259,N_7927,N_7024);
and U11260 (N_11260,N_7723,N_9705);
or U11261 (N_11261,N_6222,N_9224);
xor U11262 (N_11262,N_6093,N_9753);
and U11263 (N_11263,N_6680,N_6346);
and U11264 (N_11264,N_8637,N_8982);
or U11265 (N_11265,N_7958,N_9272);
nor U11266 (N_11266,N_6189,N_5630);
xnor U11267 (N_11267,N_8152,N_5791);
or U11268 (N_11268,N_8437,N_8110);
or U11269 (N_11269,N_8835,N_8466);
and U11270 (N_11270,N_6071,N_7981);
nor U11271 (N_11271,N_7624,N_5704);
xor U11272 (N_11272,N_9412,N_7549);
nor U11273 (N_11273,N_8986,N_5198);
nand U11274 (N_11274,N_6358,N_9801);
nand U11275 (N_11275,N_7743,N_5022);
and U11276 (N_11276,N_5337,N_5555);
xnor U11277 (N_11277,N_7885,N_9503);
and U11278 (N_11278,N_8125,N_6437);
or U11279 (N_11279,N_5090,N_9712);
or U11280 (N_11280,N_6913,N_7782);
nor U11281 (N_11281,N_7874,N_9803);
nand U11282 (N_11282,N_7237,N_5471);
and U11283 (N_11283,N_5398,N_7722);
nor U11284 (N_11284,N_8880,N_8753);
xor U11285 (N_11285,N_7544,N_5741);
xor U11286 (N_11286,N_6827,N_6715);
or U11287 (N_11287,N_9411,N_8278);
nor U11288 (N_11288,N_7848,N_7937);
xnor U11289 (N_11289,N_5435,N_7450);
nand U11290 (N_11290,N_9455,N_6843);
and U11291 (N_11291,N_7163,N_6027);
or U11292 (N_11292,N_7183,N_6435);
nor U11293 (N_11293,N_7248,N_8702);
or U11294 (N_11294,N_9778,N_8530);
or U11295 (N_11295,N_8561,N_7078);
nand U11296 (N_11296,N_8917,N_5192);
nand U11297 (N_11297,N_8582,N_8717);
or U11298 (N_11298,N_6026,N_9519);
xnor U11299 (N_11299,N_6471,N_5401);
and U11300 (N_11300,N_9884,N_7715);
or U11301 (N_11301,N_5567,N_6173);
nand U11302 (N_11302,N_9790,N_8428);
and U11303 (N_11303,N_6398,N_7188);
and U11304 (N_11304,N_5991,N_8737);
and U11305 (N_11305,N_9298,N_6933);
nor U11306 (N_11306,N_5899,N_6013);
or U11307 (N_11307,N_8063,N_5222);
xor U11308 (N_11308,N_8133,N_9490);
xor U11309 (N_11309,N_9296,N_5182);
nor U11310 (N_11310,N_6556,N_5660);
and U11311 (N_11311,N_5909,N_5870);
xnor U11312 (N_11312,N_8235,N_9609);
xor U11313 (N_11313,N_6960,N_6866);
and U11314 (N_11314,N_7875,N_6665);
nor U11315 (N_11315,N_9804,N_7403);
and U11316 (N_11316,N_8583,N_5323);
nor U11317 (N_11317,N_5806,N_7116);
nor U11318 (N_11318,N_9350,N_8144);
and U11319 (N_11319,N_9614,N_6992);
nor U11320 (N_11320,N_9662,N_9305);
nand U11321 (N_11321,N_9681,N_6961);
nand U11322 (N_11322,N_8668,N_5966);
and U11323 (N_11323,N_7883,N_5736);
or U11324 (N_11324,N_6056,N_6002);
nand U11325 (N_11325,N_6051,N_9132);
or U11326 (N_11326,N_7994,N_6793);
xor U11327 (N_11327,N_9741,N_8394);
and U11328 (N_11328,N_9387,N_6214);
nor U11329 (N_11329,N_8460,N_8123);
or U11330 (N_11330,N_6945,N_9035);
or U11331 (N_11331,N_7600,N_7574);
and U11332 (N_11332,N_7377,N_6605);
nor U11333 (N_11333,N_6718,N_7118);
nor U11334 (N_11334,N_6278,N_8512);
or U11335 (N_11335,N_8261,N_7127);
nor U11336 (N_11336,N_8355,N_9492);
nor U11337 (N_11337,N_6110,N_6354);
nor U11338 (N_11338,N_9425,N_5355);
nor U11339 (N_11339,N_5766,N_6570);
nand U11340 (N_11340,N_9839,N_8613);
xnor U11341 (N_11341,N_7391,N_9280);
nor U11342 (N_11342,N_8054,N_9018);
nor U11343 (N_11343,N_6188,N_8002);
or U11344 (N_11344,N_6974,N_7368);
and U11345 (N_11345,N_6769,N_8174);
nor U11346 (N_11346,N_5919,N_5226);
or U11347 (N_11347,N_5910,N_5846);
or U11348 (N_11348,N_5302,N_8249);
or U11349 (N_11349,N_6084,N_8366);
nand U11350 (N_11350,N_7617,N_7953);
and U11351 (N_11351,N_5685,N_9195);
xor U11352 (N_11352,N_9899,N_9017);
xor U11353 (N_11353,N_7915,N_5894);
xor U11354 (N_11354,N_8761,N_7025);
or U11355 (N_11355,N_9856,N_5213);
nand U11356 (N_11356,N_9524,N_9330);
nor U11357 (N_11357,N_6881,N_7208);
or U11358 (N_11358,N_5808,N_6327);
xnor U11359 (N_11359,N_5450,N_6865);
xnor U11360 (N_11360,N_7946,N_7950);
nor U11361 (N_11361,N_8888,N_5017);
nor U11362 (N_11362,N_8149,N_8795);
xor U11363 (N_11363,N_9604,N_7022);
xnor U11364 (N_11364,N_8543,N_5439);
nand U11365 (N_11365,N_7531,N_8707);
nand U11366 (N_11366,N_6795,N_5170);
and U11367 (N_11367,N_9683,N_5580);
and U11368 (N_11368,N_5632,N_6549);
xor U11369 (N_11369,N_8590,N_9608);
xor U11370 (N_11370,N_8655,N_9099);
nor U11371 (N_11371,N_6886,N_7523);
nand U11372 (N_11372,N_7398,N_6972);
or U11373 (N_11373,N_8627,N_7535);
nor U11374 (N_11374,N_6825,N_5935);
xor U11375 (N_11375,N_8321,N_5166);
nor U11376 (N_11376,N_9577,N_5734);
nor U11377 (N_11377,N_8019,N_8245);
nand U11378 (N_11378,N_8011,N_6172);
or U11379 (N_11379,N_5404,N_6439);
or U11380 (N_11380,N_6096,N_6746);
xnor U11381 (N_11381,N_9472,N_6716);
and U11382 (N_11382,N_5760,N_8963);
nor U11383 (N_11383,N_7005,N_8039);
or U11384 (N_11384,N_8378,N_8879);
nor U11385 (N_11385,N_8490,N_5694);
or U11386 (N_11386,N_9960,N_7446);
or U11387 (N_11387,N_7075,N_5656);
or U11388 (N_11388,N_7513,N_6914);
and U11389 (N_11389,N_7494,N_7633);
or U11390 (N_11390,N_6473,N_8109);
nand U11391 (N_11391,N_6143,N_6757);
nand U11392 (N_11392,N_9987,N_5205);
xor U11393 (N_11393,N_8268,N_6645);
xor U11394 (N_11394,N_5133,N_6511);
or U11395 (N_11395,N_7291,N_7539);
nand U11396 (N_11396,N_7434,N_7471);
nor U11397 (N_11397,N_9164,N_8372);
xnor U11398 (N_11398,N_6648,N_8189);
nor U11399 (N_11399,N_5765,N_6003);
nor U11400 (N_11400,N_7276,N_6856);
and U11401 (N_11401,N_6402,N_9159);
and U11402 (N_11402,N_8038,N_9805);
nor U11403 (N_11403,N_5267,N_9552);
nor U11404 (N_11404,N_6821,N_5512);
and U11405 (N_11405,N_9030,N_8346);
nor U11406 (N_11406,N_5665,N_6203);
or U11407 (N_11407,N_6342,N_5651);
or U11408 (N_11408,N_5402,N_7086);
nand U11409 (N_11409,N_7677,N_8427);
xnor U11410 (N_11410,N_8497,N_7090);
nand U11411 (N_11411,N_6255,N_7178);
nand U11412 (N_11412,N_7755,N_6015);
or U11413 (N_11413,N_7485,N_8168);
and U11414 (N_11414,N_6195,N_8747);
or U11415 (N_11415,N_7466,N_7285);
nand U11416 (N_11416,N_6572,N_7970);
xor U11417 (N_11417,N_6221,N_9212);
and U11418 (N_11418,N_8482,N_7238);
and U11419 (N_11419,N_6852,N_5693);
and U11420 (N_11420,N_6041,N_8285);
and U11421 (N_11421,N_6363,N_5446);
nor U11422 (N_11422,N_7773,N_7905);
nor U11423 (N_11423,N_9005,N_8440);
xor U11424 (N_11424,N_5103,N_8419);
or U11425 (N_11425,N_7135,N_9877);
xor U11426 (N_11426,N_9747,N_7814);
nand U11427 (N_11427,N_7470,N_8432);
xnor U11428 (N_11428,N_6848,N_8907);
and U11429 (N_11429,N_5117,N_5317);
xor U11430 (N_11430,N_5805,N_8163);
nor U11431 (N_11431,N_6454,N_5408);
nand U11432 (N_11432,N_8295,N_7210);
and U11433 (N_11433,N_5963,N_9525);
xnor U11434 (N_11434,N_9070,N_8614);
nand U11435 (N_11435,N_6146,N_5689);
and U11436 (N_11436,N_5809,N_6403);
xor U11437 (N_11437,N_7373,N_8887);
or U11438 (N_11438,N_8045,N_8873);
nor U11439 (N_11439,N_9549,N_8298);
nand U11440 (N_11440,N_7660,N_9646);
xor U11441 (N_11441,N_8224,N_9528);
xnor U11442 (N_11442,N_7992,N_6240);
nor U11443 (N_11443,N_9736,N_9707);
or U11444 (N_11444,N_9441,N_9870);
xnor U11445 (N_11445,N_7241,N_9291);
and U11446 (N_11446,N_9255,N_5232);
nand U11447 (N_11447,N_6053,N_7225);
or U11448 (N_11448,N_5279,N_6296);
or U11449 (N_11449,N_8469,N_6458);
nor U11450 (N_11450,N_9738,N_6894);
xnor U11451 (N_11451,N_8287,N_8206);
or U11452 (N_11452,N_7956,N_8518);
nand U11453 (N_11453,N_7982,N_9157);
nand U11454 (N_11454,N_5403,N_9865);
or U11455 (N_11455,N_7067,N_6291);
or U11456 (N_11456,N_5095,N_5558);
xor U11457 (N_11457,N_8111,N_8797);
nand U11458 (N_11458,N_9661,N_9998);
nor U11459 (N_11459,N_7146,N_6970);
nor U11460 (N_11460,N_6585,N_9980);
nand U11461 (N_11461,N_9827,N_6125);
and U11462 (N_11462,N_6516,N_6503);
nand U11463 (N_11463,N_8685,N_9073);
nor U11464 (N_11464,N_8930,N_6119);
nand U11465 (N_11465,N_6284,N_9016);
or U11466 (N_11466,N_7445,N_5586);
or U11467 (N_11467,N_9802,N_7454);
nor U11468 (N_11468,N_7855,N_7089);
xor U11469 (N_11469,N_5300,N_9873);
nor U11470 (N_11470,N_6314,N_7004);
xor U11471 (N_11471,N_9463,N_6787);
or U11472 (N_11472,N_7133,N_9100);
xor U11473 (N_11473,N_6934,N_8202);
and U11474 (N_11474,N_6258,N_9460);
and U11475 (N_11475,N_6696,N_9912);
xor U11476 (N_11476,N_6802,N_8755);
nor U11477 (N_11477,N_7639,N_7218);
nor U11478 (N_11478,N_9886,N_8725);
nand U11479 (N_11479,N_6413,N_9572);
and U11480 (N_11480,N_8212,N_5030);
and U11481 (N_11481,N_9769,N_7419);
xnor U11482 (N_11482,N_5260,N_8703);
or U11483 (N_11483,N_8128,N_5510);
or U11484 (N_11484,N_9555,N_8669);
nor U11485 (N_11485,N_6212,N_6553);
or U11486 (N_11486,N_8273,N_7784);
and U11487 (N_11487,N_9440,N_8242);
xnor U11488 (N_11488,N_9115,N_5056);
xnor U11489 (N_11489,N_7284,N_7073);
nand U11490 (N_11490,N_8555,N_9727);
xnor U11491 (N_11491,N_5712,N_6168);
and U11492 (N_11492,N_8533,N_6755);
nor U11493 (N_11493,N_5584,N_9221);
xor U11494 (N_11494,N_9039,N_5380);
xnor U11495 (N_11495,N_9706,N_8990);
xnor U11496 (N_11496,N_5739,N_9501);
and U11497 (N_11497,N_8732,N_8031);
nor U11498 (N_11498,N_8946,N_7423);
xor U11499 (N_11499,N_5818,N_9136);
and U11500 (N_11500,N_9430,N_8409);
nand U11501 (N_11501,N_8480,N_8911);
and U11502 (N_11502,N_7512,N_6163);
nor U11503 (N_11503,N_7242,N_7621);
xor U11504 (N_11504,N_5938,N_8158);
nor U11505 (N_11505,N_7280,N_8151);
nor U11506 (N_11506,N_5475,N_9232);
xnor U11507 (N_11507,N_7384,N_5367);
or U11508 (N_11508,N_6227,N_9276);
or U11509 (N_11509,N_6331,N_9982);
nor U11510 (N_11510,N_9234,N_6297);
or U11511 (N_11511,N_8803,N_9179);
or U11512 (N_11512,N_7348,N_9367);
and U11513 (N_11513,N_7511,N_6983);
nand U11514 (N_11514,N_7829,N_9227);
nand U11515 (N_11515,N_5206,N_5429);
xor U11516 (N_11516,N_9557,N_8276);
nor U11517 (N_11517,N_6807,N_9842);
nor U11518 (N_11518,N_8638,N_7746);
nand U11519 (N_11519,N_6604,N_7706);
or U11520 (N_11520,N_8458,N_9168);
nand U11521 (N_11521,N_8381,N_7775);
or U11522 (N_11522,N_5089,N_7359);
or U11523 (N_11523,N_8253,N_7311);
or U11524 (N_11524,N_8571,N_6199);
nand U11525 (N_11525,N_9499,N_5176);
xnor U11526 (N_11526,N_6016,N_6184);
nand U11527 (N_11527,N_5688,N_8406);
nor U11528 (N_11528,N_5012,N_9258);
xor U11529 (N_11529,N_8442,N_5047);
xor U11530 (N_11530,N_7872,N_7694);
xnor U11531 (N_11531,N_7771,N_9658);
nor U11532 (N_11532,N_9733,N_5216);
or U11533 (N_11533,N_9626,N_5352);
nor U11534 (N_11534,N_5349,N_7465);
or U11535 (N_11535,N_8564,N_5140);
nand U11536 (N_11536,N_7244,N_9541);
xnor U11537 (N_11537,N_8605,N_9173);
xor U11538 (N_11538,N_5725,N_6115);
or U11539 (N_11539,N_5330,N_8906);
nand U11540 (N_11540,N_6660,N_9041);
and U11541 (N_11541,N_6020,N_8418);
xnor U11542 (N_11542,N_8023,N_7307);
xnor U11543 (N_11543,N_6597,N_7263);
and U11544 (N_11544,N_9302,N_6640);
xnor U11545 (N_11545,N_9749,N_8779);
and U11546 (N_11546,N_6622,N_8320);
or U11547 (N_11547,N_9480,N_7630);
nand U11548 (N_11548,N_7407,N_5102);
and U11549 (N_11549,N_7720,N_6551);
and U11550 (N_11550,N_7543,N_8567);
xor U11551 (N_11551,N_8513,N_9381);
and U11552 (N_11552,N_7013,N_9728);
nor U11553 (N_11553,N_7099,N_6305);
or U11554 (N_11554,N_6343,N_7292);
and U11555 (N_11555,N_6654,N_9106);
and U11556 (N_11556,N_9603,N_9942);
nand U11557 (N_11557,N_6124,N_7716);
xor U11558 (N_11558,N_5283,N_8150);
xnor U11559 (N_11559,N_7416,N_9938);
nor U11560 (N_11560,N_8885,N_5779);
nor U11561 (N_11561,N_5046,N_7593);
nor U11562 (N_11562,N_5537,N_9761);
nor U11563 (N_11563,N_8813,N_9896);
and U11564 (N_11564,N_9845,N_6251);
or U11565 (N_11565,N_9470,N_7596);
or U11566 (N_11566,N_7893,N_9700);
and U11567 (N_11567,N_9435,N_8430);
nor U11568 (N_11568,N_8976,N_6791);
and U11569 (N_11569,N_7692,N_6683);
nand U11570 (N_11570,N_7174,N_8286);
xor U11571 (N_11571,N_7606,N_9967);
nand U11572 (N_11572,N_8196,N_6220);
and U11573 (N_11573,N_7251,N_8621);
and U11574 (N_11574,N_7199,N_8182);
and U11575 (N_11575,N_9497,N_7921);
and U11576 (N_11576,N_6087,N_6377);
nor U11577 (N_11577,N_6824,N_5091);
or U11578 (N_11578,N_9992,N_6555);
nand U11579 (N_11579,N_8796,N_6862);
nor U11580 (N_11580,N_7002,N_8426);
nand U11581 (N_11581,N_5970,N_9780);
or U11582 (N_11582,N_8363,N_6589);
xor U11583 (N_11583,N_6520,N_8776);
nor U11584 (N_11584,N_5111,N_5669);
and U11585 (N_11585,N_7871,N_8504);
and U11586 (N_11586,N_9158,N_7296);
nor U11587 (N_11587,N_5196,N_7137);
nand U11588 (N_11588,N_7638,N_6532);
or U11589 (N_11589,N_8713,N_7464);
xor U11590 (N_11590,N_8271,N_7828);
xor U11591 (N_11591,N_7295,N_8012);
or U11592 (N_11592,N_6182,N_8024);
nand U11593 (N_11593,N_7033,N_5281);
xor U11594 (N_11594,N_9592,N_6103);
or U11595 (N_11595,N_6841,N_6427);
or U11596 (N_11596,N_8508,N_8013);
nand U11597 (N_11597,N_7841,N_6117);
nor U11598 (N_11598,N_5605,N_7197);
xnor U11599 (N_11599,N_8473,N_9326);
or U11600 (N_11600,N_7038,N_5122);
and U11601 (N_11601,N_8709,N_8890);
xor U11602 (N_11602,N_7772,N_6133);
and U11603 (N_11603,N_7334,N_5447);
nor U11604 (N_11604,N_5674,N_6357);
xor U11605 (N_11605,N_7662,N_6104);
nand U11606 (N_11606,N_9675,N_7839);
or U11607 (N_11607,N_5075,N_6370);
or U11608 (N_11608,N_9691,N_8741);
nand U11609 (N_11609,N_9113,N_7324);
or U11610 (N_11610,N_9247,N_6269);
nor U11611 (N_11611,N_6399,N_6142);
and U11612 (N_11612,N_7306,N_8723);
nand U11613 (N_11613,N_8511,N_9606);
nor U11614 (N_11614,N_5619,N_6238);
and U11615 (N_11615,N_9459,N_9225);
xnor U11616 (N_11616,N_7252,N_5593);
or U11617 (N_11617,N_8730,N_6396);
or U11618 (N_11618,N_5256,N_8745);
nor U11619 (N_11619,N_6761,N_6476);
nand U11620 (N_11620,N_9418,N_7650);
nand U11621 (N_11621,N_5905,N_6175);
or U11622 (N_11622,N_7747,N_8839);
and U11623 (N_11623,N_8610,N_7961);
nand U11624 (N_11624,N_8547,N_6768);
nand U11625 (N_11625,N_8562,N_9861);
and U11626 (N_11626,N_7951,N_9824);
nor U11627 (N_11627,N_8720,N_7019);
nor U11628 (N_11628,N_5596,N_5635);
and U11629 (N_11629,N_5626,N_8371);
nand U11630 (N_11630,N_5824,N_8535);
nor U11631 (N_11631,N_6426,N_6932);
xor U11632 (N_11632,N_9075,N_5230);
nor U11633 (N_11633,N_5211,N_5058);
and U11634 (N_11634,N_6765,N_5691);
nor U11635 (N_11635,N_6523,N_6681);
xor U11636 (N_11636,N_5109,N_5800);
xnor U11637 (N_11637,N_7436,N_7274);
and U11638 (N_11638,N_7889,N_5898);
xor U11639 (N_11639,N_5968,N_7949);
nor U11640 (N_11640,N_5010,N_7977);
and U11641 (N_11641,N_5032,N_5743);
xor U11642 (N_11642,N_5296,N_8340);
or U11643 (N_11643,N_8453,N_6581);
nor U11644 (N_11644,N_6750,N_6978);
and U11645 (N_11645,N_6160,N_9782);
nand U11646 (N_11646,N_9259,N_8354);
nor U11647 (N_11647,N_9222,N_7862);
and U11648 (N_11648,N_9808,N_8925);
nand U11649 (N_11649,N_7079,N_9561);
xor U11650 (N_11650,N_5360,N_7754);
nand U11651 (N_11651,N_7132,N_6482);
nand U11652 (N_11652,N_7439,N_9994);
or U11653 (N_11653,N_7612,N_5344);
or U11654 (N_11654,N_8102,N_5191);
nor U11655 (N_11655,N_6542,N_9935);
xnor U11656 (N_11656,N_6537,N_7991);
or U11657 (N_11657,N_6929,N_9218);
or U11658 (N_11658,N_7672,N_6290);
xnor U11659 (N_11659,N_8691,N_6282);
and U11660 (N_11660,N_6044,N_5813);
nor U11661 (N_11661,N_8950,N_6194);
xnor U11662 (N_11662,N_8368,N_8288);
and U11663 (N_11663,N_8626,N_8481);
or U11664 (N_11664,N_5542,N_7734);
or U11665 (N_11665,N_9737,N_8257);
or U11666 (N_11666,N_5348,N_7804);
nor U11667 (N_11667,N_6738,N_6132);
nand U11668 (N_11668,N_9286,N_5379);
nor U11669 (N_11669,N_7425,N_9920);
or U11670 (N_11670,N_8748,N_9787);
nand U11671 (N_11671,N_5745,N_9793);
nand U11672 (N_11672,N_7185,N_6019);
or U11673 (N_11673,N_8293,N_6068);
or U11674 (N_11674,N_5003,N_9250);
nand U11675 (N_11675,N_9127,N_7059);
and U11676 (N_11676,N_5788,N_8831);
or U11677 (N_11677,N_9339,N_8211);
nand U11678 (N_11678,N_6441,N_5639);
or U11679 (N_11679,N_5393,N_6704);
nand U11680 (N_11680,N_9462,N_6275);
nand U11681 (N_11681,N_9495,N_8636);
and U11682 (N_11682,N_6038,N_9312);
or U11683 (N_11683,N_6231,N_9590);
and U11684 (N_11684,N_6639,N_5682);
or U11685 (N_11685,N_6412,N_9589);
or U11686 (N_11686,N_5937,N_6712);
and U11687 (N_11687,N_8411,N_5961);
nor U11688 (N_11688,N_5377,N_8503);
nor U11689 (N_11689,N_5424,N_9077);
nor U11690 (N_11690,N_6900,N_6744);
nand U11691 (N_11691,N_7011,N_6946);
nand U11692 (N_11692,N_8307,N_8344);
nand U11693 (N_11693,N_7726,N_5907);
nor U11694 (N_11694,N_9857,N_8953);
and U11695 (N_11695,N_9181,N_6434);
xor U11696 (N_11696,N_8859,N_8937);
and U11697 (N_11697,N_5470,N_5396);
xnor U11698 (N_11698,N_6927,N_6438);
or U11699 (N_11699,N_9147,N_9871);
nand U11700 (N_11700,N_6292,N_9019);
xnor U11701 (N_11701,N_6667,N_8065);
and U11702 (N_11702,N_5928,N_9233);
nand U11703 (N_11703,N_5994,N_9581);
and U11704 (N_11704,N_5118,N_5463);
nand U11705 (N_11705,N_7934,N_7595);
nor U11706 (N_11706,N_9685,N_8177);
xnor U11707 (N_11707,N_6268,N_9970);
nor U11708 (N_11708,N_9388,N_6513);
nor U11709 (N_11709,N_5130,N_7047);
xor U11710 (N_11710,N_7827,N_6748);
or U11711 (N_11711,N_8413,N_5602);
nor U11712 (N_11712,N_7207,N_7060);
nand U11713 (N_11713,N_5491,N_8759);
nor U11714 (N_11714,N_5711,N_9347);
xor U11715 (N_11715,N_7257,N_7495);
nand U11716 (N_11716,N_5814,N_7691);
xor U11717 (N_11717,N_8124,N_8806);
nor U11718 (N_11718,N_8101,N_7834);
and U11719 (N_11719,N_7050,N_5253);
or U11720 (N_11720,N_9151,N_5340);
or U11721 (N_11721,N_9413,N_5146);
xnor U11722 (N_11722,N_6365,N_7217);
or U11723 (N_11723,N_5523,N_7381);
nand U11724 (N_11724,N_9632,N_5336);
nand U11725 (N_11725,N_6317,N_7901);
nor U11726 (N_11726,N_8517,N_6936);
xor U11727 (N_11727,N_8704,N_7735);
or U11728 (N_11728,N_5700,N_8617);
nor U11729 (N_11729,N_5699,N_6339);
nand U11730 (N_11730,N_7191,N_6510);
nand U11731 (N_11731,N_6812,N_6808);
nor U11732 (N_11732,N_9335,N_8097);
nor U11733 (N_11733,N_6499,N_9034);
or U11734 (N_11734,N_8325,N_5822);
nor U11735 (N_11735,N_6007,N_6909);
and U11736 (N_11736,N_8597,N_7421);
nand U11737 (N_11737,N_6219,N_7068);
and U11738 (N_11738,N_6955,N_9722);
and U11739 (N_11739,N_9409,N_6616);
nand U11740 (N_11740,N_9213,N_6985);
nand U11741 (N_11741,N_6701,N_5661);
nand U11742 (N_11742,N_6475,N_5035);
nand U11743 (N_11743,N_8784,N_8291);
and U11744 (N_11744,N_7380,N_8489);
xnor U11745 (N_11745,N_9031,N_5856);
and U11746 (N_11746,N_9443,N_6379);
and U11747 (N_11747,N_6533,N_7971);
xor U11748 (N_11748,N_5640,N_7880);
or U11749 (N_11749,N_6854,N_8750);
and U11750 (N_11750,N_8783,N_6623);
nor U11751 (N_11751,N_9341,N_9378);
or U11752 (N_11752,N_9973,N_9477);
nand U11753 (N_11753,N_6780,N_5871);
nand U11754 (N_11754,N_6419,N_7582);
and U11755 (N_11755,N_8314,N_5138);
nor U11756 (N_11756,N_8542,N_8719);
nand U11757 (N_11757,N_7985,N_5572);
and U11758 (N_11758,N_7742,N_8006);
or U11759 (N_11759,N_8251,N_9154);
nor U11760 (N_11760,N_6707,N_9178);
and U11761 (N_11761,N_5947,N_5932);
nor U11762 (N_11762,N_6740,N_6661);
nor U11763 (N_11763,N_7415,N_7615);
and U11764 (N_11764,N_9636,N_8591);
nor U11765 (N_11765,N_9287,N_7978);
and U11766 (N_11766,N_7572,N_9927);
nand U11767 (N_11767,N_6560,N_7697);
and U11768 (N_11768,N_6580,N_7793);
nand U11769 (N_11769,N_7256,N_9850);
or U11770 (N_11770,N_8464,N_9565);
nand U11771 (N_11771,N_5332,N_5815);
xnor U11772 (N_11772,N_9152,N_7481);
nor U11773 (N_11773,N_9391,N_5023);
nand U11774 (N_11774,N_9776,N_6315);
xnor U11775 (N_11775,N_6122,N_6206);
and U11776 (N_11776,N_7808,N_5720);
nor U11777 (N_11777,N_7387,N_8451);
nor U11778 (N_11778,N_8947,N_5024);
and U11779 (N_11779,N_8616,N_6579);
xor U11780 (N_11780,N_7144,N_8772);
or U11781 (N_11781,N_9624,N_8598);
nor U11782 (N_11782,N_6070,N_6169);
and U11783 (N_11783,N_9745,N_6692);
or U11784 (N_11784,N_7753,N_6079);
or U11785 (N_11785,N_7084,N_8624);
xnor U11786 (N_11786,N_8868,N_7266);
nor U11787 (N_11787,N_5986,N_5242);
xor U11788 (N_11788,N_7564,N_5942);
nor U11789 (N_11789,N_8075,N_7724);
nor U11790 (N_11790,N_6670,N_5782);
xor U11791 (N_11791,N_9299,N_7536);
and U11792 (N_11792,N_7288,N_7542);
xnor U11793 (N_11793,N_5033,N_5744);
and U11794 (N_11794,N_7700,N_9535);
xnor U11795 (N_11795,N_6141,N_6905);
and U11796 (N_11796,N_7537,N_5847);
nand U11797 (N_11797,N_9078,N_5481);
xnor U11798 (N_11798,N_6137,N_9243);
nand U11799 (N_11799,N_8122,N_5372);
or U11800 (N_11800,N_9242,N_7194);
xnor U11801 (N_11801,N_9108,N_8388);
xor U11802 (N_11802,N_5680,N_6023);
xnor U11803 (N_11803,N_6920,N_9939);
nor U11804 (N_11804,N_6100,N_7036);
and U11805 (N_11805,N_7281,N_5787);
or U11806 (N_11806,N_5107,N_9398);
xor U11807 (N_11807,N_6350,N_5855);
or U11808 (N_11808,N_5065,N_9010);
nor U11809 (N_11809,N_6155,N_8129);
xnor U11810 (N_11810,N_5541,N_8957);
nor U11811 (N_11811,N_7701,N_8267);
xnor U11812 (N_11812,N_8383,N_8672);
nand U11813 (N_11813,N_8324,N_7598);
or U11814 (N_11814,N_7565,N_7371);
nand U11815 (N_11815,N_7680,N_7815);
and U11816 (N_11816,N_9037,N_7331);
nand U11817 (N_11817,N_5915,N_5850);
or U11818 (N_11818,N_8851,N_7714);
and U11819 (N_11819,N_8988,N_8436);
xnor U11820 (N_11820,N_5304,N_6925);
nor U11821 (N_11821,N_7082,N_7413);
or U11822 (N_11822,N_6452,N_9968);
nand U11823 (N_11823,N_6693,N_8651);
nor U11824 (N_11824,N_7711,N_7478);
nand U11825 (N_11825,N_7709,N_9182);
or U11826 (N_11826,N_6608,N_6423);
xor U11827 (N_11827,N_6728,N_6721);
or U11828 (N_11828,N_9484,N_9981);
and U11829 (N_11829,N_8058,N_8773);
nand U11830 (N_11830,N_8040,N_7749);
nand U11831 (N_11831,N_7605,N_8036);
or U11832 (N_11832,N_9053,N_6790);
or U11833 (N_11833,N_5259,N_9809);
xor U11834 (N_11834,N_8999,N_7626);
nand U11835 (N_11835,N_9109,N_9860);
nor U11836 (N_11836,N_9910,N_6094);
and U11837 (N_11837,N_6489,N_6018);
xor U11838 (N_11838,N_6784,N_9944);
xnor U11839 (N_11839,N_8296,N_5830);
and U11840 (N_11840,N_5227,N_6607);
xnor U11841 (N_11841,N_8476,N_7675);
or U11842 (N_11842,N_7438,N_8554);
xor U11843 (N_11843,N_6990,N_8763);
or U11844 (N_11844,N_5597,N_6567);
and U11845 (N_11845,N_9086,N_5582);
or U11846 (N_11846,N_9176,N_9946);
xnor U11847 (N_11847,N_8246,N_5097);
or U11848 (N_11848,N_5936,N_6888);
nand U11849 (N_11849,N_7206,N_5505);
or U11850 (N_11850,N_9520,N_9283);
nand U11851 (N_11851,N_6166,N_6165);
nor U11852 (N_11852,N_7960,N_9188);
nand U11853 (N_11853,N_5041,N_5869);
xor U11854 (N_11854,N_6994,N_6736);
or U11855 (N_11855,N_7119,N_7233);
nand U11856 (N_11856,N_8069,N_7069);
xnor U11857 (N_11857,N_5060,N_8106);
nor U11858 (N_11858,N_9767,N_9990);
or U11859 (N_11859,N_7583,N_7876);
and U11860 (N_11860,N_5983,N_6418);
or U11861 (N_11861,N_9930,N_6384);
nand U11862 (N_11862,N_8237,N_9851);
xnor U11863 (N_11863,N_7224,N_8089);
xnor U11864 (N_11864,N_9622,N_9466);
and U11865 (N_11865,N_9122,N_9148);
or U11866 (N_11866,N_9846,N_5189);
nand U11867 (N_11867,N_5202,N_6593);
xnor U11868 (N_11868,N_7283,N_7998);
xnor U11869 (N_11869,N_9550,N_7823);
xor U11870 (N_11870,N_5311,N_8653);
and U11871 (N_11871,N_8190,N_8724);
nor U11872 (N_11872,N_6678,N_7293);
xnor U11873 (N_11873,N_9130,N_7400);
nor U11874 (N_11874,N_5265,N_7442);
nor U11875 (N_11875,N_7664,N_7822);
or U11876 (N_11876,N_7489,N_6360);
or U11877 (N_11877,N_6863,N_8878);
and U11878 (N_11878,N_9081,N_8532);
nor U11879 (N_11879,N_8896,N_5031);
xnor U11880 (N_11880,N_6487,N_6131);
nor U11881 (N_11881,N_9693,N_6392);
or U11882 (N_11882,N_7575,N_8351);
nor U11883 (N_11883,N_8902,N_9489);
nand U11884 (N_11884,N_5436,N_9832);
or U11885 (N_11885,N_8660,N_8087);
nor U11886 (N_11886,N_9906,N_6033);
xnor U11887 (N_11887,N_6931,N_7310);
nand U11888 (N_11888,N_7042,N_8452);
xnor U11889 (N_11889,N_7873,N_9543);
and U11890 (N_11890,N_8131,N_6416);
nor U11891 (N_11891,N_6969,N_7947);
nor U11892 (N_11892,N_9651,N_5881);
xnor U11893 (N_11893,N_5709,N_7553);
or U11894 (N_11894,N_8579,N_9567);
nor U11895 (N_11895,N_8525,N_8729);
and U11896 (N_11896,N_5748,N_7155);
nor U11897 (N_11897,N_6486,N_7164);
or U11898 (N_11898,N_5233,N_9428);
or U11899 (N_11899,N_7016,N_6031);
nor U11900 (N_11900,N_7462,N_6263);
and U11901 (N_11901,N_9823,N_6530);
or U11902 (N_11902,N_9051,N_8735);
nor U11903 (N_11903,N_7561,N_9085);
xnor U11904 (N_11904,N_7114,N_7394);
nand U11905 (N_11905,N_5835,N_5827);
nor U11906 (N_11906,N_5078,N_5345);
nor U11907 (N_11907,N_6118,N_7402);
nor U11908 (N_11908,N_5885,N_5636);
xnor U11909 (N_11909,N_7613,N_7096);
or U11910 (N_11910,N_5499,N_8705);
nor U11911 (N_11911,N_5009,N_9794);
nand U11912 (N_11912,N_8239,N_8358);
nand U11913 (N_11913,N_5400,N_6371);
xor U11914 (N_11914,N_8786,N_7770);
nand U11915 (N_11915,N_7779,N_7172);
nand U11916 (N_11916,N_8306,N_6658);
xnor U11917 (N_11917,N_9602,N_6817);
or U11918 (N_11918,N_6626,N_8310);
nand U11919 (N_11919,N_5493,N_8292);
or U11920 (N_11920,N_9593,N_6082);
xnor U11921 (N_11921,N_9465,N_6028);
or U11922 (N_11922,N_6457,N_9488);
nand U11923 (N_11923,N_6455,N_9066);
nand U11924 (N_11924,N_9438,N_8670);
or U11925 (N_11925,N_6550,N_8948);
xor U11926 (N_11926,N_8978,N_5836);
nand U11927 (N_11927,N_7364,N_5353);
nor U11928 (N_11928,N_8721,N_8557);
xnor U11929 (N_11929,N_9375,N_5375);
nor U11930 (N_11930,N_9665,N_9194);
nand U11931 (N_11931,N_8465,N_5993);
nor U11932 (N_11932,N_7322,N_5134);
nand U11933 (N_11933,N_8808,N_5981);
nor U11934 (N_11934,N_6928,N_7787);
xnor U11935 (N_11935,N_9742,N_5167);
xnor U11936 (N_11936,N_6201,N_9575);
nor U11937 (N_11937,N_6975,N_5610);
xor U11938 (N_11938,N_9507,N_7308);
xnor U11939 (N_11939,N_9160,N_7551);
nor U11940 (N_11940,N_8641,N_9083);
nand U11941 (N_11941,N_6192,N_9436);
nor U11942 (N_11942,N_5492,N_8016);
nor U11943 (N_11943,N_7895,N_5219);
nor U11944 (N_11944,N_5996,N_5209);
or U11945 (N_11945,N_9187,N_8944);
nor U11946 (N_11946,N_6629,N_8631);
xnor U11947 (N_11947,N_5405,N_6694);
xnor U11948 (N_11948,N_9889,N_7014);
nand U11949 (N_11949,N_7043,N_7301);
and U11950 (N_11950,N_9327,N_7725);
or U11951 (N_11951,N_8162,N_8749);
xnor U11952 (N_11952,N_9429,N_9277);
and U11953 (N_11953,N_7176,N_5601);
nand U11954 (N_11954,N_9828,N_7223);
nor U11955 (N_11955,N_5801,N_8933);
or U11956 (N_11956,N_5478,N_7000);
or U11957 (N_11957,N_6880,N_5974);
nor U11958 (N_11958,N_7355,N_7169);
or U11959 (N_11959,N_9613,N_8811);
nor U11960 (N_11960,N_7383,N_9491);
nand U11961 (N_11961,N_7430,N_9713);
or U11962 (N_11962,N_7239,N_5530);
xnor U11963 (N_11963,N_8135,N_8188);
nor U11964 (N_11964,N_9815,N_7048);
and U11965 (N_11965,N_9309,N_5277);
or U11966 (N_11966,N_5250,N_8035);
or U11967 (N_11967,N_9513,N_6318);
or U11968 (N_11968,N_6046,N_6364);
nand U11969 (N_11969,N_9784,N_5960);
xor U11970 (N_11970,N_8080,N_6602);
nand U11971 (N_11971,N_6252,N_9349);
and U11972 (N_11972,N_9067,N_9995);
and U11973 (N_11973,N_9678,N_5428);
or U11974 (N_11974,N_5962,N_6273);
nand U11975 (N_11975,N_6484,N_8311);
nand U11976 (N_11976,N_9209,N_7123);
or U11977 (N_11977,N_5524,N_9033);
xnor U11978 (N_11978,N_7556,N_8585);
or U11979 (N_11979,N_8794,N_5068);
xor U11980 (N_11980,N_9082,N_6851);
xnor U11981 (N_11981,N_9093,N_8364);
or U11982 (N_11982,N_9835,N_5978);
nand U11983 (N_11983,N_6176,N_9914);
nor U11984 (N_11984,N_5508,N_9079);
nor U11985 (N_11985,N_6065,N_9110);
nor U11986 (N_11986,N_7578,N_8969);
or U11987 (N_11987,N_8205,N_5564);
nor U11988 (N_11988,N_9714,N_7399);
nor U11989 (N_11989,N_6577,N_6587);
nand U11990 (N_11990,N_9105,N_5521);
nor U11991 (N_11991,N_9587,N_8280);
xor U11992 (N_11992,N_5342,N_8891);
and U11993 (N_11993,N_6554,N_9135);
nand U11994 (N_11994,N_9417,N_9494);
nand U11995 (N_11995,N_8807,N_9214);
nor U11996 (N_11996,N_7162,N_8341);
nand U11997 (N_11997,N_7472,N_7684);
nand U11998 (N_11998,N_6507,N_6627);
nand U11999 (N_11999,N_9951,N_7870);
xor U12000 (N_12000,N_6135,N_9294);
nor U12001 (N_12001,N_8956,N_5613);
nand U12002 (N_12002,N_5895,N_6114);
nor U12003 (N_12003,N_9885,N_7088);
nor U12004 (N_12004,N_9036,N_9988);
nand U12005 (N_12005,N_9508,N_8734);
nor U12006 (N_12006,N_7299,N_8782);
and U12007 (N_12007,N_6233,N_9580);
nor U12008 (N_12008,N_5965,N_9735);
nand U12009 (N_12009,N_5049,N_6968);
or U12010 (N_12010,N_5727,N_8327);
or U12011 (N_12011,N_7758,N_6152);
nand U12012 (N_12012,N_7627,N_8821);
nand U12013 (N_12013,N_8243,N_7547);
and U12014 (N_12014,N_7806,N_7603);
nand U12015 (N_12015,N_6892,N_9426);
or U12016 (N_12016,N_7080,N_9262);
nand U12017 (N_12017,N_8213,N_8417);
xnor U12018 (N_12018,N_6809,N_6347);
or U12019 (N_12019,N_5287,N_9958);
nor U12020 (N_12020,N_9475,N_9446);
nand U12021 (N_12021,N_8215,N_9826);
and U12022 (N_12022,N_6536,N_5756);
nand U12023 (N_12023,N_6205,N_9400);
nor U12024 (N_12024,N_9310,N_7759);
xnor U12025 (N_12025,N_6077,N_6264);
nor U12026 (N_12026,N_7943,N_9189);
and U12027 (N_12027,N_7236,N_8908);
and U12028 (N_12028,N_7566,N_6369);
nand U12029 (N_12029,N_8743,N_8791);
or U12030 (N_12030,N_6261,N_5273);
nor U12031 (N_12031,N_5245,N_9348);
or U12032 (N_12032,N_7063,N_9248);
and U12033 (N_12033,N_6901,N_6459);
nor U12034 (N_12034,N_8673,N_5929);
nor U12035 (N_12035,N_9752,N_8927);
xor U12036 (N_12036,N_9303,N_5477);
and U12037 (N_12037,N_6611,N_8875);
or U12038 (N_12038,N_6494,N_6979);
nand U12039 (N_12039,N_5364,N_9949);
nor U12040 (N_12040,N_7456,N_9937);
nor U12041 (N_12041,N_9876,N_5014);
nor U12042 (N_12042,N_6614,N_6834);
nor U12043 (N_12043,N_5319,N_9777);
nor U12044 (N_12044,N_6323,N_8027);
xnor U12045 (N_12045,N_5165,N_5488);
and U12046 (N_12046,N_7375,N_6632);
nand U12047 (N_12047,N_7262,N_8233);
and U12048 (N_12048,N_6574,N_5945);
and U12049 (N_12049,N_5415,N_6430);
nor U12050 (N_12050,N_9304,N_7648);
nor U12051 (N_12051,N_6239,N_6988);
nor U12052 (N_12052,N_5178,N_6619);
xnor U12053 (N_12053,N_9663,N_6045);
or U12054 (N_12054,N_5149,N_9457);
and U12055 (N_12055,N_8074,N_7451);
xor U12056 (N_12056,N_8874,N_6257);
nand U12057 (N_12057,N_6121,N_6129);
nor U12058 (N_12058,N_6190,N_5184);
nor U12059 (N_12059,N_9532,N_7142);
nor U12060 (N_12060,N_7548,N_6797);
xor U12061 (N_12061,N_8459,N_8962);
nand U12062 (N_12062,N_9511,N_6548);
and U12063 (N_12063,N_8640,N_6898);
nor U12064 (N_12064,N_8744,N_9959);
nor U12065 (N_12065,N_7541,N_8867);
xnor U12066 (N_12066,N_9139,N_9694);
xnor U12067 (N_12067,N_8284,N_6414);
or U12068 (N_12068,N_7193,N_6649);
nand U12069 (N_12069,N_7738,N_9601);
nand U12070 (N_12070,N_9566,N_9810);
nor U12071 (N_12071,N_6937,N_5154);
xor U12072 (N_12072,N_5482,N_5526);
xor U12073 (N_12073,N_8633,N_7339);
and U12074 (N_12074,N_9357,N_8180);
or U12075 (N_12075,N_5239,N_8921);
nand U12076 (N_12076,N_8599,N_9196);
and U12077 (N_12077,N_6368,N_9001);
nand U12078 (N_12078,N_5235,N_5174);
xor U12079 (N_12079,N_5249,N_7576);
xor U12080 (N_12080,N_5714,N_6890);
or U12081 (N_12081,N_5257,N_8064);
or U12082 (N_12082,N_9517,N_7287);
or U12083 (N_12083,N_8335,N_5114);
or U12084 (N_12084,N_9579,N_7030);
nand U12085 (N_12085,N_5285,N_6973);
or U12086 (N_12086,N_8164,N_5368);
or U12087 (N_12087,N_6226,N_5874);
and U12088 (N_12088,N_9740,N_7678);
or U12089 (N_12089,N_6373,N_5417);
nor U12090 (N_12090,N_6180,N_6891);
nor U12091 (N_12091,N_6421,N_7866);
nand U12092 (N_12092,N_7001,N_8577);
xor U12093 (N_12093,N_8576,N_5152);
nor U12094 (N_12094,N_7037,N_8003);
and U12095 (N_12095,N_6465,N_8534);
xnor U12096 (N_12096,N_6708,N_8461);
nor U12097 (N_12097,N_5282,N_5063);
or U12098 (N_12098,N_9163,N_5085);
xor U12099 (N_12099,N_8793,N_5581);
and U12100 (N_12100,N_7026,N_7962);
nor U12101 (N_12101,N_8312,N_6777);
and U12102 (N_12102,N_9395,N_9721);
xnor U12103 (N_12103,N_5308,N_6470);
or U12104 (N_12104,N_8334,N_7693);
and U12105 (N_12105,N_5798,N_8894);
or U12106 (N_12106,N_8515,N_9991);
or U12107 (N_12107,N_5664,N_9698);
nand U12108 (N_12108,N_9966,N_8478);
nand U12109 (N_12109,N_5783,N_5775);
and U12110 (N_12110,N_9431,N_6167);
and U12111 (N_12111,N_6958,N_8390);
and U12112 (N_12112,N_9205,N_9729);
or U12113 (N_12113,N_9251,N_6558);
xor U12114 (N_12114,N_5148,N_5955);
and U12115 (N_12115,N_6663,N_7835);
nor U12116 (N_12116,N_5793,N_9726);
nor U12117 (N_12117,N_9155,N_9153);
or U12118 (N_12118,N_8926,N_6057);
nor U12119 (N_12119,N_6857,N_7180);
xor U12120 (N_12120,N_7897,N_5061);
and U12121 (N_12121,N_8979,N_7683);
xor U12122 (N_12122,N_9320,N_9432);
nand U12123 (N_12123,N_6918,N_8698);
and U12124 (N_12124,N_6312,N_6677);
or U12125 (N_12125,N_5545,N_5361);
nor U12126 (N_12126,N_5142,N_9962);
nor U12127 (N_12127,N_5064,N_6300);
nor U12128 (N_12128,N_8244,N_8053);
nand U12129 (N_12129,N_8328,N_9230);
or U12130 (N_12130,N_7856,N_6778);
xor U12131 (N_12131,N_9940,N_8994);
nor U12132 (N_12132,N_8715,N_5421);
and U12133 (N_12133,N_8767,N_8654);
or U12134 (N_12134,N_6066,N_8226);
or U12135 (N_12135,N_6519,N_7213);
nor U12136 (N_12136,N_6641,N_5879);
or U12137 (N_12137,N_9275,N_7426);
xor U12138 (N_12138,N_5326,N_8584);
and U12139 (N_12139,N_6017,N_9548);
xor U12140 (N_12140,N_7642,N_5382);
xnor U12141 (N_12141,N_9288,N_6907);
or U12142 (N_12142,N_7106,N_8619);
nor U12143 (N_12143,N_8401,N_6276);
and U12144 (N_12144,N_7356,N_9892);
or U12145 (N_12145,N_9062,N_8593);
nand U12146 (N_12146,N_8219,N_7571);
or U12147 (N_12147,N_7637,N_9957);
and U12148 (N_12148,N_7015,N_9597);
and U12149 (N_12149,N_8223,N_7204);
xnor U12150 (N_12150,N_6493,N_8199);
nand U12151 (N_12151,N_8752,N_8130);
nor U12152 (N_12152,N_9883,N_9352);
xor U12153 (N_12153,N_5556,N_6353);
xor U12154 (N_12154,N_6872,N_5121);
or U12155 (N_12155,N_6837,N_7051);
nand U12156 (N_12156,N_7912,N_9872);
nand U12157 (N_12157,N_5690,N_7783);
or U12158 (N_12158,N_7021,N_6676);
or U12159 (N_12159,N_5362,N_5641);
xnor U12160 (N_12160,N_7246,N_5092);
nand U12161 (N_12161,N_5525,N_8662);
and U12162 (N_12162,N_6541,N_7087);
xor U12163 (N_12163,N_6666,N_6763);
nor U12164 (N_12164,N_5034,N_7428);
and U12165 (N_12165,N_6980,N_5244);
nand U12166 (N_12166,N_6270,N_7917);
xor U12167 (N_12167,N_5623,N_7441);
xor U12168 (N_12168,N_5269,N_5501);
xor U12169 (N_12169,N_8606,N_5828);
or U12170 (N_12170,N_8923,N_8209);
and U12171 (N_12171,N_6213,N_5573);
nand U12172 (N_12172,N_8792,N_6253);
or U12173 (N_12173,N_5440,N_8408);
xnor U12174 (N_12174,N_5799,N_5706);
nor U12175 (N_12175,N_8435,N_9096);
nand U12176 (N_12176,N_9245,N_6745);
and U12177 (N_12177,N_6237,N_5969);
nor U12178 (N_12178,N_8870,N_5892);
xnor U12179 (N_12179,N_5862,N_7791);
xor U12180 (N_12180,N_7125,N_6847);
xor U12181 (N_12181,N_6751,N_8484);
or U12182 (N_12182,N_5655,N_9785);
nor U12183 (N_12183,N_8780,N_6179);
xor U12184 (N_12184,N_8540,N_9585);
and U12185 (N_12185,N_9586,N_8037);
nor U12186 (N_12186,N_7467,N_7673);
and U12187 (N_12187,N_7350,N_5717);
xnor U12188 (N_12188,N_5848,N_6224);
nor U12189 (N_12189,N_8728,N_7820);
nand U12190 (N_12190,N_8886,N_5084);
and U12191 (N_12191,N_7320,N_6267);
nand U12192 (N_12192,N_5716,N_8198);
nor U12193 (N_12193,N_8519,N_9373);
nor U12194 (N_12194,N_5252,N_7601);
nand U12195 (N_12195,N_8804,N_7586);
nor U12196 (N_12196,N_5275,N_8264);
nor U12197 (N_12197,N_8132,N_8017);
and U12198 (N_12198,N_5042,N_7569);
or U12199 (N_12199,N_5081,N_6869);
or U12200 (N_12200,N_8679,N_6241);
xor U12201 (N_12201,N_5129,N_9916);
nand U12202 (N_12202,N_7792,N_6786);
and U12203 (N_12203,N_8681,N_6022);
or U12204 (N_12204,N_5959,N_8822);
xnor U12205 (N_12205,N_7519,N_6868);
and U12206 (N_12206,N_5207,N_7699);
and U12207 (N_12207,N_9498,N_8421);
or U12208 (N_12208,N_7345,N_8139);
xnor U12209 (N_12209,N_7832,N_6431);
and U12210 (N_12210,N_8402,N_9366);
or U12211 (N_12211,N_5841,N_8996);
and U12212 (N_12212,N_5161,N_5217);
nand U12213 (N_12213,N_5896,N_8675);
nor U12214 (N_12214,N_6309,N_7671);
and U12215 (N_12215,N_5649,N_8632);
nand U12216 (N_12216,N_9664,N_7811);
and U12217 (N_12217,N_8545,N_6145);
nor U12218 (N_12218,N_6565,N_6839);
xnor U12219 (N_12219,N_8059,N_5008);
nor U12220 (N_12220,N_8847,N_6372);
and U12221 (N_12221,N_7580,N_7028);
xnor U12222 (N_12222,N_9150,N_8551);
nand U12223 (N_12223,N_7290,N_7843);
or U12224 (N_12224,N_7452,N_7354);
nor U12225 (N_12225,N_5757,N_9859);
or U12226 (N_12226,N_7640,N_9812);
or U12227 (N_12227,N_9731,N_8105);
and U12228 (N_12228,N_6383,N_7916);
or U12229 (N_12229,N_5877,N_9746);
and U12230 (N_12230,N_8210,N_8361);
nor U12231 (N_12231,N_8546,N_7674);
or U12232 (N_12232,N_5701,N_8541);
nand U12233 (N_12233,N_9709,N_9199);
nand U12234 (N_12234,N_8683,N_5498);
and U12235 (N_12235,N_7708,N_8272);
nand U12236 (N_12236,N_5502,N_6004);
or U12237 (N_12237,N_8416,N_7591);
xnor U12238 (N_12238,N_8961,N_8343);
nor U12239 (N_12239,N_7343,N_6410);
nand U12240 (N_12240,N_7145,N_6306);
and U12241 (N_12241,N_6771,N_7669);
nor U12242 (N_12242,N_5037,N_5977);
and U12243 (N_12243,N_7776,N_6388);
xor U12244 (N_12244,N_8165,N_6174);
xor U12245 (N_12245,N_8892,N_6559);
and U12246 (N_12246,N_5004,N_5426);
or U12247 (N_12247,N_8204,N_7646);
or U12248 (N_12248,N_5027,N_8931);
or U12249 (N_12249,N_7054,N_8537);
and U12250 (N_12250,N_6229,N_7259);
and U12251 (N_12251,N_8396,N_5221);
nor U12252 (N_12252,N_8060,N_9449);
and U12253 (N_12253,N_5119,N_7842);
xor U12254 (N_12254,N_5732,N_7170);
and U12255 (N_12255,N_7679,N_6330);
and U12256 (N_12256,N_6617,N_7076);
and U12257 (N_12257,N_7480,N_7111);
or U12258 (N_12258,N_7818,N_9530);
and U12259 (N_12259,N_7260,N_7066);
xor U12260 (N_12260,N_6394,N_8486);
and U12261 (N_12261,N_8120,N_9496);
and U12262 (N_12262,N_9770,N_9923);
and U12263 (N_12263,N_6922,N_6208);
nand U12264 (N_12264,N_9688,N_9682);
and U12265 (N_12265,N_9300,N_5231);
and U12266 (N_12266,N_7486,N_5926);
xnor U12267 (N_12267,N_7552,N_8256);
xnor U12268 (N_12268,N_7179,N_9002);
and U12269 (N_12269,N_7780,N_8347);
or U12270 (N_12270,N_7685,N_6381);
or U12271 (N_12271,N_6164,N_5859);
or U12272 (N_12272,N_6242,N_5922);
nor U12273 (N_12273,N_6157,N_5921);
nor U12274 (N_12274,N_8615,N_6779);
nand U12275 (N_12275,N_9020,N_7344);
nor U12276 (N_12276,N_8093,N_9789);
nand U12277 (N_12277,N_5321,N_5886);
and U12278 (N_12278,N_7763,N_5468);
nor U12279 (N_12279,N_5527,N_9890);
xor U12280 (N_12280,N_8832,N_6846);
xnor U12281 (N_12281,N_6432,N_5956);
or U12282 (N_12282,N_6525,N_7227);
nand U12283 (N_12283,N_7198,N_5094);
nand U12284 (N_12284,N_7655,N_9564);
or U12285 (N_12285,N_9022,N_9915);
and U12286 (N_12286,N_5773,N_8825);
nor U12287 (N_12287,N_9763,N_6794);
xnor U12288 (N_12288,N_8943,N_5677);
nor U12289 (N_12289,N_8970,N_5051);
nand U12290 (N_12290,N_8222,N_7794);
nand U12291 (N_12291,N_5175,N_7761);
nor U12292 (N_12292,N_8769,N_8057);
nand U12293 (N_12293,N_5692,N_5243);
or U12294 (N_12294,N_6217,N_9545);
or U12295 (N_12295,N_7879,N_8117);
xor U12296 (N_12296,N_7826,N_7698);
and U12297 (N_12297,N_7094,N_8445);
xor U12298 (N_12298,N_6703,N_7372);
nand U12299 (N_12299,N_8694,N_7147);
and U12300 (N_12300,N_7729,N_6842);
and U12301 (N_12301,N_9072,N_5327);
or U12302 (N_12302,N_8099,N_9766);
or U12303 (N_12303,N_7534,N_9853);
nand U12304 (N_12304,N_7974,N_6050);
nand U12305 (N_12305,N_9765,N_6885);
nand U12306 (N_12306,N_8801,N_6448);
nand U12307 (N_12307,N_6211,N_8830);
nor U12308 (N_12308,N_5762,N_7105);
or U12309 (N_12309,N_9500,N_7138);
or U12310 (N_12310,N_8757,N_8553);
nand U12311 (N_12311,N_6191,N_7682);
nand U12312 (N_12312,N_7493,N_7559);
and U12313 (N_12313,N_7620,N_5280);
or U12314 (N_12314,N_6810,N_9253);
xnor U12315 (N_12315,N_7177,N_6957);
nand U12316 (N_12316,N_9244,N_8025);
nor U12317 (N_12317,N_8509,N_5298);
nand U12318 (N_12318,N_9493,N_7899);
xnor U12319 (N_12319,N_7182,N_9786);
nand U12320 (N_12320,N_5197,N_9479);
and U12321 (N_12321,N_5059,N_8639);
nand U12322 (N_12322,N_5594,N_9257);
or U12323 (N_12323,N_7367,N_6760);
and U12324 (N_12324,N_9527,N_6830);
xnor U12325 (N_12325,N_7790,N_5591);
nand U12326 (N_12326,N_9166,N_7386);
nor U12327 (N_12327,N_6092,N_8301);
xor U12328 (N_12328,N_8185,N_8570);
and U12329 (N_12329,N_6924,N_5020);
nand U12330 (N_12330,N_8148,N_8762);
and U12331 (N_12331,N_6341,N_5413);
or U12332 (N_12332,N_6088,N_7614);
and U12333 (N_12333,N_9695,N_5503);
or U12334 (N_12334,N_5159,N_9634);
xnor U12335 (N_12335,N_9703,N_7809);
and U12336 (N_12336,N_8200,N_8876);
and U12337 (N_12337,N_5849,N_5214);
or U12338 (N_12338,N_8391,N_8113);
and U12339 (N_12339,N_5790,N_5120);
xor U12340 (N_12340,N_7903,N_7031);
and U12341 (N_12341,N_9759,N_8171);
xnor U12342 (N_12342,N_6479,N_8903);
nor U12343 (N_12343,N_5433,N_7728);
nor U12344 (N_12344,N_8941,N_7965);
or U12345 (N_12345,N_6386,N_9677);
nor U12346 (N_12346,N_6903,N_5587);
nor U12347 (N_12347,N_8014,N_5579);
or U12348 (N_12348,N_7975,N_9841);
xor U12349 (N_12349,N_6469,N_5271);
nand U12350 (N_12350,N_6279,N_7140);
or U12351 (N_12351,N_9231,N_5561);
and U12352 (N_12352,N_5070,N_9666);
xor U12353 (N_12353,N_7939,N_5026);
or U12354 (N_12354,N_6917,N_5606);
or U12355 (N_12355,N_5395,N_8758);
nor U12356 (N_12356,N_9306,N_6538);
xor U12357 (N_12357,N_6996,N_6246);
nand U12358 (N_12358,N_9027,N_6083);
or U12359 (N_12359,N_7337,N_6591);
nand U12360 (N_12360,N_9370,N_6075);
xnor U12361 (N_12361,N_5088,N_5011);
nor U12362 (N_12362,N_6265,N_7935);
xnor U12363 (N_12363,N_9481,N_9167);
nor U12364 (N_12364,N_7877,N_5195);
nand U12365 (N_12365,N_6874,N_5314);
nor U12366 (N_12366,N_7686,N_6472);
nor U12367 (N_12367,N_9390,N_5767);
nand U12368 (N_12368,N_5819,N_5378);
nand U12369 (N_12369,N_6569,N_8042);
nor U12370 (N_12370,N_9091,N_7584);
nor U12371 (N_12371,N_5116,N_9483);
or U12372 (N_12372,N_5681,N_5797);
xor U12373 (N_12373,N_8443,N_8618);
or U12374 (N_12374,N_5861,N_8586);
and U12375 (N_12375,N_9045,N_7469);
nand U12376 (N_12376,N_5618,N_8522);
and U12377 (N_12377,N_5278,N_8676);
xor U12378 (N_12378,N_8565,N_5076);
nand U12379 (N_12379,N_9764,N_7563);
xor U12380 (N_12380,N_5973,N_6259);
nor U12381 (N_12381,N_7010,N_7504);
or U12382 (N_12382,N_7309,N_5096);
xnor U12383 (N_12383,N_8143,N_6564);
nor U12384 (N_12384,N_7957,N_8373);
nor U12385 (N_12385,N_5484,N_5254);
and U12386 (N_12386,N_5341,N_9011);
and U12387 (N_12387,N_5098,N_6303);
or U12388 (N_12388,N_5309,N_7365);
nor U12389 (N_12389,N_8078,N_7298);
nand U12390 (N_12390,N_5543,N_5509);
or U12391 (N_12391,N_7342,N_5670);
and U12392 (N_12392,N_7532,N_9118);
nor U12393 (N_12393,N_8516,N_7768);
xor U12394 (N_12394,N_5733,N_9359);
and U12395 (N_12395,N_8919,N_7730);
or U12396 (N_12396,N_5181,N_8332);
xor U12397 (N_12397,N_8884,N_8004);
and U12398 (N_12398,N_6518,N_7092);
or U12399 (N_12399,N_8330,N_7813);
nand U12400 (N_12400,N_5442,N_5101);
xnor U12401 (N_12401,N_5394,N_6923);
xor U12402 (N_12402,N_8230,N_5455);
nand U12403 (N_12403,N_5952,N_6322);
nor U12404 (N_12404,N_9686,N_9023);
and U12405 (N_12405,N_8678,N_7211);
and U12406 (N_12406,N_8269,N_8145);
and U12407 (N_12407,N_6803,N_8471);
nor U12408 (N_12408,N_6899,N_6014);
nand U12409 (N_12409,N_9619,N_9318);
and U12410 (N_12410,N_7349,N_9635);
nor U12411 (N_12411,N_8972,N_6126);
nand U12412 (N_12412,N_8692,N_7976);
nor U12413 (N_12413,N_8331,N_9263);
nor U12414 (N_12414,N_7201,N_7392);
nor U12415 (N_12415,N_9068,N_7496);
nand U12416 (N_12416,N_5160,N_9560);
xor U12417 (N_12417,N_6207,N_8882);
and U12418 (N_12418,N_7707,N_8802);
or U12419 (N_12419,N_5638,N_9953);
xnor U12420 (N_12420,N_7625,N_5079);
and U12421 (N_12421,N_6344,N_6078);
xor U12422 (N_12422,N_7522,N_5611);
nor U12423 (N_12423,N_9762,N_5648);
and U12424 (N_12424,N_8007,N_8500);
nand U12425 (N_12425,N_6878,N_5590);
nor U12426 (N_12426,N_8768,N_9281);
or U12427 (N_12427,N_9971,N_8995);
nor U12428 (N_12428,N_5752,N_6076);
nand U12429 (N_12429,N_9140,N_5381);
nor U12430 (N_12430,N_9618,N_5832);
nand U12431 (N_12431,N_5164,N_6397);
nor U12432 (N_12432,N_6355,N_8446);
nor U12433 (N_12433,N_7945,N_9123);
and U12434 (N_12434,N_9506,N_6112);
nand U12435 (N_12435,N_7858,N_7165);
xnor U12436 (N_12436,N_9909,N_8342);
xor U12437 (N_12437,N_6424,N_5496);
or U12438 (N_12438,N_6930,N_8043);
nand U12439 (N_12439,N_7936,N_7482);
and U12440 (N_12440,N_9623,N_7528);
nand U12441 (N_12441,N_6528,N_6478);
xor U12442 (N_12442,N_9522,N_8056);
nand U12443 (N_12443,N_6919,N_5136);
and U12444 (N_12444,N_6951,N_5740);
nand U12445 (N_12445,N_9888,N_6111);
nor U12446 (N_12446,N_7710,N_6391);
and U12447 (N_12447,N_9261,N_8021);
xor U12448 (N_12448,N_7362,N_9215);
nor U12449 (N_12449,N_9708,N_6324);
or U12450 (N_12450,N_7379,N_8952);
nand U12451 (N_12451,N_7663,N_6531);
xnor U12452 (N_12452,N_5071,N_6308);
nand U12453 (N_12453,N_5987,N_5422);
and U12454 (N_12454,N_6805,N_9771);
nand U12455 (N_12455,N_6764,N_8142);
and U12456 (N_12456,N_5419,N_9684);
or U12457 (N_12457,N_8895,N_7836);
and U12458 (N_12458,N_6047,N_5875);
nand U12459 (N_12459,N_5350,N_5293);
nand U12460 (N_12460,N_7369,N_8098);
nor U12461 (N_12461,N_5266,N_7988);
and U12462 (N_12462,N_6575,N_6149);
nand U12463 (N_12463,N_8289,N_8339);
nand U12464 (N_12464,N_9361,N_8333);
xnor U12465 (N_12465,N_9518,N_7657);
nand U12466 (N_12466,N_8677,N_9836);
or U12467 (N_12467,N_7796,N_5820);
xnor U12468 (N_12468,N_8716,N_8071);
and U12469 (N_12469,N_8690,N_7987);
or U12470 (N_12470,N_9394,N_5839);
and U12471 (N_12471,N_5276,N_5028);
or U12472 (N_12472,N_8686,N_9464);
xor U12473 (N_12473,N_5087,N_7143);
nor U12474 (N_12474,N_7358,N_5807);
or U12475 (N_12475,N_6178,N_9719);
or U12476 (N_12476,N_5077,N_5186);
nor U12477 (N_12477,N_6500,N_5844);
or U12478 (N_12478,N_6713,N_6535);
or U12479 (N_12479,N_7502,N_6249);
or U12480 (N_12480,N_8746,N_9795);
and U12481 (N_12481,N_9945,N_6295);
nand U12482 (N_12482,N_7628,N_8386);
xnor U12483 (N_12483,N_9120,N_9961);
or U12484 (N_12484,N_5927,N_9716);
xnor U12485 (N_12485,N_7318,N_7649);
nand U12486 (N_12486,N_5539,N_8646);
or U12487 (N_12487,N_9562,N_7505);
or U12488 (N_12488,N_5933,N_7668);
nor U12489 (N_12489,N_7608,N_8893);
nor U12490 (N_12490,N_9399,N_7222);
nor U12491 (N_12491,N_6287,N_7347);
and U12492 (N_12492,N_8095,N_8722);
and U12493 (N_12493,N_5749,N_8774);
xor U12494 (N_12494,N_6030,N_9578);
or U12495 (N_12495,N_7886,N_8764);
nor U12496 (N_12496,N_9570,N_9573);
and U12497 (N_12497,N_6783,N_5557);
and U12498 (N_12498,N_9996,N_7687);
and U12499 (N_12499,N_7884,N_7995);
and U12500 (N_12500,N_8168,N_5196);
xor U12501 (N_12501,N_6645,N_8887);
and U12502 (N_12502,N_7709,N_5482);
xnor U12503 (N_12503,N_5391,N_9821);
or U12504 (N_12504,N_5369,N_9812);
nor U12505 (N_12505,N_5711,N_7268);
nand U12506 (N_12506,N_6350,N_7590);
and U12507 (N_12507,N_7773,N_9638);
or U12508 (N_12508,N_8513,N_5726);
and U12509 (N_12509,N_8757,N_8811);
xor U12510 (N_12510,N_7083,N_6889);
nand U12511 (N_12511,N_7380,N_6528);
nand U12512 (N_12512,N_6883,N_6793);
nand U12513 (N_12513,N_8602,N_8731);
nor U12514 (N_12514,N_6200,N_9826);
or U12515 (N_12515,N_7065,N_5094);
nor U12516 (N_12516,N_8770,N_8738);
and U12517 (N_12517,N_9070,N_7465);
nand U12518 (N_12518,N_7642,N_5583);
nor U12519 (N_12519,N_6424,N_5754);
or U12520 (N_12520,N_7977,N_8709);
and U12521 (N_12521,N_7356,N_9756);
or U12522 (N_12522,N_8285,N_5704);
xnor U12523 (N_12523,N_6843,N_6301);
xnor U12524 (N_12524,N_6749,N_9674);
nor U12525 (N_12525,N_8461,N_9490);
and U12526 (N_12526,N_8159,N_8898);
nor U12527 (N_12527,N_5215,N_6470);
and U12528 (N_12528,N_8964,N_8004);
or U12529 (N_12529,N_5611,N_5997);
nand U12530 (N_12530,N_5925,N_6065);
nor U12531 (N_12531,N_6567,N_5836);
or U12532 (N_12532,N_6274,N_7385);
and U12533 (N_12533,N_5464,N_8928);
nand U12534 (N_12534,N_6630,N_9533);
or U12535 (N_12535,N_8577,N_6582);
and U12536 (N_12536,N_5104,N_8319);
and U12537 (N_12537,N_7138,N_5085);
nand U12538 (N_12538,N_6465,N_8087);
or U12539 (N_12539,N_5535,N_7992);
nand U12540 (N_12540,N_5431,N_7128);
or U12541 (N_12541,N_6349,N_5089);
or U12542 (N_12542,N_8898,N_6635);
nand U12543 (N_12543,N_8555,N_7154);
or U12544 (N_12544,N_8087,N_8920);
nor U12545 (N_12545,N_8398,N_8234);
nand U12546 (N_12546,N_7711,N_7070);
nor U12547 (N_12547,N_6541,N_5208);
nor U12548 (N_12548,N_5205,N_8878);
nor U12549 (N_12549,N_7548,N_7661);
nand U12550 (N_12550,N_7117,N_8779);
nand U12551 (N_12551,N_5896,N_6357);
and U12552 (N_12552,N_8205,N_5278);
nor U12553 (N_12553,N_9620,N_5802);
nor U12554 (N_12554,N_7626,N_6626);
or U12555 (N_12555,N_7662,N_5465);
nor U12556 (N_12556,N_6795,N_6352);
nand U12557 (N_12557,N_5654,N_7158);
xnor U12558 (N_12558,N_5070,N_5451);
nor U12559 (N_12559,N_6366,N_6988);
nand U12560 (N_12560,N_8824,N_8205);
nand U12561 (N_12561,N_8641,N_9725);
and U12562 (N_12562,N_6446,N_6445);
and U12563 (N_12563,N_7854,N_7102);
nor U12564 (N_12564,N_8487,N_8091);
nor U12565 (N_12565,N_7241,N_7563);
and U12566 (N_12566,N_9631,N_7838);
or U12567 (N_12567,N_6893,N_6788);
and U12568 (N_12568,N_8096,N_8198);
and U12569 (N_12569,N_9756,N_6748);
or U12570 (N_12570,N_7453,N_5094);
nand U12571 (N_12571,N_7064,N_9781);
or U12572 (N_12572,N_9258,N_5543);
and U12573 (N_12573,N_5229,N_5818);
nand U12574 (N_12574,N_9249,N_7407);
xor U12575 (N_12575,N_6622,N_6536);
xor U12576 (N_12576,N_8944,N_7180);
xnor U12577 (N_12577,N_8641,N_5302);
xor U12578 (N_12578,N_5867,N_8818);
nand U12579 (N_12579,N_9219,N_6518);
xnor U12580 (N_12580,N_9242,N_8825);
nor U12581 (N_12581,N_7326,N_5433);
xor U12582 (N_12582,N_8225,N_9959);
xnor U12583 (N_12583,N_8107,N_6681);
nor U12584 (N_12584,N_7251,N_8733);
and U12585 (N_12585,N_8506,N_8925);
nand U12586 (N_12586,N_7629,N_9000);
and U12587 (N_12587,N_9191,N_8186);
nand U12588 (N_12588,N_9549,N_6402);
nand U12589 (N_12589,N_5738,N_8929);
and U12590 (N_12590,N_9886,N_5769);
nor U12591 (N_12591,N_9672,N_6525);
xor U12592 (N_12592,N_7680,N_7283);
and U12593 (N_12593,N_5856,N_8629);
and U12594 (N_12594,N_8117,N_7406);
nor U12595 (N_12595,N_6646,N_6514);
and U12596 (N_12596,N_7998,N_7742);
nor U12597 (N_12597,N_6054,N_6065);
nand U12598 (N_12598,N_7913,N_7787);
or U12599 (N_12599,N_7862,N_7266);
or U12600 (N_12600,N_7448,N_7037);
or U12601 (N_12601,N_7459,N_5679);
xor U12602 (N_12602,N_6134,N_7319);
xnor U12603 (N_12603,N_8562,N_5953);
and U12604 (N_12604,N_7330,N_8079);
or U12605 (N_12605,N_7224,N_5884);
or U12606 (N_12606,N_9977,N_9637);
nand U12607 (N_12607,N_6691,N_7197);
xor U12608 (N_12608,N_7588,N_7153);
xor U12609 (N_12609,N_9921,N_8404);
or U12610 (N_12610,N_6622,N_9766);
nor U12611 (N_12611,N_9339,N_8997);
xor U12612 (N_12612,N_5875,N_6465);
and U12613 (N_12613,N_8608,N_9365);
xnor U12614 (N_12614,N_5976,N_6451);
nand U12615 (N_12615,N_5494,N_5515);
or U12616 (N_12616,N_9753,N_9105);
and U12617 (N_12617,N_8154,N_8668);
and U12618 (N_12618,N_5419,N_8447);
nor U12619 (N_12619,N_6607,N_9422);
xnor U12620 (N_12620,N_8724,N_5652);
nand U12621 (N_12621,N_5846,N_7556);
and U12622 (N_12622,N_6731,N_7176);
or U12623 (N_12623,N_5466,N_9127);
nor U12624 (N_12624,N_9449,N_6184);
or U12625 (N_12625,N_5244,N_7788);
or U12626 (N_12626,N_5721,N_6117);
xor U12627 (N_12627,N_7267,N_5019);
nor U12628 (N_12628,N_9729,N_6995);
or U12629 (N_12629,N_8023,N_5523);
nor U12630 (N_12630,N_8412,N_8212);
nor U12631 (N_12631,N_5386,N_8589);
xnor U12632 (N_12632,N_5908,N_8956);
xor U12633 (N_12633,N_6169,N_9008);
and U12634 (N_12634,N_9728,N_7003);
nor U12635 (N_12635,N_8866,N_8513);
and U12636 (N_12636,N_7603,N_5842);
and U12637 (N_12637,N_7298,N_7292);
nor U12638 (N_12638,N_8043,N_7054);
xor U12639 (N_12639,N_7980,N_8430);
nor U12640 (N_12640,N_6230,N_5382);
nand U12641 (N_12641,N_5470,N_7108);
nor U12642 (N_12642,N_8094,N_7450);
and U12643 (N_12643,N_5001,N_9171);
or U12644 (N_12644,N_5255,N_9345);
and U12645 (N_12645,N_5777,N_7656);
and U12646 (N_12646,N_9593,N_5624);
nor U12647 (N_12647,N_5768,N_8739);
nor U12648 (N_12648,N_7857,N_9182);
nand U12649 (N_12649,N_6377,N_8488);
nor U12650 (N_12650,N_6388,N_6984);
xor U12651 (N_12651,N_5992,N_6432);
nand U12652 (N_12652,N_9166,N_8714);
nand U12653 (N_12653,N_5806,N_8758);
nor U12654 (N_12654,N_9000,N_8084);
and U12655 (N_12655,N_8412,N_5924);
nor U12656 (N_12656,N_9340,N_6305);
nand U12657 (N_12657,N_7598,N_8239);
nand U12658 (N_12658,N_7792,N_8740);
and U12659 (N_12659,N_7984,N_9572);
nor U12660 (N_12660,N_9223,N_6608);
nor U12661 (N_12661,N_8401,N_7852);
xor U12662 (N_12662,N_6642,N_5088);
nand U12663 (N_12663,N_8398,N_5112);
and U12664 (N_12664,N_8511,N_9662);
xnor U12665 (N_12665,N_5676,N_5074);
or U12666 (N_12666,N_6466,N_6724);
nor U12667 (N_12667,N_5539,N_5008);
and U12668 (N_12668,N_9940,N_6082);
xnor U12669 (N_12669,N_6227,N_9913);
xnor U12670 (N_12670,N_7321,N_7085);
and U12671 (N_12671,N_8252,N_8384);
or U12672 (N_12672,N_7709,N_9058);
nor U12673 (N_12673,N_9203,N_8029);
nand U12674 (N_12674,N_7667,N_6707);
or U12675 (N_12675,N_7630,N_9499);
nor U12676 (N_12676,N_6541,N_7790);
and U12677 (N_12677,N_9589,N_5452);
or U12678 (N_12678,N_9760,N_5710);
nor U12679 (N_12679,N_6517,N_5964);
xnor U12680 (N_12680,N_5285,N_5786);
nor U12681 (N_12681,N_8826,N_8573);
and U12682 (N_12682,N_7593,N_8413);
nor U12683 (N_12683,N_9518,N_9274);
nor U12684 (N_12684,N_9791,N_5853);
nand U12685 (N_12685,N_9350,N_8232);
nand U12686 (N_12686,N_6604,N_6791);
xor U12687 (N_12687,N_5398,N_9456);
or U12688 (N_12688,N_8543,N_9111);
xor U12689 (N_12689,N_6324,N_6267);
nor U12690 (N_12690,N_9636,N_8033);
or U12691 (N_12691,N_6411,N_9278);
and U12692 (N_12692,N_7530,N_7600);
nor U12693 (N_12693,N_9608,N_6981);
nand U12694 (N_12694,N_6524,N_6130);
nor U12695 (N_12695,N_5686,N_5941);
xor U12696 (N_12696,N_7189,N_9130);
xor U12697 (N_12697,N_6239,N_9072);
xnor U12698 (N_12698,N_6050,N_8896);
and U12699 (N_12699,N_9510,N_9849);
and U12700 (N_12700,N_5177,N_6979);
and U12701 (N_12701,N_5909,N_6766);
nor U12702 (N_12702,N_8869,N_5257);
nand U12703 (N_12703,N_9913,N_5354);
nor U12704 (N_12704,N_6577,N_9491);
nor U12705 (N_12705,N_7783,N_7727);
nor U12706 (N_12706,N_6205,N_5932);
or U12707 (N_12707,N_5458,N_8040);
xnor U12708 (N_12708,N_5162,N_6222);
xor U12709 (N_12709,N_8713,N_5360);
xnor U12710 (N_12710,N_6445,N_9702);
and U12711 (N_12711,N_8906,N_9788);
nor U12712 (N_12712,N_5236,N_6261);
and U12713 (N_12713,N_7942,N_7281);
or U12714 (N_12714,N_7358,N_8228);
and U12715 (N_12715,N_8609,N_6263);
or U12716 (N_12716,N_9496,N_6362);
nand U12717 (N_12717,N_6628,N_5505);
or U12718 (N_12718,N_9522,N_8533);
nor U12719 (N_12719,N_6970,N_9168);
xnor U12720 (N_12720,N_5463,N_7577);
xor U12721 (N_12721,N_6839,N_9110);
xor U12722 (N_12722,N_8414,N_5977);
nand U12723 (N_12723,N_6770,N_8384);
or U12724 (N_12724,N_6777,N_5657);
and U12725 (N_12725,N_6074,N_7297);
nor U12726 (N_12726,N_5621,N_8364);
and U12727 (N_12727,N_7171,N_9782);
and U12728 (N_12728,N_8529,N_6628);
and U12729 (N_12729,N_7981,N_9341);
nor U12730 (N_12730,N_6336,N_8979);
or U12731 (N_12731,N_6080,N_5805);
xnor U12732 (N_12732,N_6171,N_5214);
xnor U12733 (N_12733,N_8754,N_6982);
nand U12734 (N_12734,N_5850,N_7816);
or U12735 (N_12735,N_8933,N_9161);
and U12736 (N_12736,N_6430,N_5146);
nand U12737 (N_12737,N_7848,N_8769);
nand U12738 (N_12738,N_6227,N_5029);
nand U12739 (N_12739,N_7505,N_5031);
xnor U12740 (N_12740,N_6449,N_9655);
and U12741 (N_12741,N_9373,N_6858);
nand U12742 (N_12742,N_7694,N_8082);
nor U12743 (N_12743,N_6055,N_8215);
or U12744 (N_12744,N_7932,N_7847);
nor U12745 (N_12745,N_9167,N_5240);
nor U12746 (N_12746,N_9861,N_7774);
xor U12747 (N_12747,N_8319,N_7870);
xnor U12748 (N_12748,N_5659,N_9953);
nor U12749 (N_12749,N_7830,N_7463);
nor U12750 (N_12750,N_8908,N_5514);
xnor U12751 (N_12751,N_5771,N_9835);
and U12752 (N_12752,N_6761,N_6750);
nand U12753 (N_12753,N_8665,N_7582);
and U12754 (N_12754,N_8700,N_5383);
xnor U12755 (N_12755,N_9852,N_6057);
and U12756 (N_12756,N_6299,N_8887);
nor U12757 (N_12757,N_5253,N_7917);
or U12758 (N_12758,N_9654,N_5222);
nor U12759 (N_12759,N_5072,N_9892);
and U12760 (N_12760,N_7513,N_9438);
nand U12761 (N_12761,N_5394,N_6877);
nor U12762 (N_12762,N_8199,N_9975);
or U12763 (N_12763,N_9751,N_8634);
xor U12764 (N_12764,N_6580,N_9546);
xnor U12765 (N_12765,N_5458,N_5738);
nor U12766 (N_12766,N_8335,N_7808);
xor U12767 (N_12767,N_8431,N_9482);
xnor U12768 (N_12768,N_8261,N_7304);
and U12769 (N_12769,N_8097,N_8731);
nand U12770 (N_12770,N_9197,N_8822);
or U12771 (N_12771,N_6460,N_5329);
nor U12772 (N_12772,N_5979,N_8211);
nand U12773 (N_12773,N_6077,N_5656);
xor U12774 (N_12774,N_5766,N_9595);
or U12775 (N_12775,N_7531,N_6973);
nand U12776 (N_12776,N_6992,N_8180);
nor U12777 (N_12777,N_6283,N_8192);
nand U12778 (N_12778,N_8084,N_5138);
or U12779 (N_12779,N_5171,N_8870);
and U12780 (N_12780,N_5314,N_6417);
nor U12781 (N_12781,N_6937,N_5688);
and U12782 (N_12782,N_6623,N_9964);
and U12783 (N_12783,N_7422,N_8436);
xor U12784 (N_12784,N_6775,N_7007);
xnor U12785 (N_12785,N_7339,N_8806);
nor U12786 (N_12786,N_7425,N_8512);
or U12787 (N_12787,N_8816,N_9360);
or U12788 (N_12788,N_6626,N_6927);
nor U12789 (N_12789,N_6445,N_8149);
and U12790 (N_12790,N_8796,N_7838);
or U12791 (N_12791,N_9565,N_5416);
or U12792 (N_12792,N_5559,N_8574);
nand U12793 (N_12793,N_7021,N_7914);
and U12794 (N_12794,N_7575,N_8349);
or U12795 (N_12795,N_9630,N_8451);
nor U12796 (N_12796,N_6826,N_9424);
nor U12797 (N_12797,N_7722,N_6089);
or U12798 (N_12798,N_5132,N_6608);
nor U12799 (N_12799,N_7859,N_8154);
and U12800 (N_12800,N_8320,N_8836);
nand U12801 (N_12801,N_5253,N_6865);
nand U12802 (N_12802,N_9499,N_9161);
and U12803 (N_12803,N_5399,N_7331);
nor U12804 (N_12804,N_6401,N_6227);
xor U12805 (N_12805,N_9558,N_7432);
or U12806 (N_12806,N_7679,N_6006);
nand U12807 (N_12807,N_6172,N_6597);
and U12808 (N_12808,N_8345,N_9950);
nor U12809 (N_12809,N_6240,N_9125);
nand U12810 (N_12810,N_6005,N_6300);
and U12811 (N_12811,N_9372,N_6925);
nand U12812 (N_12812,N_5842,N_6131);
and U12813 (N_12813,N_9442,N_9848);
or U12814 (N_12814,N_6084,N_5450);
and U12815 (N_12815,N_6426,N_8872);
or U12816 (N_12816,N_6195,N_9319);
nand U12817 (N_12817,N_7500,N_6899);
or U12818 (N_12818,N_8075,N_7463);
nand U12819 (N_12819,N_9790,N_7955);
and U12820 (N_12820,N_7305,N_5440);
xor U12821 (N_12821,N_8332,N_8568);
nor U12822 (N_12822,N_8105,N_6141);
and U12823 (N_12823,N_7506,N_8270);
nor U12824 (N_12824,N_5745,N_9596);
nor U12825 (N_12825,N_5658,N_7196);
xor U12826 (N_12826,N_9551,N_9065);
and U12827 (N_12827,N_9650,N_9140);
xor U12828 (N_12828,N_6369,N_8346);
nor U12829 (N_12829,N_9355,N_9930);
or U12830 (N_12830,N_8536,N_9930);
and U12831 (N_12831,N_5631,N_6705);
or U12832 (N_12832,N_6724,N_6534);
nor U12833 (N_12833,N_8624,N_6520);
and U12834 (N_12834,N_6438,N_8218);
xor U12835 (N_12835,N_7891,N_6208);
xnor U12836 (N_12836,N_7218,N_6711);
nand U12837 (N_12837,N_7607,N_7465);
or U12838 (N_12838,N_9476,N_8496);
and U12839 (N_12839,N_9697,N_5463);
and U12840 (N_12840,N_6157,N_9993);
nand U12841 (N_12841,N_8591,N_9467);
and U12842 (N_12842,N_8742,N_5678);
nor U12843 (N_12843,N_8211,N_6006);
and U12844 (N_12844,N_7362,N_5493);
xnor U12845 (N_12845,N_8736,N_9435);
nand U12846 (N_12846,N_9505,N_6935);
nand U12847 (N_12847,N_8451,N_6845);
nor U12848 (N_12848,N_8140,N_8601);
nand U12849 (N_12849,N_9600,N_9619);
or U12850 (N_12850,N_5558,N_8509);
nand U12851 (N_12851,N_5520,N_9427);
nor U12852 (N_12852,N_8379,N_8018);
and U12853 (N_12853,N_9406,N_8912);
and U12854 (N_12854,N_6998,N_9523);
nor U12855 (N_12855,N_5200,N_9959);
xnor U12856 (N_12856,N_6049,N_7864);
or U12857 (N_12857,N_6276,N_9767);
and U12858 (N_12858,N_6437,N_8429);
or U12859 (N_12859,N_8633,N_7094);
xnor U12860 (N_12860,N_5422,N_5697);
nor U12861 (N_12861,N_7768,N_9641);
nand U12862 (N_12862,N_7851,N_9127);
nor U12863 (N_12863,N_9416,N_9750);
xor U12864 (N_12864,N_9336,N_6075);
nand U12865 (N_12865,N_9981,N_6340);
or U12866 (N_12866,N_7675,N_9762);
xor U12867 (N_12867,N_8769,N_8606);
and U12868 (N_12868,N_7919,N_5553);
nand U12869 (N_12869,N_6545,N_7539);
nor U12870 (N_12870,N_5973,N_5548);
nand U12871 (N_12871,N_8009,N_7778);
nand U12872 (N_12872,N_8084,N_6082);
or U12873 (N_12873,N_9306,N_9559);
nand U12874 (N_12874,N_6417,N_9257);
nor U12875 (N_12875,N_9384,N_6466);
xor U12876 (N_12876,N_5584,N_8751);
and U12877 (N_12877,N_9662,N_7582);
and U12878 (N_12878,N_9806,N_6066);
or U12879 (N_12879,N_6114,N_9911);
nand U12880 (N_12880,N_6120,N_5218);
nor U12881 (N_12881,N_5323,N_7091);
or U12882 (N_12882,N_8530,N_5937);
nand U12883 (N_12883,N_6717,N_8230);
and U12884 (N_12884,N_8995,N_8268);
nand U12885 (N_12885,N_5420,N_6260);
nand U12886 (N_12886,N_7529,N_9325);
or U12887 (N_12887,N_7635,N_5726);
xor U12888 (N_12888,N_6553,N_5373);
nor U12889 (N_12889,N_8737,N_8708);
and U12890 (N_12890,N_7597,N_5739);
nor U12891 (N_12891,N_7206,N_6464);
and U12892 (N_12892,N_8190,N_8412);
nor U12893 (N_12893,N_7063,N_9895);
nand U12894 (N_12894,N_9886,N_8688);
nor U12895 (N_12895,N_7929,N_7587);
xor U12896 (N_12896,N_5088,N_6315);
xor U12897 (N_12897,N_7733,N_9317);
and U12898 (N_12898,N_8005,N_5608);
xnor U12899 (N_12899,N_8833,N_7576);
and U12900 (N_12900,N_5857,N_7921);
nand U12901 (N_12901,N_6118,N_6507);
and U12902 (N_12902,N_6048,N_7810);
nand U12903 (N_12903,N_6366,N_5840);
xor U12904 (N_12904,N_6478,N_9135);
and U12905 (N_12905,N_7162,N_5673);
xnor U12906 (N_12906,N_7176,N_9139);
xor U12907 (N_12907,N_9421,N_5611);
nand U12908 (N_12908,N_7026,N_7929);
or U12909 (N_12909,N_8032,N_8832);
nor U12910 (N_12910,N_5749,N_6875);
nor U12911 (N_12911,N_5839,N_9435);
and U12912 (N_12912,N_8010,N_6268);
xnor U12913 (N_12913,N_5396,N_8068);
and U12914 (N_12914,N_9449,N_5970);
or U12915 (N_12915,N_5738,N_9407);
xnor U12916 (N_12916,N_9488,N_5120);
xnor U12917 (N_12917,N_9710,N_6282);
and U12918 (N_12918,N_5067,N_5140);
nor U12919 (N_12919,N_9460,N_6132);
xnor U12920 (N_12920,N_9808,N_9601);
or U12921 (N_12921,N_5781,N_6899);
xor U12922 (N_12922,N_6546,N_8140);
or U12923 (N_12923,N_7143,N_7132);
or U12924 (N_12924,N_9006,N_5895);
or U12925 (N_12925,N_6900,N_5327);
xnor U12926 (N_12926,N_6295,N_9038);
and U12927 (N_12927,N_7411,N_6247);
xnor U12928 (N_12928,N_5811,N_6173);
xnor U12929 (N_12929,N_7482,N_8560);
xor U12930 (N_12930,N_5250,N_8388);
nand U12931 (N_12931,N_7626,N_7439);
xor U12932 (N_12932,N_9044,N_8463);
nor U12933 (N_12933,N_7787,N_7010);
and U12934 (N_12934,N_7808,N_6648);
and U12935 (N_12935,N_9975,N_7514);
and U12936 (N_12936,N_9722,N_5043);
and U12937 (N_12937,N_6261,N_7829);
nor U12938 (N_12938,N_6184,N_8602);
or U12939 (N_12939,N_8433,N_8742);
and U12940 (N_12940,N_6455,N_6203);
nor U12941 (N_12941,N_7145,N_7765);
xnor U12942 (N_12942,N_8054,N_8824);
xor U12943 (N_12943,N_9936,N_9970);
and U12944 (N_12944,N_5303,N_6562);
nand U12945 (N_12945,N_8817,N_6646);
or U12946 (N_12946,N_9968,N_7404);
nand U12947 (N_12947,N_5126,N_5887);
xnor U12948 (N_12948,N_7471,N_5283);
and U12949 (N_12949,N_9392,N_6216);
or U12950 (N_12950,N_5899,N_9478);
or U12951 (N_12951,N_5926,N_6065);
or U12952 (N_12952,N_7839,N_6013);
nand U12953 (N_12953,N_9734,N_7364);
or U12954 (N_12954,N_6624,N_8944);
nor U12955 (N_12955,N_9005,N_6806);
and U12956 (N_12956,N_8221,N_7243);
xor U12957 (N_12957,N_9726,N_9169);
or U12958 (N_12958,N_7776,N_9654);
and U12959 (N_12959,N_8944,N_9397);
nand U12960 (N_12960,N_6524,N_9764);
xor U12961 (N_12961,N_5092,N_9357);
and U12962 (N_12962,N_9434,N_5490);
nor U12963 (N_12963,N_7662,N_8797);
xnor U12964 (N_12964,N_6754,N_8449);
nor U12965 (N_12965,N_5214,N_8131);
nand U12966 (N_12966,N_8860,N_7886);
nand U12967 (N_12967,N_8559,N_9976);
nor U12968 (N_12968,N_6096,N_9319);
nor U12969 (N_12969,N_5733,N_9725);
and U12970 (N_12970,N_9275,N_8758);
or U12971 (N_12971,N_5926,N_6255);
and U12972 (N_12972,N_5519,N_9648);
and U12973 (N_12973,N_6843,N_5527);
or U12974 (N_12974,N_6978,N_8752);
nor U12975 (N_12975,N_6378,N_7718);
xor U12976 (N_12976,N_9976,N_8726);
xor U12977 (N_12977,N_7737,N_8486);
xnor U12978 (N_12978,N_8746,N_8735);
or U12979 (N_12979,N_5733,N_9634);
or U12980 (N_12980,N_7359,N_8179);
or U12981 (N_12981,N_9921,N_7813);
and U12982 (N_12982,N_5458,N_6286);
nand U12983 (N_12983,N_8308,N_8812);
nor U12984 (N_12984,N_6839,N_8897);
and U12985 (N_12985,N_8829,N_6380);
and U12986 (N_12986,N_5784,N_8172);
xor U12987 (N_12987,N_9521,N_5781);
xor U12988 (N_12988,N_8717,N_8445);
xor U12989 (N_12989,N_6444,N_9463);
xnor U12990 (N_12990,N_7906,N_8065);
nand U12991 (N_12991,N_6279,N_9381);
or U12992 (N_12992,N_9512,N_7171);
nand U12993 (N_12993,N_8050,N_7378);
nor U12994 (N_12994,N_5853,N_8954);
and U12995 (N_12995,N_8438,N_7404);
or U12996 (N_12996,N_5576,N_9058);
or U12997 (N_12997,N_6303,N_5186);
xor U12998 (N_12998,N_5488,N_7547);
nor U12999 (N_12999,N_5070,N_5850);
or U13000 (N_13000,N_5214,N_5217);
or U13001 (N_13001,N_9386,N_9271);
xnor U13002 (N_13002,N_8903,N_7152);
nand U13003 (N_13003,N_9062,N_6615);
and U13004 (N_13004,N_7078,N_7256);
nand U13005 (N_13005,N_8111,N_9307);
or U13006 (N_13006,N_6369,N_5769);
xnor U13007 (N_13007,N_7510,N_5171);
and U13008 (N_13008,N_9659,N_6356);
nand U13009 (N_13009,N_9667,N_6131);
nand U13010 (N_13010,N_5161,N_9740);
and U13011 (N_13011,N_8072,N_5834);
xor U13012 (N_13012,N_8484,N_7606);
or U13013 (N_13013,N_5340,N_6075);
and U13014 (N_13014,N_5072,N_5701);
xor U13015 (N_13015,N_5667,N_7911);
nand U13016 (N_13016,N_9080,N_9312);
nand U13017 (N_13017,N_5973,N_9427);
nor U13018 (N_13018,N_8683,N_5289);
xnor U13019 (N_13019,N_7497,N_7120);
xor U13020 (N_13020,N_9728,N_6880);
nor U13021 (N_13021,N_9894,N_7437);
xor U13022 (N_13022,N_8743,N_7464);
nand U13023 (N_13023,N_7421,N_8045);
or U13024 (N_13024,N_6005,N_6943);
and U13025 (N_13025,N_9654,N_5203);
nor U13026 (N_13026,N_5934,N_6254);
and U13027 (N_13027,N_6770,N_6417);
and U13028 (N_13028,N_6440,N_5542);
and U13029 (N_13029,N_5149,N_6630);
nor U13030 (N_13030,N_6138,N_7683);
xor U13031 (N_13031,N_8774,N_9521);
nor U13032 (N_13032,N_5503,N_5824);
nor U13033 (N_13033,N_6620,N_7701);
or U13034 (N_13034,N_8800,N_7053);
nand U13035 (N_13035,N_6936,N_6893);
nand U13036 (N_13036,N_5675,N_6860);
or U13037 (N_13037,N_8742,N_6116);
and U13038 (N_13038,N_5406,N_6878);
nand U13039 (N_13039,N_6719,N_6568);
or U13040 (N_13040,N_7983,N_7773);
nor U13041 (N_13041,N_9312,N_6172);
and U13042 (N_13042,N_7040,N_9435);
nor U13043 (N_13043,N_6727,N_9611);
xnor U13044 (N_13044,N_5807,N_7767);
or U13045 (N_13045,N_5783,N_6328);
xor U13046 (N_13046,N_6022,N_7726);
nand U13047 (N_13047,N_7657,N_9513);
nand U13048 (N_13048,N_7184,N_8585);
nor U13049 (N_13049,N_8084,N_8938);
or U13050 (N_13050,N_8101,N_6908);
nor U13051 (N_13051,N_9591,N_7818);
or U13052 (N_13052,N_9988,N_7601);
or U13053 (N_13053,N_8644,N_5215);
nor U13054 (N_13054,N_9010,N_6041);
nor U13055 (N_13055,N_7361,N_8839);
or U13056 (N_13056,N_5092,N_7150);
xnor U13057 (N_13057,N_5983,N_5971);
or U13058 (N_13058,N_6788,N_5944);
nor U13059 (N_13059,N_9535,N_8976);
and U13060 (N_13060,N_7742,N_8153);
or U13061 (N_13061,N_6129,N_7351);
nor U13062 (N_13062,N_8533,N_9747);
xnor U13063 (N_13063,N_5165,N_8374);
nand U13064 (N_13064,N_5513,N_8075);
nor U13065 (N_13065,N_6881,N_5584);
nor U13066 (N_13066,N_7902,N_7669);
xnor U13067 (N_13067,N_5775,N_7350);
nor U13068 (N_13068,N_6875,N_8780);
nand U13069 (N_13069,N_6188,N_8937);
or U13070 (N_13070,N_5232,N_6197);
nand U13071 (N_13071,N_6966,N_8123);
nor U13072 (N_13072,N_5434,N_6154);
nor U13073 (N_13073,N_6865,N_9057);
or U13074 (N_13074,N_6794,N_6144);
and U13075 (N_13075,N_8674,N_5849);
xnor U13076 (N_13076,N_7857,N_9401);
and U13077 (N_13077,N_8790,N_6758);
and U13078 (N_13078,N_9943,N_8871);
nand U13079 (N_13079,N_6373,N_9052);
nand U13080 (N_13080,N_7791,N_8828);
or U13081 (N_13081,N_7037,N_9602);
nand U13082 (N_13082,N_8401,N_9432);
nor U13083 (N_13083,N_9205,N_5216);
nor U13084 (N_13084,N_7362,N_8468);
nor U13085 (N_13085,N_9609,N_6425);
xnor U13086 (N_13086,N_6310,N_7136);
nor U13087 (N_13087,N_8852,N_8656);
xor U13088 (N_13088,N_7272,N_9055);
nor U13089 (N_13089,N_7897,N_5198);
and U13090 (N_13090,N_5995,N_5339);
xor U13091 (N_13091,N_6630,N_9513);
nor U13092 (N_13092,N_5729,N_7160);
or U13093 (N_13093,N_5826,N_7334);
nand U13094 (N_13094,N_9052,N_5319);
nor U13095 (N_13095,N_6557,N_5147);
nand U13096 (N_13096,N_6042,N_7898);
xor U13097 (N_13097,N_8952,N_6952);
and U13098 (N_13098,N_5525,N_6506);
or U13099 (N_13099,N_6544,N_6477);
xor U13100 (N_13100,N_8858,N_7833);
or U13101 (N_13101,N_5194,N_5723);
nand U13102 (N_13102,N_7575,N_7236);
or U13103 (N_13103,N_8164,N_8117);
or U13104 (N_13104,N_8854,N_6480);
nand U13105 (N_13105,N_6049,N_8196);
nor U13106 (N_13106,N_5823,N_9174);
and U13107 (N_13107,N_6146,N_9094);
and U13108 (N_13108,N_9939,N_9940);
xor U13109 (N_13109,N_5448,N_6125);
xor U13110 (N_13110,N_5004,N_6811);
nand U13111 (N_13111,N_8821,N_8061);
nand U13112 (N_13112,N_5521,N_5539);
or U13113 (N_13113,N_8590,N_8714);
xor U13114 (N_13114,N_9957,N_8556);
nor U13115 (N_13115,N_9036,N_9491);
nand U13116 (N_13116,N_9110,N_8730);
and U13117 (N_13117,N_8988,N_6180);
nand U13118 (N_13118,N_8199,N_6158);
xor U13119 (N_13119,N_6312,N_5795);
and U13120 (N_13120,N_9393,N_7643);
xnor U13121 (N_13121,N_7826,N_9779);
or U13122 (N_13122,N_5156,N_6917);
xor U13123 (N_13123,N_6382,N_8382);
nand U13124 (N_13124,N_8447,N_8965);
nor U13125 (N_13125,N_5565,N_9643);
xnor U13126 (N_13126,N_9563,N_5308);
nor U13127 (N_13127,N_5075,N_8670);
xor U13128 (N_13128,N_6934,N_5709);
nand U13129 (N_13129,N_5614,N_6350);
xnor U13130 (N_13130,N_9001,N_9075);
nor U13131 (N_13131,N_6216,N_9386);
and U13132 (N_13132,N_6707,N_7823);
and U13133 (N_13133,N_5062,N_8822);
xor U13134 (N_13134,N_5402,N_6260);
xor U13135 (N_13135,N_6945,N_6249);
and U13136 (N_13136,N_5390,N_7466);
or U13137 (N_13137,N_5805,N_5775);
nand U13138 (N_13138,N_7082,N_6954);
nand U13139 (N_13139,N_5920,N_6141);
nand U13140 (N_13140,N_9630,N_6844);
and U13141 (N_13141,N_8167,N_9012);
nor U13142 (N_13142,N_6847,N_9108);
nor U13143 (N_13143,N_9762,N_8275);
nand U13144 (N_13144,N_8842,N_8602);
xnor U13145 (N_13145,N_8325,N_9299);
nor U13146 (N_13146,N_9669,N_7071);
nor U13147 (N_13147,N_8453,N_5624);
nor U13148 (N_13148,N_7378,N_9348);
nor U13149 (N_13149,N_9180,N_7353);
or U13150 (N_13150,N_9471,N_8233);
nor U13151 (N_13151,N_5722,N_6473);
and U13152 (N_13152,N_5147,N_5018);
or U13153 (N_13153,N_6546,N_5652);
and U13154 (N_13154,N_5067,N_7406);
nand U13155 (N_13155,N_9645,N_9900);
nor U13156 (N_13156,N_7297,N_5190);
nor U13157 (N_13157,N_9502,N_7098);
nand U13158 (N_13158,N_5112,N_8185);
nand U13159 (N_13159,N_6173,N_5922);
nor U13160 (N_13160,N_6416,N_8866);
nand U13161 (N_13161,N_9633,N_6972);
and U13162 (N_13162,N_5820,N_7154);
and U13163 (N_13163,N_9456,N_5739);
nand U13164 (N_13164,N_6610,N_8103);
and U13165 (N_13165,N_6993,N_8312);
or U13166 (N_13166,N_6246,N_6135);
and U13167 (N_13167,N_8710,N_5140);
or U13168 (N_13168,N_5269,N_5213);
xor U13169 (N_13169,N_8465,N_7424);
nor U13170 (N_13170,N_5985,N_6990);
nand U13171 (N_13171,N_5649,N_8503);
and U13172 (N_13172,N_7744,N_7780);
nand U13173 (N_13173,N_7286,N_8779);
nor U13174 (N_13174,N_9947,N_8822);
nor U13175 (N_13175,N_5709,N_8356);
nand U13176 (N_13176,N_7753,N_7388);
nor U13177 (N_13177,N_8217,N_6275);
and U13178 (N_13178,N_9098,N_9724);
xor U13179 (N_13179,N_8412,N_6479);
or U13180 (N_13180,N_6579,N_8288);
nor U13181 (N_13181,N_9184,N_8616);
nor U13182 (N_13182,N_5390,N_6212);
nand U13183 (N_13183,N_7453,N_8984);
or U13184 (N_13184,N_9094,N_9572);
and U13185 (N_13185,N_9291,N_7542);
or U13186 (N_13186,N_5531,N_5604);
nand U13187 (N_13187,N_7834,N_9925);
and U13188 (N_13188,N_5742,N_9259);
and U13189 (N_13189,N_5216,N_8629);
nor U13190 (N_13190,N_8382,N_6117);
xnor U13191 (N_13191,N_6203,N_8026);
xor U13192 (N_13192,N_7028,N_7025);
or U13193 (N_13193,N_8260,N_5740);
nor U13194 (N_13194,N_6979,N_7731);
nand U13195 (N_13195,N_5284,N_5087);
nor U13196 (N_13196,N_6693,N_7243);
or U13197 (N_13197,N_6380,N_7115);
xor U13198 (N_13198,N_6625,N_9088);
nor U13199 (N_13199,N_6779,N_7968);
xor U13200 (N_13200,N_8987,N_5051);
nand U13201 (N_13201,N_8590,N_6374);
or U13202 (N_13202,N_6107,N_6127);
and U13203 (N_13203,N_6168,N_6737);
and U13204 (N_13204,N_9889,N_9463);
nor U13205 (N_13205,N_7607,N_6776);
and U13206 (N_13206,N_9155,N_9889);
xnor U13207 (N_13207,N_5442,N_8308);
xor U13208 (N_13208,N_8836,N_7137);
nor U13209 (N_13209,N_7613,N_9002);
xnor U13210 (N_13210,N_5955,N_5498);
xor U13211 (N_13211,N_8517,N_7019);
or U13212 (N_13212,N_9863,N_8200);
xnor U13213 (N_13213,N_8596,N_9075);
or U13214 (N_13214,N_9197,N_6100);
or U13215 (N_13215,N_6999,N_9121);
and U13216 (N_13216,N_6832,N_7112);
xor U13217 (N_13217,N_5178,N_7409);
or U13218 (N_13218,N_9084,N_5671);
nand U13219 (N_13219,N_8010,N_6532);
nor U13220 (N_13220,N_9669,N_8014);
nand U13221 (N_13221,N_6950,N_7845);
nor U13222 (N_13222,N_6716,N_6203);
xor U13223 (N_13223,N_7384,N_6809);
xor U13224 (N_13224,N_5894,N_9013);
nand U13225 (N_13225,N_7832,N_7331);
nor U13226 (N_13226,N_6985,N_7024);
and U13227 (N_13227,N_9618,N_7901);
nor U13228 (N_13228,N_8674,N_5320);
and U13229 (N_13229,N_5911,N_5339);
xor U13230 (N_13230,N_6436,N_6470);
xnor U13231 (N_13231,N_5191,N_5634);
nand U13232 (N_13232,N_7916,N_9143);
and U13233 (N_13233,N_9568,N_8160);
nand U13234 (N_13234,N_6097,N_7620);
or U13235 (N_13235,N_5204,N_5855);
and U13236 (N_13236,N_6917,N_8686);
or U13237 (N_13237,N_9786,N_7394);
or U13238 (N_13238,N_9186,N_7171);
and U13239 (N_13239,N_7557,N_9119);
nand U13240 (N_13240,N_9664,N_6441);
xor U13241 (N_13241,N_9781,N_7339);
and U13242 (N_13242,N_5664,N_6449);
nor U13243 (N_13243,N_8473,N_8853);
nor U13244 (N_13244,N_9656,N_5001);
and U13245 (N_13245,N_9842,N_8533);
nor U13246 (N_13246,N_9533,N_8740);
and U13247 (N_13247,N_9079,N_6312);
nand U13248 (N_13248,N_7517,N_5477);
or U13249 (N_13249,N_8135,N_6349);
nor U13250 (N_13250,N_8458,N_8770);
nand U13251 (N_13251,N_6663,N_6697);
and U13252 (N_13252,N_5378,N_8589);
xor U13253 (N_13253,N_5226,N_9608);
nor U13254 (N_13254,N_6252,N_7895);
xnor U13255 (N_13255,N_7396,N_9187);
or U13256 (N_13256,N_5670,N_7175);
nand U13257 (N_13257,N_7731,N_5542);
and U13258 (N_13258,N_7672,N_7747);
nand U13259 (N_13259,N_9032,N_6733);
nand U13260 (N_13260,N_6353,N_9067);
or U13261 (N_13261,N_5746,N_9822);
xor U13262 (N_13262,N_8726,N_8613);
xnor U13263 (N_13263,N_7951,N_7009);
and U13264 (N_13264,N_7241,N_9894);
xnor U13265 (N_13265,N_6026,N_7884);
xor U13266 (N_13266,N_6887,N_5995);
or U13267 (N_13267,N_8316,N_8065);
nand U13268 (N_13268,N_6661,N_8660);
nand U13269 (N_13269,N_5456,N_7134);
nand U13270 (N_13270,N_5789,N_5529);
xnor U13271 (N_13271,N_7258,N_9044);
nand U13272 (N_13272,N_9810,N_8727);
nor U13273 (N_13273,N_9569,N_5063);
or U13274 (N_13274,N_5147,N_6117);
and U13275 (N_13275,N_6389,N_6813);
and U13276 (N_13276,N_5865,N_7617);
nor U13277 (N_13277,N_5722,N_7497);
xnor U13278 (N_13278,N_5786,N_9852);
and U13279 (N_13279,N_5985,N_7900);
or U13280 (N_13280,N_9383,N_8278);
nand U13281 (N_13281,N_8465,N_5033);
xnor U13282 (N_13282,N_5038,N_5593);
or U13283 (N_13283,N_5792,N_9752);
nand U13284 (N_13284,N_8718,N_7375);
nor U13285 (N_13285,N_8823,N_9547);
nor U13286 (N_13286,N_5337,N_7429);
nand U13287 (N_13287,N_8478,N_7820);
or U13288 (N_13288,N_8864,N_9082);
nand U13289 (N_13289,N_6919,N_7601);
and U13290 (N_13290,N_7503,N_6545);
nor U13291 (N_13291,N_6639,N_9485);
xor U13292 (N_13292,N_8642,N_6504);
or U13293 (N_13293,N_6062,N_9685);
or U13294 (N_13294,N_7441,N_8113);
or U13295 (N_13295,N_9558,N_6628);
or U13296 (N_13296,N_9291,N_8124);
and U13297 (N_13297,N_8955,N_6733);
nor U13298 (N_13298,N_7422,N_8414);
and U13299 (N_13299,N_7244,N_7870);
nor U13300 (N_13300,N_9173,N_8629);
or U13301 (N_13301,N_5559,N_7987);
and U13302 (N_13302,N_7224,N_7232);
xor U13303 (N_13303,N_6319,N_5113);
and U13304 (N_13304,N_7368,N_8669);
and U13305 (N_13305,N_6142,N_5805);
and U13306 (N_13306,N_5788,N_7518);
xor U13307 (N_13307,N_8583,N_9258);
xor U13308 (N_13308,N_7005,N_8293);
and U13309 (N_13309,N_7784,N_9423);
nor U13310 (N_13310,N_7434,N_9088);
nor U13311 (N_13311,N_6867,N_8905);
or U13312 (N_13312,N_9106,N_9278);
and U13313 (N_13313,N_9301,N_6891);
nand U13314 (N_13314,N_9976,N_6175);
or U13315 (N_13315,N_5742,N_9658);
or U13316 (N_13316,N_6458,N_8271);
or U13317 (N_13317,N_6311,N_8422);
and U13318 (N_13318,N_7638,N_8465);
or U13319 (N_13319,N_9399,N_9818);
nor U13320 (N_13320,N_6036,N_6763);
nor U13321 (N_13321,N_6466,N_6087);
or U13322 (N_13322,N_6294,N_6325);
or U13323 (N_13323,N_5658,N_5587);
or U13324 (N_13324,N_8834,N_6485);
and U13325 (N_13325,N_9875,N_8062);
or U13326 (N_13326,N_5383,N_5846);
xnor U13327 (N_13327,N_7858,N_8230);
and U13328 (N_13328,N_5435,N_6274);
nand U13329 (N_13329,N_7688,N_8303);
xor U13330 (N_13330,N_6216,N_5651);
nand U13331 (N_13331,N_8676,N_6690);
or U13332 (N_13332,N_9551,N_7941);
or U13333 (N_13333,N_9033,N_8885);
nand U13334 (N_13334,N_8317,N_8144);
or U13335 (N_13335,N_8622,N_7709);
or U13336 (N_13336,N_5303,N_9243);
nor U13337 (N_13337,N_7508,N_6727);
and U13338 (N_13338,N_9274,N_5854);
xnor U13339 (N_13339,N_9813,N_5258);
xnor U13340 (N_13340,N_7131,N_7809);
xnor U13341 (N_13341,N_6550,N_5526);
or U13342 (N_13342,N_5218,N_5195);
or U13343 (N_13343,N_8649,N_5791);
nor U13344 (N_13344,N_6427,N_6782);
and U13345 (N_13345,N_7426,N_9944);
xnor U13346 (N_13346,N_5057,N_6895);
nor U13347 (N_13347,N_6060,N_8016);
xor U13348 (N_13348,N_7270,N_7836);
nand U13349 (N_13349,N_7801,N_6540);
and U13350 (N_13350,N_5803,N_9697);
or U13351 (N_13351,N_9875,N_7732);
xnor U13352 (N_13352,N_9714,N_5430);
nand U13353 (N_13353,N_9531,N_9350);
or U13354 (N_13354,N_8374,N_5733);
and U13355 (N_13355,N_5389,N_9289);
and U13356 (N_13356,N_7954,N_8062);
xnor U13357 (N_13357,N_5936,N_9020);
nor U13358 (N_13358,N_6581,N_7406);
nor U13359 (N_13359,N_8888,N_7013);
or U13360 (N_13360,N_8870,N_6346);
xor U13361 (N_13361,N_7644,N_9242);
nand U13362 (N_13362,N_7048,N_7443);
or U13363 (N_13363,N_9617,N_7901);
or U13364 (N_13364,N_6131,N_6153);
or U13365 (N_13365,N_7155,N_5354);
nand U13366 (N_13366,N_8394,N_8935);
and U13367 (N_13367,N_9288,N_8846);
and U13368 (N_13368,N_7750,N_5864);
and U13369 (N_13369,N_5067,N_6998);
and U13370 (N_13370,N_7352,N_9812);
or U13371 (N_13371,N_7983,N_8667);
xor U13372 (N_13372,N_6727,N_5520);
and U13373 (N_13373,N_6838,N_7767);
and U13374 (N_13374,N_8827,N_8308);
nor U13375 (N_13375,N_5683,N_7213);
xor U13376 (N_13376,N_6690,N_9283);
nand U13377 (N_13377,N_8073,N_8287);
or U13378 (N_13378,N_7486,N_9257);
and U13379 (N_13379,N_9387,N_8997);
xnor U13380 (N_13380,N_6945,N_8410);
xnor U13381 (N_13381,N_9427,N_9052);
xnor U13382 (N_13382,N_8780,N_5347);
and U13383 (N_13383,N_6024,N_6364);
and U13384 (N_13384,N_6073,N_8838);
nand U13385 (N_13385,N_8459,N_7578);
xnor U13386 (N_13386,N_9016,N_8780);
nand U13387 (N_13387,N_8609,N_7631);
or U13388 (N_13388,N_5889,N_8843);
and U13389 (N_13389,N_7113,N_6258);
and U13390 (N_13390,N_8368,N_5589);
xor U13391 (N_13391,N_8856,N_6347);
xnor U13392 (N_13392,N_9315,N_6131);
or U13393 (N_13393,N_8334,N_5056);
xor U13394 (N_13394,N_9132,N_5144);
xor U13395 (N_13395,N_7783,N_8947);
or U13396 (N_13396,N_9332,N_5018);
xnor U13397 (N_13397,N_9482,N_6683);
xor U13398 (N_13398,N_7413,N_7174);
nor U13399 (N_13399,N_7897,N_7485);
or U13400 (N_13400,N_9050,N_8991);
nor U13401 (N_13401,N_6280,N_5325);
and U13402 (N_13402,N_5705,N_8072);
or U13403 (N_13403,N_6055,N_6490);
nor U13404 (N_13404,N_5724,N_9876);
nand U13405 (N_13405,N_5412,N_8671);
or U13406 (N_13406,N_7011,N_9743);
or U13407 (N_13407,N_6378,N_5649);
nor U13408 (N_13408,N_5808,N_6315);
and U13409 (N_13409,N_7966,N_8784);
xnor U13410 (N_13410,N_7962,N_5469);
or U13411 (N_13411,N_5989,N_9658);
or U13412 (N_13412,N_9348,N_8587);
and U13413 (N_13413,N_7997,N_9430);
and U13414 (N_13414,N_8635,N_9377);
nand U13415 (N_13415,N_8584,N_9121);
nand U13416 (N_13416,N_8420,N_5221);
nand U13417 (N_13417,N_8816,N_7857);
nor U13418 (N_13418,N_9862,N_5218);
xnor U13419 (N_13419,N_6643,N_8232);
nor U13420 (N_13420,N_6432,N_5191);
nand U13421 (N_13421,N_5996,N_9007);
xnor U13422 (N_13422,N_5922,N_7388);
and U13423 (N_13423,N_9038,N_9956);
xor U13424 (N_13424,N_9559,N_6033);
xnor U13425 (N_13425,N_8564,N_8022);
and U13426 (N_13426,N_5573,N_9088);
and U13427 (N_13427,N_7707,N_9513);
nor U13428 (N_13428,N_6176,N_7403);
nand U13429 (N_13429,N_7118,N_8424);
xnor U13430 (N_13430,N_5583,N_7377);
nand U13431 (N_13431,N_7153,N_6166);
nand U13432 (N_13432,N_6355,N_6931);
nor U13433 (N_13433,N_8630,N_8632);
nor U13434 (N_13434,N_8154,N_6330);
nor U13435 (N_13435,N_5184,N_6667);
and U13436 (N_13436,N_9831,N_8573);
and U13437 (N_13437,N_5650,N_7690);
nand U13438 (N_13438,N_6509,N_9854);
xnor U13439 (N_13439,N_7302,N_5239);
nand U13440 (N_13440,N_5215,N_8162);
and U13441 (N_13441,N_7532,N_6578);
or U13442 (N_13442,N_6368,N_5605);
nand U13443 (N_13443,N_6497,N_6836);
nor U13444 (N_13444,N_7768,N_6240);
nor U13445 (N_13445,N_7195,N_9553);
xnor U13446 (N_13446,N_6356,N_8996);
or U13447 (N_13447,N_9028,N_8366);
nor U13448 (N_13448,N_6660,N_7364);
or U13449 (N_13449,N_8188,N_8600);
and U13450 (N_13450,N_9116,N_7525);
nand U13451 (N_13451,N_7470,N_7862);
nor U13452 (N_13452,N_9225,N_7778);
xnor U13453 (N_13453,N_9409,N_5046);
nand U13454 (N_13454,N_5960,N_9360);
and U13455 (N_13455,N_9041,N_6503);
nor U13456 (N_13456,N_8670,N_7797);
nand U13457 (N_13457,N_6549,N_9941);
xnor U13458 (N_13458,N_9243,N_6484);
nand U13459 (N_13459,N_6923,N_8186);
nor U13460 (N_13460,N_6309,N_5473);
nor U13461 (N_13461,N_5934,N_8199);
or U13462 (N_13462,N_5683,N_8011);
xor U13463 (N_13463,N_8635,N_9681);
xnor U13464 (N_13464,N_8932,N_9020);
xor U13465 (N_13465,N_9252,N_6741);
and U13466 (N_13466,N_6474,N_5580);
and U13467 (N_13467,N_8430,N_7844);
or U13468 (N_13468,N_8399,N_9894);
or U13469 (N_13469,N_7547,N_5432);
xnor U13470 (N_13470,N_8071,N_5882);
and U13471 (N_13471,N_9835,N_9789);
or U13472 (N_13472,N_5536,N_5575);
xnor U13473 (N_13473,N_8978,N_5933);
and U13474 (N_13474,N_9684,N_9673);
xor U13475 (N_13475,N_9703,N_7538);
xnor U13476 (N_13476,N_5023,N_5929);
or U13477 (N_13477,N_5921,N_8945);
nand U13478 (N_13478,N_9535,N_9934);
xnor U13479 (N_13479,N_9062,N_6160);
or U13480 (N_13480,N_9167,N_7843);
and U13481 (N_13481,N_5512,N_8084);
nor U13482 (N_13482,N_6503,N_8887);
xnor U13483 (N_13483,N_7448,N_8004);
nand U13484 (N_13484,N_5250,N_6854);
and U13485 (N_13485,N_8069,N_6844);
xor U13486 (N_13486,N_9713,N_6410);
or U13487 (N_13487,N_7686,N_8916);
nand U13488 (N_13488,N_9770,N_9817);
nor U13489 (N_13489,N_6632,N_5455);
and U13490 (N_13490,N_5697,N_8317);
nor U13491 (N_13491,N_5013,N_5366);
nor U13492 (N_13492,N_9031,N_8919);
or U13493 (N_13493,N_8683,N_6883);
or U13494 (N_13494,N_9763,N_5874);
or U13495 (N_13495,N_7880,N_6537);
nand U13496 (N_13496,N_7021,N_8320);
xnor U13497 (N_13497,N_5832,N_8207);
xor U13498 (N_13498,N_8516,N_7610);
nand U13499 (N_13499,N_6046,N_8265);
or U13500 (N_13500,N_6101,N_5786);
and U13501 (N_13501,N_9739,N_5647);
nand U13502 (N_13502,N_7169,N_8955);
and U13503 (N_13503,N_6393,N_5712);
nand U13504 (N_13504,N_6324,N_7268);
nand U13505 (N_13505,N_5755,N_5589);
or U13506 (N_13506,N_9514,N_6447);
nor U13507 (N_13507,N_6177,N_6423);
nand U13508 (N_13508,N_9265,N_9595);
nor U13509 (N_13509,N_8578,N_8540);
nand U13510 (N_13510,N_8835,N_9121);
nand U13511 (N_13511,N_9439,N_8587);
xnor U13512 (N_13512,N_5093,N_8676);
and U13513 (N_13513,N_5970,N_5659);
and U13514 (N_13514,N_9940,N_7227);
xor U13515 (N_13515,N_8665,N_7038);
and U13516 (N_13516,N_6812,N_8836);
and U13517 (N_13517,N_6423,N_9947);
nand U13518 (N_13518,N_7479,N_8399);
and U13519 (N_13519,N_6093,N_6969);
nor U13520 (N_13520,N_5431,N_6676);
nand U13521 (N_13521,N_7212,N_5214);
and U13522 (N_13522,N_5850,N_6218);
xor U13523 (N_13523,N_6689,N_7696);
xor U13524 (N_13524,N_7035,N_8094);
nand U13525 (N_13525,N_9966,N_6553);
nand U13526 (N_13526,N_6681,N_5825);
or U13527 (N_13527,N_7696,N_5970);
nor U13528 (N_13528,N_8115,N_9146);
or U13529 (N_13529,N_8696,N_6440);
nor U13530 (N_13530,N_7919,N_9687);
nand U13531 (N_13531,N_7125,N_5195);
nand U13532 (N_13532,N_7729,N_8108);
xor U13533 (N_13533,N_8911,N_5241);
or U13534 (N_13534,N_8860,N_9085);
nor U13535 (N_13535,N_7108,N_9415);
nand U13536 (N_13536,N_5348,N_7688);
xor U13537 (N_13537,N_8955,N_5886);
or U13538 (N_13538,N_9241,N_6634);
and U13539 (N_13539,N_5895,N_5572);
nor U13540 (N_13540,N_7172,N_8712);
xor U13541 (N_13541,N_8461,N_7849);
xor U13542 (N_13542,N_5561,N_5027);
nor U13543 (N_13543,N_5333,N_5233);
nand U13544 (N_13544,N_7283,N_5634);
nand U13545 (N_13545,N_5523,N_7075);
nand U13546 (N_13546,N_8277,N_8750);
xor U13547 (N_13547,N_6457,N_6061);
and U13548 (N_13548,N_7793,N_9361);
xnor U13549 (N_13549,N_9825,N_9887);
xor U13550 (N_13550,N_9446,N_5191);
or U13551 (N_13551,N_7765,N_7997);
nor U13552 (N_13552,N_5632,N_8452);
nand U13553 (N_13553,N_6646,N_7222);
nand U13554 (N_13554,N_7067,N_6462);
nor U13555 (N_13555,N_8487,N_9139);
xor U13556 (N_13556,N_7409,N_9199);
nor U13557 (N_13557,N_6070,N_7102);
nand U13558 (N_13558,N_5391,N_7857);
xnor U13559 (N_13559,N_9594,N_7407);
or U13560 (N_13560,N_9579,N_9442);
nand U13561 (N_13561,N_9830,N_6862);
nor U13562 (N_13562,N_8057,N_9954);
xor U13563 (N_13563,N_6864,N_6328);
and U13564 (N_13564,N_5474,N_7745);
and U13565 (N_13565,N_6451,N_9434);
nand U13566 (N_13566,N_7269,N_9927);
and U13567 (N_13567,N_8663,N_8568);
nor U13568 (N_13568,N_9132,N_9504);
xnor U13569 (N_13569,N_8712,N_7541);
xnor U13570 (N_13570,N_6918,N_6199);
and U13571 (N_13571,N_9400,N_7513);
and U13572 (N_13572,N_5547,N_9517);
or U13573 (N_13573,N_6569,N_8469);
xnor U13574 (N_13574,N_6756,N_7874);
or U13575 (N_13575,N_9168,N_8404);
xor U13576 (N_13576,N_6052,N_7377);
or U13577 (N_13577,N_7386,N_8139);
or U13578 (N_13578,N_7241,N_7104);
and U13579 (N_13579,N_5392,N_6502);
and U13580 (N_13580,N_6162,N_5583);
nand U13581 (N_13581,N_6149,N_8579);
or U13582 (N_13582,N_8476,N_7968);
or U13583 (N_13583,N_8092,N_6643);
xor U13584 (N_13584,N_7750,N_5585);
or U13585 (N_13585,N_6858,N_8034);
and U13586 (N_13586,N_9627,N_8528);
nor U13587 (N_13587,N_7965,N_8723);
or U13588 (N_13588,N_7033,N_6911);
nand U13589 (N_13589,N_7513,N_8455);
and U13590 (N_13590,N_8981,N_9593);
nor U13591 (N_13591,N_5996,N_6679);
and U13592 (N_13592,N_6311,N_5272);
xor U13593 (N_13593,N_7745,N_7324);
xnor U13594 (N_13594,N_5196,N_5150);
nand U13595 (N_13595,N_5795,N_6039);
xor U13596 (N_13596,N_6765,N_8058);
and U13597 (N_13597,N_5223,N_9412);
xor U13598 (N_13598,N_5633,N_6289);
nor U13599 (N_13599,N_8591,N_6634);
xnor U13600 (N_13600,N_9042,N_6668);
and U13601 (N_13601,N_5220,N_7642);
and U13602 (N_13602,N_7337,N_7508);
nor U13603 (N_13603,N_6983,N_7728);
nand U13604 (N_13604,N_5830,N_6129);
xor U13605 (N_13605,N_9290,N_8266);
or U13606 (N_13606,N_9993,N_7598);
or U13607 (N_13607,N_7356,N_5572);
xnor U13608 (N_13608,N_6357,N_7387);
xor U13609 (N_13609,N_5214,N_7564);
nand U13610 (N_13610,N_5831,N_5418);
xor U13611 (N_13611,N_7228,N_8691);
xnor U13612 (N_13612,N_8448,N_7089);
xor U13613 (N_13613,N_5562,N_9013);
xor U13614 (N_13614,N_5555,N_6456);
and U13615 (N_13615,N_5437,N_6080);
and U13616 (N_13616,N_7496,N_7921);
and U13617 (N_13617,N_7522,N_8241);
and U13618 (N_13618,N_8146,N_6398);
and U13619 (N_13619,N_6930,N_9654);
or U13620 (N_13620,N_5564,N_9540);
or U13621 (N_13621,N_9675,N_8320);
nor U13622 (N_13622,N_8940,N_7100);
and U13623 (N_13623,N_6177,N_6349);
nand U13624 (N_13624,N_5910,N_8411);
nand U13625 (N_13625,N_6310,N_5152);
and U13626 (N_13626,N_5792,N_8497);
and U13627 (N_13627,N_7990,N_7344);
xnor U13628 (N_13628,N_7055,N_6851);
or U13629 (N_13629,N_8591,N_8608);
or U13630 (N_13630,N_5490,N_8883);
and U13631 (N_13631,N_9594,N_6772);
or U13632 (N_13632,N_6357,N_8766);
xor U13633 (N_13633,N_6693,N_8054);
xor U13634 (N_13634,N_6917,N_7577);
nand U13635 (N_13635,N_6348,N_9596);
nand U13636 (N_13636,N_7171,N_5272);
or U13637 (N_13637,N_9669,N_5077);
nor U13638 (N_13638,N_7060,N_8377);
or U13639 (N_13639,N_7027,N_6998);
xor U13640 (N_13640,N_5670,N_5366);
nor U13641 (N_13641,N_9203,N_6685);
nor U13642 (N_13642,N_5185,N_6217);
and U13643 (N_13643,N_8744,N_8734);
nor U13644 (N_13644,N_9603,N_9914);
nor U13645 (N_13645,N_8610,N_6609);
and U13646 (N_13646,N_7602,N_9212);
nand U13647 (N_13647,N_8314,N_8843);
nand U13648 (N_13648,N_5214,N_8444);
xnor U13649 (N_13649,N_5175,N_5353);
nor U13650 (N_13650,N_7478,N_5964);
or U13651 (N_13651,N_9066,N_5062);
or U13652 (N_13652,N_5823,N_6017);
nand U13653 (N_13653,N_8332,N_9380);
and U13654 (N_13654,N_5067,N_7742);
xor U13655 (N_13655,N_7072,N_8426);
xnor U13656 (N_13656,N_8077,N_9957);
and U13657 (N_13657,N_5116,N_5067);
or U13658 (N_13658,N_5183,N_5547);
or U13659 (N_13659,N_6614,N_6071);
and U13660 (N_13660,N_9663,N_8927);
nor U13661 (N_13661,N_6493,N_9317);
xor U13662 (N_13662,N_9735,N_6152);
nor U13663 (N_13663,N_8452,N_8682);
nand U13664 (N_13664,N_9005,N_5727);
nor U13665 (N_13665,N_7740,N_9597);
xnor U13666 (N_13666,N_8704,N_7910);
or U13667 (N_13667,N_7226,N_5356);
xnor U13668 (N_13668,N_9733,N_6994);
or U13669 (N_13669,N_8573,N_9662);
nor U13670 (N_13670,N_6469,N_7963);
nor U13671 (N_13671,N_8062,N_8847);
xor U13672 (N_13672,N_8549,N_9378);
or U13673 (N_13673,N_6373,N_6798);
and U13674 (N_13674,N_9684,N_8031);
or U13675 (N_13675,N_5807,N_7569);
or U13676 (N_13676,N_5130,N_6978);
or U13677 (N_13677,N_5913,N_6301);
nor U13678 (N_13678,N_6565,N_8211);
or U13679 (N_13679,N_7042,N_5489);
xnor U13680 (N_13680,N_9529,N_8501);
nor U13681 (N_13681,N_6023,N_5221);
or U13682 (N_13682,N_6504,N_9188);
and U13683 (N_13683,N_9794,N_8428);
or U13684 (N_13684,N_9789,N_6915);
nor U13685 (N_13685,N_6824,N_8732);
nor U13686 (N_13686,N_7796,N_5082);
and U13687 (N_13687,N_5394,N_5785);
xor U13688 (N_13688,N_5342,N_6041);
and U13689 (N_13689,N_9714,N_7056);
or U13690 (N_13690,N_6613,N_6823);
and U13691 (N_13691,N_8139,N_5728);
nand U13692 (N_13692,N_9358,N_8185);
nand U13693 (N_13693,N_6622,N_6062);
nand U13694 (N_13694,N_5384,N_8756);
or U13695 (N_13695,N_8217,N_9474);
or U13696 (N_13696,N_7389,N_8735);
xnor U13697 (N_13697,N_6340,N_8436);
nand U13698 (N_13698,N_9158,N_8668);
xnor U13699 (N_13699,N_6284,N_9512);
and U13700 (N_13700,N_8658,N_6730);
nand U13701 (N_13701,N_8240,N_6803);
nand U13702 (N_13702,N_7871,N_6499);
nor U13703 (N_13703,N_5787,N_8248);
or U13704 (N_13704,N_8916,N_6035);
nor U13705 (N_13705,N_6383,N_8352);
nand U13706 (N_13706,N_5200,N_9649);
xnor U13707 (N_13707,N_7095,N_9723);
nand U13708 (N_13708,N_6198,N_6507);
and U13709 (N_13709,N_5338,N_9573);
nand U13710 (N_13710,N_9018,N_9649);
nand U13711 (N_13711,N_5665,N_9966);
xnor U13712 (N_13712,N_8854,N_7725);
nand U13713 (N_13713,N_9040,N_8445);
xor U13714 (N_13714,N_7244,N_7028);
or U13715 (N_13715,N_5587,N_8177);
nor U13716 (N_13716,N_6342,N_7092);
and U13717 (N_13717,N_8808,N_6111);
nor U13718 (N_13718,N_6243,N_9596);
or U13719 (N_13719,N_8323,N_5699);
and U13720 (N_13720,N_7840,N_6715);
xor U13721 (N_13721,N_8694,N_8970);
or U13722 (N_13722,N_5935,N_9293);
nand U13723 (N_13723,N_5801,N_7557);
nor U13724 (N_13724,N_5956,N_7382);
nand U13725 (N_13725,N_9434,N_7863);
nand U13726 (N_13726,N_7336,N_5111);
nand U13727 (N_13727,N_8403,N_9938);
nand U13728 (N_13728,N_9126,N_8591);
nand U13729 (N_13729,N_8376,N_5272);
nand U13730 (N_13730,N_6665,N_5461);
nor U13731 (N_13731,N_8197,N_5577);
nor U13732 (N_13732,N_6986,N_8470);
nand U13733 (N_13733,N_5425,N_5682);
and U13734 (N_13734,N_9637,N_6844);
xnor U13735 (N_13735,N_6566,N_8579);
or U13736 (N_13736,N_9645,N_9543);
nor U13737 (N_13737,N_7090,N_8793);
or U13738 (N_13738,N_6286,N_6497);
xor U13739 (N_13739,N_9290,N_5105);
nand U13740 (N_13740,N_5983,N_6449);
and U13741 (N_13741,N_8019,N_6033);
and U13742 (N_13742,N_5085,N_6120);
nor U13743 (N_13743,N_9018,N_7636);
nor U13744 (N_13744,N_9450,N_7217);
nand U13745 (N_13745,N_6233,N_5624);
nor U13746 (N_13746,N_7061,N_6059);
and U13747 (N_13747,N_8271,N_8866);
or U13748 (N_13748,N_7737,N_5486);
nand U13749 (N_13749,N_6574,N_8297);
nand U13750 (N_13750,N_5275,N_6839);
or U13751 (N_13751,N_9645,N_7970);
nor U13752 (N_13752,N_7476,N_6426);
xnor U13753 (N_13753,N_6710,N_9532);
nor U13754 (N_13754,N_6050,N_7587);
xnor U13755 (N_13755,N_9539,N_5552);
or U13756 (N_13756,N_6034,N_7454);
or U13757 (N_13757,N_7441,N_9273);
or U13758 (N_13758,N_7063,N_8637);
xor U13759 (N_13759,N_7700,N_9389);
xnor U13760 (N_13760,N_5024,N_6223);
nand U13761 (N_13761,N_6577,N_7704);
nand U13762 (N_13762,N_5008,N_5325);
or U13763 (N_13763,N_9378,N_6139);
nand U13764 (N_13764,N_9342,N_9938);
nand U13765 (N_13765,N_8051,N_6718);
nand U13766 (N_13766,N_8431,N_9187);
nor U13767 (N_13767,N_8531,N_5143);
nor U13768 (N_13768,N_6747,N_9063);
xnor U13769 (N_13769,N_5659,N_6466);
or U13770 (N_13770,N_7766,N_6475);
or U13771 (N_13771,N_9495,N_7554);
xor U13772 (N_13772,N_5546,N_6926);
and U13773 (N_13773,N_5736,N_7276);
nand U13774 (N_13774,N_7373,N_5312);
and U13775 (N_13775,N_9413,N_6016);
nor U13776 (N_13776,N_5978,N_7285);
and U13777 (N_13777,N_6426,N_5375);
nor U13778 (N_13778,N_6008,N_6659);
nand U13779 (N_13779,N_6477,N_7452);
nand U13780 (N_13780,N_9054,N_6555);
nor U13781 (N_13781,N_6328,N_7298);
nor U13782 (N_13782,N_7989,N_6760);
or U13783 (N_13783,N_5974,N_5718);
nand U13784 (N_13784,N_7333,N_6971);
xor U13785 (N_13785,N_8870,N_7915);
nor U13786 (N_13786,N_5092,N_5752);
and U13787 (N_13787,N_8596,N_8200);
and U13788 (N_13788,N_7677,N_8962);
xnor U13789 (N_13789,N_7802,N_6956);
or U13790 (N_13790,N_9176,N_8938);
nand U13791 (N_13791,N_6331,N_8137);
nand U13792 (N_13792,N_9035,N_5629);
and U13793 (N_13793,N_7558,N_5467);
and U13794 (N_13794,N_9860,N_7162);
nor U13795 (N_13795,N_7987,N_6102);
and U13796 (N_13796,N_8292,N_9650);
xor U13797 (N_13797,N_8531,N_9808);
or U13798 (N_13798,N_7031,N_7350);
and U13799 (N_13799,N_6327,N_6690);
xor U13800 (N_13800,N_7629,N_9469);
and U13801 (N_13801,N_5801,N_9994);
nor U13802 (N_13802,N_7548,N_5485);
xnor U13803 (N_13803,N_5933,N_8257);
and U13804 (N_13804,N_9454,N_5183);
nand U13805 (N_13805,N_6189,N_6204);
nand U13806 (N_13806,N_9917,N_7038);
nand U13807 (N_13807,N_9947,N_6143);
nand U13808 (N_13808,N_7050,N_5716);
or U13809 (N_13809,N_9277,N_5523);
or U13810 (N_13810,N_6181,N_5473);
nand U13811 (N_13811,N_8475,N_7545);
and U13812 (N_13812,N_7201,N_9078);
and U13813 (N_13813,N_6825,N_6846);
or U13814 (N_13814,N_5746,N_7889);
and U13815 (N_13815,N_8546,N_9324);
nand U13816 (N_13816,N_6491,N_8165);
and U13817 (N_13817,N_8921,N_5296);
nand U13818 (N_13818,N_5471,N_7800);
xor U13819 (N_13819,N_7780,N_6195);
or U13820 (N_13820,N_8493,N_5418);
or U13821 (N_13821,N_8522,N_7367);
nand U13822 (N_13822,N_9472,N_9900);
nand U13823 (N_13823,N_6306,N_7576);
xor U13824 (N_13824,N_5873,N_6644);
and U13825 (N_13825,N_6038,N_5584);
xnor U13826 (N_13826,N_8310,N_6854);
xnor U13827 (N_13827,N_6146,N_9724);
or U13828 (N_13828,N_8656,N_8401);
or U13829 (N_13829,N_9205,N_7620);
or U13830 (N_13830,N_7072,N_8471);
nor U13831 (N_13831,N_7974,N_8919);
nor U13832 (N_13832,N_9608,N_8851);
and U13833 (N_13833,N_9030,N_9104);
nor U13834 (N_13834,N_5198,N_8429);
nand U13835 (N_13835,N_7712,N_6445);
nand U13836 (N_13836,N_7761,N_8928);
and U13837 (N_13837,N_9857,N_7236);
or U13838 (N_13838,N_9518,N_5764);
nor U13839 (N_13839,N_5808,N_8396);
xnor U13840 (N_13840,N_9124,N_8299);
xor U13841 (N_13841,N_7149,N_9631);
xor U13842 (N_13842,N_9331,N_8012);
nor U13843 (N_13843,N_5091,N_6062);
and U13844 (N_13844,N_8656,N_6093);
xor U13845 (N_13845,N_7088,N_6803);
or U13846 (N_13846,N_6092,N_7200);
xnor U13847 (N_13847,N_5791,N_8930);
or U13848 (N_13848,N_8391,N_7785);
nand U13849 (N_13849,N_5070,N_8421);
nor U13850 (N_13850,N_5517,N_8288);
xor U13851 (N_13851,N_7381,N_9644);
xor U13852 (N_13852,N_8890,N_9258);
or U13853 (N_13853,N_5075,N_9351);
or U13854 (N_13854,N_8414,N_9636);
xor U13855 (N_13855,N_5388,N_8167);
and U13856 (N_13856,N_9741,N_5851);
xor U13857 (N_13857,N_5881,N_9257);
xor U13858 (N_13858,N_7346,N_9058);
nand U13859 (N_13859,N_6503,N_9889);
nand U13860 (N_13860,N_9418,N_5987);
nor U13861 (N_13861,N_6494,N_6719);
and U13862 (N_13862,N_5255,N_9817);
or U13863 (N_13863,N_9144,N_6314);
xor U13864 (N_13864,N_8826,N_9093);
nand U13865 (N_13865,N_7341,N_8587);
xnor U13866 (N_13866,N_7305,N_5831);
xor U13867 (N_13867,N_7416,N_5930);
or U13868 (N_13868,N_9947,N_5698);
nand U13869 (N_13869,N_5015,N_9295);
nand U13870 (N_13870,N_9205,N_6152);
nand U13871 (N_13871,N_6050,N_6871);
or U13872 (N_13872,N_8519,N_7361);
nor U13873 (N_13873,N_7581,N_8427);
nand U13874 (N_13874,N_5223,N_7762);
or U13875 (N_13875,N_9375,N_8771);
nor U13876 (N_13876,N_6243,N_5509);
xnor U13877 (N_13877,N_7489,N_9710);
xor U13878 (N_13878,N_7269,N_6081);
nand U13879 (N_13879,N_7460,N_8481);
nand U13880 (N_13880,N_7647,N_9558);
xnor U13881 (N_13881,N_6115,N_8365);
nand U13882 (N_13882,N_9126,N_8036);
and U13883 (N_13883,N_7205,N_8879);
and U13884 (N_13884,N_8946,N_8387);
and U13885 (N_13885,N_6859,N_9727);
xor U13886 (N_13886,N_9500,N_5698);
xnor U13887 (N_13887,N_6423,N_5898);
nor U13888 (N_13888,N_9428,N_9524);
or U13889 (N_13889,N_7188,N_5980);
and U13890 (N_13890,N_6353,N_6653);
and U13891 (N_13891,N_8591,N_9356);
nor U13892 (N_13892,N_8693,N_9080);
xnor U13893 (N_13893,N_6512,N_5893);
nor U13894 (N_13894,N_9564,N_5760);
nor U13895 (N_13895,N_6471,N_8995);
or U13896 (N_13896,N_5406,N_6475);
or U13897 (N_13897,N_8359,N_5286);
or U13898 (N_13898,N_5687,N_6698);
nor U13899 (N_13899,N_5947,N_9653);
and U13900 (N_13900,N_8035,N_8027);
nand U13901 (N_13901,N_8424,N_5744);
nand U13902 (N_13902,N_9747,N_6568);
or U13903 (N_13903,N_7300,N_9585);
nand U13904 (N_13904,N_8417,N_5517);
and U13905 (N_13905,N_6016,N_8488);
or U13906 (N_13906,N_5164,N_5526);
or U13907 (N_13907,N_5222,N_9756);
xnor U13908 (N_13908,N_7664,N_6398);
or U13909 (N_13909,N_5794,N_8767);
nor U13910 (N_13910,N_7534,N_7036);
nand U13911 (N_13911,N_6359,N_9838);
xor U13912 (N_13912,N_5694,N_9963);
nand U13913 (N_13913,N_9601,N_8073);
xnor U13914 (N_13914,N_5596,N_5446);
nor U13915 (N_13915,N_6043,N_6379);
nand U13916 (N_13916,N_8650,N_5074);
xnor U13917 (N_13917,N_7211,N_6161);
nor U13918 (N_13918,N_8544,N_8142);
nand U13919 (N_13919,N_6494,N_9018);
or U13920 (N_13920,N_7732,N_9737);
and U13921 (N_13921,N_5551,N_9496);
or U13922 (N_13922,N_6445,N_6554);
or U13923 (N_13923,N_8821,N_6007);
nand U13924 (N_13924,N_6379,N_9949);
nand U13925 (N_13925,N_6174,N_6528);
and U13926 (N_13926,N_7951,N_7534);
xor U13927 (N_13927,N_6095,N_6612);
and U13928 (N_13928,N_9493,N_6002);
xor U13929 (N_13929,N_5412,N_5917);
nor U13930 (N_13930,N_7159,N_6370);
or U13931 (N_13931,N_9521,N_7268);
nand U13932 (N_13932,N_6249,N_5658);
xor U13933 (N_13933,N_8764,N_7988);
nor U13934 (N_13934,N_6740,N_5294);
xnor U13935 (N_13935,N_9065,N_8572);
nand U13936 (N_13936,N_9190,N_9230);
xnor U13937 (N_13937,N_6215,N_8876);
nor U13938 (N_13938,N_6585,N_6614);
xor U13939 (N_13939,N_6925,N_7031);
xnor U13940 (N_13940,N_6471,N_5665);
and U13941 (N_13941,N_8153,N_8520);
xor U13942 (N_13942,N_9117,N_6934);
xnor U13943 (N_13943,N_7332,N_9921);
or U13944 (N_13944,N_5879,N_5946);
xor U13945 (N_13945,N_5339,N_7013);
and U13946 (N_13946,N_6745,N_6166);
nor U13947 (N_13947,N_8401,N_9721);
nand U13948 (N_13948,N_7677,N_6040);
nand U13949 (N_13949,N_7021,N_7318);
xnor U13950 (N_13950,N_9743,N_5198);
or U13951 (N_13951,N_5618,N_7641);
nand U13952 (N_13952,N_8460,N_6487);
nor U13953 (N_13953,N_8454,N_5709);
or U13954 (N_13954,N_7405,N_6948);
nand U13955 (N_13955,N_8269,N_7391);
and U13956 (N_13956,N_6676,N_9159);
nand U13957 (N_13957,N_9746,N_7246);
nand U13958 (N_13958,N_7976,N_8560);
xor U13959 (N_13959,N_9080,N_8649);
xor U13960 (N_13960,N_9423,N_7175);
or U13961 (N_13961,N_9947,N_6163);
nor U13962 (N_13962,N_7381,N_8686);
and U13963 (N_13963,N_5736,N_7150);
and U13964 (N_13964,N_8017,N_7513);
xor U13965 (N_13965,N_7170,N_6946);
or U13966 (N_13966,N_8212,N_9078);
or U13967 (N_13967,N_9992,N_9423);
and U13968 (N_13968,N_5292,N_8789);
xor U13969 (N_13969,N_5989,N_7622);
nor U13970 (N_13970,N_6752,N_9835);
and U13971 (N_13971,N_5865,N_5090);
nand U13972 (N_13972,N_9288,N_9278);
nor U13973 (N_13973,N_8608,N_7939);
nor U13974 (N_13974,N_8759,N_9751);
xnor U13975 (N_13975,N_9310,N_6191);
and U13976 (N_13976,N_8991,N_7960);
and U13977 (N_13977,N_9435,N_6143);
or U13978 (N_13978,N_7436,N_6600);
nand U13979 (N_13979,N_9792,N_9404);
and U13980 (N_13980,N_9622,N_5357);
nor U13981 (N_13981,N_7415,N_6193);
or U13982 (N_13982,N_7754,N_5372);
nor U13983 (N_13983,N_5480,N_5231);
and U13984 (N_13984,N_9744,N_7530);
nor U13985 (N_13985,N_6296,N_9365);
or U13986 (N_13986,N_8313,N_9156);
or U13987 (N_13987,N_7671,N_7712);
and U13988 (N_13988,N_6245,N_9323);
xnor U13989 (N_13989,N_5011,N_6228);
nand U13990 (N_13990,N_7196,N_8274);
or U13991 (N_13991,N_7279,N_5575);
xor U13992 (N_13992,N_8817,N_5845);
nor U13993 (N_13993,N_5657,N_8445);
nor U13994 (N_13994,N_9427,N_8839);
nor U13995 (N_13995,N_5558,N_5085);
and U13996 (N_13996,N_9673,N_5094);
nor U13997 (N_13997,N_8294,N_7947);
and U13998 (N_13998,N_9613,N_6702);
xor U13999 (N_13999,N_8428,N_9640);
or U14000 (N_14000,N_7598,N_5078);
nand U14001 (N_14001,N_6634,N_7807);
nand U14002 (N_14002,N_6358,N_6952);
and U14003 (N_14003,N_5512,N_5601);
and U14004 (N_14004,N_5033,N_6684);
and U14005 (N_14005,N_6120,N_6064);
nand U14006 (N_14006,N_6525,N_5486);
or U14007 (N_14007,N_8249,N_9690);
and U14008 (N_14008,N_9248,N_8135);
and U14009 (N_14009,N_8818,N_5379);
nand U14010 (N_14010,N_6580,N_9975);
nor U14011 (N_14011,N_5553,N_9691);
nand U14012 (N_14012,N_5532,N_7964);
nor U14013 (N_14013,N_7759,N_5745);
xor U14014 (N_14014,N_6870,N_5685);
nor U14015 (N_14015,N_6735,N_8304);
nand U14016 (N_14016,N_7843,N_8022);
xor U14017 (N_14017,N_9114,N_9950);
or U14018 (N_14018,N_9156,N_9044);
and U14019 (N_14019,N_7610,N_8707);
and U14020 (N_14020,N_8477,N_9365);
nand U14021 (N_14021,N_8153,N_8008);
nand U14022 (N_14022,N_8395,N_9054);
nor U14023 (N_14023,N_8299,N_8770);
nand U14024 (N_14024,N_5719,N_5123);
nand U14025 (N_14025,N_5635,N_5143);
nand U14026 (N_14026,N_9959,N_9628);
and U14027 (N_14027,N_7546,N_8652);
nor U14028 (N_14028,N_6688,N_6956);
or U14029 (N_14029,N_6881,N_8487);
or U14030 (N_14030,N_8586,N_8288);
and U14031 (N_14031,N_8226,N_7250);
nand U14032 (N_14032,N_7110,N_6923);
nand U14033 (N_14033,N_5009,N_5893);
or U14034 (N_14034,N_7023,N_5507);
nor U14035 (N_14035,N_5823,N_8620);
or U14036 (N_14036,N_5264,N_8289);
and U14037 (N_14037,N_6551,N_8300);
xnor U14038 (N_14038,N_9548,N_6355);
or U14039 (N_14039,N_5306,N_7003);
xor U14040 (N_14040,N_8663,N_9509);
xor U14041 (N_14041,N_7275,N_6633);
or U14042 (N_14042,N_9536,N_5828);
and U14043 (N_14043,N_7033,N_8882);
nor U14044 (N_14044,N_9466,N_5143);
or U14045 (N_14045,N_7220,N_5732);
nand U14046 (N_14046,N_5951,N_9506);
nand U14047 (N_14047,N_5363,N_9167);
nor U14048 (N_14048,N_6989,N_9804);
nor U14049 (N_14049,N_6815,N_6285);
nor U14050 (N_14050,N_9252,N_9075);
xor U14051 (N_14051,N_5421,N_7616);
or U14052 (N_14052,N_9589,N_9575);
nand U14053 (N_14053,N_5684,N_5282);
nand U14054 (N_14054,N_8651,N_9497);
nor U14055 (N_14055,N_9923,N_7485);
or U14056 (N_14056,N_5801,N_5456);
or U14057 (N_14057,N_7101,N_6229);
or U14058 (N_14058,N_6267,N_8321);
and U14059 (N_14059,N_7063,N_9538);
or U14060 (N_14060,N_6767,N_7291);
and U14061 (N_14061,N_5023,N_8058);
and U14062 (N_14062,N_9197,N_7369);
xor U14063 (N_14063,N_9433,N_8868);
nand U14064 (N_14064,N_9159,N_8474);
nor U14065 (N_14065,N_8231,N_8973);
xor U14066 (N_14066,N_9820,N_7069);
xor U14067 (N_14067,N_7623,N_7694);
and U14068 (N_14068,N_9619,N_5859);
or U14069 (N_14069,N_8826,N_6874);
nor U14070 (N_14070,N_8911,N_6415);
and U14071 (N_14071,N_5991,N_9406);
or U14072 (N_14072,N_8961,N_8099);
nor U14073 (N_14073,N_5075,N_9048);
nand U14074 (N_14074,N_5441,N_6205);
nand U14075 (N_14075,N_6896,N_8761);
or U14076 (N_14076,N_8484,N_9516);
nand U14077 (N_14077,N_8872,N_6326);
and U14078 (N_14078,N_5694,N_6085);
and U14079 (N_14079,N_9842,N_6231);
and U14080 (N_14080,N_8808,N_6163);
nor U14081 (N_14081,N_9230,N_7261);
nand U14082 (N_14082,N_6442,N_7838);
or U14083 (N_14083,N_8336,N_5550);
and U14084 (N_14084,N_9312,N_9989);
nor U14085 (N_14085,N_8637,N_5887);
and U14086 (N_14086,N_9705,N_9541);
nor U14087 (N_14087,N_7458,N_5930);
xnor U14088 (N_14088,N_7126,N_5716);
or U14089 (N_14089,N_9381,N_6907);
or U14090 (N_14090,N_7679,N_6811);
or U14091 (N_14091,N_5119,N_7330);
xnor U14092 (N_14092,N_5271,N_7455);
xnor U14093 (N_14093,N_9685,N_7142);
or U14094 (N_14094,N_5229,N_9140);
and U14095 (N_14095,N_9477,N_8690);
or U14096 (N_14096,N_7370,N_6100);
xor U14097 (N_14097,N_7568,N_5103);
or U14098 (N_14098,N_8376,N_6378);
nand U14099 (N_14099,N_5243,N_6836);
nand U14100 (N_14100,N_7900,N_6412);
nor U14101 (N_14101,N_5815,N_6598);
or U14102 (N_14102,N_8165,N_7129);
and U14103 (N_14103,N_5317,N_5331);
or U14104 (N_14104,N_9843,N_9899);
nand U14105 (N_14105,N_7966,N_5117);
and U14106 (N_14106,N_5841,N_6788);
nand U14107 (N_14107,N_6745,N_6693);
nor U14108 (N_14108,N_9537,N_6671);
nor U14109 (N_14109,N_5032,N_7204);
nor U14110 (N_14110,N_8460,N_5391);
xnor U14111 (N_14111,N_8253,N_9290);
nand U14112 (N_14112,N_6952,N_5354);
and U14113 (N_14113,N_9716,N_7810);
nor U14114 (N_14114,N_5621,N_7606);
nand U14115 (N_14115,N_5231,N_6068);
nand U14116 (N_14116,N_5082,N_7641);
nand U14117 (N_14117,N_7887,N_8897);
nand U14118 (N_14118,N_8099,N_7877);
xnor U14119 (N_14119,N_7786,N_8936);
xor U14120 (N_14120,N_8434,N_8856);
nand U14121 (N_14121,N_9640,N_7270);
and U14122 (N_14122,N_6756,N_6516);
or U14123 (N_14123,N_8675,N_8735);
and U14124 (N_14124,N_8233,N_8523);
or U14125 (N_14125,N_5198,N_8775);
nand U14126 (N_14126,N_7369,N_6678);
and U14127 (N_14127,N_8599,N_6092);
nor U14128 (N_14128,N_8349,N_7404);
or U14129 (N_14129,N_6114,N_6566);
xnor U14130 (N_14130,N_7380,N_9931);
xor U14131 (N_14131,N_7691,N_9857);
nor U14132 (N_14132,N_8542,N_5167);
xor U14133 (N_14133,N_9179,N_6802);
nor U14134 (N_14134,N_8644,N_6817);
nor U14135 (N_14135,N_5572,N_5469);
and U14136 (N_14136,N_8472,N_5624);
nor U14137 (N_14137,N_7365,N_8489);
nand U14138 (N_14138,N_8003,N_9201);
nor U14139 (N_14139,N_9969,N_9931);
nand U14140 (N_14140,N_8427,N_5082);
or U14141 (N_14141,N_9503,N_6092);
xor U14142 (N_14142,N_8340,N_6286);
or U14143 (N_14143,N_9901,N_6206);
and U14144 (N_14144,N_5588,N_8936);
or U14145 (N_14145,N_6654,N_7179);
or U14146 (N_14146,N_8272,N_5486);
and U14147 (N_14147,N_8939,N_8764);
nand U14148 (N_14148,N_8307,N_9001);
nand U14149 (N_14149,N_9793,N_5713);
or U14150 (N_14150,N_9766,N_7371);
nand U14151 (N_14151,N_8474,N_6952);
nor U14152 (N_14152,N_8609,N_9565);
nand U14153 (N_14153,N_9593,N_5636);
or U14154 (N_14154,N_7911,N_8274);
or U14155 (N_14155,N_7705,N_8759);
or U14156 (N_14156,N_9972,N_6063);
nor U14157 (N_14157,N_9862,N_6828);
or U14158 (N_14158,N_8120,N_7900);
xor U14159 (N_14159,N_6206,N_6624);
nand U14160 (N_14160,N_7965,N_5677);
nand U14161 (N_14161,N_9720,N_5911);
nand U14162 (N_14162,N_9690,N_6688);
and U14163 (N_14163,N_6703,N_5642);
nor U14164 (N_14164,N_8875,N_8967);
or U14165 (N_14165,N_9651,N_7602);
and U14166 (N_14166,N_5103,N_9894);
nor U14167 (N_14167,N_8401,N_9673);
or U14168 (N_14168,N_6630,N_9538);
or U14169 (N_14169,N_7239,N_5732);
nand U14170 (N_14170,N_5106,N_7164);
nor U14171 (N_14171,N_7623,N_5228);
nor U14172 (N_14172,N_7290,N_8907);
or U14173 (N_14173,N_6699,N_7801);
and U14174 (N_14174,N_5607,N_8738);
and U14175 (N_14175,N_7347,N_9465);
nor U14176 (N_14176,N_5662,N_9243);
or U14177 (N_14177,N_6899,N_7884);
nor U14178 (N_14178,N_9302,N_7818);
nor U14179 (N_14179,N_8953,N_8412);
nor U14180 (N_14180,N_8786,N_5729);
nand U14181 (N_14181,N_7377,N_6020);
nand U14182 (N_14182,N_7890,N_8813);
nand U14183 (N_14183,N_9572,N_8822);
nand U14184 (N_14184,N_6184,N_5346);
xnor U14185 (N_14185,N_5999,N_6174);
nor U14186 (N_14186,N_7851,N_6958);
nand U14187 (N_14187,N_8728,N_5607);
or U14188 (N_14188,N_7625,N_9023);
xor U14189 (N_14189,N_5120,N_7403);
or U14190 (N_14190,N_5672,N_8687);
xnor U14191 (N_14191,N_6264,N_6676);
and U14192 (N_14192,N_5962,N_8249);
xor U14193 (N_14193,N_9987,N_8435);
xor U14194 (N_14194,N_5375,N_6775);
xnor U14195 (N_14195,N_6260,N_9426);
or U14196 (N_14196,N_6638,N_5649);
nor U14197 (N_14197,N_7936,N_6992);
nor U14198 (N_14198,N_5377,N_6181);
or U14199 (N_14199,N_7912,N_5976);
nor U14200 (N_14200,N_6192,N_8276);
xor U14201 (N_14201,N_7952,N_7681);
nor U14202 (N_14202,N_6289,N_6142);
or U14203 (N_14203,N_7995,N_6343);
and U14204 (N_14204,N_5908,N_5544);
and U14205 (N_14205,N_6451,N_7239);
nor U14206 (N_14206,N_5143,N_5387);
or U14207 (N_14207,N_7560,N_8670);
and U14208 (N_14208,N_9762,N_8586);
nand U14209 (N_14209,N_8310,N_7958);
or U14210 (N_14210,N_9549,N_5874);
or U14211 (N_14211,N_7744,N_9954);
xor U14212 (N_14212,N_8025,N_7966);
nor U14213 (N_14213,N_5639,N_5406);
and U14214 (N_14214,N_9418,N_8709);
or U14215 (N_14215,N_5366,N_5912);
nand U14216 (N_14216,N_9723,N_5254);
nand U14217 (N_14217,N_6015,N_9113);
nand U14218 (N_14218,N_5616,N_5998);
nor U14219 (N_14219,N_5104,N_9514);
and U14220 (N_14220,N_6670,N_9928);
and U14221 (N_14221,N_6764,N_7360);
xnor U14222 (N_14222,N_9470,N_8174);
nor U14223 (N_14223,N_9154,N_7161);
nand U14224 (N_14224,N_8977,N_8556);
nor U14225 (N_14225,N_9747,N_6691);
xnor U14226 (N_14226,N_9923,N_8450);
nand U14227 (N_14227,N_9959,N_9461);
nand U14228 (N_14228,N_9556,N_6775);
xnor U14229 (N_14229,N_8349,N_5688);
nor U14230 (N_14230,N_6092,N_7408);
xor U14231 (N_14231,N_7939,N_6255);
or U14232 (N_14232,N_9588,N_5872);
or U14233 (N_14233,N_7888,N_9338);
or U14234 (N_14234,N_6940,N_7347);
xor U14235 (N_14235,N_6230,N_5105);
nor U14236 (N_14236,N_5635,N_7133);
xor U14237 (N_14237,N_5782,N_5215);
nor U14238 (N_14238,N_5609,N_9350);
and U14239 (N_14239,N_5802,N_8665);
or U14240 (N_14240,N_9014,N_8694);
or U14241 (N_14241,N_8671,N_5016);
xnor U14242 (N_14242,N_9385,N_9537);
and U14243 (N_14243,N_8410,N_7403);
nand U14244 (N_14244,N_7257,N_9890);
and U14245 (N_14245,N_6705,N_5303);
or U14246 (N_14246,N_6409,N_8277);
nand U14247 (N_14247,N_5495,N_9303);
nand U14248 (N_14248,N_5753,N_5809);
nand U14249 (N_14249,N_9274,N_9643);
xnor U14250 (N_14250,N_7261,N_7058);
or U14251 (N_14251,N_6024,N_5634);
nor U14252 (N_14252,N_5560,N_5220);
or U14253 (N_14253,N_5949,N_5458);
and U14254 (N_14254,N_7647,N_5282);
or U14255 (N_14255,N_6438,N_9636);
nor U14256 (N_14256,N_6786,N_5098);
nand U14257 (N_14257,N_9170,N_9281);
or U14258 (N_14258,N_7640,N_7566);
nand U14259 (N_14259,N_8778,N_7736);
xor U14260 (N_14260,N_5996,N_8389);
nor U14261 (N_14261,N_8589,N_7791);
and U14262 (N_14262,N_7905,N_8417);
nand U14263 (N_14263,N_7719,N_5634);
nand U14264 (N_14264,N_5966,N_8219);
nand U14265 (N_14265,N_6573,N_6239);
or U14266 (N_14266,N_8580,N_5913);
and U14267 (N_14267,N_6262,N_9169);
nand U14268 (N_14268,N_7477,N_8918);
and U14269 (N_14269,N_8478,N_8610);
or U14270 (N_14270,N_6080,N_8140);
and U14271 (N_14271,N_9956,N_8830);
xor U14272 (N_14272,N_6213,N_8555);
nor U14273 (N_14273,N_5062,N_7660);
xnor U14274 (N_14274,N_9742,N_9975);
nand U14275 (N_14275,N_6173,N_5241);
or U14276 (N_14276,N_8876,N_7566);
xor U14277 (N_14277,N_7003,N_7998);
nor U14278 (N_14278,N_9014,N_7915);
and U14279 (N_14279,N_5125,N_5369);
nor U14280 (N_14280,N_6101,N_8572);
nor U14281 (N_14281,N_7797,N_8956);
xor U14282 (N_14282,N_7345,N_7065);
nand U14283 (N_14283,N_6122,N_8382);
nand U14284 (N_14284,N_6171,N_8142);
nor U14285 (N_14285,N_9866,N_7505);
and U14286 (N_14286,N_9829,N_5427);
xor U14287 (N_14287,N_5313,N_7987);
xor U14288 (N_14288,N_8819,N_7872);
and U14289 (N_14289,N_9638,N_5929);
and U14290 (N_14290,N_7694,N_9346);
nand U14291 (N_14291,N_5428,N_7544);
xnor U14292 (N_14292,N_5435,N_6698);
or U14293 (N_14293,N_5146,N_9071);
nand U14294 (N_14294,N_9011,N_5797);
or U14295 (N_14295,N_6558,N_6563);
or U14296 (N_14296,N_5995,N_8911);
and U14297 (N_14297,N_9228,N_6528);
and U14298 (N_14298,N_9582,N_5102);
and U14299 (N_14299,N_8649,N_7594);
and U14300 (N_14300,N_5008,N_8430);
or U14301 (N_14301,N_5879,N_5729);
or U14302 (N_14302,N_7633,N_5007);
nor U14303 (N_14303,N_8503,N_9302);
nand U14304 (N_14304,N_9577,N_9970);
and U14305 (N_14305,N_5012,N_9576);
or U14306 (N_14306,N_7233,N_6535);
or U14307 (N_14307,N_9430,N_5221);
xnor U14308 (N_14308,N_6390,N_8657);
and U14309 (N_14309,N_5561,N_6678);
nor U14310 (N_14310,N_5595,N_5926);
xor U14311 (N_14311,N_5068,N_6521);
nand U14312 (N_14312,N_6315,N_5111);
or U14313 (N_14313,N_6218,N_5170);
or U14314 (N_14314,N_7168,N_9108);
nand U14315 (N_14315,N_7526,N_9519);
nand U14316 (N_14316,N_7472,N_9981);
nor U14317 (N_14317,N_8546,N_5028);
and U14318 (N_14318,N_6099,N_8606);
and U14319 (N_14319,N_9520,N_8885);
nand U14320 (N_14320,N_8426,N_6121);
xor U14321 (N_14321,N_7853,N_6310);
nor U14322 (N_14322,N_6743,N_5656);
xor U14323 (N_14323,N_8792,N_7673);
and U14324 (N_14324,N_8277,N_5661);
nand U14325 (N_14325,N_6923,N_5443);
and U14326 (N_14326,N_9636,N_8331);
nand U14327 (N_14327,N_8406,N_9510);
xnor U14328 (N_14328,N_8238,N_5766);
and U14329 (N_14329,N_7166,N_5517);
nor U14330 (N_14330,N_5501,N_9067);
nand U14331 (N_14331,N_8714,N_8344);
nand U14332 (N_14332,N_6483,N_9709);
nor U14333 (N_14333,N_5528,N_9915);
nor U14334 (N_14334,N_6437,N_5288);
and U14335 (N_14335,N_9173,N_5884);
and U14336 (N_14336,N_9072,N_8476);
nor U14337 (N_14337,N_8276,N_7464);
nand U14338 (N_14338,N_6960,N_9919);
or U14339 (N_14339,N_6757,N_9544);
xor U14340 (N_14340,N_8474,N_8026);
nor U14341 (N_14341,N_8150,N_9854);
or U14342 (N_14342,N_6561,N_6689);
nand U14343 (N_14343,N_6347,N_7858);
and U14344 (N_14344,N_7878,N_9592);
and U14345 (N_14345,N_5011,N_8748);
nor U14346 (N_14346,N_8660,N_8510);
or U14347 (N_14347,N_8488,N_6068);
xor U14348 (N_14348,N_9881,N_7313);
nand U14349 (N_14349,N_6799,N_6076);
and U14350 (N_14350,N_6390,N_7090);
nand U14351 (N_14351,N_5924,N_5606);
or U14352 (N_14352,N_5222,N_9517);
and U14353 (N_14353,N_7756,N_7713);
nor U14354 (N_14354,N_5378,N_7457);
nand U14355 (N_14355,N_5600,N_6455);
or U14356 (N_14356,N_6661,N_9105);
nor U14357 (N_14357,N_8484,N_5568);
nor U14358 (N_14358,N_9858,N_8563);
or U14359 (N_14359,N_7258,N_6297);
and U14360 (N_14360,N_5252,N_9397);
nor U14361 (N_14361,N_7300,N_8335);
nor U14362 (N_14362,N_5447,N_9895);
xor U14363 (N_14363,N_7227,N_5985);
xor U14364 (N_14364,N_5573,N_8001);
nand U14365 (N_14365,N_8519,N_8205);
nor U14366 (N_14366,N_6885,N_7973);
xnor U14367 (N_14367,N_9460,N_5828);
xnor U14368 (N_14368,N_9012,N_9380);
and U14369 (N_14369,N_5496,N_5657);
nor U14370 (N_14370,N_8827,N_9767);
or U14371 (N_14371,N_5395,N_5524);
or U14372 (N_14372,N_6904,N_7855);
xnor U14373 (N_14373,N_5528,N_7544);
or U14374 (N_14374,N_9795,N_5793);
xor U14375 (N_14375,N_8689,N_8317);
nand U14376 (N_14376,N_7181,N_8370);
and U14377 (N_14377,N_5623,N_5524);
nand U14378 (N_14378,N_7583,N_6813);
xnor U14379 (N_14379,N_6042,N_6933);
and U14380 (N_14380,N_7699,N_8482);
nand U14381 (N_14381,N_5627,N_7136);
xor U14382 (N_14382,N_8528,N_8908);
and U14383 (N_14383,N_6826,N_5371);
nand U14384 (N_14384,N_7292,N_8377);
xnor U14385 (N_14385,N_7769,N_5661);
or U14386 (N_14386,N_8752,N_6348);
nand U14387 (N_14387,N_5864,N_6269);
nand U14388 (N_14388,N_7290,N_9308);
nor U14389 (N_14389,N_9189,N_9160);
nand U14390 (N_14390,N_7875,N_7588);
xor U14391 (N_14391,N_9335,N_6236);
nor U14392 (N_14392,N_6066,N_5262);
xor U14393 (N_14393,N_7151,N_6294);
and U14394 (N_14394,N_9567,N_5015);
nor U14395 (N_14395,N_8636,N_7453);
xor U14396 (N_14396,N_8915,N_7211);
or U14397 (N_14397,N_9410,N_8471);
xor U14398 (N_14398,N_7003,N_5502);
and U14399 (N_14399,N_8311,N_6891);
or U14400 (N_14400,N_5216,N_6156);
nor U14401 (N_14401,N_6911,N_9769);
and U14402 (N_14402,N_7860,N_6390);
nor U14403 (N_14403,N_5525,N_9059);
and U14404 (N_14404,N_8023,N_6685);
nor U14405 (N_14405,N_5966,N_5160);
xor U14406 (N_14406,N_8108,N_7412);
xnor U14407 (N_14407,N_6796,N_5905);
or U14408 (N_14408,N_8679,N_9095);
xnor U14409 (N_14409,N_8522,N_6740);
or U14410 (N_14410,N_6975,N_6937);
xor U14411 (N_14411,N_7682,N_7831);
and U14412 (N_14412,N_6626,N_9285);
and U14413 (N_14413,N_5906,N_9541);
or U14414 (N_14414,N_6382,N_7688);
or U14415 (N_14415,N_9280,N_5165);
and U14416 (N_14416,N_7970,N_7914);
and U14417 (N_14417,N_7989,N_5465);
nand U14418 (N_14418,N_7241,N_7322);
and U14419 (N_14419,N_8133,N_6668);
or U14420 (N_14420,N_9863,N_7616);
nor U14421 (N_14421,N_8679,N_7214);
and U14422 (N_14422,N_5087,N_5623);
xnor U14423 (N_14423,N_9515,N_5555);
nand U14424 (N_14424,N_9889,N_5639);
and U14425 (N_14425,N_8126,N_7931);
and U14426 (N_14426,N_6809,N_9508);
nor U14427 (N_14427,N_9494,N_8783);
xor U14428 (N_14428,N_6301,N_6118);
nor U14429 (N_14429,N_5167,N_5595);
nand U14430 (N_14430,N_8094,N_5421);
or U14431 (N_14431,N_8900,N_5735);
nand U14432 (N_14432,N_7683,N_8915);
and U14433 (N_14433,N_7612,N_8565);
nor U14434 (N_14434,N_7085,N_6648);
nor U14435 (N_14435,N_7184,N_5157);
xnor U14436 (N_14436,N_6311,N_8683);
xor U14437 (N_14437,N_7614,N_7547);
or U14438 (N_14438,N_9570,N_7141);
nand U14439 (N_14439,N_7985,N_9826);
xnor U14440 (N_14440,N_6893,N_6117);
and U14441 (N_14441,N_7727,N_5008);
nor U14442 (N_14442,N_9804,N_8909);
nor U14443 (N_14443,N_7982,N_9228);
and U14444 (N_14444,N_9817,N_7631);
or U14445 (N_14445,N_8693,N_9238);
xor U14446 (N_14446,N_6634,N_6742);
nor U14447 (N_14447,N_6683,N_9370);
or U14448 (N_14448,N_7281,N_9169);
xor U14449 (N_14449,N_5238,N_9999);
nor U14450 (N_14450,N_6277,N_8993);
or U14451 (N_14451,N_7871,N_9066);
and U14452 (N_14452,N_8698,N_5229);
or U14453 (N_14453,N_7943,N_8326);
nand U14454 (N_14454,N_5762,N_7543);
nor U14455 (N_14455,N_6774,N_8267);
xor U14456 (N_14456,N_9156,N_7986);
xor U14457 (N_14457,N_8555,N_9575);
xor U14458 (N_14458,N_7469,N_9521);
or U14459 (N_14459,N_7722,N_6091);
nor U14460 (N_14460,N_6211,N_7165);
xor U14461 (N_14461,N_7707,N_8223);
nand U14462 (N_14462,N_8600,N_6710);
nor U14463 (N_14463,N_9850,N_6969);
and U14464 (N_14464,N_7783,N_5864);
xor U14465 (N_14465,N_8452,N_6071);
nand U14466 (N_14466,N_6200,N_7764);
nand U14467 (N_14467,N_5489,N_8352);
nor U14468 (N_14468,N_8651,N_7166);
xnor U14469 (N_14469,N_5656,N_5263);
xor U14470 (N_14470,N_8357,N_8072);
nor U14471 (N_14471,N_7472,N_6001);
or U14472 (N_14472,N_5615,N_6656);
nand U14473 (N_14473,N_5921,N_8118);
and U14474 (N_14474,N_9540,N_6717);
nand U14475 (N_14475,N_5558,N_9967);
nand U14476 (N_14476,N_5622,N_5334);
xor U14477 (N_14477,N_6948,N_8476);
nor U14478 (N_14478,N_5128,N_9121);
nand U14479 (N_14479,N_8289,N_6142);
nand U14480 (N_14480,N_8320,N_6361);
or U14481 (N_14481,N_8775,N_9342);
xor U14482 (N_14482,N_5793,N_6901);
and U14483 (N_14483,N_6072,N_9586);
xnor U14484 (N_14484,N_5838,N_6516);
or U14485 (N_14485,N_6535,N_8586);
or U14486 (N_14486,N_9681,N_5146);
nand U14487 (N_14487,N_9391,N_6104);
and U14488 (N_14488,N_7001,N_5187);
nor U14489 (N_14489,N_8216,N_6564);
or U14490 (N_14490,N_8551,N_5387);
or U14491 (N_14491,N_5655,N_6011);
nand U14492 (N_14492,N_6945,N_6553);
nand U14493 (N_14493,N_6033,N_9812);
xnor U14494 (N_14494,N_7273,N_8530);
and U14495 (N_14495,N_8865,N_6046);
and U14496 (N_14496,N_7379,N_8942);
nor U14497 (N_14497,N_5956,N_8894);
or U14498 (N_14498,N_8920,N_8558);
nor U14499 (N_14499,N_7039,N_5392);
nor U14500 (N_14500,N_8683,N_5113);
xnor U14501 (N_14501,N_5339,N_5195);
nor U14502 (N_14502,N_6669,N_5211);
xnor U14503 (N_14503,N_9114,N_8271);
xor U14504 (N_14504,N_9875,N_7846);
and U14505 (N_14505,N_9495,N_9781);
xnor U14506 (N_14506,N_5871,N_7191);
xor U14507 (N_14507,N_8643,N_8973);
and U14508 (N_14508,N_9021,N_9030);
or U14509 (N_14509,N_6051,N_7059);
or U14510 (N_14510,N_6890,N_9734);
nor U14511 (N_14511,N_9650,N_7691);
nor U14512 (N_14512,N_5995,N_8359);
xor U14513 (N_14513,N_8783,N_8657);
and U14514 (N_14514,N_7023,N_5171);
nor U14515 (N_14515,N_7710,N_7394);
nor U14516 (N_14516,N_8439,N_5091);
xnor U14517 (N_14517,N_9856,N_6246);
nand U14518 (N_14518,N_8702,N_9523);
and U14519 (N_14519,N_8306,N_7988);
and U14520 (N_14520,N_5981,N_6899);
nand U14521 (N_14521,N_7531,N_7052);
and U14522 (N_14522,N_8203,N_9663);
nand U14523 (N_14523,N_8486,N_6134);
or U14524 (N_14524,N_6002,N_8539);
nor U14525 (N_14525,N_6374,N_5781);
or U14526 (N_14526,N_9012,N_5670);
nor U14527 (N_14527,N_8276,N_6039);
nor U14528 (N_14528,N_6177,N_6697);
nand U14529 (N_14529,N_7549,N_8742);
nand U14530 (N_14530,N_8782,N_7491);
nand U14531 (N_14531,N_7505,N_6544);
or U14532 (N_14532,N_5844,N_7453);
and U14533 (N_14533,N_9014,N_9703);
and U14534 (N_14534,N_9909,N_8349);
nand U14535 (N_14535,N_5079,N_9917);
and U14536 (N_14536,N_8853,N_8438);
nand U14537 (N_14537,N_6460,N_6613);
nor U14538 (N_14538,N_6821,N_9332);
nand U14539 (N_14539,N_6900,N_7682);
xor U14540 (N_14540,N_7991,N_9648);
or U14541 (N_14541,N_9107,N_6327);
or U14542 (N_14542,N_5519,N_5749);
xnor U14543 (N_14543,N_8026,N_9601);
nor U14544 (N_14544,N_9269,N_8360);
nand U14545 (N_14545,N_9877,N_8472);
and U14546 (N_14546,N_7535,N_7129);
nor U14547 (N_14547,N_6875,N_5383);
nand U14548 (N_14548,N_7798,N_7849);
nor U14549 (N_14549,N_6887,N_9125);
nand U14550 (N_14550,N_6052,N_7021);
xor U14551 (N_14551,N_7882,N_6198);
or U14552 (N_14552,N_7179,N_8280);
and U14553 (N_14553,N_9696,N_6213);
or U14554 (N_14554,N_8895,N_9342);
nand U14555 (N_14555,N_5988,N_7355);
or U14556 (N_14556,N_9252,N_6871);
nor U14557 (N_14557,N_8538,N_9131);
or U14558 (N_14558,N_5441,N_5826);
or U14559 (N_14559,N_7453,N_6137);
xor U14560 (N_14560,N_7018,N_5572);
or U14561 (N_14561,N_5344,N_9478);
or U14562 (N_14562,N_9795,N_6605);
or U14563 (N_14563,N_6647,N_7859);
xor U14564 (N_14564,N_8438,N_8755);
or U14565 (N_14565,N_6118,N_7672);
xnor U14566 (N_14566,N_9665,N_5685);
or U14567 (N_14567,N_6856,N_9945);
or U14568 (N_14568,N_6352,N_5198);
nand U14569 (N_14569,N_9106,N_8706);
and U14570 (N_14570,N_5765,N_8586);
or U14571 (N_14571,N_9215,N_9219);
or U14572 (N_14572,N_9667,N_5318);
or U14573 (N_14573,N_7888,N_7919);
xnor U14574 (N_14574,N_7238,N_8875);
or U14575 (N_14575,N_5746,N_5533);
nand U14576 (N_14576,N_8955,N_8254);
and U14577 (N_14577,N_6909,N_7120);
or U14578 (N_14578,N_9830,N_5122);
or U14579 (N_14579,N_5768,N_8962);
or U14580 (N_14580,N_8992,N_8045);
or U14581 (N_14581,N_5725,N_5976);
and U14582 (N_14582,N_9484,N_8605);
xnor U14583 (N_14583,N_6641,N_8746);
and U14584 (N_14584,N_6997,N_5479);
xnor U14585 (N_14585,N_5861,N_6894);
xor U14586 (N_14586,N_9973,N_6730);
or U14587 (N_14587,N_5225,N_9638);
and U14588 (N_14588,N_5080,N_8233);
nand U14589 (N_14589,N_8341,N_6501);
xnor U14590 (N_14590,N_9703,N_9939);
nand U14591 (N_14591,N_6235,N_7484);
and U14592 (N_14592,N_5503,N_8863);
xnor U14593 (N_14593,N_6269,N_5389);
and U14594 (N_14594,N_9085,N_8364);
and U14595 (N_14595,N_7599,N_6114);
and U14596 (N_14596,N_8908,N_5512);
nor U14597 (N_14597,N_8324,N_7251);
xor U14598 (N_14598,N_6584,N_5826);
or U14599 (N_14599,N_5179,N_8865);
nor U14600 (N_14600,N_8629,N_8734);
and U14601 (N_14601,N_7832,N_9267);
xor U14602 (N_14602,N_5177,N_8845);
or U14603 (N_14603,N_7432,N_7304);
or U14604 (N_14604,N_6795,N_9139);
or U14605 (N_14605,N_5267,N_5060);
or U14606 (N_14606,N_5041,N_8722);
and U14607 (N_14607,N_5898,N_7492);
nor U14608 (N_14608,N_9746,N_6247);
or U14609 (N_14609,N_9501,N_7872);
nand U14610 (N_14610,N_9885,N_6830);
xnor U14611 (N_14611,N_7106,N_7186);
or U14612 (N_14612,N_8753,N_8274);
and U14613 (N_14613,N_6963,N_7118);
xnor U14614 (N_14614,N_5512,N_6007);
or U14615 (N_14615,N_8345,N_5619);
and U14616 (N_14616,N_7397,N_6592);
or U14617 (N_14617,N_5367,N_5044);
or U14618 (N_14618,N_5990,N_6128);
xnor U14619 (N_14619,N_9575,N_9875);
and U14620 (N_14620,N_6606,N_8883);
nor U14621 (N_14621,N_9640,N_6477);
nand U14622 (N_14622,N_9203,N_9213);
and U14623 (N_14623,N_8409,N_8634);
and U14624 (N_14624,N_6001,N_9189);
nand U14625 (N_14625,N_6264,N_5732);
or U14626 (N_14626,N_5360,N_9549);
or U14627 (N_14627,N_6992,N_9151);
and U14628 (N_14628,N_8077,N_9461);
nand U14629 (N_14629,N_5412,N_6006);
or U14630 (N_14630,N_8784,N_6549);
nor U14631 (N_14631,N_9276,N_7969);
and U14632 (N_14632,N_8393,N_6654);
and U14633 (N_14633,N_5691,N_6276);
nand U14634 (N_14634,N_9293,N_8540);
or U14635 (N_14635,N_5994,N_9471);
nor U14636 (N_14636,N_5883,N_9105);
and U14637 (N_14637,N_6268,N_5797);
nor U14638 (N_14638,N_9994,N_9788);
xor U14639 (N_14639,N_8125,N_5045);
and U14640 (N_14640,N_5211,N_5314);
nand U14641 (N_14641,N_7764,N_9125);
nand U14642 (N_14642,N_9303,N_5168);
xor U14643 (N_14643,N_9243,N_9690);
xnor U14644 (N_14644,N_8878,N_5009);
nand U14645 (N_14645,N_9413,N_6727);
and U14646 (N_14646,N_6111,N_7945);
nor U14647 (N_14647,N_6750,N_9623);
xor U14648 (N_14648,N_8523,N_5423);
xor U14649 (N_14649,N_5640,N_7504);
nand U14650 (N_14650,N_6620,N_9681);
and U14651 (N_14651,N_5364,N_6523);
and U14652 (N_14652,N_7859,N_5724);
nor U14653 (N_14653,N_9100,N_5715);
or U14654 (N_14654,N_6646,N_5061);
or U14655 (N_14655,N_8376,N_5248);
and U14656 (N_14656,N_9324,N_7234);
nand U14657 (N_14657,N_7316,N_5633);
xnor U14658 (N_14658,N_5426,N_5935);
and U14659 (N_14659,N_5508,N_6425);
nor U14660 (N_14660,N_9819,N_9378);
and U14661 (N_14661,N_6799,N_5217);
nor U14662 (N_14662,N_6771,N_8849);
and U14663 (N_14663,N_6313,N_5971);
or U14664 (N_14664,N_8094,N_5016);
xnor U14665 (N_14665,N_9980,N_5115);
nor U14666 (N_14666,N_9313,N_7434);
nand U14667 (N_14667,N_9049,N_9381);
nand U14668 (N_14668,N_5546,N_6343);
and U14669 (N_14669,N_9230,N_9878);
or U14670 (N_14670,N_8066,N_7173);
nor U14671 (N_14671,N_6784,N_7713);
xnor U14672 (N_14672,N_8898,N_8420);
xnor U14673 (N_14673,N_7765,N_9190);
nor U14674 (N_14674,N_6847,N_6455);
nand U14675 (N_14675,N_6724,N_5445);
nand U14676 (N_14676,N_6002,N_5003);
and U14677 (N_14677,N_7267,N_9060);
xnor U14678 (N_14678,N_9931,N_6422);
nand U14679 (N_14679,N_7640,N_5891);
and U14680 (N_14680,N_5969,N_5547);
xor U14681 (N_14681,N_5353,N_8330);
nand U14682 (N_14682,N_7529,N_7835);
xor U14683 (N_14683,N_6865,N_8332);
or U14684 (N_14684,N_8155,N_9029);
xor U14685 (N_14685,N_9854,N_8795);
xnor U14686 (N_14686,N_9781,N_8406);
nand U14687 (N_14687,N_6326,N_8338);
and U14688 (N_14688,N_5705,N_8788);
and U14689 (N_14689,N_5605,N_5732);
and U14690 (N_14690,N_8740,N_8609);
or U14691 (N_14691,N_8243,N_5718);
nand U14692 (N_14692,N_9694,N_5144);
xor U14693 (N_14693,N_5519,N_7704);
and U14694 (N_14694,N_5046,N_8292);
or U14695 (N_14695,N_9407,N_9622);
nand U14696 (N_14696,N_9248,N_8915);
xor U14697 (N_14697,N_9471,N_8055);
xnor U14698 (N_14698,N_8950,N_9440);
and U14699 (N_14699,N_5807,N_9688);
and U14700 (N_14700,N_5686,N_8951);
xnor U14701 (N_14701,N_6847,N_9857);
nand U14702 (N_14702,N_5271,N_8303);
xnor U14703 (N_14703,N_7572,N_6539);
or U14704 (N_14704,N_9270,N_9888);
nand U14705 (N_14705,N_8886,N_6912);
xor U14706 (N_14706,N_7110,N_9730);
xor U14707 (N_14707,N_5152,N_5289);
or U14708 (N_14708,N_6525,N_6262);
xnor U14709 (N_14709,N_6705,N_8531);
xor U14710 (N_14710,N_8316,N_9782);
xnor U14711 (N_14711,N_5358,N_9122);
or U14712 (N_14712,N_9525,N_8427);
or U14713 (N_14713,N_8878,N_9495);
nor U14714 (N_14714,N_7089,N_8644);
nand U14715 (N_14715,N_5173,N_7135);
nor U14716 (N_14716,N_7062,N_6619);
nor U14717 (N_14717,N_6858,N_9615);
and U14718 (N_14718,N_8319,N_7571);
nor U14719 (N_14719,N_7980,N_9476);
and U14720 (N_14720,N_9992,N_5653);
and U14721 (N_14721,N_5941,N_5958);
nand U14722 (N_14722,N_7036,N_9700);
and U14723 (N_14723,N_8243,N_7433);
xnor U14724 (N_14724,N_7763,N_7087);
xor U14725 (N_14725,N_7215,N_9332);
nand U14726 (N_14726,N_6505,N_5851);
nor U14727 (N_14727,N_8002,N_7505);
nor U14728 (N_14728,N_6390,N_9803);
xnor U14729 (N_14729,N_7110,N_9847);
nor U14730 (N_14730,N_5326,N_6752);
and U14731 (N_14731,N_5644,N_8675);
and U14732 (N_14732,N_5976,N_6562);
or U14733 (N_14733,N_5298,N_9884);
xnor U14734 (N_14734,N_9703,N_7848);
nor U14735 (N_14735,N_7009,N_5807);
nor U14736 (N_14736,N_9259,N_6177);
and U14737 (N_14737,N_8382,N_7192);
nand U14738 (N_14738,N_5689,N_6918);
and U14739 (N_14739,N_6931,N_5348);
and U14740 (N_14740,N_9381,N_6379);
nand U14741 (N_14741,N_6304,N_7926);
or U14742 (N_14742,N_6864,N_7190);
nor U14743 (N_14743,N_7158,N_5209);
and U14744 (N_14744,N_5024,N_7467);
and U14745 (N_14745,N_6885,N_6135);
and U14746 (N_14746,N_8483,N_5446);
nand U14747 (N_14747,N_5503,N_7133);
nand U14748 (N_14748,N_8473,N_5735);
or U14749 (N_14749,N_5634,N_8365);
nor U14750 (N_14750,N_9538,N_6988);
and U14751 (N_14751,N_8955,N_8359);
xnor U14752 (N_14752,N_5938,N_8894);
xnor U14753 (N_14753,N_8824,N_5067);
or U14754 (N_14754,N_6974,N_6540);
nor U14755 (N_14755,N_7018,N_9025);
and U14756 (N_14756,N_6541,N_6368);
nor U14757 (N_14757,N_6021,N_5053);
nor U14758 (N_14758,N_6520,N_5446);
xnor U14759 (N_14759,N_8984,N_6294);
xor U14760 (N_14760,N_8810,N_9901);
nor U14761 (N_14761,N_5131,N_6152);
nor U14762 (N_14762,N_6410,N_7689);
and U14763 (N_14763,N_9316,N_7172);
nand U14764 (N_14764,N_6617,N_9250);
nand U14765 (N_14765,N_8617,N_5685);
or U14766 (N_14766,N_8721,N_8573);
nand U14767 (N_14767,N_9232,N_5499);
nand U14768 (N_14768,N_6023,N_9190);
nand U14769 (N_14769,N_6407,N_9879);
and U14770 (N_14770,N_7555,N_5409);
nor U14771 (N_14771,N_5098,N_9907);
and U14772 (N_14772,N_7011,N_6408);
nor U14773 (N_14773,N_5453,N_8905);
or U14774 (N_14774,N_9554,N_8303);
nand U14775 (N_14775,N_7350,N_8174);
nand U14776 (N_14776,N_5315,N_9707);
xnor U14777 (N_14777,N_5410,N_5654);
xnor U14778 (N_14778,N_8170,N_7955);
nor U14779 (N_14779,N_9454,N_8133);
nand U14780 (N_14780,N_6250,N_7478);
nor U14781 (N_14781,N_9376,N_6553);
nand U14782 (N_14782,N_9350,N_6804);
xor U14783 (N_14783,N_5466,N_8231);
and U14784 (N_14784,N_8903,N_6049);
nor U14785 (N_14785,N_8898,N_5720);
nand U14786 (N_14786,N_8862,N_7005);
xnor U14787 (N_14787,N_6842,N_5580);
and U14788 (N_14788,N_6507,N_6611);
nor U14789 (N_14789,N_5308,N_6385);
nand U14790 (N_14790,N_5560,N_6919);
and U14791 (N_14791,N_9813,N_8040);
or U14792 (N_14792,N_8608,N_9280);
or U14793 (N_14793,N_7631,N_6991);
or U14794 (N_14794,N_7211,N_5580);
or U14795 (N_14795,N_5868,N_5604);
nor U14796 (N_14796,N_9889,N_5409);
nand U14797 (N_14797,N_8202,N_5930);
xnor U14798 (N_14798,N_7451,N_6129);
and U14799 (N_14799,N_5229,N_7855);
or U14800 (N_14800,N_7147,N_7941);
or U14801 (N_14801,N_7718,N_6955);
nand U14802 (N_14802,N_6378,N_6690);
and U14803 (N_14803,N_8393,N_7020);
or U14804 (N_14804,N_9176,N_6009);
nand U14805 (N_14805,N_7306,N_8747);
nor U14806 (N_14806,N_9232,N_9527);
nand U14807 (N_14807,N_9749,N_7123);
nor U14808 (N_14808,N_8315,N_6608);
or U14809 (N_14809,N_9478,N_6903);
nand U14810 (N_14810,N_9206,N_6500);
xor U14811 (N_14811,N_6730,N_7521);
and U14812 (N_14812,N_5751,N_5253);
nand U14813 (N_14813,N_8420,N_7458);
nand U14814 (N_14814,N_7154,N_7877);
nand U14815 (N_14815,N_5266,N_7019);
xnor U14816 (N_14816,N_5297,N_9720);
nor U14817 (N_14817,N_8444,N_9649);
xnor U14818 (N_14818,N_7269,N_8578);
xor U14819 (N_14819,N_7571,N_7261);
or U14820 (N_14820,N_6048,N_5792);
nand U14821 (N_14821,N_8788,N_5690);
xor U14822 (N_14822,N_8800,N_7935);
nand U14823 (N_14823,N_8344,N_6207);
nand U14824 (N_14824,N_6062,N_6921);
xor U14825 (N_14825,N_6621,N_6973);
nand U14826 (N_14826,N_9565,N_5768);
nor U14827 (N_14827,N_6741,N_6916);
or U14828 (N_14828,N_6699,N_7082);
xnor U14829 (N_14829,N_6208,N_9089);
nand U14830 (N_14830,N_7422,N_6663);
nor U14831 (N_14831,N_7038,N_8153);
xnor U14832 (N_14832,N_5138,N_8169);
nor U14833 (N_14833,N_7024,N_5321);
nand U14834 (N_14834,N_9374,N_5976);
or U14835 (N_14835,N_5245,N_9006);
or U14836 (N_14836,N_8094,N_9978);
nor U14837 (N_14837,N_6398,N_8966);
or U14838 (N_14838,N_5800,N_6336);
nor U14839 (N_14839,N_7701,N_9316);
nand U14840 (N_14840,N_5527,N_8174);
or U14841 (N_14841,N_9236,N_7436);
xor U14842 (N_14842,N_7225,N_7064);
nand U14843 (N_14843,N_5495,N_8840);
nor U14844 (N_14844,N_6506,N_6018);
or U14845 (N_14845,N_9575,N_6346);
nand U14846 (N_14846,N_7692,N_8296);
nor U14847 (N_14847,N_7950,N_5501);
nor U14848 (N_14848,N_6436,N_6932);
and U14849 (N_14849,N_6694,N_5125);
nand U14850 (N_14850,N_9915,N_9179);
xnor U14851 (N_14851,N_6885,N_7900);
and U14852 (N_14852,N_7319,N_6669);
nand U14853 (N_14853,N_5749,N_9693);
or U14854 (N_14854,N_9224,N_8012);
nor U14855 (N_14855,N_8970,N_5851);
or U14856 (N_14856,N_8586,N_9345);
nand U14857 (N_14857,N_7015,N_5302);
and U14858 (N_14858,N_5734,N_8253);
and U14859 (N_14859,N_5181,N_7376);
and U14860 (N_14860,N_5198,N_6268);
nand U14861 (N_14861,N_6624,N_9373);
nor U14862 (N_14862,N_9571,N_8177);
and U14863 (N_14863,N_5582,N_9552);
and U14864 (N_14864,N_6102,N_6205);
xnor U14865 (N_14865,N_9778,N_5870);
and U14866 (N_14866,N_8371,N_9354);
xnor U14867 (N_14867,N_5546,N_6782);
and U14868 (N_14868,N_9381,N_5642);
xnor U14869 (N_14869,N_5554,N_6470);
and U14870 (N_14870,N_9309,N_7117);
and U14871 (N_14871,N_7234,N_8068);
and U14872 (N_14872,N_7185,N_9641);
nand U14873 (N_14873,N_7762,N_9155);
xor U14874 (N_14874,N_6065,N_6654);
xor U14875 (N_14875,N_7226,N_5956);
xnor U14876 (N_14876,N_5356,N_8632);
and U14877 (N_14877,N_5049,N_6163);
xor U14878 (N_14878,N_6305,N_6072);
nand U14879 (N_14879,N_6067,N_5680);
nor U14880 (N_14880,N_8520,N_7673);
nor U14881 (N_14881,N_7994,N_5136);
nand U14882 (N_14882,N_8779,N_9174);
nor U14883 (N_14883,N_6413,N_5064);
xnor U14884 (N_14884,N_7011,N_6207);
and U14885 (N_14885,N_6450,N_9731);
nor U14886 (N_14886,N_9740,N_7614);
xor U14887 (N_14887,N_6569,N_8262);
xor U14888 (N_14888,N_8721,N_6283);
or U14889 (N_14889,N_7154,N_5933);
xor U14890 (N_14890,N_9194,N_9311);
and U14891 (N_14891,N_8650,N_9030);
or U14892 (N_14892,N_7423,N_6146);
or U14893 (N_14893,N_8639,N_7126);
xnor U14894 (N_14894,N_7108,N_8907);
or U14895 (N_14895,N_5187,N_9546);
nor U14896 (N_14896,N_7941,N_8580);
or U14897 (N_14897,N_8295,N_8164);
nand U14898 (N_14898,N_9053,N_8854);
nand U14899 (N_14899,N_5291,N_8634);
or U14900 (N_14900,N_9211,N_7053);
nor U14901 (N_14901,N_5934,N_5167);
nand U14902 (N_14902,N_9368,N_5036);
or U14903 (N_14903,N_7564,N_6579);
xnor U14904 (N_14904,N_5352,N_6240);
or U14905 (N_14905,N_9844,N_8279);
or U14906 (N_14906,N_5625,N_9799);
or U14907 (N_14907,N_7193,N_9751);
or U14908 (N_14908,N_8426,N_8977);
nor U14909 (N_14909,N_8088,N_7256);
and U14910 (N_14910,N_6352,N_5392);
nor U14911 (N_14911,N_6962,N_8189);
or U14912 (N_14912,N_9370,N_8590);
nand U14913 (N_14913,N_5759,N_9251);
nor U14914 (N_14914,N_6947,N_8582);
nor U14915 (N_14915,N_6187,N_6238);
nor U14916 (N_14916,N_9783,N_7746);
nor U14917 (N_14917,N_9449,N_5328);
xnor U14918 (N_14918,N_7118,N_5832);
nor U14919 (N_14919,N_9215,N_8065);
and U14920 (N_14920,N_9372,N_7820);
nor U14921 (N_14921,N_8729,N_9959);
and U14922 (N_14922,N_8683,N_8260);
xor U14923 (N_14923,N_8353,N_8168);
and U14924 (N_14924,N_9891,N_7193);
or U14925 (N_14925,N_8083,N_6715);
xor U14926 (N_14926,N_7104,N_6893);
nand U14927 (N_14927,N_9126,N_5582);
xnor U14928 (N_14928,N_8472,N_5021);
and U14929 (N_14929,N_6713,N_8182);
and U14930 (N_14930,N_7839,N_9327);
nor U14931 (N_14931,N_9472,N_9631);
nor U14932 (N_14932,N_9026,N_6891);
and U14933 (N_14933,N_9923,N_7171);
nand U14934 (N_14934,N_5122,N_7841);
xor U14935 (N_14935,N_8135,N_9787);
and U14936 (N_14936,N_5357,N_7126);
nand U14937 (N_14937,N_9171,N_7699);
nor U14938 (N_14938,N_7083,N_8752);
and U14939 (N_14939,N_8597,N_5706);
nand U14940 (N_14940,N_5221,N_9322);
or U14941 (N_14941,N_9207,N_7961);
and U14942 (N_14942,N_7049,N_5092);
nand U14943 (N_14943,N_5269,N_7863);
nand U14944 (N_14944,N_9470,N_5550);
and U14945 (N_14945,N_5761,N_9936);
or U14946 (N_14946,N_6017,N_5031);
and U14947 (N_14947,N_8709,N_5909);
xnor U14948 (N_14948,N_8600,N_5556);
nand U14949 (N_14949,N_7655,N_5901);
nor U14950 (N_14950,N_5645,N_8508);
and U14951 (N_14951,N_9865,N_5715);
nand U14952 (N_14952,N_9478,N_8862);
nand U14953 (N_14953,N_6923,N_8333);
nor U14954 (N_14954,N_6444,N_8500);
or U14955 (N_14955,N_5992,N_7701);
and U14956 (N_14956,N_8781,N_5636);
nand U14957 (N_14957,N_9397,N_5095);
nand U14958 (N_14958,N_9700,N_5244);
or U14959 (N_14959,N_5719,N_8685);
or U14960 (N_14960,N_7481,N_9472);
xnor U14961 (N_14961,N_9241,N_9170);
xor U14962 (N_14962,N_8342,N_8152);
or U14963 (N_14963,N_9815,N_5995);
nor U14964 (N_14964,N_9296,N_5430);
xor U14965 (N_14965,N_9370,N_9148);
nand U14966 (N_14966,N_7792,N_5313);
or U14967 (N_14967,N_8562,N_7072);
or U14968 (N_14968,N_8052,N_7033);
xnor U14969 (N_14969,N_6576,N_7779);
xor U14970 (N_14970,N_5230,N_6623);
nor U14971 (N_14971,N_7606,N_6488);
nand U14972 (N_14972,N_7002,N_7405);
xnor U14973 (N_14973,N_7989,N_7426);
or U14974 (N_14974,N_7687,N_7158);
xnor U14975 (N_14975,N_8783,N_9434);
nor U14976 (N_14976,N_8301,N_6044);
and U14977 (N_14977,N_8442,N_6426);
or U14978 (N_14978,N_7063,N_8260);
or U14979 (N_14979,N_7760,N_6722);
and U14980 (N_14980,N_5560,N_8477);
or U14981 (N_14981,N_8629,N_5958);
nand U14982 (N_14982,N_6666,N_9467);
nand U14983 (N_14983,N_8231,N_8449);
and U14984 (N_14984,N_8196,N_5993);
and U14985 (N_14985,N_9016,N_6534);
nand U14986 (N_14986,N_5329,N_5203);
nand U14987 (N_14987,N_6994,N_7531);
nand U14988 (N_14988,N_6296,N_9621);
xnor U14989 (N_14989,N_6623,N_9878);
nor U14990 (N_14990,N_8981,N_6006);
nor U14991 (N_14991,N_7892,N_6599);
nor U14992 (N_14992,N_6978,N_8283);
or U14993 (N_14993,N_9945,N_9643);
nand U14994 (N_14994,N_8058,N_6440);
xor U14995 (N_14995,N_9613,N_8605);
xor U14996 (N_14996,N_8873,N_5323);
nand U14997 (N_14997,N_7377,N_8717);
nor U14998 (N_14998,N_8604,N_6499);
xnor U14999 (N_14999,N_6087,N_5078);
xor U15000 (N_15000,N_13719,N_12558);
and U15001 (N_15001,N_14221,N_14542);
xnor U15002 (N_15002,N_10478,N_14808);
nand U15003 (N_15003,N_12096,N_10231);
nor U15004 (N_15004,N_13607,N_11640);
and U15005 (N_15005,N_14656,N_14637);
and U15006 (N_15006,N_10534,N_11642);
xor U15007 (N_15007,N_13395,N_14075);
or U15008 (N_15008,N_10361,N_10699);
or U15009 (N_15009,N_14074,N_10044);
and U15010 (N_15010,N_14940,N_12434);
or U15011 (N_15011,N_10099,N_13286);
or U15012 (N_15012,N_11403,N_14514);
and U15013 (N_15013,N_14689,N_11304);
xnor U15014 (N_15014,N_11918,N_12553);
xor U15015 (N_15015,N_10449,N_10100);
and U15016 (N_15016,N_13392,N_11977);
nand U15017 (N_15017,N_11035,N_10342);
nor U15018 (N_15018,N_11370,N_10981);
nor U15019 (N_15019,N_10089,N_10520);
or U15020 (N_15020,N_12311,N_10603);
nand U15021 (N_15021,N_11654,N_13554);
xnor U15022 (N_15022,N_10200,N_10193);
nand U15023 (N_15023,N_12134,N_14740);
xnor U15024 (N_15024,N_12640,N_11248);
or U15025 (N_15025,N_14247,N_13322);
or U15026 (N_15026,N_13971,N_12573);
or U15027 (N_15027,N_14550,N_13780);
and U15028 (N_15028,N_10023,N_12926);
nand U15029 (N_15029,N_12199,N_11697);
and U15030 (N_15030,N_13296,N_14695);
or U15031 (N_15031,N_14963,N_12921);
nor U15032 (N_15032,N_13752,N_11633);
xor U15033 (N_15033,N_12923,N_10959);
nor U15034 (N_15034,N_13933,N_14754);
or U15035 (N_15035,N_12473,N_10207);
nor U15036 (N_15036,N_10442,N_11952);
nor U15037 (N_15037,N_13939,N_11657);
xnor U15038 (N_15038,N_12151,N_12601);
nand U15039 (N_15039,N_13037,N_13685);
nor U15040 (N_15040,N_11429,N_11177);
and U15041 (N_15041,N_10000,N_14967);
nor U15042 (N_15042,N_11186,N_13421);
nand U15043 (N_15043,N_13211,N_11155);
and U15044 (N_15044,N_13239,N_14323);
or U15045 (N_15045,N_11891,N_12362);
or U15046 (N_15046,N_10014,N_12121);
nand U15047 (N_15047,N_11306,N_11480);
and U15048 (N_15048,N_11754,N_12300);
nor U15049 (N_15049,N_11361,N_14841);
nand U15050 (N_15050,N_11572,N_13107);
nand U15051 (N_15051,N_10568,N_12585);
xnor U15052 (N_15052,N_10715,N_14017);
xnor U15053 (N_15053,N_12470,N_13809);
or U15054 (N_15054,N_13687,N_13579);
nor U15055 (N_15055,N_12119,N_12825);
nand U15056 (N_15056,N_14164,N_10798);
nand U15057 (N_15057,N_11011,N_13544);
nand U15058 (N_15058,N_11969,N_10587);
and U15059 (N_15059,N_13690,N_14518);
or U15060 (N_15060,N_10060,N_11335);
nand U15061 (N_15061,N_14393,N_13154);
nor U15062 (N_15062,N_11010,N_11620);
nor U15063 (N_15063,N_10188,N_14035);
nor U15064 (N_15064,N_13701,N_14724);
and U15065 (N_15065,N_14556,N_11066);
xor U15066 (N_15066,N_14315,N_11913);
and U15067 (N_15067,N_12847,N_10775);
xnor U15068 (N_15068,N_11415,N_10918);
nor U15069 (N_15069,N_10781,N_12692);
xnor U15070 (N_15070,N_13472,N_14988);
xnor U15071 (N_15071,N_10007,N_11297);
nand U15072 (N_15072,N_12721,N_10021);
or U15073 (N_15073,N_14582,N_14823);
nand U15074 (N_15074,N_13815,N_10818);
xor U15075 (N_15075,N_13217,N_11794);
nand U15076 (N_15076,N_14507,N_13490);
xnor U15077 (N_15077,N_14567,N_11265);
nand U15078 (N_15078,N_13750,N_11027);
or U15079 (N_15079,N_12531,N_14520);
or U15080 (N_15080,N_13161,N_14917);
or U15081 (N_15081,N_11289,N_14326);
xnor U15082 (N_15082,N_12077,N_14054);
nand U15083 (N_15083,N_13077,N_10469);
or U15084 (N_15084,N_13941,N_14274);
nor U15085 (N_15085,N_14147,N_12645);
nor U15086 (N_15086,N_14552,N_14465);
and U15087 (N_15087,N_12145,N_10867);
nand U15088 (N_15088,N_10773,N_13022);
xnor U15089 (N_15089,N_10495,N_11598);
and U15090 (N_15090,N_13728,N_12809);
nand U15091 (N_15091,N_13848,N_13367);
nand U15092 (N_15092,N_13174,N_11185);
or U15093 (N_15093,N_10426,N_11854);
xnor U15094 (N_15094,N_13813,N_10653);
or U15095 (N_15095,N_11139,N_14061);
xnor U15096 (N_15096,N_11823,N_14226);
nor U15097 (N_15097,N_13835,N_11147);
xor U15098 (N_15098,N_10430,N_14802);
or U15099 (N_15099,N_11603,N_10698);
nand U15100 (N_15100,N_12856,N_14821);
nor U15101 (N_15101,N_13073,N_10151);
nor U15102 (N_15102,N_14447,N_14392);
nand U15103 (N_15103,N_13720,N_10514);
nor U15104 (N_15104,N_12070,N_10196);
xnor U15105 (N_15105,N_12292,N_11454);
or U15106 (N_15106,N_11243,N_12678);
and U15107 (N_15107,N_12644,N_12715);
nor U15108 (N_15108,N_13783,N_13309);
nand U15109 (N_15109,N_12051,N_14446);
and U15110 (N_15110,N_13333,N_11498);
nand U15111 (N_15111,N_10459,N_11832);
nor U15112 (N_15112,N_11128,N_14743);
and U15113 (N_15113,N_10085,N_12159);
or U15114 (N_15114,N_12377,N_10289);
xor U15115 (N_15115,N_14885,N_14363);
xor U15116 (N_15116,N_14258,N_13441);
xnor U15117 (N_15117,N_14050,N_12885);
and U15118 (N_15118,N_14261,N_10790);
xnor U15119 (N_15119,N_12332,N_11451);
or U15120 (N_15120,N_14768,N_12616);
and U15121 (N_15121,N_10287,N_10812);
nor U15122 (N_15122,N_10064,N_12412);
and U15123 (N_15123,N_13857,N_14161);
or U15124 (N_15124,N_12891,N_14372);
nand U15125 (N_15125,N_11946,N_12308);
nand U15126 (N_15126,N_10174,N_13257);
and U15127 (N_15127,N_14271,N_14709);
or U15128 (N_15128,N_12592,N_10864);
xor U15129 (N_15129,N_11099,N_10148);
nor U15130 (N_15130,N_11921,N_13341);
and U15131 (N_15131,N_12727,N_13007);
nor U15132 (N_15132,N_14620,N_14111);
xor U15133 (N_15133,N_14858,N_12491);
xor U15134 (N_15134,N_14073,N_12829);
and U15135 (N_15135,N_11092,N_11531);
or U15136 (N_15136,N_14647,N_14364);
nand U15137 (N_15137,N_12965,N_10857);
and U15138 (N_15138,N_12057,N_10283);
nand U15139 (N_15139,N_12111,N_13775);
nor U15140 (N_15140,N_14855,N_12361);
xor U15141 (N_15141,N_11847,N_11455);
xor U15142 (N_15142,N_10397,N_14448);
nand U15143 (N_15143,N_10106,N_10737);
xnor U15144 (N_15144,N_12661,N_12498);
and U15145 (N_15145,N_11637,N_14998);
nor U15146 (N_15146,N_11967,N_12050);
xnor U15147 (N_15147,N_10136,N_14551);
nand U15148 (N_15148,N_12277,N_12078);
or U15149 (N_15149,N_12161,N_14286);
xor U15150 (N_15150,N_10721,N_12665);
nor U15151 (N_15151,N_11367,N_10847);
and U15152 (N_15152,N_13470,N_14635);
nand U15153 (N_15153,N_13893,N_13051);
xor U15154 (N_15154,N_11971,N_14104);
and U15155 (N_15155,N_12203,N_13834);
nand U15156 (N_15156,N_14375,N_14122);
or U15157 (N_15157,N_14527,N_10935);
and U15158 (N_15158,N_14391,N_11477);
xor U15159 (N_15159,N_13888,N_13624);
or U15160 (N_15160,N_11436,N_10871);
xor U15161 (N_15161,N_10876,N_10239);
xor U15162 (N_15162,N_10576,N_14734);
nand U15163 (N_15163,N_12671,N_12194);
nand U15164 (N_15164,N_10635,N_14160);
nand U15165 (N_15165,N_14617,N_13374);
nand U15166 (N_15166,N_14409,N_10719);
or U15167 (N_15167,N_10001,N_14394);
or U15168 (N_15168,N_10938,N_10630);
nand U15169 (N_15169,N_10175,N_12945);
nor U15170 (N_15170,N_14208,N_11703);
or U15171 (N_15171,N_12632,N_12060);
nor U15172 (N_15172,N_10802,N_10811);
nand U15173 (N_15173,N_14360,N_14048);
or U15174 (N_15174,N_10108,N_12480);
nor U15175 (N_15175,N_14726,N_11905);
xnor U15176 (N_15176,N_11793,N_12245);
or U15177 (N_15177,N_11242,N_10685);
nor U15178 (N_15178,N_13859,N_11101);
or U15179 (N_15179,N_14825,N_10796);
xor U15180 (N_15180,N_13638,N_12983);
and U15181 (N_15181,N_12198,N_14771);
xor U15182 (N_15182,N_13203,N_13935);
nand U15183 (N_15183,N_14675,N_10845);
nor U15184 (N_15184,N_13418,N_11281);
nor U15185 (N_15185,N_12544,N_12790);
or U15186 (N_15186,N_11356,N_13986);
nand U15187 (N_15187,N_10149,N_14499);
and U15188 (N_15188,N_12477,N_10625);
xnor U15189 (N_15189,N_11029,N_10232);
and U15190 (N_15190,N_11524,N_13363);
and U15191 (N_15191,N_11881,N_10394);
nor U15192 (N_15192,N_12172,N_13737);
nand U15193 (N_15193,N_10946,N_12022);
nand U15194 (N_15194,N_10580,N_10022);
xnor U15195 (N_15195,N_14806,N_10643);
nor U15196 (N_15196,N_13116,N_13186);
and U15197 (N_15197,N_14452,N_11091);
xor U15198 (N_15198,N_11475,N_10974);
and U15199 (N_15199,N_11715,N_13310);
nand U15200 (N_15200,N_13485,N_11539);
or U15201 (N_15201,N_10199,N_11956);
xor U15202 (N_15202,N_14264,N_12455);
nor U15203 (N_15203,N_12086,N_14099);
nor U15204 (N_15204,N_10450,N_11643);
xor U15205 (N_15205,N_11548,N_10674);
nor U15206 (N_15206,N_12808,N_13486);
nor U15207 (N_15207,N_12869,N_11689);
or U15208 (N_15208,N_12981,N_11233);
xnor U15209 (N_15209,N_12631,N_13634);
xor U15210 (N_15210,N_12520,N_14679);
xnor U15211 (N_15211,N_10105,N_12577);
or U15212 (N_15212,N_10835,N_11677);
nand U15213 (N_15213,N_14445,N_13012);
and U15214 (N_15214,N_12739,N_11473);
and U15215 (N_15215,N_10244,N_12810);
nor U15216 (N_15216,N_12504,N_14662);
nand U15217 (N_15217,N_10889,N_14463);
and U15218 (N_15218,N_13112,N_13901);
xnor U15219 (N_15219,N_11288,N_11486);
and U15220 (N_15220,N_13265,N_14432);
nand U15221 (N_15221,N_11492,N_10906);
nor U15222 (N_15222,N_14300,N_14838);
nor U15223 (N_15223,N_14913,N_10440);
xnor U15224 (N_15224,N_12834,N_11217);
xor U15225 (N_15225,N_10567,N_12201);
and U15226 (N_15226,N_10662,N_11904);
or U15227 (N_15227,N_13021,N_10858);
and U15228 (N_15228,N_14900,N_11109);
or U15229 (N_15229,N_13703,N_11647);
or U15230 (N_15230,N_12454,N_12506);
xor U15231 (N_15231,N_12700,N_12024);
or U15232 (N_15232,N_14131,N_12364);
xnor U15233 (N_15233,N_12509,N_11980);
xnor U15234 (N_15234,N_10343,N_13376);
and U15235 (N_15235,N_11467,N_11716);
nor U15236 (N_15236,N_12688,N_12272);
nor U15237 (N_15237,N_11118,N_11404);
and U15238 (N_15238,N_12797,N_13169);
nor U15239 (N_15239,N_13000,N_10577);
and U15240 (N_15240,N_10051,N_12903);
xnor U15241 (N_15241,N_12030,N_14015);
or U15242 (N_15242,N_11230,N_11330);
nor U15243 (N_15243,N_10664,N_10086);
nand U15244 (N_15244,N_14605,N_11982);
or U15245 (N_15245,N_14985,N_14805);
or U15246 (N_15246,N_10045,N_10985);
nand U15247 (N_15247,N_10899,N_12539);
and U15248 (N_15248,N_12246,N_13276);
and U15249 (N_15249,N_10789,N_10128);
nand U15250 (N_15250,N_12497,N_11063);
nor U15251 (N_15251,N_11141,N_10153);
or U15252 (N_15252,N_10349,N_12262);
nor U15253 (N_15253,N_12327,N_10513);
and U15254 (N_15254,N_10947,N_12551);
nor U15255 (N_15255,N_10205,N_14705);
or U15256 (N_15256,N_12943,N_13229);
xnor U15257 (N_15257,N_14043,N_13015);
and U15258 (N_15258,N_10024,N_14165);
xor U15259 (N_15259,N_14882,N_14046);
nor U15260 (N_15260,N_13659,N_10327);
nand U15261 (N_15261,N_14005,N_11622);
nand U15262 (N_15262,N_14177,N_13457);
nor U15263 (N_15263,N_11266,N_14758);
nand U15264 (N_15264,N_12540,N_13358);
and U15265 (N_15265,N_13724,N_11499);
or U15266 (N_15266,N_14856,N_13832);
and U15267 (N_15267,N_14748,N_13619);
nand U15268 (N_15268,N_10376,N_10941);
and U15269 (N_15269,N_11252,N_10113);
xor U15270 (N_15270,N_13176,N_12113);
or U15271 (N_15271,N_10137,N_11607);
or U15272 (N_15272,N_11318,N_14545);
xor U15273 (N_15273,N_12851,N_11742);
nor U15274 (N_15274,N_14842,N_13066);
or U15275 (N_15275,N_11782,N_14419);
or U15276 (N_15276,N_12791,N_12526);
or U15277 (N_15277,N_12735,N_10581);
or U15278 (N_15278,N_11987,N_12171);
and U15279 (N_15279,N_12398,N_11414);
or U15280 (N_15280,N_11025,N_10543);
or U15281 (N_15281,N_10868,N_14175);
nor U15282 (N_15282,N_11775,N_10438);
or U15283 (N_15283,N_12970,N_14737);
nand U15284 (N_15284,N_11138,N_14906);
xor U15285 (N_15285,N_11746,N_13039);
or U15286 (N_15286,N_11048,N_13975);
and U15287 (N_15287,N_11383,N_10360);
nor U15288 (N_15288,N_13318,N_12521);
or U15289 (N_15289,N_12674,N_12280);
xnor U15290 (N_15290,N_10395,N_12352);
xnor U15291 (N_15291,N_10917,N_14385);
xnor U15292 (N_15292,N_10055,N_11618);
nand U15293 (N_15293,N_13964,N_13702);
nor U15294 (N_15294,N_12679,N_13604);
or U15295 (N_15295,N_12984,N_14715);
or U15296 (N_15296,N_12140,N_14349);
nor U15297 (N_15297,N_12603,N_14510);
nand U15298 (N_15298,N_10339,N_13671);
xnor U15299 (N_15299,N_12156,N_14627);
and U15300 (N_15300,N_14253,N_12732);
or U15301 (N_15301,N_14348,N_14693);
or U15302 (N_15302,N_11639,N_13467);
nand U15303 (N_15303,N_10624,N_14596);
nand U15304 (N_15304,N_13969,N_14473);
nor U15305 (N_15305,N_12693,N_14890);
xor U15306 (N_15306,N_12074,N_13155);
or U15307 (N_15307,N_13498,N_11222);
and U15308 (N_15308,N_12927,N_11857);
xnor U15309 (N_15309,N_12507,N_10413);
and U15310 (N_15310,N_13303,N_11108);
nand U15311 (N_15311,N_14251,N_14555);
xnor U15312 (N_15312,N_11839,N_11024);
xor U15313 (N_15313,N_11296,N_11047);
and U15314 (N_15314,N_11562,N_10731);
nor U15315 (N_15315,N_13869,N_12550);
and U15316 (N_15316,N_11036,N_10486);
or U15317 (N_15317,N_12493,N_12500);
nor U15318 (N_15318,N_12565,N_11442);
nor U15319 (N_15319,N_11419,N_13080);
nand U15320 (N_15320,N_11820,N_11870);
and U15321 (N_15321,N_12196,N_10875);
xnor U15322 (N_15322,N_11725,N_11001);
and U15323 (N_15323,N_10431,N_13111);
and U15324 (N_15324,N_10317,N_13827);
xor U15325 (N_15325,N_12125,N_11632);
nor U15326 (N_15326,N_12605,N_14663);
or U15327 (N_15327,N_11340,N_14664);
nor U15328 (N_15328,N_14149,N_10301);
xnor U15329 (N_15329,N_14714,N_12816);
and U15330 (N_15330,N_14310,N_11378);
or U15331 (N_15331,N_12863,N_13676);
or U15332 (N_15332,N_11979,N_13043);
nand U15333 (N_15333,N_11930,N_12483);
xor U15334 (N_15334,N_12962,N_11223);
nand U15335 (N_15335,N_12376,N_13740);
xor U15336 (N_15336,N_10268,N_10842);
nor U15337 (N_15337,N_12578,N_13016);
nand U15338 (N_15338,N_12282,N_14884);
and U15339 (N_15339,N_10237,N_12994);
and U15340 (N_15340,N_14505,N_10043);
nor U15341 (N_15341,N_13948,N_10226);
and U15342 (N_15342,N_12225,N_10973);
nor U15343 (N_15343,N_14036,N_14873);
nand U15344 (N_15344,N_10248,N_12005);
nand U15345 (N_15345,N_11376,N_14130);
xor U15346 (N_15346,N_12942,N_10228);
xnor U15347 (N_15347,N_14969,N_12518);
xor U15348 (N_15348,N_13650,N_12424);
xor U15349 (N_15349,N_10649,N_13336);
or U15350 (N_15350,N_11788,N_14457);
or U15351 (N_15351,N_11947,N_11317);
xnor U15352 (N_15352,N_10261,N_10822);
and U15353 (N_15353,N_13062,N_13705);
and U15354 (N_15354,N_12484,N_14876);
or U15355 (N_15355,N_10987,N_13573);
or U15356 (N_15356,N_12011,N_14396);
nor U15357 (N_15357,N_10124,N_13072);
and U15358 (N_15358,N_10986,N_13299);
nand U15359 (N_15359,N_14612,N_14281);
and U15360 (N_15360,N_13526,N_12185);
or U15361 (N_15361,N_12288,N_11268);
xor U15362 (N_15362,N_12597,N_12363);
nand U15363 (N_15363,N_13426,N_12010);
xor U15364 (N_15364,N_14321,N_12378);
and U15365 (N_15365,N_11079,N_10502);
and U15366 (N_15366,N_11608,N_11549);
and U15367 (N_15367,N_13584,N_11807);
xor U15368 (N_15368,N_14824,N_12935);
nand U15369 (N_15369,N_10690,N_10995);
nor U15370 (N_15370,N_14216,N_12023);
nand U15371 (N_15371,N_12803,N_13110);
or U15372 (N_15372,N_11624,N_10177);
xnor U15373 (N_15373,N_12705,N_10526);
nor U15374 (N_15374,N_13314,N_12662);
nand U15375 (N_15375,N_10952,N_12479);
nand U15376 (N_15376,N_14205,N_13681);
nor U15377 (N_15377,N_13556,N_14456);
xor U15378 (N_15378,N_14930,N_10275);
nand U15379 (N_15379,N_14710,N_12044);
xor U15380 (N_15380,N_14211,N_14925);
and U15381 (N_15381,N_10211,N_12669);
nor U15382 (N_15382,N_11919,N_13099);
xor U15383 (N_15383,N_11687,N_14318);
or U15384 (N_15384,N_14924,N_10574);
and U15385 (N_15385,N_12838,N_11594);
xnor U15386 (N_15386,N_10245,N_10879);
or U15387 (N_15387,N_11965,N_12155);
nor U15388 (N_15388,N_10640,N_10996);
or U15389 (N_15389,N_13905,N_13629);
and U15390 (N_15390,N_12021,N_10214);
nand U15391 (N_15391,N_12559,N_12069);
or U15392 (N_15392,N_14927,N_11395);
xor U15393 (N_15393,N_10632,N_10542);
or U15394 (N_15394,N_14287,N_14626);
and U15395 (N_15395,N_10537,N_10622);
and U15396 (N_15396,N_10262,N_13583);
or U15397 (N_15397,N_13951,N_12525);
and U15398 (N_15398,N_11257,N_13384);
nor U15399 (N_15399,N_12012,N_10689);
or U15400 (N_15400,N_13818,N_14524);
nor U15401 (N_15401,N_11274,N_11055);
and U15402 (N_15402,N_11371,N_13113);
or U15403 (N_15403,N_12109,N_14333);
nor U15404 (N_15404,N_12654,N_12492);
and U15405 (N_15405,N_14041,N_12120);
xnor U15406 (N_15406,N_14680,N_11738);
or U15407 (N_15407,N_13292,N_14966);
and U15408 (N_15408,N_10766,N_12373);
nor U15409 (N_15409,N_12313,N_11332);
and U15410 (N_15410,N_11529,N_14257);
nor U15411 (N_15411,N_11342,N_12396);
nand U15412 (N_15412,N_10084,N_11999);
and U15413 (N_15413,N_12205,N_14943);
nor U15414 (N_15414,N_10920,N_13478);
or U15415 (N_15415,N_13797,N_12515);
nor U15416 (N_15416,N_14098,N_10681);
nor U15417 (N_15417,N_13782,N_14494);
or U15418 (N_15418,N_13093,N_10712);
and U15419 (N_15419,N_10994,N_13916);
nand U15420 (N_15420,N_12989,N_12514);
nand U15421 (N_15421,N_14214,N_12426);
and U15422 (N_15422,N_12606,N_13708);
nor U15423 (N_15423,N_13123,N_11450);
xnor U15424 (N_15424,N_12355,N_11150);
nor U15425 (N_15425,N_14954,N_14652);
and U15426 (N_15426,N_12763,N_11908);
and U15427 (N_15427,N_11595,N_11723);
and U15428 (N_15428,N_14283,N_10955);
xnor U15429 (N_15429,N_13536,N_13406);
nor U15430 (N_15430,N_14931,N_13483);
or U15431 (N_15431,N_11142,N_13393);
and U15432 (N_15432,N_13897,N_14210);
xor U15433 (N_15433,N_12835,N_12167);
xnor U15434 (N_15434,N_10372,N_10963);
nand U15435 (N_15435,N_12574,N_14334);
xnor U15436 (N_15436,N_11465,N_13098);
xor U15437 (N_15437,N_14889,N_12114);
xor U15438 (N_15438,N_13805,N_10532);
xor U15439 (N_15439,N_14135,N_13448);
and U15440 (N_15440,N_11253,N_13293);
nor U15441 (N_15441,N_10611,N_13562);
and U15442 (N_15442,N_14573,N_13697);
and U15443 (N_15443,N_13953,N_12160);
and U15444 (N_15444,N_14250,N_11320);
xor U15445 (N_15445,N_11666,N_10391);
xor U15446 (N_15446,N_14894,N_12370);
nor U15447 (N_15447,N_11251,N_11924);
and U15448 (N_15448,N_10210,N_14156);
nor U15449 (N_15449,N_14068,N_10516);
nor U15450 (N_15450,N_14475,N_13873);
nor U15451 (N_15451,N_10252,N_14004);
and U15452 (N_15452,N_13236,N_10885);
xor U15453 (N_15453,N_13987,N_11733);
nor U15454 (N_15454,N_10700,N_13182);
xor U15455 (N_15455,N_10894,N_11538);
nor U15456 (N_15456,N_13529,N_12919);
or U15457 (N_15457,N_13183,N_14720);
nor U15458 (N_15458,N_10346,N_14798);
xnor U15459 (N_15459,N_11254,N_12569);
nor U15460 (N_15460,N_12707,N_14862);
nand U15461 (N_15461,N_10213,N_11246);
and U15462 (N_15462,N_11729,N_14614);
or U15463 (N_15463,N_10280,N_14633);
and U15464 (N_15464,N_14389,N_11482);
xnor U15465 (N_15465,N_11043,N_14667);
or U15466 (N_15466,N_10745,N_12457);
or U15467 (N_15467,N_12960,N_11551);
nand U15468 (N_15468,N_14123,N_12859);
or U15469 (N_15469,N_14294,N_14938);
and U15470 (N_15470,N_11479,N_13365);
xor U15471 (N_15471,N_11286,N_10227);
xnor U15472 (N_15472,N_13577,N_10316);
or U15473 (N_15473,N_13716,N_13268);
and U15474 (N_15474,N_13669,N_12048);
nand U15475 (N_15475,N_13789,N_12297);
or U15476 (N_15476,N_10524,N_12058);
nor U15477 (N_15477,N_14342,N_13026);
xnor U15478 (N_15478,N_10236,N_12898);
and U15479 (N_15479,N_10671,N_12886);
and U15480 (N_15480,N_12772,N_11227);
or U15481 (N_15481,N_14417,N_11213);
and U15482 (N_15482,N_12094,N_14140);
xnor U15483 (N_15483,N_10883,N_11509);
nand U15484 (N_15484,N_10950,N_11571);
xor U15485 (N_15485,N_14012,N_14528);
nor U15486 (N_15486,N_13890,N_12754);
xor U15487 (N_15487,N_10890,N_12418);
nand U15488 (N_15488,N_12013,N_13230);
and U15489 (N_15489,N_14229,N_10650);
nor U15490 (N_15490,N_10765,N_13718);
xor U15491 (N_15491,N_11179,N_11062);
nand U15492 (N_15492,N_13534,N_11061);
or U15493 (N_15493,N_13497,N_13514);
and U15494 (N_15494,N_14192,N_13757);
and U15495 (N_15495,N_13076,N_10159);
nor U15496 (N_15496,N_12306,N_14599);
or U15497 (N_15497,N_12449,N_13585);
and U15498 (N_15498,N_12897,N_10102);
or U15499 (N_15499,N_11948,N_13244);
nor U15500 (N_15500,N_13221,N_10993);
or U15501 (N_15501,N_12007,N_13704);
xor U15502 (N_15502,N_14462,N_12931);
nand U15503 (N_15503,N_10535,N_14944);
xnor U15504 (N_15504,N_11617,N_14209);
xor U15505 (N_15505,N_11544,N_12893);
xor U15506 (N_15506,N_10753,N_13680);
nor U15507 (N_15507,N_14727,N_14765);
xnor U15508 (N_15508,N_14412,N_13977);
nand U15509 (N_15509,N_12852,N_13994);
xor U15510 (N_15510,N_10760,N_11435);
nand U15511 (N_15511,N_12743,N_10800);
or U15512 (N_15512,N_14284,N_14430);
nor U15513 (N_15513,N_11559,N_10063);
nand U15514 (N_15514,N_13100,N_12231);
nor U15515 (N_15515,N_12102,N_13427);
or U15516 (N_15516,N_10415,N_13868);
or U15517 (N_15517,N_13555,N_11893);
xnor U15518 (N_15518,N_12649,N_11669);
nand U15519 (N_15519,N_14269,N_12647);
xnor U15520 (N_15520,N_14901,N_10824);
nor U15521 (N_15521,N_11874,N_10460);
nand U15522 (N_15522,N_13260,N_13435);
xor U15523 (N_15523,N_13689,N_11761);
nor U15524 (N_15524,N_12805,N_12414);
nand U15525 (N_15525,N_10109,N_11084);
nand U15526 (N_15526,N_11316,N_10296);
nor U15527 (N_15527,N_14543,N_13606);
or U15528 (N_15528,N_13751,N_10929);
or U15529 (N_15529,N_14782,N_14827);
and U15530 (N_15530,N_12736,N_11074);
and U15531 (N_15531,N_10588,N_10758);
and U15532 (N_15532,N_10667,N_10065);
nand U15533 (N_15533,N_14583,N_13966);
or U15534 (N_15534,N_13068,N_12845);
nor U15535 (N_15535,N_11690,N_10432);
nand U15536 (N_15536,N_10479,N_10597);
nor U15537 (N_15537,N_14467,N_14792);
nor U15538 (N_15538,N_11341,N_12485);
or U15539 (N_15539,N_13989,N_11827);
xor U15540 (N_15540,N_14291,N_11817);
and U15541 (N_15541,N_10954,N_14248);
or U15542 (N_15542,N_13610,N_13988);
nand U15543 (N_15543,N_13445,N_13008);
xor U15544 (N_15544,N_13919,N_14402);
and U15545 (N_15545,N_11845,N_13014);
nand U15546 (N_15546,N_14960,N_12933);
and U15547 (N_15547,N_13499,N_11256);
nand U15548 (N_15548,N_13207,N_11705);
nor U15549 (N_15549,N_14290,N_12435);
xor U15550 (N_15550,N_14387,N_11115);
xnor U15551 (N_15551,N_11925,N_10217);
or U15552 (N_15552,N_12741,N_12738);
and U15553 (N_15553,N_11393,N_11573);
nor U15554 (N_15554,N_12655,N_11495);
or U15555 (N_15555,N_14584,N_11802);
nor U15556 (N_15556,N_13135,N_12093);
nand U15557 (N_15557,N_13044,N_12438);
xnor U15558 (N_15558,N_14153,N_10747);
and U15559 (N_15559,N_12350,N_11162);
xnor U15560 (N_15560,N_11993,N_11636);
xnor U15561 (N_15561,N_12687,N_12046);
xor U15562 (N_15562,N_12193,N_12423);
nand U15563 (N_15563,N_11030,N_12554);
xnor U15564 (N_15564,N_12234,N_13743);
nor U15565 (N_15565,N_13308,N_12142);
nor U15566 (N_15566,N_12811,N_12830);
xnor U15567 (N_15567,N_11887,N_13925);
xnor U15568 (N_15568,N_12165,N_10742);
or U15569 (N_15569,N_10971,N_11379);
nor U15570 (N_15570,N_13428,N_10634);
and U15571 (N_15571,N_13453,N_13460);
and U15572 (N_15572,N_13698,N_11410);
nor U15573 (N_15573,N_10851,N_13343);
and U15574 (N_15574,N_13291,N_10922);
or U15575 (N_15575,N_14224,N_11300);
nor U15576 (N_15576,N_10246,N_14517);
nor U15577 (N_15577,N_11597,N_12080);
and U15578 (N_15578,N_13850,N_13833);
and U15579 (N_15579,N_13920,N_12588);
xnor U15580 (N_15580,N_13807,N_14874);
or U15581 (N_15581,N_12917,N_13668);
and U15582 (N_15582,N_12501,N_11464);
and U15583 (N_15583,N_11671,N_12883);
or U15584 (N_15584,N_14794,N_11773);
nand U15585 (N_15585,N_10648,N_12636);
xor U15586 (N_15586,N_14683,N_12706);
nand U15587 (N_15587,N_11020,N_12330);
xnor U15588 (N_15588,N_14981,N_12928);
nand U15589 (N_15589,N_10945,N_10098);
xor U15590 (N_15590,N_14624,N_11623);
or U15591 (N_15591,N_13147,N_11273);
xnor U15592 (N_15592,N_14469,N_11522);
and U15593 (N_15593,N_14576,N_10221);
and U15594 (N_15594,N_13097,N_13515);
or U15595 (N_15595,N_12978,N_10255);
xor U15596 (N_15596,N_10320,N_14502);
and U15597 (N_15597,N_13501,N_13178);
and U15598 (N_15598,N_14189,N_12663);
xnor U15599 (N_15599,N_13722,N_10723);
and U15600 (N_15600,N_10780,N_10791);
nand U15601 (N_15601,N_14541,N_14811);
nand U15602 (N_15602,N_11570,N_14833);
xnor U15603 (N_15603,N_12420,N_12133);
nor U15604 (N_15604,N_13642,N_13173);
and U15605 (N_15605,N_12686,N_14807);
nor U15606 (N_15606,N_11910,N_14057);
nand U15607 (N_15607,N_14819,N_13349);
xor U15608 (N_15608,N_10797,N_11113);
nand U15609 (N_15609,N_13403,N_10553);
and U15610 (N_15610,N_10999,N_11587);
and U15611 (N_15611,N_13005,N_13576);
xnor U15612 (N_15612,N_13364,N_10152);
xor U15613 (N_15613,N_11542,N_14195);
xnor U15614 (N_15614,N_11724,N_12218);
xor U15615 (N_15615,N_14566,N_11806);
nand U15616 (N_15616,N_14176,N_14026);
xor U15617 (N_15617,N_10825,N_12682);
or U15618 (N_15618,N_13205,N_13620);
or U15619 (N_15619,N_13535,N_10638);
and U15620 (N_15620,N_11172,N_12312);
xnor U15621 (N_15621,N_10919,N_12633);
nand U15622 (N_15622,N_13052,N_14403);
or U15623 (N_15623,N_14852,N_11159);
xnor U15624 (N_15624,N_13799,N_10080);
and U15625 (N_15625,N_10891,N_14201);
nor U15626 (N_15626,N_12673,N_12325);
xnor U15627 (N_15627,N_12996,N_13542);
xnor U15628 (N_15628,N_10185,N_14105);
nor U15629 (N_15629,N_10220,N_10130);
and U15630 (N_15630,N_10846,N_13240);
and U15631 (N_15631,N_12922,N_10202);
nand U15632 (N_15632,N_11900,N_12238);
nand U15633 (N_15633,N_11850,N_10276);
or U15634 (N_15634,N_11884,N_12416);
nor U15635 (N_15635,N_11757,N_13302);
nand U15636 (N_15636,N_10897,N_12918);
or U15637 (N_15637,N_10592,N_13510);
and U15638 (N_15638,N_10484,N_14145);
or U15639 (N_15639,N_13956,N_11518);
and U15640 (N_15640,N_12294,N_10499);
nand U15641 (N_15641,N_10302,N_14526);
nand U15642 (N_15642,N_12773,N_10840);
nor U15643 (N_15643,N_11994,N_13172);
xnor U15644 (N_15644,N_10770,N_14317);
or U15645 (N_15645,N_14092,N_14871);
nor U15646 (N_15646,N_12264,N_10616);
and U15647 (N_15647,N_13375,N_14180);
nor U15648 (N_15648,N_13450,N_14482);
and U15649 (N_15649,N_10498,N_13755);
nor U15650 (N_15650,N_12162,N_14414);
xor U15651 (N_15651,N_12235,N_14243);
nor U15652 (N_15652,N_10071,N_12836);
and U15653 (N_15653,N_11694,N_14909);
and U15654 (N_15654,N_11585,N_10453);
nor U15655 (N_15655,N_12768,N_14312);
and U15656 (N_15656,N_13191,N_13649);
or U15657 (N_15657,N_13042,N_10240);
and U15658 (N_15658,N_13399,N_11886);
xor U15659 (N_15659,N_12146,N_14231);
xor U15660 (N_15660,N_11466,N_11207);
and U15661 (N_15661,N_10076,N_10249);
or U15662 (N_15662,N_13481,N_11611);
xor U15663 (N_15663,N_14435,N_12036);
xor U15664 (N_15664,N_11278,N_13712);
and U15665 (N_15665,N_10269,N_12725);
nand U15666 (N_15666,N_11593,N_10732);
and U15667 (N_15667,N_11546,N_14001);
nor U15668 (N_15668,N_10072,N_12658);
nor U15669 (N_15669,N_14359,N_13731);
nand U15670 (N_15670,N_14066,N_14707);
xor U15671 (N_15671,N_14719,N_10501);
xor U15672 (N_15672,N_14700,N_10122);
or U15673 (N_15673,N_13241,N_13480);
or U15674 (N_15674,N_13158,N_11397);
nor U15675 (N_15675,N_14653,N_13753);
nand U15676 (N_15676,N_14265,N_13684);
and U15677 (N_15677,N_14158,N_14094);
or U15678 (N_15678,N_10852,N_11519);
xor U15679 (N_15679,N_13565,N_11319);
nor U15680 (N_15680,N_10010,N_13761);
and U15681 (N_15681,N_10554,N_13851);
nand U15682 (N_15682,N_13288,N_11602);
or U15683 (N_15683,N_13006,N_13222);
nor U15684 (N_15684,N_12443,N_10808);
nand U15685 (N_15685,N_14593,N_11143);
or U15686 (N_15686,N_12714,N_13770);
nor U15687 (N_15687,N_11433,N_14832);
or U15688 (N_15688,N_10035,N_11350);
and U15689 (N_15689,N_14461,N_11869);
nand U15690 (N_15690,N_11777,N_13086);
nor U15691 (N_15691,N_14923,N_10139);
nand U15692 (N_15692,N_11621,N_11567);
nor U15693 (N_15693,N_13165,N_14492);
or U15694 (N_15694,N_10272,N_10115);
and U15695 (N_15695,N_12190,N_13034);
xor U15696 (N_15696,N_13656,N_11338);
xor U15697 (N_15697,N_12173,N_13463);
nor U15698 (N_15698,N_12634,N_14449);
or U15699 (N_15699,N_13345,N_13134);
or U15700 (N_15700,N_12958,N_10670);
or U15701 (N_15701,N_13844,N_12912);
nor U15702 (N_15702,N_14783,N_13495);
nand U15703 (N_15703,N_10752,N_14571);
or U15704 (N_15704,N_10591,N_11204);
and U15705 (N_15705,N_12524,N_10006);
or U15706 (N_15706,N_13630,N_13330);
nor U15707 (N_15707,N_13575,N_10563);
or U15708 (N_15708,N_10849,N_12907);
xnor U15709 (N_15709,N_10002,N_14301);
nand U15710 (N_15710,N_13710,N_12395);
and U15711 (N_15711,N_13955,N_12757);
nor U15712 (N_15712,N_10464,N_10490);
nand U15713 (N_15713,N_12316,N_14322);
nor U15714 (N_15714,N_10546,N_14139);
nor U15715 (N_15715,N_11943,N_11423);
xor U15716 (N_15716,N_13422,N_10830);
nand U15717 (N_15717,N_12062,N_14163);
or U15718 (N_15718,N_14867,N_11131);
nand U15719 (N_15719,N_13400,N_12459);
xor U15720 (N_15720,N_13496,N_10794);
xor U15721 (N_15721,N_14521,N_12072);
or U15722 (N_15722,N_11135,N_12100);
nor U15723 (N_15723,N_14947,N_11709);
and U15724 (N_15724,N_13787,N_13910);
xor U15725 (N_15725,N_12372,N_13865);
nor U15726 (N_15726,N_14769,N_10475);
nand U15727 (N_15727,N_10077,N_13803);
xor U15728 (N_15728,N_12356,N_12122);
or U15729 (N_15729,N_10146,N_10740);
and U15730 (N_15730,N_11203,N_13778);
nand U15731 (N_15731,N_10677,N_13083);
nor U15732 (N_15732,N_13348,N_11298);
nor U15733 (N_15733,N_13746,N_11954);
nand U15734 (N_15734,N_14386,N_13921);
xnor U15735 (N_15735,N_12227,N_12860);
xor U15736 (N_15736,N_11226,N_11045);
nand U15737 (N_15737,N_13886,N_11774);
nand U15738 (N_15738,N_14304,N_11805);
xnor U15739 (N_15739,N_12930,N_11556);
xnor U15740 (N_15740,N_13880,N_12123);
and U15741 (N_15741,N_11420,N_12948);
nor U15742 (N_15742,N_10458,N_14878);
nand U15743 (N_15743,N_10003,N_10103);
nand U15744 (N_15744,N_11659,N_11660);
nor U15745 (N_15745,N_10882,N_13298);
and U15746 (N_15746,N_13040,N_14897);
nand U15747 (N_15747,N_14877,N_11122);
nor U15748 (N_15748,N_11914,N_13992);
and U15749 (N_15749,N_13171,N_11629);
or U15750 (N_15750,N_13396,N_13891);
and U15751 (N_15751,N_14003,N_12635);
or U15752 (N_15752,N_14117,N_11962);
xor U15753 (N_15753,N_13711,N_12009);
nand U15754 (N_15754,N_10839,N_12762);
nand U15755 (N_15755,N_13249,N_11899);
or U15756 (N_15756,N_13602,N_13070);
or U15757 (N_15757,N_13386,N_12348);
and U15758 (N_15758,N_13861,N_11708);
nand U15759 (N_15759,N_13227,N_11895);
nor U15760 (N_15760,N_14948,N_10522);
nand U15761 (N_15761,N_11153,N_13608);
or U15762 (N_15762,N_11759,N_11126);
or U15763 (N_15763,N_12224,N_10046);
xnor U15764 (N_15764,N_10019,N_10154);
or U15765 (N_15765,N_11440,N_11250);
xnor U15766 (N_15766,N_14970,N_13934);
or U15767 (N_15767,N_13644,N_12379);
xor U15768 (N_15768,N_10834,N_13802);
nor U15769 (N_15769,N_14083,N_10556);
and U15770 (N_15770,N_11344,N_11958);
nor U15771 (N_15771,N_12040,N_12138);
and U15772 (N_15772,N_10527,N_14536);
xnor U15773 (N_15773,N_13029,N_14818);
and U15774 (N_15774,N_12625,N_11547);
nand U15775 (N_15775,N_12314,N_12581);
and U15776 (N_15776,N_11554,N_11828);
nand U15777 (N_15777,N_12268,N_13922);
nor U15778 (N_15778,N_12648,N_11129);
and U15779 (N_15779,N_11182,N_13993);
xnor U15780 (N_15780,N_10013,N_13474);
nor U15781 (N_15781,N_14178,N_11683);
nand U15782 (N_15782,N_13282,N_11301);
and U15783 (N_15783,N_14863,N_14801);
nor U15784 (N_15784,N_10170,N_14779);
and U15785 (N_15785,N_11221,N_11872);
or U15786 (N_15786,N_11124,N_12124);
xor U15787 (N_15787,N_10983,N_13632);
or U15788 (N_15788,N_10138,N_11966);
and U15789 (N_15789,N_14788,N_12095);
and U15790 (N_15790,N_11836,N_11458);
or U15791 (N_15791,N_10988,N_14904);
xor U15792 (N_15792,N_13796,N_12614);
and U15793 (N_15793,N_13137,N_11601);
or U15794 (N_15794,N_14659,N_13101);
or U15795 (N_15795,N_11770,N_10550);
nand U15796 (N_15796,N_11214,N_11331);
nor U15797 (N_15797,N_10201,N_12924);
xnor U15798 (N_15798,N_13709,N_13144);
or U15799 (N_15799,N_14421,N_12502);
or U15800 (N_15800,N_13908,N_14000);
or U15801 (N_15801,N_13381,N_12854);
and U15802 (N_15802,N_14657,N_10887);
nor U15803 (N_15803,N_13870,N_10548);
nand U15804 (N_15804,N_12701,N_11391);
and U15805 (N_15805,N_14275,N_12104);
nor U15806 (N_15806,N_11231,N_11837);
nor U15807 (N_15807,N_10411,N_12932);
or U15808 (N_15808,N_13204,N_14308);
xor U15809 (N_15809,N_14643,N_11533);
xor U15810 (N_15810,N_11497,N_11491);
nand U15811 (N_15811,N_10961,N_10416);
nor U15812 (N_15812,N_11046,N_10730);
or U15813 (N_15813,N_10441,N_14500);
nor U15814 (N_15814,N_12241,N_10295);
or U15815 (N_15815,N_13605,N_11211);
xor U15816 (N_15816,N_13316,N_10477);
nor U15817 (N_15817,N_13202,N_11280);
nand U15818 (N_15818,N_12278,N_14879);
xor U15819 (N_15819,N_12799,N_11493);
xor U15820 (N_15820,N_10485,N_10618);
xor U15821 (N_15821,N_13440,N_13959);
and U15822 (N_15822,N_10436,N_11628);
and U15823 (N_15823,N_10884,N_14080);
nor U15824 (N_15824,N_14581,N_10056);
and U15825 (N_15825,N_13615,N_11719);
and U15826 (N_15826,N_14548,N_14096);
xnor U15827 (N_15827,N_11290,N_11767);
nand U15828 (N_15828,N_10016,N_10823);
and U15829 (N_15829,N_11923,N_12759);
or U15830 (N_15830,N_12385,N_13876);
or U15831 (N_15831,N_10350,N_11950);
nor U15832 (N_15832,N_13667,N_12971);
nor U15833 (N_15833,N_11661,N_11137);
or U15834 (N_15834,N_14618,N_10480);
and U15835 (N_15835,N_14113,N_13357);
and U15836 (N_15836,N_14427,N_14951);
xor U15837 (N_15837,N_12699,N_11205);
xnor U15838 (N_15838,N_12444,N_14644);
nand U15839 (N_15839,N_13617,N_14936);
or U15840 (N_15840,N_14957,N_11144);
and U15841 (N_15841,N_12815,N_13636);
nor U15842 (N_15842,N_11665,N_13200);
xor U15843 (N_15843,N_13092,N_10601);
nand U15844 (N_15844,N_13679,N_11012);
xor U15845 (N_15845,N_11976,N_11032);
or U15846 (N_15846,N_13795,N_13943);
nand U15847 (N_15847,N_12656,N_14891);
nor U15848 (N_15848,N_13009,N_14400);
xor U15849 (N_15849,N_13011,N_12784);
and U15850 (N_15850,N_10860,N_13614);
or U15851 (N_15851,N_11056,N_12242);
nand U15852 (N_15852,N_14685,N_13160);
nand U15853 (N_15853,N_13637,N_10218);
or U15854 (N_15854,N_10399,N_12253);
xnor U15855 (N_15855,N_13972,N_13027);
nand U15856 (N_15856,N_12295,N_11523);
or U15857 (N_15857,N_10126,N_11329);
nor U15858 (N_15858,N_13433,N_11955);
and U15859 (N_15859,N_10405,N_13852);
or U15860 (N_15860,N_14255,N_12323);
or U15861 (N_15861,N_14276,N_10344);
or U15862 (N_15862,N_14553,N_13913);
nor U15863 (N_15863,N_11578,N_14854);
and U15864 (N_15864,N_11680,N_14674);
nand U15865 (N_15865,N_12117,N_13139);
xor U15866 (N_15866,N_11916,N_13819);
xor U15867 (N_15867,N_13640,N_11399);
and U15868 (N_15868,N_14831,N_11555);
nor U15869 (N_15869,N_11553,N_11604);
or U15870 (N_15870,N_10815,N_14346);
and U15871 (N_15871,N_14712,N_12744);
nor U15872 (N_15872,N_13766,N_14225);
or U15873 (N_15873,N_10570,N_14546);
or U15874 (N_15874,N_14628,N_12613);
xor U15875 (N_15875,N_11051,N_13145);
and U15876 (N_15876,N_12680,N_11557);
or U15877 (N_15877,N_11149,N_14977);
and U15878 (N_15878,N_10422,N_14196);
nor U15879 (N_15879,N_10804,N_12406);
or U15880 (N_15880,N_14489,N_10821);
nand U15881 (N_15881,N_11478,N_11763);
nand U15882 (N_15882,N_10762,N_11086);
nand U15883 (N_15883,N_14745,N_11873);
or U15884 (N_15884,N_12003,N_14634);
or U15885 (N_15885,N_13214,N_14212);
xor U15886 (N_15886,N_14064,N_13837);
nor U15887 (N_15887,N_10445,N_12310);
nor U15888 (N_15888,N_12256,N_11789);
xor U15889 (N_15889,N_12849,N_11206);
nor U15890 (N_15890,N_14861,N_10647);
nand U15891 (N_15891,N_11154,N_12118);
xor U15892 (N_15892,N_14508,N_10672);
nand U15893 (N_15893,N_11682,N_11975);
or U15894 (N_15894,N_10163,N_14725);
nand U15895 (N_15895,N_10299,N_14677);
nand U15896 (N_15896,N_12800,N_14179);
xor U15897 (N_15897,N_11405,N_13166);
xor U15898 (N_15898,N_12026,N_13654);
nand U15899 (N_15899,N_14126,N_12445);
or U15900 (N_15900,N_13095,N_13695);
and U15901 (N_15901,N_14641,N_11068);
and U15902 (N_15902,N_12236,N_12775);
nand U15903 (N_15903,N_13305,N_13315);
nand U15904 (N_15904,N_10410,N_12328);
or U15905 (N_15905,N_14812,N_14907);
nor U15906 (N_15906,N_10305,N_10466);
or U15907 (N_15907,N_11398,N_10615);
nor U15908 (N_15908,N_13380,N_13447);
xor U15909 (N_15909,N_12170,N_14137);
and U15910 (N_15910,N_12404,N_13465);
xnor U15911 (N_15911,N_10297,N_12555);
nand U15912 (N_15912,N_10040,N_14757);
nand U15913 (N_15913,N_10768,N_11022);
and U15914 (N_15914,N_10260,N_14747);
xnor U15915 (N_15915,N_10104,N_14155);
and U15916 (N_15916,N_12955,N_11815);
nand U15917 (N_15917,N_13129,N_10409);
xnor U15918 (N_15918,N_14922,N_11859);
and U15919 (N_15919,N_10363,N_11877);
nor U15920 (N_15920,N_11566,N_11581);
nor U15921 (N_15921,N_14384,N_12589);
nand U15922 (N_15922,N_13652,N_11041);
nand U15923 (N_15923,N_11136,N_14813);
and U15924 (N_15924,N_10491,N_12599);
nand U15925 (N_15925,N_12986,N_11152);
or U15926 (N_15926,N_14320,N_10345);
nand U15927 (N_15927,N_11651,N_10759);
xnor U15928 (N_15928,N_14405,N_11922);
nor U15929 (N_15929,N_14613,N_12063);
nor U15930 (N_15930,N_10708,N_10826);
xor U15931 (N_15931,N_12284,N_10724);
xnor U15932 (N_15932,N_12365,N_11228);
nand U15933 (N_15933,N_13225,N_12972);
nor U15934 (N_15934,N_13126,N_12820);
and U15935 (N_15935,N_14522,N_11858);
and U15936 (N_15936,N_10171,N_12557);
xor U15937 (N_15937,N_10258,N_12371);
and U15938 (N_15938,N_10366,N_10037);
or U15939 (N_15939,N_12879,N_13439);
nor U15940 (N_15940,N_13432,N_11474);
or U15941 (N_15941,N_11841,N_10703);
xor U15942 (N_15942,N_12664,N_10582);
xor U15943 (N_15943,N_12819,N_11076);
nand U15944 (N_15944,N_11307,N_11866);
nor U15945 (N_15945,N_10982,N_14611);
nand U15946 (N_15946,N_13075,N_12756);
nand U15947 (N_15947,N_14650,N_10369);
and U15948 (N_15948,N_13409,N_12781);
xnor U15949 (N_15949,N_10629,N_12066);
and U15950 (N_15950,N_14646,N_11078);
and U15951 (N_15951,N_10536,N_14609);
nor U15952 (N_15952,N_10254,N_12433);
and U15953 (N_15953,N_11575,N_11600);
xor U15954 (N_15954,N_13898,N_10434);
xor U15955 (N_15955,N_10127,N_10352);
nand U15956 (N_15956,N_11707,N_12857);
xnor U15957 (N_15957,N_11801,N_14902);
and U15958 (N_15958,N_14241,N_10306);
xnor U15959 (N_15959,N_10850,N_12019);
nand U15960 (N_15960,N_11194,N_10117);
xor U15961 (N_15961,N_11530,N_11333);
nor U15962 (N_15962,N_11550,N_14961);
xor U15963 (N_15963,N_12568,N_10468);
nor U15964 (N_15964,N_11730,N_12976);
nor U15965 (N_15965,N_10530,N_11102);
xnor U15966 (N_15966,N_13522,N_13519);
or U15967 (N_15967,N_11931,N_13088);
and U15968 (N_15968,N_14299,N_12874);
or U15969 (N_15969,N_14239,N_12399);
nor U15970 (N_15970,N_10838,N_11019);
xnor U15971 (N_15971,N_13338,N_14826);
xor U15972 (N_15972,N_10803,N_13121);
and U15973 (N_15973,N_12765,N_10560);
nand U15974 (N_15974,N_13477,N_10027);
nor U15975 (N_15975,N_11785,N_14999);
nand U15976 (N_15976,N_12780,N_13623);
nor U15977 (N_15977,N_14547,N_14383);
nand U15978 (N_15978,N_14442,N_13420);
or U15979 (N_15979,N_11443,N_14512);
nand U15980 (N_15980,N_13826,N_12908);
and U15981 (N_15981,N_14694,N_11996);
or U15982 (N_15982,N_12250,N_11166);
nor U15983 (N_15983,N_13351,N_10523);
and U15984 (N_15984,N_10166,N_13907);
xnor U15985 (N_15985,N_10461,N_11487);
nand U15986 (N_15986,N_13729,N_14351);
or U15987 (N_15987,N_14534,N_13324);
nor U15988 (N_15988,N_10709,N_12582);
nand U15989 (N_15989,N_14762,N_14756);
nand U15990 (N_15990,N_11731,N_12894);
and U15991 (N_15991,N_12934,N_14640);
nand U15992 (N_15992,N_13030,N_12624);
or U15993 (N_15993,N_10328,N_14621);
nand U15994 (N_15994,N_11516,N_14623);
or U15995 (N_15995,N_13456,N_10337);
or U15996 (N_15996,N_10609,N_12702);
or U15997 (N_15997,N_13328,N_11146);
nor U15998 (N_15998,N_11528,N_14682);
nand U15999 (N_15999,N_12818,N_14557);
xnor U16000 (N_16000,N_14173,N_12150);
xnor U16001 (N_16001,N_11123,N_12839);
nand U16002 (N_16002,N_12015,N_13767);
and U16003 (N_16003,N_12950,N_14103);
or U16004 (N_16004,N_14731,N_11098);
or U16005 (N_16005,N_14314,N_11328);
or U16006 (N_16006,N_12823,N_11720);
and U16007 (N_16007,N_13301,N_13114);
nand U16008 (N_16008,N_14666,N_13253);
nand U16009 (N_16009,N_13372,N_12572);
nor U16010 (N_16010,N_12347,N_11501);
and U16011 (N_16011,N_13732,N_10859);
nand U16012 (N_16012,N_14222,N_14759);
nand U16013 (N_16013,N_12027,N_14352);
nor U16014 (N_16014,N_10738,N_10281);
nor U16015 (N_16015,N_10924,N_11125);
or U16016 (N_16016,N_13791,N_10614);
nor U16017 (N_16017,N_10754,N_10332);
nand U16018 (N_16018,N_13354,N_13226);
or U16019 (N_16019,N_12877,N_12054);
xnor U16020 (N_16020,N_12837,N_10079);
and U16021 (N_16021,N_14022,N_10388);
nor U16022 (N_16022,N_11840,N_12166);
nand U16023 (N_16023,N_11711,N_13130);
and U16024 (N_16024,N_10418,N_12450);
and U16025 (N_16025,N_12925,N_11911);
nand U16026 (N_16026,N_12182,N_10605);
nor U16027 (N_16027,N_13290,N_11772);
and U16028 (N_16028,N_11885,N_11013);
nand U16029 (N_16029,N_11229,N_14407);
nor U16030 (N_16030,N_13284,N_12583);
xnor U16031 (N_16031,N_14956,N_14007);
nand U16032 (N_16032,N_11552,N_13997);
and U16033 (N_16033,N_13942,N_11664);
xor U16034 (N_16034,N_11485,N_13691);
xor U16035 (N_16035,N_14579,N_14217);
or U16036 (N_16036,N_12002,N_13373);
nor U16037 (N_16037,N_10158,N_14688);
nor U16038 (N_16038,N_13558,N_10810);
nand U16039 (N_16039,N_14564,N_10286);
nor U16040 (N_16040,N_12999,N_10042);
nor U16041 (N_16041,N_13466,N_11615);
and U16042 (N_16042,N_14678,N_13047);
nand U16043 (N_16043,N_14606,N_11347);
nand U16044 (N_16044,N_12646,N_12252);
nor U16045 (N_16045,N_14102,N_10284);
nand U16046 (N_16046,N_13004,N_10763);
xor U16047 (N_16047,N_14244,N_14051);
nor U16048 (N_16048,N_12591,N_13567);
nand U16049 (N_16049,N_12427,N_13513);
and U16050 (N_16050,N_14121,N_10176);
nand U16051 (N_16051,N_10161,N_11745);
or U16052 (N_16052,N_12143,N_14132);
and U16053 (N_16053,N_12571,N_11853);
or U16054 (N_16054,N_10979,N_14602);
and U16055 (N_16055,N_10285,N_11812);
nand U16056 (N_16056,N_14648,N_10335);
xor U16057 (N_16057,N_11007,N_14138);
or U16058 (N_16058,N_13970,N_13360);
xnor U16059 (N_16059,N_10336,N_10642);
xnor U16060 (N_16060,N_11835,N_10334);
and U16061 (N_16061,N_10722,N_11644);
or U16062 (N_16062,N_12035,N_10748);
nand U16063 (N_16063,N_10820,N_14716);
and U16064 (N_16064,N_13625,N_12299);
or U16065 (N_16065,N_11846,N_12431);
nor U16066 (N_16066,N_10874,N_14112);
and U16067 (N_16067,N_11609,N_14232);
or U16068 (N_16068,N_12411,N_12528);
nor U16069 (N_16069,N_11195,N_14058);
and U16070 (N_16070,N_14056,N_12405);
xor U16071 (N_16071,N_14368,N_12503);
or U16072 (N_16072,N_12778,N_14660);
nor U16073 (N_16073,N_11198,N_11541);
nand U16074 (N_16074,N_11670,N_11704);
xor U16075 (N_16075,N_14767,N_12622);
xnor U16076 (N_16076,N_14506,N_10351);
nor U16077 (N_16077,N_12488,N_13405);
nand U16078 (N_16078,N_10900,N_12032);
nand U16079 (N_16079,N_11355,N_10697);
and U16080 (N_16080,N_10364,N_10545);
nand U16081 (N_16081,N_13258,N_12523);
nor U16082 (N_16082,N_11563,N_13540);
nand U16083 (N_16083,N_12728,N_12968);
nand U16084 (N_16084,N_14169,N_11941);
or U16085 (N_16085,N_14327,N_10243);
xor U16086 (N_16086,N_12108,N_11236);
or U16087 (N_16087,N_12892,N_10510);
and U16088 (N_16088,N_14107,N_13232);
and U16089 (N_16089,N_12549,N_14063);
and U16090 (N_16090,N_13773,N_10187);
nand U16091 (N_16091,N_12349,N_13487);
or U16092 (N_16092,N_11038,N_14357);
nand U16093 (N_16093,N_14658,N_13127);
nor U16094 (N_16094,N_14992,N_14533);
nor U16095 (N_16095,N_14501,N_11635);
nor U16096 (N_16096,N_12563,N_13781);
nor U16097 (N_16097,N_13476,N_10401);
xor U16098 (N_16098,N_10565,N_10092);
nand U16099 (N_16099,N_12627,N_13682);
nor U16100 (N_16100,N_13451,N_11384);
and U16101 (N_16101,N_14330,N_12180);
nand U16102 (N_16102,N_12333,N_14919);
nand U16103 (N_16103,N_13771,N_12233);
nor U16104 (N_16104,N_10507,N_12712);
or U16105 (N_16105,N_11360,N_10143);
nand U16106 (N_16106,N_11520,N_14006);
or U16107 (N_16107,N_13369,N_14468);
or U16108 (N_16108,N_11471,N_11726);
nand U16109 (N_16109,N_11781,N_13281);
and U16110 (N_16110,N_12643,N_12876);
nor U16111 (N_16111,N_11416,N_12821);
or U16112 (N_16112,N_11005,N_12345);
nand U16113 (N_16113,N_13507,N_13839);
or U16114 (N_16114,N_10118,N_14784);
and U16115 (N_16115,N_13482,N_13321);
or U16116 (N_16116,N_11973,N_11107);
nor U16117 (N_16117,N_14515,N_10167);
or U16118 (N_16118,N_13944,N_11508);
or U16119 (N_16119,N_14335,N_14150);
nor U16120 (N_16120,N_14381,N_12824);
or U16121 (N_16121,N_13146,N_10512);
nor U16122 (N_16122,N_13601,N_12342);
xor U16123 (N_16123,N_11284,N_13353);
xnor U16124 (N_16124,N_13312,N_10209);
nor U16125 (N_16125,N_12001,N_12047);
and U16126 (N_16126,N_14629,N_12267);
nor U16127 (N_16127,N_14834,N_11238);
xor U16128 (N_16128,N_10880,N_14272);
and U16129 (N_16129,N_13996,N_13164);
nor U16130 (N_16130,N_10841,N_10482);
nor U16131 (N_16131,N_13242,N_11484);
nor U16132 (N_16132,N_12628,N_11998);
and U16133 (N_16133,N_13087,N_13816);
or U16134 (N_16134,N_11765,N_12338);
nand U16135 (N_16135,N_13909,N_11851);
nor U16136 (N_16136,N_13696,N_10787);
or U16137 (N_16137,N_11762,N_13163);
nor U16138 (N_16138,N_13115,N_10263);
or U16139 (N_16139,N_12899,N_10011);
nor U16140 (N_16140,N_13377,N_11656);
and U16141 (N_16141,N_12512,N_13055);
xnor U16142 (N_16142,N_11995,N_10427);
nor U16143 (N_16143,N_14921,N_13385);
nand U16144 (N_16144,N_14845,N_12988);
xnor U16145 (N_16145,N_11829,N_11259);
or U16146 (N_16146,N_12200,N_13674);
and U16147 (N_16147,N_14458,N_13185);
or U16148 (N_16148,N_13824,N_12749);
nand U16149 (N_16149,N_13587,N_11650);
or U16150 (N_16150,N_10476,N_11894);
and U16151 (N_16151,N_13438,N_12068);
or U16152 (N_16152,N_10462,N_13181);
nor U16153 (N_16153,N_11717,N_12429);
or U16154 (N_16154,N_13666,N_13598);
nand U16155 (N_16155,N_14847,N_11305);
nand U16156 (N_16156,N_11083,N_13231);
nand U16157 (N_16157,N_11121,N_12496);
or U16158 (N_16158,N_14866,N_13715);
and U16159 (N_16159,N_10097,N_13001);
nand U16160 (N_16160,N_12341,N_10916);
xnor U16161 (N_16161,N_10756,N_14124);
nand U16162 (N_16162,N_10050,N_14839);
or U16163 (N_16163,N_12793,N_13105);
nand U16164 (N_16164,N_10144,N_10123);
nand U16165 (N_16165,N_11396,N_13259);
and U16166 (N_16166,N_11425,N_13228);
and U16167 (N_16167,N_13754,N_13902);
nand U16168 (N_16168,N_13626,N_13817);
nor U16169 (N_16169,N_11786,N_14908);
or U16170 (N_16170,N_14128,N_13218);
nor U16171 (N_16171,N_11985,N_11963);
xor U16172 (N_16172,N_13928,N_11935);
or U16173 (N_16173,N_10412,N_12533);
xnor U16174 (N_16174,N_10658,N_12034);
nand U16175 (N_16175,N_13206,N_13103);
nor U16176 (N_16176,N_13836,N_12266);
and U16177 (N_16177,N_14814,N_11018);
nor U16178 (N_16178,N_11831,N_11702);
xor U16179 (N_16179,N_13840,N_12453);
or U16180 (N_16180,N_10687,N_14840);
nand U16181 (N_16181,N_13122,N_10844);
and U16182 (N_16182,N_12340,N_11359);
xnor U16183 (N_16183,N_11838,N_14388);
and U16184 (N_16184,N_10521,N_10259);
nor U16185 (N_16185,N_14994,N_12812);
and U16186 (N_16186,N_13549,N_11303);
xor U16187 (N_16187,N_11933,N_11819);
xor U16188 (N_16188,N_10125,N_10686);
nand U16189 (N_16189,N_13069,N_12868);
nand U16190 (N_16190,N_12959,N_10873);
nor U16191 (N_16191,N_14021,N_10623);
nor U16192 (N_16192,N_13527,N_11119);
nor U16193 (N_16193,N_14649,N_11472);
or U16194 (N_16194,N_13618,N_10180);
or U16195 (N_16195,N_11090,N_13853);
nand U16196 (N_16196,N_13389,N_14437);
or U16197 (N_16197,N_14796,N_12522);
nor U16198 (N_16198,N_13511,N_10373);
xor U16199 (N_16199,N_14892,N_13462);
nand U16200 (N_16200,N_11627,N_11861);
or U16201 (N_16201,N_11470,N_10303);
or U16202 (N_16202,N_14453,N_10381);
or U16203 (N_16203,N_14072,N_10446);
xor U16204 (N_16204,N_12667,N_10833);
nand U16205 (N_16205,N_14116,N_13162);
and U16206 (N_16206,N_12556,N_14843);
nand U16207 (N_16207,N_13882,N_14764);
or U16208 (N_16208,N_12430,N_11844);
nand U16209 (N_16209,N_12938,N_11849);
nand U16210 (N_16210,N_10799,N_13963);
and U16211 (N_16211,N_14692,N_14181);
or U16212 (N_16212,N_11313,N_14496);
nand U16213 (N_16213,N_10910,N_10931);
or U16214 (N_16214,N_13199,N_13762);
nand U16215 (N_16215,N_14410,N_12135);
or U16216 (N_16216,N_10313,N_12228);
nor U16217 (N_16217,N_10741,N_11165);
xor U16218 (N_16218,N_10311,N_13843);
nor U16219 (N_16219,N_12178,N_10696);
nand U16220 (N_16220,N_11343,N_13104);
nand U16221 (N_16221,N_14238,N_13455);
and U16222 (N_16222,N_10212,N_12008);
nor U16223 (N_16223,N_12782,N_11446);
xor U16224 (N_16224,N_10178,N_14270);
or U16225 (N_16225,N_14355,N_12615);
and U16226 (N_16226,N_11323,N_14741);
or U16227 (N_16227,N_14345,N_12296);
nand U16228 (N_16228,N_13653,N_13738);
and U16229 (N_16229,N_11756,N_14371);
and U16230 (N_16230,N_13657,N_10452);
or U16231 (N_16231,N_10607,N_14760);
and U16232 (N_16232,N_11270,N_14776);
or U16233 (N_16233,N_11928,N_12844);
nand U16234 (N_16234,N_13238,N_14971);
and U16235 (N_16235,N_14213,N_13157);
nor U16236 (N_16236,N_10250,N_10222);
and U16237 (N_16237,N_12103,N_14095);
nand U16238 (N_16238,N_13190,N_11006);
and U16239 (N_16239,N_12850,N_10493);
xor U16240 (N_16240,N_14065,N_12476);
xor U16241 (N_16241,N_12608,N_14198);
or U16242 (N_16242,N_12576,N_11276);
nand U16243 (N_16243,N_11039,N_13334);
nand U16244 (N_16244,N_11161,N_11698);
nand U16245 (N_16245,N_14406,N_14895);
nand U16246 (N_16246,N_14763,N_12319);
or U16247 (N_16247,N_13945,N_13023);
and U16248 (N_16248,N_10133,N_13918);
and U16249 (N_16249,N_14549,N_14916);
nor U16250 (N_16250,N_11699,N_12116);
xnor U16251 (N_16251,N_12841,N_10009);
and U16252 (N_16252,N_10968,N_10028);
nand U16253 (N_16253,N_11085,N_13149);
nor U16254 (N_16254,N_12401,N_14120);
nor U16255 (N_16255,N_10074,N_14397);
and U16256 (N_16256,N_10326,N_10854);
and U16257 (N_16257,N_13949,N_12081);
nand U16258 (N_16258,N_11014,N_10353);
and U16259 (N_16259,N_13443,N_13627);
or U16260 (N_16260,N_12997,N_14804);
and U16261 (N_16261,N_13936,N_14718);
and U16262 (N_16262,N_10069,N_11505);
or U16263 (N_16263,N_11052,N_10562);
nand U16264 (N_16264,N_13054,N_14703);
xor U16265 (N_16265,N_13518,N_11282);
nor U16266 (N_16266,N_12320,N_12331);
nand U16267 (N_16267,N_14721,N_13250);
nor U16268 (N_16268,N_14729,N_11937);
or U16269 (N_16269,N_12391,N_14829);
or U16270 (N_16270,N_14109,N_14498);
and U16271 (N_16271,N_13167,N_13063);
and U16272 (N_16272,N_10549,N_10215);
xor U16273 (N_16273,N_10093,N_13270);
nand U16274 (N_16274,N_12905,N_14440);
and U16275 (N_16275,N_14860,N_13235);
or U16276 (N_16276,N_11599,N_11822);
nor U16277 (N_16277,N_13142,N_14869);
and U16278 (N_16278,N_14110,N_11314);
and U16279 (N_16279,N_10367,N_11712);
xor U16280 (N_16280,N_13713,N_14562);
nand U16281 (N_16281,N_13747,N_12675);
nor U16282 (N_16282,N_13790,N_13930);
and U16283 (N_16283,N_10292,N_14670);
nor U16284 (N_16284,N_13973,N_13082);
or U16285 (N_16285,N_14684,N_10406);
and U16286 (N_16286,N_12513,N_10714);
nor U16287 (N_16287,N_13564,N_11890);
nand U16288 (N_16288,N_12575,N_12748);
or U16289 (N_16289,N_13347,N_14933);
and U16290 (N_16290,N_11970,N_10377);
nor U16291 (N_16291,N_11164,N_11490);
nor U16292 (N_16292,N_12357,N_11310);
and U16293 (N_16293,N_13950,N_13210);
nand U16294 (N_16294,N_12566,N_11613);
nand U16295 (N_16295,N_12711,N_11727);
nor U16296 (N_16296,N_11174,N_12065);
nor U16297 (N_16297,N_11220,N_12867);
nor U16298 (N_16298,N_14042,N_10467);
xor U16299 (N_16299,N_13611,N_10005);
nor U16300 (N_16300,N_13894,N_14965);
nand U16301 (N_16301,N_14219,N_11082);
nand U16302 (N_16302,N_11192,N_14292);
nand U16303 (N_16303,N_12004,N_10324);
xnor U16304 (N_16304,N_13279,N_14973);
nor U16305 (N_16305,N_12244,N_12770);
nor U16306 (N_16306,N_10385,N_11734);
nor U16307 (N_16307,N_10251,N_13903);
xnor U16308 (N_16308,N_10934,N_10735);
and U16309 (N_16309,N_12374,N_13237);
and U16310 (N_16310,N_12611,N_10315);
nor U16311 (N_16311,N_12499,N_12274);
and U16312 (N_16312,N_14795,N_12324);
nor U16313 (N_16313,N_13133,N_12360);
nand U16314 (N_16314,N_10483,N_12642);
xor U16315 (N_16315,N_13120,N_10749);
or U16316 (N_16316,N_10788,N_14875);
xor U16317 (N_16317,N_13699,N_13020);
or U16318 (N_16318,N_12064,N_14990);
nand U16319 (N_16319,N_13700,N_10831);
xor U16320 (N_16320,N_14174,N_10355);
and U16321 (N_16321,N_10049,N_11009);
nand U16322 (N_16322,N_11736,N_10116);
nand U16323 (N_16323,N_13484,N_11990);
nor U16324 (N_16324,N_11112,N_14070);
and U16325 (N_16325,N_11710,N_11771);
nor U16326 (N_16326,N_12261,N_11511);
xnor U16327 (N_16327,N_10181,N_12460);
xnor U16328 (N_16328,N_12321,N_13036);
nand U16329 (N_16329,N_11120,N_11021);
or U16330 (N_16330,N_10266,N_10767);
and U16331 (N_16331,N_10600,N_12458);
xnor U16332 (N_16332,N_11427,N_13213);
xnor U16333 (N_16333,N_13946,N_12795);
xnor U16334 (N_16334,N_13317,N_12163);
or U16335 (N_16335,N_10140,N_11500);
xnor U16336 (N_16336,N_11476,N_12018);
or U16337 (N_16337,N_10515,N_11073);
xnor U16338 (N_16338,N_13523,N_11312);
xor U16339 (N_16339,N_10041,N_10359);
nand U16340 (N_16340,N_10162,N_10114);
nand U16341 (N_16341,N_14423,N_14585);
xor U16342 (N_16342,N_14577,N_13820);
or U16343 (N_16343,N_13494,N_11616);
or U16344 (N_16344,N_11513,N_14370);
or U16345 (N_16345,N_10750,N_10318);
nor U16346 (N_16346,N_12911,N_14338);
or U16347 (N_16347,N_12164,N_11067);
xnor U16348 (N_16348,N_11856,N_13085);
and U16349 (N_16349,N_14415,N_14167);
nor U16350 (N_16350,N_10423,N_13248);
xnor U16351 (N_16351,N_11605,N_13361);
nor U16352 (N_16352,N_13401,N_11675);
nor U16353 (N_16353,N_14146,N_13694);
xnor U16354 (N_16354,N_11196,N_10015);
nand U16355 (N_16355,N_10264,N_13064);
nand U16356 (N_16356,N_10081,N_11558);
and U16357 (N_16357,N_10817,N_11903);
xnor U16358 (N_16358,N_13633,N_11889);
or U16359 (N_16359,N_10684,N_10913);
or U16360 (N_16360,N_11017,N_13019);
or U16361 (N_16361,N_14240,N_12570);
nor U16362 (N_16362,N_10646,N_11190);
and U16363 (N_16363,N_13726,N_14915);
and U16364 (N_16364,N_12761,N_11406);
nand U16365 (N_16365,N_14019,N_13459);
xnor U16366 (N_16366,N_10392,N_11826);
and U16367 (N_16367,N_14339,N_12771);
nor U16368 (N_16368,N_14118,N_13061);
xnor U16369 (N_16369,N_10778,N_12548);
nor U16370 (N_16370,N_13561,N_11267);
nor U16371 (N_16371,N_11326,N_10552);
xor U16372 (N_16372,N_14898,N_12866);
nand U16373 (N_16373,N_14511,N_10633);
nor U16374 (N_16374,N_13119,N_13983);
xor U16375 (N_16375,N_10589,N_10183);
nand U16376 (N_16376,N_12315,N_11674);
nor U16377 (N_16377,N_12181,N_13326);
and U16378 (N_16378,N_12567,N_10256);
or U16379 (N_16379,N_12630,N_10312);
nor U16380 (N_16380,N_11200,N_10606);
and U16381 (N_16381,N_12289,N_13168);
nand U16382 (N_16382,N_14436,N_13356);
and U16383 (N_16383,N_13900,N_13096);
nor U16384 (N_16384,N_13962,N_10713);
nor U16385 (N_16385,N_11783,N_11679);
xnor U16386 (N_16386,N_13355,N_10375);
and U16387 (N_16387,N_11299,N_12920);
nand U16388 (N_16388,N_14911,N_13670);
nand U16389 (N_16389,N_14199,N_11089);
nand U16390 (N_16390,N_13736,N_13590);
or U16391 (N_16391,N_13774,N_13430);
xor U16392 (N_16392,N_14100,N_12409);
nand U16393 (N_16393,N_14416,N_10881);
xnor U16394 (N_16394,N_10673,N_13545);
xnor U16395 (N_16395,N_14190,N_12144);
and U16396 (N_16396,N_12760,N_13745);
xnor U16397 (N_16397,N_14033,N_14361);
xnor U16398 (N_16398,N_14144,N_10861);
nor U16399 (N_16399,N_14607,N_12301);
nor U16400 (N_16400,N_12240,N_14989);
and U16401 (N_16401,N_13557,N_10457);
nand U16402 (N_16402,N_14565,N_14976);
xor U16403 (N_16403,N_12469,N_11208);
and U16404 (N_16404,N_14610,N_12098);
or U16405 (N_16405,N_13858,N_11814);
and U16406 (N_16406,N_11163,N_12188);
xor U16407 (N_16407,N_10525,N_12806);
and U16408 (N_16408,N_14793,N_11380);
nor U16409 (N_16409,N_10980,N_13509);
and U16410 (N_16410,N_12186,N_11057);
xnor U16411 (N_16411,N_13371,N_14595);
nand U16412 (N_16412,N_12684,N_14964);
and U16413 (N_16413,N_11855,N_13031);
nor U16414 (N_16414,N_11132,N_13424);
or U16415 (N_16415,N_14002,N_12452);
or U16416 (N_16416,N_11357,N_14702);
nand U16417 (N_16417,N_14324,N_11610);
or U16418 (N_16418,N_11065,N_12676);
nor U16419 (N_16419,N_12481,N_10494);
nor U16420 (N_16420,N_14332,N_13981);
or U16421 (N_16421,N_13603,N_14735);
xor U16422 (N_16422,N_10111,N_11496);
xor U16423 (N_16423,N_10094,N_14013);
xnor U16424 (N_16424,N_11561,N_10886);
nand U16425 (N_16425,N_12833,N_10135);
xnor U16426 (N_16426,N_14929,N_10694);
or U16427 (N_16427,N_10956,N_14481);
or U16428 (N_16428,N_12487,N_10702);
nor U16429 (N_16429,N_11879,N_13967);
nand U16430 (N_16430,N_10927,N_10958);
or U16431 (N_16431,N_11833,N_14151);
xor U16432 (N_16432,N_13153,N_11240);
or U16433 (N_16433,N_11506,N_14235);
nor U16434 (N_16434,N_11945,N_10509);
and U16435 (N_16435,N_12537,N_10271);
xor U16436 (N_16436,N_10975,N_14968);
xor U16437 (N_16437,N_12329,N_12831);
or U16438 (N_16438,N_13337,N_10718);
nor U16439 (N_16439,N_13520,N_11579);
xor U16440 (N_16440,N_14282,N_11521);
xor U16441 (N_16441,N_11592,N_11188);
nand U16442 (N_16442,N_12639,N_10656);
xnor U16443 (N_16443,N_10197,N_10421);
nor U16444 (N_16444,N_11438,N_10783);
or U16445 (N_16445,N_11302,N_11526);
nor U16446 (N_16446,N_12901,N_10017);
xor U16447 (N_16447,N_13194,N_12486);
xor U16448 (N_16448,N_10253,N_11158);
nor U16449 (N_16449,N_12386,N_12407);
nand U16450 (N_16450,N_11087,N_13528);
or U16451 (N_16451,N_11368,N_13914);
xor U16452 (N_16452,N_14045,N_13808);
and U16453 (N_16453,N_10408,N_13533);
xor U16454 (N_16454,N_12217,N_11358);
or U16455 (N_16455,N_14574,N_13862);
or U16456 (N_16456,N_10575,N_14262);
and U16457 (N_16457,N_10047,N_12529);
xor U16458 (N_16458,N_10184,N_12394);
nor U16459 (N_16459,N_11094,N_13366);
or U16460 (N_16460,N_11239,N_14329);
xnor U16461 (N_16461,N_13074,N_14563);
nand U16462 (N_16462,N_10288,N_11077);
or U16463 (N_16463,N_10474,N_14182);
nor U16464 (N_16464,N_12428,N_12107);
or U16465 (N_16465,N_11510,N_13383);
xor U16466 (N_16466,N_13177,N_13278);
xor U16467 (N_16467,N_13842,N_14958);
xnor U16468 (N_16468,N_12729,N_14942);
or U16469 (N_16469,N_10856,N_14509);
xor U16470 (N_16470,N_10704,N_10241);
nor U16471 (N_16471,N_13581,N_14307);
and U16472 (N_16472,N_10270,N_13655);
or U16473 (N_16473,N_11327,N_12904);
nor U16474 (N_16474,N_13313,N_10892);
nor U16475 (N_16475,N_14690,N_11984);
nand U16476 (N_16476,N_11537,N_11407);
or U16477 (N_16477,N_12753,N_14206);
nor U16478 (N_16478,N_12666,N_13404);
nand U16479 (N_16479,N_12255,N_11897);
and U16480 (N_16480,N_10206,N_11365);
or U16481 (N_16481,N_14319,N_13397);
nand U16482 (N_16482,N_11070,N_10273);
or U16483 (N_16483,N_14537,N_11287);
xor U16484 (N_16484,N_13425,N_12612);
nor U16485 (N_16485,N_12650,N_13209);
and U16486 (N_16486,N_13821,N_13906);
nor U16487 (N_16487,N_13464,N_14848);
and U16488 (N_16488,N_10121,N_13414);
and U16489 (N_16489,N_13940,N_13407);
xor U16490 (N_16490,N_13734,N_14297);
xor U16491 (N_16491,N_10338,N_13580);
and U16492 (N_16492,N_14935,N_14987);
and U16493 (N_16493,N_13877,N_11543);
xor U16494 (N_16494,N_13911,N_12963);
or U16495 (N_16495,N_10923,N_10511);
and U16496 (N_16496,N_11974,N_10384);
xnor U16497 (N_16497,N_14280,N_14454);
nand U16498 (N_16498,N_10505,N_13568);
nand U16499 (N_16499,N_11218,N_11294);
or U16500 (N_16500,N_14544,N_14233);
nor U16501 (N_16501,N_11283,N_12530);
or U16502 (N_16502,N_13024,N_11883);
or U16503 (N_16503,N_13505,N_12746);
xnor U16504 (N_16504,N_14249,N_10274);
xor U16505 (N_16505,N_13049,N_13442);
and U16506 (N_16506,N_13524,N_14234);
nand U16507 (N_16507,N_14945,N_14485);
nand U16508 (N_16508,N_13320,N_10805);
and U16509 (N_16509,N_13046,N_11718);
and U16510 (N_16510,N_10307,N_10659);
xnor U16511 (N_16511,N_12375,N_13025);
xor U16512 (N_16512,N_12619,N_13609);
nand U16513 (N_16513,N_12461,N_14742);
xnor U16514 (N_16514,N_14353,N_12990);
xor U16515 (N_16515,N_12287,N_11584);
or U16516 (N_16516,N_11686,N_12691);
nand U16517 (N_16517,N_14390,N_13124);
nor U16518 (N_16518,N_12090,N_10620);
and U16519 (N_16519,N_13976,N_14398);
or U16520 (N_16520,N_13056,N_11502);
nor U16521 (N_16521,N_12388,N_13663);
or U16522 (N_16522,N_14746,N_11311);
and U16523 (N_16523,N_14918,N_13600);
or U16524 (N_16524,N_14439,N_11648);
and U16525 (N_16525,N_10110,N_11663);
xor U16526 (N_16526,N_12979,N_11008);
xnor U16527 (N_16527,N_11049,N_10348);
xnor U16528 (N_16528,N_14252,N_12519);
xnor U16529 (N_16529,N_11972,N_11421);
nand U16530 (N_16530,N_13489,N_14591);
xnor U16531 (N_16531,N_11127,N_13423);
nor U16532 (N_16532,N_11058,N_13643);
xor U16533 (N_16533,N_13065,N_13245);
xor U16534 (N_16534,N_14797,N_14328);
or U16535 (N_16535,N_11915,N_12814);
and U16536 (N_16536,N_11448,N_14816);
xor U16537 (N_16537,N_10096,N_10083);
or U16538 (N_16538,N_10470,N_14401);
or U16539 (N_16539,N_12787,N_11751);
and U16540 (N_16540,N_12752,N_11494);
and U16541 (N_16541,N_10444,N_12626);
nand U16542 (N_16542,N_12099,N_14039);
nor U16543 (N_16543,N_13931,N_10179);
xnor U16544 (N_16544,N_12967,N_12794);
nor U16545 (N_16545,N_12204,N_14404);
nand U16546 (N_16546,N_13675,N_13175);
nand U16547 (N_16547,N_11932,N_13999);
xor U16548 (N_16548,N_10517,N_14487);
xor U16549 (N_16549,N_11706,N_11428);
nand U16550 (N_16550,N_12158,N_14114);
xor U16551 (N_16551,N_12947,N_12448);
nor U16552 (N_16552,N_12861,N_13271);
nor U16553 (N_16553,N_10341,N_11157);
or U16554 (N_16554,N_13416,N_14770);
nor U16555 (N_16555,N_10358,N_12042);
nand U16556 (N_16556,N_13566,N_14223);
nand U16557 (N_16557,N_14020,N_11808);
or U16558 (N_16558,N_10862,N_10029);
xnor U16559 (N_16559,N_14828,N_13398);
and U16560 (N_16560,N_10020,N_12029);
nor U16561 (N_16561,N_13998,N_13990);
nor U16562 (N_16562,N_11821,N_10816);
xor U16563 (N_16563,N_13454,N_14455);
nand U16564 (N_16564,N_13084,N_12964);
xnor U16565 (N_16565,N_13261,N_13304);
nor U16566 (N_16566,N_13179,N_11424);
or U16567 (N_16567,N_11574,N_10637);
or U16568 (N_16568,N_12213,N_10141);
or U16569 (N_16569,N_11830,N_10428);
nand U16570 (N_16570,N_10970,N_14638);
or U16571 (N_16571,N_10048,N_13431);
nand U16572 (N_16572,N_13812,N_14868);
xnor U16573 (N_16573,N_12351,N_10095);
nand U16574 (N_16574,N_13140,N_13570);
and U16575 (N_16575,N_10528,N_14236);
or U16576 (N_16576,N_11722,N_11612);
or U16577 (N_16577,N_11408,N_12593);
xor U16578 (N_16578,N_12489,N_11468);
nand U16579 (N_16579,N_14732,N_11768);
or U16580 (N_16580,N_10293,N_10940);
and U16581 (N_16581,N_12344,N_12546);
or U16582 (N_16582,N_12745,N_10707);
nor U16583 (N_16583,N_11279,N_12105);
nor U16584 (N_16584,N_14263,N_14723);
xor U16585 (N_16585,N_13264,N_10617);
xor U16586 (N_16586,N_13879,N_12187);
xnor U16587 (N_16587,N_13547,N_12718);
nor U16588 (N_16588,N_12381,N_13707);
xor U16589 (N_16589,N_13759,N_10942);
nand U16590 (N_16590,N_14561,N_14038);
nor U16591 (N_16591,N_12392,N_12197);
nor U16592 (N_16592,N_10242,N_10792);
nor U16593 (N_16593,N_12694,N_14676);
nand U16594 (N_16594,N_14932,N_10356);
and U16595 (N_16595,N_13899,N_12410);
nor U16596 (N_16596,N_14431,N_14830);
nand U16597 (N_16597,N_14651,N_10456);
xnor U16598 (N_16598,N_10626,N_12073);
and U16599 (N_16599,N_14295,N_14254);
nor U16600 (N_16600,N_13723,N_12226);
or U16601 (N_16601,N_14744,N_12061);
nor U16602 (N_16602,N_14302,N_12056);
nand U16603 (N_16603,N_10828,N_14495);
or U16604 (N_16604,N_13810,N_11151);
or U16605 (N_16605,N_10836,N_12464);
nand U16606 (N_16606,N_14093,N_14625);
nand U16607 (N_16607,N_10669,N_14975);
nand U16608 (N_16608,N_14787,N_12991);
xor U16609 (N_16609,N_12257,N_12130);
or U16610 (N_16610,N_11692,N_14946);
nor U16611 (N_16611,N_13342,N_11469);
and U16612 (N_16612,N_13078,N_10801);
and U16613 (N_16613,N_12258,N_11418);
nor U16614 (N_16614,N_10654,N_10331);
and U16615 (N_16615,N_12254,N_10583);
xnor U16616 (N_16616,N_10371,N_11324);
nand U16617 (N_16617,N_13541,N_13323);
nand U16618 (N_16618,N_11769,N_14369);
or U16619 (N_16619,N_11388,N_10572);
and U16620 (N_16620,N_10026,N_13307);
or U16621 (N_16621,N_11431,N_13332);
nand U16622 (N_16622,N_11105,N_10529);
nor U16623 (N_16623,N_13493,N_14928);
xor U16624 (N_16624,N_14859,N_10915);
and U16625 (N_16625,N_10949,N_11452);
xor U16626 (N_16626,N_10368,N_10683);
and U16627 (N_16627,N_12685,N_12541);
or U16628 (N_16628,N_11517,N_10279);
xnor U16629 (N_16629,N_12629,N_14354);
and U16630 (N_16630,N_11981,N_11614);
and U16631 (N_16631,N_13768,N_10726);
nand U16632 (N_16632,N_11004,N_10157);
or U16633 (N_16633,N_14108,N_12872);
or U16634 (N_16634,N_13772,N_14750);
nor U16635 (N_16635,N_12888,N_11545);
or U16636 (N_16636,N_12290,N_13800);
and U16637 (N_16637,N_11339,N_12230);
or U16638 (N_16638,N_13503,N_13251);
and U16639 (N_16639,N_11199,N_14950);
and U16640 (N_16640,N_11483,N_10976);
nor U16641 (N_16641,N_14097,N_11936);
xor U16642 (N_16642,N_14673,N_10291);
and U16643 (N_16643,N_11210,N_13058);
nor U16644 (N_16644,N_11912,N_13280);
xor U16645 (N_16645,N_13965,N_10657);
nand U16646 (N_16646,N_11755,N_13937);
or U16647 (N_16647,N_11752,N_11978);
xnor U16648 (N_16648,N_11002,N_14598);
xnor U16649 (N_16649,N_11892,N_12913);
xnor U16650 (N_16650,N_14539,N_11906);
or U16651 (N_16651,N_12532,N_13553);
nand U16652 (N_16652,N_12087,N_11983);
and U16653 (N_16653,N_13212,N_11183);
or U16654 (N_16654,N_10561,N_10407);
nor U16655 (N_16655,N_10652,N_11173);
and U16656 (N_16656,N_13300,N_13159);
nor U16657 (N_16657,N_12082,N_12956);
xor U16658 (N_16658,N_13822,N_13957);
nand U16659 (N_16659,N_10068,N_11753);
xnor U16660 (N_16660,N_12696,N_11586);
nor U16661 (N_16661,N_12609,N_14903);
or U16662 (N_16662,N_11261,N_13591);
and U16663 (N_16663,N_11787,N_11100);
or U16664 (N_16664,N_13329,N_11901);
or U16665 (N_16665,N_14752,N_12998);
nand U16666 (N_16666,N_11292,N_11540);
nor U16667 (N_16667,N_13184,N_14279);
xnor U16668 (N_16668,N_12697,N_14084);
nand U16669 (N_16669,N_11235,N_13436);
and U16670 (N_16670,N_13923,N_14870);
nand U16671 (N_16671,N_10663,N_13382);
xnor U16672 (N_16672,N_13041,N_14422);
nor U16673 (N_16673,N_14085,N_14608);
nand U16674 (N_16674,N_12045,N_10594);
and U16675 (N_16675,N_14325,N_11439);
xnor U16676 (N_16676,N_13141,N_13262);
xor U16677 (N_16677,N_12698,N_13801);
and U16678 (N_16678,N_11232,N_10508);
xor U16679 (N_16679,N_10928,N_10419);
and U16680 (N_16680,N_11362,N_14986);
xor U16681 (N_16681,N_11875,N_11799);
nor U16682 (N_16682,N_13875,N_11175);
nand U16683 (N_16683,N_14127,N_11054);
nand U16684 (N_16684,N_12335,N_11949);
or U16685 (N_16685,N_12237,N_13285);
or U16686 (N_16686,N_13980,N_11034);
xnor U16687 (N_16687,N_12317,N_12059);
nor U16688 (N_16688,N_10277,N_10330);
nand U16689 (N_16689,N_11293,N_12037);
nor U16690 (N_16690,N_12796,N_14630);
or U16691 (N_16691,N_11219,N_14170);
and U16692 (N_16692,N_14978,N_12425);
and U16693 (N_16693,N_11225,N_10504);
nand U16694 (N_16694,N_10544,N_11641);
xnor U16695 (N_16695,N_13926,N_12221);
and U16696 (N_16696,N_10235,N_12862);
or U16697 (N_16697,N_10641,N_12265);
and U16698 (N_16698,N_11181,N_13756);
xor U16699 (N_16699,N_10463,N_10160);
or U16700 (N_16700,N_14078,N_12747);
nor U16701 (N_16701,N_13552,N_10290);
nor U16702 (N_16702,N_11658,N_11693);
or U16703 (N_16703,N_14791,N_11688);
xnor U16704 (N_16704,N_13136,N_11535);
xnor U16705 (N_16705,N_12657,N_12017);
nor U16706 (N_16706,N_12343,N_13672);
and U16707 (N_16707,N_12792,N_13635);
xnor U16708 (N_16708,N_14661,N_12538);
nor U16709 (N_16709,N_12890,N_12954);
nor U16710 (N_16710,N_13335,N_14554);
xnor U16711 (N_16711,N_13198,N_11631);
or U16712 (N_16712,N_11031,N_10692);
xor U16713 (N_16713,N_13924,N_14781);
nor U16714 (N_16714,N_12183,N_14491);
nand U16715 (N_16715,N_14687,N_10720);
and U16716 (N_16716,N_13247,N_14148);
xnor U16717 (N_16717,N_10389,N_10965);
xor U16718 (N_16718,N_14493,N_12049);
nand U16719 (N_16719,N_10564,N_12067);
nor U16720 (N_16720,N_12769,N_12211);
and U16721 (N_16721,N_10112,N_11927);
nor U16722 (N_16722,N_13370,N_13032);
nand U16723 (N_16723,N_10678,N_14237);
and U16724 (N_16724,N_14367,N_13860);
nor U16725 (N_16725,N_14529,N_13002);
and U16726 (N_16726,N_14686,N_10693);
xor U16727 (N_16727,N_13531,N_13749);
nor U16728 (N_16728,N_10613,N_12307);
or U16729 (N_16729,N_13492,N_10433);
or U16730 (N_16730,N_10937,N_10691);
xnor U16731 (N_16731,N_11673,N_12653);
and U16732 (N_16732,N_13612,N_14444);
and U16733 (N_16733,N_12039,N_10129);
and U16734 (N_16734,N_14497,N_11059);
and U16735 (N_16735,N_12767,N_11140);
xor U16736 (N_16736,N_11606,N_14157);
nand U16737 (N_16737,N_12710,N_11040);
xnor U16738 (N_16738,N_12855,N_12939);
xnor U16739 (N_16739,N_13410,N_10538);
and U16740 (N_16740,N_12101,N_12870);
and U16741 (N_16741,N_13543,N_13665);
and U16742 (N_16742,N_14592,N_12951);
nand U16743 (N_16743,N_13208,N_11072);
or U16744 (N_16744,N_10717,N_11386);
and U16745 (N_16745,N_10447,N_14486);
and U16746 (N_16746,N_10012,N_11037);
nor U16747 (N_16747,N_13197,N_10972);
xor U16748 (N_16748,N_13686,N_14880);
or U16749 (N_16749,N_13995,N_11308);
xor U16750 (N_16750,N_13727,N_13359);
xor U16751 (N_16751,N_10030,N_14242);
nand U16752 (N_16752,N_12390,N_12895);
nor U16753 (N_16753,N_13658,N_10506);
or U16754 (N_16754,N_10744,N_14905);
nor U16755 (N_16755,N_11354,N_10777);
nor U16756 (N_16756,N_11209,N_14029);
and U16757 (N_16757,N_12220,N_13327);
nor U16758 (N_16758,N_11655,N_10370);
nand U16759 (N_16759,N_12358,N_11275);
nor U16760 (N_16760,N_14162,N_10612);
or U16761 (N_16761,N_11460,N_12214);
or U16762 (N_16762,N_13094,N_14711);
and U16763 (N_16763,N_12887,N_11168);
xnor U16764 (N_16764,N_14450,N_10984);
xnor U16765 (N_16765,N_14377,N_11026);
or U16766 (N_16766,N_11167,N_14278);
or U16767 (N_16767,N_10120,N_14071);
nor U16768 (N_16768,N_11960,N_11791);
xor U16769 (N_16769,N_14955,N_13411);
or U16770 (N_16770,N_11681,N_10150);
and U16771 (N_16771,N_12880,N_13594);
or U16772 (N_16772,N_11457,N_11959);
or U16773 (N_16773,N_11672,N_14373);
xnor U16774 (N_16774,N_14306,N_11878);
xor U16775 (N_16775,N_10793,N_14159);
xnor U16776 (N_16776,N_13683,N_14464);
or U16777 (N_16777,N_12153,N_14230);
or U16778 (N_16778,N_10425,N_10282);
nor U16779 (N_16779,N_14197,N_12020);
or U16780 (N_16780,N_11645,N_12383);
nand U16781 (N_16781,N_14736,N_11264);
nor U16782 (N_16782,N_10234,N_13871);
nor U16783 (N_16783,N_10936,N_12600);
or U16784 (N_16784,N_13461,N_12339);
nand U16785 (N_16785,N_14088,N_13325);
or U16786 (N_16786,N_10165,N_10455);
nand U16787 (N_16787,N_10198,N_10172);
nand U16788 (N_16788,N_13578,N_12916);
nor U16789 (N_16789,N_14184,N_12232);
nand U16790 (N_16790,N_14778,N_11426);
xnor U16791 (N_16791,N_10964,N_12038);
or U16792 (N_16792,N_14774,N_10991);
and U16793 (N_16793,N_11591,N_11315);
xor U16794 (N_16794,N_14340,N_14730);
nand U16795 (N_16795,N_10374,N_14817);
nand U16796 (N_16796,N_11336,N_13788);
nor U16797 (N_16797,N_12936,N_14119);
nand U16798 (N_16798,N_13854,N_13596);
nand U16799 (N_16799,N_14803,N_10977);
nor U16800 (N_16800,N_11800,N_11422);
or U16801 (N_16801,N_11382,N_11865);
or U16802 (N_16802,N_11411,N_11868);
nor U16803 (N_16803,N_13661,N_11345);
and U16804 (N_16804,N_12536,N_10247);
and U16805 (N_16805,N_14974,N_12695);
nand U16806 (N_16806,N_12251,N_10855);
and U16807 (N_16807,N_13180,N_12914);
nor U16808 (N_16808,N_10319,N_10557);
or U16809 (N_16809,N_12179,N_12961);
nor U16810 (N_16810,N_12641,N_14883);
or U16811 (N_16811,N_12408,N_10400);
or U16812 (N_16812,N_13915,N_12789);
nand U16813 (N_16813,N_14844,N_13413);
nand U16814 (N_16814,N_13769,N_11096);
and U16815 (N_16815,N_10396,N_10819);
xor U16816 (N_16816,N_11534,N_12463);
xnor U16817 (N_16817,N_12053,N_10869);
nand U16818 (N_16818,N_13593,N_12309);
or U16819 (N_16819,N_14030,N_11685);
or U16820 (N_16820,N_12263,N_11961);
nand U16821 (N_16821,N_10059,N_10645);
nor U16822 (N_16822,N_14365,N_10164);
or U16823 (N_16823,N_11696,N_12937);
and U16824 (N_16824,N_13106,N_12875);
nor U16825 (N_16825,N_12304,N_10733);
xor U16826 (N_16826,N_14008,N_10904);
or U16827 (N_16827,N_13741,N_11430);
nor U16828 (N_16828,N_12704,N_11880);
xnor U16829 (N_16829,N_11189,N_13346);
nor U16830 (N_16830,N_12564,N_13823);
and U16831 (N_16831,N_11750,N_14594);
nand U16832 (N_16832,N_13079,N_13419);
nor U16833 (N_16833,N_10727,N_11272);
and U16834 (N_16834,N_12561,N_10559);
or U16835 (N_16835,N_12547,N_13091);
xnor U16836 (N_16836,N_14037,N_11060);
nor U16837 (N_16837,N_11461,N_10223);
nor U16838 (N_16838,N_13798,N_12802);
and U16839 (N_16839,N_14293,N_11249);
nand U16840 (N_16840,N_10155,N_14079);
xor U16841 (N_16841,N_10785,N_10393);
or U16842 (N_16842,N_12243,N_14538);
nand U16843 (N_16843,N_14451,N_13266);
nor U16844 (N_16844,N_12016,N_14337);
nor U16845 (N_16845,N_12467,N_13143);
and U16846 (N_16846,N_12384,N_14273);
and U16847 (N_16847,N_10300,N_10666);
and U16848 (N_16848,N_11489,N_13648);
and U16849 (N_16849,N_13784,N_14597);
or U16850 (N_16850,N_10786,N_11867);
and U16851 (N_16851,N_10267,N_11117);
or U16852 (N_16852,N_11564,N_14172);
or U16853 (N_16853,N_13102,N_10189);
xnor U16854 (N_16854,N_12148,N_13517);
xnor U16855 (N_16855,N_10957,N_10169);
xor U16856 (N_16856,N_13776,N_13792);
or U16857 (N_16857,N_12260,N_10898);
and U16858 (N_16858,N_11713,N_12733);
nand U16859 (N_16859,N_12724,N_14215);
or U16860 (N_16860,N_12368,N_14188);
or U16861 (N_16861,N_10225,N_14984);
or U16862 (N_16862,N_12586,N_12380);
xnor U16863 (N_16863,N_12025,N_14590);
or U16864 (N_16864,N_12222,N_10070);
nand U16865 (N_16865,N_12157,N_12084);
nor U16866 (N_16866,N_14313,N_14952);
nor U16867 (N_16867,N_10437,N_13283);
nand U16868 (N_16868,N_10896,N_14069);
and U16869 (N_16869,N_10191,N_10091);
or U16870 (N_16870,N_13978,N_11095);
xnor U16871 (N_16871,N_10132,N_10481);
or U16872 (N_16872,N_13295,N_11277);
xnor U16873 (N_16873,N_10390,N_11569);
and U16874 (N_16874,N_10989,N_14141);
xor U16875 (N_16875,N_14519,N_13378);
or U16876 (N_16876,N_12878,N_11271);
xnor U16877 (N_16877,N_10067,N_10706);
or U16878 (N_16878,N_13512,N_12511);
nor U16879 (N_16879,N_14418,N_12858);
and U16880 (N_16880,N_10679,N_14277);
or U16881 (N_16881,N_10569,N_11590);
xnor U16882 (N_16882,N_11373,N_13287);
xnor U16883 (N_16883,N_12478,N_11902);
or U16884 (N_16884,N_12354,N_12944);
xnor U16885 (N_16885,N_13272,N_14309);
nand U16886 (N_16886,N_14753,N_12359);
nor U16887 (N_16887,N_12462,N_10866);
and U16888 (N_16888,N_13532,N_11381);
and U16889 (N_16889,N_11412,N_13003);
or U16890 (N_16890,N_13613,N_13765);
xor U16891 (N_16891,N_11876,N_12969);
nand U16892 (N_16892,N_14134,N_10734);
and U16893 (N_16893,N_13866,N_11369);
xor U16894 (N_16894,N_11237,N_11589);
nor U16895 (N_16895,N_11997,N_14851);
nor U16896 (N_16896,N_12421,N_11269);
xnor U16897 (N_16897,N_11258,N_12652);
nand U16898 (N_16898,N_12750,N_13391);
nor U16899 (N_16899,N_12827,N_14023);
nor U16900 (N_16900,N_12598,N_12884);
and U16901 (N_16901,N_11780,N_12089);
nand U16902 (N_16902,N_10147,N_12177);
or U16903 (N_16903,N_13927,N_10602);
or U16904 (N_16904,N_11776,N_10182);
xor U16905 (N_16905,N_12896,N_10298);
xnor U16906 (N_16906,N_12209,N_11816);
and U16907 (N_16907,N_14820,N_10173);
nand U16908 (N_16908,N_13469,N_13018);
and U16909 (N_16909,N_10644,N_10661);
nand U16910 (N_16910,N_10751,N_10619);
and U16911 (N_16911,N_11080,N_14331);
or U16912 (N_16912,N_10082,N_11843);
nor U16913 (N_16913,N_13849,N_12456);
nor U16914 (N_16914,N_10531,N_10710);
nor U16915 (N_16915,N_13415,N_11187);
and U16916 (N_16916,N_11372,N_14031);
nor U16917 (N_16917,N_10186,N_10939);
or U16918 (N_16918,N_12723,N_12681);
and U16919 (N_16919,N_12618,N_13831);
nor U16920 (N_16920,N_12677,N_14645);
nand U16921 (N_16921,N_11825,N_12326);
or U16922 (N_16922,N_11432,N_10608);
nand U16923 (N_16923,N_13263,N_11532);
nor U16924 (N_16924,N_12505,N_13571);
or U16925 (N_16925,N_13616,N_13651);
xnor U16926 (N_16926,N_14459,N_12207);
nand U16927 (N_16927,N_14979,N_14669);
and U16928 (N_16928,N_14154,N_12584);
xnor U16929 (N_16929,N_10604,N_10586);
nand U16930 (N_16930,N_11463,N_10932);
nor U16931 (N_16931,N_10036,N_12822);
nand U16932 (N_16932,N_11626,N_11760);
nand U16933 (N_16933,N_12014,N_10496);
nand U16934 (N_16934,N_12889,N_13132);
or U16935 (N_16935,N_11863,N_14136);
or U16936 (N_16936,N_11728,N_14142);
or U16937 (N_16937,N_10101,N_12417);
and U16938 (N_16938,N_11103,N_13735);
and U16939 (N_16939,N_14053,N_13491);
and U16940 (N_16940,N_13589,N_13297);
and U16941 (N_16941,N_14886,N_13151);
nor U16942 (N_16942,N_13344,N_12281);
or U16943 (N_16943,N_14786,N_11130);
nor U16944 (N_16944,N_10134,N_10230);
xor U16945 (N_16945,N_11988,N_11653);
or U16946 (N_16946,N_11247,N_10925);
or U16947 (N_16947,N_10776,N_13804);
nor U16948 (N_16948,N_12910,N_13764);
or U16949 (N_16949,N_11322,N_12734);
xnor U16950 (N_16950,N_11434,N_12873);
nand U16951 (N_16951,N_10746,N_14558);
nand U16952 (N_16952,N_14568,N_13252);
and U16953 (N_16953,N_10621,N_10930);
xnor U16954 (N_16954,N_14697,N_10417);
nand U16955 (N_16955,N_12987,N_14671);
or U16956 (N_16956,N_10908,N_12709);
nor U16957 (N_16957,N_14972,N_11462);
or U16958 (N_16958,N_11321,N_11784);
nor U16959 (N_16959,N_10933,N_12785);
nor U16960 (N_16960,N_13863,N_11536);
or U16961 (N_16961,N_14356,N_12906);
or U16962 (N_16962,N_10329,N_11758);
or U16963 (N_16963,N_14395,N_12336);
nor U16964 (N_16964,N_13234,N_13128);
nand U16965 (N_16965,N_14115,N_13148);
and U16966 (N_16966,N_14059,N_14780);
and U16967 (N_16967,N_14289,N_11042);
nor U16968 (N_16968,N_10761,N_13479);
nor U16969 (N_16969,N_11735,N_13108);
nand U16970 (N_16970,N_14586,N_10978);
and U16971 (N_16971,N_12291,N_11064);
nand U16972 (N_16972,N_14525,N_12206);
or U16973 (N_16973,N_11234,N_11385);
xor U16974 (N_16974,N_11201,N_10323);
or U16975 (N_16975,N_11691,N_11016);
nand U16976 (N_16976,N_11170,N_13530);
nor U16977 (N_16977,N_12853,N_13721);
nor U16978 (N_16978,N_12607,N_11795);
nand U16979 (N_16979,N_12977,N_12730);
nand U16980 (N_16980,N_10593,N_11938);
and U16981 (N_16981,N_13896,N_14516);
or U16982 (N_16982,N_14490,N_14713);
and U16983 (N_16983,N_12400,N_14631);
or U16984 (N_16984,N_14316,N_10848);
nor U16985 (N_16985,N_12131,N_13748);
xor U16986 (N_16986,N_11695,N_14503);
xor U16987 (N_16987,N_14010,N_13779);
or U16988 (N_16988,N_12840,N_14009);
nand U16989 (N_16989,N_10190,N_10688);
nand U16990 (N_16990,N_12248,N_11583);
or U16991 (N_16991,N_13350,N_13294);
or U16992 (N_16992,N_12842,N_12174);
nor U16993 (N_16993,N_14082,N_10921);
nor U16994 (N_16994,N_10639,N_10901);
xor U16995 (N_16995,N_13961,N_12154);
nand U16996 (N_16996,N_12403,N_11810);
nand U16997 (N_16997,N_13388,N_11244);
or U16998 (N_16998,N_13739,N_11184);
nor U16999 (N_16999,N_12742,N_13985);
nand U17000 (N_17000,N_11560,N_12285);
nor U17001 (N_17001,N_14425,N_10807);
or U17002 (N_17002,N_14246,N_11824);
nand U17003 (N_17003,N_13254,N_11676);
xor U17004 (N_17004,N_14914,N_10471);
xor U17005 (N_17005,N_10784,N_14488);
nor U17006 (N_17006,N_13814,N_11652);
or U17007 (N_17007,N_12269,N_14532);
xor U17008 (N_17008,N_12817,N_12929);
nand U17009 (N_17009,N_12028,N_11514);
xnor U17010 (N_17010,N_10701,N_11818);
nand U17011 (N_17011,N_10208,N_14204);
xor U17012 (N_17012,N_10728,N_14636);
xnor U17013 (N_17013,N_10387,N_10057);
nand U17014 (N_17014,N_10034,N_12191);
and U17015 (N_17015,N_13830,N_10905);
nand U17016 (N_17016,N_13688,N_11334);
and U17017 (N_17017,N_14766,N_10769);
xnor U17018 (N_17018,N_14853,N_11402);
nor U17019 (N_17019,N_14480,N_10309);
nand U17020 (N_17020,N_14777,N_14420);
nor U17021 (N_17021,N_10168,N_13744);
nor U17022 (N_17022,N_10304,N_12672);
xnor U17023 (N_17023,N_14850,N_14995);
nor U17024 (N_17024,N_14809,N_10503);
nor U17025 (N_17025,N_12303,N_11180);
nand U17026 (N_17026,N_11003,N_14622);
nor U17027 (N_17027,N_12293,N_10764);
or U17028 (N_17028,N_14086,N_13267);
nor U17029 (N_17029,N_13929,N_10233);
xnor U17030 (N_17030,N_13446,N_10651);
or U17031 (N_17031,N_11848,N_10806);
and U17032 (N_17032,N_12594,N_10877);
and U17033 (N_17033,N_12189,N_10145);
nor U17034 (N_17034,N_11263,N_11811);
and U17035 (N_17035,N_10454,N_12720);
nor U17036 (N_17036,N_10827,N_13195);
or U17037 (N_17037,N_12129,N_13188);
nand U17038 (N_17038,N_13597,N_10294);
nand U17039 (N_17039,N_14028,N_11986);
xor U17040 (N_17040,N_11747,N_13872);
nor U17041 (N_17041,N_10194,N_14060);
xnor U17042 (N_17042,N_10943,N_11525);
xnor U17043 (N_17043,N_10420,N_14696);
nand U17044 (N_17044,N_13216,N_13563);
nor U17045 (N_17045,N_11804,N_12210);
xnor U17046 (N_17046,N_12239,N_14305);
xor U17047 (N_17047,N_14789,N_13504);
xnor U17048 (N_17048,N_12788,N_14642);
nor U17049 (N_17049,N_11951,N_12900);
xnor U17050 (N_17050,N_14800,N_10705);
or U17051 (N_17051,N_10655,N_13525);
or U17052 (N_17052,N_12777,N_10893);
nand U17053 (N_17053,N_12472,N_14296);
nor U17054 (N_17054,N_10472,N_10872);
nor U17055 (N_17055,N_12085,N_13013);
and U17056 (N_17056,N_13660,N_10004);
xor U17057 (N_17057,N_13150,N_10951);
nand U17058 (N_17058,N_13885,N_12079);
nand U17059 (N_17059,N_10967,N_12941);
nand U17060 (N_17060,N_13500,N_14267);
nand U17061 (N_17061,N_13725,N_13932);
and U17062 (N_17062,N_10636,N_11576);
nand U17063 (N_17063,N_11156,N_13340);
xor U17064 (N_17064,N_12141,N_13582);
or U17065 (N_17065,N_13968,N_14433);
nor U17066 (N_17066,N_10052,N_14091);
nor U17067 (N_17067,N_10018,N_14575);
and U17068 (N_17068,N_13057,N_14202);
xnor U17069 (N_17069,N_13599,N_12137);
and U17070 (N_17070,N_11798,N_14560);
xor U17071 (N_17071,N_13917,N_13954);
and U17072 (N_17072,N_11337,N_14288);
xor U17073 (N_17073,N_10062,N_14535);
nand U17074 (N_17074,N_12415,N_14424);
nand U17075 (N_17075,N_14106,N_14129);
or U17076 (N_17076,N_13539,N_11721);
xor U17077 (N_17077,N_11700,N_10382);
xor U17078 (N_17078,N_11044,N_14785);
or U17079 (N_17079,N_10107,N_14311);
nand U17080 (N_17080,N_12229,N_10403);
xor U17081 (N_17081,N_11015,N_13733);
xnor U17082 (N_17082,N_14380,N_14245);
nand U17083 (N_17083,N_13255,N_14672);
xor U17084 (N_17084,N_12992,N_11625);
xnor U17085 (N_17085,N_11834,N_10066);
or U17086 (N_17086,N_14962,N_12726);
nor U17087 (N_17087,N_11920,N_11898);
and U17088 (N_17088,N_13352,N_12909);
xnor U17089 (N_17089,N_10966,N_10911);
nand U17090 (N_17090,N_11392,N_12843);
and U17091 (N_17091,N_12346,N_10555);
nor U17092 (N_17092,N_10843,N_13960);
and U17093 (N_17093,N_14799,N_14836);
nor U17094 (N_17094,N_12367,N_14587);
or U17095 (N_17095,N_14413,N_10953);
and U17096 (N_17096,N_12740,N_11968);
nand U17097 (N_17097,N_14849,N_12846);
nor U17098 (N_17098,N_10631,N_11864);
or U17099 (N_17099,N_13138,N_10061);
and U17100 (N_17100,N_13592,N_13991);
xor U17101 (N_17101,N_14865,N_12075);
nor U17102 (N_17102,N_12076,N_10675);
nand U17103 (N_17103,N_13828,N_12952);
xor U17104 (N_17104,N_11860,N_14755);
and U17105 (N_17105,N_13895,N_13777);
xnor U17106 (N_17106,N_14220,N_11375);
nor U17107 (N_17107,N_14438,N_14881);
or U17108 (N_17108,N_13559,N_13277);
or U17109 (N_17109,N_13067,N_10757);
xor U17110 (N_17110,N_12276,N_14937);
nand U17111 (N_17111,N_12413,N_11352);
nor U17112 (N_17112,N_14691,N_12974);
nor U17113 (N_17113,N_10414,N_14570);
nand U17114 (N_17114,N_14559,N_12660);
xnor U17115 (N_17115,N_14580,N_10053);
or U17116 (N_17116,N_11000,N_14034);
xnor U17117 (N_17117,N_13109,N_14193);
nand U17118 (N_17118,N_12440,N_11619);
xor U17119 (N_17119,N_14285,N_11888);
nor U17120 (N_17120,N_13289,N_10383);
nand U17121 (N_17121,N_12587,N_10829);
or U17122 (N_17122,N_11577,N_14336);
and U17123 (N_17123,N_11255,N_12219);
or U17124 (N_17124,N_11939,N_13786);
or U17125 (N_17125,N_14588,N_12620);
or U17126 (N_17126,N_11743,N_13958);
nand U17127 (N_17127,N_14953,N_13841);
nor U17128 (N_17128,N_14888,N_10566);
nand U17129 (N_17129,N_12737,N_14569);
xor U17130 (N_17130,N_12279,N_11363);
nand U17131 (N_17131,N_14531,N_11409);
nor U17132 (N_17132,N_12055,N_11133);
nor U17133 (N_17133,N_11374,N_10357);
nor U17134 (N_17134,N_14478,N_11202);
and U17135 (N_17135,N_12397,N_13417);
xnor U17136 (N_17136,N_10492,N_11749);
and U17137 (N_17137,N_13368,N_14014);
and U17138 (N_17138,N_11349,N_12508);
or U17139 (N_17139,N_12215,N_11353);
xor U17140 (N_17140,N_12447,N_14483);
xnor U17141 (N_17141,N_13048,N_13362);
xor U17142 (N_17142,N_12275,N_12689);
and U17143 (N_17143,N_10216,N_12353);
and U17144 (N_17144,N_13794,N_12975);
nand U17145 (N_17145,N_12801,N_14822);
nor U17146 (N_17146,N_12579,N_11871);
xnor U17147 (N_17147,N_13233,N_14443);
or U17148 (N_17148,N_10039,N_11842);
nor U17149 (N_17149,N_10224,N_14751);
nand U17150 (N_17150,N_12527,N_13730);
nand U17151 (N_17151,N_10914,N_10895);
xnor U17152 (N_17152,N_14991,N_14087);
nand U17153 (N_17153,N_14358,N_10627);
nor U17154 (N_17154,N_10310,N_12184);
nor U17155 (N_17155,N_12755,N_11580);
nand U17156 (N_17156,N_13811,N_14733);
nand U17157 (N_17157,N_14708,N_12305);
nand U17158 (N_17158,N_10579,N_14081);
xor U17159 (N_17159,N_12006,N_13059);
or U17160 (N_17160,N_12764,N_12881);
nor U17161 (N_17161,N_11193,N_12774);
nand U17162 (N_17162,N_12271,N_10878);
or U17163 (N_17163,N_12092,N_14665);
xor U17164 (N_17164,N_13475,N_11779);
nand U17165 (N_17165,N_14654,N_11028);
nor U17166 (N_17166,N_10195,N_10755);
and U17167 (N_17167,N_11481,N_13516);
or U17168 (N_17168,N_11766,N_13884);
and U17169 (N_17169,N_11940,N_11744);
or U17170 (N_17170,N_13586,N_10398);
or U17171 (N_17171,N_12946,N_14399);
nor U17172 (N_17172,N_13979,N_12915);
nor U17173 (N_17173,N_14983,N_13806);
and U17174 (N_17174,N_13887,N_12543);
xnor U17175 (N_17175,N_12731,N_13678);
and U17176 (N_17176,N_10926,N_10676);
or U17177 (N_17177,N_13117,N_12798);
nor U17178 (N_17178,N_11929,N_11714);
or U17179 (N_17179,N_11216,N_14343);
and U17180 (N_17180,N_12202,N_10404);
xor U17181 (N_17181,N_13220,N_14434);
or U17182 (N_17182,N_14018,N_11917);
nand U17183 (N_17183,N_11023,N_12132);
nor U17184 (N_17184,N_14668,N_11667);
nor U17185 (N_17185,N_10088,N_10465);
or U17186 (N_17186,N_10573,N_13693);
nand U17187 (N_17187,N_13473,N_10865);
xor U17188 (N_17188,N_13548,N_11106);
and U17189 (N_17189,N_14699,N_10340);
nor U17190 (N_17190,N_11588,N_12610);
xor U17191 (N_17191,N_11178,N_13125);
nor U17192 (N_17192,N_13402,N_14168);
nor U17193 (N_17193,N_14476,N_14171);
nor U17194 (N_17194,N_14604,N_11053);
and U17195 (N_17195,N_12259,N_11145);
nor U17196 (N_17196,N_14477,N_14016);
and U17197 (N_17197,N_12865,N_14260);
nand U17198 (N_17198,N_12091,N_14362);
nand U17199 (N_17199,N_12334,N_11992);
nor U17200 (N_17200,N_13033,N_12249);
and U17201 (N_17201,N_14810,N_11449);
nor U17202 (N_17202,N_12471,N_10333);
and U17203 (N_17203,N_14268,N_14738);
and U17204 (N_17204,N_14772,N_11507);
nor U17205 (N_17205,N_12494,N_10774);
or U17206 (N_17206,N_10325,N_12031);
and U17207 (N_17207,N_13560,N_10729);
nand U17208 (N_17208,N_10365,N_11684);
xnor U17209 (N_17209,N_10038,N_14655);
xor U17210 (N_17210,N_12302,N_11171);
nor U17211 (N_17211,N_14207,N_10540);
xnor U17212 (N_17212,N_12779,N_14047);
or U17213 (N_17213,N_10660,N_14032);
xor U17214 (N_17214,N_11377,N_13646);
nor U17215 (N_17215,N_12446,N_11445);
and U17216 (N_17216,N_14027,N_14055);
and U17217 (N_17217,N_12097,N_12465);
and U17218 (N_17218,N_10278,N_14775);
or U17219 (N_17219,N_14203,N_12590);
and U17220 (N_17220,N_14835,N_12716);
or U17221 (N_17221,N_11245,N_13269);
or U17222 (N_17222,N_12813,N_10429);
xnor U17223 (N_17223,N_10992,N_12283);
nand U17224 (N_17224,N_10711,N_10451);
nor U17225 (N_17225,N_14739,N_10488);
and U17226 (N_17226,N_10489,N_13053);
or U17227 (N_17227,N_13829,N_13639);
nand U17228 (N_17228,N_12517,N_11678);
nand U17229 (N_17229,N_12112,N_12602);
xnor U17230 (N_17230,N_12719,N_13974);
nor U17231 (N_17231,N_12683,N_13550);
nor U17232 (N_17232,N_12973,N_14441);
nand U17233 (N_17233,N_13595,N_11909);
and U17234 (N_17234,N_11325,N_12940);
nor U17235 (N_17235,N_14540,N_12369);
nand U17236 (N_17236,N_12298,N_11944);
xnor U17237 (N_17237,N_11515,N_14049);
and U17238 (N_17238,N_11527,N_11459);
xor U17239 (N_17239,N_14589,N_14912);
and U17240 (N_17240,N_12776,N_11110);
nand U17241 (N_17241,N_10743,N_13256);
nor U17242 (N_17242,N_10853,N_10813);
nand U17243 (N_17243,N_14980,N_10909);
or U17244 (N_17244,N_11215,N_13437);
nor U17245 (N_17245,N_12442,N_12273);
or U17246 (N_17246,N_12175,N_12659);
xor U17247 (N_17247,N_11813,N_13793);
or U17248 (N_17248,N_13273,N_12286);
and U17249 (N_17249,N_13673,N_12864);
or U17250 (N_17250,N_11262,N_10599);
nor U17251 (N_17251,N_12466,N_13538);
xor U17252 (N_17252,N_10238,N_12617);
nand U17253 (N_17253,N_11803,N_11792);
nor U17254 (N_17254,N_13038,N_13458);
and U17255 (N_17255,N_13224,N_13938);
and U17256 (N_17256,N_10628,N_12106);
xor U17257 (N_17257,N_13984,N_10595);
and U17258 (N_17258,N_12534,N_14504);
xnor U17259 (N_17259,N_11764,N_10551);
or U17260 (N_17260,N_13664,N_13838);
and U17261 (N_17261,N_13187,N_13412);
nor U17262 (N_17262,N_10585,N_13760);
nor U17263 (N_17263,N_14040,N_14303);
and U17264 (N_17264,N_12828,N_13551);
nand U17265 (N_17265,N_10025,N_12621);
nand U17266 (N_17266,N_10119,N_11134);
xnor U17267 (N_17267,N_12651,N_13215);
nor U17268 (N_17268,N_10347,N_10590);
nor U17269 (N_17269,N_13856,N_13785);
and U17270 (N_17270,N_12382,N_13645);
or U17271 (N_17271,N_13677,N_10944);
nor U17272 (N_17272,N_10912,N_13621);
nand U17273 (N_17273,N_13028,N_12490);
nand U17274 (N_17274,N_13246,N_12422);
xor U17275 (N_17275,N_14218,N_10962);
nor U17276 (N_17276,N_12208,N_13379);
or U17277 (N_17277,N_14949,N_11224);
or U17278 (N_17278,N_10725,N_14379);
nand U17279 (N_17279,N_10008,N_13647);
and U17280 (N_17280,N_11896,N_10903);
nor U17281 (N_17281,N_14749,N_11662);
nor U17282 (N_17282,N_14615,N_10519);
or U17283 (N_17283,N_10439,N_14426);
nand U17284 (N_17284,N_10782,N_10424);
or U17285 (N_17285,N_11088,N_12195);
and U17286 (N_17286,N_14101,N_12783);
or U17287 (N_17287,N_12848,N_13471);
nand U17288 (N_17288,N_11991,N_14378);
nor U17289 (N_17289,N_10682,N_13889);
or U17290 (N_17290,N_12168,N_13170);
and U17291 (N_17291,N_10203,N_10907);
nand U17292 (N_17292,N_13193,N_11852);
xnor U17293 (N_17293,N_14366,N_13845);
and U17294 (N_17294,N_11741,N_13982);
nor U17295 (N_17295,N_11862,N_10308);
nor U17296 (N_17296,N_13878,N_10219);
nand U17297 (N_17297,N_14616,N_11097);
xor U17298 (N_17298,N_13081,N_11114);
xor U17299 (N_17299,N_11568,N_11447);
or U17300 (N_17300,N_10990,N_12562);
nand U17301 (N_17301,N_14460,N_13569);
xnor U17302 (N_17302,N_12439,N_11739);
nor U17303 (N_17303,N_12495,N_14704);
xnor U17304 (N_17304,N_14228,N_12147);
or U17305 (N_17305,N_13864,N_10500);
nand U17306 (N_17306,N_14185,N_11456);
and U17307 (N_17307,N_14076,N_14959);
and U17308 (N_17308,N_10779,N_10487);
xnor U17309 (N_17309,N_10795,N_14639);
and U17310 (N_17310,N_14133,N_10058);
or U17311 (N_17311,N_10443,N_13429);
xnor U17312 (N_17312,N_14411,N_10558);
nor U17313 (N_17313,N_14846,N_10736);
xnor U17314 (N_17314,N_14837,N_10497);
xor U17315 (N_17315,N_13196,N_14997);
nor U17316 (N_17316,N_12985,N_13883);
or U17317 (N_17317,N_12708,N_14166);
xnor U17318 (N_17318,N_14408,N_13488);
xnor U17319 (N_17319,N_10032,N_13390);
xnor U17320 (N_17320,N_12713,N_11778);
and U17321 (N_17321,N_14717,N_10668);
nand U17322 (N_17322,N_12216,N_11646);
or U17323 (N_17323,N_14089,N_10863);
nor U17324 (N_17324,N_10997,N_10739);
nand U17325 (N_17325,N_13090,N_14934);
or U17326 (N_17326,N_10998,N_11050);
nand U17327 (N_17327,N_12083,N_14466);
nand U17328 (N_17328,N_11212,N_12468);
or U17329 (N_17329,N_12668,N_14887);
xnor U17330 (N_17330,N_10680,N_14600);
or U17331 (N_17331,N_13010,N_14429);
or U17332 (N_17332,N_14920,N_14471);
xor U17333 (N_17333,N_12152,N_12595);
and U17334 (N_17334,N_11348,N_13912);
and U17335 (N_17335,N_14011,N_12751);
and U17336 (N_17336,N_12957,N_12804);
or U17337 (N_17337,N_14893,N_14062);
xnor U17338 (N_17338,N_12516,N_13118);
nand U17339 (N_17339,N_14864,N_12758);
nand U17340 (N_17340,N_11241,N_13331);
or U17341 (N_17341,N_12128,N_10435);
nand U17342 (N_17342,N_11116,N_12580);
and U17343 (N_17343,N_12033,N_12088);
and U17344 (N_17344,N_10090,N_14350);
nor U17345 (N_17345,N_12722,N_14474);
or U17346 (N_17346,N_10518,N_10578);
nor U17347 (N_17347,N_13311,N_11797);
nor U17348 (N_17348,N_14632,N_13017);
xor U17349 (N_17349,N_11285,N_11033);
xor U17350 (N_17350,N_13628,N_14896);
nor U17351 (N_17351,N_12387,N_14790);
nand U17352 (N_17352,N_11488,N_11503);
and U17353 (N_17353,N_12322,N_10716);
xnor U17354 (N_17354,N_10265,N_12176);
xnor U17355 (N_17355,N_10533,N_12596);
xnor U17356 (N_17356,N_12115,N_14484);
and U17357 (N_17357,N_12882,N_13521);
nor U17358 (N_17358,N_12535,N_13223);
nor U17359 (N_17359,N_13131,N_10541);
xor U17360 (N_17360,N_11071,N_14428);
xor U17361 (N_17361,N_13071,N_14187);
and U17362 (N_17362,N_13408,N_11596);
nand U17363 (N_17363,N_11093,N_13546);
and U17364 (N_17364,N_14186,N_10314);
or U17365 (N_17365,N_12169,N_11176);
and U17366 (N_17366,N_13089,N_12604);
nand U17367 (N_17367,N_11453,N_12389);
nor U17368 (N_17368,N_10902,N_13434);
or U17369 (N_17369,N_14025,N_12270);
and U17370 (N_17370,N_14200,N_13572);
nor U17371 (N_17371,N_10033,N_12482);
and U17372 (N_17372,N_12475,N_12393);
and U17373 (N_17373,N_13156,N_14572);
xor U17374 (N_17374,N_10772,N_14259);
nor U17375 (N_17375,N_11882,N_12402);
xor U17376 (N_17376,N_13742,N_11400);
and U17377 (N_17377,N_14815,N_11934);
or U17378 (N_17378,N_14706,N_11441);
nor U17379 (N_17379,N_10809,N_13274);
xnor U17380 (N_17380,N_13306,N_10054);
nand U17381 (N_17381,N_10087,N_13189);
nand U17382 (N_17382,N_13588,N_10354);
or U17383 (N_17383,N_14872,N_12043);
and U17384 (N_17384,N_13275,N_12637);
and U17385 (N_17385,N_10142,N_12542);
xnor U17386 (N_17386,N_13537,N_14194);
or U17387 (N_17387,N_10448,N_10380);
nand U17388 (N_17388,N_14344,N_14298);
xor U17389 (N_17389,N_11351,N_12993);
and U17390 (N_17390,N_12437,N_14530);
or U17391 (N_17391,N_10969,N_12136);
nand U17392 (N_17392,N_13394,N_13692);
or U17393 (N_17393,N_12638,N_12432);
nand U17394 (N_17394,N_11394,N_10322);
or U17395 (N_17395,N_13502,N_10610);
nor U17396 (N_17396,N_12451,N_12126);
nand U17397 (N_17397,N_11504,N_10031);
xnor U17398 (N_17398,N_10078,N_14926);
nor U17399 (N_17399,N_13706,N_13631);
and U17400 (N_17400,N_12552,N_11069);
xor U17401 (N_17401,N_14857,N_14183);
and U17402 (N_17402,N_14479,N_10257);
nand U17403 (N_17403,N_12000,N_14143);
nand U17404 (N_17404,N_10870,N_14256);
and U17405 (N_17405,N_10837,N_13339);
and U17406 (N_17406,N_14701,N_14044);
nor U17407 (N_17407,N_10362,N_12766);
xor U17408 (N_17408,N_10814,N_13641);
or U17409 (N_17409,N_12545,N_13035);
or U17410 (N_17410,N_14681,N_11169);
nor U17411 (N_17411,N_11197,N_14698);
xnor U17412 (N_17412,N_12419,N_14266);
nand U17413 (N_17413,N_14941,N_10402);
xnor U17414 (N_17414,N_13508,N_14761);
nor U17415 (N_17415,N_10571,N_13050);
nor U17416 (N_17416,N_11191,N_13855);
or U17417 (N_17417,N_12052,N_12807);
and U17418 (N_17418,N_14603,N_12982);
xnor U17419 (N_17419,N_11565,N_13243);
or U17420 (N_17420,N_11701,N_14470);
nand U17421 (N_17421,N_10131,N_11737);
and U17422 (N_17422,N_12623,N_11081);
or U17423 (N_17423,N_11346,N_10832);
or U17424 (N_17424,N_14982,N_12212);
xor U17425 (N_17425,N_11389,N_13867);
and U17426 (N_17426,N_12966,N_11989);
nor U17427 (N_17427,N_13904,N_14619);
or U17428 (N_17428,N_11732,N_13045);
nor U17429 (N_17429,N_13192,N_14067);
nor U17430 (N_17430,N_13825,N_14899);
or U17431 (N_17431,N_14728,N_10192);
xor U17432 (N_17432,N_11907,N_10204);
xor U17433 (N_17433,N_11634,N_14382);
and U17434 (N_17434,N_10771,N_14347);
nor U17435 (N_17435,N_14578,N_11957);
xor U17436 (N_17436,N_11953,N_14993);
nand U17437 (N_17437,N_14341,N_11309);
or U17438 (N_17438,N_12110,N_13717);
or U17439 (N_17439,N_11582,N_13846);
or U17440 (N_17440,N_13892,N_12670);
nand U17441 (N_17441,N_14227,N_12366);
nor U17442 (N_17442,N_12139,N_11512);
nand U17443 (N_17443,N_14773,N_14996);
xnor U17444 (N_17444,N_12826,N_11926);
or U17445 (N_17445,N_13319,N_13758);
nor U17446 (N_17446,N_10378,N_14376);
or U17447 (N_17447,N_10539,N_13452);
nor U17448 (N_17448,N_10073,N_12871);
or U17449 (N_17449,N_11075,N_14152);
nor U17450 (N_17450,N_13201,N_13881);
nor U17451 (N_17451,N_14722,N_14513);
or U17452 (N_17452,N_13763,N_12980);
or U17453 (N_17453,N_12949,N_12223);
nand U17454 (N_17454,N_14472,N_12474);
nand U17455 (N_17455,N_14077,N_13152);
nor U17456 (N_17456,N_10229,N_11649);
and U17457 (N_17457,N_12441,N_11366);
and U17458 (N_17458,N_11437,N_13714);
and U17459 (N_17459,N_14601,N_10948);
or U17460 (N_17460,N_13449,N_11387);
and U17461 (N_17461,N_11748,N_13574);
or U17462 (N_17462,N_14090,N_12902);
and U17463 (N_17463,N_11638,N_14191);
nor U17464 (N_17464,N_12703,N_10584);
nor U17465 (N_17465,N_13444,N_13219);
xor U17466 (N_17466,N_12995,N_11668);
and U17467 (N_17467,N_11390,N_13506);
nor U17468 (N_17468,N_12690,N_14910);
xnor U17469 (N_17469,N_11444,N_13847);
or U17470 (N_17470,N_13874,N_11160);
xnor U17471 (N_17471,N_10379,N_11417);
or U17472 (N_17472,N_12149,N_11364);
or U17473 (N_17473,N_12192,N_13468);
nor U17474 (N_17474,N_11630,N_13947);
or U17475 (N_17475,N_11942,N_10695);
and U17476 (N_17476,N_14374,N_11964);
or U17477 (N_17477,N_12560,N_14052);
nand U17478 (N_17478,N_12510,N_10075);
xnor U17479 (N_17479,N_11401,N_10547);
xor U17480 (N_17480,N_12436,N_13060);
or U17481 (N_17481,N_13952,N_12127);
and U17482 (N_17482,N_10665,N_12953);
or U17483 (N_17483,N_11104,N_12318);
nand U17484 (N_17484,N_10473,N_11260);
and U17485 (N_17485,N_11809,N_14024);
or U17486 (N_17486,N_11111,N_13622);
xor U17487 (N_17487,N_11295,N_10598);
or U17488 (N_17488,N_14523,N_10386);
nor U17489 (N_17489,N_13662,N_11291);
xor U17490 (N_17490,N_14125,N_12041);
or U17491 (N_17491,N_12832,N_12247);
nand U17492 (N_17492,N_12071,N_12786);
and U17493 (N_17493,N_11148,N_10960);
nor U17494 (N_17494,N_11413,N_10156);
nor U17495 (N_17495,N_11796,N_14939);
nand U17496 (N_17496,N_12717,N_12337);
xnor U17497 (N_17497,N_13387,N_11740);
or U17498 (N_17498,N_10596,N_10888);
and U17499 (N_17499,N_10321,N_11790);
xor U17500 (N_17500,N_11738,N_12007);
nor U17501 (N_17501,N_12443,N_13106);
nand U17502 (N_17502,N_13900,N_10199);
nor U17503 (N_17503,N_10063,N_11713);
or U17504 (N_17504,N_10349,N_12803);
or U17505 (N_17505,N_10048,N_13461);
nand U17506 (N_17506,N_10022,N_11095);
nor U17507 (N_17507,N_13923,N_13100);
and U17508 (N_17508,N_13582,N_14769);
nor U17509 (N_17509,N_10512,N_10043);
xnor U17510 (N_17510,N_13029,N_13836);
and U17511 (N_17511,N_14236,N_13079);
xnor U17512 (N_17512,N_13428,N_11987);
or U17513 (N_17513,N_14883,N_11943);
nor U17514 (N_17514,N_13644,N_14464);
and U17515 (N_17515,N_13169,N_12540);
or U17516 (N_17516,N_14122,N_12414);
and U17517 (N_17517,N_12739,N_13529);
xor U17518 (N_17518,N_11956,N_13829);
or U17519 (N_17519,N_12894,N_12820);
and U17520 (N_17520,N_14542,N_14115);
nand U17521 (N_17521,N_12012,N_10314);
or U17522 (N_17522,N_14271,N_14698);
or U17523 (N_17523,N_13779,N_10504);
xnor U17524 (N_17524,N_10711,N_11892);
and U17525 (N_17525,N_12580,N_14891);
xnor U17526 (N_17526,N_14719,N_12007);
or U17527 (N_17527,N_13442,N_12199);
or U17528 (N_17528,N_10381,N_12942);
nand U17529 (N_17529,N_12793,N_11586);
and U17530 (N_17530,N_13805,N_10510);
and U17531 (N_17531,N_10761,N_12052);
xor U17532 (N_17532,N_10681,N_12980);
and U17533 (N_17533,N_10635,N_11438);
nand U17534 (N_17534,N_14470,N_10461);
or U17535 (N_17535,N_10103,N_14181);
or U17536 (N_17536,N_12197,N_14628);
or U17537 (N_17537,N_12001,N_10757);
nor U17538 (N_17538,N_11921,N_12793);
xor U17539 (N_17539,N_11109,N_11888);
and U17540 (N_17540,N_13107,N_11431);
nor U17541 (N_17541,N_13271,N_13971);
and U17542 (N_17542,N_14452,N_12473);
and U17543 (N_17543,N_13471,N_12254);
or U17544 (N_17544,N_14403,N_11239);
nor U17545 (N_17545,N_10084,N_11922);
or U17546 (N_17546,N_10901,N_12785);
nand U17547 (N_17547,N_10911,N_10888);
nand U17548 (N_17548,N_10592,N_11349);
and U17549 (N_17549,N_12868,N_12822);
or U17550 (N_17550,N_14028,N_12856);
nand U17551 (N_17551,N_11259,N_12126);
or U17552 (N_17552,N_13450,N_12967);
and U17553 (N_17553,N_11962,N_12842);
or U17554 (N_17554,N_11776,N_14124);
or U17555 (N_17555,N_13906,N_11937);
or U17556 (N_17556,N_10047,N_14249);
nor U17557 (N_17557,N_13152,N_13481);
and U17558 (N_17558,N_12862,N_13378);
and U17559 (N_17559,N_11372,N_14635);
or U17560 (N_17560,N_14464,N_13464);
xor U17561 (N_17561,N_10800,N_14451);
nor U17562 (N_17562,N_13250,N_14100);
xnor U17563 (N_17563,N_13430,N_12168);
or U17564 (N_17564,N_10451,N_11363);
nand U17565 (N_17565,N_12722,N_10565);
or U17566 (N_17566,N_12950,N_12798);
nand U17567 (N_17567,N_11342,N_11299);
xnor U17568 (N_17568,N_12747,N_11282);
and U17569 (N_17569,N_11030,N_14830);
nor U17570 (N_17570,N_11043,N_14576);
nand U17571 (N_17571,N_11140,N_10600);
nand U17572 (N_17572,N_12614,N_13018);
xor U17573 (N_17573,N_11700,N_14802);
nand U17574 (N_17574,N_13209,N_10215);
nor U17575 (N_17575,N_10504,N_12010);
and U17576 (N_17576,N_12476,N_13001);
xor U17577 (N_17577,N_11212,N_12226);
nand U17578 (N_17578,N_14536,N_11615);
nor U17579 (N_17579,N_13897,N_10019);
nand U17580 (N_17580,N_11877,N_14850);
and U17581 (N_17581,N_14811,N_10607);
or U17582 (N_17582,N_13212,N_10957);
nor U17583 (N_17583,N_12810,N_12376);
and U17584 (N_17584,N_13404,N_14655);
xor U17585 (N_17585,N_14273,N_14074);
or U17586 (N_17586,N_12048,N_12755);
nor U17587 (N_17587,N_11169,N_12034);
nand U17588 (N_17588,N_10197,N_11310);
and U17589 (N_17589,N_14212,N_11036);
nor U17590 (N_17590,N_14973,N_10211);
or U17591 (N_17591,N_14400,N_14915);
nand U17592 (N_17592,N_14899,N_11118);
nand U17593 (N_17593,N_14547,N_13049);
nand U17594 (N_17594,N_10405,N_11079);
and U17595 (N_17595,N_10347,N_13290);
nor U17596 (N_17596,N_13095,N_11067);
nor U17597 (N_17597,N_11502,N_11335);
xnor U17598 (N_17598,N_13249,N_12503);
or U17599 (N_17599,N_10970,N_13729);
xnor U17600 (N_17600,N_13885,N_11021);
nand U17601 (N_17601,N_12598,N_14399);
xnor U17602 (N_17602,N_12020,N_13957);
nor U17603 (N_17603,N_11106,N_11502);
nand U17604 (N_17604,N_14120,N_11989);
and U17605 (N_17605,N_11083,N_12197);
nor U17606 (N_17606,N_13241,N_14039);
and U17607 (N_17607,N_10819,N_13700);
nand U17608 (N_17608,N_10646,N_12698);
nand U17609 (N_17609,N_12625,N_13237);
or U17610 (N_17610,N_12934,N_13585);
nand U17611 (N_17611,N_13116,N_10368);
xnor U17612 (N_17612,N_10740,N_13618);
nand U17613 (N_17613,N_13090,N_10573);
xnor U17614 (N_17614,N_14791,N_10464);
or U17615 (N_17615,N_13885,N_10831);
nand U17616 (N_17616,N_11553,N_11656);
nand U17617 (N_17617,N_10519,N_14848);
xnor U17618 (N_17618,N_13923,N_14242);
or U17619 (N_17619,N_13797,N_10154);
or U17620 (N_17620,N_11865,N_14461);
or U17621 (N_17621,N_13357,N_11663);
xnor U17622 (N_17622,N_11169,N_10933);
xor U17623 (N_17623,N_10036,N_14654);
or U17624 (N_17624,N_13053,N_13648);
nor U17625 (N_17625,N_12371,N_14823);
and U17626 (N_17626,N_11990,N_12137);
xnor U17627 (N_17627,N_14666,N_14776);
and U17628 (N_17628,N_11396,N_14046);
and U17629 (N_17629,N_11162,N_11395);
nand U17630 (N_17630,N_11865,N_10466);
and U17631 (N_17631,N_12951,N_10445);
and U17632 (N_17632,N_13805,N_13657);
nand U17633 (N_17633,N_12106,N_11257);
nor U17634 (N_17634,N_13813,N_13535);
nor U17635 (N_17635,N_11667,N_10431);
and U17636 (N_17636,N_12544,N_10303);
nand U17637 (N_17637,N_14486,N_13621);
nand U17638 (N_17638,N_11198,N_11615);
nor U17639 (N_17639,N_11965,N_12412);
nor U17640 (N_17640,N_12190,N_11248);
xnor U17641 (N_17641,N_14738,N_11387);
nand U17642 (N_17642,N_14909,N_10414);
nor U17643 (N_17643,N_10860,N_10672);
nor U17644 (N_17644,N_13039,N_10319);
or U17645 (N_17645,N_13820,N_13430);
and U17646 (N_17646,N_11209,N_14316);
nand U17647 (N_17647,N_12494,N_14491);
nand U17648 (N_17648,N_11640,N_12097);
nor U17649 (N_17649,N_11345,N_13140);
nand U17650 (N_17650,N_12705,N_13897);
xor U17651 (N_17651,N_10746,N_10755);
or U17652 (N_17652,N_12852,N_11695);
xnor U17653 (N_17653,N_11640,N_14618);
and U17654 (N_17654,N_14238,N_13663);
and U17655 (N_17655,N_12215,N_12676);
and U17656 (N_17656,N_12675,N_13794);
or U17657 (N_17657,N_14708,N_14617);
and U17658 (N_17658,N_10457,N_14469);
nand U17659 (N_17659,N_14749,N_10018);
and U17660 (N_17660,N_12085,N_12263);
and U17661 (N_17661,N_12290,N_11835);
nand U17662 (N_17662,N_10569,N_12851);
and U17663 (N_17663,N_13500,N_12027);
and U17664 (N_17664,N_13010,N_10736);
nand U17665 (N_17665,N_11899,N_14948);
and U17666 (N_17666,N_10192,N_14022);
nand U17667 (N_17667,N_12336,N_11391);
and U17668 (N_17668,N_13129,N_14229);
nor U17669 (N_17669,N_13004,N_11527);
nand U17670 (N_17670,N_12248,N_10386);
or U17671 (N_17671,N_12582,N_10519);
xor U17672 (N_17672,N_11709,N_10581);
nand U17673 (N_17673,N_14573,N_10712);
and U17674 (N_17674,N_14745,N_12402);
and U17675 (N_17675,N_12830,N_12969);
and U17676 (N_17676,N_12195,N_13856);
and U17677 (N_17677,N_10073,N_13869);
nand U17678 (N_17678,N_10911,N_10940);
nor U17679 (N_17679,N_14326,N_14548);
or U17680 (N_17680,N_13094,N_12172);
or U17681 (N_17681,N_14517,N_11673);
or U17682 (N_17682,N_10195,N_10055);
and U17683 (N_17683,N_14026,N_10737);
and U17684 (N_17684,N_10666,N_10089);
xnor U17685 (N_17685,N_10204,N_11111);
xnor U17686 (N_17686,N_10999,N_12484);
nand U17687 (N_17687,N_12029,N_13148);
and U17688 (N_17688,N_10488,N_14552);
nor U17689 (N_17689,N_12432,N_11232);
nand U17690 (N_17690,N_13264,N_10199);
and U17691 (N_17691,N_10593,N_10209);
and U17692 (N_17692,N_12283,N_11872);
nor U17693 (N_17693,N_12575,N_14876);
and U17694 (N_17694,N_12029,N_14829);
and U17695 (N_17695,N_10909,N_10815);
nor U17696 (N_17696,N_14099,N_10323);
nor U17697 (N_17697,N_14961,N_10563);
nor U17698 (N_17698,N_14146,N_12503);
nor U17699 (N_17699,N_11618,N_11684);
nor U17700 (N_17700,N_12629,N_10676);
xnor U17701 (N_17701,N_11336,N_11364);
or U17702 (N_17702,N_12269,N_10931);
and U17703 (N_17703,N_13597,N_14948);
nor U17704 (N_17704,N_10792,N_12876);
xnor U17705 (N_17705,N_14474,N_11156);
nand U17706 (N_17706,N_12209,N_10849);
nor U17707 (N_17707,N_12513,N_14362);
or U17708 (N_17708,N_13078,N_14312);
nor U17709 (N_17709,N_13779,N_13943);
nand U17710 (N_17710,N_10123,N_14762);
and U17711 (N_17711,N_11723,N_12300);
xnor U17712 (N_17712,N_10408,N_12696);
or U17713 (N_17713,N_14154,N_11105);
xnor U17714 (N_17714,N_10544,N_10920);
nor U17715 (N_17715,N_11031,N_11266);
nand U17716 (N_17716,N_14079,N_10025);
nand U17717 (N_17717,N_10457,N_10995);
xor U17718 (N_17718,N_12995,N_14174);
xor U17719 (N_17719,N_13631,N_10703);
and U17720 (N_17720,N_14403,N_10206);
and U17721 (N_17721,N_11163,N_14323);
xnor U17722 (N_17722,N_13364,N_13730);
or U17723 (N_17723,N_10416,N_14576);
and U17724 (N_17724,N_13549,N_13255);
and U17725 (N_17725,N_10397,N_14958);
nand U17726 (N_17726,N_14104,N_11611);
nand U17727 (N_17727,N_10321,N_14656);
xnor U17728 (N_17728,N_10194,N_10298);
nor U17729 (N_17729,N_12689,N_11888);
nand U17730 (N_17730,N_13221,N_11774);
nor U17731 (N_17731,N_13456,N_13559);
and U17732 (N_17732,N_13919,N_12725);
nand U17733 (N_17733,N_10819,N_10018);
xnor U17734 (N_17734,N_10141,N_11360);
nand U17735 (N_17735,N_11291,N_10772);
and U17736 (N_17736,N_12925,N_13102);
nand U17737 (N_17737,N_13432,N_10061);
nor U17738 (N_17738,N_11122,N_11069);
nor U17739 (N_17739,N_12856,N_12571);
nor U17740 (N_17740,N_11198,N_11413);
or U17741 (N_17741,N_11788,N_14358);
nor U17742 (N_17742,N_13157,N_14921);
and U17743 (N_17743,N_10781,N_12555);
xor U17744 (N_17744,N_14997,N_14941);
xor U17745 (N_17745,N_13214,N_14338);
nand U17746 (N_17746,N_10516,N_11964);
and U17747 (N_17747,N_14711,N_10531);
xor U17748 (N_17748,N_13087,N_12242);
xor U17749 (N_17749,N_12935,N_13837);
xor U17750 (N_17750,N_10406,N_14439);
and U17751 (N_17751,N_13862,N_12735);
nand U17752 (N_17752,N_12786,N_12323);
xnor U17753 (N_17753,N_12639,N_11825);
nor U17754 (N_17754,N_11869,N_14539);
nand U17755 (N_17755,N_10187,N_12364);
nor U17756 (N_17756,N_14489,N_12233);
nand U17757 (N_17757,N_10175,N_12789);
nor U17758 (N_17758,N_12444,N_12871);
xor U17759 (N_17759,N_12855,N_11282);
xor U17760 (N_17760,N_11173,N_12828);
xor U17761 (N_17761,N_12076,N_12465);
or U17762 (N_17762,N_14267,N_12337);
or U17763 (N_17763,N_13036,N_12581);
nor U17764 (N_17764,N_14864,N_13593);
nand U17765 (N_17765,N_14070,N_14226);
or U17766 (N_17766,N_14597,N_11332);
xnor U17767 (N_17767,N_13669,N_10880);
nor U17768 (N_17768,N_11531,N_14544);
xnor U17769 (N_17769,N_11559,N_12077);
nand U17770 (N_17770,N_14068,N_11311);
and U17771 (N_17771,N_12905,N_14932);
xnor U17772 (N_17772,N_12878,N_12480);
or U17773 (N_17773,N_14005,N_13215);
or U17774 (N_17774,N_12808,N_12014);
nor U17775 (N_17775,N_12210,N_11410);
or U17776 (N_17776,N_13611,N_14482);
xnor U17777 (N_17777,N_12530,N_14565);
nand U17778 (N_17778,N_12661,N_14122);
xor U17779 (N_17779,N_13142,N_14265);
and U17780 (N_17780,N_12670,N_10130);
and U17781 (N_17781,N_14828,N_11794);
and U17782 (N_17782,N_11906,N_12837);
nor U17783 (N_17783,N_10310,N_13221);
nand U17784 (N_17784,N_13154,N_14911);
nand U17785 (N_17785,N_14255,N_12719);
or U17786 (N_17786,N_11401,N_11476);
and U17787 (N_17787,N_10266,N_12982);
xor U17788 (N_17788,N_10235,N_12399);
or U17789 (N_17789,N_14690,N_14196);
and U17790 (N_17790,N_11429,N_10477);
xnor U17791 (N_17791,N_14814,N_12512);
nor U17792 (N_17792,N_11855,N_14418);
or U17793 (N_17793,N_12416,N_13610);
or U17794 (N_17794,N_12342,N_14829);
xnor U17795 (N_17795,N_14024,N_10471);
or U17796 (N_17796,N_14777,N_14195);
or U17797 (N_17797,N_13446,N_13201);
xor U17798 (N_17798,N_10888,N_10352);
nor U17799 (N_17799,N_13885,N_11972);
or U17800 (N_17800,N_13670,N_12505);
xnor U17801 (N_17801,N_10052,N_14947);
nand U17802 (N_17802,N_13390,N_13502);
and U17803 (N_17803,N_10919,N_12781);
nor U17804 (N_17804,N_10448,N_10365);
xnor U17805 (N_17805,N_11865,N_12054);
and U17806 (N_17806,N_12806,N_11106);
xor U17807 (N_17807,N_10793,N_12418);
and U17808 (N_17808,N_13984,N_12832);
or U17809 (N_17809,N_13575,N_12486);
xnor U17810 (N_17810,N_13921,N_13944);
and U17811 (N_17811,N_14070,N_10836);
and U17812 (N_17812,N_12395,N_14479);
or U17813 (N_17813,N_13246,N_11225);
xnor U17814 (N_17814,N_12909,N_14054);
and U17815 (N_17815,N_12318,N_14169);
and U17816 (N_17816,N_11900,N_13414);
or U17817 (N_17817,N_12543,N_10555);
and U17818 (N_17818,N_10644,N_10252);
or U17819 (N_17819,N_13325,N_12502);
and U17820 (N_17820,N_14076,N_14869);
nor U17821 (N_17821,N_12045,N_10870);
nand U17822 (N_17822,N_10465,N_10527);
and U17823 (N_17823,N_12851,N_14403);
and U17824 (N_17824,N_12778,N_11061);
and U17825 (N_17825,N_13525,N_11096);
and U17826 (N_17826,N_10544,N_13239);
and U17827 (N_17827,N_11795,N_11965);
and U17828 (N_17828,N_13911,N_10540);
or U17829 (N_17829,N_10151,N_12061);
nand U17830 (N_17830,N_10770,N_11224);
nor U17831 (N_17831,N_10567,N_12659);
nor U17832 (N_17832,N_14713,N_11328);
and U17833 (N_17833,N_10158,N_12633);
xor U17834 (N_17834,N_13435,N_11355);
nand U17835 (N_17835,N_11364,N_14950);
or U17836 (N_17836,N_11029,N_12476);
nor U17837 (N_17837,N_13261,N_13634);
xor U17838 (N_17838,N_11708,N_12911);
xor U17839 (N_17839,N_11892,N_12835);
nand U17840 (N_17840,N_12951,N_11826);
nor U17841 (N_17841,N_10486,N_14197);
or U17842 (N_17842,N_12686,N_11847);
xor U17843 (N_17843,N_10963,N_14849);
or U17844 (N_17844,N_14790,N_11278);
nand U17845 (N_17845,N_10224,N_11854);
nor U17846 (N_17846,N_11303,N_13883);
nor U17847 (N_17847,N_12325,N_13241);
nand U17848 (N_17848,N_11068,N_13349);
nand U17849 (N_17849,N_14589,N_12144);
xor U17850 (N_17850,N_12743,N_12391);
nand U17851 (N_17851,N_13057,N_10107);
xnor U17852 (N_17852,N_11554,N_14976);
nor U17853 (N_17853,N_11464,N_12415);
nand U17854 (N_17854,N_13408,N_14071);
nor U17855 (N_17855,N_13142,N_12774);
xnor U17856 (N_17856,N_14673,N_11012);
or U17857 (N_17857,N_10524,N_10500);
or U17858 (N_17858,N_13601,N_10052);
nand U17859 (N_17859,N_12495,N_12707);
xnor U17860 (N_17860,N_14937,N_12243);
and U17861 (N_17861,N_10729,N_10225);
or U17862 (N_17862,N_12884,N_14741);
nor U17863 (N_17863,N_13130,N_12847);
xor U17864 (N_17864,N_10934,N_13208);
nor U17865 (N_17865,N_14984,N_13393);
nand U17866 (N_17866,N_10970,N_11818);
nand U17867 (N_17867,N_13010,N_10150);
nor U17868 (N_17868,N_11354,N_13871);
nor U17869 (N_17869,N_11015,N_13054);
or U17870 (N_17870,N_11522,N_10550);
nand U17871 (N_17871,N_12657,N_13001);
xnor U17872 (N_17872,N_10613,N_11001);
nand U17873 (N_17873,N_10887,N_11973);
nand U17874 (N_17874,N_14305,N_13393);
xnor U17875 (N_17875,N_13903,N_13441);
and U17876 (N_17876,N_12820,N_12259);
or U17877 (N_17877,N_10691,N_10184);
nor U17878 (N_17878,N_13573,N_12182);
xor U17879 (N_17879,N_12436,N_11487);
nor U17880 (N_17880,N_11396,N_13664);
or U17881 (N_17881,N_14673,N_12421);
nand U17882 (N_17882,N_10016,N_14949);
nor U17883 (N_17883,N_13642,N_12541);
xnor U17884 (N_17884,N_12184,N_12135);
nand U17885 (N_17885,N_11958,N_13355);
or U17886 (N_17886,N_11371,N_13941);
and U17887 (N_17887,N_11344,N_12477);
and U17888 (N_17888,N_14925,N_10252);
xnor U17889 (N_17889,N_11512,N_14390);
nand U17890 (N_17890,N_11516,N_12107);
or U17891 (N_17891,N_14927,N_13765);
and U17892 (N_17892,N_13304,N_12371);
xor U17893 (N_17893,N_10285,N_12087);
xor U17894 (N_17894,N_10594,N_12330);
nor U17895 (N_17895,N_12912,N_13062);
and U17896 (N_17896,N_10387,N_11407);
xor U17897 (N_17897,N_13843,N_10249);
and U17898 (N_17898,N_14291,N_11529);
and U17899 (N_17899,N_11896,N_13086);
or U17900 (N_17900,N_14334,N_14258);
nand U17901 (N_17901,N_10489,N_13536);
nor U17902 (N_17902,N_11887,N_12851);
xnor U17903 (N_17903,N_13417,N_11528);
nor U17904 (N_17904,N_12397,N_13426);
nand U17905 (N_17905,N_12519,N_14807);
or U17906 (N_17906,N_13984,N_13196);
xor U17907 (N_17907,N_11852,N_14948);
and U17908 (N_17908,N_10240,N_10396);
xor U17909 (N_17909,N_10072,N_13910);
xor U17910 (N_17910,N_10118,N_13111);
or U17911 (N_17911,N_11723,N_12704);
or U17912 (N_17912,N_10849,N_14112);
nand U17913 (N_17913,N_13492,N_10994);
nor U17914 (N_17914,N_12317,N_11325);
xor U17915 (N_17915,N_11441,N_10389);
xnor U17916 (N_17916,N_10301,N_13374);
and U17917 (N_17917,N_11089,N_11301);
xor U17918 (N_17918,N_13027,N_14411);
or U17919 (N_17919,N_14224,N_13296);
and U17920 (N_17920,N_10026,N_10608);
or U17921 (N_17921,N_11928,N_11746);
nor U17922 (N_17922,N_11032,N_14439);
xnor U17923 (N_17923,N_14414,N_11788);
or U17924 (N_17924,N_13532,N_12292);
nand U17925 (N_17925,N_11635,N_11456);
nor U17926 (N_17926,N_11202,N_11342);
nand U17927 (N_17927,N_12512,N_11081);
or U17928 (N_17928,N_12726,N_13128);
and U17929 (N_17929,N_11515,N_14266);
and U17930 (N_17930,N_11757,N_11005);
nor U17931 (N_17931,N_11636,N_13883);
or U17932 (N_17932,N_10420,N_12039);
nand U17933 (N_17933,N_14959,N_14690);
or U17934 (N_17934,N_13244,N_10769);
or U17935 (N_17935,N_10032,N_13895);
nor U17936 (N_17936,N_12604,N_12064);
nor U17937 (N_17937,N_10849,N_14868);
nor U17938 (N_17938,N_10154,N_13329);
and U17939 (N_17939,N_14029,N_10956);
nor U17940 (N_17940,N_10519,N_12326);
xor U17941 (N_17941,N_13974,N_13288);
nor U17942 (N_17942,N_12839,N_10526);
or U17943 (N_17943,N_13044,N_14529);
nand U17944 (N_17944,N_14845,N_12035);
and U17945 (N_17945,N_10443,N_14856);
and U17946 (N_17946,N_13593,N_12207);
or U17947 (N_17947,N_10363,N_13441);
or U17948 (N_17948,N_12077,N_10169);
and U17949 (N_17949,N_14378,N_13248);
or U17950 (N_17950,N_14074,N_11134);
nand U17951 (N_17951,N_13396,N_11897);
xnor U17952 (N_17952,N_14064,N_10956);
or U17953 (N_17953,N_10374,N_13596);
or U17954 (N_17954,N_12810,N_14160);
nor U17955 (N_17955,N_12051,N_13806);
or U17956 (N_17956,N_11872,N_11681);
xnor U17957 (N_17957,N_11263,N_14272);
or U17958 (N_17958,N_10967,N_14777);
nor U17959 (N_17959,N_10642,N_13726);
xor U17960 (N_17960,N_14459,N_12050);
nand U17961 (N_17961,N_12219,N_12161);
xnor U17962 (N_17962,N_10328,N_13728);
or U17963 (N_17963,N_14158,N_12787);
nand U17964 (N_17964,N_11104,N_12223);
xnor U17965 (N_17965,N_11671,N_12729);
nand U17966 (N_17966,N_11260,N_13906);
xnor U17967 (N_17967,N_13614,N_12906);
and U17968 (N_17968,N_14714,N_13103);
xor U17969 (N_17969,N_11905,N_10923);
xor U17970 (N_17970,N_14982,N_14353);
or U17971 (N_17971,N_10510,N_11752);
and U17972 (N_17972,N_14108,N_11043);
and U17973 (N_17973,N_11799,N_14491);
xnor U17974 (N_17974,N_14356,N_14128);
nand U17975 (N_17975,N_13458,N_12730);
or U17976 (N_17976,N_12698,N_12492);
xnor U17977 (N_17977,N_14543,N_10180);
or U17978 (N_17978,N_11025,N_12638);
nand U17979 (N_17979,N_11957,N_14980);
nor U17980 (N_17980,N_11825,N_13017);
nor U17981 (N_17981,N_12467,N_10216);
nor U17982 (N_17982,N_10108,N_10474);
nand U17983 (N_17983,N_12895,N_12726);
nand U17984 (N_17984,N_12824,N_13970);
xor U17985 (N_17985,N_10077,N_11613);
nand U17986 (N_17986,N_10939,N_13898);
and U17987 (N_17987,N_13394,N_10913);
nor U17988 (N_17988,N_13373,N_11972);
nor U17989 (N_17989,N_14088,N_11845);
or U17990 (N_17990,N_14738,N_13274);
xnor U17991 (N_17991,N_11983,N_14058);
xor U17992 (N_17992,N_10673,N_12492);
or U17993 (N_17993,N_13458,N_14152);
and U17994 (N_17994,N_11940,N_12816);
nand U17995 (N_17995,N_14083,N_10688);
and U17996 (N_17996,N_11728,N_13719);
xor U17997 (N_17997,N_10778,N_13244);
nand U17998 (N_17998,N_14473,N_10552);
or U17999 (N_17999,N_13493,N_14099);
and U18000 (N_18000,N_13970,N_10717);
or U18001 (N_18001,N_12169,N_14779);
and U18002 (N_18002,N_14054,N_12818);
and U18003 (N_18003,N_13970,N_10237);
or U18004 (N_18004,N_10106,N_14944);
nand U18005 (N_18005,N_11822,N_12307);
nand U18006 (N_18006,N_12738,N_13434);
nand U18007 (N_18007,N_12276,N_10718);
and U18008 (N_18008,N_14112,N_12998);
nand U18009 (N_18009,N_12141,N_10895);
nor U18010 (N_18010,N_10719,N_11958);
nor U18011 (N_18011,N_10230,N_10106);
nand U18012 (N_18012,N_11982,N_12344);
nand U18013 (N_18013,N_13532,N_11130);
nand U18014 (N_18014,N_14588,N_13306);
and U18015 (N_18015,N_10118,N_13216);
nor U18016 (N_18016,N_10642,N_11328);
nand U18017 (N_18017,N_13751,N_13048);
nand U18018 (N_18018,N_14124,N_14412);
or U18019 (N_18019,N_14538,N_13109);
and U18020 (N_18020,N_13348,N_10410);
nand U18021 (N_18021,N_11275,N_10387);
nand U18022 (N_18022,N_14866,N_14645);
and U18023 (N_18023,N_12362,N_14701);
or U18024 (N_18024,N_11368,N_13939);
nor U18025 (N_18025,N_14797,N_11919);
xor U18026 (N_18026,N_11495,N_13264);
and U18027 (N_18027,N_11814,N_12622);
nor U18028 (N_18028,N_13433,N_10706);
and U18029 (N_18029,N_11576,N_14298);
xnor U18030 (N_18030,N_10292,N_14968);
xnor U18031 (N_18031,N_13181,N_11021);
nor U18032 (N_18032,N_13359,N_14090);
xor U18033 (N_18033,N_11707,N_14692);
xor U18034 (N_18034,N_11786,N_12947);
and U18035 (N_18035,N_13660,N_12746);
nand U18036 (N_18036,N_14648,N_13864);
or U18037 (N_18037,N_14325,N_13993);
nand U18038 (N_18038,N_14152,N_14151);
and U18039 (N_18039,N_10743,N_13141);
xnor U18040 (N_18040,N_10433,N_13473);
nand U18041 (N_18041,N_12318,N_11867);
or U18042 (N_18042,N_14186,N_10512);
nor U18043 (N_18043,N_10711,N_14172);
nor U18044 (N_18044,N_11579,N_12310);
and U18045 (N_18045,N_14125,N_12954);
nor U18046 (N_18046,N_14058,N_14391);
nor U18047 (N_18047,N_10541,N_11112);
or U18048 (N_18048,N_14604,N_12313);
and U18049 (N_18049,N_12039,N_12237);
nor U18050 (N_18050,N_11953,N_13805);
nand U18051 (N_18051,N_11570,N_13354);
nor U18052 (N_18052,N_14302,N_13930);
nand U18053 (N_18053,N_12595,N_13280);
nor U18054 (N_18054,N_12309,N_13988);
nor U18055 (N_18055,N_11256,N_13649);
nor U18056 (N_18056,N_14483,N_11837);
and U18057 (N_18057,N_11230,N_14800);
nand U18058 (N_18058,N_12761,N_13783);
or U18059 (N_18059,N_14285,N_14260);
or U18060 (N_18060,N_11352,N_11033);
and U18061 (N_18061,N_12755,N_13335);
nand U18062 (N_18062,N_14889,N_10566);
xnor U18063 (N_18063,N_12365,N_14248);
xor U18064 (N_18064,N_13963,N_10431);
nor U18065 (N_18065,N_13702,N_11890);
xnor U18066 (N_18066,N_14482,N_10356);
xnor U18067 (N_18067,N_10512,N_13726);
xnor U18068 (N_18068,N_11087,N_11756);
or U18069 (N_18069,N_10410,N_12229);
nand U18070 (N_18070,N_12058,N_14526);
or U18071 (N_18071,N_12626,N_13482);
xor U18072 (N_18072,N_11597,N_12537);
nand U18073 (N_18073,N_14599,N_13779);
or U18074 (N_18074,N_13977,N_11426);
and U18075 (N_18075,N_12419,N_11575);
xnor U18076 (N_18076,N_11544,N_13207);
or U18077 (N_18077,N_11085,N_10548);
or U18078 (N_18078,N_10969,N_14487);
nand U18079 (N_18079,N_12244,N_12318);
and U18080 (N_18080,N_11740,N_12228);
and U18081 (N_18081,N_10291,N_14473);
or U18082 (N_18082,N_13452,N_11857);
or U18083 (N_18083,N_14091,N_12519);
and U18084 (N_18084,N_11695,N_13186);
or U18085 (N_18085,N_12311,N_14906);
and U18086 (N_18086,N_12870,N_14732);
or U18087 (N_18087,N_10248,N_14249);
or U18088 (N_18088,N_13227,N_14105);
and U18089 (N_18089,N_14926,N_14504);
or U18090 (N_18090,N_13159,N_12985);
nor U18091 (N_18091,N_12363,N_12760);
xor U18092 (N_18092,N_10284,N_10106);
nor U18093 (N_18093,N_10365,N_14151);
or U18094 (N_18094,N_11666,N_11451);
and U18095 (N_18095,N_10602,N_14898);
and U18096 (N_18096,N_10765,N_11515);
xnor U18097 (N_18097,N_10183,N_14006);
or U18098 (N_18098,N_14969,N_12124);
or U18099 (N_18099,N_12397,N_12564);
and U18100 (N_18100,N_11672,N_14810);
nor U18101 (N_18101,N_14239,N_12527);
nor U18102 (N_18102,N_12798,N_10889);
nor U18103 (N_18103,N_10935,N_13792);
and U18104 (N_18104,N_12512,N_14672);
xnor U18105 (N_18105,N_10897,N_14985);
nor U18106 (N_18106,N_10908,N_10994);
nand U18107 (N_18107,N_14663,N_11510);
xnor U18108 (N_18108,N_11240,N_14022);
or U18109 (N_18109,N_10822,N_14511);
nand U18110 (N_18110,N_14320,N_13104);
and U18111 (N_18111,N_10145,N_12905);
and U18112 (N_18112,N_13700,N_10686);
nand U18113 (N_18113,N_14450,N_13365);
nand U18114 (N_18114,N_12449,N_10652);
nor U18115 (N_18115,N_13052,N_11356);
nand U18116 (N_18116,N_11499,N_14152);
and U18117 (N_18117,N_13024,N_13875);
xnor U18118 (N_18118,N_12593,N_14854);
and U18119 (N_18119,N_12384,N_11713);
nor U18120 (N_18120,N_11765,N_10026);
or U18121 (N_18121,N_13269,N_13467);
nor U18122 (N_18122,N_14733,N_14616);
or U18123 (N_18123,N_11516,N_10425);
and U18124 (N_18124,N_11858,N_11903);
and U18125 (N_18125,N_14951,N_14431);
or U18126 (N_18126,N_12001,N_12968);
nor U18127 (N_18127,N_13758,N_12860);
and U18128 (N_18128,N_12946,N_14369);
or U18129 (N_18129,N_14646,N_10417);
or U18130 (N_18130,N_10167,N_12885);
nand U18131 (N_18131,N_10431,N_13091);
nand U18132 (N_18132,N_14785,N_14579);
xor U18133 (N_18133,N_10890,N_12696);
and U18134 (N_18134,N_14402,N_11154);
and U18135 (N_18135,N_13471,N_12850);
or U18136 (N_18136,N_14215,N_14440);
nand U18137 (N_18137,N_13137,N_14162);
or U18138 (N_18138,N_14572,N_12569);
nor U18139 (N_18139,N_12692,N_10671);
or U18140 (N_18140,N_10833,N_12689);
and U18141 (N_18141,N_14447,N_14646);
xnor U18142 (N_18142,N_12009,N_14204);
nor U18143 (N_18143,N_12902,N_14861);
or U18144 (N_18144,N_13560,N_12737);
xnor U18145 (N_18145,N_14761,N_10896);
nor U18146 (N_18146,N_10663,N_11900);
nand U18147 (N_18147,N_12237,N_14600);
nand U18148 (N_18148,N_10257,N_11199);
xor U18149 (N_18149,N_13894,N_12347);
or U18150 (N_18150,N_14836,N_13763);
or U18151 (N_18151,N_10982,N_13655);
or U18152 (N_18152,N_10835,N_14932);
nor U18153 (N_18153,N_10744,N_13800);
xor U18154 (N_18154,N_11001,N_10816);
nand U18155 (N_18155,N_13247,N_12647);
and U18156 (N_18156,N_14403,N_11121);
or U18157 (N_18157,N_12497,N_10160);
or U18158 (N_18158,N_10235,N_13073);
nor U18159 (N_18159,N_14981,N_14183);
nand U18160 (N_18160,N_13353,N_14419);
and U18161 (N_18161,N_10579,N_13280);
nand U18162 (N_18162,N_13242,N_12061);
nand U18163 (N_18163,N_11008,N_14006);
nand U18164 (N_18164,N_11585,N_12805);
nor U18165 (N_18165,N_14886,N_11532);
xor U18166 (N_18166,N_11472,N_14646);
or U18167 (N_18167,N_12813,N_12696);
nand U18168 (N_18168,N_10546,N_12236);
or U18169 (N_18169,N_14596,N_13896);
and U18170 (N_18170,N_14637,N_11888);
nor U18171 (N_18171,N_14324,N_11168);
and U18172 (N_18172,N_10412,N_11379);
or U18173 (N_18173,N_14303,N_12634);
nor U18174 (N_18174,N_12280,N_14292);
nor U18175 (N_18175,N_10173,N_14621);
or U18176 (N_18176,N_13016,N_12017);
nand U18177 (N_18177,N_11770,N_13705);
nand U18178 (N_18178,N_12347,N_13198);
or U18179 (N_18179,N_14857,N_10770);
nand U18180 (N_18180,N_10560,N_14245);
and U18181 (N_18181,N_12247,N_10146);
nor U18182 (N_18182,N_13143,N_11782);
or U18183 (N_18183,N_12033,N_10167);
and U18184 (N_18184,N_13225,N_13709);
and U18185 (N_18185,N_11058,N_14264);
and U18186 (N_18186,N_10511,N_12437);
or U18187 (N_18187,N_14208,N_14670);
or U18188 (N_18188,N_11586,N_10988);
and U18189 (N_18189,N_11751,N_10276);
nand U18190 (N_18190,N_11435,N_12691);
xor U18191 (N_18191,N_14149,N_14507);
and U18192 (N_18192,N_10065,N_11186);
nand U18193 (N_18193,N_14035,N_12030);
nor U18194 (N_18194,N_13253,N_12856);
or U18195 (N_18195,N_12264,N_14462);
nor U18196 (N_18196,N_13761,N_12570);
nand U18197 (N_18197,N_10731,N_14570);
or U18198 (N_18198,N_11188,N_14264);
or U18199 (N_18199,N_14412,N_10852);
nand U18200 (N_18200,N_12662,N_13540);
or U18201 (N_18201,N_12222,N_14784);
and U18202 (N_18202,N_12512,N_12910);
and U18203 (N_18203,N_13993,N_13772);
nor U18204 (N_18204,N_11128,N_14715);
nand U18205 (N_18205,N_10636,N_14845);
nor U18206 (N_18206,N_12046,N_12427);
or U18207 (N_18207,N_11139,N_14791);
or U18208 (N_18208,N_10723,N_11764);
xnor U18209 (N_18209,N_10816,N_14632);
and U18210 (N_18210,N_11852,N_10892);
nand U18211 (N_18211,N_10589,N_10592);
nor U18212 (N_18212,N_12045,N_10894);
nand U18213 (N_18213,N_11814,N_12883);
nand U18214 (N_18214,N_11018,N_10720);
nor U18215 (N_18215,N_13485,N_12520);
nand U18216 (N_18216,N_10715,N_12242);
nand U18217 (N_18217,N_12417,N_11709);
or U18218 (N_18218,N_12493,N_13013);
nand U18219 (N_18219,N_14551,N_11155);
and U18220 (N_18220,N_14736,N_13751);
and U18221 (N_18221,N_13550,N_10063);
nor U18222 (N_18222,N_12019,N_13293);
and U18223 (N_18223,N_10618,N_12596);
nand U18224 (N_18224,N_10749,N_12353);
or U18225 (N_18225,N_13339,N_12130);
or U18226 (N_18226,N_12685,N_14636);
or U18227 (N_18227,N_14478,N_13841);
and U18228 (N_18228,N_14450,N_14985);
and U18229 (N_18229,N_11484,N_10075);
nor U18230 (N_18230,N_10528,N_12539);
and U18231 (N_18231,N_11549,N_10830);
nor U18232 (N_18232,N_14577,N_11516);
or U18233 (N_18233,N_13479,N_14736);
and U18234 (N_18234,N_10161,N_11015);
and U18235 (N_18235,N_14952,N_13835);
xnor U18236 (N_18236,N_10231,N_13221);
nand U18237 (N_18237,N_10732,N_11487);
or U18238 (N_18238,N_10478,N_12882);
xor U18239 (N_18239,N_10961,N_11600);
or U18240 (N_18240,N_11862,N_12788);
or U18241 (N_18241,N_14121,N_11605);
nor U18242 (N_18242,N_12893,N_12241);
or U18243 (N_18243,N_13109,N_10300);
nand U18244 (N_18244,N_11112,N_13068);
xnor U18245 (N_18245,N_11469,N_13684);
xnor U18246 (N_18246,N_10735,N_11973);
nand U18247 (N_18247,N_13224,N_11996);
nor U18248 (N_18248,N_11910,N_14544);
nor U18249 (N_18249,N_14462,N_12313);
or U18250 (N_18250,N_14116,N_12195);
nor U18251 (N_18251,N_13575,N_13192);
and U18252 (N_18252,N_12871,N_11074);
nand U18253 (N_18253,N_14172,N_13141);
nor U18254 (N_18254,N_14451,N_14102);
nand U18255 (N_18255,N_13543,N_10457);
xnor U18256 (N_18256,N_12779,N_10733);
or U18257 (N_18257,N_11774,N_14987);
or U18258 (N_18258,N_12460,N_13086);
nor U18259 (N_18259,N_11086,N_12048);
xor U18260 (N_18260,N_11641,N_13043);
xor U18261 (N_18261,N_12536,N_13179);
xnor U18262 (N_18262,N_12340,N_11614);
or U18263 (N_18263,N_13345,N_14917);
and U18264 (N_18264,N_14457,N_14710);
nor U18265 (N_18265,N_12944,N_13922);
xnor U18266 (N_18266,N_11103,N_12260);
and U18267 (N_18267,N_11694,N_10095);
nor U18268 (N_18268,N_11670,N_10243);
xor U18269 (N_18269,N_14911,N_13911);
and U18270 (N_18270,N_14312,N_13486);
nor U18271 (N_18271,N_11548,N_13823);
xor U18272 (N_18272,N_13473,N_14115);
or U18273 (N_18273,N_13451,N_10543);
and U18274 (N_18274,N_10299,N_14259);
nor U18275 (N_18275,N_14597,N_12835);
or U18276 (N_18276,N_13643,N_10992);
nand U18277 (N_18277,N_14282,N_13076);
nand U18278 (N_18278,N_12967,N_13854);
xor U18279 (N_18279,N_14015,N_13882);
or U18280 (N_18280,N_13794,N_12732);
nor U18281 (N_18281,N_14613,N_14839);
nor U18282 (N_18282,N_10696,N_14342);
or U18283 (N_18283,N_12401,N_12481);
or U18284 (N_18284,N_14228,N_12395);
or U18285 (N_18285,N_10332,N_13160);
nand U18286 (N_18286,N_10680,N_13845);
and U18287 (N_18287,N_12558,N_14132);
or U18288 (N_18288,N_14442,N_14166);
or U18289 (N_18289,N_10993,N_12597);
xor U18290 (N_18290,N_13352,N_13476);
and U18291 (N_18291,N_11301,N_11091);
or U18292 (N_18292,N_12809,N_14138);
and U18293 (N_18293,N_11229,N_12862);
nand U18294 (N_18294,N_12277,N_12465);
nand U18295 (N_18295,N_11130,N_10742);
or U18296 (N_18296,N_14245,N_11563);
nor U18297 (N_18297,N_14337,N_13207);
xor U18298 (N_18298,N_10578,N_13654);
and U18299 (N_18299,N_13507,N_13425);
xnor U18300 (N_18300,N_11514,N_10802);
nor U18301 (N_18301,N_14767,N_13448);
and U18302 (N_18302,N_12461,N_10953);
xor U18303 (N_18303,N_14470,N_11857);
xor U18304 (N_18304,N_14995,N_12738);
nor U18305 (N_18305,N_11919,N_11495);
and U18306 (N_18306,N_13250,N_12997);
nand U18307 (N_18307,N_11975,N_13594);
nor U18308 (N_18308,N_14966,N_10206);
nor U18309 (N_18309,N_14623,N_10748);
xor U18310 (N_18310,N_11609,N_11411);
xnor U18311 (N_18311,N_12055,N_12822);
and U18312 (N_18312,N_10886,N_14193);
nand U18313 (N_18313,N_14987,N_13593);
nor U18314 (N_18314,N_11280,N_14693);
xor U18315 (N_18315,N_14219,N_14954);
or U18316 (N_18316,N_10552,N_12714);
nand U18317 (N_18317,N_10274,N_10515);
xor U18318 (N_18318,N_10439,N_11888);
nand U18319 (N_18319,N_11876,N_10441);
nor U18320 (N_18320,N_13631,N_12587);
or U18321 (N_18321,N_12411,N_13465);
nor U18322 (N_18322,N_14119,N_14685);
nor U18323 (N_18323,N_10308,N_14649);
or U18324 (N_18324,N_13855,N_12708);
nor U18325 (N_18325,N_13721,N_13659);
xor U18326 (N_18326,N_12767,N_14976);
and U18327 (N_18327,N_13418,N_12112);
nand U18328 (N_18328,N_12091,N_11080);
and U18329 (N_18329,N_13859,N_14577);
and U18330 (N_18330,N_14683,N_11532);
nand U18331 (N_18331,N_14077,N_14909);
xor U18332 (N_18332,N_14454,N_11782);
or U18333 (N_18333,N_10925,N_12430);
and U18334 (N_18334,N_11023,N_14913);
and U18335 (N_18335,N_11110,N_10440);
or U18336 (N_18336,N_11576,N_11188);
and U18337 (N_18337,N_10931,N_13497);
or U18338 (N_18338,N_11238,N_11433);
nor U18339 (N_18339,N_11198,N_10884);
xor U18340 (N_18340,N_10275,N_10879);
xor U18341 (N_18341,N_11203,N_10996);
nor U18342 (N_18342,N_11728,N_14315);
and U18343 (N_18343,N_11946,N_12863);
nand U18344 (N_18344,N_14874,N_12145);
or U18345 (N_18345,N_13909,N_10732);
xor U18346 (N_18346,N_14440,N_12882);
or U18347 (N_18347,N_10057,N_10238);
or U18348 (N_18348,N_13453,N_14152);
or U18349 (N_18349,N_13674,N_12330);
nand U18350 (N_18350,N_10480,N_12679);
xnor U18351 (N_18351,N_13747,N_13402);
nand U18352 (N_18352,N_11847,N_11541);
and U18353 (N_18353,N_13980,N_14963);
and U18354 (N_18354,N_14680,N_11566);
and U18355 (N_18355,N_10861,N_14707);
nor U18356 (N_18356,N_12315,N_13744);
and U18357 (N_18357,N_14290,N_13195);
or U18358 (N_18358,N_14816,N_10216);
nor U18359 (N_18359,N_12942,N_14258);
nand U18360 (N_18360,N_14849,N_10092);
nand U18361 (N_18361,N_11591,N_14316);
or U18362 (N_18362,N_11087,N_10111);
nor U18363 (N_18363,N_12849,N_13354);
and U18364 (N_18364,N_10261,N_10268);
and U18365 (N_18365,N_12885,N_11586);
or U18366 (N_18366,N_12692,N_10792);
and U18367 (N_18367,N_12128,N_10388);
nand U18368 (N_18368,N_14200,N_11363);
and U18369 (N_18369,N_10016,N_10777);
and U18370 (N_18370,N_14684,N_11112);
nor U18371 (N_18371,N_12386,N_12334);
nor U18372 (N_18372,N_12088,N_10328);
or U18373 (N_18373,N_13588,N_12442);
nor U18374 (N_18374,N_13424,N_13817);
xor U18375 (N_18375,N_12124,N_14340);
nor U18376 (N_18376,N_13036,N_14720);
and U18377 (N_18377,N_11696,N_14088);
and U18378 (N_18378,N_14600,N_10855);
xor U18379 (N_18379,N_10629,N_10774);
or U18380 (N_18380,N_13161,N_11731);
nor U18381 (N_18381,N_12786,N_13069);
or U18382 (N_18382,N_12863,N_10917);
and U18383 (N_18383,N_11709,N_14654);
and U18384 (N_18384,N_14035,N_10664);
or U18385 (N_18385,N_10916,N_11657);
nor U18386 (N_18386,N_12657,N_12930);
xnor U18387 (N_18387,N_13676,N_10686);
nor U18388 (N_18388,N_11083,N_14576);
nand U18389 (N_18389,N_10831,N_12188);
or U18390 (N_18390,N_12959,N_14715);
nor U18391 (N_18391,N_13817,N_11143);
nand U18392 (N_18392,N_14057,N_12256);
or U18393 (N_18393,N_12081,N_14442);
and U18394 (N_18394,N_12296,N_12386);
nand U18395 (N_18395,N_14953,N_11171);
nand U18396 (N_18396,N_13597,N_14494);
nor U18397 (N_18397,N_14467,N_14282);
and U18398 (N_18398,N_12985,N_11815);
and U18399 (N_18399,N_13427,N_11986);
and U18400 (N_18400,N_12191,N_13196);
nor U18401 (N_18401,N_10900,N_13885);
xnor U18402 (N_18402,N_14273,N_11638);
and U18403 (N_18403,N_14811,N_11935);
and U18404 (N_18404,N_12690,N_12152);
and U18405 (N_18405,N_13749,N_10208);
or U18406 (N_18406,N_11588,N_14322);
or U18407 (N_18407,N_12474,N_10427);
nor U18408 (N_18408,N_10269,N_12752);
and U18409 (N_18409,N_13779,N_12753);
nand U18410 (N_18410,N_14282,N_12191);
or U18411 (N_18411,N_14769,N_11616);
nor U18412 (N_18412,N_11033,N_12013);
xor U18413 (N_18413,N_13701,N_13629);
nor U18414 (N_18414,N_12796,N_12450);
nor U18415 (N_18415,N_10757,N_13783);
xor U18416 (N_18416,N_14285,N_14182);
nor U18417 (N_18417,N_12555,N_14372);
or U18418 (N_18418,N_14861,N_13072);
nand U18419 (N_18419,N_12877,N_13654);
xor U18420 (N_18420,N_14867,N_11613);
nor U18421 (N_18421,N_14989,N_14876);
xor U18422 (N_18422,N_12103,N_11252);
nor U18423 (N_18423,N_14761,N_14564);
nand U18424 (N_18424,N_12291,N_12241);
and U18425 (N_18425,N_13013,N_10708);
or U18426 (N_18426,N_10600,N_14228);
nor U18427 (N_18427,N_12569,N_14492);
or U18428 (N_18428,N_11684,N_12218);
xnor U18429 (N_18429,N_10567,N_13738);
nor U18430 (N_18430,N_13771,N_10779);
nor U18431 (N_18431,N_12805,N_11838);
xor U18432 (N_18432,N_10175,N_12622);
and U18433 (N_18433,N_14655,N_14918);
nand U18434 (N_18434,N_12503,N_10545);
nor U18435 (N_18435,N_10145,N_14120);
nand U18436 (N_18436,N_12608,N_11336);
nand U18437 (N_18437,N_11892,N_14200);
nor U18438 (N_18438,N_14409,N_13401);
xor U18439 (N_18439,N_11867,N_10536);
nand U18440 (N_18440,N_10958,N_14463);
and U18441 (N_18441,N_13248,N_12022);
xor U18442 (N_18442,N_12524,N_14941);
and U18443 (N_18443,N_11813,N_12206);
nor U18444 (N_18444,N_14186,N_11889);
nor U18445 (N_18445,N_13351,N_14948);
or U18446 (N_18446,N_10969,N_12033);
nand U18447 (N_18447,N_13558,N_14616);
and U18448 (N_18448,N_12987,N_13689);
xnor U18449 (N_18449,N_13794,N_11786);
nand U18450 (N_18450,N_10624,N_14795);
and U18451 (N_18451,N_14824,N_14417);
or U18452 (N_18452,N_14996,N_13478);
nor U18453 (N_18453,N_10190,N_13961);
nand U18454 (N_18454,N_13996,N_11923);
xnor U18455 (N_18455,N_10065,N_14060);
and U18456 (N_18456,N_13090,N_11302);
xor U18457 (N_18457,N_12153,N_13028);
or U18458 (N_18458,N_14181,N_10581);
nor U18459 (N_18459,N_13015,N_14863);
xnor U18460 (N_18460,N_10521,N_10742);
and U18461 (N_18461,N_11778,N_13349);
and U18462 (N_18462,N_11671,N_10113);
nor U18463 (N_18463,N_10832,N_13900);
or U18464 (N_18464,N_12184,N_12762);
nand U18465 (N_18465,N_13736,N_14103);
or U18466 (N_18466,N_12180,N_13378);
xnor U18467 (N_18467,N_11834,N_14168);
and U18468 (N_18468,N_11478,N_10735);
or U18469 (N_18469,N_13358,N_12188);
nor U18470 (N_18470,N_12470,N_11646);
or U18471 (N_18471,N_14044,N_14121);
nand U18472 (N_18472,N_10444,N_12450);
nand U18473 (N_18473,N_10727,N_14160);
xnor U18474 (N_18474,N_10446,N_11484);
xnor U18475 (N_18475,N_13589,N_11351);
or U18476 (N_18476,N_14865,N_14365);
or U18477 (N_18477,N_14217,N_11207);
or U18478 (N_18478,N_12543,N_14171);
and U18479 (N_18479,N_14631,N_11030);
and U18480 (N_18480,N_10689,N_10496);
nand U18481 (N_18481,N_10345,N_12173);
nand U18482 (N_18482,N_14499,N_11509);
nor U18483 (N_18483,N_12174,N_13976);
nor U18484 (N_18484,N_12342,N_10858);
xor U18485 (N_18485,N_14097,N_10626);
nand U18486 (N_18486,N_12690,N_14605);
xor U18487 (N_18487,N_11156,N_10519);
xor U18488 (N_18488,N_13236,N_10825);
and U18489 (N_18489,N_13933,N_12814);
nor U18490 (N_18490,N_11736,N_11795);
xor U18491 (N_18491,N_13447,N_14177);
nor U18492 (N_18492,N_11981,N_13976);
nor U18493 (N_18493,N_11677,N_12814);
and U18494 (N_18494,N_10065,N_14855);
xor U18495 (N_18495,N_13134,N_13870);
nand U18496 (N_18496,N_10503,N_11991);
and U18497 (N_18497,N_11993,N_14306);
nor U18498 (N_18498,N_10629,N_12475);
and U18499 (N_18499,N_10871,N_10653);
nor U18500 (N_18500,N_10533,N_11887);
nand U18501 (N_18501,N_13434,N_11085);
nor U18502 (N_18502,N_14477,N_12600);
nand U18503 (N_18503,N_13903,N_10209);
xnor U18504 (N_18504,N_10360,N_13807);
and U18505 (N_18505,N_11185,N_12810);
and U18506 (N_18506,N_10805,N_13370);
nor U18507 (N_18507,N_11296,N_13365);
nor U18508 (N_18508,N_10735,N_12037);
nand U18509 (N_18509,N_13399,N_14017);
xor U18510 (N_18510,N_10798,N_11461);
nand U18511 (N_18511,N_12663,N_13142);
xor U18512 (N_18512,N_12226,N_10080);
nor U18513 (N_18513,N_11950,N_14371);
or U18514 (N_18514,N_11108,N_11636);
and U18515 (N_18515,N_11112,N_12037);
nor U18516 (N_18516,N_13532,N_13673);
xor U18517 (N_18517,N_11820,N_11392);
or U18518 (N_18518,N_13906,N_12102);
nand U18519 (N_18519,N_10930,N_13621);
nor U18520 (N_18520,N_13465,N_14357);
xor U18521 (N_18521,N_13387,N_10555);
xor U18522 (N_18522,N_13419,N_14028);
xor U18523 (N_18523,N_14262,N_10352);
or U18524 (N_18524,N_14306,N_12417);
or U18525 (N_18525,N_12217,N_12480);
nor U18526 (N_18526,N_14050,N_10696);
or U18527 (N_18527,N_14469,N_13707);
nand U18528 (N_18528,N_13463,N_13936);
nor U18529 (N_18529,N_12784,N_13971);
nand U18530 (N_18530,N_12739,N_10371);
xnor U18531 (N_18531,N_10266,N_13518);
nand U18532 (N_18532,N_10268,N_10755);
and U18533 (N_18533,N_12184,N_11185);
or U18534 (N_18534,N_11185,N_11532);
or U18535 (N_18535,N_13433,N_12352);
xor U18536 (N_18536,N_14511,N_10572);
and U18537 (N_18537,N_11745,N_13907);
nand U18538 (N_18538,N_10952,N_13370);
nand U18539 (N_18539,N_10339,N_10988);
and U18540 (N_18540,N_10308,N_14663);
or U18541 (N_18541,N_12219,N_12385);
xor U18542 (N_18542,N_12609,N_10488);
nor U18543 (N_18543,N_10137,N_12690);
or U18544 (N_18544,N_13772,N_12903);
or U18545 (N_18545,N_11982,N_12915);
and U18546 (N_18546,N_10951,N_14041);
or U18547 (N_18547,N_14780,N_12857);
and U18548 (N_18548,N_14415,N_14628);
nand U18549 (N_18549,N_12139,N_14911);
xor U18550 (N_18550,N_10612,N_11688);
xor U18551 (N_18551,N_12669,N_14220);
nor U18552 (N_18552,N_12204,N_12577);
nor U18553 (N_18553,N_14200,N_14723);
xor U18554 (N_18554,N_10544,N_13444);
nand U18555 (N_18555,N_10686,N_14970);
nor U18556 (N_18556,N_11406,N_13157);
nor U18557 (N_18557,N_14272,N_14690);
or U18558 (N_18558,N_10032,N_14168);
and U18559 (N_18559,N_13675,N_10085);
or U18560 (N_18560,N_13466,N_11493);
nor U18561 (N_18561,N_14903,N_14775);
or U18562 (N_18562,N_14085,N_11385);
or U18563 (N_18563,N_14708,N_13157);
nand U18564 (N_18564,N_10715,N_14016);
xor U18565 (N_18565,N_10097,N_11395);
nand U18566 (N_18566,N_10780,N_13408);
nor U18567 (N_18567,N_12442,N_10373);
or U18568 (N_18568,N_12488,N_11721);
nand U18569 (N_18569,N_13511,N_12948);
and U18570 (N_18570,N_10971,N_13539);
nand U18571 (N_18571,N_11009,N_14770);
and U18572 (N_18572,N_11088,N_12025);
nand U18573 (N_18573,N_11542,N_12325);
nand U18574 (N_18574,N_13826,N_12081);
nor U18575 (N_18575,N_10627,N_13821);
nor U18576 (N_18576,N_13560,N_10646);
nor U18577 (N_18577,N_11123,N_13229);
or U18578 (N_18578,N_10944,N_13344);
nor U18579 (N_18579,N_10262,N_11017);
nand U18580 (N_18580,N_13612,N_11124);
nor U18581 (N_18581,N_13558,N_11372);
xor U18582 (N_18582,N_10579,N_10819);
xnor U18583 (N_18583,N_14705,N_12870);
and U18584 (N_18584,N_13431,N_14430);
nor U18585 (N_18585,N_10942,N_12703);
and U18586 (N_18586,N_11880,N_13903);
or U18587 (N_18587,N_10064,N_11190);
and U18588 (N_18588,N_13739,N_11033);
nor U18589 (N_18589,N_12027,N_13933);
or U18590 (N_18590,N_10886,N_11090);
nand U18591 (N_18591,N_14354,N_14260);
xnor U18592 (N_18592,N_14240,N_12913);
nand U18593 (N_18593,N_11928,N_13228);
xnor U18594 (N_18594,N_11302,N_11896);
nand U18595 (N_18595,N_11707,N_10952);
and U18596 (N_18596,N_14293,N_14675);
and U18597 (N_18597,N_10479,N_13761);
nand U18598 (N_18598,N_12029,N_10393);
nor U18599 (N_18599,N_14401,N_11596);
nor U18600 (N_18600,N_11564,N_13071);
nor U18601 (N_18601,N_11232,N_10382);
xor U18602 (N_18602,N_13682,N_14633);
nand U18603 (N_18603,N_12726,N_14403);
xnor U18604 (N_18604,N_11834,N_12448);
or U18605 (N_18605,N_10012,N_10948);
and U18606 (N_18606,N_14156,N_10402);
xor U18607 (N_18607,N_10840,N_11873);
nand U18608 (N_18608,N_11207,N_11784);
nand U18609 (N_18609,N_10954,N_10520);
nor U18610 (N_18610,N_12142,N_11534);
nor U18611 (N_18611,N_10234,N_10780);
or U18612 (N_18612,N_14765,N_10562);
nor U18613 (N_18613,N_11808,N_11805);
and U18614 (N_18614,N_14409,N_12148);
or U18615 (N_18615,N_11465,N_14717);
nor U18616 (N_18616,N_11899,N_10376);
xnor U18617 (N_18617,N_13026,N_11989);
xnor U18618 (N_18618,N_11798,N_10823);
or U18619 (N_18619,N_14604,N_11693);
and U18620 (N_18620,N_10475,N_13178);
nand U18621 (N_18621,N_11103,N_10091);
or U18622 (N_18622,N_11231,N_12145);
xnor U18623 (N_18623,N_11042,N_13404);
or U18624 (N_18624,N_10139,N_10615);
and U18625 (N_18625,N_13594,N_14801);
nor U18626 (N_18626,N_13751,N_11846);
or U18627 (N_18627,N_13195,N_14692);
and U18628 (N_18628,N_13191,N_11064);
and U18629 (N_18629,N_13007,N_13771);
or U18630 (N_18630,N_11989,N_10515);
and U18631 (N_18631,N_14232,N_12229);
nand U18632 (N_18632,N_12715,N_14516);
nand U18633 (N_18633,N_10345,N_14442);
and U18634 (N_18634,N_10402,N_13977);
nor U18635 (N_18635,N_11702,N_11442);
nor U18636 (N_18636,N_11668,N_11330);
or U18637 (N_18637,N_14680,N_12566);
and U18638 (N_18638,N_14099,N_13992);
and U18639 (N_18639,N_12375,N_10439);
xor U18640 (N_18640,N_14813,N_12205);
nand U18641 (N_18641,N_10882,N_14695);
or U18642 (N_18642,N_10980,N_11768);
nor U18643 (N_18643,N_14551,N_13009);
and U18644 (N_18644,N_11722,N_12868);
and U18645 (N_18645,N_12509,N_13966);
and U18646 (N_18646,N_12038,N_10214);
and U18647 (N_18647,N_12560,N_13891);
or U18648 (N_18648,N_14612,N_12572);
nand U18649 (N_18649,N_11877,N_11513);
and U18650 (N_18650,N_12288,N_10540);
nand U18651 (N_18651,N_13688,N_11304);
or U18652 (N_18652,N_10658,N_14166);
xnor U18653 (N_18653,N_14815,N_10758);
and U18654 (N_18654,N_11828,N_13175);
and U18655 (N_18655,N_10808,N_13204);
and U18656 (N_18656,N_14262,N_13506);
nand U18657 (N_18657,N_10756,N_12346);
and U18658 (N_18658,N_13949,N_11066);
or U18659 (N_18659,N_10275,N_11363);
or U18660 (N_18660,N_12521,N_12196);
nor U18661 (N_18661,N_10229,N_11841);
nand U18662 (N_18662,N_10686,N_10890);
and U18663 (N_18663,N_14326,N_13448);
and U18664 (N_18664,N_12110,N_13839);
nor U18665 (N_18665,N_11064,N_12537);
and U18666 (N_18666,N_11438,N_11108);
nor U18667 (N_18667,N_13559,N_12975);
xnor U18668 (N_18668,N_12235,N_10871);
and U18669 (N_18669,N_14440,N_10058);
nand U18670 (N_18670,N_10977,N_10422);
or U18671 (N_18671,N_11520,N_12124);
nand U18672 (N_18672,N_10593,N_12463);
xor U18673 (N_18673,N_13493,N_11914);
nor U18674 (N_18674,N_11045,N_12493);
nor U18675 (N_18675,N_11142,N_10058);
nor U18676 (N_18676,N_11797,N_12164);
or U18677 (N_18677,N_14529,N_10791);
nor U18678 (N_18678,N_11622,N_10492);
nand U18679 (N_18679,N_14353,N_12821);
nand U18680 (N_18680,N_11605,N_12870);
nand U18681 (N_18681,N_12491,N_12077);
and U18682 (N_18682,N_11468,N_13561);
nor U18683 (N_18683,N_13907,N_12985);
nor U18684 (N_18684,N_12968,N_12863);
nor U18685 (N_18685,N_13541,N_12166);
xnor U18686 (N_18686,N_13881,N_12806);
xnor U18687 (N_18687,N_10259,N_11282);
xor U18688 (N_18688,N_14578,N_13481);
nor U18689 (N_18689,N_11348,N_14112);
and U18690 (N_18690,N_14249,N_11255);
nor U18691 (N_18691,N_10319,N_13253);
or U18692 (N_18692,N_12430,N_10369);
nor U18693 (N_18693,N_14058,N_11399);
nand U18694 (N_18694,N_14869,N_13966);
nand U18695 (N_18695,N_11955,N_12474);
nor U18696 (N_18696,N_13406,N_10300);
nand U18697 (N_18697,N_10489,N_10577);
or U18698 (N_18698,N_10872,N_13909);
nand U18699 (N_18699,N_11237,N_12226);
nand U18700 (N_18700,N_14286,N_12474);
or U18701 (N_18701,N_13438,N_10442);
and U18702 (N_18702,N_11133,N_14802);
and U18703 (N_18703,N_13287,N_14840);
xor U18704 (N_18704,N_14291,N_12988);
and U18705 (N_18705,N_11285,N_14155);
and U18706 (N_18706,N_14896,N_10616);
or U18707 (N_18707,N_14243,N_14596);
and U18708 (N_18708,N_11250,N_14622);
or U18709 (N_18709,N_12719,N_12804);
xor U18710 (N_18710,N_13130,N_11704);
nor U18711 (N_18711,N_13140,N_12885);
or U18712 (N_18712,N_14641,N_12015);
and U18713 (N_18713,N_10938,N_12928);
nor U18714 (N_18714,N_11496,N_11845);
xnor U18715 (N_18715,N_11173,N_13568);
or U18716 (N_18716,N_14942,N_12990);
xnor U18717 (N_18717,N_12417,N_13982);
or U18718 (N_18718,N_12220,N_11775);
and U18719 (N_18719,N_13201,N_13067);
nor U18720 (N_18720,N_12616,N_14484);
or U18721 (N_18721,N_12759,N_12212);
nor U18722 (N_18722,N_11980,N_13121);
or U18723 (N_18723,N_14113,N_11726);
xor U18724 (N_18724,N_11890,N_12972);
or U18725 (N_18725,N_13765,N_14316);
nand U18726 (N_18726,N_13668,N_14321);
and U18727 (N_18727,N_14768,N_11989);
xnor U18728 (N_18728,N_13001,N_11327);
and U18729 (N_18729,N_10948,N_12046);
nand U18730 (N_18730,N_10442,N_12421);
or U18731 (N_18731,N_14228,N_11440);
or U18732 (N_18732,N_12039,N_12960);
or U18733 (N_18733,N_14739,N_10562);
nor U18734 (N_18734,N_12664,N_12998);
and U18735 (N_18735,N_11305,N_12254);
nor U18736 (N_18736,N_14958,N_14652);
xnor U18737 (N_18737,N_13028,N_10415);
xnor U18738 (N_18738,N_10988,N_13503);
or U18739 (N_18739,N_13513,N_13637);
or U18740 (N_18740,N_13000,N_10620);
nand U18741 (N_18741,N_12502,N_13612);
xnor U18742 (N_18742,N_13594,N_14025);
and U18743 (N_18743,N_13327,N_11699);
or U18744 (N_18744,N_14626,N_10781);
and U18745 (N_18745,N_14028,N_11064);
and U18746 (N_18746,N_14352,N_14199);
xor U18747 (N_18747,N_11506,N_10892);
xnor U18748 (N_18748,N_13113,N_10589);
xor U18749 (N_18749,N_11810,N_13870);
nand U18750 (N_18750,N_12709,N_11384);
or U18751 (N_18751,N_14700,N_11073);
and U18752 (N_18752,N_14300,N_14880);
or U18753 (N_18753,N_11992,N_12066);
xnor U18754 (N_18754,N_11270,N_12502);
or U18755 (N_18755,N_12306,N_10148);
nor U18756 (N_18756,N_10677,N_14729);
nor U18757 (N_18757,N_12877,N_12710);
or U18758 (N_18758,N_10360,N_12172);
nand U18759 (N_18759,N_13006,N_11298);
xnor U18760 (N_18760,N_12726,N_14135);
xor U18761 (N_18761,N_14918,N_13955);
xor U18762 (N_18762,N_13982,N_10264);
and U18763 (N_18763,N_10153,N_14044);
nand U18764 (N_18764,N_12736,N_12489);
and U18765 (N_18765,N_11370,N_11344);
or U18766 (N_18766,N_13259,N_12187);
nor U18767 (N_18767,N_12624,N_10748);
xnor U18768 (N_18768,N_11031,N_10418);
and U18769 (N_18769,N_11239,N_11369);
xor U18770 (N_18770,N_14810,N_12693);
xor U18771 (N_18771,N_13683,N_10584);
and U18772 (N_18772,N_10241,N_14997);
or U18773 (N_18773,N_13372,N_13924);
and U18774 (N_18774,N_13024,N_12556);
xnor U18775 (N_18775,N_10655,N_10241);
and U18776 (N_18776,N_10566,N_10767);
nand U18777 (N_18777,N_10553,N_14709);
xor U18778 (N_18778,N_11446,N_11560);
nor U18779 (N_18779,N_13420,N_14358);
nor U18780 (N_18780,N_14638,N_11920);
xnor U18781 (N_18781,N_10097,N_14123);
xor U18782 (N_18782,N_14507,N_14991);
and U18783 (N_18783,N_14790,N_10657);
nand U18784 (N_18784,N_13148,N_14970);
nor U18785 (N_18785,N_14531,N_13704);
xor U18786 (N_18786,N_13723,N_11534);
or U18787 (N_18787,N_14694,N_11891);
xnor U18788 (N_18788,N_11642,N_14883);
and U18789 (N_18789,N_11930,N_13013);
or U18790 (N_18790,N_12449,N_14830);
and U18791 (N_18791,N_11328,N_13577);
nand U18792 (N_18792,N_10722,N_12045);
or U18793 (N_18793,N_13085,N_10325);
or U18794 (N_18794,N_10321,N_14324);
and U18795 (N_18795,N_11380,N_12146);
xor U18796 (N_18796,N_14480,N_13388);
xnor U18797 (N_18797,N_14718,N_11841);
xor U18798 (N_18798,N_11042,N_13625);
or U18799 (N_18799,N_13846,N_14874);
nand U18800 (N_18800,N_10514,N_13387);
xor U18801 (N_18801,N_14421,N_12727);
or U18802 (N_18802,N_14405,N_13432);
nand U18803 (N_18803,N_12243,N_14157);
or U18804 (N_18804,N_11218,N_12520);
xor U18805 (N_18805,N_10843,N_10782);
or U18806 (N_18806,N_13372,N_13088);
nand U18807 (N_18807,N_11333,N_11866);
and U18808 (N_18808,N_11054,N_13257);
and U18809 (N_18809,N_14363,N_10393);
nand U18810 (N_18810,N_12760,N_10858);
nor U18811 (N_18811,N_10510,N_11371);
nor U18812 (N_18812,N_11485,N_13926);
nor U18813 (N_18813,N_12617,N_11739);
nand U18814 (N_18814,N_14271,N_10988);
nand U18815 (N_18815,N_10454,N_13510);
nand U18816 (N_18816,N_13840,N_11322);
xnor U18817 (N_18817,N_14498,N_10474);
xnor U18818 (N_18818,N_10093,N_10294);
xor U18819 (N_18819,N_11207,N_12237);
xor U18820 (N_18820,N_10546,N_10595);
nor U18821 (N_18821,N_12079,N_12027);
nand U18822 (N_18822,N_13677,N_10728);
nor U18823 (N_18823,N_10668,N_11800);
or U18824 (N_18824,N_11546,N_11824);
nand U18825 (N_18825,N_12250,N_14862);
nor U18826 (N_18826,N_14392,N_13790);
xor U18827 (N_18827,N_10562,N_10640);
or U18828 (N_18828,N_14114,N_11227);
nor U18829 (N_18829,N_12867,N_12952);
xnor U18830 (N_18830,N_12530,N_10720);
nand U18831 (N_18831,N_11796,N_13558);
or U18832 (N_18832,N_14521,N_11036);
nand U18833 (N_18833,N_14108,N_13894);
and U18834 (N_18834,N_12412,N_13318);
or U18835 (N_18835,N_12711,N_12266);
and U18836 (N_18836,N_14365,N_12662);
and U18837 (N_18837,N_14254,N_11120);
or U18838 (N_18838,N_13953,N_11922);
nor U18839 (N_18839,N_11253,N_14174);
xnor U18840 (N_18840,N_10748,N_11577);
nand U18841 (N_18841,N_10375,N_11984);
nand U18842 (N_18842,N_11757,N_10362);
nor U18843 (N_18843,N_11281,N_13581);
nand U18844 (N_18844,N_11295,N_14802);
nor U18845 (N_18845,N_14761,N_11840);
or U18846 (N_18846,N_14477,N_14428);
nand U18847 (N_18847,N_11058,N_10010);
and U18848 (N_18848,N_12543,N_11280);
nand U18849 (N_18849,N_13173,N_13683);
nor U18850 (N_18850,N_12843,N_12727);
or U18851 (N_18851,N_14639,N_14440);
and U18852 (N_18852,N_13447,N_10773);
or U18853 (N_18853,N_11485,N_14829);
nor U18854 (N_18854,N_13456,N_11915);
or U18855 (N_18855,N_11417,N_14949);
nand U18856 (N_18856,N_11424,N_12176);
nor U18857 (N_18857,N_13824,N_13469);
xnor U18858 (N_18858,N_11904,N_12752);
and U18859 (N_18859,N_10651,N_11190);
nand U18860 (N_18860,N_11558,N_14645);
and U18861 (N_18861,N_11612,N_10001);
and U18862 (N_18862,N_13802,N_10917);
and U18863 (N_18863,N_13939,N_11918);
nand U18864 (N_18864,N_13999,N_13085);
or U18865 (N_18865,N_13320,N_14557);
xor U18866 (N_18866,N_12942,N_11228);
and U18867 (N_18867,N_11498,N_10553);
nand U18868 (N_18868,N_14522,N_12570);
and U18869 (N_18869,N_11665,N_14872);
or U18870 (N_18870,N_13571,N_10347);
or U18871 (N_18871,N_11690,N_13768);
and U18872 (N_18872,N_11906,N_10745);
nand U18873 (N_18873,N_10908,N_14020);
and U18874 (N_18874,N_11952,N_12321);
or U18875 (N_18875,N_11508,N_14397);
or U18876 (N_18876,N_14930,N_10695);
nand U18877 (N_18877,N_11186,N_12739);
and U18878 (N_18878,N_14398,N_10800);
or U18879 (N_18879,N_12223,N_10956);
or U18880 (N_18880,N_12851,N_10466);
or U18881 (N_18881,N_10670,N_12795);
xnor U18882 (N_18882,N_13757,N_13810);
nand U18883 (N_18883,N_12420,N_11371);
xor U18884 (N_18884,N_14753,N_10924);
nand U18885 (N_18885,N_13404,N_13373);
xnor U18886 (N_18886,N_13003,N_11621);
or U18887 (N_18887,N_11506,N_12037);
or U18888 (N_18888,N_11896,N_13831);
or U18889 (N_18889,N_10602,N_13650);
nand U18890 (N_18890,N_14097,N_13109);
nand U18891 (N_18891,N_11336,N_14299);
nand U18892 (N_18892,N_13132,N_11782);
xnor U18893 (N_18893,N_13001,N_14867);
nor U18894 (N_18894,N_10056,N_12477);
and U18895 (N_18895,N_13281,N_14785);
or U18896 (N_18896,N_10279,N_14018);
and U18897 (N_18897,N_13917,N_13447);
and U18898 (N_18898,N_12958,N_12247);
nor U18899 (N_18899,N_12711,N_14783);
and U18900 (N_18900,N_10852,N_10257);
nor U18901 (N_18901,N_10085,N_11331);
nor U18902 (N_18902,N_10201,N_13261);
xnor U18903 (N_18903,N_13783,N_12058);
xnor U18904 (N_18904,N_11591,N_10586);
nand U18905 (N_18905,N_11482,N_13085);
nand U18906 (N_18906,N_11536,N_10708);
or U18907 (N_18907,N_12391,N_10087);
nand U18908 (N_18908,N_12448,N_13188);
or U18909 (N_18909,N_11548,N_11291);
nand U18910 (N_18910,N_10383,N_13904);
xnor U18911 (N_18911,N_11094,N_14052);
nor U18912 (N_18912,N_14513,N_14629);
xor U18913 (N_18913,N_11622,N_13299);
nand U18914 (N_18914,N_10322,N_13489);
nand U18915 (N_18915,N_11768,N_13888);
nand U18916 (N_18916,N_10917,N_11581);
nand U18917 (N_18917,N_14596,N_10059);
nand U18918 (N_18918,N_14037,N_11434);
or U18919 (N_18919,N_12775,N_12185);
and U18920 (N_18920,N_11808,N_14865);
xnor U18921 (N_18921,N_13990,N_12302);
xor U18922 (N_18922,N_11582,N_12363);
xnor U18923 (N_18923,N_13928,N_14600);
nand U18924 (N_18924,N_10144,N_12805);
or U18925 (N_18925,N_12250,N_11611);
xnor U18926 (N_18926,N_13973,N_13526);
and U18927 (N_18927,N_11948,N_13378);
xor U18928 (N_18928,N_14706,N_11296);
xor U18929 (N_18929,N_14984,N_13646);
or U18930 (N_18930,N_13344,N_14827);
xor U18931 (N_18931,N_10951,N_13420);
or U18932 (N_18932,N_11455,N_10250);
nand U18933 (N_18933,N_12944,N_11730);
nor U18934 (N_18934,N_10622,N_10956);
or U18935 (N_18935,N_13492,N_13764);
or U18936 (N_18936,N_10265,N_14864);
or U18937 (N_18937,N_13541,N_10776);
and U18938 (N_18938,N_12841,N_12612);
xnor U18939 (N_18939,N_14043,N_11821);
or U18940 (N_18940,N_11493,N_14822);
xnor U18941 (N_18941,N_13513,N_13362);
or U18942 (N_18942,N_11970,N_12737);
nand U18943 (N_18943,N_13173,N_13665);
nor U18944 (N_18944,N_12894,N_11633);
xnor U18945 (N_18945,N_13114,N_10195);
nor U18946 (N_18946,N_12475,N_12826);
nor U18947 (N_18947,N_14114,N_12391);
nor U18948 (N_18948,N_14368,N_12063);
nor U18949 (N_18949,N_14804,N_14954);
and U18950 (N_18950,N_11200,N_10855);
nor U18951 (N_18951,N_13685,N_10185);
nand U18952 (N_18952,N_14470,N_10791);
or U18953 (N_18953,N_12787,N_10425);
nor U18954 (N_18954,N_12278,N_14628);
nor U18955 (N_18955,N_12209,N_11083);
xnor U18956 (N_18956,N_13044,N_11156);
nor U18957 (N_18957,N_10597,N_14114);
and U18958 (N_18958,N_11299,N_10543);
nor U18959 (N_18959,N_14596,N_12360);
xnor U18960 (N_18960,N_11761,N_10355);
nor U18961 (N_18961,N_11892,N_13843);
and U18962 (N_18962,N_10416,N_12381);
nor U18963 (N_18963,N_13945,N_10750);
and U18964 (N_18964,N_12191,N_12024);
or U18965 (N_18965,N_13939,N_12249);
and U18966 (N_18966,N_11217,N_13270);
xor U18967 (N_18967,N_13771,N_12834);
nor U18968 (N_18968,N_12777,N_14057);
or U18969 (N_18969,N_10371,N_12500);
nor U18970 (N_18970,N_10166,N_14704);
xor U18971 (N_18971,N_11941,N_14415);
xnor U18972 (N_18972,N_14619,N_11576);
or U18973 (N_18973,N_14949,N_11507);
nor U18974 (N_18974,N_13788,N_12938);
and U18975 (N_18975,N_14807,N_10772);
nor U18976 (N_18976,N_14615,N_14366);
nand U18977 (N_18977,N_13163,N_10670);
and U18978 (N_18978,N_14971,N_14646);
nand U18979 (N_18979,N_11154,N_14031);
nor U18980 (N_18980,N_11385,N_11511);
or U18981 (N_18981,N_14330,N_14339);
nor U18982 (N_18982,N_12235,N_12339);
nor U18983 (N_18983,N_13332,N_14439);
nor U18984 (N_18984,N_10791,N_12094);
and U18985 (N_18985,N_12897,N_14556);
nand U18986 (N_18986,N_11088,N_14233);
nor U18987 (N_18987,N_12913,N_13989);
and U18988 (N_18988,N_10485,N_11224);
nand U18989 (N_18989,N_12976,N_14164);
or U18990 (N_18990,N_12230,N_11694);
nor U18991 (N_18991,N_12116,N_14117);
and U18992 (N_18992,N_12726,N_13874);
or U18993 (N_18993,N_14623,N_10152);
or U18994 (N_18994,N_13425,N_14142);
xor U18995 (N_18995,N_12226,N_13764);
and U18996 (N_18996,N_11630,N_13157);
nor U18997 (N_18997,N_10861,N_10068);
and U18998 (N_18998,N_14204,N_11794);
xnor U18999 (N_18999,N_12748,N_12171);
xor U19000 (N_19000,N_13822,N_13977);
or U19001 (N_19001,N_14283,N_14147);
xor U19002 (N_19002,N_14163,N_11695);
or U19003 (N_19003,N_12487,N_11016);
nor U19004 (N_19004,N_14938,N_11371);
nor U19005 (N_19005,N_13478,N_10975);
nand U19006 (N_19006,N_11712,N_12421);
or U19007 (N_19007,N_12708,N_12951);
or U19008 (N_19008,N_11225,N_13376);
and U19009 (N_19009,N_13621,N_13854);
or U19010 (N_19010,N_11061,N_10833);
or U19011 (N_19011,N_10328,N_11278);
xor U19012 (N_19012,N_11065,N_10808);
nor U19013 (N_19013,N_11205,N_10330);
and U19014 (N_19014,N_12005,N_14658);
or U19015 (N_19015,N_12034,N_14163);
nand U19016 (N_19016,N_10406,N_13347);
xnor U19017 (N_19017,N_13284,N_11847);
and U19018 (N_19018,N_11586,N_12165);
nor U19019 (N_19019,N_11401,N_12055);
xnor U19020 (N_19020,N_12502,N_14876);
nor U19021 (N_19021,N_13384,N_10225);
and U19022 (N_19022,N_11626,N_10553);
nand U19023 (N_19023,N_10322,N_11071);
xor U19024 (N_19024,N_13495,N_10960);
nand U19025 (N_19025,N_12118,N_13815);
nand U19026 (N_19026,N_12504,N_12604);
or U19027 (N_19027,N_11114,N_14981);
nand U19028 (N_19028,N_13277,N_11716);
and U19029 (N_19029,N_10131,N_14299);
nor U19030 (N_19030,N_11030,N_10648);
xor U19031 (N_19031,N_14840,N_10792);
nor U19032 (N_19032,N_11584,N_10361);
xnor U19033 (N_19033,N_13610,N_13738);
nor U19034 (N_19034,N_10356,N_11581);
and U19035 (N_19035,N_14117,N_11211);
or U19036 (N_19036,N_13631,N_13575);
xor U19037 (N_19037,N_14159,N_13468);
xor U19038 (N_19038,N_14701,N_12871);
nor U19039 (N_19039,N_13877,N_13814);
xor U19040 (N_19040,N_11329,N_12572);
or U19041 (N_19041,N_13520,N_11165);
nor U19042 (N_19042,N_12039,N_13290);
nand U19043 (N_19043,N_10592,N_14403);
or U19044 (N_19044,N_14943,N_11428);
nand U19045 (N_19045,N_13887,N_12178);
nor U19046 (N_19046,N_11501,N_13634);
xnor U19047 (N_19047,N_12877,N_14864);
nor U19048 (N_19048,N_11082,N_12985);
or U19049 (N_19049,N_14272,N_13698);
xor U19050 (N_19050,N_11152,N_13781);
nor U19051 (N_19051,N_12850,N_14612);
xor U19052 (N_19052,N_10349,N_10001);
or U19053 (N_19053,N_10039,N_10112);
nor U19054 (N_19054,N_14431,N_12511);
nor U19055 (N_19055,N_12507,N_12720);
nand U19056 (N_19056,N_13862,N_11686);
or U19057 (N_19057,N_13618,N_14179);
nor U19058 (N_19058,N_11401,N_10661);
or U19059 (N_19059,N_13934,N_11561);
and U19060 (N_19060,N_12343,N_10258);
or U19061 (N_19061,N_12468,N_13669);
or U19062 (N_19062,N_11395,N_12814);
and U19063 (N_19063,N_11949,N_12453);
or U19064 (N_19064,N_14145,N_10911);
or U19065 (N_19065,N_14156,N_13773);
nand U19066 (N_19066,N_13578,N_10421);
and U19067 (N_19067,N_11688,N_14110);
nand U19068 (N_19068,N_13493,N_13473);
and U19069 (N_19069,N_10280,N_11153);
nand U19070 (N_19070,N_11228,N_14865);
nand U19071 (N_19071,N_12195,N_12321);
nor U19072 (N_19072,N_12309,N_10879);
xor U19073 (N_19073,N_13646,N_14051);
nand U19074 (N_19074,N_10285,N_14889);
xor U19075 (N_19075,N_10170,N_13206);
nand U19076 (N_19076,N_10100,N_12380);
xor U19077 (N_19077,N_13390,N_12145);
or U19078 (N_19078,N_11487,N_12764);
xnor U19079 (N_19079,N_10680,N_11115);
and U19080 (N_19080,N_12394,N_11033);
xnor U19081 (N_19081,N_11739,N_14095);
nor U19082 (N_19082,N_11656,N_14740);
and U19083 (N_19083,N_13444,N_11409);
and U19084 (N_19084,N_13581,N_11879);
and U19085 (N_19085,N_10860,N_10852);
and U19086 (N_19086,N_13880,N_11897);
or U19087 (N_19087,N_14266,N_11969);
or U19088 (N_19088,N_13049,N_12741);
nand U19089 (N_19089,N_12727,N_12045);
nor U19090 (N_19090,N_11719,N_12029);
and U19091 (N_19091,N_12538,N_10750);
xnor U19092 (N_19092,N_13305,N_14483);
nor U19093 (N_19093,N_10303,N_13596);
or U19094 (N_19094,N_14547,N_13926);
nor U19095 (N_19095,N_14090,N_10541);
nand U19096 (N_19096,N_12478,N_14652);
and U19097 (N_19097,N_10004,N_14768);
and U19098 (N_19098,N_11971,N_10342);
and U19099 (N_19099,N_10349,N_11071);
or U19100 (N_19100,N_11249,N_14909);
nor U19101 (N_19101,N_10518,N_12840);
and U19102 (N_19102,N_12544,N_14438);
and U19103 (N_19103,N_11716,N_11132);
nor U19104 (N_19104,N_11029,N_10474);
or U19105 (N_19105,N_14171,N_10209);
and U19106 (N_19106,N_13685,N_10794);
nor U19107 (N_19107,N_13345,N_13434);
nor U19108 (N_19108,N_12618,N_12772);
nor U19109 (N_19109,N_14452,N_13710);
and U19110 (N_19110,N_13069,N_13119);
nor U19111 (N_19111,N_10946,N_14122);
nand U19112 (N_19112,N_11229,N_14234);
and U19113 (N_19113,N_13049,N_11570);
nor U19114 (N_19114,N_10681,N_13549);
xor U19115 (N_19115,N_13468,N_12929);
and U19116 (N_19116,N_11479,N_13449);
and U19117 (N_19117,N_13541,N_10055);
or U19118 (N_19118,N_14988,N_11130);
or U19119 (N_19119,N_12504,N_14965);
or U19120 (N_19120,N_13431,N_12043);
nand U19121 (N_19121,N_14900,N_12219);
or U19122 (N_19122,N_12135,N_10629);
xnor U19123 (N_19123,N_12041,N_14048);
xnor U19124 (N_19124,N_13127,N_14392);
and U19125 (N_19125,N_10796,N_11575);
xor U19126 (N_19126,N_11342,N_13162);
and U19127 (N_19127,N_13326,N_13729);
and U19128 (N_19128,N_14475,N_13823);
nand U19129 (N_19129,N_12706,N_11071);
nor U19130 (N_19130,N_13209,N_10238);
nand U19131 (N_19131,N_10709,N_11268);
nand U19132 (N_19132,N_12897,N_14645);
xor U19133 (N_19133,N_12324,N_10124);
and U19134 (N_19134,N_12680,N_12160);
xor U19135 (N_19135,N_13154,N_12345);
and U19136 (N_19136,N_13290,N_13024);
xor U19137 (N_19137,N_14007,N_10609);
nand U19138 (N_19138,N_13274,N_11961);
or U19139 (N_19139,N_12177,N_12766);
nor U19140 (N_19140,N_11338,N_11528);
or U19141 (N_19141,N_10319,N_14066);
nor U19142 (N_19142,N_14647,N_11499);
xor U19143 (N_19143,N_14269,N_14919);
and U19144 (N_19144,N_14337,N_13189);
nand U19145 (N_19145,N_12716,N_12906);
and U19146 (N_19146,N_14610,N_13247);
and U19147 (N_19147,N_11592,N_11024);
or U19148 (N_19148,N_10232,N_11461);
and U19149 (N_19149,N_13927,N_11182);
xor U19150 (N_19150,N_13787,N_10697);
nand U19151 (N_19151,N_11386,N_13792);
and U19152 (N_19152,N_12017,N_13152);
or U19153 (N_19153,N_11048,N_13024);
or U19154 (N_19154,N_13313,N_13895);
xnor U19155 (N_19155,N_14104,N_14186);
nor U19156 (N_19156,N_13512,N_14538);
nor U19157 (N_19157,N_10472,N_11076);
and U19158 (N_19158,N_10675,N_10225);
nor U19159 (N_19159,N_10887,N_14914);
nand U19160 (N_19160,N_13112,N_14073);
and U19161 (N_19161,N_12355,N_12219);
nand U19162 (N_19162,N_13550,N_12224);
nand U19163 (N_19163,N_11479,N_14894);
xnor U19164 (N_19164,N_12184,N_12833);
nor U19165 (N_19165,N_12027,N_10222);
and U19166 (N_19166,N_13527,N_13112);
nor U19167 (N_19167,N_12908,N_10312);
xnor U19168 (N_19168,N_12362,N_10613);
nor U19169 (N_19169,N_12804,N_13286);
nand U19170 (N_19170,N_13115,N_13193);
xnor U19171 (N_19171,N_12524,N_10091);
xnor U19172 (N_19172,N_10463,N_13620);
nor U19173 (N_19173,N_14169,N_12410);
and U19174 (N_19174,N_11831,N_11543);
nor U19175 (N_19175,N_11687,N_14456);
and U19176 (N_19176,N_13704,N_13881);
nor U19177 (N_19177,N_13640,N_14700);
xnor U19178 (N_19178,N_14426,N_12301);
or U19179 (N_19179,N_12103,N_13793);
or U19180 (N_19180,N_12385,N_11832);
nand U19181 (N_19181,N_11069,N_12295);
nor U19182 (N_19182,N_10305,N_13531);
nand U19183 (N_19183,N_10580,N_12414);
and U19184 (N_19184,N_13643,N_11395);
nand U19185 (N_19185,N_12462,N_12577);
and U19186 (N_19186,N_12725,N_11547);
or U19187 (N_19187,N_11929,N_11159);
nand U19188 (N_19188,N_12053,N_10948);
or U19189 (N_19189,N_10717,N_11586);
nand U19190 (N_19190,N_14393,N_10768);
xor U19191 (N_19191,N_10828,N_13365);
xnor U19192 (N_19192,N_14533,N_11197);
nand U19193 (N_19193,N_10659,N_11695);
xnor U19194 (N_19194,N_14333,N_14918);
nor U19195 (N_19195,N_11785,N_14271);
xnor U19196 (N_19196,N_13804,N_10259);
nor U19197 (N_19197,N_11764,N_13934);
nor U19198 (N_19198,N_14295,N_10574);
and U19199 (N_19199,N_14519,N_14501);
xor U19200 (N_19200,N_12012,N_13339);
nand U19201 (N_19201,N_14212,N_10981);
xor U19202 (N_19202,N_13620,N_13573);
and U19203 (N_19203,N_14990,N_11781);
and U19204 (N_19204,N_12220,N_12366);
xor U19205 (N_19205,N_10586,N_12808);
nand U19206 (N_19206,N_10695,N_12721);
nor U19207 (N_19207,N_10807,N_10244);
and U19208 (N_19208,N_12204,N_13422);
or U19209 (N_19209,N_10006,N_10310);
and U19210 (N_19210,N_10183,N_14278);
nand U19211 (N_19211,N_10166,N_12240);
and U19212 (N_19212,N_14928,N_10762);
and U19213 (N_19213,N_10059,N_14753);
xnor U19214 (N_19214,N_10312,N_10847);
and U19215 (N_19215,N_14034,N_14020);
and U19216 (N_19216,N_12466,N_13818);
or U19217 (N_19217,N_10312,N_12979);
xor U19218 (N_19218,N_12874,N_14536);
and U19219 (N_19219,N_10885,N_11741);
nor U19220 (N_19220,N_14887,N_12326);
xnor U19221 (N_19221,N_10257,N_13388);
nand U19222 (N_19222,N_13144,N_10137);
nor U19223 (N_19223,N_12468,N_12856);
nand U19224 (N_19224,N_13242,N_13261);
nor U19225 (N_19225,N_14568,N_12770);
nand U19226 (N_19226,N_14211,N_10085);
nor U19227 (N_19227,N_13276,N_11381);
xnor U19228 (N_19228,N_10143,N_10704);
nor U19229 (N_19229,N_10554,N_11544);
and U19230 (N_19230,N_11964,N_11061);
xnor U19231 (N_19231,N_10345,N_10808);
or U19232 (N_19232,N_11946,N_14747);
or U19233 (N_19233,N_10554,N_10109);
nand U19234 (N_19234,N_10438,N_10296);
and U19235 (N_19235,N_13286,N_13636);
xnor U19236 (N_19236,N_11754,N_12570);
xor U19237 (N_19237,N_12601,N_13265);
or U19238 (N_19238,N_14122,N_12089);
nand U19239 (N_19239,N_14312,N_13134);
nand U19240 (N_19240,N_12350,N_13959);
xor U19241 (N_19241,N_10818,N_10583);
xor U19242 (N_19242,N_13163,N_10839);
and U19243 (N_19243,N_10950,N_11010);
and U19244 (N_19244,N_14340,N_11424);
nand U19245 (N_19245,N_13476,N_13105);
nand U19246 (N_19246,N_13963,N_13579);
nand U19247 (N_19247,N_14879,N_14411);
and U19248 (N_19248,N_10658,N_10919);
nand U19249 (N_19249,N_13352,N_14715);
xor U19250 (N_19250,N_12618,N_12182);
nand U19251 (N_19251,N_13889,N_11631);
xnor U19252 (N_19252,N_12486,N_13323);
or U19253 (N_19253,N_14155,N_14289);
and U19254 (N_19254,N_10691,N_14367);
or U19255 (N_19255,N_14755,N_10095);
nor U19256 (N_19256,N_13490,N_12536);
or U19257 (N_19257,N_12923,N_10677);
and U19258 (N_19258,N_11554,N_10900);
nand U19259 (N_19259,N_11655,N_11620);
nor U19260 (N_19260,N_12033,N_13906);
nand U19261 (N_19261,N_14156,N_14018);
or U19262 (N_19262,N_14000,N_13608);
nand U19263 (N_19263,N_13970,N_11865);
nand U19264 (N_19264,N_11987,N_13970);
nor U19265 (N_19265,N_14642,N_13769);
nor U19266 (N_19266,N_11417,N_11859);
and U19267 (N_19267,N_12148,N_10901);
nand U19268 (N_19268,N_10950,N_11308);
or U19269 (N_19269,N_10002,N_12003);
nor U19270 (N_19270,N_10465,N_12642);
xnor U19271 (N_19271,N_11764,N_12185);
or U19272 (N_19272,N_11652,N_12005);
or U19273 (N_19273,N_11200,N_10549);
nand U19274 (N_19274,N_13788,N_14215);
or U19275 (N_19275,N_12645,N_13303);
and U19276 (N_19276,N_10440,N_11929);
xnor U19277 (N_19277,N_11414,N_14447);
nand U19278 (N_19278,N_10575,N_12066);
nand U19279 (N_19279,N_14201,N_11539);
nor U19280 (N_19280,N_10221,N_10873);
or U19281 (N_19281,N_12130,N_12052);
nor U19282 (N_19282,N_13469,N_14900);
nand U19283 (N_19283,N_14355,N_14545);
nand U19284 (N_19284,N_13663,N_13514);
xor U19285 (N_19285,N_10454,N_11273);
and U19286 (N_19286,N_14648,N_13974);
xor U19287 (N_19287,N_13191,N_14068);
and U19288 (N_19288,N_13829,N_12173);
or U19289 (N_19289,N_10257,N_12369);
and U19290 (N_19290,N_11712,N_11335);
nand U19291 (N_19291,N_14313,N_12421);
nand U19292 (N_19292,N_10043,N_13664);
and U19293 (N_19293,N_13825,N_13125);
nand U19294 (N_19294,N_13712,N_10510);
xor U19295 (N_19295,N_12449,N_11065);
xnor U19296 (N_19296,N_11370,N_10807);
nand U19297 (N_19297,N_13123,N_12565);
nor U19298 (N_19298,N_11266,N_13762);
nor U19299 (N_19299,N_10176,N_13250);
and U19300 (N_19300,N_11240,N_13705);
or U19301 (N_19301,N_13414,N_12069);
nand U19302 (N_19302,N_11225,N_11190);
xnor U19303 (N_19303,N_12487,N_13074);
and U19304 (N_19304,N_13202,N_11754);
and U19305 (N_19305,N_10443,N_14356);
nand U19306 (N_19306,N_14224,N_12397);
or U19307 (N_19307,N_10912,N_10154);
nand U19308 (N_19308,N_14689,N_14134);
or U19309 (N_19309,N_11346,N_10961);
or U19310 (N_19310,N_11310,N_14356);
and U19311 (N_19311,N_13357,N_11455);
and U19312 (N_19312,N_13810,N_12707);
nand U19313 (N_19313,N_10637,N_12649);
or U19314 (N_19314,N_13833,N_12810);
nor U19315 (N_19315,N_14579,N_13118);
and U19316 (N_19316,N_14408,N_14133);
and U19317 (N_19317,N_11387,N_12084);
nand U19318 (N_19318,N_12692,N_11606);
nand U19319 (N_19319,N_11587,N_10272);
nand U19320 (N_19320,N_10281,N_11358);
nor U19321 (N_19321,N_11956,N_12055);
and U19322 (N_19322,N_13180,N_11085);
or U19323 (N_19323,N_11802,N_10560);
xnor U19324 (N_19324,N_10735,N_12829);
and U19325 (N_19325,N_10460,N_14706);
xnor U19326 (N_19326,N_11383,N_14308);
nand U19327 (N_19327,N_14987,N_13661);
and U19328 (N_19328,N_11570,N_13886);
nor U19329 (N_19329,N_14377,N_14504);
or U19330 (N_19330,N_13446,N_10000);
xor U19331 (N_19331,N_13986,N_14594);
nor U19332 (N_19332,N_12400,N_10138);
and U19333 (N_19333,N_12776,N_12183);
nor U19334 (N_19334,N_13724,N_14672);
or U19335 (N_19335,N_12958,N_12045);
nor U19336 (N_19336,N_13413,N_11386);
or U19337 (N_19337,N_12147,N_12031);
and U19338 (N_19338,N_10473,N_11939);
nand U19339 (N_19339,N_13488,N_12606);
and U19340 (N_19340,N_10477,N_13449);
nand U19341 (N_19341,N_12723,N_11764);
or U19342 (N_19342,N_14067,N_12944);
xnor U19343 (N_19343,N_14582,N_13227);
and U19344 (N_19344,N_13202,N_10128);
xor U19345 (N_19345,N_11149,N_12847);
xnor U19346 (N_19346,N_11988,N_13982);
xnor U19347 (N_19347,N_12053,N_10387);
xnor U19348 (N_19348,N_14899,N_12764);
nor U19349 (N_19349,N_12679,N_13560);
nand U19350 (N_19350,N_12527,N_14686);
xor U19351 (N_19351,N_12776,N_10445);
and U19352 (N_19352,N_14003,N_14255);
nand U19353 (N_19353,N_10578,N_12523);
nand U19354 (N_19354,N_12786,N_13424);
and U19355 (N_19355,N_12753,N_11112);
nand U19356 (N_19356,N_10564,N_14402);
and U19357 (N_19357,N_14020,N_12721);
xor U19358 (N_19358,N_13021,N_10043);
or U19359 (N_19359,N_12785,N_12195);
nand U19360 (N_19360,N_12450,N_11643);
nand U19361 (N_19361,N_12484,N_10020);
or U19362 (N_19362,N_10461,N_14971);
nor U19363 (N_19363,N_10455,N_12542);
nand U19364 (N_19364,N_11307,N_11585);
and U19365 (N_19365,N_13902,N_10383);
xor U19366 (N_19366,N_14625,N_10361);
nor U19367 (N_19367,N_11451,N_13233);
and U19368 (N_19368,N_14097,N_10388);
nor U19369 (N_19369,N_14414,N_12909);
or U19370 (N_19370,N_13163,N_10089);
xnor U19371 (N_19371,N_10970,N_13430);
nor U19372 (N_19372,N_13784,N_13097);
or U19373 (N_19373,N_12878,N_10133);
or U19374 (N_19374,N_10862,N_14048);
nand U19375 (N_19375,N_14964,N_12407);
nand U19376 (N_19376,N_10149,N_10564);
or U19377 (N_19377,N_10862,N_13352);
nor U19378 (N_19378,N_14226,N_10694);
and U19379 (N_19379,N_10155,N_12406);
nand U19380 (N_19380,N_13394,N_12498);
nor U19381 (N_19381,N_12401,N_12001);
and U19382 (N_19382,N_12698,N_14618);
xor U19383 (N_19383,N_14852,N_11011);
and U19384 (N_19384,N_11802,N_10361);
or U19385 (N_19385,N_13372,N_11096);
nand U19386 (N_19386,N_12161,N_14179);
xnor U19387 (N_19387,N_12180,N_12185);
and U19388 (N_19388,N_10785,N_12108);
xnor U19389 (N_19389,N_10868,N_12575);
nor U19390 (N_19390,N_11161,N_11527);
or U19391 (N_19391,N_12054,N_14310);
nand U19392 (N_19392,N_14391,N_12846);
nor U19393 (N_19393,N_14710,N_14362);
nand U19394 (N_19394,N_14093,N_10745);
nor U19395 (N_19395,N_13828,N_10121);
nand U19396 (N_19396,N_11516,N_12163);
and U19397 (N_19397,N_11512,N_11897);
xnor U19398 (N_19398,N_11946,N_14552);
xor U19399 (N_19399,N_13527,N_13641);
xnor U19400 (N_19400,N_11422,N_13763);
nand U19401 (N_19401,N_12747,N_10944);
nor U19402 (N_19402,N_10248,N_12499);
nand U19403 (N_19403,N_10104,N_14287);
and U19404 (N_19404,N_13051,N_13240);
nor U19405 (N_19405,N_11986,N_14953);
or U19406 (N_19406,N_10080,N_12658);
nor U19407 (N_19407,N_12613,N_12978);
or U19408 (N_19408,N_12861,N_13984);
and U19409 (N_19409,N_11263,N_10421);
or U19410 (N_19410,N_11562,N_10671);
nand U19411 (N_19411,N_11295,N_12157);
or U19412 (N_19412,N_13793,N_11336);
nand U19413 (N_19413,N_14133,N_12204);
xnor U19414 (N_19414,N_11923,N_12600);
or U19415 (N_19415,N_12441,N_12989);
nor U19416 (N_19416,N_14884,N_10092);
and U19417 (N_19417,N_12034,N_10069);
and U19418 (N_19418,N_11585,N_11249);
and U19419 (N_19419,N_14032,N_12962);
and U19420 (N_19420,N_14896,N_13231);
and U19421 (N_19421,N_14226,N_12141);
nor U19422 (N_19422,N_13929,N_13451);
nand U19423 (N_19423,N_11412,N_12933);
or U19424 (N_19424,N_14058,N_10719);
xnor U19425 (N_19425,N_10471,N_12502);
or U19426 (N_19426,N_12466,N_10961);
and U19427 (N_19427,N_13488,N_10417);
nor U19428 (N_19428,N_14657,N_12444);
or U19429 (N_19429,N_13394,N_12672);
nand U19430 (N_19430,N_12143,N_12988);
nor U19431 (N_19431,N_14043,N_14869);
or U19432 (N_19432,N_12600,N_10188);
and U19433 (N_19433,N_10916,N_11092);
or U19434 (N_19434,N_11466,N_14132);
or U19435 (N_19435,N_11882,N_14467);
nand U19436 (N_19436,N_11895,N_14611);
xnor U19437 (N_19437,N_14068,N_14535);
or U19438 (N_19438,N_11132,N_14960);
xnor U19439 (N_19439,N_12614,N_12825);
and U19440 (N_19440,N_14960,N_11650);
nor U19441 (N_19441,N_13601,N_10400);
and U19442 (N_19442,N_10281,N_13756);
nor U19443 (N_19443,N_14672,N_10412);
nand U19444 (N_19444,N_13389,N_11991);
or U19445 (N_19445,N_11730,N_14959);
xnor U19446 (N_19446,N_11273,N_14052);
xnor U19447 (N_19447,N_11185,N_10580);
and U19448 (N_19448,N_13361,N_10266);
nor U19449 (N_19449,N_12989,N_12022);
xnor U19450 (N_19450,N_12620,N_10704);
and U19451 (N_19451,N_10694,N_13928);
or U19452 (N_19452,N_13586,N_11744);
and U19453 (N_19453,N_13725,N_13355);
and U19454 (N_19454,N_14555,N_13583);
xnor U19455 (N_19455,N_10293,N_14765);
and U19456 (N_19456,N_12638,N_10138);
or U19457 (N_19457,N_14426,N_13818);
nor U19458 (N_19458,N_11783,N_10248);
and U19459 (N_19459,N_11002,N_14227);
or U19460 (N_19460,N_13509,N_11803);
nand U19461 (N_19461,N_13579,N_12566);
nor U19462 (N_19462,N_11227,N_12584);
and U19463 (N_19463,N_13560,N_12304);
and U19464 (N_19464,N_10554,N_14872);
or U19465 (N_19465,N_13070,N_11160);
nor U19466 (N_19466,N_13924,N_12109);
xnor U19467 (N_19467,N_11189,N_11645);
nand U19468 (N_19468,N_13540,N_13094);
nor U19469 (N_19469,N_10881,N_14364);
nor U19470 (N_19470,N_13991,N_11218);
and U19471 (N_19471,N_11167,N_12529);
and U19472 (N_19472,N_11284,N_10670);
nand U19473 (N_19473,N_10983,N_10636);
nand U19474 (N_19474,N_10239,N_14238);
or U19475 (N_19475,N_11745,N_11795);
xor U19476 (N_19476,N_11849,N_13688);
and U19477 (N_19477,N_10964,N_14082);
nand U19478 (N_19478,N_13803,N_12945);
and U19479 (N_19479,N_10960,N_10873);
nor U19480 (N_19480,N_11223,N_10288);
or U19481 (N_19481,N_12309,N_13469);
or U19482 (N_19482,N_13441,N_10168);
or U19483 (N_19483,N_14411,N_14130);
xnor U19484 (N_19484,N_13970,N_11746);
nor U19485 (N_19485,N_11422,N_13503);
nor U19486 (N_19486,N_11744,N_13557);
xnor U19487 (N_19487,N_13917,N_10216);
or U19488 (N_19488,N_14396,N_10726);
nor U19489 (N_19489,N_11104,N_13291);
or U19490 (N_19490,N_13927,N_11512);
nor U19491 (N_19491,N_13163,N_14899);
and U19492 (N_19492,N_13411,N_10262);
xor U19493 (N_19493,N_13970,N_14762);
or U19494 (N_19494,N_12942,N_14087);
or U19495 (N_19495,N_14968,N_10499);
nand U19496 (N_19496,N_12513,N_11529);
nor U19497 (N_19497,N_12593,N_12904);
nor U19498 (N_19498,N_12419,N_14679);
and U19499 (N_19499,N_10837,N_14980);
nand U19500 (N_19500,N_14405,N_12947);
nor U19501 (N_19501,N_10264,N_13049);
or U19502 (N_19502,N_13167,N_13396);
nor U19503 (N_19503,N_11335,N_10448);
xor U19504 (N_19504,N_13706,N_10816);
xnor U19505 (N_19505,N_11743,N_12225);
nor U19506 (N_19506,N_14667,N_10897);
nand U19507 (N_19507,N_12598,N_12844);
nor U19508 (N_19508,N_14813,N_11672);
nor U19509 (N_19509,N_10883,N_10383);
or U19510 (N_19510,N_10460,N_11214);
xor U19511 (N_19511,N_12421,N_14566);
and U19512 (N_19512,N_10768,N_12127);
or U19513 (N_19513,N_11908,N_11317);
xnor U19514 (N_19514,N_13522,N_12933);
and U19515 (N_19515,N_11586,N_13131);
nor U19516 (N_19516,N_11969,N_13323);
or U19517 (N_19517,N_13963,N_11900);
nor U19518 (N_19518,N_12505,N_14256);
or U19519 (N_19519,N_14276,N_10775);
or U19520 (N_19520,N_11204,N_12612);
nand U19521 (N_19521,N_13356,N_11594);
or U19522 (N_19522,N_14878,N_10023);
or U19523 (N_19523,N_13908,N_12496);
or U19524 (N_19524,N_13334,N_14423);
nor U19525 (N_19525,N_14641,N_10972);
nor U19526 (N_19526,N_11082,N_12956);
or U19527 (N_19527,N_13144,N_11874);
or U19528 (N_19528,N_10238,N_11573);
and U19529 (N_19529,N_10454,N_10790);
nand U19530 (N_19530,N_14824,N_12780);
nor U19531 (N_19531,N_13220,N_14114);
xnor U19532 (N_19532,N_13778,N_10213);
nor U19533 (N_19533,N_13399,N_13957);
or U19534 (N_19534,N_13690,N_10914);
nand U19535 (N_19535,N_11691,N_11417);
or U19536 (N_19536,N_13075,N_10731);
xnor U19537 (N_19537,N_13447,N_11203);
or U19538 (N_19538,N_10573,N_12317);
xor U19539 (N_19539,N_10462,N_13531);
or U19540 (N_19540,N_11423,N_10693);
or U19541 (N_19541,N_12613,N_12591);
nor U19542 (N_19542,N_14361,N_13953);
or U19543 (N_19543,N_12349,N_13951);
nand U19544 (N_19544,N_12057,N_12335);
nand U19545 (N_19545,N_14356,N_14555);
or U19546 (N_19546,N_13800,N_10248);
nand U19547 (N_19547,N_12031,N_13720);
nor U19548 (N_19548,N_10109,N_12610);
xnor U19549 (N_19549,N_14250,N_10394);
xor U19550 (N_19550,N_14937,N_13205);
and U19551 (N_19551,N_10138,N_10708);
or U19552 (N_19552,N_13696,N_11937);
xnor U19553 (N_19553,N_12858,N_12634);
or U19554 (N_19554,N_13376,N_13477);
xor U19555 (N_19555,N_12190,N_13808);
or U19556 (N_19556,N_10729,N_11527);
nor U19557 (N_19557,N_10251,N_13759);
or U19558 (N_19558,N_13276,N_10646);
nand U19559 (N_19559,N_10467,N_12058);
and U19560 (N_19560,N_13121,N_11556);
or U19561 (N_19561,N_12504,N_11933);
nand U19562 (N_19562,N_12247,N_10442);
xor U19563 (N_19563,N_11917,N_12466);
and U19564 (N_19564,N_13763,N_12365);
xor U19565 (N_19565,N_12722,N_14117);
nand U19566 (N_19566,N_11356,N_14715);
and U19567 (N_19567,N_10970,N_14744);
nand U19568 (N_19568,N_11671,N_12626);
nor U19569 (N_19569,N_13976,N_13609);
nor U19570 (N_19570,N_12716,N_14681);
nand U19571 (N_19571,N_14894,N_14171);
and U19572 (N_19572,N_13966,N_11264);
or U19573 (N_19573,N_14804,N_13741);
or U19574 (N_19574,N_14206,N_13417);
or U19575 (N_19575,N_10621,N_13616);
and U19576 (N_19576,N_14053,N_13028);
nor U19577 (N_19577,N_11248,N_14882);
or U19578 (N_19578,N_14011,N_14399);
xnor U19579 (N_19579,N_10720,N_11138);
nor U19580 (N_19580,N_14584,N_13387);
xor U19581 (N_19581,N_11876,N_11837);
and U19582 (N_19582,N_11793,N_12349);
and U19583 (N_19583,N_12530,N_14436);
nor U19584 (N_19584,N_12242,N_14514);
xnor U19585 (N_19585,N_11762,N_13820);
or U19586 (N_19586,N_10210,N_14587);
and U19587 (N_19587,N_10086,N_11499);
xor U19588 (N_19588,N_12295,N_10057);
xor U19589 (N_19589,N_11747,N_12810);
nor U19590 (N_19590,N_11972,N_12672);
nor U19591 (N_19591,N_14002,N_12167);
or U19592 (N_19592,N_13340,N_10559);
and U19593 (N_19593,N_12004,N_11254);
or U19594 (N_19594,N_11435,N_13030);
and U19595 (N_19595,N_13338,N_11043);
xor U19596 (N_19596,N_10865,N_13158);
and U19597 (N_19597,N_12218,N_11018);
or U19598 (N_19598,N_10371,N_11603);
nor U19599 (N_19599,N_12799,N_10209);
xor U19600 (N_19600,N_11639,N_13491);
nor U19601 (N_19601,N_14233,N_12262);
xor U19602 (N_19602,N_11723,N_12481);
xnor U19603 (N_19603,N_12402,N_12438);
or U19604 (N_19604,N_14966,N_10402);
nand U19605 (N_19605,N_14516,N_13752);
xnor U19606 (N_19606,N_11530,N_13857);
and U19607 (N_19607,N_10581,N_13198);
or U19608 (N_19608,N_14236,N_10578);
nor U19609 (N_19609,N_11830,N_13886);
or U19610 (N_19610,N_13461,N_13491);
nor U19611 (N_19611,N_13789,N_10908);
nor U19612 (N_19612,N_11718,N_12326);
nand U19613 (N_19613,N_10530,N_13651);
xnor U19614 (N_19614,N_13289,N_10615);
nand U19615 (N_19615,N_14095,N_11679);
nor U19616 (N_19616,N_13148,N_12632);
xnor U19617 (N_19617,N_12963,N_10181);
or U19618 (N_19618,N_12559,N_12849);
xnor U19619 (N_19619,N_10655,N_12342);
nand U19620 (N_19620,N_10234,N_11847);
and U19621 (N_19621,N_11730,N_10852);
xnor U19622 (N_19622,N_14744,N_11788);
or U19623 (N_19623,N_13661,N_12688);
or U19624 (N_19624,N_10977,N_10570);
nor U19625 (N_19625,N_10126,N_10481);
or U19626 (N_19626,N_11215,N_10983);
xnor U19627 (N_19627,N_13086,N_10345);
nand U19628 (N_19628,N_10868,N_14703);
xnor U19629 (N_19629,N_12719,N_11462);
or U19630 (N_19630,N_13409,N_14871);
or U19631 (N_19631,N_12263,N_13111);
nor U19632 (N_19632,N_13918,N_11693);
xnor U19633 (N_19633,N_10187,N_10900);
nor U19634 (N_19634,N_13866,N_12137);
and U19635 (N_19635,N_11447,N_10226);
nor U19636 (N_19636,N_12053,N_10587);
nand U19637 (N_19637,N_12789,N_12193);
nor U19638 (N_19638,N_10898,N_13509);
nor U19639 (N_19639,N_12492,N_10905);
nor U19640 (N_19640,N_13266,N_10037);
xor U19641 (N_19641,N_14688,N_11405);
or U19642 (N_19642,N_11041,N_10831);
nand U19643 (N_19643,N_14780,N_12130);
nand U19644 (N_19644,N_14529,N_13065);
nor U19645 (N_19645,N_14496,N_14743);
xnor U19646 (N_19646,N_12675,N_10557);
nor U19647 (N_19647,N_10954,N_13331);
nand U19648 (N_19648,N_10430,N_13496);
xor U19649 (N_19649,N_10723,N_10662);
or U19650 (N_19650,N_10492,N_10085);
xnor U19651 (N_19651,N_14947,N_13665);
and U19652 (N_19652,N_12281,N_11965);
nand U19653 (N_19653,N_13167,N_10290);
and U19654 (N_19654,N_14877,N_14730);
nand U19655 (N_19655,N_12364,N_10070);
or U19656 (N_19656,N_12080,N_10325);
nand U19657 (N_19657,N_14728,N_14033);
and U19658 (N_19658,N_10424,N_11692);
nor U19659 (N_19659,N_12622,N_10160);
nand U19660 (N_19660,N_14754,N_10603);
nand U19661 (N_19661,N_14988,N_11832);
nand U19662 (N_19662,N_10644,N_13049);
xnor U19663 (N_19663,N_11163,N_14147);
or U19664 (N_19664,N_14564,N_13740);
or U19665 (N_19665,N_14085,N_11348);
or U19666 (N_19666,N_12542,N_11712);
and U19667 (N_19667,N_14869,N_11331);
nand U19668 (N_19668,N_13485,N_12888);
nand U19669 (N_19669,N_10822,N_10086);
xnor U19670 (N_19670,N_13664,N_14682);
xnor U19671 (N_19671,N_14936,N_10973);
and U19672 (N_19672,N_10417,N_14971);
xnor U19673 (N_19673,N_10481,N_12983);
nor U19674 (N_19674,N_13685,N_12586);
or U19675 (N_19675,N_10494,N_12581);
or U19676 (N_19676,N_10039,N_14030);
xnor U19677 (N_19677,N_13599,N_14389);
nor U19678 (N_19678,N_13123,N_13977);
xor U19679 (N_19679,N_14177,N_11802);
or U19680 (N_19680,N_11063,N_14172);
nand U19681 (N_19681,N_11236,N_10529);
nor U19682 (N_19682,N_13328,N_10892);
nor U19683 (N_19683,N_12794,N_10619);
nand U19684 (N_19684,N_11683,N_12419);
nand U19685 (N_19685,N_12193,N_14440);
nand U19686 (N_19686,N_13735,N_14839);
and U19687 (N_19687,N_14524,N_10218);
or U19688 (N_19688,N_10856,N_13735);
nand U19689 (N_19689,N_12903,N_10786);
xor U19690 (N_19690,N_13997,N_10479);
xnor U19691 (N_19691,N_10150,N_14161);
nand U19692 (N_19692,N_12568,N_11630);
xnor U19693 (N_19693,N_12110,N_11766);
or U19694 (N_19694,N_13286,N_14871);
and U19695 (N_19695,N_14164,N_11077);
nor U19696 (N_19696,N_14849,N_11801);
nor U19697 (N_19697,N_10666,N_12756);
and U19698 (N_19698,N_13525,N_14221);
xor U19699 (N_19699,N_14107,N_11564);
and U19700 (N_19700,N_14604,N_10205);
nand U19701 (N_19701,N_14260,N_12648);
nor U19702 (N_19702,N_13805,N_14319);
nand U19703 (N_19703,N_11435,N_13063);
nor U19704 (N_19704,N_10248,N_10296);
xnor U19705 (N_19705,N_10679,N_11187);
nand U19706 (N_19706,N_13848,N_11896);
xnor U19707 (N_19707,N_12055,N_10652);
and U19708 (N_19708,N_11045,N_10051);
or U19709 (N_19709,N_12814,N_14356);
or U19710 (N_19710,N_14630,N_11843);
xnor U19711 (N_19711,N_12349,N_10901);
and U19712 (N_19712,N_10148,N_14211);
and U19713 (N_19713,N_12482,N_14685);
or U19714 (N_19714,N_10131,N_12503);
and U19715 (N_19715,N_12233,N_11217);
nand U19716 (N_19716,N_11870,N_14631);
and U19717 (N_19717,N_14430,N_13621);
nor U19718 (N_19718,N_11232,N_10284);
nand U19719 (N_19719,N_13891,N_13595);
and U19720 (N_19720,N_13659,N_13673);
or U19721 (N_19721,N_12455,N_11032);
nand U19722 (N_19722,N_10479,N_14829);
nand U19723 (N_19723,N_12131,N_11490);
xor U19724 (N_19724,N_14138,N_11919);
and U19725 (N_19725,N_14307,N_14945);
or U19726 (N_19726,N_14362,N_13245);
and U19727 (N_19727,N_14972,N_11321);
and U19728 (N_19728,N_13405,N_14187);
nor U19729 (N_19729,N_11867,N_14151);
nor U19730 (N_19730,N_11235,N_13227);
nor U19731 (N_19731,N_12931,N_13248);
xor U19732 (N_19732,N_14128,N_13834);
nor U19733 (N_19733,N_13453,N_10470);
nand U19734 (N_19734,N_10212,N_10514);
nand U19735 (N_19735,N_11868,N_14535);
and U19736 (N_19736,N_13851,N_14836);
or U19737 (N_19737,N_11373,N_13773);
nand U19738 (N_19738,N_12969,N_10199);
nor U19739 (N_19739,N_11335,N_12914);
nand U19740 (N_19740,N_14856,N_14707);
xor U19741 (N_19741,N_14655,N_12829);
xnor U19742 (N_19742,N_13361,N_13685);
and U19743 (N_19743,N_12517,N_12315);
or U19744 (N_19744,N_13987,N_14750);
or U19745 (N_19745,N_12331,N_13947);
nor U19746 (N_19746,N_11552,N_10055);
nand U19747 (N_19747,N_14555,N_13228);
and U19748 (N_19748,N_10887,N_11197);
and U19749 (N_19749,N_12028,N_13178);
or U19750 (N_19750,N_11477,N_14527);
and U19751 (N_19751,N_13432,N_11142);
and U19752 (N_19752,N_14337,N_11512);
and U19753 (N_19753,N_13242,N_13171);
or U19754 (N_19754,N_14145,N_11755);
nor U19755 (N_19755,N_11538,N_12394);
or U19756 (N_19756,N_10259,N_11359);
or U19757 (N_19757,N_11900,N_10475);
or U19758 (N_19758,N_14724,N_14061);
and U19759 (N_19759,N_10032,N_14079);
xnor U19760 (N_19760,N_10411,N_13457);
nand U19761 (N_19761,N_11524,N_12433);
or U19762 (N_19762,N_14553,N_13599);
nand U19763 (N_19763,N_11684,N_10193);
and U19764 (N_19764,N_11489,N_14123);
and U19765 (N_19765,N_10541,N_14827);
or U19766 (N_19766,N_13254,N_13946);
or U19767 (N_19767,N_13059,N_12285);
nand U19768 (N_19768,N_13536,N_13403);
or U19769 (N_19769,N_11487,N_11949);
nor U19770 (N_19770,N_13196,N_14579);
or U19771 (N_19771,N_11710,N_10005);
nor U19772 (N_19772,N_13681,N_11531);
or U19773 (N_19773,N_11599,N_12666);
and U19774 (N_19774,N_10722,N_14259);
nor U19775 (N_19775,N_13133,N_12990);
or U19776 (N_19776,N_14733,N_14059);
nand U19777 (N_19777,N_11503,N_10144);
or U19778 (N_19778,N_12556,N_13517);
and U19779 (N_19779,N_13511,N_13376);
or U19780 (N_19780,N_13133,N_14944);
xor U19781 (N_19781,N_12320,N_13381);
nor U19782 (N_19782,N_13896,N_11738);
xor U19783 (N_19783,N_10345,N_14682);
nor U19784 (N_19784,N_11609,N_12926);
or U19785 (N_19785,N_11008,N_12909);
nand U19786 (N_19786,N_10988,N_11216);
nand U19787 (N_19787,N_13399,N_10384);
nor U19788 (N_19788,N_11997,N_11603);
nand U19789 (N_19789,N_10470,N_10393);
and U19790 (N_19790,N_13838,N_11087);
nand U19791 (N_19791,N_13946,N_14172);
and U19792 (N_19792,N_14563,N_10023);
nor U19793 (N_19793,N_10327,N_14031);
nand U19794 (N_19794,N_14359,N_12329);
nor U19795 (N_19795,N_12105,N_12733);
and U19796 (N_19796,N_11504,N_13557);
and U19797 (N_19797,N_11467,N_14440);
nor U19798 (N_19798,N_11253,N_13035);
xnor U19799 (N_19799,N_10469,N_10842);
xnor U19800 (N_19800,N_14041,N_10579);
xnor U19801 (N_19801,N_10407,N_12600);
nand U19802 (N_19802,N_14902,N_11895);
xnor U19803 (N_19803,N_10290,N_11057);
nor U19804 (N_19804,N_12054,N_11553);
nand U19805 (N_19805,N_12605,N_11110);
or U19806 (N_19806,N_13039,N_14479);
nor U19807 (N_19807,N_13602,N_14813);
and U19808 (N_19808,N_14495,N_12863);
or U19809 (N_19809,N_12952,N_13639);
or U19810 (N_19810,N_13522,N_14102);
and U19811 (N_19811,N_10739,N_13955);
nand U19812 (N_19812,N_13253,N_10352);
nand U19813 (N_19813,N_12113,N_12518);
and U19814 (N_19814,N_12583,N_10636);
xnor U19815 (N_19815,N_14213,N_11372);
nand U19816 (N_19816,N_10952,N_10220);
xor U19817 (N_19817,N_12798,N_10598);
xnor U19818 (N_19818,N_10876,N_14647);
xor U19819 (N_19819,N_11795,N_11773);
and U19820 (N_19820,N_11138,N_13986);
and U19821 (N_19821,N_11852,N_14187);
and U19822 (N_19822,N_13892,N_13884);
or U19823 (N_19823,N_10777,N_10424);
nand U19824 (N_19824,N_12552,N_11796);
or U19825 (N_19825,N_12754,N_13988);
nand U19826 (N_19826,N_13138,N_14738);
nand U19827 (N_19827,N_13356,N_14507);
or U19828 (N_19828,N_10444,N_14774);
nand U19829 (N_19829,N_13000,N_13965);
and U19830 (N_19830,N_14724,N_11273);
xor U19831 (N_19831,N_10806,N_14606);
nor U19832 (N_19832,N_11324,N_14366);
and U19833 (N_19833,N_11810,N_10636);
and U19834 (N_19834,N_11932,N_14347);
nand U19835 (N_19835,N_11369,N_11816);
nand U19836 (N_19836,N_13399,N_11631);
nor U19837 (N_19837,N_11779,N_10963);
nor U19838 (N_19838,N_12503,N_11478);
xor U19839 (N_19839,N_11772,N_12591);
nor U19840 (N_19840,N_11965,N_14684);
or U19841 (N_19841,N_11862,N_12617);
nand U19842 (N_19842,N_12658,N_14496);
nand U19843 (N_19843,N_13110,N_10781);
or U19844 (N_19844,N_10869,N_11527);
nor U19845 (N_19845,N_10618,N_12399);
or U19846 (N_19846,N_14921,N_11582);
nand U19847 (N_19847,N_14687,N_14346);
and U19848 (N_19848,N_11756,N_12815);
xnor U19849 (N_19849,N_14061,N_10423);
nand U19850 (N_19850,N_11814,N_11727);
xnor U19851 (N_19851,N_10841,N_14537);
nand U19852 (N_19852,N_10796,N_11967);
xor U19853 (N_19853,N_10663,N_10722);
or U19854 (N_19854,N_14640,N_10791);
nor U19855 (N_19855,N_13534,N_14078);
xnor U19856 (N_19856,N_14178,N_13204);
or U19857 (N_19857,N_12630,N_10702);
nor U19858 (N_19858,N_10606,N_13457);
and U19859 (N_19859,N_12344,N_11450);
xor U19860 (N_19860,N_13446,N_12884);
nor U19861 (N_19861,N_11869,N_10280);
and U19862 (N_19862,N_14797,N_13881);
nand U19863 (N_19863,N_10878,N_13079);
nand U19864 (N_19864,N_12198,N_11412);
or U19865 (N_19865,N_11456,N_12786);
xnor U19866 (N_19866,N_13858,N_13449);
and U19867 (N_19867,N_13228,N_14243);
nor U19868 (N_19868,N_10263,N_14201);
or U19869 (N_19869,N_11105,N_12857);
nand U19870 (N_19870,N_14405,N_10182);
xnor U19871 (N_19871,N_13580,N_10544);
and U19872 (N_19872,N_12264,N_12341);
xor U19873 (N_19873,N_12446,N_13971);
xnor U19874 (N_19874,N_10839,N_12231);
nand U19875 (N_19875,N_13684,N_13913);
nor U19876 (N_19876,N_14419,N_12167);
nor U19877 (N_19877,N_13005,N_13284);
nor U19878 (N_19878,N_14291,N_11276);
or U19879 (N_19879,N_14295,N_11368);
nor U19880 (N_19880,N_10855,N_14404);
or U19881 (N_19881,N_12053,N_10503);
nand U19882 (N_19882,N_14264,N_14509);
nand U19883 (N_19883,N_12621,N_13523);
nand U19884 (N_19884,N_14887,N_13973);
nor U19885 (N_19885,N_10518,N_11089);
and U19886 (N_19886,N_12220,N_10898);
nor U19887 (N_19887,N_14197,N_10293);
nor U19888 (N_19888,N_12487,N_10993);
nand U19889 (N_19889,N_11811,N_12559);
nor U19890 (N_19890,N_14841,N_14939);
nand U19891 (N_19891,N_14016,N_11271);
xor U19892 (N_19892,N_13678,N_14803);
nand U19893 (N_19893,N_12396,N_12094);
xnor U19894 (N_19894,N_13744,N_13033);
or U19895 (N_19895,N_14597,N_13080);
and U19896 (N_19896,N_13871,N_14161);
nand U19897 (N_19897,N_10122,N_11928);
and U19898 (N_19898,N_13274,N_11466);
xnor U19899 (N_19899,N_10562,N_12750);
xor U19900 (N_19900,N_10658,N_13672);
nand U19901 (N_19901,N_13474,N_11081);
nand U19902 (N_19902,N_11097,N_14466);
nor U19903 (N_19903,N_14622,N_12686);
nand U19904 (N_19904,N_13039,N_14305);
xnor U19905 (N_19905,N_10742,N_11578);
xor U19906 (N_19906,N_10115,N_11167);
nor U19907 (N_19907,N_11062,N_11676);
or U19908 (N_19908,N_11443,N_13291);
and U19909 (N_19909,N_12345,N_14777);
or U19910 (N_19910,N_12659,N_14016);
or U19911 (N_19911,N_13435,N_11681);
and U19912 (N_19912,N_13835,N_13824);
nor U19913 (N_19913,N_13267,N_12333);
nand U19914 (N_19914,N_10727,N_10419);
and U19915 (N_19915,N_12380,N_11997);
and U19916 (N_19916,N_13494,N_12114);
nor U19917 (N_19917,N_14665,N_13293);
nor U19918 (N_19918,N_12005,N_10429);
nand U19919 (N_19919,N_11206,N_12039);
nand U19920 (N_19920,N_12311,N_10981);
and U19921 (N_19921,N_10622,N_12655);
xor U19922 (N_19922,N_13075,N_10115);
nand U19923 (N_19923,N_11789,N_11433);
xnor U19924 (N_19924,N_10162,N_10920);
and U19925 (N_19925,N_10092,N_12402);
xnor U19926 (N_19926,N_12764,N_13818);
and U19927 (N_19927,N_11703,N_13054);
nor U19928 (N_19928,N_10719,N_10316);
nor U19929 (N_19929,N_12915,N_11840);
nand U19930 (N_19930,N_13598,N_10706);
nor U19931 (N_19931,N_14246,N_10040);
or U19932 (N_19932,N_13518,N_13446);
or U19933 (N_19933,N_13218,N_10289);
or U19934 (N_19934,N_11289,N_11083);
or U19935 (N_19935,N_12620,N_12235);
xor U19936 (N_19936,N_14357,N_13103);
xor U19937 (N_19937,N_10043,N_11135);
nand U19938 (N_19938,N_10583,N_13507);
nor U19939 (N_19939,N_12554,N_13403);
xnor U19940 (N_19940,N_11717,N_14293);
nor U19941 (N_19941,N_10807,N_14006);
nand U19942 (N_19942,N_14017,N_14766);
or U19943 (N_19943,N_12119,N_12521);
and U19944 (N_19944,N_12668,N_14944);
nor U19945 (N_19945,N_14118,N_14829);
and U19946 (N_19946,N_13369,N_13601);
or U19947 (N_19947,N_10042,N_12869);
or U19948 (N_19948,N_11480,N_14463);
and U19949 (N_19949,N_14110,N_10586);
nand U19950 (N_19950,N_11253,N_14658);
xor U19951 (N_19951,N_10010,N_10240);
and U19952 (N_19952,N_12703,N_11108);
and U19953 (N_19953,N_12786,N_14778);
and U19954 (N_19954,N_10588,N_11148);
or U19955 (N_19955,N_10055,N_13107);
and U19956 (N_19956,N_13140,N_12417);
nor U19957 (N_19957,N_12629,N_14938);
xnor U19958 (N_19958,N_11143,N_12155);
nor U19959 (N_19959,N_10131,N_12656);
nand U19960 (N_19960,N_10480,N_13962);
and U19961 (N_19961,N_11561,N_14797);
xnor U19962 (N_19962,N_14570,N_11148);
or U19963 (N_19963,N_12588,N_12272);
and U19964 (N_19964,N_12890,N_10292);
or U19965 (N_19965,N_13095,N_13966);
nor U19966 (N_19966,N_12495,N_13933);
and U19967 (N_19967,N_11870,N_13334);
nor U19968 (N_19968,N_14577,N_14006);
nand U19969 (N_19969,N_10573,N_13685);
xor U19970 (N_19970,N_12608,N_11053);
nor U19971 (N_19971,N_12987,N_11267);
or U19972 (N_19972,N_13731,N_14199);
xor U19973 (N_19973,N_12386,N_11221);
nand U19974 (N_19974,N_14842,N_11626);
nor U19975 (N_19975,N_14946,N_14851);
nor U19976 (N_19976,N_14028,N_12338);
or U19977 (N_19977,N_12105,N_14151);
nor U19978 (N_19978,N_11455,N_11512);
nand U19979 (N_19979,N_13471,N_11113);
xor U19980 (N_19980,N_11325,N_13767);
xor U19981 (N_19981,N_10270,N_12230);
xnor U19982 (N_19982,N_13909,N_12502);
nor U19983 (N_19983,N_11893,N_12958);
nor U19984 (N_19984,N_14155,N_12730);
nor U19985 (N_19985,N_11513,N_10877);
nor U19986 (N_19986,N_12346,N_11594);
nand U19987 (N_19987,N_11267,N_11134);
nand U19988 (N_19988,N_11188,N_14128);
nand U19989 (N_19989,N_11117,N_14883);
nand U19990 (N_19990,N_12496,N_14956);
nor U19991 (N_19991,N_10641,N_10422);
and U19992 (N_19992,N_11216,N_13775);
or U19993 (N_19993,N_14250,N_13251);
nand U19994 (N_19994,N_14219,N_13173);
xnor U19995 (N_19995,N_14942,N_10994);
nor U19996 (N_19996,N_11524,N_10592);
nand U19997 (N_19997,N_12867,N_14569);
xor U19998 (N_19998,N_13741,N_10038);
nor U19999 (N_19999,N_11876,N_14332);
or U20000 (N_20000,N_18009,N_16989);
and U20001 (N_20001,N_18059,N_15354);
xnor U20002 (N_20002,N_19726,N_17762);
nand U20003 (N_20003,N_17833,N_19633);
nand U20004 (N_20004,N_19513,N_18698);
nor U20005 (N_20005,N_15924,N_17914);
and U20006 (N_20006,N_17014,N_18315);
or U20007 (N_20007,N_19781,N_16199);
or U20008 (N_20008,N_17897,N_16786);
nand U20009 (N_20009,N_16245,N_15119);
nand U20010 (N_20010,N_18632,N_18561);
xnor U20011 (N_20011,N_19165,N_16191);
xnor U20012 (N_20012,N_16031,N_16576);
and U20013 (N_20013,N_16793,N_15501);
xnor U20014 (N_20014,N_17487,N_19709);
and U20015 (N_20015,N_16707,N_18734);
nor U20016 (N_20016,N_18126,N_19368);
nand U20017 (N_20017,N_16243,N_18015);
xnor U20018 (N_20018,N_17994,N_19126);
or U20019 (N_20019,N_15810,N_17184);
and U20020 (N_20020,N_17848,N_15601);
nor U20021 (N_20021,N_17212,N_19842);
or U20022 (N_20022,N_17176,N_19637);
nor U20023 (N_20023,N_17609,N_16290);
nand U20024 (N_20024,N_18820,N_18569);
or U20025 (N_20025,N_16858,N_19993);
or U20026 (N_20026,N_15172,N_15013);
xnor U20027 (N_20027,N_16028,N_15240);
and U20028 (N_20028,N_18308,N_15811);
nor U20029 (N_20029,N_16265,N_15914);
nor U20030 (N_20030,N_18165,N_16526);
and U20031 (N_20031,N_16422,N_17866);
nand U20032 (N_20032,N_18671,N_16886);
nand U20033 (N_20033,N_17168,N_16991);
and U20034 (N_20034,N_15068,N_16156);
and U20035 (N_20035,N_16273,N_16530);
xor U20036 (N_20036,N_15908,N_16435);
nand U20037 (N_20037,N_16518,N_19973);
and U20038 (N_20038,N_16445,N_18025);
and U20039 (N_20039,N_15826,N_16878);
or U20040 (N_20040,N_19622,N_15479);
nand U20041 (N_20041,N_16682,N_15786);
or U20042 (N_20042,N_19505,N_18726);
or U20043 (N_20043,N_17805,N_15436);
and U20044 (N_20044,N_17399,N_15935);
and U20045 (N_20045,N_19546,N_17594);
nor U20046 (N_20046,N_17954,N_18081);
or U20047 (N_20047,N_16630,N_15129);
nand U20048 (N_20048,N_19558,N_16167);
nor U20049 (N_20049,N_16078,N_16798);
nand U20050 (N_20050,N_18916,N_17813);
and U20051 (N_20051,N_18251,N_19946);
and U20052 (N_20052,N_18658,N_16342);
nand U20053 (N_20053,N_17383,N_16140);
nor U20054 (N_20054,N_16559,N_17429);
nand U20055 (N_20055,N_17831,N_19584);
or U20056 (N_20056,N_19020,N_16838);
xnor U20057 (N_20057,N_17923,N_16366);
and U20058 (N_20058,N_15791,N_17968);
xor U20059 (N_20059,N_17462,N_15413);
nand U20060 (N_20060,N_16824,N_16351);
or U20061 (N_20061,N_19043,N_19522);
nand U20062 (N_20062,N_17922,N_19421);
xor U20063 (N_20063,N_16086,N_16928);
nand U20064 (N_20064,N_15528,N_15160);
or U20065 (N_20065,N_16169,N_15142);
and U20066 (N_20066,N_16355,N_19838);
nand U20067 (N_20067,N_18495,N_16238);
or U20068 (N_20068,N_15046,N_16799);
or U20069 (N_20069,N_17064,N_17534);
and U20070 (N_20070,N_16549,N_15855);
and U20071 (N_20071,N_19554,N_19200);
and U20072 (N_20072,N_15925,N_18090);
nor U20073 (N_20073,N_15599,N_17421);
xor U20074 (N_20074,N_16396,N_17082);
or U20075 (N_20075,N_18945,N_16249);
xnor U20076 (N_20076,N_16834,N_18362);
and U20077 (N_20077,N_15262,N_17250);
nor U20078 (N_20078,N_19444,N_16353);
nor U20079 (N_20079,N_15126,N_18737);
and U20080 (N_20080,N_18605,N_18548);
nor U20081 (N_20081,N_18514,N_16157);
nand U20082 (N_20082,N_16606,N_19605);
xor U20083 (N_20083,N_18778,N_17556);
nand U20084 (N_20084,N_18089,N_19283);
xnor U20085 (N_20085,N_19237,N_19198);
xnor U20086 (N_20086,N_18976,N_15752);
nor U20087 (N_20087,N_18442,N_16041);
nor U20088 (N_20088,N_17856,N_19601);
or U20089 (N_20089,N_15514,N_15330);
or U20090 (N_20090,N_17052,N_17048);
and U20091 (N_20091,N_19231,N_19386);
or U20092 (N_20092,N_15133,N_17449);
xor U20093 (N_20093,N_17989,N_17215);
and U20094 (N_20094,N_16742,N_19476);
xor U20095 (N_20095,N_17069,N_15636);
and U20096 (N_20096,N_16462,N_18859);
nor U20097 (N_20097,N_16634,N_17226);
nor U20098 (N_20098,N_15638,N_18369);
and U20099 (N_20099,N_19492,N_19398);
xnor U20100 (N_20100,N_16547,N_17007);
xor U20101 (N_20101,N_15266,N_15841);
or U20102 (N_20102,N_16125,N_15536);
or U20103 (N_20103,N_16531,N_16487);
nor U20104 (N_20104,N_18982,N_16474);
and U20105 (N_20105,N_18249,N_19260);
nor U20106 (N_20106,N_16190,N_17379);
or U20107 (N_20107,N_15645,N_19806);
and U20108 (N_20108,N_17141,N_18659);
and U20109 (N_20109,N_16754,N_15952);
nor U20110 (N_20110,N_15264,N_15081);
or U20111 (N_20111,N_18274,N_19006);
xnor U20112 (N_20112,N_17160,N_18669);
or U20113 (N_20113,N_17512,N_17471);
and U20114 (N_20114,N_17896,N_19538);
nand U20115 (N_20115,N_18870,N_16274);
and U20116 (N_20116,N_15340,N_16962);
nor U20117 (N_20117,N_18591,N_18790);
nand U20118 (N_20118,N_16228,N_16189);
nand U20119 (N_20119,N_15852,N_17294);
and U20120 (N_20120,N_15828,N_18691);
and U20121 (N_20121,N_16034,N_19818);
nor U20122 (N_20122,N_17157,N_16451);
xnor U20123 (N_20123,N_15593,N_16821);
and U20124 (N_20124,N_19009,N_18085);
xnor U20125 (N_20125,N_17652,N_19755);
or U20126 (N_20126,N_19834,N_16850);
nor U20127 (N_20127,N_18088,N_15726);
and U20128 (N_20128,N_15432,N_19096);
or U20129 (N_20129,N_15541,N_15858);
and U20130 (N_20130,N_16323,N_17400);
nand U20131 (N_20131,N_18879,N_18335);
or U20132 (N_20132,N_15485,N_15230);
nand U20133 (N_20133,N_15152,N_15916);
xnor U20134 (N_20134,N_17349,N_19338);
nand U20135 (N_20135,N_19581,N_17941);
or U20136 (N_20136,N_15490,N_15722);
xor U20137 (N_20137,N_18707,N_17960);
or U20138 (N_20138,N_15381,N_17834);
or U20139 (N_20139,N_18023,N_17140);
nor U20140 (N_20140,N_15894,N_18831);
nand U20141 (N_20141,N_18364,N_15701);
xor U20142 (N_20142,N_16399,N_16168);
and U20143 (N_20143,N_15538,N_18505);
nor U20144 (N_20144,N_18163,N_19955);
and U20145 (N_20145,N_16807,N_16649);
xnor U20146 (N_20146,N_18533,N_15323);
nand U20147 (N_20147,N_19322,N_16889);
and U20148 (N_20148,N_18921,N_18153);
and U20149 (N_20149,N_18437,N_15205);
and U20150 (N_20150,N_17962,N_17242);
and U20151 (N_20151,N_16144,N_16002);
or U20152 (N_20152,N_15798,N_15387);
and U20153 (N_20153,N_15375,N_15865);
nand U20154 (N_20154,N_15734,N_19877);
xnor U20155 (N_20155,N_19761,N_19341);
and U20156 (N_20156,N_19108,N_17439);
nand U20157 (N_20157,N_15754,N_19613);
nor U20158 (N_20158,N_17790,N_19156);
nor U20159 (N_20159,N_18462,N_15024);
and U20160 (N_20160,N_16218,N_17861);
or U20161 (N_20161,N_18942,N_18801);
and U20162 (N_20162,N_15074,N_17729);
and U20163 (N_20163,N_18557,N_15910);
and U20164 (N_20164,N_17966,N_19887);
xnor U20165 (N_20165,N_18575,N_18094);
nor U20166 (N_20166,N_18809,N_18936);
and U20167 (N_20167,N_16550,N_18823);
nand U20168 (N_20168,N_19238,N_15080);
nor U20169 (N_20169,N_19248,N_18397);
nor U20170 (N_20170,N_18325,N_16759);
nand U20171 (N_20171,N_17980,N_17751);
or U20172 (N_20172,N_17531,N_15114);
and U20173 (N_20173,N_18227,N_16113);
nor U20174 (N_20174,N_17889,N_19769);
nor U20175 (N_20175,N_18050,N_19595);
nor U20176 (N_20176,N_17171,N_16483);
and U20177 (N_20177,N_18123,N_15980);
nor U20178 (N_20178,N_16450,N_16865);
and U20179 (N_20179,N_19753,N_16470);
or U20180 (N_20180,N_17820,N_19590);
nor U20181 (N_20181,N_17728,N_18917);
nor U20182 (N_20182,N_19742,N_19236);
and U20183 (N_20183,N_17000,N_17047);
nand U20184 (N_20184,N_17901,N_16769);
xnor U20185 (N_20185,N_19649,N_19913);
nor U20186 (N_20186,N_19155,N_17338);
and U20187 (N_20187,N_18337,N_19139);
nand U20188 (N_20188,N_19115,N_16502);
or U20189 (N_20189,N_18560,N_18565);
and U20190 (N_20190,N_15419,N_19975);
nand U20191 (N_20191,N_15449,N_16418);
nor U20192 (N_20192,N_16348,N_18600);
or U20193 (N_20193,N_16874,N_19378);
or U20194 (N_20194,N_19128,N_18861);
or U20195 (N_20195,N_17500,N_17243);
or U20196 (N_20196,N_18811,N_15179);
nor U20197 (N_20197,N_15579,N_18226);
nor U20198 (N_20198,N_15878,N_15030);
xor U20199 (N_20199,N_18950,N_15648);
xnor U20200 (N_20200,N_16693,N_15989);
xor U20201 (N_20201,N_18262,N_16772);
and U20202 (N_20202,N_15655,N_17555);
nand U20203 (N_20203,N_16272,N_19258);
nand U20204 (N_20204,N_19187,N_15048);
or U20205 (N_20205,N_18865,N_19631);
nor U20206 (N_20206,N_15972,N_15590);
and U20207 (N_20207,N_16567,N_15769);
and U20208 (N_20208,N_19738,N_19798);
nand U20209 (N_20209,N_15026,N_18405);
xor U20210 (N_20210,N_19962,N_15736);
nor U20211 (N_20211,N_18990,N_17010);
or U20212 (N_20212,N_19579,N_15446);
xor U20213 (N_20213,N_16556,N_15797);
nand U20214 (N_20214,N_17905,N_15524);
nand U20215 (N_20215,N_18963,N_17104);
xnor U20216 (N_20216,N_18073,N_18520);
or U20217 (N_20217,N_16854,N_19981);
nand U20218 (N_20218,N_17291,N_16967);
xnor U20219 (N_20219,N_19387,N_17528);
xnor U20220 (N_20220,N_18832,N_19242);
and U20221 (N_20221,N_15635,N_16747);
xnor U20222 (N_20222,N_18516,N_18633);
nand U20223 (N_20223,N_18834,N_18645);
xnor U20224 (N_20224,N_17667,N_15960);
nor U20225 (N_20225,N_15134,N_19944);
or U20226 (N_20226,N_18989,N_16101);
xor U20227 (N_20227,N_17043,N_15516);
and U20228 (N_20228,N_16334,N_16994);
or U20229 (N_20229,N_16611,N_16760);
xor U20230 (N_20230,N_19045,N_19971);
xnor U20231 (N_20231,N_17716,N_17722);
xor U20232 (N_20232,N_19344,N_19473);
or U20233 (N_20233,N_15058,N_18266);
or U20234 (N_20234,N_17492,N_15421);
or U20235 (N_20235,N_18768,N_18665);
nor U20236 (N_20236,N_19446,N_15695);
nand U20237 (N_20237,N_18889,N_18955);
or U20238 (N_20238,N_15233,N_16204);
nor U20239 (N_20239,N_17319,N_19431);
xnor U20240 (N_20240,N_17423,N_15539);
nand U20241 (N_20241,N_18711,N_15245);
or U20242 (N_20242,N_15480,N_18424);
and U20243 (N_20243,N_19662,N_19166);
nor U20244 (N_20244,N_17763,N_16667);
nand U20245 (N_20245,N_16395,N_16489);
xnor U20246 (N_20246,N_19771,N_16115);
and U20247 (N_20247,N_15303,N_19550);
and U20248 (N_20248,N_15214,N_18212);
and U20249 (N_20249,N_18544,N_15212);
nand U20250 (N_20250,N_15385,N_18223);
or U20251 (N_20251,N_18291,N_17666);
and U20252 (N_20252,N_16347,N_15084);
and U20253 (N_20253,N_18987,N_19196);
and U20254 (N_20254,N_15429,N_18733);
xnor U20255 (N_20255,N_18935,N_17198);
xnor U20256 (N_20256,N_19162,N_19385);
or U20257 (N_20257,N_16969,N_17008);
or U20258 (N_20258,N_18136,N_18128);
nand U20259 (N_20259,N_19744,N_16847);
or U20260 (N_20260,N_16719,N_15241);
or U20261 (N_20261,N_18087,N_18345);
and U20262 (N_20262,N_16280,N_17299);
nand U20263 (N_20263,N_16105,N_19556);
and U20264 (N_20264,N_18531,N_17774);
or U20265 (N_20265,N_19240,N_15039);
and U20266 (N_20266,N_17267,N_19369);
nor U20267 (N_20267,N_17680,N_15656);
or U20268 (N_20268,N_19690,N_16553);
nor U20269 (N_20269,N_16261,N_19869);
or U20270 (N_20270,N_18339,N_18205);
or U20271 (N_20271,N_18751,N_15149);
and U20272 (N_20272,N_15368,N_16340);
and U20273 (N_20273,N_16027,N_15380);
xor U20274 (N_20274,N_17650,N_17339);
nor U20275 (N_20275,N_15162,N_19669);
and U20276 (N_20276,N_16770,N_16388);
nand U20277 (N_20277,N_18101,N_17653);
xor U20278 (N_20278,N_17920,N_18293);
xnor U20279 (N_20279,N_17705,N_17692);
and U20280 (N_20280,N_16701,N_18439);
nand U20281 (N_20281,N_16458,N_15905);
nand U20282 (N_20282,N_19987,N_16235);
or U20283 (N_20283,N_19185,N_17187);
nor U20284 (N_20284,N_16880,N_19297);
nor U20285 (N_20285,N_18947,N_19434);
xnor U20286 (N_20286,N_17668,N_19364);
nor U20287 (N_20287,N_19880,N_18482);
nand U20288 (N_20288,N_19527,N_17882);
nand U20289 (N_20289,N_19339,N_18474);
or U20290 (N_20290,N_17418,N_17314);
xor U20291 (N_20291,N_18352,N_18190);
xor U20292 (N_20292,N_19775,N_18688);
or U20293 (N_20293,N_17624,N_16011);
nand U20294 (N_20294,N_15711,N_16364);
nor U20295 (N_20295,N_19016,N_18735);
or U20296 (N_20296,N_18766,N_19611);
nor U20297 (N_20297,N_16308,N_19990);
xnor U20298 (N_20298,N_17659,N_16575);
and U20299 (N_20299,N_15073,N_19026);
xnor U20300 (N_20300,N_18968,N_16780);
or U20301 (N_20301,N_19285,N_19934);
nor U20302 (N_20302,N_19206,N_18109);
nor U20303 (N_20303,N_19326,N_19278);
xor U20304 (N_20304,N_18347,N_18067);
or U20305 (N_20305,N_19114,N_15629);
nand U20306 (N_20306,N_15888,N_17024);
nand U20307 (N_20307,N_17527,N_18783);
and U20308 (N_20308,N_16892,N_15349);
nor U20309 (N_20309,N_18164,N_17511);
and U20310 (N_20310,N_15954,N_19168);
and U20311 (N_20311,N_17988,N_19901);
nand U20312 (N_20312,N_17095,N_16151);
xor U20313 (N_20313,N_18385,N_19794);
nand U20314 (N_20314,N_17554,N_16869);
nand U20315 (N_20315,N_16134,N_18620);
nor U20316 (N_20316,N_17929,N_16866);
nand U20317 (N_20317,N_15738,N_15299);
xnor U20318 (N_20318,N_19507,N_17658);
and U20319 (N_20319,N_15886,N_15132);
nor U20320 (N_20320,N_15519,N_18703);
nor U20321 (N_20321,N_19409,N_15622);
or U20322 (N_20322,N_15145,N_16241);
or U20323 (N_20323,N_17295,N_17493);
or U20324 (N_20324,N_19273,N_18946);
and U20325 (N_20325,N_17185,N_16851);
nor U20326 (N_20326,N_19050,N_15244);
xor U20327 (N_20327,N_18056,N_16279);
or U20328 (N_20328,N_18286,N_19158);
nor U20329 (N_20329,N_15667,N_16494);
nor U20330 (N_20330,N_15424,N_15127);
and U20331 (N_20331,N_18463,N_17484);
and U20332 (N_20332,N_16995,N_16110);
nor U20333 (N_20333,N_17045,N_18106);
or U20334 (N_20334,N_16753,N_19508);
and U20335 (N_20335,N_16790,N_18305);
and U20336 (N_20336,N_19014,N_16216);
or U20337 (N_20337,N_17661,N_19843);
or U20338 (N_20338,N_15596,N_18209);
xnor U20339 (N_20339,N_19257,N_19047);
or U20340 (N_20340,N_18594,N_15877);
nand U20341 (N_20341,N_17823,N_19792);
xnor U20342 (N_20342,N_15720,N_17231);
nand U20343 (N_20343,N_16424,N_18730);
xor U20344 (N_20344,N_19589,N_18393);
or U20345 (N_20345,N_18431,N_16372);
nor U20346 (N_20346,N_15566,N_16876);
xor U20347 (N_20347,N_16463,N_15343);
and U20348 (N_20348,N_16416,N_16820);
xnor U20349 (N_20349,N_18203,N_19697);
nor U20350 (N_20350,N_18629,N_18608);
and U20351 (N_20351,N_15056,N_19562);
nand U20352 (N_20352,N_15966,N_17997);
and U20353 (N_20353,N_15123,N_16224);
nand U20354 (N_20354,N_18327,N_18784);
and U20355 (N_20355,N_16705,N_16839);
nor U20356 (N_20356,N_15203,N_17396);
nor U20357 (N_20357,N_17489,N_18619);
or U20358 (N_20358,N_18721,N_16525);
nor U20359 (N_20359,N_16519,N_16049);
nor U20360 (N_20360,N_19621,N_17842);
nand U20361 (N_20361,N_16400,N_19524);
nand U20362 (N_20362,N_18804,N_16501);
or U20363 (N_20363,N_15307,N_16205);
nand U20364 (N_20364,N_17902,N_17748);
xor U20365 (N_20365,N_15334,N_18845);
xor U20366 (N_20366,N_15112,N_19347);
and U20367 (N_20367,N_18958,N_16877);
nor U20368 (N_20368,N_15053,N_16040);
nor U20369 (N_20369,N_18785,N_17051);
nor U20370 (N_20370,N_16923,N_17323);
nand U20371 (N_20371,N_16259,N_17083);
nand U20372 (N_20372,N_19317,N_15361);
nand U20373 (N_20373,N_19077,N_16785);
and U20374 (N_20374,N_19053,N_15871);
nand U20375 (N_20375,N_16072,N_18863);
and U20376 (N_20376,N_17227,N_19432);
nand U20377 (N_20377,N_19182,N_15627);
nor U20378 (N_20378,N_19447,N_19241);
and U20379 (N_20379,N_19396,N_15760);
nand U20380 (N_20380,N_17928,N_17384);
and U20381 (N_20381,N_19692,N_15669);
or U20382 (N_20382,N_15092,N_17180);
nor U20383 (N_20383,N_16180,N_18360);
nor U20384 (N_20384,N_18466,N_16673);
nand U20385 (N_20385,N_18547,N_15365);
nor U20386 (N_20386,N_18398,N_18399);
nor U20387 (N_20387,N_15344,N_16337);
nand U20388 (N_20388,N_18595,N_15192);
xor U20389 (N_20389,N_15876,N_16875);
nand U20390 (N_20390,N_18668,N_17860);
or U20391 (N_20391,N_19864,N_15746);
and U20392 (N_20392,N_19786,N_15500);
nand U20393 (N_20393,N_15922,N_18167);
or U20394 (N_20394,N_19705,N_15728);
nor U20395 (N_20395,N_17362,N_17906);
and U20396 (N_20396,N_15772,N_19404);
nand U20397 (N_20397,N_19342,N_18937);
nand U20398 (N_20398,N_15758,N_17284);
nor U20399 (N_20399,N_17266,N_17166);
and U20400 (N_20400,N_18815,N_16058);
nor U20401 (N_20401,N_15891,N_19064);
nand U20402 (N_20402,N_15766,N_18752);
nor U20403 (N_20403,N_16260,N_18539);
nor U20404 (N_20404,N_15806,N_19092);
and U20405 (N_20405,N_19259,N_15603);
or U20406 (N_20406,N_17119,N_18195);
or U20407 (N_20407,N_16005,N_17070);
nor U20408 (N_20408,N_19749,N_17735);
nand U20409 (N_20409,N_18422,N_19923);
or U20410 (N_20410,N_19885,N_19376);
or U20411 (N_20411,N_19334,N_15450);
and U20412 (N_20412,N_15540,N_17279);
or U20413 (N_20413,N_15971,N_18610);
or U20414 (N_20414,N_16263,N_18792);
or U20415 (N_20415,N_18161,N_18746);
or U20416 (N_20416,N_16499,N_19866);
and U20417 (N_20417,N_16116,N_16479);
and U20418 (N_20418,N_19687,N_16762);
nand U20419 (N_20419,N_19216,N_18553);
nand U20420 (N_20420,N_18927,N_19974);
and U20421 (N_20421,N_19003,N_19251);
nor U20422 (N_20422,N_19418,N_16150);
nand U20423 (N_20423,N_18744,N_19416);
or U20424 (N_20424,N_18184,N_15866);
nand U20425 (N_20425,N_16440,N_19573);
nor U20426 (N_20426,N_18687,N_19180);
or U20427 (N_20427,N_16979,N_18064);
or U20428 (N_20428,N_18493,N_16871);
or U20429 (N_20429,N_18760,N_19942);
xnor U20430 (N_20430,N_15584,N_16225);
nand U20431 (N_20431,N_17733,N_16376);
and U20432 (N_20432,N_16903,N_16695);
or U20433 (N_20433,N_18871,N_18674);
nand U20434 (N_20434,N_19281,N_17887);
nand U20435 (N_20435,N_17621,N_19666);
nand U20436 (N_20436,N_15146,N_15243);
and U20437 (N_20437,N_17755,N_18856);
xnor U20438 (N_20438,N_19295,N_17483);
xnor U20439 (N_20439,N_16295,N_15598);
or U20440 (N_20440,N_16117,N_19881);
nand U20441 (N_20441,N_15225,N_16711);
or U20442 (N_20442,N_18018,N_19337);
or U20443 (N_20443,N_15833,N_18238);
nand U20444 (N_20444,N_19069,N_17604);
nand U20445 (N_20445,N_16133,N_19463);
nor U20446 (N_20446,N_16666,N_17101);
xnor U20447 (N_20447,N_19644,N_18559);
nand U20448 (N_20448,N_19498,N_17347);
or U20449 (N_20449,N_15136,N_19090);
nand U20450 (N_20450,N_16981,N_18851);
xnor U20451 (N_20451,N_19325,N_15776);
and U20452 (N_20452,N_17590,N_16867);
nand U20453 (N_20453,N_19907,N_19719);
nand U20454 (N_20454,N_16025,N_18130);
or U20455 (N_20455,N_19487,N_17036);
xor U20456 (N_20456,N_16944,N_18459);
xnor U20457 (N_20457,N_18827,N_18006);
xor U20458 (N_20458,N_16936,N_18366);
nand U20459 (N_20459,N_16738,N_16748);
or U20460 (N_20460,N_16596,N_15059);
or U20461 (N_20461,N_15255,N_17220);
nor U20462 (N_20462,N_18214,N_17791);
xor U20463 (N_20463,N_16370,N_18627);
or U20464 (N_20464,N_15729,N_17642);
and U20465 (N_20465,N_16375,N_15571);
and U20466 (N_20466,N_15995,N_19125);
and U20467 (N_20467,N_16650,N_17038);
and U20468 (N_20468,N_19530,N_19673);
or U20469 (N_20469,N_18607,N_19360);
nor U20470 (N_20470,N_17461,N_15724);
nand U20471 (N_20471,N_19335,N_16062);
xnor U20472 (N_20472,N_18105,N_19262);
nand U20473 (N_20473,N_18762,N_18017);
nor U20474 (N_20474,N_16047,N_18704);
or U20475 (N_20475,N_19723,N_17208);
or U20476 (N_20476,N_17127,N_19677);
nor U20477 (N_20477,N_17352,N_19356);
nor U20478 (N_20478,N_15895,N_15577);
and U20479 (N_20479,N_19226,N_19645);
and U20480 (N_20480,N_17948,N_18417);
xnor U20481 (N_20481,N_17845,N_19087);
and U20482 (N_20482,N_16159,N_16590);
xor U20483 (N_20483,N_16581,N_15606);
and U20484 (N_20484,N_15427,N_19711);
or U20485 (N_20485,N_16929,N_18225);
xnor U20486 (N_20486,N_18319,N_17759);
xnor U20487 (N_20487,N_18798,N_16633);
or U20488 (N_20488,N_18825,N_17093);
or U20489 (N_20489,N_19056,N_19411);
xnor U20490 (N_20490,N_15312,N_19233);
nor U20491 (N_20491,N_18512,N_18450);
and U20492 (N_20492,N_19703,N_16070);
and U20493 (N_20493,N_19983,N_19460);
or U20494 (N_20494,N_19557,N_16552);
nand U20495 (N_20495,N_15759,N_19620);
xor U20496 (N_20496,N_16848,N_17712);
xor U20497 (N_20497,N_17702,N_15659);
xnor U20498 (N_20498,N_16817,N_15252);
xnor U20499 (N_20499,N_15078,N_19675);
and U20500 (N_20500,N_18156,N_15787);
or U20501 (N_20501,N_16024,N_15176);
nor U20502 (N_20502,N_19586,N_17075);
or U20503 (N_20503,N_19531,N_18074);
nand U20504 (N_20504,N_15719,N_17537);
or U20505 (N_20505,N_15840,N_16870);
nand U20506 (N_20506,N_17046,N_19038);
nand U20507 (N_20507,N_15364,N_16032);
nor U20508 (N_20508,N_19807,N_17268);
xnor U20509 (N_20509,N_19247,N_19395);
or U20510 (N_20510,N_17998,N_17937);
and U20511 (N_20511,N_18464,N_15277);
nand U20512 (N_20512,N_19821,N_19791);
xnor U20513 (N_20513,N_19480,N_19564);
nor U20514 (N_20514,N_17246,N_19919);
or U20515 (N_20515,N_18230,N_17363);
or U20516 (N_20516,N_19999,N_15180);
or U20517 (N_20517,N_15200,N_18538);
or U20518 (N_20518,N_16276,N_17067);
nand U20519 (N_20519,N_19729,N_19861);
nand U20520 (N_20520,N_17721,N_15699);
and U20521 (N_20521,N_19081,N_17524);
nand U20522 (N_20522,N_18000,N_15947);
nor U20523 (N_20523,N_17033,N_17434);
xnor U20524 (N_20524,N_16935,N_19865);
and U20525 (N_20525,N_16973,N_16727);
nand U20526 (N_20526,N_19735,N_16778);
or U20527 (N_20527,N_15019,N_16941);
nor U20528 (N_20528,N_18492,N_16773);
xor U20529 (N_20529,N_16832,N_16812);
or U20530 (N_20530,N_15371,N_19737);
xor U20531 (N_20531,N_15529,N_17482);
and U20532 (N_20532,N_16099,N_19203);
xnor U20533 (N_20533,N_15016,N_17356);
nor U20534 (N_20534,N_17739,N_16781);
nor U20535 (N_20535,N_17145,N_19095);
and U20536 (N_20536,N_19488,N_15543);
or U20537 (N_20537,N_16262,N_18646);
nand U20538 (N_20538,N_15892,N_18941);
xnor U20539 (N_20539,N_15911,N_16537);
and U20540 (N_20540,N_15282,N_19549);
or U20541 (N_20541,N_19871,N_19765);
xnor U20542 (N_20542,N_17009,N_19272);
or U20543 (N_20543,N_18664,N_16597);
nor U20544 (N_20544,N_17156,N_18055);
and U20545 (N_20545,N_18786,N_18476);
nor U20546 (N_20546,N_17520,N_18530);
or U20547 (N_20547,N_18791,N_16325);
nand U20548 (N_20548,N_18993,N_17073);
xor U20549 (N_20549,N_19074,N_19793);
xor U20550 (N_20550,N_19129,N_15434);
and U20551 (N_20551,N_17129,N_18586);
nor U20552 (N_20552,N_15100,N_19788);
nor U20553 (N_20553,N_15700,N_17592);
or U20554 (N_20554,N_17687,N_17699);
and U20555 (N_20555,N_17466,N_18158);
nand U20556 (N_20556,N_18211,N_18451);
and U20557 (N_20557,N_19147,N_16696);
xor U20558 (N_20558,N_19355,N_18813);
or U20559 (N_20559,N_16532,N_16919);
nand U20560 (N_20560,N_18676,N_17214);
xnor U20561 (N_20561,N_17063,N_15077);
or U20562 (N_20562,N_15567,N_18841);
nand U20563 (N_20563,N_19503,N_15285);
nor U20564 (N_20564,N_17086,N_19435);
xor U20565 (N_20565,N_15228,N_16541);
and U20566 (N_20566,N_15642,N_19269);
nand U20567 (N_20567,N_18890,N_18970);
xnor U20568 (N_20568,N_16933,N_15270);
and U20569 (N_20569,N_17765,N_17252);
xnor U20570 (N_20570,N_19664,N_16795);
and U20571 (N_20571,N_17999,N_18853);
xor U20572 (N_20572,N_16584,N_18881);
nand U20573 (N_20573,N_19193,N_16339);
nor U20574 (N_20574,N_16872,N_15997);
nand U20575 (N_20575,N_15353,N_16560);
xor U20576 (N_20576,N_15658,N_16697);
nor U20577 (N_20577,N_15652,N_18732);
or U20578 (N_20578,N_16401,N_16186);
nor U20579 (N_20579,N_19921,N_16411);
nor U20580 (N_20580,N_17839,N_15672);
or U20581 (N_20581,N_19676,N_17382);
or U20582 (N_20582,N_18564,N_15415);
xor U20583 (N_20583,N_17787,N_17378);
xor U20584 (N_20584,N_15739,N_18061);
xnor U20585 (N_20585,N_16053,N_19250);
and U20586 (N_20586,N_15904,N_17432);
and U20587 (N_20587,N_16642,N_16736);
or U20588 (N_20588,N_16913,N_16258);
nor U20589 (N_20589,N_18192,N_19540);
or U20590 (N_20590,N_18295,N_18342);
xnor U20591 (N_20591,N_15012,N_15496);
or U20592 (N_20592,N_18742,N_18876);
nand U20593 (N_20593,N_15899,N_15713);
xnor U20594 (N_20594,N_16840,N_15508);
or U20595 (N_20595,N_17256,N_19466);
xnor U20596 (N_20596,N_18383,N_18628);
nor U20597 (N_20597,N_16800,N_15578);
nor U20598 (N_20598,N_17177,N_17239);
nor U20599 (N_20599,N_16543,N_16819);
or U20600 (N_20600,N_16495,N_18765);
nand U20601 (N_20601,N_15725,N_15341);
nor U20602 (N_20602,N_19164,N_15259);
and U20603 (N_20603,N_16749,N_16562);
nand U20604 (N_20604,N_17785,N_16794);
nand U20605 (N_20605,N_17921,N_15920);
and U20606 (N_20606,N_15442,N_17094);
and U20607 (N_20607,N_15651,N_18263);
and U20608 (N_20608,N_18913,N_17867);
or U20609 (N_20609,N_15624,N_15850);
nand U20610 (N_20610,N_15350,N_15022);
nor U20611 (N_20611,N_15513,N_16148);
xor U20612 (N_20612,N_17028,N_16327);
nor U20613 (N_20613,N_19560,N_15064);
nor U20614 (N_20614,N_18057,N_15497);
xnor U20615 (N_20615,N_16946,N_17199);
nand U20616 (N_20616,N_16955,N_17933);
and U20617 (N_20617,N_18418,N_15909);
nand U20618 (N_20618,N_16951,N_16587);
and U20619 (N_20619,N_18518,N_16573);
nor U20620 (N_20620,N_15360,N_18440);
or U20621 (N_20621,N_16731,N_16554);
xor U20622 (N_20622,N_17830,N_19433);
nor U20623 (N_20623,N_19770,N_17431);
nand U20624 (N_20624,N_15358,N_19350);
nand U20625 (N_20625,N_17569,N_15226);
nand U20626 (N_20626,N_18489,N_16548);
xor U20627 (N_20627,N_18139,N_17174);
nand U20628 (N_20628,N_15633,N_15052);
or U20629 (N_20629,N_15410,N_16291);
and U20630 (N_20630,N_19679,N_19483);
or U20631 (N_20631,N_19320,N_15352);
or U20632 (N_20632,N_16383,N_15055);
and U20633 (N_20633,N_17518,N_19234);
nand U20634 (N_20634,N_17855,N_17758);
or U20635 (N_20635,N_17032,N_15780);
or U20636 (N_20636,N_15166,N_17975);
and U20637 (N_20637,N_19181,N_19977);
and U20638 (N_20638,N_17022,N_18661);
and U20639 (N_20639,N_15408,N_18452);
nand U20640 (N_20640,N_18977,N_18596);
xnor U20641 (N_20641,N_18381,N_17163);
or U20642 (N_20642,N_18833,N_17367);
xor U20643 (N_20643,N_17292,N_16322);
and U20644 (N_20644,N_19657,N_15632);
or U20645 (N_20645,N_18245,N_19706);
or U20646 (N_20646,N_16803,N_19169);
nor U20647 (N_20647,N_19683,N_16409);
or U20648 (N_20648,N_19448,N_17258);
or U20649 (N_20649,N_15804,N_18117);
and U20650 (N_20650,N_16881,N_15171);
or U20651 (N_20651,N_18256,N_18292);
or U20652 (N_20652,N_19345,N_17131);
nor U20653 (N_20653,N_16578,N_16934);
and U20654 (N_20654,N_19668,N_16947);
nor U20655 (N_20655,N_16608,N_18083);
and U20656 (N_20656,N_17898,N_16108);
and U20657 (N_20657,N_19936,N_18176);
or U20658 (N_20658,N_15710,N_16623);
and U20659 (N_20659,N_17322,N_17983);
nand U20660 (N_20660,N_16367,N_18320);
nand U20661 (N_20661,N_17812,N_18621);
and U20662 (N_20662,N_15174,N_16333);
nor U20663 (N_20663,N_17553,N_16240);
or U20664 (N_20664,N_18975,N_15553);
nand U20665 (N_20665,N_18477,N_15903);
and U20666 (N_20666,N_17583,N_17688);
and U20667 (N_20667,N_15957,N_15223);
nand U20668 (N_20668,N_16741,N_15605);
or U20669 (N_20669,N_17843,N_18330);
nand U20670 (N_20670,N_17793,N_15304);
and U20671 (N_20671,N_19072,N_18408);
nand U20672 (N_20672,N_16956,N_15477);
xor U20673 (N_20673,N_15721,N_15859);
or U20674 (N_20674,N_17618,N_16659);
nand U20675 (N_20675,N_15531,N_18697);
xor U20676 (N_20676,N_15156,N_19964);
xor U20677 (N_20677,N_15491,N_16632);
xnor U20678 (N_20678,N_17803,N_19456);
or U20679 (N_20679,N_17570,N_19486);
nand U20680 (N_20680,N_15236,N_17125);
nor U20681 (N_20681,N_15573,N_18578);
xor U20682 (N_20682,N_17329,N_16591);
xnor U20683 (N_20683,N_18283,N_19321);
xor U20684 (N_20684,N_16296,N_16811);
nor U20685 (N_20685,N_18396,N_16456);
nor U20686 (N_20686,N_16917,N_17505);
nor U20687 (N_20687,N_18540,N_15781);
and U20688 (N_20688,N_15001,N_16358);
nand U20689 (N_20689,N_19388,N_15836);
and U20690 (N_20690,N_15140,N_18324);
or U20691 (N_20691,N_18582,N_15662);
nand U20692 (N_20692,N_16061,N_15591);
or U20693 (N_20693,N_17674,N_16129);
xnor U20694 (N_20694,N_15499,N_15657);
xnor U20695 (N_20695,N_19058,N_18636);
or U20696 (N_20696,N_15099,N_17771);
nor U20697 (N_20697,N_16890,N_15939);
nand U20698 (N_20698,N_17625,N_16831);
or U20699 (N_20699,N_19478,N_19359);
nor U20700 (N_20700,N_16536,N_19220);
or U20701 (N_20701,N_15765,N_19629);
and U20702 (N_20702,N_17477,N_16209);
nand U20703 (N_20703,N_17216,N_17282);
and U20704 (N_20704,N_16905,N_15884);
and U20705 (N_20705,N_16277,N_17133);
nand U20706 (N_20706,N_18624,N_16505);
xnor U20707 (N_20707,N_16460,N_16313);
or U20708 (N_20708,N_19438,N_18349);
nor U20709 (N_20709,N_19840,N_17300);
or U20710 (N_20710,N_19314,N_16635);
xnor U20711 (N_20711,N_18277,N_15696);
xor U20712 (N_20712,N_16616,N_17143);
nand U20713 (N_20713,N_18488,N_17217);
or U20714 (N_20714,N_17139,N_17944);
nor U20715 (N_20715,N_19229,N_17990);
or U20716 (N_20716,N_16195,N_16478);
nand U20717 (N_20717,N_16615,N_19106);
xnor U20718 (N_20718,N_18490,N_16746);
xor U20719 (N_20719,N_16257,N_15423);
or U20720 (N_20720,N_17516,N_17390);
nand U20721 (N_20721,N_19812,N_16570);
xnor U20722 (N_20722,N_16896,N_15926);
and U20723 (N_20723,N_15617,N_17211);
or U20724 (N_20724,N_15986,N_16433);
xnor U20725 (N_20725,N_15452,N_17281);
nor U20726 (N_20726,N_19702,N_17006);
or U20727 (N_20727,N_16836,N_15495);
and U20728 (N_20728,N_16301,N_18837);
and U20729 (N_20729,N_19373,N_16201);
nor U20730 (N_20730,N_17596,N_16266);
or U20731 (N_20731,N_16911,N_15934);
and U20732 (N_20732,N_18830,N_17469);
and U20733 (N_20733,N_15556,N_19585);
or U20734 (N_20734,N_18534,N_19626);
nor U20735 (N_20735,N_17496,N_18983);
and U20736 (N_20736,N_18897,N_18053);
and U20737 (N_20737,N_15463,N_15562);
nor U20738 (N_20738,N_15021,N_15944);
and U20739 (N_20739,N_18773,N_19306);
xor U20740 (N_20740,N_19979,N_16540);
and U20741 (N_20741,N_19704,N_17497);
nor U20742 (N_20742,N_18551,N_17137);
nand U20743 (N_20743,N_15558,N_15979);
nor U20744 (N_20744,N_15561,N_17162);
and U20745 (N_20745,N_17269,N_15388);
nor U20746 (N_20746,N_15647,N_16879);
nor U20747 (N_20747,N_18086,N_18019);
xor U20748 (N_20748,N_19614,N_17873);
or U20749 (N_20749,N_16906,N_19094);
xnor U20750 (N_20750,N_18037,N_18857);
and U20751 (N_20751,N_15936,N_19380);
and U20752 (N_20752,N_16963,N_16307);
or U20753 (N_20753,N_17459,N_17110);
nor U20754 (N_20754,N_16709,N_18186);
nand U20755 (N_20755,N_19963,N_19820);
xor U20756 (N_20756,N_18480,N_18051);
or U20757 (N_20757,N_17891,N_19496);
xor U20758 (N_20758,N_15938,N_19174);
nor U20759 (N_20759,N_16298,N_17796);
and U20760 (N_20760,N_15807,N_19961);
and U20761 (N_20761,N_16582,N_15088);
xnor U20762 (N_20762,N_16909,N_19232);
and U20763 (N_20763,N_16442,N_17235);
and U20764 (N_20764,N_18446,N_19826);
or U20765 (N_20765,N_15321,N_15879);
nor U20766 (N_20766,N_19635,N_17320);
nand U20767 (N_20767,N_19222,N_18468);
or U20768 (N_20768,N_19551,N_19802);
nand U20769 (N_20769,N_15454,N_15441);
nor U20770 (N_20770,N_17610,N_17951);
and U20771 (N_20771,N_15329,N_18447);
or U20772 (N_20772,N_18157,N_17513);
or U20773 (N_20773,N_16686,N_17971);
nor U20774 (N_20774,N_17982,N_18503);
nor U20775 (N_20775,N_18739,N_19417);
and U20776 (N_20776,N_17580,N_15276);
or U20777 (N_20777,N_15912,N_17271);
or U20778 (N_20778,N_19516,N_18906);
or U20779 (N_20779,N_19493,N_17021);
xor U20780 (N_20780,N_19479,N_18307);
xnor U20781 (N_20781,N_17607,N_18441);
and U20782 (N_20782,N_17877,N_17470);
nand U20783 (N_20783,N_16164,N_19996);
or U20784 (N_20784,N_17875,N_16314);
nor U20785 (N_20785,N_18054,N_17708);
xnor U20786 (N_20786,N_16815,N_18208);
xnor U20787 (N_20787,N_18239,N_15535);
nor U20788 (N_20788,N_19470,N_19583);
nand U20789 (N_20789,N_19348,N_19068);
xnor U20790 (N_20790,N_18370,N_15318);
xnor U20791 (N_20791,N_16160,N_18012);
nor U20792 (N_20792,N_18718,N_18866);
nor U20793 (N_20793,N_16402,N_16200);
or U20794 (N_20794,N_19394,N_16067);
and U20795 (N_20795,N_18522,N_17325);
and U20796 (N_20796,N_18457,N_17773);
and U20797 (N_20797,N_17274,N_17940);
nor U20798 (N_20798,N_19302,N_17837);
nand U20799 (N_20799,N_19136,N_15475);
or U20800 (N_20800,N_15272,N_18338);
nor U20801 (N_20801,N_16345,N_18272);
and U20802 (N_20802,N_17696,N_19437);
or U20803 (N_20803,N_19824,N_19930);
or U20804 (N_20804,N_15305,N_15990);
or U20805 (N_20805,N_17561,N_17460);
or U20806 (N_20806,N_15619,N_19904);
and U20807 (N_20807,N_17040,N_15274);
nand U20808 (N_20808,N_18852,N_15254);
xor U20809 (N_20809,N_16637,N_16949);
or U20810 (N_20810,N_15317,N_18717);
and U20811 (N_20811,N_18643,N_17730);
and U20812 (N_20812,N_16221,N_18332);
and U20813 (N_20813,N_19795,N_17710);
nand U20814 (N_20814,N_15880,N_18098);
xor U20815 (N_20815,N_16750,N_15355);
nor U20816 (N_20816,N_19526,N_16755);
nand U20817 (N_20817,N_15515,N_19183);
nand U20818 (N_20818,N_19952,N_16533);
and U20819 (N_20819,N_17600,N_17822);
and U20820 (N_20820,N_17579,N_17501);
or U20821 (N_20821,N_17465,N_15735);
nand U20822 (N_20822,N_17634,N_16627);
and U20823 (N_20823,N_18537,N_19027);
xor U20824 (N_20824,N_17368,N_16278);
xnor U20825 (N_20825,N_17457,N_16703);
nand U20826 (N_20826,N_19785,N_19715);
nor U20827 (N_20827,N_18250,N_15121);
nand U20828 (N_20828,N_17738,N_18681);
xor U20829 (N_20829,N_18297,N_18653);
nor U20830 (N_20830,N_19052,N_16497);
or U20831 (N_20831,N_18780,N_17049);
or U20832 (N_20832,N_19299,N_18115);
xor U20833 (N_20833,N_15999,N_16508);
nand U20834 (N_20834,N_19195,N_19529);
xor U20835 (N_20835,N_19701,N_19132);
nand U20836 (N_20836,N_16510,N_17241);
or U20837 (N_20837,N_19728,N_17391);
nor U20838 (N_20838,N_17386,N_18151);
nand U20839 (N_20839,N_19566,N_18922);
or U20840 (N_20840,N_18114,N_18821);
or U20841 (N_20841,N_17189,N_15837);
nand U20842 (N_20842,N_19717,N_15587);
or U20843 (N_20843,N_15682,N_19602);
or U20844 (N_20844,N_19111,N_19490);
nor U20845 (N_20845,N_17880,N_18150);
xnor U20846 (N_20846,N_18298,N_16904);
nand U20847 (N_20847,N_18581,N_17844);
or U20848 (N_20848,N_15007,N_17878);
nor U20849 (N_20849,N_15197,N_19528);
or U20850 (N_20850,N_18219,N_19157);
and U20851 (N_20851,N_17117,N_16622);
and U20852 (N_20852,N_15470,N_17879);
nand U20853 (N_20853,N_17315,N_16841);
and U20854 (N_20854,N_16381,N_15671);
xnor U20855 (N_20855,N_19365,N_19249);
nand U20856 (N_20856,N_18670,N_19160);
nor U20857 (N_20857,N_19091,N_17099);
xnor U20858 (N_20858,N_15196,N_16178);
xnor U20859 (N_20859,N_16710,N_19822);
and U20860 (N_20860,N_17332,N_18874);
nand U20861 (N_20861,N_18222,N_17353);
or U20862 (N_20862,N_18677,N_15681);
and U20863 (N_20863,N_18065,N_15788);
nand U20864 (N_20864,N_16830,N_17925);
nand U20865 (N_20865,N_19844,N_15994);
and U20866 (N_20866,N_16978,N_15626);
xor U20867 (N_20867,N_15414,N_16453);
and U20868 (N_20868,N_17814,N_18217);
xor U20869 (N_20869,N_16119,N_16758);
and U20870 (N_20870,N_18340,N_19767);
and U20871 (N_20871,N_15473,N_17026);
xnor U20872 (N_20872,N_19949,N_18835);
and U20873 (N_20873,N_17535,N_19451);
nand U20874 (N_20874,N_15592,N_17023);
or U20875 (N_20875,N_15322,N_18886);
and U20876 (N_20876,N_15173,N_16426);
nor U20877 (N_20877,N_17149,N_18079);
xor U20878 (N_20878,N_17961,N_15041);
nor U20879 (N_20879,N_18781,N_16184);
nand U20880 (N_20880,N_16008,N_19734);
and U20881 (N_20881,N_17087,N_19215);
and U20882 (N_20882,N_18840,N_19831);
nand U20883 (N_20883,N_17230,N_17761);
nor U20884 (N_20884,N_18682,N_18965);
nor U20885 (N_20885,N_16293,N_16491);
nor U20886 (N_20886,N_18078,N_16672);
or U20887 (N_20887,N_17911,N_19829);
xor U20888 (N_20888,N_15289,N_17280);
and U20889 (N_20889,N_16720,N_17646);
or U20890 (N_20890,N_19291,N_15392);
nand U20891 (N_20891,N_15443,N_17832);
xor U20892 (N_20892,N_15534,N_15369);
nand U20893 (N_20893,N_15600,N_17351);
nand U20894 (N_20894,N_16048,N_15187);
nand U20895 (N_20895,N_18590,N_15666);
and U20896 (N_20896,N_18252,N_19495);
nand U20897 (N_20897,N_18433,N_17371);
or U20898 (N_20898,N_17895,N_15067);
and U20899 (N_20899,N_17438,N_19199);
or U20900 (N_20900,N_17359,N_19275);
and U20901 (N_20901,N_19217,N_18731);
or U20902 (N_20902,N_15199,N_19707);
nand U20903 (N_20903,N_19214,N_15814);
xor U20904 (N_20904,N_18002,N_19803);
xnor U20905 (N_20905,N_19333,N_18483);
nor U20906 (N_20906,N_17532,N_17996);
or U20907 (N_20907,N_19909,N_15843);
or U20908 (N_20908,N_19651,N_19773);
nand U20909 (N_20909,N_16198,N_16572);
and U20910 (N_20910,N_18042,N_19401);
or U20911 (N_20911,N_19750,N_19854);
and U20912 (N_20912,N_17985,N_19502);
nor U20913 (N_20913,N_17700,N_15346);
or U20914 (N_20914,N_15094,N_19918);
or U20915 (N_20915,N_16176,N_19415);
or U20916 (N_20916,N_19445,N_19804);
nand U20917 (N_20917,N_18905,N_16669);
and U20918 (N_20918,N_16352,N_19148);
or U20919 (N_20919,N_15825,N_16846);
xnor U20920 (N_20920,N_19908,N_19592);
xnor U20921 (N_20921,N_15559,N_15768);
nand U20922 (N_20922,N_18390,N_15337);
nor U20923 (N_20923,N_19796,N_17302);
nand U20924 (N_20924,N_15893,N_15653);
or U20925 (N_20925,N_16683,N_18959);
and U20926 (N_20926,N_19970,N_18456);
and U20927 (N_20927,N_17454,N_17341);
and U20928 (N_20928,N_19874,N_19693);
xor U20929 (N_20929,N_16545,N_17935);
xor U20930 (N_20930,N_19856,N_19457);
or U20931 (N_20931,N_19209,N_19895);
nor U20932 (N_20932,N_18084,N_17455);
nor U20933 (N_20933,N_16529,N_19390);
nor U20934 (N_20934,N_16739,N_15771);
xnor U20935 (N_20935,N_19372,N_17435);
xor U20936 (N_20936,N_15991,N_19357);
nand U20937 (N_20937,N_17183,N_16765);
nand U20938 (N_20938,N_18678,N_19436);
or U20939 (N_20939,N_18873,N_18413);
or U20940 (N_20940,N_18160,N_18925);
nand U20941 (N_20941,N_15431,N_15332);
and U20942 (N_20942,N_19892,N_19658);
nor U20943 (N_20943,N_16391,N_19615);
or U20944 (N_20944,N_18162,N_18981);
nand U20945 (N_20945,N_19443,N_15854);
or U20946 (N_20946,N_19960,N_18625);
nor U20947 (N_20947,N_15649,N_16469);
xor U20948 (N_20948,N_15774,N_18550);
nor U20949 (N_20949,N_19266,N_15309);
or U20950 (N_20950,N_19227,N_17138);
and U20951 (N_20951,N_17614,N_17192);
xor U20952 (N_20952,N_19980,N_17308);
and U20953 (N_20953,N_17207,N_19428);
or U20954 (N_20954,N_19362,N_19413);
and U20955 (N_20955,N_17616,N_18654);
or U20956 (N_20956,N_16085,N_19696);
xnor U20957 (N_20957,N_17337,N_17203);
nand U20958 (N_20958,N_15887,N_15229);
xor U20959 (N_20959,N_17035,N_17084);
nor U20960 (N_20960,N_17136,N_18066);
nand U20961 (N_20961,N_15767,N_18213);
and U20962 (N_20962,N_16255,N_19288);
or U20963 (N_20963,N_18141,N_16579);
nor U20964 (N_20964,N_18777,N_16421);
xor U20965 (N_20965,N_16123,N_18599);
or U20966 (N_20966,N_19632,N_17910);
and U20967 (N_20967,N_17724,N_16132);
and U20968 (N_20968,N_18901,N_16055);
or U20969 (N_20969,N_17611,N_18617);
nand U20970 (N_20970,N_15654,N_19265);
nor U20971 (N_20971,N_15435,N_17358);
or U20972 (N_20972,N_15420,N_16665);
or U20973 (N_20973,N_17725,N_18666);
nand U20974 (N_20974,N_16714,N_17623);
nor U20975 (N_20975,N_15135,N_19268);
nand U20976 (N_20976,N_17883,N_19627);
nand U20977 (N_20977,N_19412,N_17573);
nand U20978 (N_20978,N_16419,N_17365);
or U20979 (N_20979,N_17786,N_18882);
nand U20980 (N_20980,N_18720,N_19046);
nor U20981 (N_20981,N_15673,N_18069);
nand U20982 (N_20982,N_19698,N_19407);
nor U20983 (N_20983,N_19660,N_15646);
nand U20984 (N_20984,N_16521,N_17893);
or U20985 (N_20985,N_16222,N_18570);
and U20986 (N_20986,N_19568,N_18471);
and U20987 (N_20987,N_18984,N_19577);
nand U20988 (N_20988,N_19034,N_17525);
nor U20989 (N_20989,N_18063,N_19972);
nand U20990 (N_20990,N_17154,N_17370);
xnor U20991 (N_20991,N_17078,N_15474);
and U20992 (N_20992,N_16481,N_16103);
xnor U20993 (N_20993,N_17956,N_18358);
nand U20994 (N_20994,N_16361,N_15813);
or U20995 (N_20995,N_16188,N_15342);
and U20996 (N_20996,N_19948,N_19167);
or U20997 (N_20997,N_18536,N_18683);
or U20998 (N_20998,N_17445,N_19509);
or U20999 (N_20999,N_17781,N_15839);
and U21000 (N_21000,N_15327,N_18727);
and U21001 (N_21001,N_17336,N_16744);
nor U21002 (N_21002,N_15488,N_18010);
nand U21003 (N_21003,N_16398,N_16429);
xor U21004 (N_21004,N_18255,N_18257);
nor U21005 (N_21005,N_19464,N_16074);
xnor U21006 (N_21006,N_17595,N_15875);
and U21007 (N_21007,N_15550,N_15393);
xor U21008 (N_21008,N_19015,N_16916);
or U21009 (N_21009,N_16428,N_19305);
xnor U21010 (N_21010,N_18155,N_16417);
xor U21011 (N_21011,N_18973,N_15399);
nor U21012 (N_21012,N_18519,N_18120);
xnor U21013 (N_21013,N_19894,N_15251);
or U21014 (N_21014,N_15595,N_18923);
and U21015 (N_21015,N_15976,N_15006);
nand U21016 (N_21016,N_17683,N_15631);
nand U21017 (N_21017,N_17909,N_17001);
and U21018 (N_21018,N_18836,N_16302);
nand U21019 (N_21019,N_18122,N_15247);
xnor U21020 (N_21020,N_19927,N_17240);
and U21021 (N_21021,N_17098,N_15822);
or U21022 (N_21022,N_16163,N_18004);
or U21023 (N_21023,N_16362,N_17678);
or U21024 (N_21024,N_16065,N_15456);
or U21025 (N_21025,N_18129,N_17478);
nand U21026 (N_21026,N_15628,N_16970);
xor U21027 (N_21027,N_15359,N_19768);
nand U21028 (N_21028,N_17124,N_16270);
and U21029 (N_21029,N_18204,N_17627);
nor U21030 (N_21030,N_19188,N_19264);
and U21031 (N_21031,N_18939,N_18328);
nor U21032 (N_21032,N_16730,N_17123);
nand U21033 (N_21033,N_16885,N_15025);
or U21034 (N_21034,N_16174,N_17430);
nor U21035 (N_21035,N_18003,N_15065);
nand U21036 (N_21036,N_19298,N_16809);
or U21037 (N_21037,N_15493,N_16141);
or U21038 (N_21038,N_15520,N_17182);
xnor U21039 (N_21039,N_16899,N_18386);
nor U21040 (N_21040,N_18598,N_15018);
nor U21041 (N_21041,N_18716,N_19358);
and U21042 (N_21042,N_15630,N_18651);
and U21043 (N_21043,N_19004,N_15691);
xor U21044 (N_21044,N_15931,N_15201);
and U21045 (N_21045,N_18816,N_16500);
xor U21046 (N_21046,N_18072,N_18154);
or U21047 (N_21047,N_15464,N_17313);
xnor U21048 (N_21048,N_17852,N_16535);
or U21049 (N_21049,N_19915,N_15469);
or U21050 (N_21050,N_15868,N_19191);
xnor U21051 (N_21051,N_16984,N_15718);
nand U21052 (N_21052,N_16406,N_16004);
xor U21053 (N_21053,N_16842,N_19179);
or U21054 (N_21054,N_17389,N_18449);
nor U21055 (N_21055,N_19029,N_15396);
nor U21056 (N_21056,N_16544,N_16009);
nor U21057 (N_21057,N_19603,N_17345);
xnor U21058 (N_21058,N_17085,N_16166);
nor U21059 (N_21059,N_17585,N_17750);
nor U21060 (N_21060,N_18640,N_15188);
and U21061 (N_21061,N_19353,N_19084);
xor U21062 (N_21062,N_16153,N_17599);
xnor U21063 (N_21063,N_18800,N_16980);
xnor U21064 (N_21064,N_16386,N_19780);
and U21065 (N_21065,N_19891,N_16037);
nand U21066 (N_21066,N_19286,N_15812);
and U21067 (N_21067,N_16096,N_16480);
or U21068 (N_21068,N_19030,N_18623);
and U21069 (N_21069,N_17890,N_19066);
nor U21070 (N_21070,N_18008,N_16154);
and U21071 (N_21071,N_17706,N_19741);
or U21072 (N_21072,N_15816,N_18988);
nor U21073 (N_21073,N_18243,N_16664);
xor U21074 (N_21074,N_16763,N_17004);
or U21075 (N_21075,N_16764,N_18187);
nor U21076 (N_21076,N_18542,N_16443);
or U21077 (N_21077,N_16791,N_15020);
or U21078 (N_21078,N_18414,N_15727);
nor U21079 (N_21079,N_15557,N_15169);
xnor U21080 (N_21080,N_18168,N_19931);
nor U21081 (N_21081,N_15708,N_15753);
nor U21082 (N_21082,N_17330,N_15217);
xor U21083 (N_21083,N_15336,N_15779);
or U21084 (N_21084,N_19008,N_18380);
and U21085 (N_21085,N_17309,N_19400);
xnor U21086 (N_21086,N_19559,N_18022);
nor U21087 (N_21087,N_15182,N_17870);
or U21088 (N_21088,N_16438,N_17238);
and U21089 (N_21089,N_16482,N_15940);
nor U21090 (N_21090,N_17364,N_19083);
and U21091 (N_21091,N_18007,N_16859);
xor U21092 (N_21092,N_19089,N_17472);
nand U21093 (N_21093,N_15181,N_17949);
xnor U21094 (N_21094,N_17826,N_18387);
xnor U21095 (N_21095,N_16993,N_15356);
nand U21096 (N_21096,N_18710,N_17836);
nand U21097 (N_21097,N_18563,N_16081);
and U21098 (N_21098,N_19420,N_16699);
or U21099 (N_21099,N_16231,N_19879);
nor U21100 (N_21100,N_18996,N_16894);
nand U21101 (N_21101,N_18743,N_16385);
and U21102 (N_21102,N_15644,N_18708);
and U21103 (N_21103,N_15032,N_18552);
nor U21104 (N_21104,N_17859,N_16629);
and U21105 (N_21105,N_16636,N_15686);
or U21106 (N_21106,N_17732,N_17572);
and U21107 (N_21107,N_17924,N_15527);
or U21108 (N_21108,N_17639,N_15613);
nand U21109 (N_21109,N_19117,N_19145);
nand U21110 (N_21110,N_18843,N_17817);
nor U21111 (N_21111,N_19178,N_17888);
or U21112 (N_21112,N_19039,N_18159);
nand U21113 (N_21113,N_17065,N_17649);
xnor U21114 (N_21114,N_16109,N_19361);
nor U21115 (N_21115,N_16229,N_15547);
and U21116 (N_21116,N_15191,N_18673);
nor U21117 (N_21117,N_19113,N_18699);
nand U21118 (N_21118,N_17747,N_16193);
and U21119 (N_21119,N_16861,N_18663);
xor U21120 (N_21120,N_17723,N_16823);
xnor U21121 (N_21121,N_16021,N_17264);
xor U21122 (N_21122,N_18789,N_16410);
and U21123 (N_21123,N_16843,N_15504);
nor U21124 (N_21124,N_19967,N_15948);
nor U21125 (N_21125,N_17620,N_17981);
nand U21126 (N_21126,N_16439,N_16248);
and U21127 (N_21127,N_19426,N_19910);
xor U21128 (N_21128,N_18199,N_16729);
xnor U21129 (N_21129,N_16771,N_15853);
xor U21130 (N_21130,N_15498,N_18858);
or U21131 (N_21131,N_16321,N_15366);
nand U21132 (N_21132,N_15206,N_19580);
or U21133 (N_21133,N_18756,N_16050);
or U21134 (N_21134,N_17113,N_15071);
nor U21135 (N_21135,N_16604,N_15883);
and U21136 (N_21136,N_19452,N_16998);
and U21137 (N_21137,N_19057,N_15612);
nand U21138 (N_21138,N_19569,N_16454);
nor U21139 (N_21139,N_19670,N_16986);
and U21140 (N_21140,N_17740,N_16360);
nor U21141 (N_21141,N_18032,N_15546);
and U21142 (N_21142,N_16655,N_19205);
and U21143 (N_21143,N_18893,N_15800);
nand U21144 (N_21144,N_16952,N_15465);
nand U21145 (N_21145,N_16042,N_19110);
xor U21146 (N_21146,N_18895,N_15730);
nand U21147 (N_21147,N_17201,N_19712);
and U21148 (N_21148,N_18690,N_16808);
nor U21149 (N_21149,N_15572,N_19612);
or U21150 (N_21150,N_19255,N_16845);
nand U21151 (N_21151,N_19774,N_19736);
nor U21152 (N_21152,N_15325,N_18404);
xnor U21153 (N_21153,N_19797,N_16639);
nor U21154 (N_21154,N_18914,N_19071);
nor U21155 (N_21155,N_16640,N_18986);
xor U21156 (N_21156,N_18592,N_18144);
nand U21157 (N_21157,N_17191,N_19565);
xor U21158 (N_21158,N_18102,N_17357);
and U21159 (N_21159,N_18755,N_16523);
nand U21160 (N_21160,N_19727,N_16676);
nor U21161 (N_21161,N_15751,N_18500);
nand U21162 (N_21162,N_17521,N_18172);
and U21163 (N_21163,N_17428,N_19517);
nor U21164 (N_21164,N_18336,N_16610);
xor U21165 (N_21165,N_16444,N_15110);
or U21166 (N_21166,N_17407,N_16960);
or U21167 (N_21167,N_19103,N_17387);
nand U21168 (N_21168,N_16987,N_18011);
and U21169 (N_21169,N_19992,N_17629);
and U21170 (N_21170,N_18147,N_16475);
nand U21171 (N_21171,N_15848,N_19153);
or U21172 (N_21172,N_18313,N_17109);
xnor U21173 (N_21173,N_16335,N_15004);
xnor U21174 (N_21174,N_17398,N_19988);
and U21175 (N_21175,N_17779,N_19184);
nand U21176 (N_21176,N_16592,N_17794);
nor U21177 (N_21177,N_17417,N_16054);
or U21178 (N_21178,N_18535,N_19925);
nand U21179 (N_21179,N_15845,N_16091);
nand U21180 (N_21180,N_19001,N_19124);
xnor U21181 (N_21181,N_16131,N_16612);
xor U21182 (N_21182,N_18026,N_17193);
and U21183 (N_21183,N_19759,N_18793);
nor U21184 (N_21184,N_17275,N_18660);
nand U21185 (N_21185,N_15898,N_17829);
nand U21186 (N_21186,N_16256,N_17995);
nor U21187 (N_21187,N_16350,N_19772);
and U21188 (N_21188,N_19049,N_19343);
xnor U21189 (N_21189,N_16292,N_19604);
xor U21190 (N_21190,N_15002,N_15017);
nor U21191 (N_21191,N_18967,N_18107);
nor U21192 (N_21192,N_16558,N_16810);
nor U21193 (N_21193,N_17159,N_18103);
and U21194 (N_21194,N_18883,N_16974);
nand U21195 (N_21195,N_18903,N_19212);
and U21196 (N_21196,N_19582,N_17118);
nand U21197 (N_21197,N_15213,N_18029);
and U21198 (N_21198,N_17130,N_16527);
nand U21199 (N_21199,N_16268,N_16835);
and U21200 (N_21200,N_19746,N_15987);
or U21201 (N_21201,N_16057,N_16196);
or U21202 (N_21202,N_17079,N_19739);
and U21203 (N_21203,N_15040,N_17374);
xnor U21204 (N_21204,N_18124,N_16514);
xnor U21205 (N_21205,N_18181,N_19484);
xnor U21206 (N_21206,N_15731,N_19471);
xor U21207 (N_21207,N_17560,N_17446);
and U21208 (N_21208,N_18944,N_17795);
nor U21209 (N_21209,N_19300,N_19123);
and U21210 (N_21210,N_19763,N_18384);
nor U21211 (N_21211,N_18215,N_19985);
and U21212 (N_21212,N_17055,N_18021);
or U21213 (N_21213,N_19965,N_19163);
and U21214 (N_21214,N_17310,N_15037);
and U21215 (N_21215,N_16788,N_18341);
nand U21216 (N_21216,N_18504,N_15009);
or U21217 (N_21217,N_16208,N_16864);
nand U21218 (N_21218,N_19201,N_16179);
nand U21219 (N_21219,N_18487,N_19847);
or U21220 (N_21220,N_18373,N_16740);
nand U21221 (N_21221,N_18615,N_16887);
xnor U21222 (N_21222,N_19732,N_15762);
and U21223 (N_21223,N_15554,N_17544);
nand U21224 (N_21224,N_16713,N_19916);
or U21225 (N_21225,N_16857,N_15440);
or U21226 (N_21226,N_17249,N_16246);
or U21227 (N_21227,N_17536,N_15005);
nor U21228 (N_21228,N_17858,N_18478);
nor U21229 (N_21229,N_17233,N_15919);
xnor U21230 (N_21230,N_18806,N_19600);
xnor U21231 (N_21231,N_16064,N_16718);
nand U21232 (N_21232,N_16751,N_18951);
or U21233 (N_21233,N_19628,N_15755);
and U21234 (N_21234,N_19561,N_19544);
xor U21235 (N_21235,N_18618,N_18421);
nand U21236 (N_21236,N_16555,N_19730);
nand U21237 (N_21237,N_16377,N_16593);
nand U21238 (N_21238,N_16619,N_16441);
nor U21239 (N_21239,N_19754,N_15310);
or U21240 (N_21240,N_19811,N_18887);
nand U21241 (N_21241,N_17566,N_16063);
xor U21242 (N_21242,N_18401,N_16551);
nor U21243 (N_21243,N_16106,N_18244);
or U21244 (N_21244,N_15790,N_19817);
or U21245 (N_21245,N_17991,N_19441);
and U21246 (N_21246,N_16563,N_15157);
nand U21247 (N_21247,N_17297,N_17144);
nand U21248 (N_21248,N_16379,N_19876);
nor U21249 (N_21249,N_15761,N_16203);
or U21250 (N_21250,N_19537,N_17042);
or U21251 (N_21251,N_18912,N_19455);
or U21252 (N_21252,N_16253,N_18631);
nand U21253 (N_21253,N_17355,N_15882);
and U21254 (N_21254,N_18991,N_17270);
nand U21255 (N_21255,N_19086,N_19716);
or U21256 (N_21256,N_19691,N_18429);
nand U21257 (N_21257,N_17662,N_17591);
xnor U21258 (N_21258,N_16953,N_16155);
or U21259 (N_21259,N_16656,N_16090);
and U21260 (N_21260,N_19012,N_16346);
or U21261 (N_21261,N_19868,N_19751);
or U21262 (N_21262,N_19327,N_17091);
nor U21263 (N_21263,N_15338,N_19926);
xor U21264 (N_21264,N_17402,N_19747);
xnor U21265 (N_21265,N_15794,N_17675);
nand U21266 (N_21266,N_16586,N_18509);
and U21267 (N_21267,N_17451,N_16114);
or U21268 (N_21268,N_19017,N_15401);
and U21269 (N_21269,N_19674,N_15279);
nor U21270 (N_21270,N_17494,N_15057);
nand U21271 (N_21271,N_15036,N_17286);
xnor U21272 (N_21272,N_16645,N_15249);
nand U21273 (N_21273,N_15958,N_19596);
xor U21274 (N_21274,N_17190,N_16092);
nor U21275 (N_21275,N_15585,N_15367);
or U21276 (N_21276,N_15709,N_17293);
and U21277 (N_21277,N_15857,N_17644);
xnor U21278 (N_21278,N_19539,N_19519);
nand U21279 (N_21279,N_18310,N_15237);
xor U21280 (N_21280,N_17444,N_16601);
nand U21281 (N_21281,N_19482,N_19532);
xor U21282 (N_21282,N_15675,N_15148);
nand U21283 (N_21283,N_15102,N_18571);
nor U21284 (N_21284,N_18507,N_19667);
xor U21285 (N_21285,N_17376,N_18046);
xnor U21286 (N_21286,N_18301,N_16922);
and U21287 (N_21287,N_15743,N_17694);
and U21288 (N_21288,N_15522,N_19567);
nor U21289 (N_21289,N_18265,N_18499);
nand U21290 (N_21290,N_19648,N_18234);
xnor U21291 (N_21291,N_19440,N_15941);
and U21292 (N_21292,N_18964,N_16833);
or U21293 (N_21293,N_16286,N_15215);
or U21294 (N_21294,N_15615,N_16687);
nand U21295 (N_21295,N_16732,N_19896);
nor U21296 (N_21296,N_18794,N_17631);
nor U21297 (N_21297,N_15526,N_16447);
or U21298 (N_21298,N_19223,N_15260);
nor U21299 (N_21299,N_18524,N_16211);
nand U21300 (N_21300,N_15565,N_19825);
nor U21301 (N_21301,N_16084,N_15418);
nor U21302 (N_21302,N_17547,N_17783);
or U21303 (N_21303,N_18350,N_15328);
nor U21304 (N_21304,N_19722,N_17711);
or U21305 (N_21305,N_17565,N_19659);
nor U21306 (N_21306,N_15974,N_19943);
xor U21307 (N_21307,N_19366,N_18312);
and U21308 (N_21308,N_16577,N_16359);
nor U21309 (N_21309,N_15060,N_15287);
nand U21310 (N_21310,N_18034,N_17574);
nor U21311 (N_21311,N_16958,N_18724);
nor U21312 (N_21312,N_17311,N_19097);
and U21313 (N_21313,N_19647,N_15186);
nor U21314 (N_21314,N_18585,N_15457);
nor U21315 (N_21315,N_17603,N_17321);
nor U21316 (N_21316,N_17930,N_15639);
nand U21317 (N_21317,N_19541,N_19423);
nand U21318 (N_21318,N_19002,N_15570);
or U21319 (N_21319,N_18111,N_17606);
xor U21320 (N_21320,N_17259,N_19958);
and U21321 (N_21321,N_15139,N_18013);
or U21322 (N_21322,N_18894,N_18810);
and U21323 (N_21323,N_18484,N_19594);
xor U21324 (N_21324,N_17657,N_17677);
nor U21325 (N_21325,N_19700,N_16075);
xor U21326 (N_21326,N_18391,N_18077);
and U21327 (N_21327,N_18848,N_19617);
nor U21328 (N_21328,N_18299,N_15785);
or U21329 (N_21329,N_15792,N_19024);
nand U21330 (N_21330,N_15151,N_16624);
nand U21331 (N_21331,N_16143,N_19989);
xnor U21332 (N_21332,N_17481,N_18803);
or U21333 (N_21333,N_16975,N_18494);
and U21334 (N_21334,N_17760,N_16088);
and U21335 (N_21335,N_19663,N_19033);
or U21336 (N_21336,N_17645,N_17436);
and U21337 (N_21337,N_15165,N_16120);
and U21338 (N_21338,N_15300,N_16651);
and U21339 (N_21339,N_18572,N_19849);
or U21340 (N_21340,N_19213,N_15660);
and U21341 (N_21341,N_19953,N_17522);
or U21342 (N_21342,N_16585,N_19375);
nand U21343 (N_21343,N_18479,N_16728);
or U21344 (N_21344,N_17577,N_19500);
nand U21345 (N_21345,N_19450,N_17304);
nand U21346 (N_21346,N_18672,N_17393);
or U21347 (N_21347,N_15564,N_17588);
xnor U21348 (N_21348,N_18723,N_16446);
nand U21349 (N_21349,N_19120,N_18930);
xor U21350 (N_21350,N_17821,N_19758);
and U21351 (N_21351,N_17993,N_18100);
and U21352 (N_21352,N_17146,N_16856);
and U21353 (N_21353,N_17060,N_17348);
nand U21354 (N_21354,N_17745,N_15083);
nor U21355 (N_21355,N_16675,N_15511);
xnor U21356 (N_21356,N_18269,N_15583);
and U21357 (N_21357,N_17543,N_16883);
xor U21358 (N_21358,N_18191,N_19671);
nand U21359 (N_21359,N_19591,N_18071);
xor U21360 (N_21360,N_19756,N_17828);
nand U21361 (N_21361,N_17169,N_19023);
nor U21362 (N_21362,N_19261,N_18268);
nand U21363 (N_21363,N_15131,N_15802);
nor U21364 (N_21364,N_17167,N_15548);
nor U21365 (N_21365,N_15589,N_17697);
nor U21366 (N_21366,N_15314,N_19170);
xor U21367 (N_21367,N_16648,N_16757);
and U21368 (N_21368,N_19654,N_17403);
or U21369 (N_21369,N_17245,N_18322);
nor U21370 (N_21370,N_16574,N_17647);
xor U21371 (N_21371,N_16957,N_19536);
nor U21372 (N_21372,N_18481,N_19575);
and U21373 (N_21373,N_15978,N_19890);
or U21374 (N_21374,N_17871,N_18043);
or U21375 (N_21375,N_17969,N_17799);
or U21376 (N_21376,N_15963,N_19636);
or U21377 (N_21377,N_16948,N_16171);
xor U21378 (N_21378,N_17685,N_15363);
and U21379 (N_21379,N_16289,N_16380);
xor U21380 (N_21380,N_16234,N_16394);
nand U21381 (N_21381,N_18467,N_19391);
nand U21382 (N_21382,N_19823,N_17850);
nand U21383 (N_21383,N_17530,N_17846);
xnor U21384 (N_21384,N_16561,N_18118);
xor U21385 (N_21385,N_16897,N_15732);
and U21386 (N_21386,N_19828,N_17155);
nor U21387 (N_21387,N_17802,N_17602);
or U21388 (N_21388,N_19256,N_17768);
and U21389 (N_21389,N_15184,N_15471);
nand U21390 (N_21390,N_15750,N_19638);
xnor U21391 (N_21391,N_16390,N_16030);
or U21392 (N_21392,N_19403,N_18508);
or U21393 (N_21393,N_19102,N_15339);
xnor U21394 (N_21394,N_16431,N_18943);
xor U21395 (N_21395,N_19606,N_15684);
nor U21396 (N_21396,N_15221,N_15115);
nor U21397 (N_21397,N_19929,N_17224);
xor U21398 (N_21398,N_18016,N_15194);
or U21399 (N_21399,N_15290,N_16496);
and U21400 (N_21400,N_15164,N_16828);
and U21401 (N_21401,N_18171,N_15849);
xor U21402 (N_21402,N_18207,N_16317);
nor U21403 (N_21403,N_18807,N_19695);
or U21404 (N_21404,N_16512,N_16745);
nand U21405 (N_21405,N_17058,N_19025);
and U21406 (N_21406,N_18253,N_17946);
nand U21407 (N_21407,N_17331,N_15095);
nand U21408 (N_21408,N_17448,N_15690);
xor U21409 (N_21409,N_19510,N_19044);
and U21410 (N_21410,N_15773,N_16373);
or U21411 (N_21411,N_15253,N_18041);
and U21412 (N_21412,N_15988,N_15637);
or U21413 (N_21413,N_15202,N_17132);
xor U21414 (N_21414,N_17031,N_17538);
or U21415 (N_21415,N_16269,N_17415);
or U21416 (N_21416,N_15993,N_18601);
xor U21417 (N_21417,N_19713,N_17927);
or U21418 (N_21418,N_17806,N_19467);
nor U21419 (N_21419,N_16852,N_16822);
nor U21420 (N_21420,N_16829,N_19725);
xor U21421 (N_21421,N_16660,N_15805);
nor U21422 (N_21422,N_15677,N_16569);
or U21423 (N_21423,N_17965,N_18880);
xor U21424 (N_21424,N_15679,N_17424);
xor U21425 (N_21425,N_17719,N_19787);
or U21426 (N_21426,N_19572,N_17643);
and U21427 (N_21427,N_18052,N_18954);
and U21428 (N_21428,N_17987,N_17088);
and U21429 (N_21429,N_18435,N_19998);
nor U21430 (N_21430,N_17637,N_16921);
nand U21431 (N_21431,N_17851,N_16706);
nor U21432 (N_21432,N_17673,N_16059);
nand U21433 (N_21433,N_15552,N_17608);
and U21434 (N_21434,N_16374,N_18202);
xnor U21435 (N_21435,N_19878,N_18918);
nand U21436 (N_21436,N_16014,N_15964);
xor U21437 (N_21437,N_15116,N_19211);
xor U21438 (N_21438,N_17749,N_15483);
and U21439 (N_21439,N_19219,N_16486);
nand U21440 (N_21440,N_17307,N_18206);
xor U21441 (N_21441,N_17422,N_18410);
or U21442 (N_21442,N_17651,N_16618);
nor U21443 (N_21443,N_18031,N_19054);
or U21444 (N_21444,N_15778,N_18597);
or U21445 (N_21445,N_19112,N_16507);
and U21446 (N_21446,N_17612,N_15847);
or U21447 (N_21447,N_16073,N_17213);
xor U21448 (N_21448,N_19599,N_17978);
nor U21449 (N_21449,N_19640,N_16513);
or U21450 (N_21450,N_16663,N_17054);
nor U21451 (N_21451,N_18997,N_17342);
nand U21452 (N_21452,N_19619,N_17720);
xnor U21453 (N_21453,N_16694,N_17426);
nand U21454 (N_21454,N_17102,N_19292);
xor U21455 (N_21455,N_15832,N_18028);
and U21456 (N_21456,N_16522,N_16467);
xor U21457 (N_21457,N_16511,N_16122);
nor U21458 (N_21458,N_19277,N_17979);
nand U21459 (N_21459,N_17225,N_17408);
nor U21460 (N_21460,N_17681,N_18036);
nand U21461 (N_21461,N_15096,N_18513);
and U21462 (N_21462,N_18001,N_15158);
nor U21463 (N_21463,N_15238,N_19239);
or U21464 (N_21464,N_19315,N_16961);
xnor U21465 (N_21465,N_17458,N_19607);
nand U21466 (N_21466,N_18695,N_16227);
or U21467 (N_21467,N_18502,N_18379);
or U21468 (N_21468,N_18024,N_15326);
and U21469 (N_21469,N_15298,N_18082);
and U21470 (N_21470,N_19313,N_18075);
xnor U21471 (N_21471,N_16332,N_18368);
xor U21472 (N_21472,N_16281,N_15478);
and U21473 (N_21473,N_17654,N_16060);
xnor U21474 (N_21474,N_16983,N_18884);
nand U21475 (N_21475,N_19381,N_17373);
nand U21476 (N_21476,N_16102,N_19870);
nor U21477 (N_21477,N_19062,N_18241);
and U21478 (N_21478,N_17413,N_19959);
nand U21479 (N_21479,N_19543,N_16976);
nor U21480 (N_21480,N_17835,N_16232);
and U21481 (N_21481,N_15054,N_18860);
or U21482 (N_21482,N_17253,N_18776);
or U21483 (N_21483,N_16893,N_17917);
nor U21484 (N_21484,N_16580,N_19055);
and U21485 (N_21485,N_19363,N_15977);
and U21486 (N_21486,N_15130,N_15820);
xnor U21487 (N_21487,N_19104,N_15345);
nand U21488 (N_21488,N_18314,N_19542);
xnor U21489 (N_21489,N_15372,N_18258);
nor U21490 (N_21490,N_17188,N_16657);
xnor U21491 (N_21491,N_18888,N_19414);
nor U21492 (N_21492,N_17263,N_15239);
or U21493 (N_21493,N_18169,N_18838);
xor U21494 (N_21494,N_16776,N_16568);
or U21495 (N_21495,N_18904,N_15451);
nor U21496 (N_21496,N_16207,N_18657);
xor U21497 (N_21497,N_17664,N_17780);
and U21498 (N_21498,N_19011,N_19883);
nand U21499 (N_21499,N_19845,N_18566);
nor U21500 (N_21500,N_18080,N_18093);
xnor U21501 (N_21501,N_19905,N_19497);
or U21502 (N_21502,N_15231,N_17232);
nor U21503 (N_21503,N_18420,N_18407);
nor U21504 (N_21504,N_17648,N_19309);
and U21505 (N_21505,N_16324,N_18885);
nor U21506 (N_21506,N_19462,N_17754);
or U21507 (N_21507,N_15687,N_16662);
and U21508 (N_21508,N_16363,N_16223);
and U21509 (N_21509,N_19065,N_18545);
xnor U21510 (N_21510,N_16309,N_19501);
xor U21511 (N_21511,N_15398,N_18999);
or U21512 (N_21512,N_17456,N_17908);
xnor U21513 (N_21513,N_19511,N_18472);
or U21514 (N_21514,N_17170,N_18259);
nor U21515 (N_21515,N_19809,N_19766);
and U21516 (N_21516,N_16052,N_15970);
or U21517 (N_21517,N_15195,N_15426);
nor U21518 (N_21518,N_15049,N_17605);
and U21519 (N_21519,N_19425,N_15444);
or U21520 (N_21520,N_16766,N_18960);
and U21521 (N_21521,N_17427,N_17255);
xor U21522 (N_21522,N_18924,N_18758);
and U21523 (N_21523,N_16464,N_16752);
nand U21524 (N_21524,N_16288,N_16413);
nand U21525 (N_21525,N_16192,N_17976);
or U21526 (N_21526,N_18796,N_18795);
or U21527 (N_21527,N_15246,N_16679);
and U21528 (N_21528,N_16940,N_16855);
and U21529 (N_21529,N_17206,N_18271);
nor U21530 (N_21530,N_15044,N_17476);
nor U21531 (N_21531,N_17958,N_18892);
xor U21532 (N_21532,N_15143,N_18152);
and U21533 (N_21533,N_15098,N_16145);
nor U21534 (N_21534,N_19152,N_19808);
xnor U21535 (N_21535,N_18125,N_17467);
nand U21536 (N_21536,N_18044,N_17097);
nor U21537 (N_21537,N_18388,N_18148);
nand U21538 (N_21538,N_18900,N_18040);
xnor U21539 (N_21539,N_15864,N_16007);
nor U21540 (N_21540,N_16035,N_15872);
or U21541 (N_21541,N_19161,N_19578);
or U21542 (N_21542,N_17622,N_17874);
and U21543 (N_21543,N_17020,N_15216);
nor U21544 (N_21544,N_16329,N_16283);
nor U21545 (N_21545,N_19439,N_17701);
nand U21546 (N_21546,N_17411,N_18648);
nand U21547 (N_21547,N_16459,N_19246);
nor U21548 (N_21548,N_16182,N_17361);
nor U21549 (N_21549,N_17942,N_15035);
nand U21550 (N_21550,N_19010,N_15090);
xor U21551 (N_21551,N_16853,N_16504);
xor U21552 (N_21552,N_18354,N_15362);
nor U21553 (N_21553,N_16080,N_18686);
and U21554 (N_21554,N_16026,N_17504);
nand U21555 (N_21555,N_16915,N_17260);
xnor U21556 (N_21556,N_18611,N_15394);
nor U21557 (N_21557,N_17894,N_18378);
or U21558 (N_21558,N_18276,N_18588);
xor U21559 (N_21559,N_15286,N_15232);
or U21560 (N_21560,N_15042,N_19718);
or U21561 (N_21561,N_19175,N_17571);
and U21562 (N_21562,N_15302,N_15744);
nor U21563 (N_21563,N_16185,N_18248);
xor U21564 (N_21564,N_19067,N_15551);
nand U21565 (N_21565,N_16724,N_15000);
nand U21566 (N_21566,N_18216,N_15378);
nand U21567 (N_21567,N_17092,N_16966);
or U21568 (N_21568,N_16524,N_17100);
nand U21569 (N_21569,N_18189,N_15703);
nor U21570 (N_21570,N_15803,N_17112);
or U21571 (N_21571,N_17134,N_17955);
nand U21572 (N_21572,N_15167,N_18135);
nand U21573 (N_21573,N_19159,N_19099);
or U21574 (N_21574,N_19310,N_18725);
nor U21575 (N_21575,N_19346,N_19202);
nand U21576 (N_21576,N_17334,N_16602);
and U21577 (N_21577,N_16015,N_16690);
nand U21578 (N_21578,N_19427,N_15961);
nor U21579 (N_21579,N_17943,N_15723);
or U21580 (N_21580,N_17380,N_18432);
and U21581 (N_21581,N_18182,N_15953);
nand U21582 (N_21582,N_19790,N_18119);
and U21583 (N_21583,N_17913,N_18178);
xor U21584 (N_21584,N_18146,N_16023);
xor U21585 (N_21585,N_18603,N_17071);
xnor U21586 (N_21586,N_19902,N_16565);
xnor U21587 (N_21587,N_15650,N_16437);
nand U21588 (N_21588,N_17209,N_18416);
xor U21589 (N_21589,N_16111,N_19323);
nand U21590 (N_21590,N_16628,N_15204);
nor U21591 (N_21591,N_17770,N_18142);
and U21592 (N_21592,N_15087,N_15507);
nand U21593 (N_21593,N_15124,N_17636);
nand U21594 (N_21594,N_17414,N_18679);
xor U21595 (N_21595,N_19041,N_17753);
and U21596 (N_21596,N_15224,N_17630);
nor U21597 (N_21597,N_17746,N_18517);
or U21598 (N_21598,N_18910,N_17970);
nand U21599 (N_21599,N_19252,N_19846);
or U21600 (N_21600,N_16528,N_16079);
xnor U21601 (N_21601,N_17800,N_17290);
or U21602 (N_21602,N_17804,N_16723);
xor U21603 (N_21603,N_19154,N_17517);
nand U21604 (N_21604,N_19714,N_18501);
xor U21605 (N_21605,N_17818,N_18824);
nor U21606 (N_21606,N_19491,N_15161);
nor U21607 (N_21607,N_15370,N_15714);
or U21608 (N_21608,N_15693,N_18637);
or U21609 (N_21609,N_16403,N_19282);
nand U21610 (N_21610,N_19138,N_19454);
nand U21611 (N_21611,N_19776,N_19013);
xnor U21612 (N_21612,N_17298,N_15486);
nor U21613 (N_21613,N_17548,N_18929);
nand U21614 (N_21614,N_16571,N_16888);
and U21615 (N_21615,N_15357,N_19442);
xor U21616 (N_21616,N_15097,N_19351);
nor U21617 (N_21617,N_15235,N_17503);
xnor U21618 (N_21618,N_15416,N_17452);
nor U21619 (N_21619,N_15063,N_15683);
nor U21620 (N_21620,N_19950,N_17816);
nor U21621 (N_21621,N_19135,N_18898);
xor U21622 (N_21622,N_17597,N_18953);
nor U21623 (N_21623,N_16704,N_18180);
xor U21624 (N_21624,N_16121,N_18747);
or U21625 (N_21625,N_16789,N_15448);
nor U21626 (N_21626,N_16165,N_18318);
xor U21627 (N_21627,N_15320,N_16432);
xor U21628 (N_21628,N_15447,N_17542);
nor U21629 (N_21629,N_19922,N_19192);
and U21630 (N_21630,N_15051,N_18455);
xor U21631 (N_21631,N_18194,N_16708);
xor U21632 (N_21632,N_19449,N_15640);
nor U21633 (N_21633,N_16033,N_19588);
nand U21634 (N_21634,N_16999,N_19848);
nor U21635 (N_21635,N_16420,N_15985);
nor U21636 (N_21636,N_19274,N_15890);
xor U21637 (N_21637,N_16783,N_17122);
or U21638 (N_21638,N_18174,N_18994);
nand U21639 (N_21639,N_17312,N_19656);
or U21640 (N_21640,N_15028,N_19518);
nor U21641 (N_21641,N_17074,N_17172);
nand U21642 (N_21642,N_16484,N_18701);
nand U21643 (N_21643,N_19563,N_18267);
and U21644 (N_21644,N_17346,N_16264);
nand U21645 (N_21645,N_17498,N_18772);
nand U21646 (N_21646,N_16546,N_15268);
xnor U21647 (N_21647,N_17491,N_15284);
and U21648 (N_21648,N_19597,N_18280);
nand U21649 (N_21649,N_16213,N_19289);
xor U21650 (N_21650,N_19688,N_16397);
and U21651 (N_21651,N_15834,N_15950);
nor U21652 (N_21652,N_16692,N_15502);
nand U21653 (N_21653,N_18966,N_16219);
nor U21654 (N_21654,N_17016,N_16461);
nor U21655 (N_21655,N_17050,N_17265);
nor U21656 (N_21656,N_19468,N_17788);
xor U21657 (N_21657,N_18278,N_19810);
or U21658 (N_21658,N_18218,N_18814);
nor U21659 (N_21659,N_18344,N_16382);
or U21660 (N_21660,N_17107,N_17617);
and U21661 (N_21661,N_17236,N_17690);
or U21662 (N_21662,N_15634,N_15190);
and U21663 (N_21663,N_16784,N_15594);
or U21664 (N_21664,N_19784,N_16056);
xnor U21665 (N_21665,N_18091,N_15742);
or U21666 (N_21666,N_18188,N_15915);
and U21667 (N_21667,N_16797,N_15210);
or U21668 (N_21668,N_18375,N_17388);
nand U21669 (N_21669,N_17468,N_17377);
nand U21670 (N_21670,N_18974,N_19254);
nand U21671 (N_21671,N_19893,N_18060);
nor U21672 (N_21672,N_16356,N_18185);
nand U21673 (N_21673,N_19287,N_19051);
and U21674 (N_21674,N_19245,N_18382);
xnor U21675 (N_21675,N_15430,N_15616);
nand U21676 (N_21676,N_18099,N_16674);
or U21677 (N_21677,N_16415,N_17615);
nand U21678 (N_21678,N_17824,N_16226);
and U21679 (N_21679,N_15120,N_19966);
nand U21680 (N_21680,N_15159,N_16215);
and U21681 (N_21681,N_18850,N_18712);
or U21682 (N_21682,N_17128,N_15296);
and U21683 (N_21683,N_19903,N_17333);
nor U21684 (N_21684,N_19279,N_16247);
and U21685 (N_21685,N_18409,N_17229);
nor U21686 (N_21686,N_19898,N_15107);
nor U21687 (N_21687,N_18233,N_17854);
and U21688 (N_21688,N_15147,N_19225);
xor U21689 (N_21689,N_16920,N_15468);
nor U21690 (N_21690,N_15942,N_16862);
nand U21691 (N_21691,N_19935,N_19146);
nand U21692 (N_21692,N_15402,N_19331);
and U21693 (N_21693,N_15609,N_17486);
nand U21694 (N_21694,N_19382,N_17731);
nor U21695 (N_21695,N_17447,N_18443);
and U21696 (N_21696,N_18453,N_18498);
or U21697 (N_21697,N_16237,N_19116);
and U21698 (N_21698,N_17717,N_17782);
nand U21699 (N_21699,N_18229,N_19340);
nand U21700 (N_21700,N_18133,N_19475);
nor U21701 (N_21701,N_18197,N_15144);
or U21702 (N_21702,N_16404,N_17847);
xnor U21703 (N_21703,N_18279,N_15295);
xnor U21704 (N_21704,N_18558,N_15455);
nand U21705 (N_21705,N_17714,N_18329);
nand U21706 (N_21706,N_17433,N_18839);
and U21707 (N_21707,N_16654,N_15439);
xor U21708 (N_21708,N_18579,N_18326);
nor U21709 (N_21709,N_17360,N_16044);
nand U21710 (N_21710,N_18574,N_19917);
or U21711 (N_21711,N_18076,N_19140);
nand U21712 (N_21712,N_16100,N_17247);
nand U21713 (N_21713,N_17576,N_17228);
and U21714 (N_21714,N_17412,N_16104);
nand U21715 (N_21715,N_16239,N_16520);
nand U21716 (N_21716,N_16087,N_19655);
or U21717 (N_21717,N_18515,N_16734);
nor U21718 (N_21718,N_19646,N_15869);
nand U21719 (N_21719,N_16792,N_19079);
and U21720 (N_21720,N_19101,N_19994);
or U21721 (N_21721,N_19686,N_15503);
or U21722 (N_21722,N_19681,N_17056);
nor U21723 (N_21723,N_15101,N_17589);
or U21724 (N_21724,N_18113,N_19835);
nor U21725 (N_21725,N_18630,N_15458);
xnor U21726 (N_21726,N_16369,N_17772);
or U21727 (N_21727,N_16768,N_18196);
nand U21728 (N_21728,N_19624,N_17903);
or U21729 (N_21729,N_15581,N_18962);
nor U21730 (N_21730,N_18562,N_18062);
nand U21731 (N_21731,N_19472,N_19499);
nor U21732 (N_21732,N_19059,N_18287);
xnor U21733 (N_21733,N_17709,N_17672);
nand U21734 (N_21734,N_17153,N_17568);
and U21735 (N_21735,N_15965,N_16688);
and U21736 (N_21736,N_16620,N_16312);
nor U21737 (N_21737,N_19906,N_19945);
and U21738 (N_21738,N_16476,N_15586);
nand U21739 (N_21739,N_16127,N_18047);
and U21740 (N_21740,N_17945,N_17340);
nand U21741 (N_21741,N_16220,N_15409);
nand U21742 (N_21742,N_15661,N_18644);
xnor U21743 (N_21743,N_16509,N_16449);
and U21744 (N_21744,N_17303,N_19888);
nand U21745 (N_21745,N_16534,N_19682);
nand U21746 (N_21746,N_18849,N_17509);
and U21747 (N_21747,N_18411,N_17090);
nor U21748 (N_21748,N_18577,N_18235);
nand U21749 (N_21749,N_18902,N_17317);
nand U21750 (N_21750,N_17559,N_15433);
or U21751 (N_21751,N_18321,N_15269);
nor U21752 (N_21752,N_16996,N_15900);
and U21753 (N_21753,N_19900,N_18872);
nor U21754 (N_21754,N_16310,N_19312);
or U21755 (N_21755,N_19863,N_19533);
or U21756 (N_21756,N_17404,N_15670);
or U21757 (N_21757,N_17257,N_15198);
or U21758 (N_21758,N_18911,N_16539);
or U21759 (N_21759,N_17881,N_18926);
xnor U21760 (N_21760,N_17593,N_18854);
xor U21761 (N_21761,N_19947,N_16212);
nand U21762 (N_21762,N_18170,N_17394);
nand U21763 (N_21763,N_16452,N_15062);
and U21764 (N_21764,N_15082,N_16142);
nor U21765 (N_21765,N_15856,N_19762);
or U21766 (N_21766,N_15404,N_18284);
or U21767 (N_21767,N_17633,N_16436);
and U21768 (N_21768,N_15509,N_15967);
or U21769 (N_21769,N_17953,N_17039);
or U21770 (N_21770,N_15576,N_18532);
nand U21771 (N_21771,N_17691,N_15747);
and U21772 (N_21772,N_16330,N_16796);
xor U21773 (N_21773,N_18116,N_16082);
nor U21774 (N_21774,N_19672,N_15799);
or U21775 (N_21775,N_19859,N_16787);
nand U21776 (N_21776,N_16774,N_15932);
xnor U21777 (N_21777,N_17972,N_17533);
or U21778 (N_21778,N_15177,N_15819);
nand U21779 (N_21779,N_16083,N_17912);
and U21780 (N_21780,N_17473,N_16964);
nor U21781 (N_21781,N_16098,N_19779);
nor U21782 (N_21782,N_16093,N_17655);
or U21783 (N_21783,N_17752,N_15861);
or U21784 (N_21784,N_18580,N_17736);
nand U21785 (N_21785,N_17076,N_19850);
or U21786 (N_21786,N_19940,N_19678);
and U21787 (N_21787,N_16644,N_19235);
xor U21788 (N_21788,N_19643,N_18808);
and U21789 (N_21789,N_15085,N_18694);
or U21790 (N_21790,N_17499,N_19576);
and U21791 (N_21791,N_18878,N_15829);
and U21792 (N_21792,N_17395,N_18638);
nor U21793 (N_21793,N_15984,N_17663);
nand U21794 (N_21794,N_16427,N_15011);
and U21795 (N_21795,N_15460,N_17581);
or U21796 (N_21796,N_17707,N_18346);
or U21797 (N_21797,N_15998,N_15611);
nor U21798 (N_21798,N_18014,N_16473);
xnor U21799 (N_21799,N_16468,N_17409);
nor U21800 (N_21800,N_18949,N_18068);
and U21801 (N_21801,N_18523,N_19141);
nor U21802 (N_21802,N_16311,N_19005);
or U21803 (N_21803,N_19740,N_19882);
or U21804 (N_21804,N_19379,N_15066);
xor U21805 (N_21805,N_17165,N_15117);
or U21806 (N_21806,N_19037,N_17204);
nand U21807 (N_21807,N_18817,N_16001);
or U21808 (N_21808,N_15694,N_19778);
or U21809 (N_21809,N_15740,N_16681);
or U21810 (N_21810,N_17053,N_17778);
nand U21811 (N_21811,N_19133,N_17862);
nand U21812 (N_21812,N_16733,N_17557);
xnor U21813 (N_21813,N_16349,N_18750);
nand U21814 (N_21814,N_17327,N_18104);
xor U21815 (N_21815,N_17984,N_16197);
and U21816 (N_21816,N_19485,N_16251);
or U21817 (N_21817,N_15842,N_16985);
nor U21818 (N_21818,N_19853,N_15906);
or U21819 (N_21819,N_15425,N_17222);
and U21820 (N_21820,N_18033,N_17237);
xor U21821 (N_21821,N_15846,N_18058);
or U21822 (N_21822,N_17142,N_18377);
nor U21823 (N_21823,N_15072,N_17196);
nand U21824 (N_21824,N_15688,N_19553);
or U21825 (N_21825,N_19858,N_15949);
and U21826 (N_21826,N_15668,N_17613);
nor U21827 (N_21827,N_18693,N_15692);
nor U21828 (N_21828,N_18877,N_15031);
or U21829 (N_21829,N_15874,N_16837);
or U21830 (N_21830,N_15489,N_19316);
xor U21831 (N_21831,N_17974,N_15168);
or U21832 (N_21832,N_19075,N_15817);
and U21833 (N_21833,N_17546,N_17181);
nand U21834 (N_21834,N_15306,N_15308);
xor U21835 (N_21835,N_19458,N_18527);
nand U21836 (N_21836,N_19410,N_19623);
nor U21837 (N_21837,N_17756,N_17066);
and U21838 (N_21838,N_16202,N_18496);
or U21839 (N_21839,N_15467,N_18506);
nor U21840 (N_21840,N_15261,N_15607);
nand U21841 (N_21841,N_19642,N_15333);
and U21842 (N_21842,N_16954,N_17179);
nor U21843 (N_21843,N_15863,N_16089);
nand U21844 (N_21844,N_16968,N_18460);
xnor U21845 (N_21845,N_15597,N_18715);
or U21846 (N_21846,N_19397,N_19392);
xnor U21847 (N_21847,N_19465,N_18097);
nor U21848 (N_21848,N_17289,N_16813);
nand U21849 (N_21849,N_19035,N_15763);
xor U21850 (N_21850,N_16932,N_18220);
nor U21851 (N_21851,N_18583,N_18254);
nor U21852 (N_21852,N_18112,N_15288);
nor U21853 (N_21853,N_16715,N_19587);
nor U21854 (N_21854,N_17150,N_16621);
and U21855 (N_21855,N_18395,N_19991);
or U21856 (N_21856,N_16726,N_18465);
nand U21857 (N_21857,N_19082,N_17601);
and U21858 (N_21858,N_19534,N_19073);
xor U21859 (N_21859,N_18242,N_17704);
or U21860 (N_21860,N_17938,N_18049);
nor U21861 (N_21861,N_18940,N_17372);
nand U21862 (N_21862,N_15275,N_15218);
or U21863 (N_21863,N_17869,N_17776);
or U21864 (N_21864,N_18127,N_16898);
and U21865 (N_21865,N_19836,N_15045);
or U21866 (N_21866,N_15870,N_16414);
xor U21867 (N_21867,N_19422,N_19743);
nor U21868 (N_21868,N_15620,N_17947);
nor U21869 (N_21869,N_15283,N_18546);
xnor U21870 (N_21870,N_16036,N_15537);
and U21871 (N_21871,N_18869,N_19889);
or U21872 (N_21872,N_19752,N_18928);
and U21873 (N_21873,N_15163,N_17495);
and U21874 (N_21874,N_17278,N_18826);
or U21875 (N_21875,N_16825,N_19294);
nand U21876 (N_21876,N_17737,N_17841);
nor U21877 (N_21877,N_15756,N_17784);
xor U21878 (N_21878,N_18769,N_18303);
and U21879 (N_21879,N_17743,N_16939);
nor U21880 (N_21880,N_17366,N_19862);
or U21881 (N_21881,N_19021,N_16387);
or U21882 (N_21882,N_19461,N_16671);
nand U21883 (N_21883,N_19134,N_18260);
and U21884 (N_21884,N_19308,N_19284);
and U21885 (N_21885,N_19978,N_16516);
xor U21886 (N_21886,N_17121,N_18622);
nor U21887 (N_21887,N_17963,N_18285);
nor U21888 (N_21888,N_16700,N_15220);
or U21889 (N_21889,N_16583,N_16515);
and U21890 (N_21890,N_19652,N_19523);
xor U21891 (N_21891,N_16407,N_19118);
and U21892 (N_21892,N_15775,N_17272);
xor U21893 (N_21893,N_18719,N_15280);
xor U21894 (N_21894,N_18430,N_17081);
and U21895 (N_21895,N_17015,N_17276);
or U21896 (N_21896,N_15770,N_17344);
xnor U21897 (N_21897,N_15685,N_17419);
or U21898 (N_21898,N_19127,N_19070);
xnor U21899 (N_21899,N_15015,N_16017);
nand U21900 (N_21900,N_18454,N_16412);
and U21901 (N_21901,N_18371,N_15982);
or U21902 (N_21902,N_16285,N_16638);
and U21903 (N_21903,N_18475,N_16737);
and U21904 (N_21904,N_18907,N_18149);
and U21905 (N_21905,N_17025,N_16680);
nand U21906 (N_21906,N_16194,N_17775);
or U21907 (N_21907,N_19733,N_15749);
and U21908 (N_21908,N_15705,N_17453);
xnor U21909 (N_21909,N_19815,N_15185);
xor U21910 (N_21910,N_15506,N_15189);
or U21911 (N_21911,N_16175,N_19253);
and U21912 (N_21912,N_15823,N_15664);
or U21913 (N_21913,N_15716,N_17195);
and U21914 (N_21914,N_15462,N_17111);
and U21915 (N_21915,N_16045,N_17916);
nor U21916 (N_21916,N_19007,N_15913);
nor U21917 (N_21917,N_19699,N_17899);
nor U21918 (N_21918,N_19290,N_19109);
and U21919 (N_21919,N_18470,N_19852);
xor U21920 (N_21920,N_19571,N_15981);
nor U21921 (N_21921,N_17967,N_17019);
xor U21922 (N_21922,N_18394,N_18296);
or U21923 (N_21923,N_15917,N_18855);
nor U21924 (N_21924,N_16517,N_15250);
nand U21925 (N_21925,N_16884,N_16071);
nand U21926 (N_21926,N_17385,N_19521);
and U21927 (N_21927,N_19814,N_15927);
or U21928 (N_21928,N_19630,N_19204);
or U21929 (N_21929,N_17977,N_18306);
xor U21930 (N_21930,N_19639,N_15574);
nor U21931 (N_21931,N_18511,N_15523);
or U21932 (N_21932,N_19911,N_17202);
and U21933 (N_21933,N_18779,N_18131);
or U21934 (N_21934,N_16425,N_16294);
nand U21935 (N_21935,N_18415,N_19093);
xnor U21936 (N_21936,N_18173,N_18589);
xnor U21937 (N_21937,N_16076,N_15271);
xnor U21938 (N_21938,N_17523,N_15466);
and U21939 (N_21939,N_18587,N_15311);
xor U21940 (N_21940,N_19969,N_17682);
xor U21941 (N_21941,N_15996,N_15835);
and U21942 (N_21942,N_19685,N_17656);
nor U21943 (N_21943,N_18649,N_15170);
and U21944 (N_21944,N_16146,N_18728);
nor U21945 (N_21945,N_19042,N_15968);
xnor U21946 (N_21946,N_15623,N_18193);
and U21947 (N_21947,N_16670,N_17679);
xnor U21948 (N_21948,N_16668,N_19481);
and U21949 (N_21949,N_19525,N_17013);
or U21950 (N_21950,N_16128,N_16354);
or U21951 (N_21951,N_17529,N_15793);
xor U21952 (N_21952,N_18934,N_19506);
nand U21953 (N_21953,N_19800,N_16217);
or U21954 (N_21954,N_17480,N_17089);
nand U21955 (N_21955,N_15377,N_15951);
or U21956 (N_21956,N_17034,N_16173);
xor U21957 (N_21957,N_15405,N_15860);
xor U21958 (N_21958,N_18020,N_19171);
or U21959 (N_21959,N_15267,N_16725);
nor U21960 (N_21960,N_15604,N_19884);
nor U21961 (N_21961,N_18684,N_18200);
nor U21962 (N_21962,N_15155,N_18497);
xnor U21963 (N_21963,N_16691,N_18995);
nand U21964 (N_21964,N_16343,N_15389);
xnor U21965 (N_21965,N_18175,N_18745);
nor U21966 (N_21966,N_18685,N_17715);
nand U21967 (N_21967,N_15712,N_18788);
or U21968 (N_21968,N_17173,N_18915);
and U21969 (N_21969,N_19263,N_19399);
and U21970 (N_21970,N_17037,N_19799);
xnor U21971 (N_21971,N_16392,N_19731);
xnor U21972 (N_21972,N_15897,N_17305);
nand U21973 (N_21973,N_19920,N_19319);
and U21974 (N_21974,N_17343,N_19968);
nor U21975 (N_21975,N_18908,N_18179);
and U21976 (N_21976,N_16698,N_16661);
and U21977 (N_21977,N_16614,N_18819);
or U21978 (N_21978,N_17463,N_19142);
and U21979 (N_21979,N_16284,N_16646);
nand U21980 (N_21980,N_18070,N_19837);
nor U21981 (N_21981,N_19271,N_17219);
xor U21982 (N_21982,N_17350,N_17003);
nand U21983 (N_21983,N_15921,N_16609);
nand U21984 (N_21984,N_15411,N_17464);
nand U21985 (N_21985,N_16161,N_17810);
nor U21986 (N_21986,N_18289,N_17012);
and U21987 (N_21987,N_15137,N_17695);
xnor U21988 (N_21988,N_15621,N_15386);
nand U21989 (N_21989,N_19832,N_18428);
nor U21990 (N_21990,N_17441,N_19875);
nor U21991 (N_21991,N_18359,N_17475);
and U21992 (N_21992,N_17218,N_15412);
and U21993 (N_21993,N_19332,N_18282);
and U21994 (N_21994,N_15560,N_15563);
xnor U21995 (N_21995,N_15257,N_19680);
xnor U21996 (N_21996,N_19367,N_17986);
and U21997 (N_21997,N_17885,N_18604);
or U21998 (N_21998,N_16318,N_17876);
and U21999 (N_21999,N_15969,N_15733);
nor U22000 (N_22000,N_16603,N_19634);
nand U22001 (N_22001,N_17797,N_15297);
nor U22002 (N_22002,N_19371,N_16914);
nor U22003 (N_22003,N_18264,N_16802);
xor U22004 (N_22004,N_19886,N_15678);
xor U22005 (N_22005,N_15263,N_17029);
xnor U22006 (N_22006,N_18132,N_15428);
and U22007 (N_22007,N_16712,N_16051);
and U22008 (N_22008,N_19459,N_16095);
xnor U22009 (N_22009,N_15663,N_17161);
or U22010 (N_22010,N_18491,N_19374);
xor U22011 (N_22011,N_15211,N_17151);
or U22012 (N_22012,N_15901,N_17002);
or U22013 (N_22013,N_19816,N_19745);
xnor U22014 (N_22014,N_17262,N_18842);
xor U22015 (N_22015,N_15698,N_17479);
nand U22016 (N_22016,N_16287,N_16162);
and U22017 (N_22017,N_16860,N_19684);
xnor U22018 (N_22018,N_19329,N_18403);
nand U22019 (N_22019,N_15207,N_16982);
nor U22020 (N_22020,N_18702,N_19857);
xnor U22021 (N_22021,N_15674,N_16242);
or U22022 (N_22022,N_17660,N_16170);
nand U22023 (N_22023,N_15689,N_16471);
or U22024 (N_22024,N_19330,N_19197);
or U22025 (N_22025,N_18626,N_17392);
nor U22026 (N_22026,N_18576,N_18584);
nor U22027 (N_22027,N_15555,N_15602);
or U22028 (N_22028,N_16950,N_15918);
or U22029 (N_22029,N_18555,N_19616);
or U22030 (N_22030,N_19119,N_16653);
and U22031 (N_22031,N_15521,N_15208);
or U22032 (N_22032,N_17853,N_19855);
and U22033 (N_22033,N_15153,N_16761);
xor U22034 (N_22034,N_16013,N_19207);
or U22035 (N_22035,N_19301,N_16303);
and U22036 (N_22036,N_16020,N_18652);
nor U22037 (N_22037,N_18609,N_15706);
or U22038 (N_22038,N_16210,N_19801);
or U22039 (N_22039,N_19708,N_15946);
or U22040 (N_22040,N_15079,N_15061);
nor U22041 (N_22041,N_19028,N_15608);
nand U22042 (N_22042,N_19230,N_16112);
and U22043 (N_22043,N_16992,N_16542);
nand U22044 (N_22044,N_15745,N_18092);
nor U22045 (N_22045,N_16365,N_17301);
and U22046 (N_22046,N_17120,N_17684);
or U22047 (N_22047,N_17369,N_19098);
or U22048 (N_22048,N_19354,N_18971);
nand U22049 (N_22049,N_19939,N_17011);
nand U22050 (N_22050,N_18525,N_19984);
and U22051 (N_22051,N_17815,N_16912);
or U22052 (N_22052,N_15697,N_17277);
xor U22053 (N_22053,N_19608,N_19172);
nor U22054 (N_22054,N_16873,N_16137);
xnor U22055 (N_22055,N_15265,N_15518);
and U22056 (N_22056,N_19618,N_18351);
and U22057 (N_22057,N_16931,N_19839);
and U22058 (N_22058,N_16806,N_19805);
nand U22059 (N_22059,N_18198,N_17892);
or U22060 (N_22060,N_18867,N_17931);
and U22061 (N_22061,N_16743,N_16181);
nand U22062 (N_22062,N_17251,N_16677);
or U22063 (N_22063,N_15789,N_16328);
nand U22064 (N_22064,N_19941,N_17992);
xnor U22065 (N_22065,N_15154,N_16594);
nor U22066 (N_22066,N_17550,N_18240);
nor U22067 (N_22067,N_15316,N_15494);
xor U22068 (N_22068,N_16882,N_15795);
nor U22069 (N_22069,N_18650,N_19208);
and U22070 (N_22070,N_16943,N_19151);
nand U22071 (N_22071,N_17080,N_16588);
or U22072 (N_22072,N_16267,N_17900);
or U22073 (N_22073,N_17619,N_15348);
and U22074 (N_22074,N_15335,N_19424);
nand U22075 (N_22075,N_15715,N_17676);
or U22076 (N_22076,N_18473,N_19383);
or U22077 (N_22077,N_18764,N_15122);
nor U22078 (N_22078,N_16589,N_15992);
or U22079 (N_22079,N_16368,N_17147);
nor U22080 (N_22080,N_19933,N_17939);
and U22081 (N_22081,N_17807,N_16827);
nor U22082 (N_22082,N_19924,N_16617);
nor U22083 (N_22083,N_17919,N_17670);
nand U22084 (N_22084,N_18992,N_15453);
and U22085 (N_22085,N_19419,N_17335);
xnor U22086 (N_22086,N_18426,N_17296);
or U22087 (N_22087,N_16595,N_15397);
xnor U22088 (N_22088,N_19867,N_15047);
nand U22089 (N_22089,N_17114,N_19176);
nand U22090 (N_22090,N_15294,N_15815);
nand U22091 (N_22091,N_16814,N_17562);
nand U22092 (N_22092,N_18402,N_18667);
xor U22093 (N_22093,N_16177,N_15027);
and U22094 (N_22094,N_19293,N_17545);
or U22095 (N_22095,N_18228,N_17027);
nand U22096 (N_22096,N_18541,N_18696);
and U22097 (N_22097,N_17742,N_17703);
nor U22098 (N_22098,N_15034,N_18899);
and U22099 (N_22099,N_15568,N_15178);
nor U22100 (N_22100,N_18635,N_19899);
nand U22101 (N_22101,N_18612,N_16756);
and U22102 (N_22102,N_16236,N_18602);
and U22103 (N_22103,N_15138,N_19764);
and U22104 (N_22104,N_16077,N_18554);
nor U22105 (N_22105,N_17287,N_19405);
nor U22106 (N_22106,N_18896,N_17811);
nand U22107 (N_22107,N_18749,N_19997);
nand U22108 (N_22108,N_16434,N_15003);
nor U22109 (N_22109,N_17635,N_18108);
and U22110 (N_22110,N_15643,N_18048);
xor U22111 (N_22111,N_19137,N_18134);
nor U22112 (N_22112,N_17072,N_17686);
xor U22113 (N_22113,N_16926,N_15070);
or U22114 (N_22114,N_15937,N_16016);
nor U22115 (N_22115,N_19210,N_18771);
nand U22116 (N_22116,N_18573,N_16902);
nand U22117 (N_22117,N_16326,N_19349);
xnor U22118 (N_22118,N_15783,N_17744);
nor U22119 (N_22119,N_16152,N_17425);
xnor U22120 (N_22120,N_15008,N_15492);
nor U22121 (N_22121,N_16357,N_19720);
nand U22122 (N_22122,N_17819,N_16046);
and U22123 (N_22123,N_17825,N_17519);
or U22124 (N_22124,N_18709,N_16039);
nand U22125 (N_22125,N_18236,N_19650);
or U22126 (N_22126,N_19873,N_16423);
xnor U22127 (N_22127,N_17767,N_16118);
or U22128 (N_22128,N_18261,N_16304);
and U22129 (N_22129,N_16250,N_15091);
xor U22130 (N_22130,N_17506,N_16775);
nand U22131 (N_22131,N_15482,N_18656);
xor U22132 (N_22132,N_19710,N_18616);
nor U22133 (N_22133,N_15043,N_18567);
xor U22134 (N_22134,N_19819,N_19063);
nor U22135 (N_22135,N_15407,N_19694);
nand U22136 (N_22136,N_19665,N_17406);
xor U22137 (N_22137,N_16006,N_17248);
nand U22138 (N_22138,N_19914,N_15717);
nor U22139 (N_22139,N_19494,N_18969);
nand U22140 (N_22140,N_18027,N_18361);
or U22141 (N_22141,N_16466,N_19512);
nand U22142 (N_22142,N_15023,N_17116);
nand U22143 (N_22143,N_17508,N_15737);
and U22144 (N_22144,N_16930,N_19897);
nor U22145 (N_22145,N_15108,N_18613);
xnor U22146 (N_22146,N_16130,N_18045);
xnor U22147 (N_22147,N_15702,N_18978);
and U22148 (N_22148,N_18689,N_16735);
xnor U22149 (N_22149,N_17410,N_16271);
or U22150 (N_22150,N_16605,N_16844);
nand U22151 (N_22151,N_18356,N_15437);
and U22152 (N_22152,N_15128,N_18317);
or U22153 (N_22153,N_16147,N_19318);
xnor U22154 (N_22154,N_17808,N_17567);
or U22155 (N_22155,N_19121,N_15505);
nand U22156 (N_22156,N_16607,N_18392);
nor U22157 (N_22157,N_18389,N_16282);
or U22158 (N_22158,N_19430,N_17669);
xnor U22159 (N_22159,N_18367,N_19548);
and U22160 (N_22160,N_16631,N_18281);
nor U22161 (N_22161,N_19336,N_15292);
or U22162 (N_22162,N_15227,N_19827);
or U22163 (N_22163,N_15103,N_19218);
nand U22164 (N_22164,N_16566,N_15324);
and U22165 (N_22165,N_19625,N_17397);
nand U22166 (N_22166,N_15885,N_15930);
nand U22167 (N_22167,N_15907,N_17178);
and U22168 (N_22168,N_16010,N_15481);
xnor U22169 (N_22169,N_19228,N_18614);
and U22170 (N_22170,N_18458,N_15209);
or U22171 (N_22171,N_15542,N_19535);
and U22172 (N_22172,N_19377,N_17641);
xnor U22173 (N_22173,N_17405,N_15234);
or U22174 (N_22174,N_18818,N_17474);
or U22175 (N_22175,N_16895,N_18875);
and U22176 (N_22176,N_15831,N_16135);
and U22177 (N_22177,N_15406,N_15851);
and U22178 (N_22178,N_18221,N_17507);
or U22179 (N_22179,N_17626,N_18948);
or U22180 (N_22180,N_16126,N_18770);
nand U22181 (N_22181,N_15614,N_16488);
and U22182 (N_22182,N_16938,N_17186);
nor U22183 (N_22183,N_17044,N_18304);
and U22184 (N_22184,N_17578,N_17959);
xor U22185 (N_22185,N_17734,N_15014);
or U22186 (N_22186,N_19276,N_16868);
nor U22187 (N_22187,N_19912,N_18448);
and U22188 (N_22188,N_16767,N_16187);
nand U22189 (N_22189,N_16826,N_18444);
nor U22190 (N_22190,N_18110,N_18767);
or U22191 (N_22191,N_18700,N_15569);
nor U22192 (N_22192,N_18641,N_17950);
xnor U22193 (N_22193,N_19995,N_18844);
nand U22194 (N_22194,N_18938,N_15384);
and U22195 (N_22195,N_17865,N_18748);
and U22196 (N_22196,N_18521,N_17288);
or U22197 (N_22197,N_16022,N_15748);
nor U22198 (N_22198,N_15943,N_17488);
nand U22199 (N_22199,N_19303,N_16678);
or U22200 (N_22200,N_15889,N_18952);
xnor U22201 (N_22201,N_18722,N_18797);
or U22202 (N_22202,N_16477,N_15824);
or U22203 (N_22203,N_19060,N_17718);
and U22204 (N_22204,N_18400,N_15301);
xor U22205 (N_22205,N_15809,N_15106);
nand U22206 (N_22206,N_18166,N_18224);
nand U22207 (N_22207,N_17904,N_16107);
xor U22208 (N_22208,N_19872,N_16316);
and U22209 (N_22209,N_19760,N_17789);
xnor U22210 (N_22210,N_18121,N_17849);
xor U22211 (N_22211,N_15069,N_15956);
nor U22212 (N_22212,N_16598,N_15973);
nand U22213 (N_22213,N_15782,N_16069);
nand U22214 (N_22214,N_18039,N_16901);
nor U22215 (N_22215,N_19951,N_16233);
nand U22216 (N_22216,N_15319,N_15517);
nor U22217 (N_22217,N_15818,N_16988);
nand U22218 (N_22218,N_17126,N_15777);
or U22219 (N_22219,N_17194,N_16942);
and U22220 (N_22220,N_16971,N_19552);
nor U22221 (N_22221,N_16647,N_15575);
xnor U22222 (N_22222,N_15680,N_17777);
xnor U22223 (N_22223,N_15959,N_18210);
or U22224 (N_22224,N_18137,N_17175);
or U22225 (N_22225,N_16389,N_19189);
nor U22226 (N_22226,N_18436,N_18738);
or U22227 (N_22227,N_15347,N_18331);
or U22228 (N_22228,N_16997,N_19721);
nand U22229 (N_22229,N_18787,N_19280);
nand U22230 (N_22230,N_15076,N_19311);
and U22231 (N_22231,N_19928,N_16506);
nor U22232 (N_22232,N_18647,N_16320);
nand U22233 (N_22233,N_19076,N_17726);
nand U22234 (N_22234,N_16599,N_16094);
nand U22235 (N_22235,N_15933,N_17285);
or U22236 (N_22236,N_19130,N_18634);
nor U22237 (N_22237,N_19080,N_15038);
nor U22238 (N_22238,N_17210,N_17502);
xnor U22239 (N_22239,N_18932,N_18556);
or U22240 (N_22240,N_19957,N_16405);
and U22241 (N_22241,N_16779,N_19267);
xor U22242 (N_22242,N_16493,N_17437);
or U22243 (N_22243,N_19019,N_15383);
nor U22244 (N_22244,N_18761,N_18956);
xor U22245 (N_22245,N_17514,N_19131);
or U22246 (N_22246,N_19724,N_17440);
or U22247 (N_22247,N_15086,N_19088);
xor U22248 (N_22248,N_16925,N_18425);
and U22249 (N_22249,N_18363,N_18692);
and U22250 (N_22250,N_15400,N_19610);
or U22251 (N_22251,N_16918,N_17838);
or U22252 (N_22252,N_17628,N_18486);
xnor U22253 (N_22253,N_16625,N_17964);
xnor U22254 (N_22254,N_15676,N_18005);
or U22255 (N_22255,N_16492,N_16658);
nand U22256 (N_22256,N_15955,N_17857);
nor U22257 (N_22257,N_15844,N_16183);
nand U22258 (N_22258,N_18847,N_18316);
and U22259 (N_22259,N_18232,N_16685);
and U22260 (N_22260,N_18247,N_18680);
nand U22261 (N_22261,N_18201,N_17864);
and U22262 (N_22262,N_16538,N_17077);
or U22263 (N_22263,N_17884,N_16214);
and U22264 (N_22264,N_19186,N_15256);
and U22265 (N_22265,N_17316,N_19296);
nand U22266 (N_22266,N_18275,N_17598);
nand U22267 (N_22267,N_19477,N_17443);
and U22268 (N_22268,N_18300,N_17401);
xnor U22269 (N_22269,N_18957,N_16910);
and U22270 (N_22270,N_17318,N_17932);
xor U22271 (N_22271,N_19976,N_18775);
nand U22272 (N_22272,N_16722,N_18355);
and U22273 (N_22273,N_18713,N_18675);
or U22274 (N_22274,N_17059,N_18757);
nand U22275 (N_22275,N_18753,N_15382);
nand U22276 (N_22276,N_18802,N_17490);
nand U22277 (N_22277,N_17326,N_17057);
or U22278 (N_22278,N_16012,N_17926);
nand U22279 (N_22279,N_19100,N_18662);
nor U22280 (N_22280,N_18593,N_16805);
and U22281 (N_22281,N_16252,N_18740);
and U22282 (N_22282,N_17062,N_17205);
nor U22283 (N_22283,N_15827,N_19048);
or U22284 (N_22284,N_15530,N_19022);
nor U22285 (N_22285,N_18526,N_15141);
xnor U22286 (N_22286,N_16038,N_19598);
and U22287 (N_22287,N_17584,N_18288);
nand U22288 (N_22288,N_19040,N_17324);
nand U22289 (N_22289,N_18138,N_15929);
xnor U22290 (N_22290,N_19190,N_16068);
and U22291 (N_22291,N_15033,N_18461);
xor U22292 (N_22292,N_18642,N_19851);
nand U22293 (N_22293,N_19307,N_18961);
nand U22294 (N_22294,N_17872,N_18919);
nand U22295 (N_22295,N_16503,N_17375);
nand U22296 (N_22296,N_18864,N_15219);
nor U22297 (N_22297,N_19324,N_19149);
and U22298 (N_22298,N_15438,N_17540);
and U22299 (N_22299,N_19000,N_19032);
xnor U22300 (N_22300,N_15983,N_19609);
and U22301 (N_22301,N_17798,N_19937);
nand U22302 (N_22302,N_15588,N_18799);
or U22303 (N_22303,N_16465,N_15896);
nor U22304 (N_22304,N_16136,N_19150);
nand U22305 (N_22305,N_16927,N_18290);
or U22306 (N_22306,N_18920,N_15315);
xnor U22307 (N_22307,N_19244,N_16716);
xor U22308 (N_22308,N_19932,N_15104);
xor U22309 (N_22309,N_15532,N_19555);
xnor U22310 (N_22310,N_16448,N_18376);
nand U22311 (N_22311,N_16849,N_15484);
and U22312 (N_22312,N_15830,N_19408);
and U22313 (N_22313,N_18972,N_16275);
or U22314 (N_22314,N_16371,N_15331);
and U22315 (N_22315,N_15821,N_18419);
nand U22316 (N_22316,N_18705,N_17727);
or U22317 (N_22317,N_19221,N_15422);
or U22318 (N_22318,N_18828,N_15525);
xor U22319 (N_22319,N_17936,N_16907);
or U22320 (N_22320,N_19547,N_16600);
and U22321 (N_22321,N_15403,N_15975);
nand U22322 (N_22322,N_16315,N_16331);
nand U22323 (N_22323,N_19748,N_17689);
xnor U22324 (N_22324,N_15741,N_18774);
and U22325 (N_22325,N_15273,N_17018);
nor U22326 (N_22326,N_15258,N_16804);
xnor U22327 (N_22327,N_19570,N_17665);
nand U22328 (N_22328,N_16254,N_18035);
nor U22329 (N_22329,N_18333,N_18469);
or U22330 (N_22330,N_17416,N_18549);
nor U22331 (N_22331,N_19504,N_16305);
or U22332 (N_22332,N_17801,N_16689);
or U22333 (N_22333,N_16457,N_15111);
xnor U22334 (N_22334,N_18412,N_18143);
nor U22335 (N_22335,N_15618,N_18334);
nand U22336 (N_22336,N_17106,N_16299);
nand U22337 (N_22337,N_17868,N_16149);
and U22338 (N_22338,N_15902,N_16652);
or U22339 (N_22339,N_18302,N_18985);
xor U22340 (N_22340,N_18754,N_19661);
nor U22341 (N_22341,N_17539,N_17907);
or U22342 (N_22342,N_19545,N_19370);
or U22343 (N_22343,N_17764,N_15313);
or U22344 (N_22344,N_17510,N_18606);
nor U22345 (N_22345,N_18427,N_16924);
or U22346 (N_22346,N_18323,N_17918);
xnor U22347 (N_22347,N_17792,N_16702);
xnor U22348 (N_22348,N_18829,N_19393);
or U22349 (N_22349,N_15391,N_16393);
xnor U22350 (N_22350,N_18510,N_18528);
nor U22351 (N_22351,N_18706,N_18655);
or U22352 (N_22352,N_15862,N_15395);
or U22353 (N_22353,N_17886,N_19830);
nor U22354 (N_22354,N_15764,N_18812);
and U22355 (N_22355,N_18846,N_15487);
nand U22356 (N_22356,N_17671,N_19954);
xor U22357 (N_22357,N_19406,N_19593);
or U22358 (N_22358,N_18485,N_19986);
nor U22359 (N_22359,N_15625,N_17809);
nand U22360 (N_22360,N_16891,N_15109);
xnor U22361 (N_22361,N_18357,N_16626);
or U22362 (N_22362,N_17558,N_17957);
xor U22363 (N_22363,N_19982,N_17261);
or U22364 (N_22364,N_19173,N_17103);
xor U22365 (N_22365,N_15390,N_15445);
nand U22366 (N_22366,N_16863,N_17115);
and U22367 (N_22367,N_16158,N_16472);
and U22368 (N_22368,N_19304,N_17328);
xnor U22369 (N_22369,N_16043,N_17244);
xnor U22370 (N_22370,N_15808,N_16717);
or U22371 (N_22371,N_18177,N_19389);
xor U22372 (N_22372,N_16138,N_16564);
and U22373 (N_22373,N_16965,N_16319);
nor U22374 (N_22374,N_17769,N_17306);
or U22375 (N_22375,N_16344,N_19789);
nand U22376 (N_22376,N_19352,N_19469);
nor U22377 (N_22377,N_15610,N_15351);
xnor U22378 (N_22378,N_17221,N_17283);
xnor U22379 (N_22379,N_16336,N_17973);
nand U22380 (N_22380,N_18891,N_16066);
xor U22381 (N_22381,N_19031,N_17549);
or U22382 (N_22382,N_18434,N_18822);
and U22383 (N_22383,N_17164,N_19757);
nand U22384 (N_22384,N_17200,N_18096);
nand U22385 (N_22385,N_18979,N_16959);
nor U22386 (N_22386,N_18438,N_16782);
nor U22387 (N_22387,N_17197,N_18406);
and U22388 (N_22388,N_18348,N_18140);
and U22389 (N_22389,N_19429,N_15549);
nand U22390 (N_22390,N_15193,N_19122);
nor U22391 (N_22391,N_15089,N_16300);
and U22392 (N_22392,N_17552,N_15707);
or U22393 (N_22393,N_17632,N_19036);
or U22394 (N_22394,N_15175,N_17840);
or U22395 (N_22395,N_16455,N_19841);
or U22396 (N_22396,N_15373,N_19224);
or U22397 (N_22397,N_17273,N_17713);
nor U22398 (N_22398,N_18309,N_19177);
nor U22399 (N_22399,N_18868,N_15928);
xor U22400 (N_22400,N_18270,N_15010);
nor U22401 (N_22401,N_16816,N_17017);
nor U22402 (N_22402,N_15962,N_16684);
xor U22403 (N_22403,N_19143,N_16139);
nand U22404 (N_22404,N_18353,N_16557);
or U22405 (N_22405,N_15580,N_18529);
or U22406 (N_22406,N_17450,N_17223);
and U22407 (N_22407,N_16643,N_18237);
xnor U22408 (N_22408,N_18862,N_17693);
nor U22409 (N_22409,N_19384,N_16777);
and U22410 (N_22410,N_17485,N_15029);
and U22411 (N_22411,N_15704,N_15293);
nand U22412 (N_22412,N_17135,N_18246);
xnor U22413 (N_22413,N_15784,N_17952);
xor U22414 (N_22414,N_17108,N_18782);
nor U22415 (N_22415,N_18231,N_15512);
xnor U22416 (N_22416,N_16908,N_15222);
or U22417 (N_22417,N_15291,N_18998);
nand U22418 (N_22418,N_15873,N_19777);
nand U22419 (N_22419,N_15075,N_17698);
or U22420 (N_22420,N_17563,N_19956);
and U22421 (N_22421,N_17152,N_15150);
or U22422 (N_22422,N_16641,N_16384);
nor U22423 (N_22423,N_18145,N_18273);
or U22424 (N_22424,N_18294,N_18933);
and U22425 (N_22425,N_19574,N_19520);
nand U22426 (N_22426,N_15801,N_15510);
xor U22427 (N_22427,N_17442,N_18931);
or U22428 (N_22428,N_19813,N_16230);
nor U22429 (N_22429,N_17254,N_15050);
xor U22430 (N_22430,N_16990,N_17587);
xnor U22431 (N_22431,N_18038,N_18365);
xor U22432 (N_22432,N_18805,N_18909);
nand U22433 (N_22433,N_19782,N_16306);
nor U22434 (N_22434,N_16937,N_16019);
nand U22435 (N_22435,N_17757,N_15278);
xnor U22436 (N_22436,N_15796,N_15248);
nand U22437 (N_22437,N_16972,N_16341);
nor U22438 (N_22438,N_15867,N_17061);
nor U22439 (N_22439,N_18095,N_16977);
nand U22440 (N_22440,N_17551,N_17741);
xor U22441 (N_22441,N_19489,N_19085);
or U22442 (N_22442,N_16490,N_16000);
nand U22443 (N_22443,N_17381,N_19515);
and U22444 (N_22444,N_17638,N_18543);
nor U22445 (N_22445,N_19641,N_19105);
or U22446 (N_22446,N_19194,N_17420);
and U22447 (N_22447,N_17148,N_15665);
or U22448 (N_22448,N_16029,N_19860);
or U22449 (N_22449,N_15242,N_17105);
or U22450 (N_22450,N_17005,N_17640);
or U22451 (N_22451,N_19402,N_17526);
nand U22452 (N_22452,N_15533,N_19938);
and U22453 (N_22453,N_19514,N_16408);
and U22454 (N_22454,N_16721,N_19061);
and U22455 (N_22455,N_16018,N_17041);
or U22456 (N_22456,N_18311,N_19833);
xor U22457 (N_22457,N_16818,N_18736);
and U22458 (N_22458,N_15417,N_19270);
nor U22459 (N_22459,N_17586,N_16900);
xnor U22460 (N_22460,N_15376,N_15472);
or U22461 (N_22461,N_18639,N_19018);
and U22462 (N_22462,N_16206,N_16338);
nand U22463 (N_22463,N_17915,N_19653);
nor U22464 (N_22464,N_15923,N_16945);
and U22465 (N_22465,N_18759,N_16498);
and U22466 (N_22466,N_17863,N_15881);
nand U22467 (N_22467,N_18568,N_15183);
nand U22468 (N_22468,N_15118,N_17575);
and U22469 (N_22469,N_17564,N_15945);
nor U22470 (N_22470,N_18714,N_17096);
nand U22471 (N_22471,N_17158,N_16244);
xor U22472 (N_22472,N_15461,N_15641);
and U22473 (N_22473,N_15093,N_18372);
or U22474 (N_22474,N_15459,N_16003);
nor U22475 (N_22475,N_17354,N_16485);
nand U22476 (N_22476,N_18374,N_19689);
xnor U22477 (N_22477,N_17766,N_18729);
and U22478 (N_22478,N_16430,N_18423);
or U22479 (N_22479,N_19783,N_15582);
nor U22480 (N_22480,N_19453,N_15125);
nor U22481 (N_22481,N_16172,N_17541);
nor U22482 (N_22482,N_15379,N_16378);
or U22483 (N_22483,N_16097,N_18343);
nor U22484 (N_22484,N_18980,N_16124);
nor U22485 (N_22485,N_18030,N_19107);
xnor U22486 (N_22486,N_19078,N_16613);
or U22487 (N_22487,N_15374,N_17234);
and U22488 (N_22488,N_17030,N_17827);
xnor U22489 (N_22489,N_17068,N_15838);
nand U22490 (N_22490,N_18763,N_19144);
and U22491 (N_22491,N_15544,N_19474);
xnor U22492 (N_22492,N_15476,N_19243);
or U22493 (N_22493,N_17934,N_18183);
or U22494 (N_22494,N_16801,N_15113);
and U22495 (N_22495,N_15105,N_18445);
and U22496 (N_22496,N_17582,N_15757);
xnor U22497 (N_22497,N_16297,N_15545);
nand U22498 (N_22498,N_19328,N_15281);
or U22499 (N_22499,N_17515,N_18741);
or U22500 (N_22500,N_17947,N_17559);
nor U22501 (N_22501,N_15166,N_17398);
nand U22502 (N_22502,N_15925,N_16519);
and U22503 (N_22503,N_15459,N_18977);
xnor U22504 (N_22504,N_17676,N_19648);
xnor U22505 (N_22505,N_18649,N_17184);
xnor U22506 (N_22506,N_16220,N_19057);
and U22507 (N_22507,N_19829,N_15825);
nand U22508 (N_22508,N_19197,N_17468);
and U22509 (N_22509,N_19260,N_17858);
and U22510 (N_22510,N_17469,N_15730);
xnor U22511 (N_22511,N_15811,N_19726);
nand U22512 (N_22512,N_19947,N_19724);
or U22513 (N_22513,N_19932,N_16162);
and U22514 (N_22514,N_17647,N_15561);
nand U22515 (N_22515,N_16599,N_16629);
and U22516 (N_22516,N_17781,N_18256);
and U22517 (N_22517,N_17307,N_18217);
and U22518 (N_22518,N_19501,N_16914);
xor U22519 (N_22519,N_15509,N_16566);
nor U22520 (N_22520,N_17377,N_15043);
and U22521 (N_22521,N_19496,N_17407);
nor U22522 (N_22522,N_19306,N_15763);
or U22523 (N_22523,N_16759,N_18006);
xor U22524 (N_22524,N_18287,N_19174);
or U22525 (N_22525,N_18188,N_17145);
xor U22526 (N_22526,N_19717,N_15809);
nand U22527 (N_22527,N_16888,N_18078);
nand U22528 (N_22528,N_18013,N_19407);
and U22529 (N_22529,N_15016,N_18447);
xor U22530 (N_22530,N_18343,N_19261);
and U22531 (N_22531,N_15626,N_18957);
nor U22532 (N_22532,N_16543,N_16316);
and U22533 (N_22533,N_15225,N_18912);
and U22534 (N_22534,N_18334,N_19150);
nor U22535 (N_22535,N_18629,N_17798);
nor U22536 (N_22536,N_17574,N_19337);
and U22537 (N_22537,N_16767,N_18882);
and U22538 (N_22538,N_18648,N_18432);
and U22539 (N_22539,N_15105,N_16299);
or U22540 (N_22540,N_18865,N_19143);
nand U22541 (N_22541,N_17959,N_19289);
xnor U22542 (N_22542,N_16816,N_18628);
xnor U22543 (N_22543,N_19379,N_16911);
nor U22544 (N_22544,N_16009,N_17331);
nand U22545 (N_22545,N_19753,N_18882);
nand U22546 (N_22546,N_19412,N_15917);
nand U22547 (N_22547,N_17490,N_19935);
xnor U22548 (N_22548,N_17667,N_19000);
or U22549 (N_22549,N_19222,N_16451);
nor U22550 (N_22550,N_19647,N_18612);
or U22551 (N_22551,N_17779,N_16637);
xnor U22552 (N_22552,N_17543,N_17096);
and U22553 (N_22553,N_16030,N_18849);
or U22554 (N_22554,N_16352,N_19425);
xnor U22555 (N_22555,N_17167,N_15408);
or U22556 (N_22556,N_16019,N_17380);
nor U22557 (N_22557,N_17347,N_15659);
xnor U22558 (N_22558,N_18490,N_18690);
and U22559 (N_22559,N_16292,N_19085);
xnor U22560 (N_22560,N_17946,N_15541);
or U22561 (N_22561,N_17357,N_19739);
and U22562 (N_22562,N_16126,N_18460);
or U22563 (N_22563,N_15437,N_18148);
or U22564 (N_22564,N_17584,N_17774);
nor U22565 (N_22565,N_17662,N_15318);
nor U22566 (N_22566,N_18000,N_17949);
nand U22567 (N_22567,N_16523,N_16029);
xor U22568 (N_22568,N_19490,N_17320);
and U22569 (N_22569,N_16811,N_18212);
and U22570 (N_22570,N_15373,N_19237);
and U22571 (N_22571,N_15689,N_19331);
nand U22572 (N_22572,N_16284,N_16069);
or U22573 (N_22573,N_17224,N_16898);
xnor U22574 (N_22574,N_19072,N_17570);
xor U22575 (N_22575,N_18455,N_19782);
and U22576 (N_22576,N_16399,N_19561);
or U22577 (N_22577,N_19820,N_17154);
and U22578 (N_22578,N_15288,N_19823);
and U22579 (N_22579,N_17493,N_17344);
xor U22580 (N_22580,N_15994,N_16940);
or U22581 (N_22581,N_17738,N_19693);
and U22582 (N_22582,N_18543,N_18401);
nor U22583 (N_22583,N_17428,N_16807);
nand U22584 (N_22584,N_16777,N_15112);
xnor U22585 (N_22585,N_19151,N_15720);
and U22586 (N_22586,N_18723,N_18849);
and U22587 (N_22587,N_15901,N_19969);
and U22588 (N_22588,N_16436,N_17874);
and U22589 (N_22589,N_16588,N_16825);
xor U22590 (N_22590,N_19709,N_17634);
xor U22591 (N_22591,N_15440,N_17442);
or U22592 (N_22592,N_17482,N_15958);
or U22593 (N_22593,N_16097,N_17255);
xnor U22594 (N_22594,N_16601,N_16054);
and U22595 (N_22595,N_17369,N_19917);
nor U22596 (N_22596,N_18895,N_16539);
nand U22597 (N_22597,N_17368,N_16633);
nor U22598 (N_22598,N_15303,N_15534);
or U22599 (N_22599,N_15694,N_17573);
nor U22600 (N_22600,N_19655,N_18192);
nand U22601 (N_22601,N_18375,N_19340);
and U22602 (N_22602,N_16913,N_18173);
nor U22603 (N_22603,N_16495,N_18435);
xor U22604 (N_22604,N_19565,N_19684);
or U22605 (N_22605,N_19356,N_18620);
and U22606 (N_22606,N_17073,N_19176);
xnor U22607 (N_22607,N_15610,N_17673);
xnor U22608 (N_22608,N_18313,N_15479);
or U22609 (N_22609,N_16789,N_19856);
or U22610 (N_22610,N_15666,N_17462);
nand U22611 (N_22611,N_16362,N_18669);
nand U22612 (N_22612,N_17150,N_19856);
and U22613 (N_22613,N_17835,N_18923);
or U22614 (N_22614,N_16436,N_19049);
or U22615 (N_22615,N_19841,N_17324);
nand U22616 (N_22616,N_17271,N_17130);
xor U22617 (N_22617,N_18123,N_16427);
and U22618 (N_22618,N_18895,N_18393);
nor U22619 (N_22619,N_18188,N_16069);
xnor U22620 (N_22620,N_16467,N_15491);
and U22621 (N_22621,N_15441,N_18504);
or U22622 (N_22622,N_15960,N_15940);
and U22623 (N_22623,N_15428,N_19556);
nor U22624 (N_22624,N_17602,N_16527);
nor U22625 (N_22625,N_16718,N_18534);
and U22626 (N_22626,N_15989,N_17829);
nand U22627 (N_22627,N_18762,N_15712);
xor U22628 (N_22628,N_18022,N_15549);
and U22629 (N_22629,N_16194,N_17080);
nand U22630 (N_22630,N_15740,N_19126);
xnor U22631 (N_22631,N_18755,N_18591);
and U22632 (N_22632,N_19160,N_16894);
and U22633 (N_22633,N_18333,N_15962);
xnor U22634 (N_22634,N_17353,N_16210);
nand U22635 (N_22635,N_19772,N_18906);
and U22636 (N_22636,N_18775,N_19433);
and U22637 (N_22637,N_19170,N_19612);
nor U22638 (N_22638,N_18620,N_17533);
xor U22639 (N_22639,N_19799,N_19546);
nand U22640 (N_22640,N_17254,N_18609);
xor U22641 (N_22641,N_17846,N_17139);
nand U22642 (N_22642,N_16818,N_15958);
nor U22643 (N_22643,N_18848,N_17282);
or U22644 (N_22644,N_15209,N_18106);
nand U22645 (N_22645,N_15950,N_17278);
and U22646 (N_22646,N_17320,N_19915);
or U22647 (N_22647,N_19200,N_19931);
nor U22648 (N_22648,N_16102,N_16982);
and U22649 (N_22649,N_15528,N_16383);
or U22650 (N_22650,N_18325,N_17251);
and U22651 (N_22651,N_17193,N_17653);
or U22652 (N_22652,N_19730,N_15790);
xor U22653 (N_22653,N_15692,N_17309);
nand U22654 (N_22654,N_17994,N_19441);
and U22655 (N_22655,N_19348,N_19517);
nor U22656 (N_22656,N_16585,N_18308);
xor U22657 (N_22657,N_16116,N_15670);
and U22658 (N_22658,N_17661,N_17841);
or U22659 (N_22659,N_15375,N_18651);
or U22660 (N_22660,N_15725,N_19978);
or U22661 (N_22661,N_19031,N_17071);
xnor U22662 (N_22662,N_19992,N_15938);
xnor U22663 (N_22663,N_19041,N_16599);
nand U22664 (N_22664,N_18523,N_18139);
and U22665 (N_22665,N_17701,N_19541);
and U22666 (N_22666,N_17479,N_17119);
and U22667 (N_22667,N_19736,N_15409);
xor U22668 (N_22668,N_18338,N_16565);
and U22669 (N_22669,N_19622,N_18731);
nand U22670 (N_22670,N_15280,N_17248);
or U22671 (N_22671,N_18149,N_19086);
nand U22672 (N_22672,N_15403,N_19055);
and U22673 (N_22673,N_16906,N_18788);
nor U22674 (N_22674,N_15342,N_19715);
xor U22675 (N_22675,N_18032,N_15119);
or U22676 (N_22676,N_15950,N_19190);
nor U22677 (N_22677,N_18598,N_19201);
nor U22678 (N_22678,N_18083,N_15131);
nor U22679 (N_22679,N_19755,N_17108);
nand U22680 (N_22680,N_18836,N_18350);
nor U22681 (N_22681,N_16121,N_16844);
or U22682 (N_22682,N_17444,N_19251);
nand U22683 (N_22683,N_15229,N_16976);
nand U22684 (N_22684,N_17929,N_16560);
and U22685 (N_22685,N_17273,N_16744);
xor U22686 (N_22686,N_18030,N_18059);
nor U22687 (N_22687,N_15394,N_17628);
xnor U22688 (N_22688,N_17939,N_17917);
nor U22689 (N_22689,N_19243,N_18187);
xnor U22690 (N_22690,N_16177,N_19274);
or U22691 (N_22691,N_19834,N_15384);
and U22692 (N_22692,N_18238,N_16211);
or U22693 (N_22693,N_15944,N_16898);
nor U22694 (N_22694,N_18825,N_16909);
or U22695 (N_22695,N_16714,N_15372);
nor U22696 (N_22696,N_19698,N_15966);
xor U22697 (N_22697,N_19720,N_18654);
and U22698 (N_22698,N_16492,N_19475);
nand U22699 (N_22699,N_15342,N_18386);
and U22700 (N_22700,N_16210,N_15519);
nor U22701 (N_22701,N_15534,N_17592);
nand U22702 (N_22702,N_17300,N_18441);
nand U22703 (N_22703,N_15504,N_19712);
or U22704 (N_22704,N_18536,N_15656);
or U22705 (N_22705,N_18226,N_19770);
xnor U22706 (N_22706,N_18197,N_18005);
nand U22707 (N_22707,N_19133,N_19751);
nor U22708 (N_22708,N_15059,N_19842);
nand U22709 (N_22709,N_15484,N_18533);
and U22710 (N_22710,N_15788,N_15208);
or U22711 (N_22711,N_18254,N_16810);
xnor U22712 (N_22712,N_17089,N_16181);
and U22713 (N_22713,N_15733,N_15010);
nor U22714 (N_22714,N_15861,N_18232);
nor U22715 (N_22715,N_17159,N_15391);
xor U22716 (N_22716,N_19826,N_16075);
and U22717 (N_22717,N_15012,N_19627);
nor U22718 (N_22718,N_19272,N_18116);
and U22719 (N_22719,N_16921,N_17221);
or U22720 (N_22720,N_19178,N_17884);
nand U22721 (N_22721,N_19260,N_18787);
or U22722 (N_22722,N_19301,N_17268);
nand U22723 (N_22723,N_15594,N_16865);
nor U22724 (N_22724,N_15958,N_17742);
xnor U22725 (N_22725,N_16576,N_17989);
xor U22726 (N_22726,N_17586,N_19798);
xnor U22727 (N_22727,N_18715,N_16429);
nand U22728 (N_22728,N_19738,N_16055);
nor U22729 (N_22729,N_19003,N_15300);
or U22730 (N_22730,N_17317,N_15287);
xor U22731 (N_22731,N_19126,N_18339);
xor U22732 (N_22732,N_18840,N_16653);
and U22733 (N_22733,N_16355,N_16810);
nor U22734 (N_22734,N_16545,N_18991);
or U22735 (N_22735,N_18456,N_19073);
nand U22736 (N_22736,N_15793,N_19739);
or U22737 (N_22737,N_17219,N_19390);
nor U22738 (N_22738,N_17935,N_16239);
nand U22739 (N_22739,N_15798,N_16238);
xor U22740 (N_22740,N_18020,N_18748);
nand U22741 (N_22741,N_16178,N_17287);
and U22742 (N_22742,N_19486,N_18020);
nor U22743 (N_22743,N_19584,N_18659);
nor U22744 (N_22744,N_18082,N_19710);
xor U22745 (N_22745,N_19889,N_19710);
nand U22746 (N_22746,N_17022,N_16256);
xor U22747 (N_22747,N_17496,N_18595);
or U22748 (N_22748,N_16834,N_16327);
xnor U22749 (N_22749,N_17910,N_19924);
nand U22750 (N_22750,N_18817,N_15881);
nor U22751 (N_22751,N_17886,N_15782);
nand U22752 (N_22752,N_18764,N_17407);
or U22753 (N_22753,N_15191,N_15307);
or U22754 (N_22754,N_18869,N_16084);
xnor U22755 (N_22755,N_16156,N_18976);
xnor U22756 (N_22756,N_18790,N_18532);
nand U22757 (N_22757,N_17731,N_15019);
nor U22758 (N_22758,N_19138,N_16847);
nor U22759 (N_22759,N_19197,N_17096);
nor U22760 (N_22760,N_15704,N_18706);
xnor U22761 (N_22761,N_16162,N_19472);
nand U22762 (N_22762,N_18536,N_19017);
and U22763 (N_22763,N_18055,N_17059);
and U22764 (N_22764,N_16445,N_18522);
and U22765 (N_22765,N_16507,N_19917);
or U22766 (N_22766,N_15197,N_19693);
or U22767 (N_22767,N_15261,N_17908);
xnor U22768 (N_22768,N_15323,N_15776);
nand U22769 (N_22769,N_19376,N_16795);
xnor U22770 (N_22770,N_17961,N_18648);
and U22771 (N_22771,N_16991,N_15583);
and U22772 (N_22772,N_19040,N_16912);
nor U22773 (N_22773,N_18801,N_19902);
and U22774 (N_22774,N_19207,N_15196);
and U22775 (N_22775,N_19302,N_15428);
nand U22776 (N_22776,N_15309,N_16132);
nand U22777 (N_22777,N_17529,N_17053);
or U22778 (N_22778,N_17990,N_17232);
nor U22779 (N_22779,N_18467,N_19317);
and U22780 (N_22780,N_17023,N_19978);
xor U22781 (N_22781,N_16557,N_17976);
and U22782 (N_22782,N_16379,N_16199);
xnor U22783 (N_22783,N_15078,N_15416);
or U22784 (N_22784,N_18416,N_17484);
and U22785 (N_22785,N_18905,N_19749);
and U22786 (N_22786,N_17597,N_16969);
nand U22787 (N_22787,N_19237,N_15121);
or U22788 (N_22788,N_15793,N_19356);
xor U22789 (N_22789,N_19105,N_16120);
nor U22790 (N_22790,N_19103,N_18140);
or U22791 (N_22791,N_16413,N_17325);
nor U22792 (N_22792,N_18134,N_19582);
xnor U22793 (N_22793,N_15647,N_16731);
and U22794 (N_22794,N_19725,N_17727);
or U22795 (N_22795,N_17053,N_17244);
xor U22796 (N_22796,N_17627,N_18222);
nor U22797 (N_22797,N_16744,N_15562);
xor U22798 (N_22798,N_19185,N_16604);
and U22799 (N_22799,N_18150,N_16813);
nor U22800 (N_22800,N_16276,N_15094);
xnor U22801 (N_22801,N_18986,N_17473);
or U22802 (N_22802,N_16495,N_17740);
nand U22803 (N_22803,N_19864,N_17645);
nor U22804 (N_22804,N_18666,N_17833);
nand U22805 (N_22805,N_16949,N_15727);
nand U22806 (N_22806,N_18418,N_19703);
xor U22807 (N_22807,N_16410,N_15935);
xnor U22808 (N_22808,N_17993,N_17391);
xnor U22809 (N_22809,N_15662,N_15732);
or U22810 (N_22810,N_18195,N_18755);
or U22811 (N_22811,N_17084,N_17752);
nand U22812 (N_22812,N_19586,N_15096);
xor U22813 (N_22813,N_16266,N_18105);
or U22814 (N_22814,N_19712,N_16626);
nor U22815 (N_22815,N_19658,N_17991);
xor U22816 (N_22816,N_18353,N_19605);
xnor U22817 (N_22817,N_18526,N_15417);
and U22818 (N_22818,N_16299,N_18791);
nor U22819 (N_22819,N_18107,N_15636);
and U22820 (N_22820,N_16383,N_15565);
nor U22821 (N_22821,N_19595,N_17329);
nand U22822 (N_22822,N_18972,N_19929);
and U22823 (N_22823,N_16472,N_16897);
or U22824 (N_22824,N_19906,N_15309);
nand U22825 (N_22825,N_16303,N_16635);
xnor U22826 (N_22826,N_17872,N_18190);
xor U22827 (N_22827,N_17609,N_18105);
nor U22828 (N_22828,N_18023,N_19576);
nand U22829 (N_22829,N_16829,N_16256);
or U22830 (N_22830,N_18952,N_17216);
or U22831 (N_22831,N_16266,N_15806);
nor U22832 (N_22832,N_15463,N_17797);
and U22833 (N_22833,N_19538,N_16389);
xnor U22834 (N_22834,N_16775,N_17205);
and U22835 (N_22835,N_19397,N_19632);
nand U22836 (N_22836,N_15020,N_15377);
xor U22837 (N_22837,N_18639,N_17947);
and U22838 (N_22838,N_16657,N_16899);
xnor U22839 (N_22839,N_17060,N_17042);
or U22840 (N_22840,N_16337,N_16615);
xor U22841 (N_22841,N_19412,N_15388);
nand U22842 (N_22842,N_19996,N_15758);
nand U22843 (N_22843,N_19010,N_19503);
or U22844 (N_22844,N_19560,N_16819);
and U22845 (N_22845,N_16263,N_16467);
nor U22846 (N_22846,N_18314,N_18647);
nand U22847 (N_22847,N_16485,N_15657);
nor U22848 (N_22848,N_18126,N_16217);
xnor U22849 (N_22849,N_19282,N_16732);
nand U22850 (N_22850,N_17038,N_16921);
xor U22851 (N_22851,N_18360,N_18404);
xor U22852 (N_22852,N_16408,N_17895);
nand U22853 (N_22853,N_18022,N_17733);
nand U22854 (N_22854,N_16056,N_16928);
nor U22855 (N_22855,N_19040,N_17342);
nor U22856 (N_22856,N_17943,N_19191);
xor U22857 (N_22857,N_15947,N_17432);
and U22858 (N_22858,N_17522,N_19544);
xor U22859 (N_22859,N_17466,N_17617);
nand U22860 (N_22860,N_15406,N_17921);
nand U22861 (N_22861,N_19539,N_17533);
and U22862 (N_22862,N_18825,N_16277);
nor U22863 (N_22863,N_19555,N_15007);
xor U22864 (N_22864,N_18573,N_18797);
or U22865 (N_22865,N_17041,N_19333);
nor U22866 (N_22866,N_16974,N_18189);
nor U22867 (N_22867,N_17440,N_16710);
or U22868 (N_22868,N_19631,N_17095);
or U22869 (N_22869,N_16906,N_16234);
and U22870 (N_22870,N_18163,N_16885);
and U22871 (N_22871,N_15621,N_15798);
nor U22872 (N_22872,N_16879,N_18314);
or U22873 (N_22873,N_17712,N_15614);
nand U22874 (N_22874,N_18270,N_17548);
nor U22875 (N_22875,N_18326,N_16906);
nand U22876 (N_22876,N_19227,N_16297);
or U22877 (N_22877,N_18836,N_16000);
xor U22878 (N_22878,N_15112,N_15348);
and U22879 (N_22879,N_19022,N_19709);
nor U22880 (N_22880,N_18524,N_18532);
nor U22881 (N_22881,N_15319,N_16891);
nor U22882 (N_22882,N_15503,N_15249);
or U22883 (N_22883,N_16456,N_17145);
nand U22884 (N_22884,N_15994,N_19066);
nor U22885 (N_22885,N_19438,N_16983);
and U22886 (N_22886,N_17208,N_19173);
xnor U22887 (N_22887,N_16019,N_16013);
xnor U22888 (N_22888,N_17107,N_16385);
nor U22889 (N_22889,N_16042,N_16162);
and U22890 (N_22890,N_19992,N_19506);
and U22891 (N_22891,N_15648,N_16657);
or U22892 (N_22892,N_18317,N_16876);
xor U22893 (N_22893,N_19865,N_19680);
nor U22894 (N_22894,N_15345,N_16643);
nor U22895 (N_22895,N_17855,N_15126);
and U22896 (N_22896,N_15671,N_17252);
or U22897 (N_22897,N_16870,N_17482);
or U22898 (N_22898,N_18309,N_17894);
nor U22899 (N_22899,N_19011,N_18313);
nor U22900 (N_22900,N_19598,N_18449);
or U22901 (N_22901,N_19123,N_19760);
or U22902 (N_22902,N_19412,N_16842);
nor U22903 (N_22903,N_15003,N_16439);
xnor U22904 (N_22904,N_16509,N_19373);
nor U22905 (N_22905,N_17063,N_17971);
xnor U22906 (N_22906,N_16062,N_18964);
nand U22907 (N_22907,N_19008,N_18770);
or U22908 (N_22908,N_15831,N_15249);
nor U22909 (N_22909,N_18397,N_15607);
nand U22910 (N_22910,N_19426,N_19907);
and U22911 (N_22911,N_19756,N_16954);
and U22912 (N_22912,N_15175,N_17898);
nand U22913 (N_22913,N_15300,N_18573);
xor U22914 (N_22914,N_16503,N_16659);
xor U22915 (N_22915,N_15474,N_19017);
or U22916 (N_22916,N_18690,N_16531);
nor U22917 (N_22917,N_15345,N_18161);
nand U22918 (N_22918,N_15940,N_17563);
xnor U22919 (N_22919,N_16912,N_16201);
nor U22920 (N_22920,N_18453,N_18392);
or U22921 (N_22921,N_16583,N_15472);
and U22922 (N_22922,N_16308,N_19808);
and U22923 (N_22923,N_19701,N_18703);
xnor U22924 (N_22924,N_19982,N_18225);
nor U22925 (N_22925,N_19883,N_18657);
nor U22926 (N_22926,N_17447,N_16430);
or U22927 (N_22927,N_19021,N_16316);
xnor U22928 (N_22928,N_16260,N_17695);
and U22929 (N_22929,N_15286,N_16379);
or U22930 (N_22930,N_17198,N_17474);
xnor U22931 (N_22931,N_15549,N_15248);
nand U22932 (N_22932,N_17883,N_17430);
nand U22933 (N_22933,N_16607,N_18158);
xnor U22934 (N_22934,N_16658,N_18575);
and U22935 (N_22935,N_17302,N_18320);
nand U22936 (N_22936,N_19674,N_16683);
or U22937 (N_22937,N_18995,N_15541);
and U22938 (N_22938,N_16160,N_16419);
and U22939 (N_22939,N_17420,N_19257);
nand U22940 (N_22940,N_18600,N_16234);
or U22941 (N_22941,N_18725,N_19382);
nand U22942 (N_22942,N_17745,N_16086);
nand U22943 (N_22943,N_17581,N_16687);
or U22944 (N_22944,N_15248,N_15386);
nor U22945 (N_22945,N_17515,N_19296);
xnor U22946 (N_22946,N_18605,N_19045);
nor U22947 (N_22947,N_15363,N_19846);
nor U22948 (N_22948,N_17690,N_15653);
nand U22949 (N_22949,N_16889,N_19370);
xor U22950 (N_22950,N_18717,N_19246);
xnor U22951 (N_22951,N_18928,N_18448);
xnor U22952 (N_22952,N_16967,N_19019);
nor U22953 (N_22953,N_15589,N_16074);
xnor U22954 (N_22954,N_17091,N_17465);
nand U22955 (N_22955,N_18213,N_19431);
nand U22956 (N_22956,N_17605,N_16091);
or U22957 (N_22957,N_18175,N_15083);
or U22958 (N_22958,N_18324,N_16317);
xnor U22959 (N_22959,N_15593,N_17982);
and U22960 (N_22960,N_17408,N_16704);
xor U22961 (N_22961,N_17826,N_17603);
and U22962 (N_22962,N_19975,N_19918);
nor U22963 (N_22963,N_17717,N_19980);
nor U22964 (N_22964,N_18962,N_18189);
nor U22965 (N_22965,N_15514,N_17982);
and U22966 (N_22966,N_18591,N_18801);
nand U22967 (N_22967,N_15559,N_17570);
nor U22968 (N_22968,N_17625,N_18850);
or U22969 (N_22969,N_18422,N_16150);
nor U22970 (N_22970,N_19800,N_18280);
or U22971 (N_22971,N_17999,N_18288);
xor U22972 (N_22972,N_15667,N_18872);
nor U22973 (N_22973,N_15068,N_15019);
and U22974 (N_22974,N_17151,N_19746);
nor U22975 (N_22975,N_16752,N_18940);
nand U22976 (N_22976,N_15075,N_15601);
nor U22977 (N_22977,N_17498,N_18125);
or U22978 (N_22978,N_17738,N_18649);
nor U22979 (N_22979,N_17812,N_18222);
nor U22980 (N_22980,N_17521,N_18423);
and U22981 (N_22981,N_19411,N_16205);
nor U22982 (N_22982,N_16479,N_16314);
nor U22983 (N_22983,N_17721,N_19129);
nand U22984 (N_22984,N_18172,N_18538);
or U22985 (N_22985,N_15092,N_17591);
xnor U22986 (N_22986,N_15503,N_15885);
or U22987 (N_22987,N_16062,N_18758);
nand U22988 (N_22988,N_17206,N_16904);
and U22989 (N_22989,N_17425,N_16826);
nor U22990 (N_22990,N_19323,N_15075);
nand U22991 (N_22991,N_15277,N_18657);
xor U22992 (N_22992,N_19634,N_19580);
xor U22993 (N_22993,N_15147,N_17805);
nand U22994 (N_22994,N_19991,N_19454);
nor U22995 (N_22995,N_19925,N_17905);
nand U22996 (N_22996,N_18047,N_15797);
nor U22997 (N_22997,N_15444,N_17208);
nand U22998 (N_22998,N_19581,N_16315);
or U22999 (N_22999,N_18316,N_18926);
nand U23000 (N_23000,N_18624,N_18512);
nor U23001 (N_23001,N_19167,N_18917);
and U23002 (N_23002,N_17028,N_15306);
nor U23003 (N_23003,N_16305,N_19784);
and U23004 (N_23004,N_17292,N_19689);
nand U23005 (N_23005,N_16561,N_18856);
nor U23006 (N_23006,N_15748,N_18866);
or U23007 (N_23007,N_16439,N_15792);
and U23008 (N_23008,N_15060,N_17442);
xnor U23009 (N_23009,N_16386,N_16777);
xnor U23010 (N_23010,N_18595,N_15658);
nand U23011 (N_23011,N_16157,N_18715);
and U23012 (N_23012,N_15178,N_19716);
and U23013 (N_23013,N_17994,N_18920);
or U23014 (N_23014,N_18179,N_15992);
or U23015 (N_23015,N_15980,N_15212);
or U23016 (N_23016,N_15986,N_18486);
nand U23017 (N_23017,N_16910,N_15541);
nand U23018 (N_23018,N_16828,N_16928);
and U23019 (N_23019,N_16533,N_16170);
and U23020 (N_23020,N_15712,N_19900);
and U23021 (N_23021,N_18757,N_15305);
xor U23022 (N_23022,N_17053,N_17287);
nand U23023 (N_23023,N_16964,N_15507);
nand U23024 (N_23024,N_18696,N_19646);
or U23025 (N_23025,N_16916,N_16044);
or U23026 (N_23026,N_17858,N_15412);
nor U23027 (N_23027,N_19875,N_18334);
and U23028 (N_23028,N_17007,N_18568);
and U23029 (N_23029,N_19931,N_18922);
xnor U23030 (N_23030,N_19406,N_16016);
nand U23031 (N_23031,N_19474,N_17009);
xnor U23032 (N_23032,N_17684,N_18735);
nand U23033 (N_23033,N_17953,N_19174);
and U23034 (N_23034,N_16963,N_17448);
nor U23035 (N_23035,N_19003,N_18807);
nor U23036 (N_23036,N_19403,N_19307);
nand U23037 (N_23037,N_18434,N_18683);
nor U23038 (N_23038,N_17284,N_17535);
and U23039 (N_23039,N_17701,N_19290);
or U23040 (N_23040,N_17540,N_18188);
or U23041 (N_23041,N_16589,N_16773);
or U23042 (N_23042,N_15789,N_15192);
and U23043 (N_23043,N_15093,N_15504);
nand U23044 (N_23044,N_19626,N_19445);
nor U23045 (N_23045,N_18547,N_19114);
and U23046 (N_23046,N_18027,N_19064);
xnor U23047 (N_23047,N_17349,N_17631);
xnor U23048 (N_23048,N_18443,N_19484);
xor U23049 (N_23049,N_18356,N_18612);
nor U23050 (N_23050,N_17344,N_19147);
nor U23051 (N_23051,N_18653,N_17151);
and U23052 (N_23052,N_16292,N_15035);
xnor U23053 (N_23053,N_19031,N_15995);
or U23054 (N_23054,N_18848,N_19461);
or U23055 (N_23055,N_19452,N_15487);
nor U23056 (N_23056,N_17534,N_19474);
nor U23057 (N_23057,N_16632,N_19222);
nor U23058 (N_23058,N_19982,N_19393);
nand U23059 (N_23059,N_17591,N_16864);
nand U23060 (N_23060,N_16245,N_16204);
nor U23061 (N_23061,N_16491,N_17364);
xor U23062 (N_23062,N_18252,N_17684);
or U23063 (N_23063,N_18904,N_17155);
xnor U23064 (N_23064,N_15632,N_18510);
nand U23065 (N_23065,N_17764,N_19495);
nand U23066 (N_23066,N_16888,N_17024);
and U23067 (N_23067,N_17696,N_18845);
or U23068 (N_23068,N_17474,N_19598);
or U23069 (N_23069,N_16573,N_15539);
or U23070 (N_23070,N_19957,N_18323);
xnor U23071 (N_23071,N_17638,N_18753);
xnor U23072 (N_23072,N_18056,N_15570);
nand U23073 (N_23073,N_17085,N_18761);
and U23074 (N_23074,N_15081,N_18725);
nand U23075 (N_23075,N_19400,N_15165);
or U23076 (N_23076,N_16516,N_18387);
and U23077 (N_23077,N_18256,N_15694);
xor U23078 (N_23078,N_16044,N_18523);
and U23079 (N_23079,N_18709,N_15194);
and U23080 (N_23080,N_18864,N_15228);
and U23081 (N_23081,N_16537,N_16658);
nand U23082 (N_23082,N_15532,N_18491);
xor U23083 (N_23083,N_19398,N_19657);
nor U23084 (N_23084,N_15444,N_17487);
xnor U23085 (N_23085,N_19527,N_18633);
and U23086 (N_23086,N_19458,N_16082);
nor U23087 (N_23087,N_17970,N_16287);
and U23088 (N_23088,N_15709,N_17970);
nand U23089 (N_23089,N_18666,N_16923);
and U23090 (N_23090,N_19633,N_16621);
nor U23091 (N_23091,N_16978,N_18012);
nand U23092 (N_23092,N_16935,N_16018);
xor U23093 (N_23093,N_19387,N_17587);
or U23094 (N_23094,N_18282,N_17884);
and U23095 (N_23095,N_18417,N_17372);
nor U23096 (N_23096,N_15024,N_19123);
and U23097 (N_23097,N_15222,N_17564);
and U23098 (N_23098,N_16844,N_15943);
and U23099 (N_23099,N_16325,N_16878);
and U23100 (N_23100,N_16798,N_16132);
xnor U23101 (N_23101,N_17329,N_19483);
xnor U23102 (N_23102,N_18330,N_15827);
nand U23103 (N_23103,N_16381,N_17792);
nand U23104 (N_23104,N_18365,N_17754);
or U23105 (N_23105,N_15360,N_18356);
xor U23106 (N_23106,N_18113,N_17892);
or U23107 (N_23107,N_19355,N_15362);
and U23108 (N_23108,N_16743,N_15150);
nor U23109 (N_23109,N_16389,N_16126);
or U23110 (N_23110,N_17886,N_19983);
nor U23111 (N_23111,N_16799,N_18537);
and U23112 (N_23112,N_18038,N_15383);
nand U23113 (N_23113,N_18541,N_15434);
and U23114 (N_23114,N_15501,N_16563);
xor U23115 (N_23115,N_16402,N_15696);
and U23116 (N_23116,N_18672,N_19684);
and U23117 (N_23117,N_18017,N_19311);
or U23118 (N_23118,N_15934,N_18666);
xor U23119 (N_23119,N_17744,N_16850);
or U23120 (N_23120,N_19296,N_16220);
nor U23121 (N_23121,N_16091,N_19859);
or U23122 (N_23122,N_18939,N_17039);
or U23123 (N_23123,N_17433,N_16066);
nor U23124 (N_23124,N_19282,N_19922);
xor U23125 (N_23125,N_16112,N_15538);
or U23126 (N_23126,N_17803,N_15184);
and U23127 (N_23127,N_19446,N_16133);
nand U23128 (N_23128,N_16786,N_17025);
nor U23129 (N_23129,N_19988,N_16654);
nor U23130 (N_23130,N_18067,N_18849);
nor U23131 (N_23131,N_19740,N_18975);
nand U23132 (N_23132,N_19353,N_19970);
or U23133 (N_23133,N_18261,N_18165);
and U23134 (N_23134,N_15755,N_16421);
nor U23135 (N_23135,N_15263,N_15971);
or U23136 (N_23136,N_15037,N_19983);
nor U23137 (N_23137,N_18686,N_18563);
xnor U23138 (N_23138,N_18026,N_16531);
or U23139 (N_23139,N_16739,N_18079);
xor U23140 (N_23140,N_16573,N_17631);
nand U23141 (N_23141,N_16765,N_19278);
xor U23142 (N_23142,N_18178,N_15631);
xnor U23143 (N_23143,N_19541,N_15082);
xor U23144 (N_23144,N_17382,N_16607);
nor U23145 (N_23145,N_15007,N_16346);
and U23146 (N_23146,N_18698,N_19117);
or U23147 (N_23147,N_17753,N_16404);
nand U23148 (N_23148,N_15861,N_16770);
and U23149 (N_23149,N_18199,N_15765);
or U23150 (N_23150,N_16517,N_19959);
nand U23151 (N_23151,N_16499,N_16733);
xor U23152 (N_23152,N_19587,N_15584);
nand U23153 (N_23153,N_19182,N_15543);
and U23154 (N_23154,N_18582,N_15413);
nor U23155 (N_23155,N_18295,N_18348);
or U23156 (N_23156,N_17846,N_18693);
and U23157 (N_23157,N_18147,N_19336);
nand U23158 (N_23158,N_19441,N_16927);
xor U23159 (N_23159,N_15471,N_15732);
nor U23160 (N_23160,N_17832,N_18720);
xor U23161 (N_23161,N_15201,N_16627);
or U23162 (N_23162,N_19800,N_19534);
nor U23163 (N_23163,N_17563,N_18948);
or U23164 (N_23164,N_19095,N_15190);
and U23165 (N_23165,N_16320,N_15845);
xnor U23166 (N_23166,N_15827,N_17628);
xnor U23167 (N_23167,N_18555,N_19611);
nand U23168 (N_23168,N_18110,N_16602);
and U23169 (N_23169,N_15549,N_19872);
or U23170 (N_23170,N_15757,N_16159);
and U23171 (N_23171,N_16507,N_19495);
xor U23172 (N_23172,N_16228,N_19204);
xnor U23173 (N_23173,N_16965,N_16341);
nor U23174 (N_23174,N_19418,N_15190);
xor U23175 (N_23175,N_15466,N_18585);
nand U23176 (N_23176,N_18346,N_16029);
or U23177 (N_23177,N_15471,N_18547);
xnor U23178 (N_23178,N_19487,N_17620);
nand U23179 (N_23179,N_19996,N_18184);
nand U23180 (N_23180,N_18106,N_16047);
and U23181 (N_23181,N_16814,N_18213);
or U23182 (N_23182,N_19899,N_15178);
and U23183 (N_23183,N_15057,N_15549);
and U23184 (N_23184,N_15044,N_15203);
and U23185 (N_23185,N_17238,N_16776);
or U23186 (N_23186,N_16458,N_17980);
nand U23187 (N_23187,N_19318,N_15211);
or U23188 (N_23188,N_18042,N_18885);
and U23189 (N_23189,N_17412,N_17800);
nand U23190 (N_23190,N_17986,N_16508);
xor U23191 (N_23191,N_16829,N_16963);
nand U23192 (N_23192,N_18211,N_16832);
nand U23193 (N_23193,N_18876,N_15736);
nor U23194 (N_23194,N_18710,N_19609);
nor U23195 (N_23195,N_18725,N_19660);
or U23196 (N_23196,N_16052,N_17640);
and U23197 (N_23197,N_17957,N_15574);
nand U23198 (N_23198,N_19842,N_17527);
nand U23199 (N_23199,N_18772,N_19041);
xnor U23200 (N_23200,N_19895,N_17286);
xnor U23201 (N_23201,N_16304,N_17997);
and U23202 (N_23202,N_16462,N_17584);
and U23203 (N_23203,N_15870,N_18275);
and U23204 (N_23204,N_19051,N_16543);
or U23205 (N_23205,N_15371,N_16904);
or U23206 (N_23206,N_18142,N_15772);
nand U23207 (N_23207,N_19582,N_17693);
or U23208 (N_23208,N_16612,N_16503);
xor U23209 (N_23209,N_17572,N_16718);
and U23210 (N_23210,N_16060,N_16025);
nand U23211 (N_23211,N_15240,N_16052);
or U23212 (N_23212,N_15314,N_17031);
xor U23213 (N_23213,N_15775,N_18219);
nor U23214 (N_23214,N_19460,N_16840);
or U23215 (N_23215,N_17156,N_18091);
nand U23216 (N_23216,N_15338,N_18728);
xor U23217 (N_23217,N_16198,N_16479);
xor U23218 (N_23218,N_19323,N_15675);
or U23219 (N_23219,N_16636,N_16821);
or U23220 (N_23220,N_19745,N_19457);
and U23221 (N_23221,N_17458,N_16152);
nor U23222 (N_23222,N_15805,N_17178);
and U23223 (N_23223,N_16781,N_17345);
nor U23224 (N_23224,N_18972,N_18542);
nand U23225 (N_23225,N_16262,N_17378);
nand U23226 (N_23226,N_16112,N_16430);
or U23227 (N_23227,N_19020,N_15774);
nand U23228 (N_23228,N_19702,N_15115);
and U23229 (N_23229,N_16435,N_19795);
and U23230 (N_23230,N_19049,N_18786);
xnor U23231 (N_23231,N_17505,N_17349);
nand U23232 (N_23232,N_19681,N_19575);
or U23233 (N_23233,N_15597,N_15915);
or U23234 (N_23234,N_17985,N_15275);
or U23235 (N_23235,N_17808,N_19699);
xor U23236 (N_23236,N_18615,N_16168);
or U23237 (N_23237,N_18527,N_17696);
nand U23238 (N_23238,N_15370,N_16471);
xnor U23239 (N_23239,N_15408,N_16140);
xnor U23240 (N_23240,N_19913,N_16658);
nand U23241 (N_23241,N_17899,N_17781);
and U23242 (N_23242,N_17428,N_16974);
nor U23243 (N_23243,N_19314,N_19066);
and U23244 (N_23244,N_15582,N_19469);
xnor U23245 (N_23245,N_18598,N_18580);
xnor U23246 (N_23246,N_17754,N_18818);
or U23247 (N_23247,N_19240,N_15251);
nor U23248 (N_23248,N_16812,N_16710);
xor U23249 (N_23249,N_16360,N_16661);
nand U23250 (N_23250,N_18094,N_17646);
and U23251 (N_23251,N_16713,N_16398);
and U23252 (N_23252,N_18732,N_19548);
nor U23253 (N_23253,N_15715,N_16278);
and U23254 (N_23254,N_15309,N_19614);
xor U23255 (N_23255,N_18872,N_17465);
and U23256 (N_23256,N_17922,N_17090);
or U23257 (N_23257,N_16952,N_18677);
nor U23258 (N_23258,N_15367,N_15046);
nor U23259 (N_23259,N_17014,N_16794);
and U23260 (N_23260,N_15346,N_18861);
or U23261 (N_23261,N_19192,N_19454);
and U23262 (N_23262,N_15402,N_19877);
nand U23263 (N_23263,N_15764,N_17525);
nor U23264 (N_23264,N_16012,N_19427);
xor U23265 (N_23265,N_17462,N_17129);
nand U23266 (N_23266,N_18707,N_18467);
xor U23267 (N_23267,N_17196,N_18661);
and U23268 (N_23268,N_19919,N_15538);
or U23269 (N_23269,N_18256,N_16977);
nand U23270 (N_23270,N_16338,N_15230);
nor U23271 (N_23271,N_19007,N_17819);
or U23272 (N_23272,N_16316,N_16417);
nor U23273 (N_23273,N_15074,N_15946);
or U23274 (N_23274,N_18736,N_16541);
or U23275 (N_23275,N_16556,N_16038);
and U23276 (N_23276,N_19502,N_18810);
xor U23277 (N_23277,N_17272,N_18341);
and U23278 (N_23278,N_15016,N_19405);
xnor U23279 (N_23279,N_16865,N_15762);
and U23280 (N_23280,N_19288,N_19379);
xnor U23281 (N_23281,N_18921,N_19706);
nor U23282 (N_23282,N_18812,N_16536);
xor U23283 (N_23283,N_19360,N_16243);
and U23284 (N_23284,N_15922,N_17075);
xnor U23285 (N_23285,N_16730,N_19744);
or U23286 (N_23286,N_16194,N_16321);
xnor U23287 (N_23287,N_17169,N_18382);
and U23288 (N_23288,N_19031,N_16907);
and U23289 (N_23289,N_15270,N_19633);
and U23290 (N_23290,N_19719,N_15480);
nor U23291 (N_23291,N_19970,N_15009);
and U23292 (N_23292,N_17557,N_19055);
xnor U23293 (N_23293,N_16986,N_17623);
nand U23294 (N_23294,N_19141,N_19904);
nand U23295 (N_23295,N_15462,N_17079);
or U23296 (N_23296,N_15545,N_15726);
xor U23297 (N_23297,N_19183,N_15959);
or U23298 (N_23298,N_18206,N_17864);
or U23299 (N_23299,N_18651,N_18114);
nand U23300 (N_23300,N_16349,N_18769);
xnor U23301 (N_23301,N_15624,N_19341);
nor U23302 (N_23302,N_16283,N_18532);
and U23303 (N_23303,N_18986,N_18624);
and U23304 (N_23304,N_16041,N_17660);
or U23305 (N_23305,N_18676,N_18956);
xnor U23306 (N_23306,N_17492,N_18060);
nand U23307 (N_23307,N_18096,N_17837);
nor U23308 (N_23308,N_16231,N_17253);
or U23309 (N_23309,N_18638,N_15051);
nand U23310 (N_23310,N_15307,N_18080);
xor U23311 (N_23311,N_18762,N_19454);
or U23312 (N_23312,N_18638,N_17298);
nand U23313 (N_23313,N_19704,N_16522);
xor U23314 (N_23314,N_16760,N_19015);
xnor U23315 (N_23315,N_15188,N_19463);
and U23316 (N_23316,N_19855,N_16756);
nor U23317 (N_23317,N_17618,N_19521);
nand U23318 (N_23318,N_16588,N_18925);
xor U23319 (N_23319,N_19695,N_16537);
xnor U23320 (N_23320,N_19624,N_18771);
xor U23321 (N_23321,N_18154,N_15144);
nand U23322 (N_23322,N_19748,N_19936);
nand U23323 (N_23323,N_17229,N_17445);
xor U23324 (N_23324,N_19410,N_18975);
nand U23325 (N_23325,N_16658,N_19381);
or U23326 (N_23326,N_18201,N_19773);
nand U23327 (N_23327,N_19316,N_19880);
and U23328 (N_23328,N_19571,N_16997);
nor U23329 (N_23329,N_18753,N_16039);
xnor U23330 (N_23330,N_19603,N_15424);
or U23331 (N_23331,N_15910,N_15652);
nand U23332 (N_23332,N_19671,N_17401);
nand U23333 (N_23333,N_15717,N_18196);
or U23334 (N_23334,N_15548,N_16681);
nand U23335 (N_23335,N_15490,N_19396);
nand U23336 (N_23336,N_19657,N_18187);
xnor U23337 (N_23337,N_19171,N_17221);
and U23338 (N_23338,N_16690,N_16298);
or U23339 (N_23339,N_16166,N_16184);
and U23340 (N_23340,N_17705,N_17600);
nor U23341 (N_23341,N_18774,N_17877);
nor U23342 (N_23342,N_16546,N_15809);
xor U23343 (N_23343,N_15700,N_15313);
nor U23344 (N_23344,N_15485,N_18274);
xnor U23345 (N_23345,N_19966,N_15194);
xor U23346 (N_23346,N_17515,N_15461);
and U23347 (N_23347,N_15430,N_15654);
and U23348 (N_23348,N_18651,N_18022);
nor U23349 (N_23349,N_18698,N_17061);
nor U23350 (N_23350,N_18980,N_17761);
nand U23351 (N_23351,N_19698,N_16906);
and U23352 (N_23352,N_19723,N_18796);
nor U23353 (N_23353,N_17538,N_15697);
nand U23354 (N_23354,N_19113,N_18906);
nor U23355 (N_23355,N_16809,N_15021);
xnor U23356 (N_23356,N_16498,N_19075);
nand U23357 (N_23357,N_15243,N_17617);
and U23358 (N_23358,N_15098,N_18896);
or U23359 (N_23359,N_19774,N_15393);
nor U23360 (N_23360,N_19376,N_15722);
and U23361 (N_23361,N_18147,N_16414);
nand U23362 (N_23362,N_19571,N_19466);
or U23363 (N_23363,N_19578,N_17432);
nand U23364 (N_23364,N_16589,N_17847);
or U23365 (N_23365,N_19517,N_15440);
nand U23366 (N_23366,N_19532,N_16519);
or U23367 (N_23367,N_16699,N_16914);
xnor U23368 (N_23368,N_15470,N_18637);
nor U23369 (N_23369,N_19588,N_17484);
nor U23370 (N_23370,N_18865,N_16610);
or U23371 (N_23371,N_16942,N_16152);
or U23372 (N_23372,N_17724,N_17323);
nand U23373 (N_23373,N_17654,N_17873);
and U23374 (N_23374,N_19777,N_18351);
nand U23375 (N_23375,N_15969,N_18436);
nand U23376 (N_23376,N_16994,N_15539);
xor U23377 (N_23377,N_17657,N_15444);
nor U23378 (N_23378,N_15413,N_15184);
xor U23379 (N_23379,N_18011,N_19476);
nor U23380 (N_23380,N_15908,N_18202);
nand U23381 (N_23381,N_17745,N_19766);
nand U23382 (N_23382,N_17394,N_16253);
xnor U23383 (N_23383,N_19864,N_19470);
nand U23384 (N_23384,N_17126,N_15039);
or U23385 (N_23385,N_18653,N_19941);
xnor U23386 (N_23386,N_18279,N_15328);
or U23387 (N_23387,N_16041,N_16109);
nor U23388 (N_23388,N_19827,N_17869);
nor U23389 (N_23389,N_17754,N_18738);
or U23390 (N_23390,N_15142,N_17362);
xnor U23391 (N_23391,N_15673,N_15921);
nor U23392 (N_23392,N_16405,N_18280);
and U23393 (N_23393,N_18608,N_17107);
nor U23394 (N_23394,N_15328,N_15195);
or U23395 (N_23395,N_16087,N_17887);
xnor U23396 (N_23396,N_18302,N_18142);
or U23397 (N_23397,N_15800,N_15011);
nand U23398 (N_23398,N_19677,N_19707);
xnor U23399 (N_23399,N_18890,N_18981);
xor U23400 (N_23400,N_19817,N_17253);
nor U23401 (N_23401,N_16212,N_19535);
nor U23402 (N_23402,N_18287,N_18495);
or U23403 (N_23403,N_18285,N_18524);
nor U23404 (N_23404,N_16491,N_18817);
nand U23405 (N_23405,N_17930,N_17377);
nand U23406 (N_23406,N_15811,N_18589);
and U23407 (N_23407,N_17121,N_16279);
nor U23408 (N_23408,N_18985,N_15381);
or U23409 (N_23409,N_17157,N_18200);
nand U23410 (N_23410,N_17952,N_17670);
or U23411 (N_23411,N_16627,N_16439);
xnor U23412 (N_23412,N_15734,N_19646);
nor U23413 (N_23413,N_19566,N_18654);
and U23414 (N_23414,N_15859,N_18147);
and U23415 (N_23415,N_16514,N_15418);
xnor U23416 (N_23416,N_16315,N_17697);
and U23417 (N_23417,N_17840,N_17790);
and U23418 (N_23418,N_17494,N_16555);
and U23419 (N_23419,N_16442,N_19246);
and U23420 (N_23420,N_19422,N_16952);
nor U23421 (N_23421,N_19513,N_18704);
and U23422 (N_23422,N_17869,N_18570);
nand U23423 (N_23423,N_18901,N_17103);
nand U23424 (N_23424,N_16854,N_15536);
nor U23425 (N_23425,N_17094,N_17519);
and U23426 (N_23426,N_16033,N_19648);
nor U23427 (N_23427,N_15651,N_17407);
or U23428 (N_23428,N_18118,N_17213);
or U23429 (N_23429,N_16742,N_18120);
or U23430 (N_23430,N_16203,N_16620);
xor U23431 (N_23431,N_19954,N_19530);
nor U23432 (N_23432,N_18072,N_16428);
or U23433 (N_23433,N_15968,N_16746);
or U23434 (N_23434,N_16205,N_18056);
and U23435 (N_23435,N_15193,N_19949);
and U23436 (N_23436,N_17983,N_16934);
xor U23437 (N_23437,N_17963,N_15861);
and U23438 (N_23438,N_17737,N_18170);
nor U23439 (N_23439,N_18771,N_16842);
nor U23440 (N_23440,N_15629,N_18575);
xnor U23441 (N_23441,N_15084,N_15816);
nand U23442 (N_23442,N_18533,N_17293);
and U23443 (N_23443,N_16964,N_15790);
nor U23444 (N_23444,N_19241,N_15674);
or U23445 (N_23445,N_19853,N_16583);
and U23446 (N_23446,N_17884,N_15819);
and U23447 (N_23447,N_16066,N_17876);
xor U23448 (N_23448,N_16180,N_17953);
nor U23449 (N_23449,N_15420,N_18750);
nand U23450 (N_23450,N_18497,N_15251);
nand U23451 (N_23451,N_19163,N_15885);
nor U23452 (N_23452,N_16814,N_19915);
xor U23453 (N_23453,N_17488,N_15938);
nor U23454 (N_23454,N_19201,N_15340);
nand U23455 (N_23455,N_17769,N_16057);
nand U23456 (N_23456,N_19879,N_17601);
nand U23457 (N_23457,N_19817,N_16423);
xnor U23458 (N_23458,N_15202,N_19714);
nand U23459 (N_23459,N_18925,N_18042);
xor U23460 (N_23460,N_17667,N_19270);
nor U23461 (N_23461,N_18269,N_17682);
or U23462 (N_23462,N_19556,N_15843);
nor U23463 (N_23463,N_18711,N_17133);
or U23464 (N_23464,N_18680,N_15366);
xnor U23465 (N_23465,N_18594,N_15718);
or U23466 (N_23466,N_18049,N_19930);
and U23467 (N_23467,N_17307,N_18557);
nand U23468 (N_23468,N_16890,N_19276);
or U23469 (N_23469,N_17192,N_18551);
or U23470 (N_23470,N_16891,N_19010);
nand U23471 (N_23471,N_17778,N_16954);
xnor U23472 (N_23472,N_16612,N_18950);
or U23473 (N_23473,N_19527,N_15514);
xnor U23474 (N_23474,N_17180,N_19954);
nor U23475 (N_23475,N_19730,N_16407);
nor U23476 (N_23476,N_19052,N_18415);
or U23477 (N_23477,N_19279,N_15511);
xor U23478 (N_23478,N_16465,N_18258);
nand U23479 (N_23479,N_15823,N_18466);
nor U23480 (N_23480,N_16504,N_19646);
nor U23481 (N_23481,N_16131,N_17336);
xnor U23482 (N_23482,N_15805,N_17405);
nor U23483 (N_23483,N_15833,N_19979);
nand U23484 (N_23484,N_19919,N_15423);
nand U23485 (N_23485,N_18180,N_19335);
and U23486 (N_23486,N_16650,N_18297);
nand U23487 (N_23487,N_16738,N_17244);
nand U23488 (N_23488,N_18973,N_16018);
xnor U23489 (N_23489,N_19084,N_19852);
and U23490 (N_23490,N_15916,N_15103);
nor U23491 (N_23491,N_15904,N_17420);
nor U23492 (N_23492,N_19160,N_16252);
and U23493 (N_23493,N_17514,N_18073);
or U23494 (N_23494,N_18007,N_16854);
or U23495 (N_23495,N_16862,N_17913);
or U23496 (N_23496,N_15504,N_19072);
xnor U23497 (N_23497,N_16500,N_16087);
and U23498 (N_23498,N_17283,N_15582);
nor U23499 (N_23499,N_15631,N_18043);
nor U23500 (N_23500,N_16919,N_17954);
or U23501 (N_23501,N_18236,N_16664);
nand U23502 (N_23502,N_19001,N_19893);
and U23503 (N_23503,N_15449,N_15206);
or U23504 (N_23504,N_15342,N_19180);
nor U23505 (N_23505,N_18477,N_16090);
nor U23506 (N_23506,N_15351,N_18132);
nand U23507 (N_23507,N_16657,N_18549);
nor U23508 (N_23508,N_16123,N_16214);
nand U23509 (N_23509,N_17959,N_16921);
or U23510 (N_23510,N_18618,N_18593);
or U23511 (N_23511,N_15732,N_19610);
and U23512 (N_23512,N_17818,N_16060);
xnor U23513 (N_23513,N_17657,N_17848);
or U23514 (N_23514,N_19129,N_16742);
nand U23515 (N_23515,N_16838,N_15098);
and U23516 (N_23516,N_18821,N_19260);
xnor U23517 (N_23517,N_17220,N_15297);
and U23518 (N_23518,N_16139,N_19564);
nor U23519 (N_23519,N_16439,N_18307);
and U23520 (N_23520,N_16112,N_19075);
and U23521 (N_23521,N_15914,N_17392);
nand U23522 (N_23522,N_18072,N_15972);
or U23523 (N_23523,N_18943,N_19429);
nor U23524 (N_23524,N_17790,N_15558);
nand U23525 (N_23525,N_19137,N_15597);
or U23526 (N_23526,N_17728,N_18661);
nor U23527 (N_23527,N_15888,N_15416);
nor U23528 (N_23528,N_17055,N_18088);
nor U23529 (N_23529,N_15173,N_19935);
nor U23530 (N_23530,N_15881,N_15045);
xnor U23531 (N_23531,N_17318,N_18414);
nand U23532 (N_23532,N_16575,N_15716);
or U23533 (N_23533,N_15931,N_15682);
nor U23534 (N_23534,N_16340,N_15662);
and U23535 (N_23535,N_17753,N_15329);
nand U23536 (N_23536,N_19934,N_16853);
nor U23537 (N_23537,N_16333,N_17816);
or U23538 (N_23538,N_17682,N_19616);
or U23539 (N_23539,N_19970,N_16499);
and U23540 (N_23540,N_19521,N_15195);
nand U23541 (N_23541,N_15073,N_16695);
nand U23542 (N_23542,N_16127,N_18403);
or U23543 (N_23543,N_19857,N_19948);
nand U23544 (N_23544,N_18339,N_15903);
or U23545 (N_23545,N_17316,N_17497);
nand U23546 (N_23546,N_17918,N_17772);
or U23547 (N_23547,N_17075,N_19067);
nor U23548 (N_23548,N_17599,N_15080);
or U23549 (N_23549,N_19893,N_16045);
and U23550 (N_23550,N_19563,N_15645);
and U23551 (N_23551,N_16719,N_17486);
xnor U23552 (N_23552,N_16370,N_17062);
xor U23553 (N_23553,N_17887,N_16632);
and U23554 (N_23554,N_16492,N_15745);
or U23555 (N_23555,N_19970,N_16491);
nor U23556 (N_23556,N_18921,N_15232);
and U23557 (N_23557,N_18867,N_17425);
and U23558 (N_23558,N_18137,N_16030);
and U23559 (N_23559,N_15645,N_18118);
and U23560 (N_23560,N_19114,N_18312);
nand U23561 (N_23561,N_15311,N_19797);
or U23562 (N_23562,N_15484,N_16872);
and U23563 (N_23563,N_16884,N_16440);
nor U23564 (N_23564,N_18850,N_18844);
nand U23565 (N_23565,N_15328,N_19506);
or U23566 (N_23566,N_17608,N_16847);
and U23567 (N_23567,N_15624,N_18400);
xnor U23568 (N_23568,N_19840,N_18935);
xnor U23569 (N_23569,N_19655,N_19171);
nor U23570 (N_23570,N_17916,N_15315);
xor U23571 (N_23571,N_17507,N_17246);
or U23572 (N_23572,N_18812,N_16862);
xor U23573 (N_23573,N_19626,N_16300);
and U23574 (N_23574,N_19524,N_16618);
and U23575 (N_23575,N_18292,N_15740);
nor U23576 (N_23576,N_16463,N_19277);
nand U23577 (N_23577,N_16438,N_18781);
and U23578 (N_23578,N_16469,N_19055);
nor U23579 (N_23579,N_19267,N_19229);
and U23580 (N_23580,N_17573,N_18695);
or U23581 (N_23581,N_17241,N_15458);
nor U23582 (N_23582,N_15990,N_15771);
nand U23583 (N_23583,N_17613,N_16220);
or U23584 (N_23584,N_16515,N_18943);
nor U23585 (N_23585,N_18596,N_19271);
or U23586 (N_23586,N_19936,N_18420);
nor U23587 (N_23587,N_15089,N_17487);
and U23588 (N_23588,N_17448,N_16763);
or U23589 (N_23589,N_17421,N_17797);
and U23590 (N_23590,N_15271,N_18137);
and U23591 (N_23591,N_15459,N_16770);
xor U23592 (N_23592,N_15611,N_15744);
xor U23593 (N_23593,N_17658,N_18165);
or U23594 (N_23594,N_19014,N_17859);
nand U23595 (N_23595,N_19256,N_18190);
or U23596 (N_23596,N_15243,N_17315);
xor U23597 (N_23597,N_17859,N_17281);
and U23598 (N_23598,N_15079,N_17473);
and U23599 (N_23599,N_17085,N_16162);
nand U23600 (N_23600,N_17023,N_15049);
or U23601 (N_23601,N_15996,N_15329);
nor U23602 (N_23602,N_19117,N_15260);
or U23603 (N_23603,N_15021,N_19678);
nor U23604 (N_23604,N_19013,N_17656);
xnor U23605 (N_23605,N_19674,N_17213);
nand U23606 (N_23606,N_15028,N_15102);
or U23607 (N_23607,N_15867,N_15315);
and U23608 (N_23608,N_15498,N_16849);
or U23609 (N_23609,N_15475,N_19803);
nor U23610 (N_23610,N_16864,N_18981);
nor U23611 (N_23611,N_17673,N_19237);
and U23612 (N_23612,N_19980,N_19890);
xnor U23613 (N_23613,N_16540,N_19042);
or U23614 (N_23614,N_15469,N_16200);
xnor U23615 (N_23615,N_17778,N_19142);
xnor U23616 (N_23616,N_17508,N_16281);
xnor U23617 (N_23617,N_15130,N_16294);
nand U23618 (N_23618,N_19308,N_18771);
nor U23619 (N_23619,N_18392,N_18148);
or U23620 (N_23620,N_18534,N_18767);
and U23621 (N_23621,N_18619,N_16706);
nand U23622 (N_23622,N_16772,N_19172);
nor U23623 (N_23623,N_16691,N_19665);
and U23624 (N_23624,N_16984,N_18079);
or U23625 (N_23625,N_15900,N_19417);
nor U23626 (N_23626,N_19804,N_19639);
or U23627 (N_23627,N_19853,N_15915);
nor U23628 (N_23628,N_15450,N_18175);
nand U23629 (N_23629,N_16440,N_16546);
xor U23630 (N_23630,N_19894,N_16145);
xor U23631 (N_23631,N_17740,N_17536);
or U23632 (N_23632,N_17961,N_19522);
or U23633 (N_23633,N_17412,N_19813);
nor U23634 (N_23634,N_17110,N_19356);
nor U23635 (N_23635,N_17252,N_16456);
xor U23636 (N_23636,N_19583,N_16387);
xnor U23637 (N_23637,N_17587,N_16999);
nor U23638 (N_23638,N_18210,N_15078);
xor U23639 (N_23639,N_15384,N_17399);
xor U23640 (N_23640,N_16388,N_17049);
xor U23641 (N_23641,N_18471,N_19639);
and U23642 (N_23642,N_18564,N_15309);
and U23643 (N_23643,N_16052,N_16820);
xnor U23644 (N_23644,N_15091,N_18219);
nand U23645 (N_23645,N_17114,N_15285);
or U23646 (N_23646,N_16299,N_19048);
and U23647 (N_23647,N_15555,N_16060);
or U23648 (N_23648,N_15377,N_17187);
xor U23649 (N_23649,N_16917,N_19739);
and U23650 (N_23650,N_18140,N_17229);
nor U23651 (N_23651,N_16739,N_18448);
xnor U23652 (N_23652,N_17321,N_19622);
and U23653 (N_23653,N_15568,N_19330);
or U23654 (N_23654,N_19394,N_16999);
and U23655 (N_23655,N_16453,N_16121);
or U23656 (N_23656,N_19656,N_17517);
and U23657 (N_23657,N_19574,N_16476);
nand U23658 (N_23658,N_15713,N_17103);
or U23659 (N_23659,N_18536,N_18035);
nand U23660 (N_23660,N_17322,N_15057);
xnor U23661 (N_23661,N_16250,N_18715);
nand U23662 (N_23662,N_18741,N_16397);
nand U23663 (N_23663,N_17807,N_18768);
or U23664 (N_23664,N_15176,N_19917);
and U23665 (N_23665,N_16888,N_18227);
and U23666 (N_23666,N_17142,N_19816);
nand U23667 (N_23667,N_15768,N_19891);
nand U23668 (N_23668,N_15539,N_17963);
and U23669 (N_23669,N_17497,N_15766);
and U23670 (N_23670,N_17131,N_16708);
or U23671 (N_23671,N_15745,N_15843);
or U23672 (N_23672,N_18838,N_16891);
or U23673 (N_23673,N_17372,N_17297);
nand U23674 (N_23674,N_15131,N_17526);
nand U23675 (N_23675,N_19659,N_18040);
and U23676 (N_23676,N_18294,N_15448);
nor U23677 (N_23677,N_18624,N_15332);
and U23678 (N_23678,N_18838,N_18073);
or U23679 (N_23679,N_17193,N_19338);
xor U23680 (N_23680,N_18522,N_19488);
nand U23681 (N_23681,N_15231,N_16014);
or U23682 (N_23682,N_17376,N_16332);
nand U23683 (N_23683,N_15127,N_18428);
or U23684 (N_23684,N_19104,N_17140);
xor U23685 (N_23685,N_19556,N_18487);
xor U23686 (N_23686,N_15538,N_17700);
nor U23687 (N_23687,N_19910,N_18956);
and U23688 (N_23688,N_19793,N_18067);
and U23689 (N_23689,N_18073,N_19469);
or U23690 (N_23690,N_17441,N_15088);
nor U23691 (N_23691,N_17919,N_17393);
and U23692 (N_23692,N_15543,N_15891);
or U23693 (N_23693,N_17628,N_17062);
or U23694 (N_23694,N_18403,N_17166);
xnor U23695 (N_23695,N_15673,N_16961);
nand U23696 (N_23696,N_18372,N_16201);
and U23697 (N_23697,N_17376,N_17739);
xor U23698 (N_23698,N_15015,N_15938);
and U23699 (N_23699,N_18565,N_19499);
xnor U23700 (N_23700,N_15967,N_15342);
xnor U23701 (N_23701,N_17276,N_16116);
nand U23702 (N_23702,N_19707,N_19131);
nor U23703 (N_23703,N_18541,N_16422);
nor U23704 (N_23704,N_15355,N_17409);
nor U23705 (N_23705,N_16198,N_19058);
nand U23706 (N_23706,N_18745,N_16303);
xnor U23707 (N_23707,N_19237,N_17134);
and U23708 (N_23708,N_19904,N_15816);
or U23709 (N_23709,N_16679,N_18978);
nor U23710 (N_23710,N_19087,N_17023);
or U23711 (N_23711,N_16649,N_16141);
nor U23712 (N_23712,N_17298,N_18287);
or U23713 (N_23713,N_18466,N_15134);
nor U23714 (N_23714,N_17924,N_19077);
nor U23715 (N_23715,N_16936,N_15631);
nand U23716 (N_23716,N_16263,N_16885);
or U23717 (N_23717,N_16788,N_17939);
nor U23718 (N_23718,N_17358,N_17649);
or U23719 (N_23719,N_18218,N_17274);
nand U23720 (N_23720,N_17091,N_16138);
nor U23721 (N_23721,N_18947,N_18093);
xor U23722 (N_23722,N_18851,N_19929);
xor U23723 (N_23723,N_17219,N_15176);
and U23724 (N_23724,N_17374,N_15142);
xnor U23725 (N_23725,N_16226,N_16358);
and U23726 (N_23726,N_18353,N_17439);
or U23727 (N_23727,N_15352,N_19439);
xnor U23728 (N_23728,N_19788,N_16798);
or U23729 (N_23729,N_15550,N_19803);
or U23730 (N_23730,N_18278,N_17611);
nand U23731 (N_23731,N_18241,N_19233);
and U23732 (N_23732,N_17249,N_15068);
or U23733 (N_23733,N_18261,N_19467);
xnor U23734 (N_23734,N_18481,N_18852);
or U23735 (N_23735,N_17960,N_19009);
nor U23736 (N_23736,N_17606,N_16759);
xnor U23737 (N_23737,N_17121,N_18600);
and U23738 (N_23738,N_19744,N_15330);
nor U23739 (N_23739,N_19745,N_15532);
xnor U23740 (N_23740,N_16225,N_16387);
nor U23741 (N_23741,N_18310,N_18803);
xnor U23742 (N_23742,N_19283,N_15009);
nor U23743 (N_23743,N_16545,N_16008);
and U23744 (N_23744,N_15175,N_18641);
xor U23745 (N_23745,N_17502,N_16756);
and U23746 (N_23746,N_19428,N_19823);
nand U23747 (N_23747,N_16451,N_18139);
nand U23748 (N_23748,N_15555,N_18259);
xor U23749 (N_23749,N_17081,N_16405);
xnor U23750 (N_23750,N_18368,N_18235);
and U23751 (N_23751,N_18690,N_16711);
and U23752 (N_23752,N_15382,N_15627);
xnor U23753 (N_23753,N_17381,N_19005);
and U23754 (N_23754,N_18941,N_18184);
or U23755 (N_23755,N_18503,N_16979);
or U23756 (N_23756,N_15212,N_18676);
nand U23757 (N_23757,N_15107,N_19493);
or U23758 (N_23758,N_18468,N_16725);
nand U23759 (N_23759,N_19676,N_18910);
nand U23760 (N_23760,N_15655,N_16610);
nor U23761 (N_23761,N_17431,N_15729);
or U23762 (N_23762,N_19833,N_19346);
or U23763 (N_23763,N_19229,N_16176);
nand U23764 (N_23764,N_17666,N_19245);
xnor U23765 (N_23765,N_18899,N_18000);
nand U23766 (N_23766,N_16379,N_16310);
or U23767 (N_23767,N_18421,N_18591);
and U23768 (N_23768,N_18758,N_18321);
nand U23769 (N_23769,N_16124,N_18241);
or U23770 (N_23770,N_18649,N_17576);
nand U23771 (N_23771,N_17069,N_19420);
xor U23772 (N_23772,N_17961,N_19069);
xor U23773 (N_23773,N_16785,N_15629);
or U23774 (N_23774,N_17763,N_16867);
and U23775 (N_23775,N_16129,N_18874);
nor U23776 (N_23776,N_16303,N_15261);
or U23777 (N_23777,N_19255,N_15196);
nand U23778 (N_23778,N_19472,N_15720);
xnor U23779 (N_23779,N_17758,N_17906);
xnor U23780 (N_23780,N_15853,N_17707);
nor U23781 (N_23781,N_19107,N_17469);
nor U23782 (N_23782,N_16247,N_18302);
xor U23783 (N_23783,N_17215,N_17828);
nand U23784 (N_23784,N_18111,N_19518);
xnor U23785 (N_23785,N_17594,N_15554);
nand U23786 (N_23786,N_18020,N_15158);
or U23787 (N_23787,N_16853,N_19289);
or U23788 (N_23788,N_15672,N_18283);
xnor U23789 (N_23789,N_17161,N_16926);
xor U23790 (N_23790,N_16247,N_17717);
or U23791 (N_23791,N_17547,N_19187);
and U23792 (N_23792,N_16980,N_18337);
nand U23793 (N_23793,N_18931,N_19407);
and U23794 (N_23794,N_18384,N_17267);
and U23795 (N_23795,N_18989,N_16830);
or U23796 (N_23796,N_18679,N_18150);
and U23797 (N_23797,N_15328,N_18447);
or U23798 (N_23798,N_15378,N_18263);
and U23799 (N_23799,N_18828,N_15593);
and U23800 (N_23800,N_17977,N_19891);
nor U23801 (N_23801,N_17747,N_15382);
and U23802 (N_23802,N_18490,N_15473);
nand U23803 (N_23803,N_17554,N_17610);
or U23804 (N_23804,N_17071,N_16059);
nor U23805 (N_23805,N_19804,N_19382);
nand U23806 (N_23806,N_17223,N_15030);
or U23807 (N_23807,N_18205,N_18689);
and U23808 (N_23808,N_16374,N_17248);
nor U23809 (N_23809,N_18735,N_18856);
and U23810 (N_23810,N_18027,N_15048);
or U23811 (N_23811,N_16346,N_16029);
nor U23812 (N_23812,N_15575,N_16267);
xnor U23813 (N_23813,N_16898,N_15945);
xnor U23814 (N_23814,N_17979,N_19914);
or U23815 (N_23815,N_15275,N_19059);
and U23816 (N_23816,N_19960,N_18850);
or U23817 (N_23817,N_19929,N_16850);
xnor U23818 (N_23818,N_19144,N_18481);
xnor U23819 (N_23819,N_15861,N_19252);
and U23820 (N_23820,N_18916,N_17193);
or U23821 (N_23821,N_17492,N_16905);
xnor U23822 (N_23822,N_19660,N_15358);
or U23823 (N_23823,N_19851,N_17352);
and U23824 (N_23824,N_19790,N_18136);
nand U23825 (N_23825,N_18100,N_16234);
or U23826 (N_23826,N_16924,N_18098);
nand U23827 (N_23827,N_15401,N_18115);
nor U23828 (N_23828,N_16835,N_19927);
and U23829 (N_23829,N_16464,N_19453);
xnor U23830 (N_23830,N_17228,N_16891);
nor U23831 (N_23831,N_16621,N_15704);
xnor U23832 (N_23832,N_19951,N_19418);
nor U23833 (N_23833,N_15276,N_17610);
nor U23834 (N_23834,N_17149,N_18247);
or U23835 (N_23835,N_17047,N_16623);
xnor U23836 (N_23836,N_19189,N_19557);
or U23837 (N_23837,N_15951,N_16877);
and U23838 (N_23838,N_19009,N_18164);
nor U23839 (N_23839,N_15172,N_18225);
xor U23840 (N_23840,N_19919,N_18767);
nand U23841 (N_23841,N_16021,N_16311);
and U23842 (N_23842,N_15649,N_17136);
or U23843 (N_23843,N_19960,N_16823);
and U23844 (N_23844,N_16783,N_17977);
and U23845 (N_23845,N_18156,N_15904);
and U23846 (N_23846,N_15338,N_15870);
or U23847 (N_23847,N_19718,N_17537);
or U23848 (N_23848,N_17571,N_19300);
xnor U23849 (N_23849,N_16684,N_15346);
xor U23850 (N_23850,N_17344,N_17312);
nand U23851 (N_23851,N_15927,N_18059);
xor U23852 (N_23852,N_19151,N_19152);
nand U23853 (N_23853,N_15328,N_16342);
nor U23854 (N_23854,N_15564,N_18053);
or U23855 (N_23855,N_15837,N_18883);
nor U23856 (N_23856,N_19060,N_19628);
xor U23857 (N_23857,N_18823,N_17407);
and U23858 (N_23858,N_16355,N_17172);
nor U23859 (N_23859,N_15896,N_19128);
nor U23860 (N_23860,N_16877,N_18032);
and U23861 (N_23861,N_15738,N_19739);
xor U23862 (N_23862,N_16870,N_17113);
and U23863 (N_23863,N_16507,N_17756);
or U23864 (N_23864,N_17028,N_15934);
or U23865 (N_23865,N_16772,N_19151);
nand U23866 (N_23866,N_15264,N_19030);
and U23867 (N_23867,N_16072,N_15185);
nand U23868 (N_23868,N_15218,N_18304);
nand U23869 (N_23869,N_16697,N_18830);
xnor U23870 (N_23870,N_17137,N_15652);
xor U23871 (N_23871,N_17163,N_16261);
and U23872 (N_23872,N_18296,N_18412);
and U23873 (N_23873,N_18079,N_19365);
nand U23874 (N_23874,N_17213,N_17301);
and U23875 (N_23875,N_16012,N_15121);
xnor U23876 (N_23876,N_15140,N_17309);
nor U23877 (N_23877,N_19428,N_16610);
or U23878 (N_23878,N_15808,N_18380);
xnor U23879 (N_23879,N_19075,N_18466);
nand U23880 (N_23880,N_17018,N_16468);
nand U23881 (N_23881,N_17502,N_19998);
and U23882 (N_23882,N_19113,N_16575);
nor U23883 (N_23883,N_19133,N_19725);
nor U23884 (N_23884,N_18292,N_15860);
nand U23885 (N_23885,N_16201,N_15190);
nor U23886 (N_23886,N_16616,N_16165);
nand U23887 (N_23887,N_16609,N_18462);
nand U23888 (N_23888,N_16974,N_16882);
nor U23889 (N_23889,N_15966,N_16116);
or U23890 (N_23890,N_19425,N_16245);
xnor U23891 (N_23891,N_15898,N_15769);
or U23892 (N_23892,N_15035,N_18876);
nor U23893 (N_23893,N_19471,N_17801);
or U23894 (N_23894,N_16623,N_17173);
xor U23895 (N_23895,N_17130,N_15219);
or U23896 (N_23896,N_15154,N_16024);
nor U23897 (N_23897,N_17489,N_16425);
or U23898 (N_23898,N_15755,N_18190);
or U23899 (N_23899,N_18523,N_16902);
or U23900 (N_23900,N_18221,N_19834);
nand U23901 (N_23901,N_15741,N_19734);
nand U23902 (N_23902,N_19277,N_18581);
nor U23903 (N_23903,N_17379,N_15408);
nor U23904 (N_23904,N_17472,N_19578);
and U23905 (N_23905,N_19692,N_17957);
nor U23906 (N_23906,N_15830,N_17185);
xor U23907 (N_23907,N_19152,N_18801);
nand U23908 (N_23908,N_18452,N_18529);
xor U23909 (N_23909,N_19198,N_18844);
and U23910 (N_23910,N_16893,N_18587);
xor U23911 (N_23911,N_16334,N_15269);
nor U23912 (N_23912,N_19445,N_16821);
or U23913 (N_23913,N_19858,N_15849);
or U23914 (N_23914,N_19498,N_17183);
and U23915 (N_23915,N_15201,N_19831);
nand U23916 (N_23916,N_15886,N_18743);
xnor U23917 (N_23917,N_18614,N_19150);
and U23918 (N_23918,N_18234,N_15898);
and U23919 (N_23919,N_19951,N_19440);
or U23920 (N_23920,N_17501,N_16270);
and U23921 (N_23921,N_18438,N_16209);
nand U23922 (N_23922,N_16197,N_19511);
nand U23923 (N_23923,N_18563,N_16563);
or U23924 (N_23924,N_16027,N_16988);
or U23925 (N_23925,N_17083,N_16709);
nand U23926 (N_23926,N_18779,N_16551);
xor U23927 (N_23927,N_19003,N_18118);
and U23928 (N_23928,N_17391,N_16576);
xor U23929 (N_23929,N_16651,N_18235);
nor U23930 (N_23930,N_17492,N_19564);
nor U23931 (N_23931,N_17878,N_17327);
nor U23932 (N_23932,N_19826,N_19582);
or U23933 (N_23933,N_19865,N_16967);
nand U23934 (N_23934,N_17293,N_19547);
or U23935 (N_23935,N_19760,N_19746);
xor U23936 (N_23936,N_18006,N_19279);
or U23937 (N_23937,N_18585,N_18040);
or U23938 (N_23938,N_19061,N_17027);
nand U23939 (N_23939,N_15004,N_17026);
and U23940 (N_23940,N_19127,N_17684);
or U23941 (N_23941,N_18921,N_17586);
xor U23942 (N_23942,N_19659,N_16294);
and U23943 (N_23943,N_16098,N_18280);
and U23944 (N_23944,N_19797,N_18134);
nor U23945 (N_23945,N_15906,N_16014);
nor U23946 (N_23946,N_17230,N_17237);
nand U23947 (N_23947,N_19550,N_18186);
or U23948 (N_23948,N_18671,N_19119);
or U23949 (N_23949,N_17464,N_17804);
xnor U23950 (N_23950,N_17331,N_18798);
or U23951 (N_23951,N_15059,N_18503);
nand U23952 (N_23952,N_18418,N_16443);
nor U23953 (N_23953,N_16445,N_15599);
nand U23954 (N_23954,N_18874,N_19750);
nor U23955 (N_23955,N_16037,N_16920);
xnor U23956 (N_23956,N_15879,N_18529);
and U23957 (N_23957,N_17793,N_16404);
nand U23958 (N_23958,N_18164,N_18242);
or U23959 (N_23959,N_15544,N_18282);
or U23960 (N_23960,N_15899,N_19743);
nor U23961 (N_23961,N_18960,N_16397);
xnor U23962 (N_23962,N_19029,N_17191);
or U23963 (N_23963,N_19013,N_16917);
xor U23964 (N_23964,N_18394,N_16427);
or U23965 (N_23965,N_18442,N_16988);
nand U23966 (N_23966,N_16618,N_17083);
and U23967 (N_23967,N_17491,N_15962);
or U23968 (N_23968,N_17546,N_18377);
nand U23969 (N_23969,N_16206,N_19785);
xnor U23970 (N_23970,N_18885,N_18069);
nand U23971 (N_23971,N_18822,N_15217);
nor U23972 (N_23972,N_18658,N_17621);
nand U23973 (N_23973,N_19954,N_16520);
nor U23974 (N_23974,N_18751,N_15462);
or U23975 (N_23975,N_18642,N_17275);
nor U23976 (N_23976,N_19066,N_17286);
nand U23977 (N_23977,N_17326,N_16217);
xnor U23978 (N_23978,N_15874,N_16999);
or U23979 (N_23979,N_19293,N_19908);
nor U23980 (N_23980,N_19303,N_19289);
or U23981 (N_23981,N_15994,N_19017);
nand U23982 (N_23982,N_19038,N_19546);
or U23983 (N_23983,N_16291,N_18035);
nand U23984 (N_23984,N_17931,N_19874);
and U23985 (N_23985,N_15252,N_15641);
or U23986 (N_23986,N_15903,N_17293);
nor U23987 (N_23987,N_17412,N_16946);
xnor U23988 (N_23988,N_17039,N_17736);
xor U23989 (N_23989,N_17343,N_17671);
xor U23990 (N_23990,N_18012,N_19331);
xnor U23991 (N_23991,N_16201,N_17794);
xnor U23992 (N_23992,N_15089,N_18712);
nor U23993 (N_23993,N_16297,N_18767);
nand U23994 (N_23994,N_15926,N_18407);
and U23995 (N_23995,N_18232,N_17303);
xor U23996 (N_23996,N_16826,N_15697);
xnor U23997 (N_23997,N_16344,N_16157);
nor U23998 (N_23998,N_16797,N_15139);
or U23999 (N_23999,N_17962,N_15191);
nor U24000 (N_24000,N_17698,N_19810);
nor U24001 (N_24001,N_16819,N_15304);
or U24002 (N_24002,N_17535,N_16090);
or U24003 (N_24003,N_18537,N_19950);
xor U24004 (N_24004,N_18841,N_19532);
nand U24005 (N_24005,N_19205,N_18605);
xor U24006 (N_24006,N_15731,N_15950);
and U24007 (N_24007,N_16321,N_18426);
and U24008 (N_24008,N_15063,N_15371);
xor U24009 (N_24009,N_18289,N_19249);
and U24010 (N_24010,N_16209,N_18885);
xnor U24011 (N_24011,N_19129,N_16896);
and U24012 (N_24012,N_18573,N_17807);
nand U24013 (N_24013,N_16388,N_17377);
nor U24014 (N_24014,N_17298,N_17392);
nor U24015 (N_24015,N_15943,N_19280);
and U24016 (N_24016,N_19684,N_17808);
xnor U24017 (N_24017,N_17868,N_18628);
or U24018 (N_24018,N_18896,N_18190);
nand U24019 (N_24019,N_19907,N_15434);
and U24020 (N_24020,N_19429,N_19939);
nand U24021 (N_24021,N_19024,N_18904);
and U24022 (N_24022,N_17138,N_17090);
nand U24023 (N_24023,N_18277,N_17071);
xor U24024 (N_24024,N_18357,N_17712);
and U24025 (N_24025,N_18841,N_18446);
xor U24026 (N_24026,N_17245,N_15408);
nand U24027 (N_24027,N_17613,N_15908);
xnor U24028 (N_24028,N_19559,N_18092);
xnor U24029 (N_24029,N_16821,N_16541);
or U24030 (N_24030,N_15803,N_17792);
and U24031 (N_24031,N_16838,N_17011);
nor U24032 (N_24032,N_19859,N_16221);
xor U24033 (N_24033,N_15276,N_17739);
and U24034 (N_24034,N_19973,N_15784);
nand U24035 (N_24035,N_19563,N_15480);
nor U24036 (N_24036,N_18466,N_16360);
xnor U24037 (N_24037,N_16334,N_15400);
nand U24038 (N_24038,N_16486,N_19897);
nor U24039 (N_24039,N_17914,N_16673);
nand U24040 (N_24040,N_18449,N_15408);
and U24041 (N_24041,N_15253,N_17214);
nand U24042 (N_24042,N_16425,N_15607);
nand U24043 (N_24043,N_19288,N_16477);
or U24044 (N_24044,N_17675,N_15456);
nor U24045 (N_24045,N_16598,N_18145);
or U24046 (N_24046,N_17580,N_17755);
and U24047 (N_24047,N_17710,N_19303);
and U24048 (N_24048,N_15631,N_19063);
nand U24049 (N_24049,N_15559,N_15945);
and U24050 (N_24050,N_17300,N_15144);
xor U24051 (N_24051,N_16811,N_18960);
and U24052 (N_24052,N_18478,N_18324);
or U24053 (N_24053,N_18303,N_17025);
or U24054 (N_24054,N_19228,N_17071);
nor U24055 (N_24055,N_17176,N_15096);
nand U24056 (N_24056,N_16597,N_19044);
nor U24057 (N_24057,N_16036,N_17111);
nand U24058 (N_24058,N_19161,N_15591);
or U24059 (N_24059,N_19533,N_18890);
xnor U24060 (N_24060,N_19045,N_17420);
or U24061 (N_24061,N_16746,N_19917);
nand U24062 (N_24062,N_19743,N_19492);
xor U24063 (N_24063,N_19065,N_18464);
xnor U24064 (N_24064,N_19255,N_18348);
xnor U24065 (N_24065,N_16393,N_19381);
xor U24066 (N_24066,N_15616,N_18746);
and U24067 (N_24067,N_18842,N_18935);
xor U24068 (N_24068,N_18651,N_18982);
or U24069 (N_24069,N_17242,N_17596);
nor U24070 (N_24070,N_18136,N_15848);
nand U24071 (N_24071,N_15437,N_15055);
or U24072 (N_24072,N_15964,N_17945);
xor U24073 (N_24073,N_16927,N_19162);
nand U24074 (N_24074,N_15929,N_15801);
xnor U24075 (N_24075,N_19047,N_16563);
nand U24076 (N_24076,N_18287,N_18375);
or U24077 (N_24077,N_16677,N_16345);
xnor U24078 (N_24078,N_19727,N_17416);
or U24079 (N_24079,N_16852,N_16131);
xor U24080 (N_24080,N_19002,N_17224);
nand U24081 (N_24081,N_17904,N_18491);
xnor U24082 (N_24082,N_15180,N_17876);
xor U24083 (N_24083,N_16736,N_16586);
or U24084 (N_24084,N_16507,N_19161);
and U24085 (N_24085,N_15945,N_19936);
xor U24086 (N_24086,N_17823,N_18145);
and U24087 (N_24087,N_17106,N_19671);
nand U24088 (N_24088,N_17329,N_17135);
and U24089 (N_24089,N_17400,N_17856);
or U24090 (N_24090,N_15044,N_16140);
or U24091 (N_24091,N_15514,N_16427);
or U24092 (N_24092,N_18305,N_17603);
xor U24093 (N_24093,N_19982,N_18655);
nand U24094 (N_24094,N_15695,N_19939);
nand U24095 (N_24095,N_18120,N_17622);
nand U24096 (N_24096,N_15672,N_19421);
or U24097 (N_24097,N_19694,N_18645);
and U24098 (N_24098,N_18356,N_18789);
nor U24099 (N_24099,N_18443,N_18780);
nor U24100 (N_24100,N_15581,N_16139);
and U24101 (N_24101,N_15341,N_16225);
nand U24102 (N_24102,N_18416,N_18785);
or U24103 (N_24103,N_19041,N_18058);
and U24104 (N_24104,N_18925,N_16700);
xnor U24105 (N_24105,N_15446,N_18408);
nor U24106 (N_24106,N_17395,N_16539);
nor U24107 (N_24107,N_17597,N_17209);
and U24108 (N_24108,N_16861,N_17548);
xnor U24109 (N_24109,N_19721,N_17710);
xnor U24110 (N_24110,N_18952,N_15985);
and U24111 (N_24111,N_16932,N_17768);
nand U24112 (N_24112,N_19981,N_15472);
nor U24113 (N_24113,N_18905,N_19399);
or U24114 (N_24114,N_18452,N_19147);
nand U24115 (N_24115,N_18469,N_15579);
or U24116 (N_24116,N_16485,N_15560);
and U24117 (N_24117,N_16093,N_17303);
nand U24118 (N_24118,N_15492,N_15063);
nor U24119 (N_24119,N_15116,N_15494);
nor U24120 (N_24120,N_17405,N_15476);
or U24121 (N_24121,N_19592,N_17492);
nor U24122 (N_24122,N_18431,N_16479);
nor U24123 (N_24123,N_15741,N_19146);
or U24124 (N_24124,N_16252,N_16888);
or U24125 (N_24125,N_18509,N_15249);
or U24126 (N_24126,N_15771,N_16934);
nor U24127 (N_24127,N_16237,N_16403);
nand U24128 (N_24128,N_16130,N_17796);
or U24129 (N_24129,N_18039,N_18230);
and U24130 (N_24130,N_17261,N_16915);
or U24131 (N_24131,N_16416,N_18323);
and U24132 (N_24132,N_17574,N_18114);
xor U24133 (N_24133,N_19988,N_15574);
or U24134 (N_24134,N_17735,N_18991);
nor U24135 (N_24135,N_17501,N_19733);
or U24136 (N_24136,N_16643,N_16791);
nand U24137 (N_24137,N_15081,N_15825);
nor U24138 (N_24138,N_15480,N_15124);
nor U24139 (N_24139,N_15881,N_15035);
nor U24140 (N_24140,N_19028,N_17133);
and U24141 (N_24141,N_18262,N_17020);
and U24142 (N_24142,N_18313,N_17791);
nor U24143 (N_24143,N_19334,N_17775);
and U24144 (N_24144,N_15596,N_19102);
and U24145 (N_24145,N_18334,N_15070);
nand U24146 (N_24146,N_19849,N_17765);
xor U24147 (N_24147,N_15207,N_15655);
or U24148 (N_24148,N_19763,N_15160);
or U24149 (N_24149,N_19324,N_17690);
or U24150 (N_24150,N_18190,N_15389);
nor U24151 (N_24151,N_16526,N_17558);
and U24152 (N_24152,N_19814,N_17817);
nor U24153 (N_24153,N_17050,N_16584);
or U24154 (N_24154,N_16157,N_16531);
xnor U24155 (N_24155,N_18800,N_19276);
nand U24156 (N_24156,N_18832,N_15589);
nand U24157 (N_24157,N_17022,N_16213);
and U24158 (N_24158,N_19214,N_19065);
or U24159 (N_24159,N_15464,N_19851);
nand U24160 (N_24160,N_15154,N_16917);
xor U24161 (N_24161,N_17217,N_16446);
xnor U24162 (N_24162,N_18607,N_15382);
xnor U24163 (N_24163,N_16606,N_18032);
nor U24164 (N_24164,N_17352,N_18315);
and U24165 (N_24165,N_19811,N_15791);
nand U24166 (N_24166,N_17174,N_19811);
xnor U24167 (N_24167,N_17983,N_19094);
and U24168 (N_24168,N_16324,N_15812);
xnor U24169 (N_24169,N_17754,N_17063);
nor U24170 (N_24170,N_18485,N_19165);
xnor U24171 (N_24171,N_19861,N_19117);
or U24172 (N_24172,N_17124,N_17872);
and U24173 (N_24173,N_18830,N_17641);
or U24174 (N_24174,N_15642,N_17644);
nand U24175 (N_24175,N_16729,N_19562);
nor U24176 (N_24176,N_17409,N_16752);
and U24177 (N_24177,N_18649,N_17510);
nand U24178 (N_24178,N_18092,N_19918);
nor U24179 (N_24179,N_15978,N_17054);
nand U24180 (N_24180,N_18650,N_18898);
and U24181 (N_24181,N_18445,N_16155);
and U24182 (N_24182,N_16316,N_16081);
nor U24183 (N_24183,N_16747,N_19560);
or U24184 (N_24184,N_15227,N_16766);
nand U24185 (N_24185,N_15364,N_17093);
xor U24186 (N_24186,N_18345,N_18869);
nor U24187 (N_24187,N_16962,N_17079);
and U24188 (N_24188,N_18395,N_17783);
and U24189 (N_24189,N_18041,N_18419);
nor U24190 (N_24190,N_18583,N_18299);
nor U24191 (N_24191,N_18029,N_18657);
nand U24192 (N_24192,N_17711,N_17045);
nand U24193 (N_24193,N_19590,N_17123);
nand U24194 (N_24194,N_19972,N_16463);
nor U24195 (N_24195,N_18632,N_17906);
nor U24196 (N_24196,N_15741,N_15376);
or U24197 (N_24197,N_16502,N_15714);
or U24198 (N_24198,N_15166,N_15071);
and U24199 (N_24199,N_16406,N_18792);
nand U24200 (N_24200,N_18689,N_15273);
nand U24201 (N_24201,N_18046,N_19309);
nor U24202 (N_24202,N_16155,N_15191);
or U24203 (N_24203,N_15339,N_19395);
nor U24204 (N_24204,N_18830,N_18070);
nand U24205 (N_24205,N_16817,N_18065);
xor U24206 (N_24206,N_19399,N_19953);
or U24207 (N_24207,N_19818,N_15771);
xnor U24208 (N_24208,N_19354,N_15025);
and U24209 (N_24209,N_19005,N_16113);
nand U24210 (N_24210,N_19830,N_16437);
xor U24211 (N_24211,N_15563,N_15402);
or U24212 (N_24212,N_15326,N_15975);
or U24213 (N_24213,N_18201,N_17887);
xnor U24214 (N_24214,N_18893,N_19084);
or U24215 (N_24215,N_17893,N_19803);
nand U24216 (N_24216,N_19170,N_15855);
or U24217 (N_24217,N_17765,N_19558);
xnor U24218 (N_24218,N_19578,N_18428);
nor U24219 (N_24219,N_16611,N_16559);
nand U24220 (N_24220,N_18827,N_17389);
xor U24221 (N_24221,N_17899,N_16159);
xnor U24222 (N_24222,N_19663,N_18217);
nand U24223 (N_24223,N_16804,N_17009);
and U24224 (N_24224,N_16703,N_15876);
nor U24225 (N_24225,N_19899,N_15759);
nor U24226 (N_24226,N_18925,N_15641);
xor U24227 (N_24227,N_18381,N_19447);
and U24228 (N_24228,N_15740,N_16710);
and U24229 (N_24229,N_15013,N_19794);
or U24230 (N_24230,N_18562,N_16064);
nand U24231 (N_24231,N_18207,N_15179);
nor U24232 (N_24232,N_18179,N_15425);
nand U24233 (N_24233,N_16831,N_16945);
xnor U24234 (N_24234,N_18622,N_18127);
nand U24235 (N_24235,N_17229,N_16879);
nor U24236 (N_24236,N_16472,N_18686);
and U24237 (N_24237,N_16674,N_17741);
and U24238 (N_24238,N_18239,N_15357);
nor U24239 (N_24239,N_17257,N_15739);
xor U24240 (N_24240,N_15530,N_15497);
and U24241 (N_24241,N_17152,N_17264);
nand U24242 (N_24242,N_15698,N_19462);
nand U24243 (N_24243,N_15193,N_15474);
nor U24244 (N_24244,N_16239,N_18491);
nor U24245 (N_24245,N_19524,N_16911);
xnor U24246 (N_24246,N_18834,N_19249);
nand U24247 (N_24247,N_19414,N_19021);
or U24248 (N_24248,N_19000,N_19586);
and U24249 (N_24249,N_18534,N_19605);
xnor U24250 (N_24250,N_19534,N_19282);
xnor U24251 (N_24251,N_19373,N_15777);
or U24252 (N_24252,N_17685,N_15111);
and U24253 (N_24253,N_15075,N_18440);
nor U24254 (N_24254,N_19159,N_18948);
nor U24255 (N_24255,N_15037,N_19068);
or U24256 (N_24256,N_17734,N_19456);
xnor U24257 (N_24257,N_16024,N_19495);
nor U24258 (N_24258,N_15238,N_16094);
nor U24259 (N_24259,N_15479,N_19582);
and U24260 (N_24260,N_19188,N_16569);
nor U24261 (N_24261,N_17742,N_16221);
nand U24262 (N_24262,N_18729,N_19762);
nand U24263 (N_24263,N_19289,N_17891);
and U24264 (N_24264,N_15979,N_19319);
nand U24265 (N_24265,N_16501,N_16253);
xnor U24266 (N_24266,N_18508,N_18210);
or U24267 (N_24267,N_17471,N_17040);
or U24268 (N_24268,N_15175,N_19843);
xnor U24269 (N_24269,N_17272,N_19687);
nand U24270 (N_24270,N_16439,N_19677);
nor U24271 (N_24271,N_18153,N_15865);
or U24272 (N_24272,N_18764,N_19600);
xor U24273 (N_24273,N_16514,N_16502);
or U24274 (N_24274,N_16692,N_18359);
nor U24275 (N_24275,N_19786,N_19314);
and U24276 (N_24276,N_19054,N_18449);
and U24277 (N_24277,N_16143,N_15625);
nand U24278 (N_24278,N_15679,N_16843);
or U24279 (N_24279,N_17428,N_15790);
xnor U24280 (N_24280,N_19635,N_15405);
or U24281 (N_24281,N_16097,N_15718);
xnor U24282 (N_24282,N_17341,N_15547);
and U24283 (N_24283,N_15758,N_17702);
nor U24284 (N_24284,N_15010,N_15535);
xor U24285 (N_24285,N_18775,N_18275);
nand U24286 (N_24286,N_17525,N_18604);
or U24287 (N_24287,N_15688,N_15354);
nor U24288 (N_24288,N_15144,N_19020);
xnor U24289 (N_24289,N_18741,N_15348);
nor U24290 (N_24290,N_19016,N_17687);
nand U24291 (N_24291,N_15050,N_15365);
nand U24292 (N_24292,N_15384,N_18865);
nor U24293 (N_24293,N_19881,N_15436);
xor U24294 (N_24294,N_18572,N_15272);
xor U24295 (N_24295,N_18815,N_18034);
and U24296 (N_24296,N_18485,N_18474);
and U24297 (N_24297,N_15998,N_17192);
xnor U24298 (N_24298,N_16613,N_17376);
or U24299 (N_24299,N_18189,N_16008);
and U24300 (N_24300,N_17897,N_15864);
xnor U24301 (N_24301,N_17735,N_18353);
nor U24302 (N_24302,N_15926,N_16577);
and U24303 (N_24303,N_16674,N_16104);
and U24304 (N_24304,N_19764,N_16417);
or U24305 (N_24305,N_18105,N_15169);
nand U24306 (N_24306,N_16157,N_18718);
or U24307 (N_24307,N_16858,N_19640);
and U24308 (N_24308,N_17084,N_15851);
or U24309 (N_24309,N_16374,N_16140);
nor U24310 (N_24310,N_15792,N_18189);
xnor U24311 (N_24311,N_17848,N_18429);
xnor U24312 (N_24312,N_19259,N_19551);
nor U24313 (N_24313,N_15771,N_16684);
xnor U24314 (N_24314,N_15485,N_19784);
or U24315 (N_24315,N_15470,N_17572);
nand U24316 (N_24316,N_16851,N_15293);
nor U24317 (N_24317,N_18170,N_18023);
nand U24318 (N_24318,N_16117,N_19032);
nand U24319 (N_24319,N_16051,N_19064);
nor U24320 (N_24320,N_16777,N_19880);
nand U24321 (N_24321,N_15870,N_18406);
nand U24322 (N_24322,N_18355,N_15649);
and U24323 (N_24323,N_16796,N_18945);
xor U24324 (N_24324,N_18972,N_19399);
xor U24325 (N_24325,N_16439,N_17450);
nor U24326 (N_24326,N_16681,N_18963);
or U24327 (N_24327,N_17393,N_16791);
nor U24328 (N_24328,N_17406,N_19211);
and U24329 (N_24329,N_16767,N_18287);
and U24330 (N_24330,N_15461,N_15421);
and U24331 (N_24331,N_16388,N_15763);
or U24332 (N_24332,N_18085,N_17750);
xnor U24333 (N_24333,N_18312,N_17505);
or U24334 (N_24334,N_19738,N_19447);
nand U24335 (N_24335,N_16143,N_19121);
and U24336 (N_24336,N_18397,N_17188);
nand U24337 (N_24337,N_17480,N_18804);
xor U24338 (N_24338,N_16733,N_16720);
and U24339 (N_24339,N_16703,N_16133);
or U24340 (N_24340,N_16170,N_16088);
nor U24341 (N_24341,N_15271,N_17206);
or U24342 (N_24342,N_19633,N_16017);
nor U24343 (N_24343,N_17487,N_19241);
or U24344 (N_24344,N_17194,N_19413);
nor U24345 (N_24345,N_18765,N_18156);
nor U24346 (N_24346,N_15218,N_15873);
nor U24347 (N_24347,N_19659,N_17185);
and U24348 (N_24348,N_16812,N_19764);
xor U24349 (N_24349,N_15009,N_17735);
and U24350 (N_24350,N_17931,N_18830);
xor U24351 (N_24351,N_19088,N_19358);
and U24352 (N_24352,N_19374,N_15414);
nand U24353 (N_24353,N_17185,N_19066);
and U24354 (N_24354,N_17603,N_19088);
nand U24355 (N_24355,N_17215,N_18548);
nor U24356 (N_24356,N_19021,N_17826);
or U24357 (N_24357,N_19984,N_15425);
nand U24358 (N_24358,N_16495,N_18348);
nand U24359 (N_24359,N_19806,N_18622);
and U24360 (N_24360,N_19802,N_17165);
nor U24361 (N_24361,N_19567,N_16731);
nand U24362 (N_24362,N_19824,N_19423);
nand U24363 (N_24363,N_15182,N_15447);
or U24364 (N_24364,N_18580,N_15109);
or U24365 (N_24365,N_17604,N_15078);
or U24366 (N_24366,N_18014,N_17775);
nor U24367 (N_24367,N_19332,N_16545);
or U24368 (N_24368,N_19883,N_18287);
xor U24369 (N_24369,N_18483,N_16879);
xor U24370 (N_24370,N_19269,N_15686);
nand U24371 (N_24371,N_16856,N_16783);
nand U24372 (N_24372,N_17729,N_16088);
or U24373 (N_24373,N_17560,N_18914);
xor U24374 (N_24374,N_17985,N_15670);
and U24375 (N_24375,N_19374,N_15320);
and U24376 (N_24376,N_19965,N_17507);
and U24377 (N_24377,N_16187,N_16008);
xnor U24378 (N_24378,N_16796,N_16529);
xnor U24379 (N_24379,N_16805,N_15595);
or U24380 (N_24380,N_16232,N_18651);
nand U24381 (N_24381,N_18988,N_16433);
nand U24382 (N_24382,N_15634,N_18955);
nor U24383 (N_24383,N_15432,N_18134);
and U24384 (N_24384,N_19845,N_17002);
xnor U24385 (N_24385,N_17368,N_17740);
or U24386 (N_24386,N_19334,N_18813);
or U24387 (N_24387,N_19397,N_19527);
nor U24388 (N_24388,N_17814,N_15560);
or U24389 (N_24389,N_15867,N_18005);
and U24390 (N_24390,N_15506,N_16440);
and U24391 (N_24391,N_18003,N_15774);
nand U24392 (N_24392,N_17496,N_17918);
and U24393 (N_24393,N_16909,N_19837);
nor U24394 (N_24394,N_18764,N_17587);
and U24395 (N_24395,N_19245,N_15669);
nand U24396 (N_24396,N_17282,N_19044);
nor U24397 (N_24397,N_18313,N_19092);
nor U24398 (N_24398,N_18228,N_17939);
nor U24399 (N_24399,N_18225,N_15137);
xor U24400 (N_24400,N_19569,N_15948);
or U24401 (N_24401,N_15292,N_16776);
nor U24402 (N_24402,N_16385,N_19223);
and U24403 (N_24403,N_19806,N_17772);
or U24404 (N_24404,N_17239,N_18630);
nor U24405 (N_24405,N_16309,N_18916);
nand U24406 (N_24406,N_15683,N_16769);
nand U24407 (N_24407,N_17572,N_16019);
xor U24408 (N_24408,N_15951,N_17639);
or U24409 (N_24409,N_15949,N_16670);
nand U24410 (N_24410,N_19107,N_18739);
and U24411 (N_24411,N_16549,N_19271);
or U24412 (N_24412,N_18616,N_17360);
nor U24413 (N_24413,N_16171,N_18904);
or U24414 (N_24414,N_16445,N_17302);
xor U24415 (N_24415,N_15467,N_19578);
or U24416 (N_24416,N_16590,N_16597);
nand U24417 (N_24417,N_19477,N_17082);
xnor U24418 (N_24418,N_18619,N_15222);
nand U24419 (N_24419,N_16336,N_18985);
xnor U24420 (N_24420,N_15735,N_16902);
nor U24421 (N_24421,N_19904,N_18923);
nand U24422 (N_24422,N_16850,N_15310);
nand U24423 (N_24423,N_17058,N_17585);
nand U24424 (N_24424,N_18761,N_15361);
or U24425 (N_24425,N_17858,N_18161);
xor U24426 (N_24426,N_16236,N_16502);
or U24427 (N_24427,N_17860,N_19709);
or U24428 (N_24428,N_19668,N_19447);
or U24429 (N_24429,N_19962,N_16824);
xor U24430 (N_24430,N_16694,N_16550);
nor U24431 (N_24431,N_15717,N_15773);
nand U24432 (N_24432,N_16139,N_18154);
nor U24433 (N_24433,N_18722,N_18782);
and U24434 (N_24434,N_18853,N_18761);
nand U24435 (N_24435,N_19213,N_18823);
or U24436 (N_24436,N_17324,N_16411);
and U24437 (N_24437,N_19819,N_16928);
nand U24438 (N_24438,N_19589,N_16517);
xnor U24439 (N_24439,N_19334,N_19621);
nand U24440 (N_24440,N_18748,N_16251);
xnor U24441 (N_24441,N_15463,N_15131);
nand U24442 (N_24442,N_16094,N_18838);
and U24443 (N_24443,N_16081,N_19639);
nor U24444 (N_24444,N_15847,N_18409);
nor U24445 (N_24445,N_15387,N_16687);
and U24446 (N_24446,N_15691,N_17817);
or U24447 (N_24447,N_15478,N_17343);
or U24448 (N_24448,N_17582,N_17284);
nor U24449 (N_24449,N_16925,N_16420);
nand U24450 (N_24450,N_17293,N_16620);
nand U24451 (N_24451,N_18292,N_19694);
and U24452 (N_24452,N_18123,N_18577);
and U24453 (N_24453,N_19334,N_16362);
or U24454 (N_24454,N_17643,N_16155);
xor U24455 (N_24455,N_16405,N_15075);
and U24456 (N_24456,N_18871,N_15613);
nand U24457 (N_24457,N_18281,N_16832);
nand U24458 (N_24458,N_17478,N_19663);
xnor U24459 (N_24459,N_19638,N_18341);
and U24460 (N_24460,N_19460,N_18287);
nor U24461 (N_24461,N_17264,N_16404);
or U24462 (N_24462,N_16367,N_19036);
nand U24463 (N_24463,N_16863,N_19451);
nor U24464 (N_24464,N_17662,N_19786);
or U24465 (N_24465,N_15063,N_18340);
xor U24466 (N_24466,N_16519,N_15030);
nor U24467 (N_24467,N_19301,N_17913);
or U24468 (N_24468,N_17451,N_19175);
or U24469 (N_24469,N_18251,N_15956);
nor U24470 (N_24470,N_15035,N_18425);
or U24471 (N_24471,N_17044,N_17642);
or U24472 (N_24472,N_16247,N_15984);
and U24473 (N_24473,N_18072,N_17346);
or U24474 (N_24474,N_19170,N_17576);
and U24475 (N_24475,N_15535,N_19105);
xnor U24476 (N_24476,N_19453,N_17732);
xor U24477 (N_24477,N_18331,N_18913);
or U24478 (N_24478,N_19459,N_15387);
and U24479 (N_24479,N_16902,N_19332);
xnor U24480 (N_24480,N_15618,N_16673);
nand U24481 (N_24481,N_17690,N_18107);
or U24482 (N_24482,N_17378,N_18055);
xnor U24483 (N_24483,N_19075,N_15223);
nor U24484 (N_24484,N_19519,N_16134);
nor U24485 (N_24485,N_18060,N_16681);
or U24486 (N_24486,N_18866,N_15296);
nor U24487 (N_24487,N_17701,N_17828);
or U24488 (N_24488,N_19511,N_18907);
nand U24489 (N_24489,N_16401,N_18780);
nor U24490 (N_24490,N_16873,N_19945);
xnor U24491 (N_24491,N_19231,N_15036);
and U24492 (N_24492,N_15861,N_17413);
or U24493 (N_24493,N_19154,N_19202);
nand U24494 (N_24494,N_16066,N_17654);
or U24495 (N_24495,N_18910,N_18152);
or U24496 (N_24496,N_19048,N_15447);
xnor U24497 (N_24497,N_18868,N_17478);
or U24498 (N_24498,N_19255,N_16418);
xnor U24499 (N_24499,N_17969,N_18671);
nand U24500 (N_24500,N_17762,N_17918);
nor U24501 (N_24501,N_19141,N_19782);
nand U24502 (N_24502,N_18996,N_19071);
nor U24503 (N_24503,N_15948,N_17889);
nand U24504 (N_24504,N_18929,N_19172);
or U24505 (N_24505,N_17924,N_16215);
xor U24506 (N_24506,N_17802,N_16168);
or U24507 (N_24507,N_15492,N_17090);
nand U24508 (N_24508,N_19433,N_19516);
nand U24509 (N_24509,N_18060,N_17006);
nor U24510 (N_24510,N_19109,N_19085);
xor U24511 (N_24511,N_18049,N_18942);
xnor U24512 (N_24512,N_16498,N_18737);
xor U24513 (N_24513,N_18567,N_17495);
and U24514 (N_24514,N_19334,N_17150);
nand U24515 (N_24515,N_15842,N_15918);
and U24516 (N_24516,N_15067,N_15734);
nor U24517 (N_24517,N_19761,N_19457);
nand U24518 (N_24518,N_19766,N_15434);
nand U24519 (N_24519,N_17096,N_18557);
and U24520 (N_24520,N_17074,N_19668);
and U24521 (N_24521,N_18332,N_15039);
xor U24522 (N_24522,N_17099,N_16324);
and U24523 (N_24523,N_16471,N_19274);
or U24524 (N_24524,N_16853,N_17885);
nand U24525 (N_24525,N_15869,N_18350);
or U24526 (N_24526,N_18457,N_16065);
nor U24527 (N_24527,N_17956,N_18522);
nand U24528 (N_24528,N_16569,N_19337);
nor U24529 (N_24529,N_17273,N_17350);
nor U24530 (N_24530,N_18340,N_17813);
nand U24531 (N_24531,N_16318,N_19330);
nand U24532 (N_24532,N_19056,N_18445);
nand U24533 (N_24533,N_19535,N_18103);
xor U24534 (N_24534,N_19125,N_15063);
xor U24535 (N_24535,N_18817,N_16090);
and U24536 (N_24536,N_18777,N_16692);
or U24537 (N_24537,N_17273,N_19508);
xnor U24538 (N_24538,N_16369,N_16422);
and U24539 (N_24539,N_19196,N_17259);
xor U24540 (N_24540,N_16192,N_15007);
nor U24541 (N_24541,N_19632,N_17325);
nand U24542 (N_24542,N_16297,N_16475);
or U24543 (N_24543,N_17282,N_18072);
xor U24544 (N_24544,N_18022,N_19293);
xor U24545 (N_24545,N_18319,N_19394);
xnor U24546 (N_24546,N_19983,N_15751);
xor U24547 (N_24547,N_17215,N_19615);
or U24548 (N_24548,N_17910,N_19007);
nand U24549 (N_24549,N_18589,N_18816);
nor U24550 (N_24550,N_16088,N_17054);
xnor U24551 (N_24551,N_16697,N_15330);
xor U24552 (N_24552,N_16858,N_17821);
or U24553 (N_24553,N_18575,N_17694);
xor U24554 (N_24554,N_17923,N_19627);
or U24555 (N_24555,N_17933,N_17812);
xor U24556 (N_24556,N_18439,N_17949);
xnor U24557 (N_24557,N_17038,N_15893);
and U24558 (N_24558,N_16818,N_15914);
or U24559 (N_24559,N_18077,N_16237);
nor U24560 (N_24560,N_15818,N_15722);
nor U24561 (N_24561,N_17077,N_17450);
xor U24562 (N_24562,N_17319,N_15129);
nand U24563 (N_24563,N_18242,N_16800);
nor U24564 (N_24564,N_15593,N_17096);
and U24565 (N_24565,N_19443,N_19191);
and U24566 (N_24566,N_17757,N_19432);
and U24567 (N_24567,N_19722,N_19257);
or U24568 (N_24568,N_15555,N_17441);
nand U24569 (N_24569,N_19773,N_19883);
nand U24570 (N_24570,N_15747,N_19733);
nor U24571 (N_24571,N_18478,N_15453);
or U24572 (N_24572,N_15134,N_17256);
nor U24573 (N_24573,N_15780,N_17459);
or U24574 (N_24574,N_19981,N_15411);
nand U24575 (N_24575,N_15831,N_16140);
nand U24576 (N_24576,N_17204,N_16192);
nand U24577 (N_24577,N_15943,N_15663);
nand U24578 (N_24578,N_17068,N_17797);
xnor U24579 (N_24579,N_18629,N_17136);
and U24580 (N_24580,N_16548,N_19150);
nand U24581 (N_24581,N_16322,N_17007);
and U24582 (N_24582,N_19085,N_16097);
and U24583 (N_24583,N_16665,N_19460);
nand U24584 (N_24584,N_15168,N_18686);
nand U24585 (N_24585,N_18757,N_16385);
or U24586 (N_24586,N_15373,N_18825);
xnor U24587 (N_24587,N_18160,N_18683);
or U24588 (N_24588,N_16969,N_15556);
and U24589 (N_24589,N_17988,N_17401);
xor U24590 (N_24590,N_17488,N_17352);
nor U24591 (N_24591,N_19963,N_16682);
xor U24592 (N_24592,N_17764,N_15355);
or U24593 (N_24593,N_19386,N_19089);
or U24594 (N_24594,N_17537,N_16261);
xor U24595 (N_24595,N_17645,N_15874);
nand U24596 (N_24596,N_19591,N_15632);
and U24597 (N_24597,N_19987,N_15204);
or U24598 (N_24598,N_18340,N_19581);
xnor U24599 (N_24599,N_15578,N_16266);
nand U24600 (N_24600,N_19905,N_18488);
xor U24601 (N_24601,N_16232,N_19546);
or U24602 (N_24602,N_17602,N_16791);
nor U24603 (N_24603,N_18269,N_17454);
or U24604 (N_24604,N_18802,N_15012);
nor U24605 (N_24605,N_15773,N_17665);
nor U24606 (N_24606,N_17505,N_17221);
nor U24607 (N_24607,N_17987,N_17103);
or U24608 (N_24608,N_19937,N_19823);
nor U24609 (N_24609,N_16332,N_18901);
and U24610 (N_24610,N_19452,N_19824);
nand U24611 (N_24611,N_18033,N_17200);
nand U24612 (N_24612,N_18730,N_16523);
xor U24613 (N_24613,N_18571,N_17050);
or U24614 (N_24614,N_17014,N_16303);
nand U24615 (N_24615,N_18219,N_19352);
or U24616 (N_24616,N_19976,N_17820);
and U24617 (N_24617,N_15168,N_15649);
nand U24618 (N_24618,N_18156,N_19215);
xor U24619 (N_24619,N_17578,N_18735);
nor U24620 (N_24620,N_17584,N_18400);
xnor U24621 (N_24621,N_15544,N_15177);
or U24622 (N_24622,N_18030,N_18268);
or U24623 (N_24623,N_17416,N_19690);
nand U24624 (N_24624,N_18341,N_18905);
and U24625 (N_24625,N_15194,N_18125);
nand U24626 (N_24626,N_15995,N_19187);
and U24627 (N_24627,N_17587,N_19648);
and U24628 (N_24628,N_15971,N_17680);
nor U24629 (N_24629,N_18947,N_18959);
nand U24630 (N_24630,N_16691,N_16829);
xnor U24631 (N_24631,N_17347,N_18040);
or U24632 (N_24632,N_15067,N_19974);
nor U24633 (N_24633,N_15322,N_18819);
nor U24634 (N_24634,N_18482,N_17818);
or U24635 (N_24635,N_17418,N_19751);
nor U24636 (N_24636,N_15743,N_15558);
xnor U24637 (N_24637,N_16898,N_19605);
nor U24638 (N_24638,N_19592,N_17415);
and U24639 (N_24639,N_16541,N_19283);
nor U24640 (N_24640,N_18543,N_19780);
or U24641 (N_24641,N_17539,N_16450);
nor U24642 (N_24642,N_16364,N_19472);
and U24643 (N_24643,N_19370,N_15109);
nor U24644 (N_24644,N_19138,N_16007);
nor U24645 (N_24645,N_19020,N_18581);
or U24646 (N_24646,N_19934,N_15031);
nor U24647 (N_24647,N_15949,N_19680);
xnor U24648 (N_24648,N_17826,N_19955);
nand U24649 (N_24649,N_19064,N_16048);
nor U24650 (N_24650,N_15878,N_19903);
xnor U24651 (N_24651,N_17926,N_15943);
and U24652 (N_24652,N_16158,N_16926);
xnor U24653 (N_24653,N_16543,N_16497);
or U24654 (N_24654,N_18315,N_17832);
nor U24655 (N_24655,N_16895,N_15195);
xor U24656 (N_24656,N_18157,N_18679);
and U24657 (N_24657,N_15412,N_17645);
xor U24658 (N_24658,N_16763,N_16015);
nor U24659 (N_24659,N_17613,N_16290);
or U24660 (N_24660,N_18450,N_19415);
or U24661 (N_24661,N_15175,N_15540);
or U24662 (N_24662,N_17833,N_16700);
and U24663 (N_24663,N_18758,N_18603);
nand U24664 (N_24664,N_18597,N_16172);
nor U24665 (N_24665,N_19181,N_15595);
nand U24666 (N_24666,N_16025,N_19695);
xnor U24667 (N_24667,N_18303,N_18491);
nand U24668 (N_24668,N_16964,N_16356);
and U24669 (N_24669,N_15654,N_18406);
xor U24670 (N_24670,N_15617,N_18492);
nor U24671 (N_24671,N_18562,N_18490);
and U24672 (N_24672,N_17867,N_15213);
nand U24673 (N_24673,N_15834,N_16009);
nand U24674 (N_24674,N_16548,N_16655);
nor U24675 (N_24675,N_17336,N_17937);
nor U24676 (N_24676,N_16143,N_19730);
and U24677 (N_24677,N_17696,N_18854);
nor U24678 (N_24678,N_16069,N_18235);
or U24679 (N_24679,N_16113,N_15116);
nand U24680 (N_24680,N_19621,N_15289);
and U24681 (N_24681,N_18029,N_15797);
and U24682 (N_24682,N_16966,N_17126);
nor U24683 (N_24683,N_15283,N_15087);
or U24684 (N_24684,N_19881,N_16002);
nor U24685 (N_24685,N_18943,N_17226);
and U24686 (N_24686,N_17315,N_16291);
xor U24687 (N_24687,N_17427,N_16977);
and U24688 (N_24688,N_17587,N_19954);
xnor U24689 (N_24689,N_16735,N_15180);
nand U24690 (N_24690,N_16266,N_17007);
nand U24691 (N_24691,N_17082,N_15797);
or U24692 (N_24692,N_18354,N_17830);
nor U24693 (N_24693,N_17171,N_16534);
or U24694 (N_24694,N_18370,N_18531);
and U24695 (N_24695,N_17594,N_19550);
or U24696 (N_24696,N_17209,N_15778);
nor U24697 (N_24697,N_17580,N_18485);
or U24698 (N_24698,N_18030,N_15387);
nand U24699 (N_24699,N_19228,N_16928);
xor U24700 (N_24700,N_15207,N_19731);
nand U24701 (N_24701,N_17237,N_17485);
nand U24702 (N_24702,N_17479,N_17246);
and U24703 (N_24703,N_16298,N_17377);
and U24704 (N_24704,N_17910,N_15487);
nor U24705 (N_24705,N_18546,N_17783);
nand U24706 (N_24706,N_16383,N_16477);
nor U24707 (N_24707,N_15493,N_19033);
nand U24708 (N_24708,N_19137,N_16787);
and U24709 (N_24709,N_18120,N_18587);
or U24710 (N_24710,N_18533,N_17279);
nand U24711 (N_24711,N_19977,N_19315);
and U24712 (N_24712,N_18443,N_19658);
xor U24713 (N_24713,N_16484,N_17735);
or U24714 (N_24714,N_18551,N_17316);
or U24715 (N_24715,N_18190,N_19970);
nand U24716 (N_24716,N_17279,N_16165);
and U24717 (N_24717,N_16492,N_16639);
or U24718 (N_24718,N_18865,N_18359);
nor U24719 (N_24719,N_17739,N_18068);
and U24720 (N_24720,N_17958,N_17870);
xnor U24721 (N_24721,N_18922,N_18610);
nand U24722 (N_24722,N_16476,N_19900);
xnor U24723 (N_24723,N_16929,N_19577);
or U24724 (N_24724,N_17159,N_19890);
and U24725 (N_24725,N_18869,N_16472);
xnor U24726 (N_24726,N_17035,N_15980);
and U24727 (N_24727,N_19464,N_17098);
nor U24728 (N_24728,N_16516,N_18934);
nand U24729 (N_24729,N_18049,N_16662);
xor U24730 (N_24730,N_19571,N_16448);
and U24731 (N_24731,N_19927,N_17674);
nor U24732 (N_24732,N_17040,N_19953);
xnor U24733 (N_24733,N_17439,N_19585);
xnor U24734 (N_24734,N_15329,N_16283);
nand U24735 (N_24735,N_16915,N_18669);
and U24736 (N_24736,N_18633,N_17522);
nor U24737 (N_24737,N_19395,N_15033);
nand U24738 (N_24738,N_15091,N_16313);
xor U24739 (N_24739,N_16443,N_19509);
nor U24740 (N_24740,N_15791,N_17691);
and U24741 (N_24741,N_18642,N_19402);
or U24742 (N_24742,N_18249,N_15179);
nor U24743 (N_24743,N_19440,N_15464);
and U24744 (N_24744,N_15599,N_19884);
and U24745 (N_24745,N_18229,N_19795);
or U24746 (N_24746,N_18817,N_16285);
nor U24747 (N_24747,N_17129,N_17343);
nor U24748 (N_24748,N_15799,N_17506);
xor U24749 (N_24749,N_17596,N_17706);
or U24750 (N_24750,N_16367,N_15909);
xor U24751 (N_24751,N_16665,N_19310);
or U24752 (N_24752,N_18458,N_17666);
or U24753 (N_24753,N_15065,N_17330);
and U24754 (N_24754,N_19280,N_16428);
xor U24755 (N_24755,N_17332,N_19107);
nor U24756 (N_24756,N_19137,N_15237);
nand U24757 (N_24757,N_15331,N_16325);
nor U24758 (N_24758,N_17499,N_15094);
and U24759 (N_24759,N_18187,N_18433);
xnor U24760 (N_24760,N_18928,N_18525);
nor U24761 (N_24761,N_16275,N_18063);
and U24762 (N_24762,N_15353,N_19812);
or U24763 (N_24763,N_17725,N_15924);
or U24764 (N_24764,N_19558,N_19694);
xnor U24765 (N_24765,N_16788,N_19258);
nor U24766 (N_24766,N_18966,N_19938);
and U24767 (N_24767,N_16994,N_19328);
xor U24768 (N_24768,N_17328,N_18153);
and U24769 (N_24769,N_15860,N_19209);
or U24770 (N_24770,N_19337,N_17237);
and U24771 (N_24771,N_15471,N_19998);
xnor U24772 (N_24772,N_18158,N_16897);
or U24773 (N_24773,N_17410,N_16939);
xnor U24774 (N_24774,N_16266,N_17506);
nor U24775 (N_24775,N_18281,N_17605);
nor U24776 (N_24776,N_18045,N_16935);
nand U24777 (N_24777,N_15983,N_18155);
xor U24778 (N_24778,N_17400,N_18613);
and U24779 (N_24779,N_15992,N_18562);
and U24780 (N_24780,N_16342,N_16905);
xnor U24781 (N_24781,N_19746,N_16535);
xor U24782 (N_24782,N_15534,N_19736);
xor U24783 (N_24783,N_15299,N_18395);
xor U24784 (N_24784,N_19456,N_15227);
nand U24785 (N_24785,N_16170,N_17787);
nor U24786 (N_24786,N_19758,N_15482);
and U24787 (N_24787,N_17214,N_15780);
xnor U24788 (N_24788,N_15908,N_17477);
and U24789 (N_24789,N_16975,N_16072);
nand U24790 (N_24790,N_18328,N_15465);
nand U24791 (N_24791,N_18605,N_18861);
nor U24792 (N_24792,N_17769,N_18319);
nand U24793 (N_24793,N_18411,N_15673);
or U24794 (N_24794,N_15650,N_18040);
nand U24795 (N_24795,N_15545,N_18141);
xor U24796 (N_24796,N_17401,N_16600);
xnor U24797 (N_24797,N_17299,N_16574);
and U24798 (N_24798,N_19325,N_17714);
or U24799 (N_24799,N_15152,N_17039);
and U24800 (N_24800,N_18361,N_17574);
nor U24801 (N_24801,N_16458,N_16552);
or U24802 (N_24802,N_15368,N_18856);
and U24803 (N_24803,N_17455,N_15504);
xnor U24804 (N_24804,N_15260,N_17483);
or U24805 (N_24805,N_17183,N_17925);
and U24806 (N_24806,N_15108,N_19700);
xnor U24807 (N_24807,N_15399,N_18126);
nand U24808 (N_24808,N_17083,N_18190);
xnor U24809 (N_24809,N_15290,N_16301);
and U24810 (N_24810,N_18495,N_17704);
nand U24811 (N_24811,N_16217,N_17361);
nor U24812 (N_24812,N_18021,N_19728);
nand U24813 (N_24813,N_19616,N_16358);
or U24814 (N_24814,N_17246,N_15067);
nand U24815 (N_24815,N_15494,N_19909);
nor U24816 (N_24816,N_16753,N_18432);
or U24817 (N_24817,N_15231,N_19446);
and U24818 (N_24818,N_16074,N_17703);
or U24819 (N_24819,N_15861,N_19088);
nand U24820 (N_24820,N_18234,N_18413);
or U24821 (N_24821,N_16588,N_16201);
nand U24822 (N_24822,N_16030,N_18408);
nor U24823 (N_24823,N_16056,N_19212);
nand U24824 (N_24824,N_15758,N_16402);
or U24825 (N_24825,N_18218,N_16908);
or U24826 (N_24826,N_15327,N_15251);
or U24827 (N_24827,N_17720,N_18591);
or U24828 (N_24828,N_19369,N_19953);
nor U24829 (N_24829,N_18772,N_19713);
xor U24830 (N_24830,N_19059,N_19719);
nor U24831 (N_24831,N_19128,N_18559);
or U24832 (N_24832,N_15948,N_18722);
or U24833 (N_24833,N_19520,N_15003);
nand U24834 (N_24834,N_17371,N_16697);
and U24835 (N_24835,N_16128,N_15877);
or U24836 (N_24836,N_18009,N_17413);
nand U24837 (N_24837,N_17044,N_19716);
nand U24838 (N_24838,N_16462,N_19533);
nor U24839 (N_24839,N_16649,N_16551);
and U24840 (N_24840,N_18310,N_16920);
and U24841 (N_24841,N_17602,N_15425);
or U24842 (N_24842,N_19491,N_16249);
or U24843 (N_24843,N_18674,N_16450);
nor U24844 (N_24844,N_16840,N_16229);
nor U24845 (N_24845,N_19822,N_16658);
xnor U24846 (N_24846,N_19792,N_18643);
or U24847 (N_24847,N_18520,N_19283);
and U24848 (N_24848,N_19770,N_16763);
xnor U24849 (N_24849,N_15068,N_19434);
nand U24850 (N_24850,N_18700,N_18300);
xor U24851 (N_24851,N_18072,N_16634);
and U24852 (N_24852,N_16054,N_19475);
nand U24853 (N_24853,N_19104,N_19122);
nand U24854 (N_24854,N_16716,N_18461);
xnor U24855 (N_24855,N_15445,N_18402);
nor U24856 (N_24856,N_16751,N_18698);
or U24857 (N_24857,N_18078,N_15261);
and U24858 (N_24858,N_19867,N_16087);
and U24859 (N_24859,N_17294,N_17395);
or U24860 (N_24860,N_17756,N_15095);
nand U24861 (N_24861,N_15307,N_19865);
xnor U24862 (N_24862,N_18586,N_15796);
xnor U24863 (N_24863,N_17614,N_15519);
xor U24864 (N_24864,N_16973,N_19614);
nor U24865 (N_24865,N_16667,N_19672);
nor U24866 (N_24866,N_18333,N_15663);
xnor U24867 (N_24867,N_16894,N_18141);
nand U24868 (N_24868,N_18625,N_15736);
and U24869 (N_24869,N_16159,N_18206);
nand U24870 (N_24870,N_16474,N_16111);
or U24871 (N_24871,N_19759,N_16167);
nand U24872 (N_24872,N_18155,N_18471);
nand U24873 (N_24873,N_19742,N_15139);
or U24874 (N_24874,N_15517,N_17774);
nor U24875 (N_24875,N_16174,N_16312);
xor U24876 (N_24876,N_18761,N_17119);
or U24877 (N_24877,N_15164,N_19065);
or U24878 (N_24878,N_15757,N_16804);
nor U24879 (N_24879,N_16224,N_15787);
and U24880 (N_24880,N_15265,N_16054);
nor U24881 (N_24881,N_17639,N_16547);
xor U24882 (N_24882,N_17398,N_17301);
nand U24883 (N_24883,N_15117,N_17862);
nor U24884 (N_24884,N_16572,N_16219);
nand U24885 (N_24885,N_15598,N_18925);
xor U24886 (N_24886,N_17274,N_16253);
xnor U24887 (N_24887,N_17812,N_15492);
nand U24888 (N_24888,N_16444,N_16788);
xnor U24889 (N_24889,N_17647,N_15136);
xnor U24890 (N_24890,N_16014,N_15181);
nand U24891 (N_24891,N_17934,N_18119);
nand U24892 (N_24892,N_16347,N_18577);
nand U24893 (N_24893,N_19177,N_17752);
xor U24894 (N_24894,N_17660,N_19861);
and U24895 (N_24895,N_15356,N_17061);
and U24896 (N_24896,N_17159,N_16094);
xor U24897 (N_24897,N_19490,N_15044);
and U24898 (N_24898,N_16169,N_18126);
xnor U24899 (N_24899,N_15141,N_15384);
or U24900 (N_24900,N_18300,N_15343);
nand U24901 (N_24901,N_17637,N_18236);
xor U24902 (N_24902,N_18533,N_19628);
and U24903 (N_24903,N_15282,N_18516);
xor U24904 (N_24904,N_16947,N_16809);
or U24905 (N_24905,N_15799,N_18727);
and U24906 (N_24906,N_18929,N_16391);
nor U24907 (N_24907,N_17849,N_16726);
nand U24908 (N_24908,N_15881,N_15991);
nand U24909 (N_24909,N_16069,N_17627);
and U24910 (N_24910,N_18240,N_18173);
xnor U24911 (N_24911,N_17493,N_19782);
nor U24912 (N_24912,N_17502,N_17018);
and U24913 (N_24913,N_17517,N_16762);
and U24914 (N_24914,N_19677,N_17271);
xnor U24915 (N_24915,N_19731,N_16826);
and U24916 (N_24916,N_19676,N_18801);
nor U24917 (N_24917,N_15867,N_15598);
nor U24918 (N_24918,N_15334,N_19365);
and U24919 (N_24919,N_18838,N_19082);
xnor U24920 (N_24920,N_18947,N_16473);
and U24921 (N_24921,N_15614,N_19269);
nand U24922 (N_24922,N_19806,N_17547);
nor U24923 (N_24923,N_19865,N_17876);
and U24924 (N_24924,N_15260,N_17238);
nor U24925 (N_24925,N_19176,N_19437);
and U24926 (N_24926,N_16925,N_15016);
nor U24927 (N_24927,N_16182,N_16268);
or U24928 (N_24928,N_15068,N_16667);
or U24929 (N_24929,N_15326,N_16201);
or U24930 (N_24930,N_16563,N_17093);
or U24931 (N_24931,N_16701,N_16200);
xor U24932 (N_24932,N_18617,N_15343);
nor U24933 (N_24933,N_19864,N_16370);
xnor U24934 (N_24934,N_17531,N_15631);
xnor U24935 (N_24935,N_15843,N_17218);
nor U24936 (N_24936,N_19200,N_15375);
xnor U24937 (N_24937,N_19423,N_16529);
or U24938 (N_24938,N_19535,N_18159);
or U24939 (N_24939,N_19454,N_19980);
nand U24940 (N_24940,N_18327,N_15512);
nor U24941 (N_24941,N_18142,N_15381);
or U24942 (N_24942,N_16497,N_19852);
and U24943 (N_24943,N_19064,N_15933);
nor U24944 (N_24944,N_16653,N_19084);
or U24945 (N_24945,N_18679,N_15873);
xnor U24946 (N_24946,N_17314,N_18585);
and U24947 (N_24947,N_15798,N_19659);
nand U24948 (N_24948,N_15908,N_17904);
or U24949 (N_24949,N_15838,N_15378);
nand U24950 (N_24950,N_18306,N_16825);
and U24951 (N_24951,N_18392,N_17592);
nor U24952 (N_24952,N_19678,N_17109);
or U24953 (N_24953,N_16182,N_19062);
nand U24954 (N_24954,N_16742,N_19298);
or U24955 (N_24955,N_15948,N_17278);
or U24956 (N_24956,N_16995,N_16605);
or U24957 (N_24957,N_15821,N_17674);
nand U24958 (N_24958,N_15666,N_19490);
nor U24959 (N_24959,N_18136,N_16157);
or U24960 (N_24960,N_17704,N_19008);
nand U24961 (N_24961,N_15589,N_16378);
nand U24962 (N_24962,N_16917,N_15578);
or U24963 (N_24963,N_19941,N_15123);
nor U24964 (N_24964,N_16418,N_18006);
nand U24965 (N_24965,N_16659,N_16381);
xor U24966 (N_24966,N_17732,N_18688);
and U24967 (N_24967,N_15731,N_18112);
nor U24968 (N_24968,N_15219,N_16066);
and U24969 (N_24969,N_17080,N_18985);
nand U24970 (N_24970,N_17653,N_17211);
xnor U24971 (N_24971,N_18788,N_18717);
xor U24972 (N_24972,N_17199,N_16181);
nor U24973 (N_24973,N_16400,N_16263);
and U24974 (N_24974,N_19412,N_19651);
or U24975 (N_24975,N_18324,N_16037);
xor U24976 (N_24976,N_15555,N_17998);
nand U24977 (N_24977,N_17717,N_16818);
and U24978 (N_24978,N_17265,N_18121);
xor U24979 (N_24979,N_18249,N_17363);
and U24980 (N_24980,N_19495,N_15271);
or U24981 (N_24981,N_17801,N_15090);
or U24982 (N_24982,N_17047,N_15033);
nor U24983 (N_24983,N_18859,N_15186);
xor U24984 (N_24984,N_16921,N_16093);
xor U24985 (N_24985,N_18921,N_15262);
xor U24986 (N_24986,N_15640,N_15190);
or U24987 (N_24987,N_19850,N_16442);
nand U24988 (N_24988,N_15700,N_15268);
xnor U24989 (N_24989,N_15116,N_18731);
and U24990 (N_24990,N_19748,N_15080);
nor U24991 (N_24991,N_19863,N_15301);
nand U24992 (N_24992,N_19291,N_15409);
xnor U24993 (N_24993,N_18680,N_19683);
xnor U24994 (N_24994,N_18217,N_17739);
nand U24995 (N_24995,N_15894,N_18806);
or U24996 (N_24996,N_18815,N_19090);
nand U24997 (N_24997,N_18272,N_19408);
xnor U24998 (N_24998,N_17659,N_18461);
and U24999 (N_24999,N_18087,N_15004);
or UO_0 (O_0,N_23941,N_21712);
nor UO_1 (O_1,N_20960,N_23423);
or UO_2 (O_2,N_24130,N_23586);
nand UO_3 (O_3,N_21483,N_24329);
and UO_4 (O_4,N_21745,N_22589);
xor UO_5 (O_5,N_24437,N_21218);
xnor UO_6 (O_6,N_22269,N_21367);
and UO_7 (O_7,N_22063,N_21938);
nand UO_8 (O_8,N_20609,N_20538);
nor UO_9 (O_9,N_20639,N_20184);
nor UO_10 (O_10,N_24044,N_23668);
and UO_11 (O_11,N_21455,N_23220);
nand UO_12 (O_12,N_22710,N_21960);
nand UO_13 (O_13,N_22544,N_22510);
nor UO_14 (O_14,N_20434,N_23042);
xnor UO_15 (O_15,N_24614,N_21309);
or UO_16 (O_16,N_22053,N_24796);
nand UO_17 (O_17,N_20642,N_21018);
and UO_18 (O_18,N_22461,N_23964);
xnor UO_19 (O_19,N_21910,N_21686);
nor UO_20 (O_20,N_22331,N_23300);
nor UO_21 (O_21,N_24232,N_21031);
nand UO_22 (O_22,N_22088,N_22062);
or UO_23 (O_23,N_23530,N_20723);
nand UO_24 (O_24,N_24394,N_23125);
xor UO_25 (O_25,N_23713,N_22697);
nor UO_26 (O_26,N_23712,N_20850);
xnor UO_27 (O_27,N_20476,N_21981);
and UO_28 (O_28,N_24009,N_24586);
nor UO_29 (O_29,N_20814,N_20893);
nor UO_30 (O_30,N_24647,N_20849);
nor UO_31 (O_31,N_24198,N_23771);
xnor UO_32 (O_32,N_20338,N_21368);
xnor UO_33 (O_33,N_21915,N_22672);
nor UO_34 (O_34,N_24295,N_22638);
nor UO_35 (O_35,N_24443,N_21462);
and UO_36 (O_36,N_22554,N_20010);
and UO_37 (O_37,N_23060,N_22590);
and UO_38 (O_38,N_20967,N_21542);
and UO_39 (O_39,N_21162,N_22270);
nor UO_40 (O_40,N_20572,N_22124);
xor UO_41 (O_41,N_21648,N_21556);
and UO_42 (O_42,N_23926,N_22962);
nor UO_43 (O_43,N_23450,N_22522);
or UO_44 (O_44,N_24734,N_24100);
xor UO_45 (O_45,N_24002,N_23947);
or UO_46 (O_46,N_22965,N_24075);
xnor UO_47 (O_47,N_21053,N_20734);
and UO_48 (O_48,N_20680,N_22006);
nor UO_49 (O_49,N_23279,N_24059);
nor UO_50 (O_50,N_21099,N_22969);
nand UO_51 (O_51,N_20043,N_20700);
nand UO_52 (O_52,N_20977,N_24165);
nand UO_53 (O_53,N_22203,N_24761);
nand UO_54 (O_54,N_20428,N_22344);
nor UO_55 (O_55,N_23293,N_20714);
and UO_56 (O_56,N_20682,N_22769);
or UO_57 (O_57,N_24216,N_22845);
nor UO_58 (O_58,N_23456,N_21216);
xor UO_59 (O_59,N_20219,N_24744);
nor UO_60 (O_60,N_23471,N_24189);
and UO_61 (O_61,N_22956,N_23349);
nand UO_62 (O_62,N_22816,N_20267);
nor UO_63 (O_63,N_22410,N_21714);
and UO_64 (O_64,N_22399,N_23266);
and UO_65 (O_65,N_23911,N_24979);
or UO_66 (O_66,N_20231,N_21963);
xor UO_67 (O_67,N_23038,N_22610);
nand UO_68 (O_68,N_24397,N_21060);
nor UO_69 (O_69,N_24867,N_21424);
xor UO_70 (O_70,N_22139,N_23663);
or UO_71 (O_71,N_20055,N_24308);
or UO_72 (O_72,N_22222,N_23968);
xnor UO_73 (O_73,N_23667,N_20891);
xor UO_74 (O_74,N_24128,N_24903);
or UO_75 (O_75,N_22333,N_20564);
nor UO_76 (O_76,N_24836,N_24309);
nand UO_77 (O_77,N_20945,N_20671);
nand UO_78 (O_78,N_22953,N_23785);
xnor UO_79 (O_79,N_22649,N_22683);
nor UO_80 (O_80,N_23055,N_24401);
nor UO_81 (O_81,N_20512,N_22308);
nand UO_82 (O_82,N_20786,N_21111);
and UO_83 (O_83,N_23736,N_21718);
nor UO_84 (O_84,N_24087,N_23270);
nand UO_85 (O_85,N_20205,N_23682);
nand UO_86 (O_86,N_20493,N_20997);
or UO_87 (O_87,N_23148,N_24465);
and UO_88 (O_88,N_21249,N_23075);
nand UO_89 (O_89,N_21756,N_21593);
xnor UO_90 (O_90,N_20106,N_24580);
or UO_91 (O_91,N_22244,N_24881);
nor UO_92 (O_92,N_23359,N_21875);
nor UO_93 (O_93,N_21588,N_24885);
xor UO_94 (O_94,N_22856,N_24337);
xnor UO_95 (O_95,N_20330,N_21548);
nand UO_96 (O_96,N_22583,N_20712);
or UO_97 (O_97,N_24967,N_23961);
and UO_98 (O_98,N_23217,N_24844);
or UO_99 (O_99,N_22411,N_24793);
nor UO_100 (O_100,N_24519,N_23443);
nand UO_101 (O_101,N_22709,N_23178);
nand UO_102 (O_102,N_21510,N_23153);
or UO_103 (O_103,N_23219,N_22384);
and UO_104 (O_104,N_23354,N_21431);
nor UO_105 (O_105,N_23717,N_24006);
or UO_106 (O_106,N_23666,N_21700);
nor UO_107 (O_107,N_23147,N_22043);
or UO_108 (O_108,N_24234,N_21208);
nand UO_109 (O_109,N_24038,N_21472);
nor UO_110 (O_110,N_22357,N_24791);
xnor UO_111 (O_111,N_23631,N_23959);
nand UO_112 (O_112,N_23620,N_21790);
and UO_113 (O_113,N_23429,N_24866);
xor UO_114 (O_114,N_22051,N_21672);
xnor UO_115 (O_115,N_24490,N_23234);
nand UO_116 (O_116,N_20166,N_24753);
or UO_117 (O_117,N_23774,N_21049);
or UO_118 (O_118,N_21059,N_23969);
nor UO_119 (O_119,N_21250,N_21450);
and UO_120 (O_120,N_24655,N_20042);
xor UO_121 (O_121,N_22689,N_23643);
or UO_122 (O_122,N_23171,N_22517);
nand UO_123 (O_123,N_23348,N_24233);
or UO_124 (O_124,N_20340,N_22827);
xor UO_125 (O_125,N_21584,N_24031);
xnor UO_126 (O_126,N_24780,N_24151);
and UO_127 (O_127,N_24719,N_21377);
or UO_128 (O_128,N_24133,N_21478);
nand UO_129 (O_129,N_21295,N_20774);
or UO_130 (O_130,N_23369,N_20618);
and UO_131 (O_131,N_20550,N_21928);
nor UO_132 (O_132,N_20212,N_23653);
or UO_133 (O_133,N_23209,N_20073);
nand UO_134 (O_134,N_22733,N_22307);
nor UO_135 (O_135,N_22225,N_20265);
nand UO_136 (O_136,N_24998,N_20364);
and UO_137 (O_137,N_22983,N_20681);
nand UO_138 (O_138,N_20819,N_20821);
nand UO_139 (O_139,N_22398,N_20225);
and UO_140 (O_140,N_20300,N_20115);
and UO_141 (O_141,N_22746,N_24116);
xnor UO_142 (O_142,N_23843,N_21345);
and UO_143 (O_143,N_20907,N_20617);
nor UO_144 (O_144,N_21738,N_23294);
or UO_145 (O_145,N_22444,N_20736);
and UO_146 (O_146,N_24702,N_21374);
xor UO_147 (O_147,N_24494,N_21573);
nor UO_148 (O_148,N_20074,N_21895);
xnor UO_149 (O_149,N_22581,N_24896);
nor UO_150 (O_150,N_24576,N_24956);
xor UO_151 (O_151,N_20366,N_20585);
xnor UO_152 (O_152,N_22970,N_22042);
or UO_153 (O_153,N_21489,N_23504);
or UO_154 (O_154,N_23155,N_21400);
xnor UO_155 (O_155,N_21457,N_22933);
or UO_156 (O_156,N_24846,N_22458);
xnor UO_157 (O_157,N_20780,N_23684);
xor UO_158 (O_158,N_24676,N_23541);
nand UO_159 (O_159,N_24313,N_23116);
nand UO_160 (O_160,N_21526,N_21505);
xnor UO_161 (O_161,N_21333,N_24563);
and UO_162 (O_162,N_24848,N_23296);
nand UO_163 (O_163,N_24681,N_20645);
nand UO_164 (O_164,N_24579,N_24657);
and UO_165 (O_165,N_21936,N_22028);
and UO_166 (O_166,N_24714,N_20095);
and UO_167 (O_167,N_24029,N_24078);
xnor UO_168 (O_168,N_22406,N_23434);
nand UO_169 (O_169,N_21105,N_21386);
xnor UO_170 (O_170,N_21007,N_24334);
or UO_171 (O_171,N_23262,N_23253);
or UO_172 (O_172,N_24854,N_22311);
xnor UO_173 (O_173,N_23345,N_22608);
nor UO_174 (O_174,N_21691,N_22240);
nor UO_175 (O_175,N_20677,N_21735);
xor UO_176 (O_176,N_24431,N_23566);
nor UO_177 (O_177,N_20531,N_23909);
nor UO_178 (O_178,N_20623,N_24514);
xnor UO_179 (O_179,N_22038,N_21382);
and UO_180 (O_180,N_24759,N_24652);
nor UO_181 (O_181,N_23996,N_23769);
nor UO_182 (O_182,N_23740,N_21114);
and UO_183 (O_183,N_21395,N_20369);
or UO_184 (O_184,N_21787,N_22516);
nand UO_185 (O_185,N_23872,N_20752);
or UO_186 (O_186,N_23536,N_20915);
nor UO_187 (O_187,N_20100,N_21256);
and UO_188 (O_188,N_21322,N_21279);
nor UO_189 (O_189,N_22732,N_21894);
nand UO_190 (O_190,N_21155,N_21914);
nand UO_191 (O_191,N_24178,N_23379);
or UO_192 (O_192,N_20549,N_21587);
nand UO_193 (O_193,N_21530,N_24725);
nor UO_194 (O_194,N_22982,N_24975);
nor UO_195 (O_195,N_22931,N_21784);
xor UO_196 (O_196,N_24414,N_22193);
xor UO_197 (O_197,N_20740,N_21062);
nand UO_198 (O_198,N_24455,N_24080);
and UO_199 (O_199,N_20876,N_20655);
xor UO_200 (O_200,N_21179,N_24727);
and UO_201 (O_201,N_21426,N_21680);
xor UO_202 (O_202,N_24858,N_24524);
nand UO_203 (O_203,N_22242,N_22105);
nor UO_204 (O_204,N_20746,N_22603);
and UO_205 (O_205,N_24730,N_24560);
and UO_206 (O_206,N_21968,N_21624);
nor UO_207 (O_207,N_24572,N_24870);
nand UO_208 (O_208,N_22415,N_21535);
and UO_209 (O_209,N_24390,N_24926);
nor UO_210 (O_210,N_21855,N_20383);
nor UO_211 (O_211,N_20005,N_20803);
nand UO_212 (O_212,N_20853,N_20435);
xnor UO_213 (O_213,N_23567,N_20889);
or UO_214 (O_214,N_20457,N_23772);
or UO_215 (O_215,N_20593,N_24473);
or UO_216 (O_216,N_21572,N_20202);
nor UO_217 (O_217,N_24668,N_21054);
nor UO_218 (O_218,N_20912,N_22747);
nor UO_219 (O_219,N_21092,N_22853);
and UO_220 (O_220,N_20255,N_23347);
nor UO_221 (O_221,N_20581,N_22945);
or UO_222 (O_222,N_22402,N_24122);
xor UO_223 (O_223,N_21101,N_20251);
and UO_224 (O_224,N_21028,N_21882);
nand UO_225 (O_225,N_22401,N_20379);
and UO_226 (O_226,N_22648,N_21673);
and UO_227 (O_227,N_22736,N_20471);
or UO_228 (O_228,N_20773,N_24330);
nor UO_229 (O_229,N_20494,N_23989);
and UO_230 (O_230,N_22570,N_21722);
xor UO_231 (O_231,N_22453,N_21922);
nor UO_232 (O_232,N_21660,N_21474);
nor UO_233 (O_233,N_22434,N_22324);
or UO_234 (O_234,N_21293,N_24598);
nor UO_235 (O_235,N_22609,N_22563);
nand UO_236 (O_236,N_24994,N_21775);
xnor UO_237 (O_237,N_20548,N_21086);
and UO_238 (O_238,N_22332,N_21750);
nor UO_239 (O_239,N_22219,N_23890);
and UO_240 (O_240,N_20007,N_22295);
or UO_241 (O_241,N_24432,N_24248);
nand UO_242 (O_242,N_20155,N_22059);
nand UO_243 (O_243,N_23627,N_24296);
xnor UO_244 (O_244,N_21183,N_22012);
nor UO_245 (O_245,N_20896,N_22126);
or UO_246 (O_246,N_21520,N_21365);
nor UO_247 (O_247,N_21363,N_24847);
xnor UO_248 (O_248,N_22941,N_22044);
nor UO_249 (O_249,N_21834,N_24677);
or UO_250 (O_250,N_22883,N_20668);
or UO_251 (O_251,N_20800,N_23309);
and UO_252 (O_252,N_20440,N_23795);
and UO_253 (O_253,N_22993,N_21291);
and UO_254 (O_254,N_22984,N_22820);
nand UO_255 (O_255,N_24489,N_21658);
nor UO_256 (O_256,N_22771,N_24521);
nor UO_257 (O_257,N_22900,N_23860);
xor UO_258 (O_258,N_24539,N_22862);
or UO_259 (O_259,N_21788,N_20670);
xor UO_260 (O_260,N_24695,N_23855);
and UO_261 (O_261,N_24005,N_21666);
nor UO_262 (O_262,N_23592,N_23021);
nor UO_263 (O_263,N_21034,N_20707);
and UO_264 (O_264,N_24747,N_21956);
and UO_265 (O_265,N_24169,N_22418);
nand UO_266 (O_266,N_21820,N_24751);
nand UO_267 (O_267,N_24193,N_23879);
nand UO_268 (O_268,N_20477,N_20611);
nand UO_269 (O_269,N_22760,N_21642);
and UO_270 (O_270,N_21926,N_21892);
and UO_271 (O_271,N_20802,N_23696);
or UO_272 (O_272,N_20273,N_24611);
xor UO_273 (O_273,N_20986,N_21888);
nand UO_274 (O_274,N_24980,N_23632);
nand UO_275 (O_275,N_24768,N_20455);
and UO_276 (O_276,N_22069,N_24673);
nand UO_277 (O_277,N_22918,N_20016);
nor UO_278 (O_278,N_24415,N_22835);
nor UO_279 (O_279,N_20976,N_20336);
xor UO_280 (O_280,N_23405,N_23120);
or UO_281 (O_281,N_22573,N_24205);
and UO_282 (O_282,N_24978,N_20710);
or UO_283 (O_283,N_21889,N_23917);
or UO_284 (O_284,N_23049,N_24860);
nand UO_285 (O_285,N_24319,N_20378);
or UO_286 (O_286,N_20018,N_20135);
nand UO_287 (O_287,N_22194,N_20067);
nand UO_288 (O_288,N_21934,N_20597);
nand UO_289 (O_289,N_21501,N_20984);
and UO_290 (O_290,N_23818,N_24594);
and UO_291 (O_291,N_20706,N_21523);
nor UO_292 (O_292,N_21688,N_21271);
nor UO_293 (O_293,N_23353,N_24255);
nor UO_294 (O_294,N_23970,N_20243);
nor UO_295 (O_295,N_23000,N_22299);
and UO_296 (O_296,N_24571,N_20091);
xor UO_297 (O_297,N_21187,N_24053);
or UO_298 (O_298,N_22076,N_21470);
xnor UO_299 (O_299,N_21194,N_24213);
nor UO_300 (O_300,N_21871,N_22750);
and UO_301 (O_301,N_24051,N_23614);
nor UO_302 (O_302,N_24821,N_23635);
and UO_303 (O_303,N_22807,N_21940);
xnor UO_304 (O_304,N_23001,N_20824);
or UO_305 (O_305,N_20316,N_21610);
nor UO_306 (O_306,N_21445,N_24850);
xor UO_307 (O_307,N_23256,N_21220);
and UO_308 (O_308,N_21169,N_21324);
nand UO_309 (O_309,N_20583,N_24621);
and UO_310 (O_310,N_21244,N_24062);
or UO_311 (O_311,N_20783,N_22146);
or UO_312 (O_312,N_20387,N_22154);
nand UO_313 (O_313,N_24593,N_22990);
and UO_314 (O_314,N_22678,N_24360);
xor UO_315 (O_315,N_22694,N_21048);
nand UO_316 (O_316,N_20266,N_24012);
or UO_317 (O_317,N_21818,N_20818);
or UO_318 (O_318,N_22768,N_21467);
or UO_319 (O_319,N_20913,N_21930);
or UO_320 (O_320,N_20761,N_23641);
or UO_321 (O_321,N_24274,N_22048);
nand UO_322 (O_322,N_21221,N_23842);
or UO_323 (O_323,N_21633,N_20835);
nor UO_324 (O_324,N_24990,N_20506);
nor UO_325 (O_325,N_20724,N_21089);
xnor UO_326 (O_326,N_20442,N_21628);
and UO_327 (O_327,N_22278,N_21631);
nor UO_328 (O_328,N_24412,N_24789);
and UO_329 (O_329,N_24762,N_23956);
xor UO_330 (O_330,N_21947,N_23494);
nand UO_331 (O_331,N_23084,N_22096);
nor UO_332 (O_332,N_20662,N_22192);
xnor UO_333 (O_333,N_23876,N_20809);
nand UO_334 (O_334,N_22874,N_21067);
nor UO_335 (O_335,N_21438,N_23849);
nor UO_336 (O_336,N_21303,N_21329);
nand UO_337 (O_337,N_23323,N_21697);
xor UO_338 (O_338,N_24946,N_21744);
or UO_339 (O_339,N_23810,N_21134);
nand UO_340 (O_340,N_20546,N_23077);
and UO_341 (O_341,N_24684,N_23221);
and UO_342 (O_342,N_24023,N_20813);
nor UO_343 (O_343,N_21824,N_24121);
nor UO_344 (O_344,N_24585,N_22375);
or UO_345 (O_345,N_20995,N_20590);
nand UO_346 (O_346,N_24426,N_21094);
nand UO_347 (O_347,N_20040,N_20154);
nor UO_348 (O_348,N_23064,N_20388);
or UO_349 (O_349,N_21172,N_23111);
and UO_350 (O_350,N_21138,N_24389);
or UO_351 (O_351,N_24500,N_23179);
nor UO_352 (O_352,N_22452,N_24823);
and UO_353 (O_353,N_20547,N_20081);
or UO_354 (O_354,N_21524,N_21879);
nand UO_355 (O_355,N_21635,N_20374);
or UO_356 (O_356,N_21181,N_22585);
nand UO_357 (O_357,N_20973,N_20906);
nor UO_358 (O_358,N_23794,N_22850);
or UO_359 (O_359,N_24067,N_21612);
xnor UO_360 (O_360,N_23441,N_21201);
xnor UO_361 (O_361,N_23339,N_20620);
or UO_362 (O_362,N_22915,N_22023);
nand UO_363 (O_363,N_23424,N_23569);
or UO_364 (O_364,N_21503,N_21334);
or UO_365 (O_365,N_21806,N_22169);
nand UO_366 (O_366,N_23612,N_22682);
nor UO_367 (O_367,N_20472,N_21786);
and UO_368 (O_368,N_21311,N_23563);
nor UO_369 (O_369,N_22572,N_20996);
or UO_370 (O_370,N_20881,N_21319);
or UO_371 (O_371,N_20794,N_22046);
and UO_372 (O_372,N_24017,N_23158);
nor UO_373 (O_373,N_23086,N_20899);
xnor UO_374 (O_374,N_20076,N_24195);
or UO_375 (O_375,N_21270,N_24887);
and UO_376 (O_376,N_21618,N_22064);
xor UO_377 (O_377,N_24092,N_22894);
and UO_378 (O_378,N_24919,N_22422);
xor UO_379 (O_379,N_20518,N_20631);
and UO_380 (O_380,N_24833,N_20036);
or UO_381 (O_381,N_24932,N_20389);
and UO_382 (O_382,N_21597,N_23767);
xnor UO_383 (O_383,N_23626,N_20156);
nand UO_384 (O_384,N_24086,N_24774);
or UO_385 (O_385,N_23479,N_21509);
or UO_386 (O_386,N_22448,N_20139);
or UO_387 (O_387,N_21619,N_20462);
and UO_388 (O_388,N_23625,N_23786);
and UO_389 (O_389,N_24943,N_22878);
or UO_390 (O_390,N_20626,N_20377);
nor UO_391 (O_391,N_24589,N_21841);
nor UO_392 (O_392,N_20197,N_23885);
or UO_393 (O_393,N_23895,N_23688);
xnor UO_394 (O_394,N_23004,N_24739);
nand UO_395 (O_395,N_22373,N_23579);
nor UO_396 (O_396,N_23224,N_20319);
nor UO_397 (O_397,N_20652,N_24875);
xor UO_398 (O_398,N_21732,N_20070);
nor UO_399 (O_399,N_20630,N_21380);
nand UO_400 (O_400,N_24982,N_21206);
xor UO_401 (O_401,N_23334,N_23858);
or UO_402 (O_402,N_22381,N_22362);
or UO_403 (O_403,N_22153,N_24587);
or UO_404 (O_404,N_24786,N_24556);
nor UO_405 (O_405,N_23466,N_20242);
and UO_406 (O_406,N_24816,N_21932);
or UO_407 (O_407,N_24693,N_21670);
and UO_408 (O_408,N_24876,N_21442);
or UO_409 (O_409,N_21639,N_20037);
nor UO_410 (O_410,N_24665,N_24378);
nand UO_411 (O_411,N_22391,N_24526);
or UO_412 (O_412,N_21435,N_23784);
xor UO_413 (O_413,N_21514,N_20708);
nor UO_414 (O_414,N_22287,N_22551);
and UO_415 (O_415,N_23199,N_23796);
nor UO_416 (O_416,N_24605,N_21717);
or UO_417 (O_417,N_23545,N_21485);
and UO_418 (O_418,N_24456,N_24889);
nand UO_419 (O_419,N_24914,N_23481);
nand UO_420 (O_420,N_21265,N_22780);
nand UO_421 (O_421,N_24974,N_21219);
nand UO_422 (O_422,N_21874,N_23887);
and UO_423 (O_423,N_22098,N_24909);
nor UO_424 (O_424,N_20788,N_24047);
nor UO_425 (O_425,N_21948,N_23830);
or UO_426 (O_426,N_22113,N_21317);
and UO_427 (O_427,N_21613,N_24779);
nor UO_428 (O_428,N_22696,N_24139);
nand UO_429 (O_429,N_23727,N_24386);
xor UO_430 (O_430,N_24852,N_20495);
nor UO_431 (O_431,N_24728,N_22637);
or UO_432 (O_432,N_24096,N_23791);
and UO_433 (O_433,N_23720,N_20123);
and UO_434 (O_434,N_20283,N_23426);
and UO_435 (O_435,N_24458,N_22852);
nand UO_436 (O_436,N_23041,N_21513);
xnor UO_437 (O_437,N_23646,N_20808);
nor UO_438 (O_438,N_23362,N_20230);
xor UO_439 (O_439,N_24737,N_24859);
and UO_440 (O_440,N_23228,N_23446);
xnor UO_441 (O_441,N_21800,N_21269);
nor UO_442 (O_442,N_23511,N_21371);
or UO_443 (O_443,N_21710,N_22557);
and UO_444 (O_444,N_22464,N_21576);
nor UO_445 (O_445,N_24527,N_22588);
xor UO_446 (O_446,N_21205,N_23694);
or UO_447 (O_447,N_23472,N_23050);
or UO_448 (O_448,N_21348,N_22786);
and UO_449 (O_449,N_20926,N_23397);
and UO_450 (O_450,N_24689,N_24423);
nor UO_451 (O_451,N_21552,N_22471);
nor UO_452 (O_452,N_23935,N_21967);
nor UO_453 (O_453,N_23062,N_24168);
nor UO_454 (O_454,N_20732,N_21952);
nor UO_455 (O_455,N_20861,N_20521);
nand UO_456 (O_456,N_20297,N_23930);
nand UO_457 (O_457,N_21158,N_21391);
nand UO_458 (O_458,N_24294,N_20644);
nor UO_459 (O_459,N_24603,N_22607);
nor UO_460 (O_460,N_21342,N_20657);
nor UO_461 (O_461,N_20659,N_21283);
xnor UO_462 (O_462,N_24032,N_23689);
nand UO_463 (O_463,N_22979,N_21707);
nand UO_464 (O_464,N_24905,N_20263);
nand UO_465 (O_465,N_20606,N_22781);
or UO_466 (O_466,N_20974,N_20114);
xnor UO_467 (O_467,N_24544,N_23222);
nor UO_468 (O_468,N_21773,N_21051);
xor UO_469 (O_469,N_20870,N_20084);
and UO_470 (O_470,N_22762,N_24505);
and UO_471 (O_471,N_24892,N_20272);
or UO_472 (O_472,N_23204,N_24757);
nand UO_473 (O_473,N_24743,N_21731);
or UO_474 (O_474,N_23624,N_24778);
or UO_475 (O_475,N_22073,N_23326);
and UO_476 (O_476,N_23358,N_21154);
nand UO_477 (O_477,N_24381,N_20610);
nor UO_478 (O_478,N_22358,N_23703);
nor UO_479 (O_479,N_21353,N_23923);
or UO_480 (O_480,N_23058,N_20622);
nor UO_481 (O_481,N_21843,N_22494);
nand UO_482 (O_482,N_22186,N_23040);
nor UO_483 (O_483,N_22512,N_21900);
xnor UO_484 (O_484,N_24879,N_23963);
or UO_485 (O_485,N_20033,N_20545);
xor UO_486 (O_486,N_21240,N_24837);
or UO_487 (O_487,N_21854,N_23240);
xor UO_488 (O_488,N_23780,N_20769);
and UO_489 (O_489,N_22364,N_22688);
nor UO_490 (O_490,N_24924,N_22070);
xnor UO_491 (O_491,N_21582,N_23406);
and UO_492 (O_492,N_23681,N_20478);
nand UO_493 (O_493,N_21195,N_24163);
nand UO_494 (O_494,N_23191,N_24601);
nor UO_495 (O_495,N_22927,N_20165);
xnor UO_496 (O_496,N_22995,N_20562);
or UO_497 (O_497,N_24829,N_21632);
xor UO_498 (O_498,N_24077,N_21844);
and UO_499 (O_499,N_24718,N_22485);
xnor UO_500 (O_500,N_24369,N_24042);
and UO_501 (O_501,N_23915,N_22966);
nand UO_502 (O_502,N_22851,N_21014);
or UO_503 (O_503,N_21159,N_21564);
or UO_504 (O_504,N_24444,N_22834);
or UO_505 (O_505,N_22178,N_24085);
nor UO_506 (O_506,N_24383,N_22256);
nand UO_507 (O_507,N_23139,N_20396);
nor UO_508 (O_508,N_20489,N_22908);
nor UO_509 (O_509,N_21768,N_24170);
nand UO_510 (O_510,N_22753,N_23521);
nand UO_511 (O_511,N_20424,N_24259);
xnor UO_512 (O_512,N_20288,N_20739);
nor UO_513 (O_513,N_24618,N_23940);
nor UO_514 (O_514,N_22802,N_23848);
xor UO_515 (O_515,N_22569,N_24127);
nand UO_516 (O_516,N_21498,N_23731);
nor UO_517 (O_517,N_23819,N_22022);
or UO_518 (O_518,N_23889,N_21289);
and UO_519 (O_519,N_24331,N_22842);
or UO_520 (O_520,N_21709,N_23574);
nand UO_521 (O_521,N_20755,N_24827);
or UO_522 (O_522,N_22929,N_20604);
nor UO_523 (O_523,N_23205,N_23182);
nand UO_524 (O_524,N_21484,N_22394);
nor UO_525 (O_525,N_22775,N_22412);
nor UO_526 (O_526,N_21925,N_22613);
and UO_527 (O_527,N_24364,N_21150);
or UO_528 (O_528,N_22437,N_24933);
and UO_529 (O_529,N_22890,N_21460);
nand UO_530 (O_530,N_21002,N_20185);
nor UO_531 (O_531,N_24619,N_20355);
or UO_532 (O_532,N_21563,N_21215);
xnor UO_533 (O_533,N_21989,N_20947);
and UO_534 (O_534,N_23711,N_24682);
and UO_535 (O_535,N_24482,N_24290);
nand UO_536 (O_536,N_20441,N_21796);
nand UO_537 (O_537,N_24615,N_20274);
xnor UO_538 (O_538,N_22863,N_20239);
nor UO_539 (O_539,N_23833,N_21823);
xnor UO_540 (O_540,N_24984,N_20296);
nand UO_541 (O_541,N_23036,N_23312);
nand UO_542 (O_542,N_23340,N_22991);
nand UO_543 (O_543,N_22283,N_24908);
nor UO_544 (O_544,N_22506,N_20674);
or UO_545 (O_545,N_22482,N_20902);
xor UO_546 (O_546,N_24841,N_20864);
nor UO_547 (O_547,N_22487,N_21698);
nor UO_548 (O_548,N_24897,N_24575);
nand UO_549 (O_549,N_23775,N_21372);
nor UO_550 (O_550,N_21668,N_21224);
nand UO_551 (O_551,N_21266,N_23273);
and UO_552 (O_552,N_24636,N_22848);
xor UO_553 (O_553,N_22148,N_22814);
and UO_554 (O_554,N_23237,N_22643);
xnor UO_555 (O_555,N_21726,N_24057);
xor UO_556 (O_556,N_24624,N_22338);
nor UO_557 (O_557,N_20480,N_22881);
xnor UO_558 (O_558,N_24538,N_21441);
or UO_559 (O_559,N_21359,N_22236);
xnor UO_560 (O_560,N_20880,N_20829);
or UO_561 (O_561,N_21822,N_22539);
xnor UO_562 (O_562,N_23235,N_21036);
nor UO_563 (O_563,N_22204,N_22879);
nor UO_564 (O_564,N_20650,N_20062);
xor UO_565 (O_565,N_22475,N_23459);
and UO_566 (O_566,N_20032,N_23672);
nand UO_567 (O_567,N_24899,N_24554);
nand UO_568 (O_568,N_24795,N_24600);
or UO_569 (O_569,N_22337,N_23214);
nand UO_570 (O_570,N_21558,N_21876);
xnor UO_571 (O_571,N_23677,N_23875);
nand UO_572 (O_572,N_24225,N_23750);
and UO_573 (O_573,N_22681,N_23281);
nor UO_574 (O_574,N_23486,N_22171);
nand UO_575 (O_575,N_24842,N_23912);
or UO_576 (O_576,N_21136,N_21749);
or UO_577 (O_577,N_21284,N_22911);
nor UO_578 (O_578,N_20147,N_24635);
xor UO_579 (O_579,N_20721,N_21197);
or UO_580 (O_580,N_24373,N_20107);
or UO_581 (O_581,N_20307,N_22841);
nand UO_582 (O_582,N_20254,N_22002);
nor UO_583 (O_583,N_22197,N_23239);
nand UO_584 (O_584,N_20661,N_21217);
or UO_585 (O_585,N_21849,N_21782);
nand UO_586 (O_586,N_23827,N_23367);
nor UO_587 (O_587,N_20425,N_23861);
nor UO_588 (O_588,N_21899,N_23480);
and UO_589 (O_589,N_23552,N_20116);
xor UO_590 (O_590,N_24229,N_21037);
xor UO_591 (O_591,N_21124,N_23793);
nor UO_592 (O_592,N_24247,N_23168);
and UO_593 (O_593,N_24028,N_24993);
or UO_594 (O_594,N_23166,N_23322);
nand UO_595 (O_595,N_20874,N_20964);
or UO_596 (O_596,N_23135,N_20726);
or UO_597 (O_597,N_20271,N_23361);
or UO_598 (O_598,N_21292,N_23828);
xor UO_599 (O_599,N_24419,N_21346);
xor UO_600 (O_600,N_23453,N_22521);
xor UO_601 (O_601,N_21022,N_23285);
nor UO_602 (O_602,N_24203,N_20569);
nor UO_603 (O_603,N_24477,N_21511);
nand UO_604 (O_604,N_20738,N_24633);
xnor UO_605 (O_605,N_23212,N_24507);
and UO_606 (O_606,N_24375,N_21559);
or UO_607 (O_607,N_21274,N_23238);
nor UO_608 (O_608,N_22885,N_21994);
nor UO_609 (O_609,N_23587,N_20765);
nand UO_610 (O_610,N_24305,N_20537);
xnor UO_611 (O_611,N_20277,N_22666);
nor UO_612 (O_612,N_23291,N_20226);
nand UO_613 (O_613,N_20994,N_24427);
nand UO_614 (O_614,N_24061,N_20632);
nor UO_615 (O_615,N_23215,N_23603);
nor UO_616 (O_616,N_24056,N_22714);
nor UO_617 (O_617,N_20727,N_20333);
nor UO_618 (O_618,N_23047,N_23485);
and UO_619 (O_619,N_24404,N_20935);
xor UO_620 (O_620,N_20499,N_21331);
and UO_621 (O_621,N_24314,N_23070);
xor UO_622 (O_622,N_24184,N_20691);
nand UO_623 (O_623,N_24830,N_21923);
nand UO_624 (O_624,N_23742,N_21664);
nor UO_625 (O_625,N_24260,N_21627);
or UO_626 (O_626,N_22158,N_21189);
and UO_627 (O_627,N_20806,N_23370);
nand UO_628 (O_628,N_22291,N_22459);
and UO_629 (O_629,N_22205,N_20485);
or UO_630 (O_630,N_20963,N_21752);
nor UO_631 (O_631,N_23059,N_20713);
nor UO_632 (O_632,N_23498,N_20787);
or UO_633 (O_633,N_23497,N_22223);
nor UO_634 (O_634,N_21596,N_20725);
and UO_635 (O_635,N_23886,N_22800);
and UO_636 (O_636,N_24559,N_20437);
nor UO_637 (O_637,N_21413,N_20851);
xor UO_638 (O_638,N_21581,N_21908);
nand UO_639 (O_639,N_22972,N_23910);
nand UO_640 (O_640,N_21369,N_20640);
xnor UO_641 (O_641,N_24724,N_24019);
nor UO_642 (O_642,N_20224,N_22377);
nor UO_643 (O_643,N_23798,N_22632);
xnor UO_644 (O_644,N_22623,N_23329);
xnor UO_645 (O_645,N_24472,N_23864);
nor UO_646 (O_646,N_23414,N_20169);
nor UO_647 (O_647,N_23507,N_24491);
nor UO_648 (O_648,N_21759,N_21041);
or UO_649 (O_649,N_21833,N_21983);
or UO_650 (O_650,N_21009,N_24691);
nand UO_651 (O_651,N_20075,N_22913);
nor UO_652 (O_652,N_23553,N_20834);
xor UO_653 (O_653,N_22695,N_24320);
nor UO_654 (O_654,N_23960,N_23371);
and UO_655 (O_655,N_22791,N_23657);
xnor UO_656 (O_656,N_21728,N_23491);
nor UO_657 (O_657,N_20779,N_20536);
nand UO_658 (O_658,N_23457,N_22912);
and UO_659 (O_659,N_22095,N_21448);
xor UO_660 (O_660,N_22700,N_22586);
nand UO_661 (O_661,N_24785,N_22598);
or UO_662 (O_662,N_20965,N_24540);
xor UO_663 (O_663,N_23639,N_24418);
nor UO_664 (O_664,N_22054,N_21263);
xor UO_665 (O_665,N_22578,N_21851);
xor UO_666 (O_666,N_22922,N_21163);
or UO_667 (O_667,N_20587,N_21196);
nor UO_668 (O_668,N_23825,N_22145);
or UO_669 (O_669,N_23402,N_21678);
and UO_670 (O_670,N_23413,N_21933);
or UO_671 (O_671,N_20352,N_24964);
and UO_672 (O_672,N_22719,N_23922);
or UO_673 (O_673,N_22473,N_21332);
nor UO_674 (O_674,N_22635,N_21601);
or UO_675 (O_675,N_21522,N_21866);
or UO_676 (O_676,N_20621,N_21427);
nor UO_677 (O_677,N_22143,N_22934);
nor UO_678 (O_678,N_24613,N_22005);
and UO_679 (O_679,N_24346,N_24348);
or UO_680 (O_680,N_20395,N_21202);
nand UO_681 (O_681,N_24790,N_24697);
and UO_682 (O_682,N_23697,N_24131);
or UO_683 (O_683,N_21273,N_22507);
or UO_684 (O_684,N_24772,N_24194);
nand UO_685 (O_685,N_21529,N_22658);
or UO_686 (O_686,N_20519,N_24787);
nand UO_687 (O_687,N_24254,N_23546);
or UO_688 (O_688,N_20467,N_22668);
xor UO_689 (O_689,N_23351,N_24284);
xor UO_690 (O_690,N_23066,N_23931);
and UO_691 (O_691,N_24073,N_21955);
xnor UO_692 (O_692,N_24877,N_20421);
and UO_693 (O_693,N_24461,N_24564);
xor UO_694 (O_694,N_20180,N_24275);
xor UO_695 (O_695,N_22917,N_23637);
nor UO_696 (O_696,N_22195,N_22707);
and UO_697 (O_697,N_24481,N_20413);
or UO_698 (O_698,N_20534,N_23645);
nand UO_699 (O_699,N_24873,N_24989);
nor UO_700 (O_700,N_24819,N_23840);
nand UO_701 (O_701,N_21663,N_21040);
or UO_702 (O_702,N_24685,N_22035);
nor UO_703 (O_703,N_21109,N_20287);
nor UO_704 (O_704,N_20795,N_21575);
nor UO_705 (O_705,N_21354,N_24453);
and UO_706 (O_706,N_23254,N_20245);
and UO_707 (O_707,N_24024,N_20673);
or UO_708 (O_708,N_20222,N_23022);
nand UO_709 (O_709,N_22537,N_21761);
nor UO_710 (O_710,N_23866,N_23244);
nor UO_711 (O_711,N_20833,N_23278);
nand UO_712 (O_712,N_23816,N_23410);
nor UO_713 (O_713,N_22880,N_20887);
xnor UO_714 (O_714,N_22206,N_23661);
or UO_715 (O_715,N_20756,N_24717);
xnor UO_716 (O_716,N_21044,N_21703);
nor UO_717 (O_717,N_24972,N_24321);
and UO_718 (O_718,N_20207,N_24565);
xor UO_719 (O_719,N_20505,N_24470);
nor UO_720 (O_720,N_24629,N_23264);
and UO_721 (O_721,N_20056,N_23690);
nor UO_722 (O_722,N_20954,N_24561);
or UO_723 (O_723,N_21126,N_23287);
or UO_724 (O_724,N_22545,N_20825);
and UO_725 (O_725,N_21423,N_24863);
nor UO_726 (O_726,N_23852,N_23372);
and UO_727 (O_727,N_23104,N_20557);
xnor UO_728 (O_728,N_21977,N_23977);
or UO_729 (O_729,N_22705,N_21419);
and UO_730 (O_730,N_20432,N_22463);
and UO_731 (O_731,N_21973,N_21580);
and UO_732 (O_732,N_24120,N_22326);
xnor UO_733 (O_733,N_23728,N_23763);
and UO_734 (O_734,N_20993,N_22368);
or UO_735 (O_735,N_23318,N_24806);
nand UO_736 (O_736,N_21415,N_21465);
nor UO_737 (O_737,N_23856,N_24632);
xor UO_738 (O_738,N_24948,N_23407);
xnor UO_739 (O_739,N_21104,N_21381);
or UO_740 (O_740,N_22756,N_23760);
and UO_741 (O_741,N_21729,N_21742);
or UO_742 (O_742,N_20920,N_22730);
nor UO_743 (O_743,N_24343,N_23467);
nand UO_744 (O_744,N_20771,N_23510);
nand UO_745 (O_745,N_22138,N_23478);
xnor UO_746 (O_746,N_23213,N_22133);
nand UO_747 (O_747,N_24034,N_24865);
and UO_748 (O_748,N_23487,N_22675);
and UO_749 (O_749,N_21638,N_21545);
nor UO_750 (O_750,N_23722,N_22989);
and UO_751 (O_751,N_20188,N_24504);
nand UO_752 (O_752,N_23927,N_22277);
xor UO_753 (O_753,N_22964,N_22187);
nand UO_754 (O_754,N_20928,N_23759);
and UO_755 (O_755,N_21937,N_21607);
or UO_756 (O_756,N_22920,N_23428);
and UO_757 (O_757,N_20999,N_20280);
or UO_758 (O_758,N_21338,N_24476);
and UO_759 (O_759,N_22264,N_20932);
or UO_760 (O_760,N_22674,N_21157);
or UO_761 (O_761,N_23762,N_22502);
nor UO_762 (O_762,N_24977,N_21487);
nand UO_763 (O_763,N_22717,N_23562);
and UO_764 (O_764,N_21515,N_20358);
or UO_765 (O_765,N_24459,N_23107);
nand UO_766 (O_766,N_23314,N_21544);
nand UO_767 (O_767,N_21502,N_22698);
xnor UO_768 (O_768,N_20624,N_22386);
xnor UO_769 (O_769,N_21405,N_21543);
xor UO_770 (O_770,N_23053,N_24738);
and UO_771 (O_771,N_23644,N_20790);
or UO_772 (O_772,N_21072,N_20305);
or UO_773 (O_773,N_22532,N_24706);
or UO_774 (O_774,N_22263,N_20529);
or UO_775 (O_775,N_22855,N_21056);
nand UO_776 (O_776,N_24606,N_23025);
or UO_777 (O_777,N_24578,N_22706);
nand UO_778 (O_778,N_21102,N_23376);
xnor UO_779 (O_779,N_21131,N_24243);
xor UO_780 (O_780,N_22818,N_23812);
or UO_781 (O_781,N_22480,N_24224);
xnor UO_782 (O_782,N_21211,N_21167);
xor UO_783 (O_783,N_21107,N_21042);
nor UO_784 (O_784,N_20404,N_24199);
or UO_785 (O_785,N_24368,N_22749);
nor UO_786 (O_786,N_23943,N_23389);
and UO_787 (O_787,N_24118,N_21885);
or UO_788 (O_788,N_22813,N_24570);
and UO_789 (O_789,N_22782,N_23835);
nand UO_790 (O_790,N_20729,N_21606);
xnor UO_791 (O_791,N_24000,N_22571);
xnor UO_792 (O_792,N_23949,N_21013);
nand UO_793 (O_793,N_22530,N_23749);
and UO_794 (O_794,N_20796,N_21763);
nand UO_795 (O_795,N_21810,N_24916);
and UO_796 (O_796,N_20414,N_22611);
xnor UO_797 (O_797,N_21602,N_23172);
and UO_798 (O_798,N_24983,N_21496);
nand UO_799 (O_799,N_23043,N_24740);
xor UO_800 (O_800,N_22273,N_21242);
nor UO_801 (O_801,N_22470,N_23594);
nand UO_802 (O_802,N_22086,N_21996);
xor UO_803 (O_803,N_24191,N_24181);
xnor UO_804 (O_804,N_24999,N_20015);
nor UO_805 (O_805,N_21999,N_21975);
or UO_806 (O_806,N_23387,N_23972);
or UO_807 (O_807,N_23869,N_22947);
and UO_808 (O_808,N_20651,N_21821);
or UO_809 (O_809,N_24172,N_24137);
nand UO_810 (O_810,N_20183,N_22072);
nand UO_811 (O_811,N_23907,N_23184);
nor UO_812 (O_812,N_24666,N_21068);
nand UO_813 (O_813,N_23522,N_23342);
nor UO_814 (O_814,N_23452,N_20985);
and UO_815 (O_815,N_21886,N_20843);
nor UO_816 (O_816,N_22060,N_22403);
nand UO_817 (O_817,N_24064,N_20174);
xor UO_818 (O_818,N_23685,N_24167);
nor UO_819 (O_819,N_20453,N_20686);
or UO_820 (O_820,N_24471,N_22102);
xnor UO_821 (O_821,N_20306,N_22624);
nand UO_822 (O_822,N_21944,N_23283);
xor UO_823 (O_823,N_23320,N_24901);
nand UO_824 (O_824,N_22641,N_22916);
xnor UO_825 (O_825,N_20048,N_23560);
or UO_826 (O_826,N_20735,N_23415);
nand UO_827 (O_827,N_21978,N_23932);
xnor UO_828 (O_828,N_23198,N_22150);
nand UO_829 (O_829,N_24049,N_20371);
nand UO_830 (O_830,N_24936,N_20636);
xor UO_831 (O_831,N_22948,N_23953);
nand UO_832 (O_832,N_23473,N_24864);
and UO_833 (O_833,N_22980,N_23299);
nand UO_834 (O_834,N_21976,N_23167);
and UO_835 (O_835,N_24711,N_20092);
and UO_836 (O_836,N_22836,N_20321);
nor UO_837 (O_837,N_20246,N_20763);
xor UO_838 (O_838,N_23097,N_24760);
or UO_839 (O_839,N_22441,N_20791);
xnor UO_840 (O_840,N_22734,N_23419);
nor UO_841 (O_841,N_20193,N_21414);
nand UO_842 (O_842,N_20104,N_23669);
and UO_843 (O_843,N_21437,N_20689);
nand UO_844 (O_844,N_23454,N_22068);
or UO_845 (O_845,N_21349,N_24813);
or UO_846 (O_846,N_22973,N_24068);
or UO_847 (O_847,N_22645,N_24179);
nand UO_848 (O_848,N_20975,N_23438);
or UO_849 (O_849,N_22425,N_22713);
nor UO_850 (O_850,N_21984,N_23606);
or UO_851 (O_851,N_23113,N_21199);
and UO_852 (O_852,N_23523,N_20816);
nand UO_853 (O_853,N_21340,N_24265);
nor UO_854 (O_854,N_21469,N_21591);
nor UO_855 (O_855,N_20801,N_22847);
nor UO_856 (O_856,N_20594,N_20167);
nor UO_857 (O_857,N_24021,N_24720);
and UO_858 (O_858,N_21739,N_23948);
nand UO_859 (O_859,N_24641,N_21471);
nor UO_860 (O_860,N_21461,N_20215);
and UO_861 (O_861,N_20595,N_20433);
nand UO_862 (O_862,N_20119,N_21969);
nor UO_863 (O_863,N_23327,N_20646);
nand UO_864 (O_864,N_22640,N_20511);
and UO_865 (O_865,N_21004,N_21918);
or UO_866 (O_866,N_22599,N_24088);
and UO_867 (O_867,N_22687,N_20758);
nand UO_868 (O_868,N_24013,N_24623);
nor UO_869 (O_869,N_24904,N_22156);
nor UO_870 (O_870,N_23551,N_22351);
or UO_871 (O_871,N_21661,N_23286);
or UO_872 (O_872,N_22898,N_22347);
nand UO_873 (O_873,N_20384,N_24945);
xnor UO_874 (O_874,N_22057,N_24242);
nand UO_875 (O_875,N_24817,N_23078);
or UO_876 (O_876,N_20279,N_24574);
xor UO_877 (O_877,N_22715,N_24736);
xor UO_878 (O_878,N_22366,N_23449);
or UO_879 (O_879,N_20951,N_23753);
and UO_880 (O_880,N_20343,N_20693);
and UO_881 (O_881,N_24413,N_22016);
nor UO_882 (O_882,N_21088,N_23400);
nor UO_883 (O_883,N_20842,N_23802);
nand UO_884 (O_884,N_24271,N_22298);
and UO_885 (O_885,N_23169,N_22826);
xnor UO_886 (O_886,N_20720,N_24258);
xnor UO_887 (O_887,N_24756,N_20301);
nand UO_888 (O_888,N_23092,N_24072);
and UO_889 (O_889,N_23559,N_22628);
xnor UO_890 (O_890,N_21616,N_24022);
xnor UO_891 (O_891,N_24487,N_21753);
and UO_892 (O_892,N_22812,N_22009);
nor UO_893 (O_893,N_23422,N_20885);
and UO_894 (O_894,N_21320,N_23385);
nand UO_895 (O_895,N_23008,N_21847);
nand UO_896 (O_896,N_22380,N_24958);
nand UO_897 (O_897,N_22552,N_22788);
and UO_898 (O_898,N_21184,N_21620);
or UO_899 (O_899,N_23265,N_20488);
or UO_900 (O_900,N_23557,N_20866);
nand UO_901 (O_901,N_24550,N_22050);
or UO_902 (O_902,N_23747,N_21394);
or UO_903 (O_903,N_22627,N_20540);
xor UO_904 (O_904,N_20807,N_23531);
nor UO_905 (O_905,N_20429,N_24475);
or UO_906 (O_906,N_21451,N_24637);
and UO_907 (O_907,N_21897,N_22456);
nor UO_908 (O_908,N_23305,N_23232);
nand UO_909 (O_909,N_20460,N_24912);
or UO_910 (O_910,N_24283,N_24555);
nand UO_911 (O_911,N_23259,N_22669);
nand UO_912 (O_912,N_22127,N_22691);
or UO_913 (O_913,N_23655,N_21836);
and UO_914 (O_914,N_20359,N_24518);
or UO_915 (O_915,N_22481,N_21433);
and UO_916 (O_916,N_20832,N_22939);
xor UO_917 (O_917,N_20871,N_23016);
nor UO_918 (O_918,N_22994,N_20209);
or UO_919 (O_919,N_21152,N_21142);
and UO_920 (O_920,N_23344,N_23460);
nor UO_921 (O_921,N_20946,N_24399);
nor UO_922 (O_922,N_23516,N_22886);
and UO_923 (O_923,N_23013,N_22772);
nor UO_924 (O_924,N_20716,N_20574);
nor UO_925 (O_925,N_23174,N_21416);
xnor UO_926 (O_926,N_21765,N_21328);
nand UO_927 (O_927,N_23505,N_20616);
nor UO_928 (O_928,N_21344,N_24285);
nor UO_929 (O_929,N_20375,N_22738);
xnor UO_930 (O_930,N_24183,N_22579);
or UO_931 (O_931,N_21468,N_22335);
xor UO_932 (O_932,N_21430,N_21006);
nand UO_933 (O_933,N_20140,N_21917);
nor UO_934 (O_934,N_24069,N_21491);
or UO_935 (O_935,N_23764,N_21170);
or UO_936 (O_936,N_20398,N_20612);
nor UO_937 (O_937,N_20372,N_21122);
xor UO_938 (O_938,N_23143,N_23508);
xor UO_939 (O_939,N_22135,N_24900);
xnor UO_940 (O_940,N_21176,N_20663);
nand UO_941 (O_941,N_21490,N_20105);
or UO_942 (O_942,N_23355,N_24256);
xnor UO_943 (O_943,N_23933,N_24588);
and UO_944 (O_944,N_23292,N_24661);
or UO_945 (O_945,N_23444,N_20006);
nand UO_946 (O_946,N_23216,N_22967);
nor UO_947 (O_947,N_24667,N_22794);
nor UO_948 (O_948,N_23122,N_20731);
xor UO_949 (O_949,N_24815,N_23518);
xnor UO_950 (O_950,N_23729,N_21832);
nor UO_951 (O_951,N_24512,N_20448);
and UO_952 (O_952,N_20957,N_22014);
nand UO_953 (O_953,N_23918,N_22279);
nand UO_954 (O_954,N_22974,N_21425);
and UO_955 (O_955,N_23079,N_20886);
xor UO_956 (O_956,N_24354,N_20194);
nor UO_957 (O_957,N_21103,N_23821);
nor UO_958 (O_958,N_22446,N_23310);
xor UO_959 (O_959,N_23384,N_20409);
nor UO_960 (O_960,N_23311,N_23462);
xor UO_961 (O_961,N_21659,N_20767);
nand UO_962 (O_962,N_21845,N_24315);
or UO_963 (O_963,N_21440,N_23211);
or UO_964 (O_964,N_22825,N_21699);
xor UO_965 (O_965,N_23356,N_23514);
xor UO_966 (O_966,N_24788,N_23616);
and UO_967 (O_967,N_24687,N_22790);
nor UO_968 (O_968,N_20528,N_23493);
or UO_969 (O_969,N_21100,N_20527);
nor UO_970 (O_970,N_24804,N_22653);
and UO_971 (O_971,N_23297,N_24824);
or UO_972 (O_972,N_22716,N_22923);
nor UO_973 (O_973,N_20014,N_23464);
or UO_974 (O_974,N_21890,N_23187);
xor UO_975 (O_975,N_20385,N_23801);
or UO_976 (O_976,N_24910,N_21883);
and UO_977 (O_977,N_22163,N_20293);
nor UO_978 (O_978,N_23882,N_22213);
xnor UO_979 (O_979,N_20085,N_23952);
nand UO_980 (O_980,N_20261,N_20058);
nand UO_981 (O_981,N_20490,N_24925);
nor UO_982 (O_982,N_24104,N_24703);
xnor UO_983 (O_983,N_22117,N_24549);
and UO_984 (O_984,N_23335,N_24834);
nand UO_985 (O_985,N_24421,N_20812);
nand UO_986 (O_986,N_22528,N_21226);
or UO_987 (O_987,N_20098,N_24942);
nand UO_988 (O_988,N_22877,N_22793);
nor UO_989 (O_989,N_24144,N_22209);
xnor UO_990 (O_990,N_21837,N_23306);
nor UO_991 (O_991,N_22977,N_22229);
or UO_992 (O_992,N_24385,N_20666);
or UO_993 (O_993,N_24750,N_22184);
and UO_994 (O_994,N_21755,N_21858);
and UO_995 (O_995,N_22876,N_21258);
and UO_996 (O_996,N_23583,N_23841);
xnor UO_997 (O_997,N_22806,N_23726);
nand UO_998 (O_998,N_20559,N_22657);
xor UO_999 (O_999,N_21654,N_20134);
or UO_1000 (O_1000,N_21130,N_23580);
nand UO_1001 (O_1001,N_20588,N_20258);
or UO_1002 (O_1002,N_22751,N_24440);
and UO_1003 (O_1003,N_22423,N_21409);
nand UO_1004 (O_1004,N_23396,N_23202);
xnor UO_1005 (O_1005,N_21743,N_20766);
or UO_1006 (O_1006,N_21825,N_20057);
nand UO_1007 (O_1007,N_21713,N_21312);
nand UO_1008 (O_1008,N_22661,N_23350);
and UO_1009 (O_1009,N_24312,N_20038);
xnor UO_1010 (O_1010,N_20071,N_24304);
nor UO_1011 (O_1011,N_20143,N_21839);
or UO_1012 (O_1012,N_22950,N_20923);
or UO_1013 (O_1013,N_22288,N_21780);
nand UO_1014 (O_1014,N_20892,N_24968);
and UO_1015 (O_1015,N_20041,N_22817);
nand UO_1016 (O_1016,N_24425,N_24447);
xnor UO_1017 (O_1017,N_21389,N_23469);
nand UO_1018 (O_1018,N_24204,N_22284);
nand UO_1019 (O_1019,N_23201,N_22239);
or UO_1020 (O_1020,N_20407,N_22003);
or UO_1021 (O_1021,N_24268,N_22686);
and UO_1022 (O_1022,N_21443,N_21396);
nand UO_1023 (O_1023,N_20148,N_23068);
nor UO_1024 (O_1024,N_24249,N_21986);
or UO_1025 (O_1025,N_23651,N_24384);
xnor UO_1026 (O_1026,N_20420,N_22957);
xor UO_1027 (O_1027,N_20029,N_21343);
xor UO_1028 (O_1028,N_24663,N_21190);
nand UO_1029 (O_1029,N_21192,N_24874);
nor UO_1030 (O_1030,N_24098,N_21390);
xnor UO_1031 (O_1031,N_21828,N_21305);
or UO_1032 (O_1032,N_23589,N_22720);
and UO_1033 (O_1033,N_22978,N_21123);
or UO_1034 (O_1034,N_22811,N_24907);
nand UO_1035 (O_1035,N_20589,N_20516);
xnor UO_1036 (O_1036,N_21376,N_20544);
and UO_1037 (O_1037,N_24318,N_24434);
or UO_1038 (O_1038,N_23973,N_21993);
xnor UO_1039 (O_1039,N_22389,N_22692);
nor UO_1040 (O_1040,N_20030,N_21799);
and UO_1041 (O_1041,N_24962,N_20186);
and UO_1042 (O_1042,N_22612,N_22177);
and UO_1043 (O_1043,N_20838,N_21852);
nand UO_1044 (O_1044,N_24569,N_23509);
or UO_1045 (O_1045,N_23321,N_22140);
nand UO_1046 (O_1046,N_21578,N_22872);
or UO_1047 (O_1047,N_22390,N_24792);
or UO_1048 (O_1048,N_23451,N_21571);
nand UO_1049 (O_1049,N_20552,N_23192);
nor UO_1050 (O_1050,N_22208,N_22220);
nor UO_1051 (O_1051,N_22013,N_22469);
or UO_1052 (O_1052,N_23787,N_23756);
or UO_1053 (O_1053,N_21856,N_20699);
or UO_1054 (O_1054,N_21865,N_23706);
nand UO_1055 (O_1055,N_20524,N_20200);
nand UO_1056 (O_1056,N_21669,N_20464);
or UO_1057 (O_1057,N_24921,N_24182);
nand UO_1058 (O_1058,N_21809,N_22428);
or UO_1059 (O_1059,N_22166,N_24054);
nand UO_1060 (O_1060,N_21232,N_24648);
xnor UO_1061 (O_1061,N_23411,N_24429);
nand UO_1062 (O_1062,N_21966,N_23275);
nor UO_1063 (O_1063,N_24679,N_23770);
or UO_1064 (O_1064,N_22067,N_21287);
xnor UO_1065 (O_1065,N_21506,N_21397);
or UO_1066 (O_1066,N_23824,N_21313);
nand UO_1067 (O_1067,N_21120,N_21921);
nand UO_1068 (O_1068,N_23618,N_22779);
xor UO_1069 (O_1069,N_22257,N_21095);
and UO_1070 (O_1070,N_22436,N_24380);
xnor UO_1071 (O_1071,N_22352,N_20335);
nand UO_1072 (O_1072,N_20762,N_23035);
nand UO_1073 (O_1073,N_21622,N_23072);
or UO_1074 (O_1074,N_20044,N_23121);
and UO_1075 (O_1075,N_24134,N_24417);
and UO_1076 (O_1076,N_23146,N_23723);
xnor UO_1077 (O_1077,N_23573,N_21962);
or UO_1078 (O_1078,N_23593,N_24422);
and UO_1079 (O_1079,N_24981,N_22602);
and UO_1080 (O_1080,N_24906,N_22618);
xor UO_1081 (O_1081,N_20248,N_22958);
and UO_1082 (O_1082,N_24405,N_21880);
xor UO_1083 (O_1083,N_21310,N_23576);
and UO_1084 (O_1084,N_22198,N_22844);
nor UO_1085 (O_1085,N_23231,N_24678);
nor UO_1086 (O_1086,N_22226,N_24478);
nor UO_1087 (O_1087,N_24152,N_23328);
or UO_1088 (O_1088,N_24102,N_23831);
nand UO_1089 (O_1089,N_20702,N_20619);
and UO_1090 (O_1090,N_22094,N_20969);
nor UO_1091 (O_1091,N_23503,N_20872);
or UO_1092 (O_1092,N_23117,N_20596);
and UO_1093 (O_1093,N_20397,N_23316);
nand UO_1094 (O_1094,N_22575,N_21276);
and UO_1095 (O_1095,N_24449,N_24856);
nand UO_1096 (O_1096,N_24201,N_24335);
or UO_1097 (O_1097,N_24132,N_21432);
nand UO_1098 (O_1098,N_24602,N_22567);
nor UO_1099 (O_1099,N_23313,N_21636);
nand UO_1100 (O_1100,N_24770,N_23360);
or UO_1101 (O_1101,N_24050,N_22000);
or UO_1102 (O_1102,N_24484,N_24428);
nor UO_1103 (O_1103,N_24653,N_24669);
or UO_1104 (O_1104,N_22925,N_24690);
xor UO_1105 (O_1105,N_21370,N_23838);
or UO_1106 (O_1106,N_20925,N_23755);
or UO_1107 (O_1107,N_24286,N_23607);
and UO_1108 (O_1108,N_20045,N_21360);
nor UO_1109 (O_1109,N_22594,N_21164);
nor UO_1110 (O_1110,N_21050,N_23003);
nand UO_1111 (O_1111,N_24721,N_23633);
nand UO_1112 (O_1112,N_23549,N_24439);
xor UO_1113 (O_1113,N_20878,N_24651);
and UO_1114 (O_1114,N_23990,N_23744);
nand UO_1115 (O_1115,N_20144,N_24462);
nand UO_1116 (O_1116,N_22180,N_21594);
or UO_1117 (O_1117,N_22888,N_22112);
and UO_1118 (O_1118,N_21486,N_22822);
and UO_1119 (O_1119,N_21681,N_24279);
nor UO_1120 (O_1120,N_21098,N_20525);
and UO_1121 (O_1121,N_20875,N_23391);
and UO_1122 (O_1122,N_21204,N_24362);
or UO_1123 (O_1123,N_22382,N_23337);
nor UO_1124 (O_1124,N_20863,N_23475);
and UO_1125 (O_1125,N_23829,N_22248);
nor UO_1126 (O_1126,N_23030,N_24307);
and UO_1127 (O_1127,N_22619,N_21797);
or UO_1128 (O_1128,N_23758,N_24025);
nor UO_1129 (O_1129,N_23483,N_20474);
xnor UO_1130 (O_1130,N_24301,N_22804);
nor UO_1131 (O_1131,N_23103,N_20049);
xor UO_1132 (O_1132,N_24162,N_20024);
nor UO_1133 (O_1133,N_20571,N_21553);
and UO_1134 (O_1134,N_23721,N_23463);
nor UO_1135 (O_1135,N_21725,N_22891);
and UO_1136 (O_1136,N_24807,N_20745);
xor UO_1137 (O_1137,N_20584,N_20256);
nor UO_1138 (O_1138,N_21589,N_20486);
nor UO_1139 (O_1139,N_24954,N_22354);
nor UO_1140 (O_1140,N_21814,N_21058);
xor UO_1141 (O_1141,N_22342,N_21198);
nor UO_1142 (O_1142,N_22798,N_20158);
xor UO_1143 (O_1143,N_20810,N_22712);
nor UO_1144 (O_1144,N_23525,N_20260);
xnor UO_1145 (O_1145,N_20391,N_20120);
nand UO_1146 (O_1146,N_21689,N_24445);
xnor UO_1147 (O_1147,N_20054,N_20473);
and UO_1148 (O_1148,N_21792,N_22543);
and UO_1149 (O_1149,N_22281,N_24280);
or UO_1150 (O_1150,N_22596,N_22238);
and UO_1151 (O_1151,N_21577,N_23269);
and UO_1152 (O_1152,N_22484,N_24662);
xor UO_1153 (O_1153,N_23338,N_22654);
and UO_1154 (O_1154,N_21603,N_23698);
and UO_1155 (O_1155,N_22860,N_20341);
xnor UO_1156 (O_1156,N_22108,N_23568);
or UO_1157 (O_1157,N_24649,N_20168);
xnor UO_1158 (O_1158,N_22742,N_23958);
nor UO_1159 (O_1159,N_21410,N_24090);
nor UO_1160 (O_1160,N_21557,N_22316);
and UO_1161 (O_1161,N_24758,N_24616);
and UO_1162 (O_1162,N_24211,N_23164);
xor UO_1163 (O_1163,N_23157,N_21733);
xor UO_1164 (O_1164,N_20406,N_20879);
nor UO_1165 (O_1165,N_23276,N_20498);
nand UO_1166 (O_1166,N_24929,N_20741);
nand UO_1167 (O_1167,N_20368,N_21203);
nor UO_1168 (O_1168,N_22840,N_20357);
nand UO_1169 (O_1169,N_22992,N_23906);
xor UO_1170 (O_1170,N_20797,N_21793);
nand UO_1171 (O_1171,N_22548,N_23251);
nor UO_1172 (O_1172,N_24158,N_24349);
or UO_1173 (O_1173,N_22690,N_23126);
xnor UO_1174 (O_1174,N_23971,N_21052);
nor UO_1175 (O_1175,N_23081,N_22555);
nand UO_1176 (O_1176,N_23331,N_20012);
or UO_1177 (O_1177,N_21262,N_23888);
or UO_1178 (O_1178,N_21133,N_22181);
nor UO_1179 (O_1179,N_21677,N_22998);
xor UO_1180 (O_1180,N_20447,N_21019);
or UO_1181 (O_1181,N_20517,N_21701);
nor UO_1182 (O_1182,N_20502,N_23302);
nor UO_1183 (O_1183,N_22361,N_24723);
or UO_1184 (O_1184,N_23439,N_20653);
nor UO_1185 (O_1185,N_24735,N_24825);
xnor UO_1186 (O_1186,N_21525,N_22685);
xor UO_1187 (O_1187,N_24140,N_21082);
or UO_1188 (O_1188,N_20635,N_24410);
xor UO_1189 (O_1189,N_23526,N_21504);
nor UO_1190 (O_1190,N_24148,N_20937);
nand UO_1191 (O_1191,N_21767,N_20649);
xnor UO_1192 (O_1192,N_22387,N_21178);
nand UO_1193 (O_1193,N_21302,N_22438);
or UO_1194 (O_1194,N_23585,N_22488);
and UO_1195 (O_1195,N_21061,N_23090);
and UO_1196 (O_1196,N_20122,N_24125);
nand UO_1197 (O_1197,N_23874,N_20465);
and UO_1198 (O_1198,N_22905,N_20730);
or UO_1199 (O_1199,N_21766,N_20322);
nor UO_1200 (O_1200,N_22642,N_23368);
xnor UO_1201 (O_1201,N_24281,N_20090);
xnor UO_1202 (O_1202,N_24686,N_23577);
or UO_1203 (O_1203,N_21241,N_21456);
or UO_1204 (O_1204,N_21075,N_20028);
or UO_1205 (O_1205,N_21392,N_21143);
and UO_1206 (O_1206,N_22617,N_22215);
and UO_1207 (O_1207,N_21679,N_23185);
xor UO_1208 (O_1208,N_20781,N_24617);
and UO_1209 (O_1209,N_22214,N_20311);
nand UO_1210 (O_1210,N_24109,N_22761);
nand UO_1211 (O_1211,N_20577,N_21495);
and UO_1212 (O_1212,N_20211,N_23983);
nand UO_1213 (O_1213,N_23642,N_21570);
nor UO_1214 (O_1214,N_20411,N_20206);
xnor UO_1215 (O_1215,N_22306,N_24659);
xnor UO_1216 (O_1216,N_21399,N_22606);
xor UO_1217 (O_1217,N_20701,N_23098);
nor UO_1218 (O_1218,N_21958,N_20563);
nor UO_1219 (O_1219,N_20751,N_24869);
nor UO_1220 (O_1220,N_23966,N_20370);
nand UO_1221 (O_1221,N_21747,N_21005);
xor UO_1222 (O_1222,N_24395,N_24071);
nand UO_1223 (O_1223,N_22864,N_22997);
or UO_1224 (O_1224,N_20658,N_20711);
xnor UO_1225 (O_1225,N_21840,N_24099);
or UO_1226 (O_1226,N_24820,N_24552);
nand UO_1227 (O_1227,N_20201,N_20856);
and UO_1228 (O_1228,N_23543,N_22741);
or UO_1229 (O_1229,N_21869,N_20728);
or UO_1230 (O_1230,N_23892,N_22370);
nor UO_1231 (O_1231,N_22625,N_23029);
nor UO_1232 (O_1232,N_24511,N_24794);
and UO_1233 (O_1233,N_21069,N_21252);
nor UO_1234 (O_1234,N_21754,N_24581);
and UO_1235 (O_1235,N_21644,N_23870);
xor UO_1236 (O_1236,N_20944,N_22029);
nand UO_1237 (O_1237,N_21209,N_23951);
xnor UO_1238 (O_1238,N_21188,N_20638);
nor UO_1239 (O_1239,N_24672,N_23105);
nand UO_1240 (O_1240,N_21035,N_20449);
nand UO_1241 (O_1241,N_20603,N_21200);
nor UO_1242 (O_1242,N_23180,N_20637);
or UO_1243 (O_1243,N_20633,N_24485);
nor UO_1244 (O_1244,N_22525,N_20737);
and UO_1245 (O_1245,N_23867,N_23965);
nand UO_1246 (O_1246,N_20079,N_20235);
xnor UO_1247 (O_1247,N_20705,N_21527);
nand UO_1248 (O_1248,N_21819,N_24045);
xor UO_1249 (O_1249,N_20164,N_21539);
nand UO_1250 (O_1250,N_21074,N_23290);
nand UO_1251 (O_1251,N_22919,N_24164);
and UO_1252 (O_1252,N_23994,N_22556);
and UO_1253 (O_1253,N_24222,N_23610);
and UO_1254 (O_1254,N_21652,N_20313);
xnor UO_1255 (O_1255,N_23925,N_21972);
or UO_1256 (O_1256,N_20942,N_22330);
or UO_1257 (O_1257,N_20958,N_24492);
nand UO_1258 (O_1258,N_24147,N_22160);
and UO_1259 (O_1259,N_20568,N_24922);
nor UO_1260 (O_1260,N_20466,N_23005);
or UO_1261 (O_1261,N_21803,N_23477);
nand UO_1262 (O_1262,N_22873,N_22334);
xnor UO_1263 (O_1263,N_22858,N_23695);
nand UO_1264 (O_1264,N_24264,N_23936);
nand UO_1265 (O_1265,N_23529,N_24340);
or UO_1266 (O_1266,N_22429,N_24202);
nor UO_1267 (O_1267,N_22119,N_23271);
nor UO_1268 (O_1268,N_22869,N_20532);
and UO_1269 (O_1269,N_24486,N_22634);
nand UO_1270 (O_1270,N_24722,N_24289);
nor UO_1271 (O_1271,N_20109,N_23893);
or UO_1272 (O_1272,N_20979,N_24712);
nor UO_1273 (O_1273,N_23236,N_20452);
nor UO_1274 (O_1274,N_21650,N_23263);
nor UO_1275 (O_1275,N_20483,N_21137);
xor UO_1276 (O_1276,N_22032,N_24696);
nor UO_1277 (O_1277,N_20744,N_23303);
nor UO_1278 (O_1278,N_22314,N_24895);
xnor UO_1279 (O_1279,N_20445,N_23789);
or UO_1280 (O_1280,N_22789,N_22999);
nand UO_1281 (O_1281,N_20468,N_21629);
or UO_1282 (O_1282,N_20647,N_22930);
nand UO_1283 (O_1283,N_22018,N_23537);
nor UO_1284 (O_1284,N_23751,N_20179);
nor UO_1285 (O_1285,N_24282,N_22805);
nor UO_1286 (O_1286,N_22671,N_23124);
or UO_1287 (O_1287,N_24210,N_22663);
or UO_1288 (O_1288,N_22479,N_22651);
nand UO_1289 (O_1289,N_24347,N_21299);
nor UO_1290 (O_1290,N_24011,N_20956);
nand UO_1291 (O_1291,N_24911,N_21193);
nand UO_1292 (O_1292,N_23363,N_21985);
or UO_1293 (O_1293,N_24654,N_20535);
or UO_1294 (O_1294,N_23420,N_20847);
and UO_1295 (O_1295,N_21626,N_21024);
nor UO_1296 (O_1296,N_20317,N_23154);
nor UO_1297 (O_1297,N_21223,N_24391);
nor UO_1298 (O_1298,N_20401,N_22356);
xnor UO_1299 (O_1299,N_21794,N_23845);
xnor UO_1300 (O_1300,N_23519,N_24111);
nor UO_1301 (O_1301,N_23561,N_21904);
and UO_1302 (O_1302,N_23019,N_20223);
xor UO_1303 (O_1303,N_22305,N_24177);
nor UO_1304 (O_1304,N_23482,N_22903);
xor UO_1305 (O_1305,N_20798,N_23837);
nand UO_1306 (O_1306,N_20696,N_24884);
nand UO_1307 (O_1307,N_23783,N_23550);
xnor UO_1308 (O_1308,N_22518,N_21434);
and UO_1309 (O_1309,N_24359,N_23834);
or UO_1310 (O_1310,N_20648,N_20232);
and UO_1311 (O_1311,N_22074,N_21171);
or UO_1312 (O_1312,N_20268,N_23392);
xor UO_1313 (O_1313,N_20709,N_23799);
nand UO_1314 (O_1314,N_24951,N_23640);
and UO_1315 (O_1315,N_21789,N_21233);
xor UO_1316 (O_1316,N_21439,N_21185);
nor UO_1317 (O_1317,N_23572,N_20050);
or UO_1318 (O_1318,N_22491,N_24235);
nor UO_1319 (O_1319,N_22740,N_20365);
nand UO_1320 (O_1320,N_24970,N_24035);
and UO_1321 (O_1321,N_22667,N_24190);
nor UO_1322 (O_1322,N_23556,N_22078);
and UO_1323 (O_1323,N_21032,N_21945);
xnor UO_1324 (O_1324,N_24344,N_22227);
xor UO_1325 (O_1325,N_21236,N_21842);
nor UO_1326 (O_1326,N_20004,N_22360);
nand UO_1327 (O_1327,N_21135,N_24135);
and UO_1328 (O_1328,N_24141,N_22652);
and UO_1329 (O_1329,N_21079,N_20002);
xor UO_1330 (O_1330,N_20592,N_24675);
nand UO_1331 (O_1331,N_20451,N_22372);
xnor UO_1332 (O_1332,N_22509,N_23193);
nor UO_1333 (O_1333,N_20159,N_23502);
nand UO_1334 (O_1334,N_24416,N_21872);
nand UO_1335 (O_1335,N_22630,N_23067);
xnor UO_1336 (O_1336,N_22123,N_21598);
nor UO_1337 (O_1337,N_23976,N_20052);
nor UO_1338 (O_1338,N_23128,N_22435);
or UO_1339 (O_1339,N_23590,N_21436);
nor UO_1340 (O_1340,N_21073,N_23884);
nand UO_1341 (O_1341,N_23258,N_23399);
or UO_1342 (O_1342,N_20203,N_23817);
and UO_1343 (O_1343,N_24124,N_20743);
nor UO_1344 (O_1344,N_24532,N_22405);
or UO_1345 (O_1345,N_22777,N_22172);
nor UO_1346 (O_1346,N_22036,N_21604);
nand UO_1347 (O_1347,N_23693,N_20692);
or UO_1348 (O_1348,N_23132,N_21641);
xnor UO_1349 (O_1349,N_24935,N_20778);
xor UO_1350 (O_1350,N_20315,N_22349);
or UO_1351 (O_1351,N_20978,N_21466);
and UO_1352 (O_1352,N_20820,N_21723);
nor UO_1353 (O_1353,N_24506,N_23375);
nand UO_1354 (O_1354,N_21549,N_24070);
and UO_1355 (O_1355,N_24424,N_23954);
nor UO_1356 (O_1356,N_20310,N_20570);
nor UO_1357 (O_1357,N_23484,N_21449);
xor UO_1358 (O_1358,N_20591,N_23797);
nor UO_1359 (O_1359,N_22110,N_21555);
or UO_1360 (O_1360,N_23319,N_21404);
nand UO_1361 (O_1361,N_21798,N_22015);
and UO_1362 (O_1362,N_21919,N_21953);
nand UO_1363 (O_1363,N_21118,N_22763);
nor UO_1364 (O_1364,N_22207,N_21770);
nand UO_1365 (O_1365,N_20077,N_24145);
and UO_1366 (O_1366,N_22085,N_24801);
nand UO_1367 (O_1367,N_24631,N_22041);
nand UO_1368 (O_1368,N_21417,N_23980);
nand UO_1369 (O_1369,N_20492,N_22460);
nor UO_1370 (O_1370,N_20332,N_24382);
or UO_1371 (O_1371,N_20940,N_21140);
nor UO_1372 (O_1372,N_20080,N_23208);
nand UO_1373 (O_1373,N_22365,N_22540);
nand UO_1374 (O_1374,N_24236,N_21860);
nand UO_1375 (O_1375,N_23591,N_24536);
xnor UO_1376 (O_1376,N_24995,N_21388);
or UO_1377 (O_1377,N_24040,N_20641);
or UO_1378 (O_1378,N_23600,N_22216);
nand UO_1379 (O_1379,N_21911,N_20931);
nand UO_1380 (O_1380,N_22090,N_23186);
and UO_1381 (O_1381,N_21898,N_23844);
or UO_1382 (O_1382,N_22476,N_23975);
or UO_1383 (O_1383,N_21939,N_20439);
or UO_1384 (O_1384,N_20393,N_22268);
or UO_1385 (O_1385,N_20053,N_23245);
nand UO_1386 (O_1386,N_23398,N_23101);
or UO_1387 (O_1387,N_23085,N_22224);
nand UO_1388 (O_1388,N_23570,N_24913);
or UO_1389 (O_1389,N_20176,N_21145);
nand UO_1390 (O_1390,N_21027,N_20025);
and UO_1391 (O_1391,N_21480,N_24374);
or UO_1392 (O_1392,N_20117,N_20660);
nand UO_1393 (O_1393,N_24091,N_22031);
nor UO_1394 (O_1394,N_22799,N_23905);
and UO_1395 (O_1395,N_20009,N_23691);
or UO_1396 (O_1396,N_22996,N_24008);
or UO_1397 (O_1397,N_23920,N_24159);
nand UO_1398 (O_1398,N_21693,N_22296);
xor UO_1399 (O_1399,N_23701,N_20855);
or UO_1400 (O_1400,N_20556,N_24082);
nand UO_1401 (O_1401,N_21941,N_20068);
xnor UO_1402 (O_1402,N_21651,N_21494);
nand UO_1403 (O_1403,N_21141,N_20125);
nor UO_1404 (O_1404,N_22170,N_24934);
or UO_1405 (O_1405,N_21909,N_21682);
xor UO_1406 (O_1406,N_24741,N_24592);
and UO_1407 (O_1407,N_21547,N_23330);
xnor UO_1408 (O_1408,N_24508,N_20415);
xnor UO_1409 (O_1409,N_21954,N_22055);
nand UO_1410 (O_1410,N_21239,N_23937);
xnor UO_1411 (O_1411,N_23138,N_22650);
xnor UO_1412 (O_1412,N_23939,N_22416);
and UO_1413 (O_1413,N_21385,N_24241);
xor UO_1414 (O_1414,N_21182,N_22228);
or UO_1415 (O_1415,N_23978,N_23017);
or UO_1416 (O_1416,N_20929,N_22261);
nor UO_1417 (O_1417,N_21634,N_23532);
nor UO_1418 (O_1418,N_23622,N_24513);
xor UO_1419 (O_1419,N_20793,N_23739);
xor UO_1420 (O_1420,N_23412,N_20386);
or UO_1421 (O_1421,N_20459,N_21827);
or UO_1422 (O_1422,N_22157,N_22558);
nor UO_1423 (O_1423,N_21168,N_20161);
or UO_1424 (O_1424,N_20605,N_24607);
nor UO_1425 (O_1425,N_24671,N_20625);
or UO_1426 (O_1426,N_22975,N_22315);
or UO_1427 (O_1427,N_21998,N_23692);
nor UO_1428 (O_1428,N_23131,N_20046);
or UO_1429 (O_1429,N_21420,N_23804);
xnor UO_1430 (O_1430,N_21421,N_21951);
and UO_1431 (O_1431,N_23374,N_23324);
xnor UO_1432 (O_1432,N_20228,N_24117);
nand UO_1433 (O_1433,N_23675,N_24400);
nand UO_1434 (O_1434,N_23388,N_24802);
nand UO_1435 (O_1435,N_23987,N_22374);
xor UO_1436 (O_1436,N_20817,N_24316);
or UO_1437 (O_1437,N_24176,N_24450);
xnor UO_1438 (O_1438,N_23039,N_21671);
or UO_1439 (O_1439,N_24351,N_23811);
and UO_1440 (O_1440,N_20703,N_20133);
or UO_1441 (O_1441,N_24891,N_22122);
and UO_1442 (O_1442,N_21884,N_21920);
nor UO_1443 (O_1443,N_20446,N_20848);
xor UO_1444 (O_1444,N_23046,N_20600);
nor UO_1445 (O_1445,N_24920,N_24940);
nor UO_1446 (O_1446,N_22906,N_23778);
and UO_1447 (O_1447,N_20138,N_23333);
nor UO_1448 (O_1448,N_23520,N_23500);
and UO_1449 (O_1449,N_21812,N_21499);
nand UO_1450 (O_1450,N_20304,N_23914);
and UO_1451 (O_1451,N_23619,N_21748);
and UO_1452 (O_1452,N_22924,N_20939);
nand UO_1453 (O_1453,N_21070,N_22867);
or UO_1454 (O_1454,N_20416,N_22621);
nand UO_1455 (O_1455,N_20921,N_23207);
nand UO_1456 (O_1456,N_23617,N_24749);
nand UO_1457 (O_1457,N_21568,N_20757);
nor UO_1458 (O_1458,N_21676,N_22285);
xnor UO_1459 (O_1459,N_21308,N_23416);
nand UO_1460 (O_1460,N_22052,N_22605);
and UO_1461 (O_1461,N_21403,N_23683);
and UO_1462 (O_1462,N_24985,N_24187);
nor UO_1463 (O_1463,N_23979,N_20582);
nand UO_1464 (O_1464,N_23853,N_23447);
xor UO_1465 (O_1465,N_22388,N_23934);
nor UO_1466 (O_1466,N_24398,N_20789);
and UO_1467 (O_1467,N_22185,N_22093);
or UO_1468 (O_1468,N_23608,N_20264);
or UO_1469 (O_1469,N_23898,N_21003);
or UO_1470 (O_1470,N_24701,N_22328);
xor UO_1471 (O_1471,N_23233,N_20066);
xnor UO_1472 (O_1472,N_24108,N_24448);
or UO_1473 (O_1473,N_24660,N_23730);
and UO_1474 (O_1474,N_22318,N_23277);
or UO_1475 (O_1475,N_21025,N_24370);
or UO_1476 (O_1476,N_20088,N_23045);
nand UO_1477 (O_1477,N_23768,N_21903);
and UO_1478 (O_1478,N_24365,N_24112);
or UO_1479 (O_1479,N_22722,N_21943);
and UO_1480 (O_1480,N_21906,N_20936);
or UO_1481 (O_1481,N_21500,N_22535);
or UO_1482 (O_1482,N_20877,N_24387);
nand UO_1483 (O_1483,N_23134,N_22008);
and UO_1484 (O_1484,N_24851,N_21802);
and UO_1485 (O_1485,N_24356,N_22499);
nand UO_1486 (O_1486,N_21300,N_20513);
and UO_1487 (O_1487,N_23110,N_24839);
or UO_1488 (O_1488,N_22200,N_24303);
xor UO_1489 (O_1489,N_21272,N_21516);
xnor UO_1490 (O_1490,N_23611,N_24704);
or UO_1491 (O_1491,N_20768,N_20615);
nor UO_1492 (O_1492,N_21355,N_22677);
xor UO_1493 (O_1493,N_20469,N_23012);
nand UO_1494 (O_1494,N_23847,N_24626);
nor UO_1495 (O_1495,N_21243,N_23149);
xnor UO_1496 (O_1496,N_22427,N_24157);
nand UO_1497 (O_1497,N_24988,N_21621);
nor UO_1498 (O_1498,N_21647,N_20380);
or UO_1499 (O_1499,N_20227,N_23488);
nor UO_1500 (O_1500,N_20672,N_22131);
and UO_1501 (O_1501,N_20142,N_24371);
and UO_1502 (O_1502,N_24411,N_23445);
and UO_1503 (O_1503,N_21492,N_24773);
xor UO_1504 (O_1504,N_20992,N_24433);
nand UO_1505 (O_1505,N_24379,N_20259);
xnor UO_1506 (O_1506,N_22508,N_21080);
nand UO_1507 (O_1507,N_22004,N_20911);
xor UO_1508 (O_1508,N_23776,N_21762);
nor UO_1509 (O_1509,N_24639,N_20826);
or UO_1510 (O_1510,N_22889,N_21454);
and UO_1511 (O_1511,N_20844,N_20948);
nand UO_1512 (O_1512,N_23704,N_23268);
nor UO_1513 (O_1513,N_21115,N_23702);
or UO_1514 (O_1514,N_21108,N_23118);
or UO_1515 (O_1515,N_24941,N_20430);
and UO_1516 (O_1516,N_24326,N_22159);
and UO_1517 (O_1517,N_23761,N_20918);
and UO_1518 (O_1518,N_21942,N_24699);
or UO_1519 (O_1519,N_20764,N_22286);
or UO_1520 (O_1520,N_22936,N_20093);
xnor UO_1521 (O_1521,N_24769,N_20431);
nor UO_1522 (O_1522,N_21029,N_22025);
or UO_1523 (O_1523,N_20565,N_20198);
or UO_1524 (O_1524,N_22454,N_24656);
nor UO_1525 (O_1525,N_22250,N_23781);
xnor UO_1526 (O_1526,N_20943,N_23082);
nand UO_1527 (O_1527,N_22445,N_21318);
nor UO_1528 (O_1528,N_20240,N_22959);
and UO_1529 (O_1529,N_21000,N_24625);
or UO_1530 (O_1530,N_23790,N_20530);
and UO_1531 (O_1531,N_22665,N_23897);
nand UO_1532 (O_1532,N_24328,N_22424);
or UO_1533 (O_1533,N_24441,N_22849);
and UO_1534 (O_1534,N_22118,N_22490);
nand UO_1535 (O_1535,N_20555,N_22084);
xor UO_1536 (O_1536,N_21229,N_21447);
xor UO_1537 (O_1537,N_23850,N_21614);
xnor UO_1538 (O_1538,N_22520,N_23383);
or UO_1539 (O_1539,N_22294,N_24288);
and UO_1540 (O_1540,N_24113,N_23063);
xnor UO_1541 (O_1541,N_21741,N_23671);
nand UO_1542 (O_1542,N_24987,N_23433);
nor UO_1543 (O_1543,N_20690,N_21238);
or UO_1544 (O_1544,N_22109,N_20656);
and UO_1545 (O_1545,N_23028,N_22744);
nor UO_1546 (O_1546,N_20324,N_22711);
and UO_1547 (O_1547,N_20717,N_22861);
xnor UO_1548 (O_1548,N_23686,N_20955);
or UO_1549 (O_1549,N_24596,N_20187);
nand UO_1550 (O_1550,N_24893,N_20627);
and UO_1551 (O_1551,N_24642,N_21815);
or UO_1552 (O_1552,N_24638,N_22449);
nor UO_1553 (O_1553,N_21149,N_21160);
xnor UO_1554 (O_1554,N_21643,N_24805);
and UO_1555 (O_1555,N_23596,N_22531);
and UO_1556 (O_1556,N_20220,N_24079);
and UO_1557 (O_1557,N_21541,N_24888);
xor UO_1558 (O_1558,N_22289,N_20952);
nand UO_1559 (O_1559,N_23476,N_20175);
nor UO_1560 (O_1560,N_23862,N_20309);
xnor UO_1561 (O_1561,N_24325,N_22597);
xor UO_1562 (O_1562,N_22935,N_22255);
nor UO_1563 (O_1563,N_22297,N_20146);
and UO_1564 (O_1564,N_21721,N_22230);
and UO_1565 (O_1565,N_22189,N_23900);
or UO_1566 (O_1566,N_21935,N_24688);
and UO_1567 (O_1567,N_21583,N_20854);
and UO_1568 (O_1568,N_22582,N_20210);
nand UO_1569 (O_1569,N_20998,N_23206);
and UO_1570 (O_1570,N_24558,N_24046);
or UO_1571 (O_1571,N_21971,N_22027);
nand UO_1572 (O_1572,N_20882,N_20097);
or UO_1573 (O_1573,N_22792,N_22149);
xnor UO_1574 (O_1574,N_22755,N_22833);
xor UO_1575 (O_1575,N_20792,N_21043);
xor UO_1576 (O_1576,N_24880,N_22854);
nand UO_1577 (O_1577,N_23765,N_23871);
nor UO_1578 (O_1578,N_22426,N_23226);
nor UO_1579 (O_1579,N_20360,N_21335);
nor UO_1580 (O_1580,N_20026,N_24640);
nor UO_1581 (O_1581,N_21657,N_23995);
nor UO_1582 (O_1582,N_24041,N_23114);
nand UO_1583 (O_1583,N_22033,N_24530);
or UO_1584 (O_1584,N_22921,N_23421);
and UO_1585 (O_1585,N_21336,N_24150);
xor UO_1586 (O_1586,N_23501,N_21165);
nor UO_1587 (O_1587,N_23813,N_21826);
or UO_1588 (O_1588,N_24597,N_21251);
or UO_1589 (O_1589,N_21294,N_22595);
nor UO_1590 (O_1590,N_24694,N_20252);
or UO_1591 (O_1591,N_23628,N_21015);
xnor UO_1592 (O_1592,N_22304,N_21314);
xor UO_1593 (O_1593,N_22321,N_22946);
or UO_1594 (O_1594,N_23255,N_20241);
or UO_1595 (O_1595,N_23805,N_20860);
nand UO_1596 (O_1596,N_24208,N_21401);
xnor UO_1597 (O_1597,N_23386,N_23942);
or UO_1598 (O_1598,N_24185,N_21777);
and UO_1599 (O_1599,N_21862,N_20262);
xor UO_1600 (O_1600,N_21225,N_21829);
or UO_1601 (O_1601,N_23745,N_24469);
and UO_1602 (O_1602,N_22327,N_21835);
or UO_1603 (O_1603,N_21147,N_20195);
nand UO_1604 (O_1604,N_23757,N_20308);
and UO_1605 (O_1605,N_22631,N_20418);
nand UO_1606 (O_1606,N_24036,N_24509);
and UO_1607 (O_1607,N_21477,N_21716);
or UO_1608 (O_1608,N_20405,N_20507);
nand UO_1609 (O_1609,N_20065,N_24628);
and UO_1610 (O_1610,N_21532,N_24729);
xor UO_1611 (O_1611,N_20289,N_23630);
nor UO_1612 (O_1612,N_22795,N_20784);
xnor UO_1613 (O_1613,N_20508,N_20350);
nand UO_1614 (O_1614,N_20695,N_21297);
nor UO_1615 (O_1615,N_20908,N_22182);
nor UO_1616 (O_1616,N_23257,N_24959);
nand UO_1617 (O_1617,N_23714,N_21459);
xnor UO_1618 (O_1618,N_24063,N_24516);
nand UO_1619 (O_1619,N_20051,N_24754);
and UO_1620 (O_1620,N_22021,N_24244);
nand UO_1621 (O_1621,N_22541,N_21579);
nand UO_1622 (O_1622,N_24209,N_24590);
xor UO_1623 (O_1623,N_23496,N_21087);
xor UO_1624 (O_1624,N_21488,N_23777);
and UO_1625 (O_1625,N_22592,N_22673);
and UO_1626 (O_1626,N_22721,N_24890);
or UO_1627 (O_1627,N_21599,N_22164);
xor UO_1628 (O_1628,N_20560,N_22188);
xnor UO_1629 (O_1629,N_20687,N_23260);
nor UO_1630 (O_1630,N_21772,N_23024);
and UO_1631 (O_1631,N_21091,N_21805);
nor UO_1632 (O_1632,N_22496,N_22561);
nand UO_1633 (O_1633,N_24186,N_24014);
nor UO_1634 (O_1634,N_22079,N_21337);
nor UO_1635 (O_1635,N_23859,N_21281);
nand UO_1636 (O_1636,N_20423,N_20299);
nand UO_1637 (O_1637,N_21227,N_23894);
and UO_1638 (O_1638,N_24076,N_20542);
or UO_1639 (O_1639,N_24783,N_22175);
and UO_1640 (O_1640,N_22797,N_22141);
and UO_1641 (O_1641,N_21665,N_21429);
nand UO_1642 (O_1642,N_20484,N_20669);
nor UO_1643 (O_1643,N_23430,N_24197);
nor UO_1644 (O_1644,N_21210,N_22770);
xnor UO_1645 (O_1645,N_22259,N_20236);
nand UO_1646 (O_1646,N_20554,N_22784);
xnor UO_1647 (O_1647,N_24207,N_20403);
nor UO_1648 (O_1648,N_20031,N_24680);
or UO_1649 (O_1649,N_20959,N_21569);
or UO_1650 (O_1650,N_20470,N_23950);
or UO_1651 (O_1651,N_20128,N_21166);
xor UO_1652 (O_1652,N_20367,N_23676);
or UO_1653 (O_1653,N_21675,N_20541);
and UO_1654 (O_1654,N_22010,N_21801);
and UO_1655 (O_1655,N_23037,N_22809);
nand UO_1656 (O_1656,N_24136,N_24630);
xor UO_1657 (O_1657,N_22301,N_22152);
xnor UO_1658 (O_1658,N_20208,N_21538);
nor UO_1659 (O_1659,N_20217,N_23127);
xnor UO_1660 (O_1660,N_22234,N_23873);
nand UO_1661 (O_1661,N_22431,N_21139);
nor UO_1662 (O_1662,N_23435,N_23241);
and UO_1663 (O_1663,N_20160,N_22034);
nand UO_1664 (O_1664,N_21760,N_23014);
and UO_1665 (O_1665,N_23647,N_23080);
nand UO_1666 (O_1666,N_20253,N_23346);
and UO_1667 (O_1667,N_22944,N_24226);
xor UO_1668 (O_1668,N_21779,N_22659);
xnor UO_1669 (O_1669,N_20580,N_22963);
or UO_1670 (O_1670,N_21479,N_24267);
nor UO_1671 (O_1671,N_24007,N_24327);
and UO_1672 (O_1672,N_22954,N_24898);
and UO_1673 (O_1673,N_24799,N_22165);
nor UO_1674 (O_1674,N_21868,N_24809);
nand UO_1675 (O_1675,N_24119,N_22383);
nor UO_1676 (O_1676,N_23088,N_21207);
nand UO_1677 (O_1677,N_23365,N_24670);
or UO_1678 (O_1678,N_22942,N_20862);
or UO_1679 (O_1679,N_23247,N_20061);
and UO_1680 (O_1680,N_22629,N_20754);
or UO_1681 (O_1681,N_23638,N_21518);
or UO_1682 (O_1682,N_22201,N_21278);
nand UO_1683 (O_1683,N_20189,N_20684);
xnor UO_1684 (O_1684,N_20909,N_21674);
xnor UO_1685 (O_1685,N_20698,N_20082);
nor UO_1686 (O_1686,N_24129,N_22837);
xnor UO_1687 (O_1687,N_21574,N_20694);
and UO_1688 (O_1688,N_21298,N_20126);
xnor UO_1689 (O_1689,N_24498,N_24831);
or UO_1690 (O_1690,N_24408,N_23304);
or UO_1691 (O_1691,N_20328,N_21033);
xor UO_1692 (O_1692,N_21708,N_22633);
or UO_1693 (O_1693,N_23679,N_22329);
or UO_1694 (O_1694,N_23051,N_24231);
nand UO_1695 (O_1695,N_23076,N_23715);
and UO_1696 (O_1696,N_23307,N_21640);
xnor UO_1697 (O_1697,N_21112,N_23656);
nor UO_1698 (O_1698,N_20078,N_24683);
and UO_1699 (O_1699,N_22235,N_23733);
and UO_1700 (O_1700,N_21356,N_23366);
xnor UO_1701 (O_1701,N_21867,N_23112);
or UO_1702 (O_1702,N_24126,N_20987);
and UO_1703 (O_1703,N_23176,N_24463);
and UO_1704 (O_1704,N_21373,N_20883);
nor UO_1705 (O_1705,N_24366,N_23901);
and UO_1706 (O_1706,N_22524,N_22871);
nand UO_1707 (O_1707,N_22823,N_20934);
and UO_1708 (O_1708,N_20285,N_22726);
or UO_1709 (O_1709,N_20190,N_21992);
or UO_1710 (O_1710,N_24361,N_24451);
or UO_1711 (O_1711,N_23584,N_21481);
or UO_1712 (O_1712,N_21023,N_22114);
nor UO_1713 (O_1713,N_23499,N_20748);
or UO_1714 (O_1714,N_22952,N_23023);
and UO_1715 (O_1715,N_22626,N_22815);
nand UO_1716 (O_1716,N_24871,N_22587);
or UO_1717 (O_1717,N_20342,N_21853);
or UO_1718 (O_1718,N_21979,N_20136);
xnor UO_1719 (O_1719,N_21327,N_22282);
and UO_1720 (O_1720,N_24479,N_23881);
xnor UO_1721 (O_1721,N_22302,N_20103);
nor UO_1722 (O_1722,N_20390,N_21191);
nor UO_1723 (O_1723,N_22489,N_24436);
nor UO_1724 (O_1724,N_23010,N_24766);
or UO_1725 (O_1725,N_22081,N_22865);
xor UO_1726 (O_1726,N_22759,N_23809);
or UO_1727 (O_1727,N_24048,N_21268);
nand UO_1728 (O_1728,N_23033,N_21307);
nand UO_1729 (O_1729,N_24219,N_20145);
or UO_1730 (O_1730,N_21383,N_24016);
nand UO_1731 (O_1731,N_24553,N_24828);
or UO_1732 (O_1732,N_22498,N_22708);
and UO_1733 (O_1733,N_23734,N_20685);
nand UO_1734 (O_1734,N_22981,N_23512);
xor UO_1735 (O_1735,N_21402,N_21304);
nand UO_1736 (O_1736,N_24971,N_20229);
nand UO_1737 (O_1737,N_23177,N_20894);
nand UO_1738 (O_1738,N_20072,N_23678);
xor UO_1739 (O_1739,N_20234,N_20497);
xor UO_1740 (O_1740,N_21384,N_20351);
or UO_1741 (O_1741,N_22241,N_20522);
xor UO_1742 (O_1742,N_20284,N_21446);
and UO_1743 (O_1743,N_23903,N_24798);
xnor UO_1744 (O_1744,N_21129,N_24644);
and UO_1745 (O_1745,N_24367,N_20573);
and UO_1746 (O_1746,N_20412,N_22393);
nand UO_1747 (O_1747,N_24591,N_23916);
and UO_1748 (O_1748,N_23524,N_20749);
xor UO_1749 (O_1749,N_23670,N_22260);
nor UO_1750 (O_1750,N_24060,N_23357);
or UO_1751 (O_1751,N_21831,N_24771);
nor UO_1752 (O_1752,N_20294,N_24551);
and UO_1753 (O_1753,N_22421,N_24228);
xor UO_1754 (O_1754,N_22111,N_22549);
nor UO_1755 (O_1755,N_23440,N_20927);
nand UO_1756 (O_1756,N_24221,N_21924);
and UO_1757 (O_1757,N_24674,N_22274);
nand UO_1758 (O_1758,N_23598,N_20118);
and UO_1759 (O_1759,N_24161,N_22679);
nor UO_1760 (O_1760,N_24372,N_20221);
and UO_1761 (O_1761,N_23597,N_21611);
and UO_1762 (O_1762,N_20312,N_20578);
nand UO_1763 (O_1763,N_20526,N_21683);
nand UO_1764 (O_1764,N_23674,N_20840);
nor UO_1765 (O_1765,N_20481,N_20988);
and UO_1766 (O_1766,N_23152,N_22604);
nand UO_1767 (O_1767,N_23878,N_21476);
nand UO_1768 (O_1768,N_23718,N_21783);
xnor UO_1769 (O_1769,N_24517,N_20163);
nor UO_1770 (O_1770,N_23648,N_21645);
and UO_1771 (O_1771,N_21724,N_21704);
nand UO_1772 (O_1772,N_24406,N_23229);
or UO_1773 (O_1773,N_22254,N_22866);
xnor UO_1774 (O_1774,N_24826,N_20846);
and UO_1775 (O_1775,N_24302,N_23929);
nand UO_1776 (O_1776,N_21186,N_20962);
nand UO_1777 (O_1777,N_23883,N_22593);
and UO_1778 (O_1778,N_22937,N_24093);
and UO_1779 (O_1779,N_22636,N_20733);
or UO_1780 (O_1780,N_21737,N_23136);
or UO_1781 (O_1781,N_23955,N_24797);
or UO_1782 (O_1782,N_21615,N_23752);
or UO_1783 (O_1783,N_23836,N_20933);
nand UO_1784 (O_1784,N_23246,N_23517);
nand UO_1785 (O_1785,N_21228,N_21325);
or UO_1786 (O_1786,N_22210,N_22859);
and UO_1787 (O_1787,N_22020,N_23863);
nand UO_1788 (O_1788,N_20172,N_23601);
nor UO_1789 (O_1789,N_21705,N_21988);
nand UO_1790 (O_1790,N_20022,N_20634);
nand UO_1791 (O_1791,N_23665,N_24277);
or UO_1792 (O_1792,N_21011,N_21121);
xnor UO_1793 (O_1793,N_24931,N_20567);
and UO_1794 (O_1794,N_24106,N_23317);
and UO_1795 (O_1795,N_21231,N_20426);
nand UO_1796 (O_1796,N_22218,N_21507);
xor UO_1797 (O_1797,N_23181,N_22914);
or UO_1798 (O_1798,N_22019,N_24142);
nor UO_1799 (O_1799,N_21275,N_24862);
nand UO_1800 (O_1800,N_22065,N_23006);
nor UO_1801 (O_1801,N_21781,N_24493);
or UO_1802 (O_1802,N_22319,N_20890);
nor UO_1803 (O_1803,N_24033,N_20614);
nor UO_1804 (O_1804,N_20865,N_21064);
nand UO_1805 (O_1805,N_22902,N_21757);
xnor UO_1806 (O_1806,N_22414,N_24052);
nand UO_1807 (O_1807,N_24291,N_21804);
nand UO_1808 (O_1808,N_24918,N_20491);
and UO_1809 (O_1809,N_22646,N_21600);
nor UO_1810 (O_1810,N_21857,N_21260);
xor UO_1811 (O_1811,N_20823,N_24584);
nand UO_1812 (O_1812,N_21656,N_23748);
xor UO_1813 (O_1813,N_22819,N_24709);
nand UO_1814 (O_1814,N_22783,N_24237);
nor UO_1815 (O_1815,N_23851,N_22082);
xor UO_1816 (O_1816,N_20898,N_20750);
and UO_1817 (O_1817,N_22729,N_21625);
nor UO_1818 (O_1818,N_23195,N_20086);
xor UO_1819 (O_1819,N_21452,N_20914);
nand UO_1820 (O_1820,N_24227,N_22801);
and UO_1821 (O_1821,N_20553,N_23636);
xnor UO_1822 (O_1822,N_20361,N_20204);
or UO_1823 (O_1823,N_23189,N_24467);
and UO_1824 (O_1824,N_23034,N_24763);
or UO_1825 (O_1825,N_23743,N_21662);
xor UO_1826 (O_1826,N_22339,N_20059);
nor UO_1827 (O_1827,N_22115,N_22129);
nor UO_1828 (O_1828,N_22796,N_21905);
nor UO_1829 (O_1829,N_20897,N_22217);
xnor UO_1830 (O_1830,N_21778,N_23766);
and UO_1831 (O_1831,N_20173,N_23408);
or UO_1832 (O_1832,N_21357,N_22501);
nor UO_1833 (O_1833,N_23188,N_23489);
or UO_1834 (O_1834,N_20281,N_24713);
xnor UO_1835 (O_1835,N_23159,N_23999);
nor UO_1836 (O_1836,N_22251,N_24488);
or UO_1837 (O_1837,N_24752,N_24939);
nand UO_1838 (O_1838,N_20278,N_23448);
or UO_1839 (O_1839,N_24323,N_22857);
nand UO_1840 (O_1840,N_22262,N_20275);
and UO_1841 (O_1841,N_20679,N_22231);
or UO_1842 (O_1842,N_20836,N_24742);
or UO_1843 (O_1843,N_22882,N_23096);
xnor UO_1844 (O_1844,N_21813,N_24775);
xnor UO_1845 (O_1845,N_20830,N_23054);
nand UO_1846 (O_1846,N_20683,N_23378);
nand UO_1847 (O_1847,N_23197,N_24991);
and UO_1848 (O_1848,N_20500,N_24745);
xnor UO_1849 (O_1849,N_24001,N_24501);
or UO_1850 (O_1850,N_22757,N_24710);
xor UO_1851 (O_1851,N_23928,N_23165);
xor UO_1852 (O_1852,N_20402,N_24522);
and UO_1853 (O_1853,N_22660,N_20759);
nand UO_1854 (O_1854,N_23108,N_23099);
nand UO_1855 (O_1855,N_22322,N_24853);
nand UO_1856 (O_1856,N_24341,N_21026);
xnor UO_1857 (O_1857,N_21144,N_24480);
nor UO_1858 (O_1858,N_20561,N_22457);
nor UO_1859 (O_1859,N_23018,N_21913);
nor UO_1860 (O_1860,N_21247,N_20991);
and UO_1861 (O_1861,N_20968,N_22737);
nor UO_1862 (O_1862,N_22735,N_24149);
and UO_1863 (O_1863,N_22355,N_22199);
and UO_1864 (O_1864,N_23007,N_22309);
xnor UO_1865 (O_1865,N_21093,N_24081);
nor UO_1866 (O_1866,N_20903,N_23658);
nor UO_1867 (O_1867,N_23401,N_20323);
and UO_1868 (O_1868,N_20504,N_22620);
xor UO_1869 (O_1869,N_22568,N_22271);
or UO_1870 (O_1870,N_21740,N_21711);
or UO_1871 (O_1871,N_22440,N_22430);
nand UO_1872 (O_1872,N_24595,N_23540);
and UO_1873 (O_1873,N_21008,N_21863);
nor UO_1874 (O_1874,N_23395,N_20664);
xor UO_1875 (O_1875,N_23394,N_20356);
and UO_1876 (O_1876,N_23352,N_23242);
nand UO_1877 (O_1877,N_24568,N_20772);
and UO_1878 (O_1878,N_24523,N_24882);
xor UO_1879 (O_1879,N_24270,N_22137);
xnor UO_1880 (O_1880,N_20110,N_24257);
and UO_1881 (O_1881,N_20011,N_24902);
nor UO_1882 (O_1882,N_23908,N_20598);
and UO_1883 (O_1883,N_22884,N_22121);
nor UO_1884 (O_1884,N_24483,N_22419);
nand UO_1885 (O_1885,N_20182,N_24153);
nor UO_1886 (O_1886,N_21096,N_21961);
and UO_1887 (O_1887,N_24103,N_21987);
nor UO_1888 (O_1888,N_24495,N_21690);
nand UO_1889 (O_1889,N_20753,N_24446);
xor UO_1890 (O_1890,N_20675,N_23708);
nor UO_1891 (O_1891,N_21083,N_23492);
or UO_1892 (O_1892,N_22275,N_22432);
or UO_1893 (O_1893,N_20233,N_21512);
nand UO_1894 (O_1894,N_22058,N_22655);
nand UO_1895 (O_1895,N_20718,N_22303);
and UO_1896 (O_1896,N_20213,N_23272);
nor UO_1897 (O_1897,N_24065,N_22601);
xor UO_1898 (O_1898,N_21696,N_20094);
nor UO_1899 (O_1899,N_22895,N_22960);
nand UO_1900 (O_1900,N_23985,N_22971);
xor UO_1901 (O_1901,N_24180,N_23223);
or UO_1902 (O_1902,N_20972,N_21734);
and UO_1903 (O_1903,N_23513,N_21957);
and UO_1904 (O_1904,N_24115,N_22417);
and UO_1905 (O_1905,N_23664,N_24692);
nor UO_1906 (O_1906,N_20444,N_21830);
nand UO_1907 (O_1907,N_22376,N_20196);
xnor UO_1908 (O_1908,N_20438,N_20153);
nor UO_1909 (O_1909,N_23857,N_24535);
xor UO_1910 (O_1910,N_24217,N_20869);
nand UO_1911 (O_1911,N_21222,N_22397);
and UO_1912 (O_1912,N_21255,N_22774);
and UO_1913 (O_1913,N_20884,N_22576);
nand UO_1914 (O_1914,N_20292,N_24474);
and UO_1915 (O_1915,N_21727,N_24317);
and UO_1916 (O_1916,N_22785,N_22442);
xnor UO_1917 (O_1917,N_20509,N_21997);
nor UO_1918 (O_1918,N_21412,N_23455);
and UO_1919 (O_1919,N_23230,N_21497);
nor UO_1920 (O_1920,N_24251,N_22584);
or UO_1921 (O_1921,N_24531,N_20867);
nand UO_1922 (O_1922,N_20970,N_23123);
nand UO_1923 (O_1923,N_24658,N_22007);
or UO_1924 (O_1924,N_23470,N_22526);
and UO_1925 (O_1925,N_20770,N_21464);
xor UO_1926 (O_1926,N_20667,N_24965);
nor UO_1927 (O_1927,N_22839,N_24966);
or UO_1928 (O_1928,N_21702,N_22504);
or UO_1929 (O_1929,N_24840,N_20628);
nand UO_1930 (O_1930,N_21117,N_23095);
and UO_1931 (O_1931,N_21730,N_24230);
xnor UO_1932 (O_1932,N_23161,N_24238);
and UO_1933 (O_1933,N_23196,N_24883);
xor UO_1934 (O_1934,N_22465,N_24332);
nand UO_1935 (O_1935,N_23074,N_21901);
xnor UO_1936 (O_1936,N_24849,N_23913);
and UO_1937 (O_1937,N_20868,N_23069);
nor UO_1938 (O_1938,N_20192,N_21418);
nor UO_1939 (O_1939,N_24143,N_20479);
nand UO_1940 (O_1940,N_23100,N_20249);
nand UO_1941 (O_1941,N_21965,N_22202);
nor UO_1942 (O_1942,N_24074,N_22745);
nor UO_1943 (O_1943,N_23659,N_21774);
nor UO_1944 (O_1944,N_24868,N_23282);
or UO_1945 (O_1945,N_24845,N_24818);
xor UO_1946 (O_1946,N_22451,N_22176);
and UO_1947 (O_1947,N_24643,N_22614);
or UO_1948 (O_1948,N_22106,N_20715);
nor UO_1949 (O_1949,N_23461,N_22348);
and UO_1950 (O_1950,N_24700,N_23599);
nor UO_1951 (O_1951,N_24973,N_22766);
xor UO_1952 (O_1952,N_23065,N_24174);
xor UO_1953 (O_1953,N_24392,N_21811);
nand UO_1954 (O_1954,N_24245,N_21110);
nor UO_1955 (O_1955,N_24430,N_24976);
nand UO_1956 (O_1956,N_21878,N_22392);
nor UO_1957 (O_1957,N_20345,N_20971);
nand UO_1958 (O_1958,N_22938,N_21896);
nor UO_1959 (O_1959,N_23839,N_20121);
and UO_1960 (O_1960,N_24767,N_23807);
xor UO_1961 (O_1961,N_24496,N_23071);
and UO_1962 (O_1962,N_20150,N_23705);
nand UO_1963 (O_1963,N_22089,N_21127);
nand UO_1964 (O_1964,N_21458,N_22343);
nor UO_1965 (O_1965,N_24223,N_21323);
xnor UO_1966 (O_1966,N_22237,N_20419);
or UO_1967 (O_1967,N_22961,N_24620);
or UO_1968 (O_1968,N_24468,N_23162);
nand UO_1969 (O_1969,N_20785,N_22765);
or UO_1970 (O_1970,N_23200,N_21116);
or UO_1971 (O_1971,N_23988,N_20900);
xnor UO_1972 (O_1972,N_21254,N_24196);
and UO_1973 (O_1973,N_20503,N_24803);
nand UO_1974 (O_1974,N_22168,N_22310);
nor UO_1975 (O_1975,N_23274,N_22536);
xnor UO_1976 (O_1976,N_23133,N_21352);
nor UO_1977 (O_1977,N_21692,N_20320);
or UO_1978 (O_1978,N_20697,N_22455);
and UO_1979 (O_1979,N_20089,N_23609);
nor UO_1980 (O_1980,N_20087,N_23707);
nand UO_1981 (O_1981,N_20859,N_21776);
xnor UO_1982 (O_1982,N_23649,N_24726);
xnor UO_1983 (O_1983,N_23308,N_22147);
nor UO_1984 (O_1984,N_20575,N_22513);
and UO_1985 (O_1985,N_22276,N_22030);
or UO_1986 (O_1986,N_24345,N_23382);
or UO_1987 (O_1987,N_22101,N_20290);
nand UO_1988 (O_1988,N_20919,N_20747);
xor UO_1989 (O_1989,N_20852,N_21362);
xnor UO_1990 (O_1990,N_21608,N_21071);
xor UO_1991 (O_1991,N_20458,N_22155);
or UO_1992 (O_1992,N_22600,N_23735);
xnor UO_1993 (O_1993,N_23089,N_23808);
or UO_1994 (O_1994,N_22191,N_23289);
and UO_1995 (O_1995,N_22580,N_24609);
and UO_1996 (O_1996,N_20291,N_22142);
or UO_1997 (O_1997,N_24698,N_24442);
nor UO_1998 (O_1998,N_22622,N_21364);
nand UO_1999 (O_1999,N_23814,N_22515);
or UO_2000 (O_2000,N_23288,N_20334);
nor UO_2001 (O_2001,N_21280,N_23588);
nand UO_2002 (O_2002,N_22676,N_22523);
xnor UO_2003 (O_2003,N_22559,N_24610);
xnor UO_2004 (O_2004,N_22943,N_21463);
nand UO_2005 (O_2005,N_24822,N_23899);
xor UO_2006 (O_2006,N_20576,N_24058);
nor UO_2007 (O_2007,N_23605,N_21850);
nand UO_2008 (O_2008,N_20337,N_23403);
or UO_2009 (O_2009,N_21567,N_20149);
or UO_2010 (O_2010,N_22107,N_21528);
xnor UO_2011 (O_2011,N_24352,N_24214);
or UO_2012 (O_2012,N_22211,N_20132);
and UO_2013 (O_2013,N_24562,N_24350);
and UO_2014 (O_2014,N_22258,N_23528);
nand UO_2015 (O_2015,N_23094,N_22926);
or UO_2016 (O_2016,N_23815,N_21358);
or UO_2017 (O_2017,N_23854,N_22134);
xor UO_2018 (O_2018,N_21695,N_22560);
or UO_2019 (O_2019,N_20427,N_20218);
xnor UO_2020 (O_2020,N_24156,N_21097);
and UO_2021 (O_2021,N_23425,N_23203);
or UO_2022 (O_2022,N_24166,N_21234);
nor UO_2023 (O_2023,N_23431,N_20665);
or UO_2024 (O_2024,N_21493,N_20177);
xor UO_2025 (O_2025,N_23613,N_23490);
nand UO_2026 (O_2026,N_20376,N_22071);
nand UO_2027 (O_2027,N_23390,N_24342);
xnor UO_2028 (O_2028,N_23571,N_22379);
and UO_2029 (O_2029,N_22091,N_20127);
nor UO_2030 (O_2030,N_20949,N_22017);
and UO_2031 (O_2031,N_21398,N_22893);
nor UO_2032 (O_2032,N_22404,N_21246);
xnor UO_2033 (O_2033,N_22542,N_23578);
or UO_2034 (O_2034,N_21473,N_24855);
nor UO_2035 (O_2035,N_23710,N_20247);
nor UO_2036 (O_2036,N_22466,N_23515);
and UO_2037 (O_2037,N_22001,N_22553);
or UO_2038 (O_2038,N_23654,N_23652);
xor UO_2039 (O_2039,N_23880,N_21949);
nand UO_2040 (O_2040,N_20777,N_22443);
nor UO_2041 (O_2041,N_20782,N_21893);
nor UO_2042 (O_2042,N_21816,N_24336);
nand UO_2043 (O_2043,N_21565,N_20295);
nor UO_2044 (O_2044,N_20613,N_21153);
and UO_2045 (O_2045,N_22728,N_24497);
and UO_2046 (O_2046,N_22420,N_24155);
nand UO_2047 (O_2047,N_20394,N_23660);
or UO_2048 (O_2048,N_22664,N_20023);
and UO_2049 (O_2049,N_22901,N_21253);
nand UO_2050 (O_2050,N_24363,N_22249);
or UO_2051 (O_2051,N_20941,N_21649);
and UO_2052 (O_2052,N_24528,N_21550);
nand UO_2053 (O_2053,N_21084,N_22100);
or UO_2054 (O_2054,N_22087,N_22829);
nand UO_2055 (O_2055,N_22092,N_20811);
xnor UO_2056 (O_2056,N_24986,N_21081);
nor UO_2057 (O_2057,N_22870,N_22533);
and UO_2058 (O_2058,N_24269,N_24297);
xor UO_2059 (O_2059,N_20108,N_23170);
xnor UO_2060 (O_2060,N_21288,N_24027);
and UO_2061 (O_2061,N_20000,N_23436);
or UO_2062 (O_2062,N_23173,N_24938);
nand UO_2063 (O_2063,N_23026,N_24253);
or UO_2064 (O_2064,N_22221,N_24708);
nor UO_2065 (O_2065,N_22550,N_23364);
or UO_2066 (O_2066,N_24731,N_23822);
nand UO_2067 (O_2067,N_22743,N_22534);
xnor UO_2068 (O_2068,N_20269,N_21038);
nor UO_2069 (O_2069,N_20888,N_21174);
nand UO_2070 (O_2070,N_21846,N_22359);
nor UO_2071 (O_2071,N_20298,N_21694);
or UO_2072 (O_2072,N_20137,N_22511);
xor UO_2073 (O_2073,N_20989,N_21630);
nor UO_2074 (O_2074,N_23806,N_24542);
and UO_2075 (O_2075,N_21406,N_20019);
nand UO_2076 (O_2076,N_23533,N_21706);
xnor UO_2077 (O_2077,N_20170,N_24262);
or UO_2078 (O_2078,N_22810,N_21715);
nand UO_2079 (O_2079,N_24240,N_21045);
xor UO_2080 (O_2080,N_20654,N_22949);
and UO_2081 (O_2081,N_22161,N_21057);
nor UO_2082 (O_2082,N_20329,N_20463);
or UO_2083 (O_2083,N_22758,N_20318);
nor UO_2084 (O_2084,N_22503,N_23823);
xnor UO_2085 (O_2085,N_24577,N_22831);
nand UO_2086 (O_2086,N_20461,N_23832);
or UO_2087 (O_2087,N_24160,N_21387);
nand UO_2088 (O_2088,N_20162,N_20579);
xor UO_2089 (O_2089,N_21592,N_23615);
and UO_2090 (O_2090,N_21540,N_23083);
and UO_2091 (O_2091,N_23002,N_23924);
xnor UO_2092 (O_2092,N_24146,N_20113);
nor UO_2093 (O_2093,N_21148,N_24407);
xnor UO_2094 (O_2094,N_21873,N_21113);
xor UO_2095 (O_2095,N_23506,N_21687);
or UO_2096 (O_2096,N_23373,N_23595);
and UO_2097 (O_2097,N_24438,N_22408);
xnor UO_2098 (O_2098,N_22462,N_22049);
or UO_2099 (O_2099,N_24969,N_23315);
and UO_2100 (O_2100,N_20804,N_23458);
or UO_2101 (O_2101,N_23984,N_23218);
nand UO_2102 (O_2102,N_22776,N_24409);
xnor UO_2103 (O_2103,N_23662,N_24376);
or UO_2104 (O_2104,N_24843,N_22896);
nor UO_2105 (O_2105,N_24537,N_24963);
or UO_2106 (O_2106,N_21546,N_20286);
or UO_2107 (O_2107,N_20533,N_23602);
nor UO_2108 (O_2108,N_23109,N_21341);
or UO_2109 (O_2109,N_20191,N_21257);
xnor UO_2110 (O_2110,N_22699,N_21063);
and UO_2111 (O_2111,N_23437,N_20003);
nor UO_2112 (O_2112,N_24039,N_24634);
and UO_2113 (O_2113,N_20845,N_21156);
and UO_2114 (O_2114,N_23468,N_21974);
and UO_2115 (O_2115,N_22838,N_24101);
and UO_2116 (O_2116,N_20678,N_23826);
nor UO_2117 (O_2117,N_22371,N_22011);
xor UO_2118 (O_2118,N_22266,N_21517);
nand UO_2119 (O_2119,N_21453,N_20543);
and UO_2120 (O_2120,N_20910,N_20141);
or UO_2121 (O_2121,N_22045,N_23048);
nor UO_2122 (O_2122,N_20276,N_23738);
xnor UO_2123 (O_2123,N_22928,N_23993);
nand UO_2124 (O_2124,N_24777,N_23102);
xnor UO_2125 (O_2125,N_24083,N_21980);
nand UO_2126 (O_2126,N_23442,N_24894);
and UO_2127 (O_2127,N_24043,N_22644);
nand UO_2128 (O_2128,N_24583,N_22132);
and UO_2129 (O_2129,N_24957,N_23754);
nand UO_2130 (O_2130,N_21590,N_22702);
nand UO_2131 (O_2131,N_21637,N_20199);
nand UO_2132 (O_2132,N_24311,N_21021);
xor UO_2133 (O_2133,N_20013,N_21964);
nor UO_2134 (O_2134,N_23716,N_22616);
nor UO_2135 (O_2135,N_21212,N_20983);
xnor UO_2136 (O_2136,N_23527,N_20152);
nor UO_2137 (O_2137,N_20354,N_22615);
or UO_2138 (O_2138,N_21379,N_23650);
nor UO_2139 (O_2139,N_23393,N_23991);
and UO_2140 (O_2140,N_22703,N_20111);
nand UO_2141 (O_2141,N_20237,N_24333);
xor UO_2142 (O_2142,N_24715,N_22363);
xnor UO_2143 (O_2143,N_20382,N_23087);
nand UO_2144 (O_2144,N_21016,N_21848);
or UO_2145 (O_2145,N_20475,N_21151);
and UO_2146 (O_2146,N_21566,N_23044);
xnor UO_2147 (O_2147,N_24355,N_20922);
or UO_2148 (O_2148,N_20047,N_24154);
nand UO_2149 (O_2149,N_22353,N_22317);
xor UO_2150 (O_2150,N_23129,N_21561);
or UO_2151 (O_2151,N_20408,N_23427);
nor UO_2152 (O_2152,N_24123,N_21180);
and UO_2153 (O_2153,N_20346,N_20953);
nor UO_2154 (O_2154,N_24298,N_20831);
xor UO_2155 (O_2155,N_23091,N_22167);
nand UO_2156 (O_2156,N_20501,N_22340);
nor UO_2157 (O_2157,N_23962,N_22514);
nor UO_2158 (O_2158,N_21296,N_20966);
and UO_2159 (O_2159,N_22345,N_21916);
nand UO_2160 (O_2160,N_22773,N_20039);
nand UO_2161 (O_2161,N_24705,N_24299);
or UO_2162 (O_2162,N_22875,N_23061);
and UO_2163 (O_2163,N_21907,N_21881);
nand UO_2164 (O_2164,N_20344,N_24937);
and UO_2165 (O_2165,N_21859,N_24138);
xnor UO_2166 (O_2166,N_22684,N_23011);
nand UO_2167 (O_2167,N_24261,N_23341);
xor UO_2168 (O_2168,N_20099,N_23891);
nor UO_2169 (O_2169,N_21982,N_21864);
and UO_2170 (O_2170,N_23629,N_22562);
and UO_2171 (O_2171,N_20643,N_24402);
xor UO_2172 (O_2172,N_21764,N_23974);
nor UO_2173 (O_2173,N_20586,N_23163);
xor UO_2174 (O_2174,N_21929,N_24755);
or UO_2175 (O_2175,N_20257,N_24377);
nand UO_2176 (O_2176,N_24322,N_21326);
or UO_2177 (O_2177,N_20422,N_20496);
nor UO_2178 (O_2178,N_22892,N_22320);
or UO_2179 (O_2179,N_22037,N_21316);
and UO_2180 (O_2180,N_24250,N_22040);
and UO_2181 (O_2181,N_20178,N_21347);
and UO_2182 (O_2182,N_20399,N_22723);
or UO_2183 (O_2183,N_21066,N_24732);
or UO_2184 (O_2184,N_21562,N_21586);
and UO_2185 (O_2185,N_21428,N_21422);
nand UO_2186 (O_2186,N_23868,N_22500);
or UO_2187 (O_2187,N_22725,N_22497);
nor UO_2188 (O_2188,N_24010,N_23474);
nor UO_2189 (O_2189,N_24781,N_20314);
nor UO_2190 (O_2190,N_24089,N_20901);
and UO_2191 (O_2191,N_22173,N_22293);
xor UO_2192 (O_2192,N_20216,N_20102);
and UO_2193 (O_2193,N_21902,N_20454);
xnor UO_2194 (O_2194,N_20805,N_22693);
and UO_2195 (O_2195,N_21807,N_22252);
nor UO_2196 (O_2196,N_21020,N_23027);
xnor UO_2197 (O_2197,N_24520,N_21177);
or UO_2198 (O_2198,N_20841,N_21077);
or UO_2199 (O_2199,N_23967,N_23160);
nand UO_2200 (O_2200,N_22325,N_20373);
or UO_2201 (O_2201,N_24927,N_21214);
or UO_2202 (O_2202,N_23902,N_24353);
and UO_2203 (O_2203,N_22245,N_22739);
nor UO_2204 (O_2204,N_21646,N_22292);
and UO_2205 (O_2205,N_21330,N_24782);
nor UO_2206 (O_2206,N_23190,N_22909);
xnor UO_2207 (O_2207,N_24930,N_23248);
nand UO_2208 (O_2208,N_23992,N_22162);
xor UO_2209 (O_2209,N_24266,N_23073);
xnor UO_2210 (O_2210,N_22400,N_21267);
and UO_2211 (O_2211,N_20348,N_23032);
and UO_2212 (O_2212,N_20981,N_21521);
xor UO_2213 (O_2213,N_22130,N_20760);
and UO_2214 (O_2214,N_22128,N_22940);
nor UO_2215 (O_2215,N_23803,N_20515);
nor UO_2216 (O_2216,N_23534,N_22439);
nor UO_2217 (O_2217,N_21771,N_24543);
and UO_2218 (O_2218,N_21719,N_24764);
and UO_2219 (O_2219,N_21655,N_22467);
nand UO_2220 (O_2220,N_21235,N_21475);
xnor UO_2221 (O_2221,N_24567,N_22120);
nor UO_2222 (O_2222,N_24435,N_20982);
or UO_2223 (O_2223,N_22821,N_22026);
nand UO_2224 (O_2224,N_20347,N_20601);
nand UO_2225 (O_2225,N_22323,N_24055);
nor UO_2226 (O_2226,N_22290,N_24338);
or UO_2227 (O_2227,N_22868,N_23997);
nand UO_2228 (O_2228,N_24664,N_20799);
nand UO_2229 (O_2229,N_20020,N_24800);
or UO_2230 (O_2230,N_20742,N_20950);
and UO_2231 (O_2231,N_23267,N_23921);
nand UO_2232 (O_2232,N_21090,N_20487);
nand UO_2233 (O_2233,N_21927,N_21282);
nor UO_2234 (O_2234,N_24861,N_21407);
nor UO_2235 (O_2235,N_21751,N_20096);
nand UO_2236 (O_2236,N_22080,N_23144);
nand UO_2237 (O_2237,N_22369,N_21408);
nor UO_2238 (O_2238,N_23409,N_24776);
or UO_2239 (O_2239,N_22061,N_21519);
nor UO_2240 (O_2240,N_21076,N_24944);
nor UO_2241 (O_2241,N_22483,N_24094);
and UO_2242 (O_2242,N_20325,N_20837);
and UO_2243 (O_2243,N_21585,N_22505);
or UO_2244 (O_2244,N_21046,N_21350);
nand UO_2245 (O_2245,N_24454,N_24886);
xnor UO_2246 (O_2246,N_20523,N_22477);
nand UO_2247 (O_2247,N_21684,N_22246);
or UO_2248 (O_2248,N_24272,N_22233);
nand UO_2249 (O_2249,N_23243,N_22846);
nand UO_2250 (O_2250,N_20362,N_21047);
xnor UO_2251 (O_2251,N_22125,N_20129);
nor UO_2252 (O_2252,N_23332,N_23792);
or UO_2253 (O_2253,N_24838,N_21132);
or UO_2254 (O_2254,N_20417,N_20539);
or UO_2255 (O_2255,N_21286,N_21970);
xnor UO_2256 (O_2256,N_24515,N_24502);
nor UO_2257 (O_2257,N_22778,N_24200);
and UO_2258 (O_2258,N_22955,N_21950);
or UO_2259 (O_2259,N_22887,N_23031);
nand UO_2260 (O_2260,N_21720,N_20008);
nor UO_2261 (O_2261,N_21551,N_21173);
or UO_2262 (O_2262,N_24952,N_20063);
xnor UO_2263 (O_2263,N_21817,N_23741);
or UO_2264 (O_2264,N_24278,N_22144);
and UO_2265 (O_2265,N_22104,N_22985);
xnor UO_2266 (O_2266,N_22396,N_20602);
nor UO_2267 (O_2267,N_20124,N_20112);
xor UO_2268 (O_2268,N_21012,N_24273);
nor UO_2269 (O_2269,N_23582,N_21378);
nand UO_2270 (O_2270,N_23284,N_23210);
nand UO_2271 (O_2271,N_20349,N_21161);
and UO_2272 (O_2272,N_21912,N_21482);
or UO_2273 (O_2273,N_21411,N_24949);
nand UO_2274 (O_2274,N_24246,N_21301);
xnor UO_2275 (O_2275,N_24292,N_20607);
nand UO_2276 (O_2276,N_21366,N_22486);
or UO_2277 (O_2277,N_22493,N_21361);
xor UO_2278 (O_2278,N_23151,N_22986);
and UO_2279 (O_2279,N_21861,N_21685);
or UO_2280 (O_2280,N_20353,N_23538);
nand UO_2281 (O_2281,N_21891,N_24812);
or UO_2282 (O_2282,N_22680,N_22174);
xor UO_2283 (O_2283,N_22099,N_21245);
nand UO_2284 (O_2284,N_21617,N_23699);
xnor UO_2285 (O_2285,N_23938,N_23404);
and UO_2286 (O_2286,N_20558,N_22824);
xor UO_2287 (O_2287,N_23555,N_20171);
nor UO_2288 (O_2288,N_22232,N_20828);
xor UO_2289 (O_2289,N_22932,N_24810);
nor UO_2290 (O_2290,N_23093,N_24573);
nor UO_2291 (O_2291,N_24114,N_21285);
xor UO_2292 (O_2292,N_20392,N_23009);
xnor UO_2293 (O_2293,N_21213,N_23377);
nand UO_2294 (O_2294,N_24953,N_23820);
xor UO_2295 (O_2295,N_22899,N_22546);
nor UO_2296 (O_2296,N_23227,N_20436);
xor UO_2297 (O_2297,N_20857,N_21175);
nand UO_2298 (O_2298,N_22367,N_21995);
xor UO_2299 (O_2299,N_21785,N_24534);
or UO_2300 (O_2300,N_24396,N_20456);
and UO_2301 (O_2301,N_24018,N_20250);
or UO_2302 (O_2302,N_23106,N_20083);
and UO_2303 (O_2303,N_23919,N_23581);
nor UO_2304 (O_2304,N_20629,N_22976);
or UO_2305 (O_2305,N_22097,N_23020);
and UO_2306 (O_2306,N_22566,N_22336);
nor UO_2307 (O_2307,N_22413,N_22409);
nand UO_2308 (O_2308,N_22247,N_24239);
xnor UO_2309 (O_2309,N_22832,N_24393);
or UO_2310 (O_2310,N_24707,N_20827);
nor UO_2311 (O_2311,N_21248,N_21758);
xnor UO_2312 (O_2312,N_23280,N_23057);
nand UO_2313 (O_2313,N_23945,N_24220);
xnor UO_2314 (O_2314,N_22433,N_20282);
nand UO_2315 (O_2315,N_20017,N_24357);
nand UO_2316 (O_2316,N_20400,N_24961);
and UO_2317 (O_2317,N_24645,N_23052);
nor UO_2318 (O_2318,N_20924,N_24097);
nor UO_2319 (O_2319,N_21306,N_21609);
or UO_2320 (O_2320,N_24004,N_20035);
nor UO_2321 (O_2321,N_24263,N_20917);
nor UO_2322 (O_2322,N_21259,N_23558);
or UO_2323 (O_2323,N_24529,N_22897);
or UO_2324 (O_2324,N_23800,N_23175);
nand UO_2325 (O_2325,N_22904,N_23547);
and UO_2326 (O_2326,N_24020,N_24403);
and UO_2327 (O_2327,N_24546,N_24765);
nor UO_2328 (O_2328,N_23261,N_24950);
xnor UO_2329 (O_2329,N_23141,N_24457);
xor UO_2330 (O_2330,N_20873,N_23982);
xnor UO_2331 (O_2331,N_21085,N_24622);
and UO_2332 (O_2332,N_20410,N_21531);
nand UO_2333 (O_2333,N_22748,N_20704);
and UO_2334 (O_2334,N_24252,N_20331);
or UO_2335 (O_2335,N_24548,N_20181);
xnor UO_2336 (O_2336,N_20916,N_21959);
or UO_2337 (O_2337,N_22136,N_21623);
xnor UO_2338 (O_2338,N_24872,N_21595);
and UO_2339 (O_2339,N_22968,N_22346);
nor UO_2340 (O_2340,N_23249,N_20566);
and UO_2341 (O_2341,N_20688,N_24095);
xor UO_2342 (O_2342,N_24878,N_21237);
nor UO_2343 (O_2343,N_23877,N_22988);
or UO_2344 (O_2344,N_21838,N_22313);
or UO_2345 (O_2345,N_22907,N_22407);
nand UO_2346 (O_2346,N_23015,N_21534);
nand UO_2347 (O_2347,N_23725,N_20270);
or UO_2348 (O_2348,N_22472,N_23621);
and UO_2349 (O_2349,N_20101,N_24923);
nor UO_2350 (O_2350,N_20130,N_20238);
and UO_2351 (O_2351,N_22564,N_22212);
and UO_2352 (O_2352,N_24358,N_24947);
and UO_2353 (O_2353,N_22265,N_22447);
xor UO_2354 (O_2354,N_22547,N_21877);
nand UO_2355 (O_2355,N_21946,N_22704);
nor UO_2356 (O_2356,N_20608,N_22300);
xnor UO_2357 (O_2357,N_22280,N_24510);
and UO_2358 (O_2358,N_23944,N_22752);
or UO_2359 (O_2359,N_21146,N_20895);
or UO_2360 (O_2360,N_20510,N_20157);
nor UO_2361 (O_2361,N_23150,N_24857);
nand UO_2362 (O_2362,N_24716,N_22656);
or UO_2363 (O_2363,N_23140,N_22066);
xor UO_2364 (O_2364,N_21667,N_21605);
nor UO_2365 (O_2365,N_23981,N_20027);
xnor UO_2366 (O_2366,N_24206,N_22253);
and UO_2367 (O_2367,N_20326,N_24300);
nand UO_2368 (O_2368,N_23773,N_22910);
and UO_2369 (O_2369,N_21991,N_24215);
or UO_2370 (O_2370,N_24835,N_23056);
or UO_2371 (O_2371,N_22196,N_22718);
and UO_2372 (O_2372,N_21315,N_21931);
or UO_2373 (O_2373,N_21795,N_24960);
xor UO_2374 (O_2374,N_20905,N_20839);
nand UO_2375 (O_2375,N_21990,N_23737);
xnor UO_2376 (O_2376,N_23782,N_23946);
xnor UO_2377 (O_2377,N_24582,N_21537);
nor UO_2378 (O_2378,N_24030,N_23115);
xnor UO_2379 (O_2379,N_22808,N_24105);
nand UO_2380 (O_2380,N_20514,N_23417);
xnor UO_2381 (O_2381,N_24533,N_23896);
nor UO_2382 (O_2382,N_21125,N_24915);
xor UO_2383 (O_2383,N_24547,N_23535);
nand UO_2384 (O_2384,N_23495,N_20327);
nor UO_2385 (O_2385,N_20822,N_24324);
nor UO_2386 (O_2386,N_21808,N_21653);
nor UO_2387 (O_2387,N_23998,N_22450);
nand UO_2388 (O_2388,N_20599,N_21393);
nor UO_2389 (O_2389,N_23194,N_24650);
nor UO_2390 (O_2390,N_21264,N_22183);
or UO_2391 (O_2391,N_24733,N_23865);
xor UO_2392 (O_2392,N_22727,N_22478);
nand UO_2393 (O_2393,N_24746,N_21444);
xor UO_2394 (O_2394,N_23680,N_24287);
or UO_2395 (O_2395,N_24814,N_20069);
and UO_2396 (O_2396,N_22670,N_24388);
nand UO_2397 (O_2397,N_23381,N_22843);
nand UO_2398 (O_2398,N_22075,N_20244);
nand UO_2399 (O_2399,N_21887,N_23137);
nor UO_2400 (O_2400,N_20021,N_23343);
nor UO_2401 (O_2401,N_22951,N_20064);
or UO_2402 (O_2402,N_22312,N_22385);
xnor UO_2403 (O_2403,N_24175,N_23380);
nand UO_2404 (O_2404,N_22647,N_22731);
nor UO_2405 (O_2405,N_20775,N_23250);
nand UO_2406 (O_2406,N_20339,N_22077);
or UO_2407 (O_2407,N_24612,N_24748);
xor UO_2408 (O_2408,N_21339,N_20551);
or UO_2409 (O_2409,N_22767,N_21791);
nor UO_2410 (O_2410,N_22272,N_20060);
nand UO_2411 (O_2411,N_23554,N_24037);
or UO_2412 (O_2412,N_24212,N_20443);
nor UO_2413 (O_2413,N_23465,N_22565);
xnor UO_2414 (O_2414,N_23904,N_21055);
nand UO_2415 (O_2415,N_20676,N_21030);
nand UO_2416 (O_2416,N_23986,N_22591);
xor UO_2417 (O_2417,N_24339,N_22083);
and UO_2418 (O_2418,N_24525,N_22639);
and UO_2419 (O_2419,N_21128,N_24015);
or UO_2420 (O_2420,N_23336,N_22474);
xnor UO_2421 (O_2421,N_24997,N_20381);
nand UO_2422 (O_2422,N_21533,N_20776);
and UO_2423 (O_2423,N_22529,N_24832);
and UO_2424 (O_2424,N_23634,N_22341);
xor UO_2425 (O_2425,N_23700,N_23719);
or UO_2426 (O_2426,N_21119,N_24464);
nor UO_2427 (O_2427,N_21078,N_24026);
nand UO_2428 (O_2428,N_24293,N_20131);
xnor UO_2429 (O_2429,N_20450,N_24996);
xor UO_2430 (O_2430,N_22395,N_23301);
and UO_2431 (O_2431,N_21017,N_24545);
or UO_2432 (O_2432,N_21560,N_24808);
nand UO_2433 (O_2433,N_22803,N_21870);
and UO_2434 (O_2434,N_22151,N_20961);
or UO_2435 (O_2435,N_24608,N_23295);
and UO_2436 (O_2436,N_20904,N_23142);
nor UO_2437 (O_2437,N_22724,N_24499);
nand UO_2438 (O_2438,N_21106,N_23779);
nand UO_2439 (O_2439,N_22828,N_24452);
xnor UO_2440 (O_2440,N_21230,N_23225);
and UO_2441 (O_2441,N_24646,N_22047);
and UO_2442 (O_2442,N_23604,N_24460);
nand UO_2443 (O_2443,N_20990,N_24171);
nand UO_2444 (O_2444,N_20858,N_22243);
and UO_2445 (O_2445,N_23539,N_20938);
xnor UO_2446 (O_2446,N_22103,N_23119);
nor UO_2447 (O_2447,N_22701,N_23565);
nor UO_2448 (O_2448,N_23564,N_21065);
or UO_2449 (O_2449,N_23957,N_23724);
nor UO_2450 (O_2450,N_24306,N_24310);
nor UO_2451 (O_2451,N_24599,N_20930);
nand UO_2452 (O_2452,N_24627,N_24811);
and UO_2453 (O_2453,N_23542,N_21736);
nor UO_2454 (O_2454,N_24992,N_24466);
or UO_2455 (O_2455,N_24557,N_22574);
xnor UO_2456 (O_2456,N_20482,N_20151);
and UO_2457 (O_2457,N_20980,N_24110);
nor UO_2458 (O_2458,N_22024,N_22787);
nor UO_2459 (O_2459,N_23145,N_23673);
or UO_2460 (O_2460,N_24928,N_24192);
or UO_2461 (O_2461,N_24218,N_21375);
and UO_2462 (O_2462,N_21001,N_23575);
nor UO_2463 (O_2463,N_24188,N_24503);
nor UO_2464 (O_2464,N_23544,N_20722);
and UO_2465 (O_2465,N_20303,N_21536);
or UO_2466 (O_2466,N_21010,N_23183);
nor UO_2467 (O_2467,N_22495,N_24955);
nor UO_2468 (O_2468,N_20214,N_24420);
or UO_2469 (O_2469,N_22764,N_23130);
or UO_2470 (O_2470,N_24784,N_23156);
nor UO_2471 (O_2471,N_21039,N_24917);
nor UO_2472 (O_2472,N_23298,N_22987);
or UO_2473 (O_2473,N_20719,N_22056);
xnor UO_2474 (O_2474,N_23788,N_22378);
or UO_2475 (O_2475,N_24107,N_22754);
or UO_2476 (O_2476,N_21351,N_22538);
and UO_2477 (O_2477,N_22350,N_24541);
nor UO_2478 (O_2478,N_22179,N_22468);
nor UO_2479 (O_2479,N_23325,N_21321);
xor UO_2480 (O_2480,N_23709,N_22039);
nand UO_2481 (O_2481,N_24066,N_23418);
and UO_2482 (O_2482,N_21290,N_22116);
or UO_2483 (O_2483,N_24566,N_21277);
nor UO_2484 (O_2484,N_21746,N_23732);
or UO_2485 (O_2485,N_21508,N_22662);
or UO_2486 (O_2486,N_24084,N_22267);
or UO_2487 (O_2487,N_23746,N_24003);
nor UO_2488 (O_2488,N_21554,N_22527);
nor UO_2489 (O_2489,N_20302,N_22190);
nand UO_2490 (O_2490,N_23548,N_20034);
nor UO_2491 (O_2491,N_24276,N_22577);
nor UO_2492 (O_2492,N_24173,N_23252);
xnor UO_2493 (O_2493,N_23846,N_22830);
nand UO_2494 (O_2494,N_21261,N_20520);
xnor UO_2495 (O_2495,N_23432,N_22492);
and UO_2496 (O_2496,N_23687,N_23623);
and UO_2497 (O_2497,N_20815,N_20001);
or UO_2498 (O_2498,N_22519,N_24604);
or UO_2499 (O_2499,N_20363,N_21769);
nor UO_2500 (O_2500,N_23807,N_22829);
and UO_2501 (O_2501,N_22213,N_23959);
and UO_2502 (O_2502,N_20139,N_21267);
and UO_2503 (O_2503,N_24914,N_24293);
and UO_2504 (O_2504,N_24455,N_22849);
xnor UO_2505 (O_2505,N_21291,N_21646);
and UO_2506 (O_2506,N_24885,N_20311);
and UO_2507 (O_2507,N_23349,N_23427);
nand UO_2508 (O_2508,N_21343,N_22252);
nand UO_2509 (O_2509,N_24739,N_23055);
and UO_2510 (O_2510,N_21462,N_22783);
nor UO_2511 (O_2511,N_20372,N_22577);
and UO_2512 (O_2512,N_23682,N_22438);
nand UO_2513 (O_2513,N_23581,N_23658);
and UO_2514 (O_2514,N_21487,N_21929);
nand UO_2515 (O_2515,N_22686,N_24703);
nor UO_2516 (O_2516,N_20243,N_23128);
or UO_2517 (O_2517,N_24282,N_21979);
nor UO_2518 (O_2518,N_21936,N_24467);
xnor UO_2519 (O_2519,N_24204,N_20524);
xnor UO_2520 (O_2520,N_23711,N_22155);
nor UO_2521 (O_2521,N_24814,N_22786);
and UO_2522 (O_2522,N_21323,N_21433);
or UO_2523 (O_2523,N_23240,N_20508);
nor UO_2524 (O_2524,N_22034,N_23895);
xor UO_2525 (O_2525,N_21264,N_23033);
nand UO_2526 (O_2526,N_20266,N_22483);
nand UO_2527 (O_2527,N_23606,N_21005);
nor UO_2528 (O_2528,N_22434,N_23127);
xnor UO_2529 (O_2529,N_23407,N_21914);
or UO_2530 (O_2530,N_22352,N_22121);
nor UO_2531 (O_2531,N_20040,N_21029);
and UO_2532 (O_2532,N_22962,N_21817);
or UO_2533 (O_2533,N_22142,N_24573);
nor UO_2534 (O_2534,N_20342,N_20409);
or UO_2535 (O_2535,N_21916,N_23807);
and UO_2536 (O_2536,N_22683,N_20546);
xor UO_2537 (O_2537,N_20833,N_24621);
nand UO_2538 (O_2538,N_24427,N_21969);
or UO_2539 (O_2539,N_23929,N_23396);
nor UO_2540 (O_2540,N_21910,N_23375);
nand UO_2541 (O_2541,N_22112,N_23617);
nand UO_2542 (O_2542,N_23794,N_23928);
or UO_2543 (O_2543,N_24376,N_20562);
nand UO_2544 (O_2544,N_24790,N_23817);
or UO_2545 (O_2545,N_23552,N_24451);
or UO_2546 (O_2546,N_20795,N_22984);
or UO_2547 (O_2547,N_21065,N_21598);
nand UO_2548 (O_2548,N_23472,N_22418);
nor UO_2549 (O_2549,N_20108,N_20605);
or UO_2550 (O_2550,N_23036,N_23534);
xnor UO_2551 (O_2551,N_22807,N_22987);
and UO_2552 (O_2552,N_21487,N_24284);
nor UO_2553 (O_2553,N_20138,N_23605);
and UO_2554 (O_2554,N_24107,N_20362);
xnor UO_2555 (O_2555,N_22670,N_21131);
nor UO_2556 (O_2556,N_23277,N_22371);
nor UO_2557 (O_2557,N_22196,N_24157);
and UO_2558 (O_2558,N_24799,N_21685);
nand UO_2559 (O_2559,N_24174,N_22447);
xnor UO_2560 (O_2560,N_23438,N_24501);
nor UO_2561 (O_2561,N_21509,N_20000);
nand UO_2562 (O_2562,N_20817,N_20766);
or UO_2563 (O_2563,N_20457,N_20204);
or UO_2564 (O_2564,N_20685,N_23600);
nand UO_2565 (O_2565,N_22412,N_22907);
or UO_2566 (O_2566,N_22807,N_24419);
nor UO_2567 (O_2567,N_23499,N_20867);
and UO_2568 (O_2568,N_22361,N_20612);
xnor UO_2569 (O_2569,N_21439,N_20632);
or UO_2570 (O_2570,N_23342,N_20823);
nor UO_2571 (O_2571,N_23467,N_23534);
nand UO_2572 (O_2572,N_24451,N_20243);
nor UO_2573 (O_2573,N_21380,N_20544);
nor UO_2574 (O_2574,N_20272,N_22465);
nor UO_2575 (O_2575,N_21227,N_23643);
or UO_2576 (O_2576,N_23844,N_20101);
and UO_2577 (O_2577,N_21032,N_20204);
xor UO_2578 (O_2578,N_24950,N_21065);
and UO_2579 (O_2579,N_20642,N_20037);
nand UO_2580 (O_2580,N_20840,N_23153);
xnor UO_2581 (O_2581,N_24519,N_20079);
nor UO_2582 (O_2582,N_24825,N_21264);
nand UO_2583 (O_2583,N_24453,N_24048);
nor UO_2584 (O_2584,N_23660,N_20578);
and UO_2585 (O_2585,N_24728,N_22360);
or UO_2586 (O_2586,N_20820,N_22435);
nor UO_2587 (O_2587,N_21315,N_23997);
nor UO_2588 (O_2588,N_22750,N_24118);
xnor UO_2589 (O_2589,N_20738,N_24235);
or UO_2590 (O_2590,N_23986,N_24990);
nand UO_2591 (O_2591,N_23125,N_20808);
nor UO_2592 (O_2592,N_21079,N_22465);
nor UO_2593 (O_2593,N_20320,N_21052);
nor UO_2594 (O_2594,N_24652,N_20391);
or UO_2595 (O_2595,N_24214,N_23144);
nand UO_2596 (O_2596,N_24176,N_21063);
nor UO_2597 (O_2597,N_22184,N_22746);
or UO_2598 (O_2598,N_24850,N_21903);
nor UO_2599 (O_2599,N_20120,N_23312);
or UO_2600 (O_2600,N_24744,N_24432);
or UO_2601 (O_2601,N_20683,N_24389);
nor UO_2602 (O_2602,N_23261,N_24307);
or UO_2603 (O_2603,N_21966,N_23443);
and UO_2604 (O_2604,N_23070,N_23409);
and UO_2605 (O_2605,N_20156,N_20516);
nor UO_2606 (O_2606,N_23576,N_22655);
or UO_2607 (O_2607,N_21710,N_22951);
or UO_2608 (O_2608,N_22779,N_23921);
xor UO_2609 (O_2609,N_22128,N_22168);
nor UO_2610 (O_2610,N_20273,N_22144);
nand UO_2611 (O_2611,N_22161,N_20024);
or UO_2612 (O_2612,N_23255,N_24805);
or UO_2613 (O_2613,N_20840,N_23126);
or UO_2614 (O_2614,N_20456,N_20116);
nand UO_2615 (O_2615,N_21915,N_24667);
nand UO_2616 (O_2616,N_20394,N_20780);
xnor UO_2617 (O_2617,N_21028,N_23094);
nand UO_2618 (O_2618,N_23922,N_20516);
xnor UO_2619 (O_2619,N_20632,N_24411);
nor UO_2620 (O_2620,N_21918,N_24467);
nor UO_2621 (O_2621,N_24523,N_22616);
nand UO_2622 (O_2622,N_20008,N_23927);
and UO_2623 (O_2623,N_23330,N_23363);
xnor UO_2624 (O_2624,N_21653,N_24739);
nor UO_2625 (O_2625,N_24877,N_24512);
nand UO_2626 (O_2626,N_20540,N_22024);
nor UO_2627 (O_2627,N_24212,N_24153);
nor UO_2628 (O_2628,N_20558,N_21381);
and UO_2629 (O_2629,N_21717,N_24170);
or UO_2630 (O_2630,N_22759,N_20880);
nand UO_2631 (O_2631,N_20758,N_20085);
nand UO_2632 (O_2632,N_22252,N_20762);
nand UO_2633 (O_2633,N_24738,N_21935);
and UO_2634 (O_2634,N_22002,N_20199);
and UO_2635 (O_2635,N_24044,N_22825);
or UO_2636 (O_2636,N_21954,N_24820);
xor UO_2637 (O_2637,N_20705,N_24133);
or UO_2638 (O_2638,N_24903,N_22953);
nor UO_2639 (O_2639,N_20863,N_23900);
and UO_2640 (O_2640,N_21206,N_21621);
xnor UO_2641 (O_2641,N_22749,N_22735);
xnor UO_2642 (O_2642,N_23496,N_20336);
xor UO_2643 (O_2643,N_20519,N_23945);
or UO_2644 (O_2644,N_21708,N_23085);
or UO_2645 (O_2645,N_20672,N_22538);
nor UO_2646 (O_2646,N_22269,N_20922);
nor UO_2647 (O_2647,N_23423,N_22930);
nor UO_2648 (O_2648,N_22757,N_22987);
xnor UO_2649 (O_2649,N_21180,N_24153);
xor UO_2650 (O_2650,N_20705,N_24681);
nand UO_2651 (O_2651,N_24597,N_24592);
nor UO_2652 (O_2652,N_21910,N_20788);
nand UO_2653 (O_2653,N_24242,N_22298);
or UO_2654 (O_2654,N_23652,N_23580);
xnor UO_2655 (O_2655,N_22359,N_21976);
nand UO_2656 (O_2656,N_23495,N_20495);
nand UO_2657 (O_2657,N_22730,N_20360);
or UO_2658 (O_2658,N_23022,N_22555);
or UO_2659 (O_2659,N_21241,N_24225);
xnor UO_2660 (O_2660,N_20212,N_24661);
nand UO_2661 (O_2661,N_20971,N_21953);
xnor UO_2662 (O_2662,N_22762,N_22732);
nand UO_2663 (O_2663,N_23038,N_24893);
and UO_2664 (O_2664,N_23050,N_22945);
and UO_2665 (O_2665,N_23941,N_21763);
nor UO_2666 (O_2666,N_20085,N_21369);
nor UO_2667 (O_2667,N_23468,N_24765);
nor UO_2668 (O_2668,N_20129,N_24342);
and UO_2669 (O_2669,N_24787,N_23822);
or UO_2670 (O_2670,N_24633,N_23199);
nand UO_2671 (O_2671,N_22891,N_22700);
nor UO_2672 (O_2672,N_22407,N_21551);
nand UO_2673 (O_2673,N_21518,N_23131);
or UO_2674 (O_2674,N_20342,N_22031);
and UO_2675 (O_2675,N_23742,N_22739);
nor UO_2676 (O_2676,N_23132,N_24714);
nor UO_2677 (O_2677,N_23477,N_21397);
nand UO_2678 (O_2678,N_20444,N_21106);
nand UO_2679 (O_2679,N_23182,N_22135);
xnor UO_2680 (O_2680,N_23492,N_20395);
nand UO_2681 (O_2681,N_21855,N_24847);
and UO_2682 (O_2682,N_24192,N_20767);
or UO_2683 (O_2683,N_24721,N_20627);
nor UO_2684 (O_2684,N_23117,N_23751);
nand UO_2685 (O_2685,N_21998,N_24150);
nor UO_2686 (O_2686,N_20111,N_23664);
and UO_2687 (O_2687,N_20384,N_21715);
xnor UO_2688 (O_2688,N_22066,N_24577);
or UO_2689 (O_2689,N_23155,N_24955);
xnor UO_2690 (O_2690,N_20430,N_20635);
xor UO_2691 (O_2691,N_24703,N_20400);
nand UO_2692 (O_2692,N_22898,N_20328);
xor UO_2693 (O_2693,N_23347,N_23865);
xor UO_2694 (O_2694,N_22528,N_23157);
xnor UO_2695 (O_2695,N_23468,N_22343);
nand UO_2696 (O_2696,N_21872,N_20542);
xnor UO_2697 (O_2697,N_24982,N_24418);
nand UO_2698 (O_2698,N_21189,N_23268);
nor UO_2699 (O_2699,N_22350,N_22970);
nor UO_2700 (O_2700,N_21729,N_21818);
or UO_2701 (O_2701,N_22556,N_23469);
nor UO_2702 (O_2702,N_23191,N_24185);
xor UO_2703 (O_2703,N_20515,N_21287);
nand UO_2704 (O_2704,N_22830,N_20682);
nor UO_2705 (O_2705,N_24729,N_22945);
xor UO_2706 (O_2706,N_22429,N_21057);
nand UO_2707 (O_2707,N_22719,N_23508);
nor UO_2708 (O_2708,N_23432,N_24161);
and UO_2709 (O_2709,N_24727,N_20747);
or UO_2710 (O_2710,N_24205,N_22286);
and UO_2711 (O_2711,N_23383,N_21349);
nand UO_2712 (O_2712,N_20922,N_23945);
or UO_2713 (O_2713,N_23626,N_23214);
xnor UO_2714 (O_2714,N_22139,N_22890);
and UO_2715 (O_2715,N_23588,N_20449);
xor UO_2716 (O_2716,N_21147,N_23466);
or UO_2717 (O_2717,N_24298,N_24512);
xor UO_2718 (O_2718,N_23793,N_24143);
and UO_2719 (O_2719,N_22934,N_20985);
or UO_2720 (O_2720,N_24984,N_24316);
and UO_2721 (O_2721,N_23784,N_21389);
and UO_2722 (O_2722,N_24063,N_21058);
nor UO_2723 (O_2723,N_24137,N_22241);
nand UO_2724 (O_2724,N_21831,N_21402);
xor UO_2725 (O_2725,N_23790,N_24964);
nor UO_2726 (O_2726,N_23214,N_22486);
xor UO_2727 (O_2727,N_20436,N_20169);
or UO_2728 (O_2728,N_21855,N_21523);
nor UO_2729 (O_2729,N_21367,N_23256);
xor UO_2730 (O_2730,N_20841,N_23138);
or UO_2731 (O_2731,N_22960,N_21598);
and UO_2732 (O_2732,N_24584,N_21118);
nand UO_2733 (O_2733,N_24270,N_22830);
nor UO_2734 (O_2734,N_20789,N_20440);
nand UO_2735 (O_2735,N_23557,N_20478);
and UO_2736 (O_2736,N_24369,N_24589);
and UO_2737 (O_2737,N_24585,N_20913);
xor UO_2738 (O_2738,N_24121,N_22495);
nor UO_2739 (O_2739,N_22153,N_23321);
nor UO_2740 (O_2740,N_24069,N_21321);
nor UO_2741 (O_2741,N_20557,N_20053);
xor UO_2742 (O_2742,N_20976,N_21558);
or UO_2743 (O_2743,N_22670,N_23598);
xnor UO_2744 (O_2744,N_24845,N_22369);
nand UO_2745 (O_2745,N_23465,N_24420);
xnor UO_2746 (O_2746,N_20032,N_22120);
or UO_2747 (O_2747,N_22899,N_21077);
nor UO_2748 (O_2748,N_24826,N_22978);
nor UO_2749 (O_2749,N_24134,N_22663);
and UO_2750 (O_2750,N_23618,N_24815);
nor UO_2751 (O_2751,N_21344,N_24290);
and UO_2752 (O_2752,N_21447,N_22211);
nand UO_2753 (O_2753,N_21033,N_20045);
nor UO_2754 (O_2754,N_20543,N_22367);
nand UO_2755 (O_2755,N_22955,N_23772);
and UO_2756 (O_2756,N_22713,N_20525);
or UO_2757 (O_2757,N_20179,N_24727);
or UO_2758 (O_2758,N_22079,N_22671);
and UO_2759 (O_2759,N_21481,N_23542);
xnor UO_2760 (O_2760,N_21946,N_21529);
nor UO_2761 (O_2761,N_23380,N_24353);
or UO_2762 (O_2762,N_22470,N_24474);
or UO_2763 (O_2763,N_24246,N_20363);
xor UO_2764 (O_2764,N_22192,N_22715);
and UO_2765 (O_2765,N_23196,N_22399);
and UO_2766 (O_2766,N_22475,N_21546);
nand UO_2767 (O_2767,N_20326,N_24948);
nor UO_2768 (O_2768,N_24490,N_22003);
and UO_2769 (O_2769,N_22319,N_22421);
xor UO_2770 (O_2770,N_20305,N_24650);
and UO_2771 (O_2771,N_21032,N_21056);
nor UO_2772 (O_2772,N_23996,N_23424);
or UO_2773 (O_2773,N_21729,N_22139);
and UO_2774 (O_2774,N_22891,N_22829);
nand UO_2775 (O_2775,N_21381,N_20848);
or UO_2776 (O_2776,N_23899,N_22812);
and UO_2777 (O_2777,N_22607,N_21892);
nand UO_2778 (O_2778,N_20350,N_23860);
or UO_2779 (O_2779,N_22326,N_23171);
nand UO_2780 (O_2780,N_24050,N_24165);
or UO_2781 (O_2781,N_23616,N_20230);
nand UO_2782 (O_2782,N_20805,N_20557);
nor UO_2783 (O_2783,N_20916,N_24955);
xnor UO_2784 (O_2784,N_24954,N_24719);
or UO_2785 (O_2785,N_23634,N_21273);
xnor UO_2786 (O_2786,N_22760,N_24944);
nor UO_2787 (O_2787,N_20273,N_23110);
or UO_2788 (O_2788,N_23839,N_21502);
or UO_2789 (O_2789,N_23512,N_21346);
or UO_2790 (O_2790,N_22022,N_24591);
nand UO_2791 (O_2791,N_24763,N_21158);
or UO_2792 (O_2792,N_23810,N_22283);
nand UO_2793 (O_2793,N_20471,N_20304);
nand UO_2794 (O_2794,N_21526,N_24423);
nand UO_2795 (O_2795,N_24752,N_24012);
or UO_2796 (O_2796,N_21973,N_23743);
or UO_2797 (O_2797,N_23012,N_22955);
nand UO_2798 (O_2798,N_21946,N_20342);
or UO_2799 (O_2799,N_22387,N_20767);
xor UO_2800 (O_2800,N_21362,N_24654);
nor UO_2801 (O_2801,N_22240,N_21355);
or UO_2802 (O_2802,N_21977,N_24144);
xor UO_2803 (O_2803,N_20245,N_22852);
and UO_2804 (O_2804,N_24271,N_22349);
or UO_2805 (O_2805,N_20657,N_23385);
xor UO_2806 (O_2806,N_20778,N_23250);
nand UO_2807 (O_2807,N_22882,N_24025);
and UO_2808 (O_2808,N_20653,N_21230);
or UO_2809 (O_2809,N_20425,N_23555);
nor UO_2810 (O_2810,N_21674,N_22427);
or UO_2811 (O_2811,N_22553,N_22710);
xnor UO_2812 (O_2812,N_23803,N_20179);
nand UO_2813 (O_2813,N_20777,N_20542);
xnor UO_2814 (O_2814,N_22057,N_22788);
and UO_2815 (O_2815,N_20965,N_23771);
and UO_2816 (O_2816,N_22022,N_23146);
or UO_2817 (O_2817,N_22352,N_22216);
xor UO_2818 (O_2818,N_20273,N_20508);
xnor UO_2819 (O_2819,N_22262,N_23128);
and UO_2820 (O_2820,N_21695,N_22906);
xor UO_2821 (O_2821,N_22319,N_23985);
nor UO_2822 (O_2822,N_20375,N_22758);
and UO_2823 (O_2823,N_21493,N_21954);
and UO_2824 (O_2824,N_23868,N_23824);
xor UO_2825 (O_2825,N_22699,N_23041);
and UO_2826 (O_2826,N_22319,N_24856);
nor UO_2827 (O_2827,N_21115,N_20947);
or UO_2828 (O_2828,N_20610,N_24583);
nand UO_2829 (O_2829,N_20409,N_21954);
nand UO_2830 (O_2830,N_21616,N_20838);
xnor UO_2831 (O_2831,N_23081,N_24353);
and UO_2832 (O_2832,N_22073,N_20556);
nand UO_2833 (O_2833,N_22182,N_21754);
nor UO_2834 (O_2834,N_24689,N_20493);
or UO_2835 (O_2835,N_23592,N_23208);
or UO_2836 (O_2836,N_24222,N_23377);
nor UO_2837 (O_2837,N_21163,N_22768);
nor UO_2838 (O_2838,N_24167,N_21865);
and UO_2839 (O_2839,N_21418,N_20270);
nand UO_2840 (O_2840,N_23085,N_20361);
and UO_2841 (O_2841,N_23267,N_24255);
nand UO_2842 (O_2842,N_23203,N_22882);
and UO_2843 (O_2843,N_21534,N_21875);
or UO_2844 (O_2844,N_21941,N_21641);
nand UO_2845 (O_2845,N_20425,N_22000);
nor UO_2846 (O_2846,N_24113,N_22290);
nor UO_2847 (O_2847,N_20218,N_23131);
or UO_2848 (O_2848,N_22190,N_22604);
nor UO_2849 (O_2849,N_22968,N_20611);
nor UO_2850 (O_2850,N_22395,N_22666);
or UO_2851 (O_2851,N_20960,N_20123);
xnor UO_2852 (O_2852,N_21678,N_24916);
xnor UO_2853 (O_2853,N_21658,N_24732);
nor UO_2854 (O_2854,N_22056,N_22253);
nand UO_2855 (O_2855,N_21270,N_24193);
or UO_2856 (O_2856,N_22590,N_20763);
and UO_2857 (O_2857,N_21990,N_21879);
nand UO_2858 (O_2858,N_20299,N_21703);
xnor UO_2859 (O_2859,N_24868,N_21828);
nand UO_2860 (O_2860,N_24869,N_23182);
xor UO_2861 (O_2861,N_24375,N_20119);
nor UO_2862 (O_2862,N_24718,N_21235);
nand UO_2863 (O_2863,N_21028,N_20301);
nor UO_2864 (O_2864,N_22717,N_22666);
nand UO_2865 (O_2865,N_23068,N_20243);
xor UO_2866 (O_2866,N_22572,N_20086);
xor UO_2867 (O_2867,N_23438,N_23435);
or UO_2868 (O_2868,N_22631,N_23773);
xnor UO_2869 (O_2869,N_21311,N_22099);
or UO_2870 (O_2870,N_20613,N_24186);
and UO_2871 (O_2871,N_20734,N_22030);
or UO_2872 (O_2872,N_22377,N_21821);
or UO_2873 (O_2873,N_21308,N_23083);
nand UO_2874 (O_2874,N_20457,N_21677);
or UO_2875 (O_2875,N_22034,N_20754);
nor UO_2876 (O_2876,N_23010,N_24915);
or UO_2877 (O_2877,N_24959,N_22546);
xnor UO_2878 (O_2878,N_24935,N_21807);
nor UO_2879 (O_2879,N_20001,N_24168);
or UO_2880 (O_2880,N_23319,N_22115);
xnor UO_2881 (O_2881,N_24961,N_21600);
nand UO_2882 (O_2882,N_22733,N_24233);
nor UO_2883 (O_2883,N_22151,N_24039);
nor UO_2884 (O_2884,N_24950,N_23722);
nand UO_2885 (O_2885,N_22243,N_21567);
and UO_2886 (O_2886,N_24445,N_24879);
xor UO_2887 (O_2887,N_20910,N_20633);
and UO_2888 (O_2888,N_21935,N_24886);
xor UO_2889 (O_2889,N_24124,N_21010);
or UO_2890 (O_2890,N_21189,N_22703);
xnor UO_2891 (O_2891,N_23012,N_21488);
nand UO_2892 (O_2892,N_24105,N_23983);
or UO_2893 (O_2893,N_24907,N_23252);
nor UO_2894 (O_2894,N_23872,N_22724);
and UO_2895 (O_2895,N_20392,N_21984);
nand UO_2896 (O_2896,N_22046,N_24577);
nand UO_2897 (O_2897,N_24951,N_22547);
xor UO_2898 (O_2898,N_23948,N_21404);
or UO_2899 (O_2899,N_20629,N_24763);
nor UO_2900 (O_2900,N_21029,N_22170);
and UO_2901 (O_2901,N_20175,N_22800);
nor UO_2902 (O_2902,N_22232,N_20943);
nand UO_2903 (O_2903,N_23963,N_24480);
xnor UO_2904 (O_2904,N_20550,N_20855);
or UO_2905 (O_2905,N_22980,N_21292);
nand UO_2906 (O_2906,N_20735,N_20190);
xor UO_2907 (O_2907,N_22565,N_24654);
or UO_2908 (O_2908,N_22390,N_24991);
or UO_2909 (O_2909,N_24336,N_23057);
or UO_2910 (O_2910,N_24999,N_20411);
or UO_2911 (O_2911,N_22803,N_22702);
nor UO_2912 (O_2912,N_23909,N_22559);
and UO_2913 (O_2913,N_20709,N_23785);
nor UO_2914 (O_2914,N_23162,N_24485);
or UO_2915 (O_2915,N_21256,N_20362);
or UO_2916 (O_2916,N_24014,N_21330);
xor UO_2917 (O_2917,N_20676,N_21723);
nand UO_2918 (O_2918,N_23660,N_23710);
nand UO_2919 (O_2919,N_21890,N_24554);
and UO_2920 (O_2920,N_21990,N_21706);
nand UO_2921 (O_2921,N_21075,N_23726);
nor UO_2922 (O_2922,N_24953,N_22553);
and UO_2923 (O_2923,N_21296,N_23775);
or UO_2924 (O_2924,N_23443,N_23280);
nand UO_2925 (O_2925,N_20327,N_22730);
nand UO_2926 (O_2926,N_23725,N_20051);
nor UO_2927 (O_2927,N_22415,N_21382);
and UO_2928 (O_2928,N_23932,N_22630);
and UO_2929 (O_2929,N_22757,N_24637);
or UO_2930 (O_2930,N_23148,N_23280);
or UO_2931 (O_2931,N_24748,N_23080);
xor UO_2932 (O_2932,N_21745,N_24914);
and UO_2933 (O_2933,N_23455,N_23609);
and UO_2934 (O_2934,N_24958,N_24678);
and UO_2935 (O_2935,N_20696,N_20946);
nor UO_2936 (O_2936,N_20717,N_23151);
nand UO_2937 (O_2937,N_20545,N_22572);
nand UO_2938 (O_2938,N_21867,N_20950);
nand UO_2939 (O_2939,N_20764,N_22464);
and UO_2940 (O_2940,N_23795,N_20158);
xor UO_2941 (O_2941,N_20239,N_22168);
nor UO_2942 (O_2942,N_23774,N_23765);
or UO_2943 (O_2943,N_24619,N_21865);
and UO_2944 (O_2944,N_21064,N_24734);
nor UO_2945 (O_2945,N_22208,N_24623);
xnor UO_2946 (O_2946,N_23273,N_23848);
xnor UO_2947 (O_2947,N_20743,N_24419);
nor UO_2948 (O_2948,N_23937,N_23391);
and UO_2949 (O_2949,N_22557,N_20475);
xor UO_2950 (O_2950,N_21863,N_23873);
nand UO_2951 (O_2951,N_20835,N_22608);
nor UO_2952 (O_2952,N_24741,N_23108);
xor UO_2953 (O_2953,N_22531,N_22280);
and UO_2954 (O_2954,N_21985,N_22581);
and UO_2955 (O_2955,N_21878,N_20427);
nor UO_2956 (O_2956,N_21597,N_22119);
nor UO_2957 (O_2957,N_22292,N_21521);
or UO_2958 (O_2958,N_21064,N_20906);
nand UO_2959 (O_2959,N_23250,N_20041);
nand UO_2960 (O_2960,N_23048,N_22907);
or UO_2961 (O_2961,N_24353,N_24166);
nor UO_2962 (O_2962,N_21512,N_23494);
nor UO_2963 (O_2963,N_20470,N_24284);
xnor UO_2964 (O_2964,N_23680,N_23838);
and UO_2965 (O_2965,N_23285,N_22459);
xor UO_2966 (O_2966,N_24324,N_23146);
nand UO_2967 (O_2967,N_20407,N_24686);
nor UO_2968 (O_2968,N_23463,N_22594);
or UO_2969 (O_2969,N_23911,N_23741);
and UO_2970 (O_2970,N_24155,N_24893);
xnor UO_2971 (O_2971,N_23460,N_20929);
and UO_2972 (O_2972,N_24790,N_21493);
nor UO_2973 (O_2973,N_21161,N_20291);
nor UO_2974 (O_2974,N_23484,N_24608);
nor UO_2975 (O_2975,N_22719,N_22151);
nor UO_2976 (O_2976,N_20823,N_21212);
xnor UO_2977 (O_2977,N_21595,N_21950);
nor UO_2978 (O_2978,N_21563,N_23475);
and UO_2979 (O_2979,N_21632,N_21758);
nand UO_2980 (O_2980,N_24989,N_23067);
and UO_2981 (O_2981,N_20269,N_22537);
nor UO_2982 (O_2982,N_23134,N_24775);
and UO_2983 (O_2983,N_21057,N_22564);
nor UO_2984 (O_2984,N_20399,N_21027);
and UO_2985 (O_2985,N_20475,N_22210);
and UO_2986 (O_2986,N_21954,N_23004);
xnor UO_2987 (O_2987,N_21429,N_20502);
xor UO_2988 (O_2988,N_21942,N_21914);
or UO_2989 (O_2989,N_23931,N_22421);
nor UO_2990 (O_2990,N_21520,N_22595);
xor UO_2991 (O_2991,N_24024,N_23791);
and UO_2992 (O_2992,N_20729,N_20663);
and UO_2993 (O_2993,N_21199,N_24826);
or UO_2994 (O_2994,N_24099,N_20679);
and UO_2995 (O_2995,N_21720,N_22404);
xor UO_2996 (O_2996,N_21626,N_23686);
or UO_2997 (O_2997,N_21861,N_24380);
nand UO_2998 (O_2998,N_21608,N_24040);
or UO_2999 (O_2999,N_20078,N_22239);
endmodule