module basic_3000_30000_3500_20_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
and U0 (N_0,In_1484,In_1669);
xor U1 (N_1,In_89,In_641);
or U2 (N_2,In_463,In_895);
xnor U3 (N_3,In_203,In_1564);
and U4 (N_4,In_2675,In_2353);
nor U5 (N_5,In_871,In_958);
nor U6 (N_6,In_468,In_2374);
nand U7 (N_7,In_2790,In_1984);
and U8 (N_8,In_883,In_113);
and U9 (N_9,In_1415,In_2034);
nand U10 (N_10,In_973,In_2513);
nand U11 (N_11,In_1418,In_1154);
nor U12 (N_12,In_1660,In_1218);
xor U13 (N_13,In_1659,In_1644);
or U14 (N_14,In_2398,In_1449);
nor U15 (N_15,In_1627,In_1972);
and U16 (N_16,In_1392,In_2476);
nor U17 (N_17,In_2424,In_111);
xor U18 (N_18,In_1251,In_1105);
nor U19 (N_19,In_1455,In_169);
xnor U20 (N_20,In_314,In_1720);
and U21 (N_21,In_1483,In_2433);
nor U22 (N_22,In_465,In_2597);
nand U23 (N_23,In_2651,In_818);
nand U24 (N_24,In_2735,In_2333);
nor U25 (N_25,In_699,In_758);
or U26 (N_26,In_1387,In_797);
and U27 (N_27,In_213,In_2257);
xor U28 (N_28,In_1638,In_2144);
or U29 (N_29,In_1945,In_2526);
and U30 (N_30,In_281,In_2452);
xnor U31 (N_31,In_832,In_2075);
nand U32 (N_32,In_2818,In_986);
and U33 (N_33,In_338,In_544);
or U34 (N_34,In_1709,In_2715);
nand U35 (N_35,In_1837,In_924);
or U36 (N_36,In_769,In_2888);
nand U37 (N_37,In_1268,In_1994);
and U38 (N_38,In_1839,In_1672);
nand U39 (N_39,In_1796,In_1464);
nand U40 (N_40,In_1042,In_1489);
and U41 (N_41,In_2755,In_2577);
and U42 (N_42,In_777,In_1577);
or U43 (N_43,In_1369,In_1857);
nand U44 (N_44,In_2509,In_2845);
xnor U45 (N_45,In_2935,In_917);
and U46 (N_46,In_1684,In_1211);
nand U47 (N_47,In_1277,In_2956);
xor U48 (N_48,In_370,In_40);
nand U49 (N_49,In_1469,In_342);
nor U50 (N_50,In_390,In_2140);
and U51 (N_51,In_1969,In_1616);
nor U52 (N_52,In_534,In_2861);
and U53 (N_53,In_1375,In_1540);
nor U54 (N_54,In_1257,In_1274);
or U55 (N_55,In_245,In_1704);
and U56 (N_56,In_2205,In_990);
or U57 (N_57,In_1065,In_2833);
and U58 (N_58,In_358,In_961);
nand U59 (N_59,In_2750,In_311);
or U60 (N_60,In_2302,In_2064);
nand U61 (N_61,In_1865,In_2278);
nor U62 (N_62,In_1031,In_2005);
and U63 (N_63,In_690,In_962);
nand U64 (N_64,In_2834,In_2732);
nand U65 (N_65,In_470,In_2434);
nand U66 (N_66,In_1447,In_1142);
xor U67 (N_67,In_2661,In_844);
nand U68 (N_68,In_603,In_2);
or U69 (N_69,In_762,In_1967);
nor U70 (N_70,In_1550,In_199);
nor U71 (N_71,In_400,In_2311);
xor U72 (N_72,In_2870,In_2060);
nand U73 (N_73,In_2958,In_964);
nand U74 (N_74,In_956,In_1498);
nor U75 (N_75,In_795,In_589);
nand U76 (N_76,In_656,In_1217);
nor U77 (N_77,In_195,In_989);
nand U78 (N_78,In_2373,In_549);
nand U79 (N_79,In_2377,In_664);
or U80 (N_80,In_524,In_200);
xnor U81 (N_81,In_2685,In_2237);
nor U82 (N_82,In_1604,In_343);
nand U83 (N_83,In_2281,In_2198);
or U84 (N_84,In_30,In_1781);
nor U85 (N_85,In_2020,In_2827);
or U86 (N_86,In_1853,In_409);
or U87 (N_87,In_673,In_318);
nand U88 (N_88,In_1408,In_2209);
and U89 (N_89,In_2017,In_2738);
xor U90 (N_90,In_253,In_2048);
and U91 (N_91,In_1301,In_136);
xor U92 (N_92,In_2025,In_2329);
xnor U93 (N_93,In_1683,In_437);
or U94 (N_94,In_263,In_750);
or U95 (N_95,In_76,In_2160);
nand U96 (N_96,In_237,In_2745);
nor U97 (N_97,In_1492,In_2059);
or U98 (N_98,In_886,In_2251);
xnor U99 (N_99,In_6,In_530);
and U100 (N_100,In_57,In_248);
nor U101 (N_101,In_2401,In_1917);
or U102 (N_102,In_2824,In_881);
or U103 (N_103,In_1749,In_1407);
xnor U104 (N_104,In_2915,In_1027);
or U105 (N_105,In_331,In_2306);
nand U106 (N_106,In_610,In_1478);
or U107 (N_107,In_1399,In_2904);
nor U108 (N_108,In_1735,In_2285);
nand U109 (N_109,In_596,In_693);
or U110 (N_110,In_1094,In_2523);
and U111 (N_111,In_885,In_1887);
nand U112 (N_112,In_1645,In_718);
and U113 (N_113,In_531,In_1283);
nor U114 (N_114,In_701,In_1838);
nand U115 (N_115,In_1727,In_1593);
nand U116 (N_116,In_462,In_2647);
or U117 (N_117,In_51,In_1231);
nor U118 (N_118,In_69,In_2829);
xor U119 (N_119,In_267,In_1115);
or U120 (N_120,In_230,In_1546);
nand U121 (N_121,In_613,In_1358);
or U122 (N_122,In_2866,In_93);
and U123 (N_123,In_384,In_775);
nand U124 (N_124,In_2400,In_1882);
and U125 (N_125,In_1794,In_2794);
xor U126 (N_126,In_893,In_2898);
and U127 (N_127,In_2563,In_735);
and U128 (N_128,In_1290,In_1880);
or U129 (N_129,In_1252,In_1092);
xnor U130 (N_130,In_1906,In_2080);
and U131 (N_131,In_322,In_256);
and U132 (N_132,In_1699,In_1336);
xor U133 (N_133,In_455,In_2351);
nand U134 (N_134,In_1964,In_1966);
or U135 (N_135,In_2649,In_1035);
xor U136 (N_136,In_2444,In_1083);
nor U137 (N_137,In_1419,In_1303);
nand U138 (N_138,In_2610,In_2923);
or U139 (N_139,In_1560,In_2803);
and U140 (N_140,In_2644,In_882);
nor U141 (N_141,In_2136,In_377);
or U142 (N_142,In_1428,In_2480);
xor U143 (N_143,In_215,In_1662);
and U144 (N_144,In_2785,In_2375);
nor U145 (N_145,In_1104,In_2936);
nand U146 (N_146,In_28,In_1767);
or U147 (N_147,In_1260,In_58);
xnor U148 (N_148,In_1904,In_1993);
or U149 (N_149,In_621,In_301);
xor U150 (N_150,In_2910,In_2038);
or U151 (N_151,In_1108,In_2763);
and U152 (N_152,In_2540,In_2742);
nor U153 (N_153,In_2843,In_1140);
or U154 (N_154,In_779,In_91);
nor U155 (N_155,In_686,In_874);
xor U156 (N_156,In_1011,In_484);
nand U157 (N_157,In_2949,In_2671);
nand U158 (N_158,In_796,In_422);
or U159 (N_159,In_2893,In_105);
nand U160 (N_160,In_2220,In_726);
nand U161 (N_161,In_2913,In_864);
or U162 (N_162,In_1587,In_1137);
xnor U163 (N_163,In_862,In_1725);
xnor U164 (N_164,In_1385,In_1068);
xnor U165 (N_165,In_442,In_937);
nor U166 (N_166,In_114,In_2903);
nor U167 (N_167,In_144,In_2907);
and U168 (N_168,In_2010,In_2464);
xnor U169 (N_169,In_653,In_46);
and U170 (N_170,In_835,In_86);
nand U171 (N_171,In_2420,In_1400);
and U172 (N_172,In_742,In_2980);
and U173 (N_173,In_2686,In_2297);
or U174 (N_174,In_2668,In_145);
nor U175 (N_175,In_1451,In_1368);
xor U176 (N_176,In_2930,In_660);
and U177 (N_177,In_642,In_2967);
or U178 (N_178,In_1681,In_532);
or U179 (N_179,In_695,In_608);
and U180 (N_180,In_566,In_509);
and U181 (N_181,In_529,In_1039);
or U182 (N_182,In_2461,In_2601);
and U183 (N_183,In_2445,In_396);
nand U184 (N_184,In_2484,In_180);
nor U185 (N_185,In_555,In_348);
nand U186 (N_186,In_2493,In_217);
or U187 (N_187,In_800,In_1192);
nor U188 (N_188,In_418,In_149);
or U189 (N_189,In_740,In_1223);
nand U190 (N_190,In_2448,In_1958);
or U191 (N_191,In_663,In_146);
and U192 (N_192,In_497,In_1536);
xor U193 (N_193,In_1122,In_1205);
nor U194 (N_194,In_2598,In_1036);
nand U195 (N_195,In_1810,In_1258);
or U196 (N_196,In_303,In_220);
nand U197 (N_197,In_1099,In_2955);
nor U198 (N_198,In_344,In_1222);
nor U199 (N_199,In_2043,In_2648);
nand U200 (N_200,In_730,In_2239);
nand U201 (N_201,In_2830,In_88);
and U202 (N_202,In_1544,In_211);
and U203 (N_203,In_234,In_2887);
and U204 (N_204,In_2109,In_2417);
or U205 (N_205,In_1112,In_1071);
and U206 (N_206,In_206,In_583);
and U207 (N_207,In_2185,In_2154);
or U208 (N_208,In_47,In_869);
and U209 (N_209,In_2699,In_2314);
nor U210 (N_210,In_363,In_1867);
and U211 (N_211,In_1708,In_731);
or U212 (N_212,In_1736,In_9);
nor U213 (N_213,In_414,In_1331);
nor U214 (N_214,In_1696,In_2243);
nor U215 (N_215,In_420,In_788);
and U216 (N_216,In_1491,In_1367);
xor U217 (N_217,In_661,In_1800);
xnor U218 (N_218,In_2875,In_1746);
and U219 (N_219,In_100,In_2547);
and U220 (N_220,In_327,In_1745);
nor U221 (N_221,In_2883,In_1895);
and U222 (N_222,In_2739,In_2708);
or U223 (N_223,In_2519,In_850);
nand U224 (N_224,In_877,In_1193);
or U225 (N_225,In_2677,In_383);
xnor U226 (N_226,In_1049,In_428);
or U227 (N_227,In_638,In_1394);
xor U228 (N_228,In_506,In_1490);
xor U229 (N_229,In_2954,In_1898);
nor U230 (N_230,In_1467,In_678);
nor U231 (N_231,In_429,In_280);
or U232 (N_232,In_1685,In_575);
nor U233 (N_233,In_1729,In_2987);
and U234 (N_234,In_243,In_2029);
xnor U235 (N_235,In_127,In_559);
xor U236 (N_236,In_2149,In_2326);
xor U237 (N_237,In_2072,In_2856);
xnor U238 (N_238,In_2757,In_410);
nor U239 (N_239,In_2238,In_360);
or U240 (N_240,In_703,In_2186);
or U241 (N_241,In_242,In_944);
nor U242 (N_242,In_514,In_1349);
nor U243 (N_243,In_2130,In_2611);
nor U244 (N_244,In_1514,In_150);
or U245 (N_245,In_102,In_987);
nand U246 (N_246,In_840,In_942);
nor U247 (N_247,In_2892,In_192);
nor U248 (N_248,In_2365,In_1983);
and U249 (N_249,In_495,In_1107);
or U250 (N_250,In_887,In_2700);
xor U251 (N_251,In_2941,In_48);
nor U252 (N_252,In_235,In_2008);
xor U253 (N_253,In_1586,In_1214);
or U254 (N_254,In_2421,In_1971);
or U255 (N_255,In_1273,In_2427);
nand U256 (N_256,In_2531,In_2582);
xor U257 (N_257,In_334,In_1959);
xor U258 (N_258,In_737,In_1138);
xor U259 (N_259,In_1089,In_1168);
and U260 (N_260,In_2174,In_1836);
or U261 (N_261,In_2858,In_2643);
and U262 (N_262,In_2355,In_352);
nor U263 (N_263,In_2983,In_2938);
nand U264 (N_264,In_1145,In_2016);
nor U265 (N_265,In_765,In_1850);
nand U266 (N_266,In_205,In_1420);
xnor U267 (N_267,In_983,In_2985);
or U268 (N_268,In_2681,In_1808);
xor U269 (N_269,In_671,In_2851);
or U270 (N_270,In_441,In_2234);
or U271 (N_271,In_369,In_1934);
nor U272 (N_272,In_2124,In_2635);
and U273 (N_273,In_1100,In_2925);
or U274 (N_274,In_2158,In_2438);
xor U275 (N_275,In_902,In_1754);
xor U276 (N_276,In_757,In_1302);
and U277 (N_277,In_2340,In_1652);
xor U278 (N_278,In_2990,In_141);
nand U279 (N_279,In_2979,In_2163);
nor U280 (N_280,In_865,In_2702);
nor U281 (N_281,In_2896,In_466);
nand U282 (N_282,In_2622,In_1238);
or U283 (N_283,In_2804,In_1789);
xor U284 (N_284,In_1481,In_1988);
and U285 (N_285,In_2069,In_1146);
or U286 (N_286,In_1430,In_1424);
xor U287 (N_287,In_1732,In_2439);
or U288 (N_288,In_1432,In_1739);
and U289 (N_289,In_1267,In_1143);
and U290 (N_290,In_1204,In_2614);
and U291 (N_291,In_1411,In_2864);
xnor U292 (N_292,In_2606,In_2951);
nor U293 (N_293,In_1907,In_2252);
xnor U294 (N_294,In_2828,In_14);
or U295 (N_295,In_1989,In_2545);
or U296 (N_296,In_503,In_491);
or U297 (N_297,In_2689,In_135);
nand U298 (N_298,In_2712,In_919);
and U299 (N_299,In_1213,In_1365);
or U300 (N_300,In_1409,In_2294);
or U301 (N_301,In_2352,In_593);
or U302 (N_302,In_505,In_2660);
xnor U303 (N_303,In_920,In_1706);
or U304 (N_304,In_1173,In_981);
and U305 (N_305,In_533,In_2569);
and U306 (N_306,In_1963,In_1236);
nand U307 (N_307,In_674,In_2137);
nand U308 (N_308,In_2203,In_710);
and U309 (N_309,In_2007,In_2659);
xor U310 (N_310,In_2092,In_1785);
or U311 (N_311,In_19,In_1396);
and U312 (N_312,In_2873,In_1172);
and U313 (N_313,In_2103,In_1435);
nand U314 (N_314,In_264,In_115);
and U315 (N_315,In_39,In_2613);
nand U316 (N_316,In_619,In_1629);
and U317 (N_317,In_2045,In_2769);
or U318 (N_318,In_724,In_1021);
or U319 (N_319,In_2612,In_2180);
or U320 (N_320,In_2259,In_475);
nand U321 (N_321,In_635,In_2429);
and U322 (N_322,In_2135,In_153);
or U323 (N_323,In_2773,In_1671);
nand U324 (N_324,In_1459,In_355);
nor U325 (N_325,In_2996,In_2662);
or U326 (N_326,In_1245,In_24);
xnor U327 (N_327,In_1817,In_1315);
nor U328 (N_328,In_1051,In_910);
nand U329 (N_329,In_967,In_411);
and U330 (N_330,In_1816,In_313);
or U331 (N_331,In_1753,In_649);
and U332 (N_332,In_1020,In_449);
nand U333 (N_333,In_2150,In_1740);
and U334 (N_334,In_1591,In_764);
nand U335 (N_335,In_493,In_907);
nor U336 (N_336,In_108,In_2319);
or U337 (N_337,In_2736,In_1686);
or U338 (N_338,In_2096,In_728);
and U339 (N_339,In_861,In_2315);
xor U340 (N_340,In_1741,In_117);
or U341 (N_341,In_2026,In_2539);
and U342 (N_342,In_1960,In_32);
nor U343 (N_343,In_1592,In_2057);
xnor U344 (N_344,In_232,In_592);
xnor U345 (N_345,In_1632,In_1869);
nor U346 (N_346,In_2552,In_451);
or U347 (N_347,In_1325,In_2431);
nand U348 (N_348,In_2615,In_20);
xor U349 (N_349,In_2003,In_2813);
nand U350 (N_350,In_561,In_2206);
nand U351 (N_351,In_2100,In_2338);
or U352 (N_352,In_1598,In_888);
and U353 (N_353,In_490,In_1650);
xor U354 (N_354,In_1731,In_616);
or U355 (N_355,In_567,In_1599);
and U356 (N_356,In_336,In_2968);
xnor U357 (N_357,In_1057,In_685);
nor U358 (N_358,In_1378,In_590);
nand U359 (N_359,In_1532,In_2703);
xor U360 (N_360,In_2188,In_1977);
nand U361 (N_361,In_74,In_1347);
nor U362 (N_362,In_1477,In_1045);
xor U363 (N_363,In_1634,In_2815);
and U364 (N_364,In_2264,In_270);
or U365 (N_365,In_2360,In_2318);
xor U366 (N_366,In_1928,In_655);
nor U367 (N_367,In_274,In_582);
xnor U368 (N_368,In_2811,In_1862);
and U369 (N_369,In_1773,In_604);
nor U370 (N_370,In_288,In_2176);
and U371 (N_371,In_1723,In_2111);
or U372 (N_372,In_792,In_2775);
nand U373 (N_373,In_1195,In_333);
xnor U374 (N_374,In_2462,In_2086);
nor U375 (N_375,In_1256,In_675);
nand U376 (N_376,In_2947,In_1298);
or U377 (N_377,In_1982,In_928);
nor U378 (N_378,In_2618,In_2854);
nor U379 (N_379,In_2256,In_972);
and U380 (N_380,In_1058,In_299);
and U381 (N_381,In_1431,In_851);
and U382 (N_382,In_78,In_1822);
nand U383 (N_383,In_1324,In_1229);
and U384 (N_384,In_1643,In_745);
nor U385 (N_385,In_1093,In_1233);
nor U386 (N_386,In_2428,In_2293);
nand U387 (N_387,In_1062,In_2877);
or U388 (N_388,In_1770,In_287);
nand U389 (N_389,In_2630,In_137);
xnor U390 (N_390,In_1539,In_408);
nor U391 (N_391,In_2113,In_969);
xor U392 (N_392,In_2802,In_798);
and U393 (N_393,In_809,In_282);
nor U394 (N_394,In_1893,In_985);
nor U395 (N_395,In_2138,In_759);
or U396 (N_396,In_1783,In_1961);
or U397 (N_397,In_717,In_2190);
or U398 (N_398,In_2976,In_1182);
and U399 (N_399,In_978,In_623);
nand U400 (N_400,In_502,In_2376);
or U401 (N_401,In_1744,In_2056);
or U402 (N_402,In_1755,In_2934);
nand U403 (N_403,In_719,In_1263);
nor U404 (N_404,In_478,In_2784);
nor U405 (N_405,In_838,In_2228);
nand U406 (N_406,In_1178,In_2741);
nand U407 (N_407,In_1621,In_1271);
and U408 (N_408,In_2665,In_1354);
xor U409 (N_409,In_2718,In_1391);
nor U410 (N_410,In_2272,In_1041);
and U411 (N_411,In_2780,In_793);
nor U412 (N_412,In_1209,In_1016);
or U413 (N_413,In_1933,In_2468);
xor U414 (N_414,In_2806,In_1828);
or U415 (N_415,In_2616,In_2194);
or U416 (N_416,In_2807,In_1525);
and U417 (N_417,In_498,In_2403);
nand U418 (N_418,In_1295,In_2078);
and U419 (N_419,In_1337,In_927);
nor U420 (N_420,In_188,In_2814);
xor U421 (N_421,In_448,In_992);
xnor U422 (N_422,In_2798,In_1653);
nor U423 (N_423,In_744,In_2178);
or U424 (N_424,In_1501,In_2962);
or U425 (N_425,In_246,In_2267);
xor U426 (N_426,In_2161,In_128);
or U427 (N_427,In_1320,In_2359);
xnor U428 (N_428,In_1284,In_1919);
nor U429 (N_429,In_2467,In_189);
nand U430 (N_430,In_1445,In_460);
and U431 (N_431,In_1473,In_366);
nor U432 (N_432,In_1373,In_1758);
nor U433 (N_433,In_2193,In_2364);
or U434 (N_434,In_1121,In_781);
nor U435 (N_435,In_553,In_1230);
nand U436 (N_436,In_2832,In_2216);
or U437 (N_437,In_1352,In_1562);
nor U438 (N_438,In_1136,In_0);
or U439 (N_439,In_799,In_1821);
nand U440 (N_440,In_525,In_648);
or U441 (N_441,In_2507,In_736);
nand U442 (N_442,In_2327,In_868);
or U443 (N_443,In_2578,In_1500);
xnor U444 (N_444,In_855,In_542);
xnor U445 (N_445,In_1050,In_644);
and U446 (N_446,In_1441,In_2179);
nand U447 (N_447,In_289,In_26);
nor U448 (N_448,In_1676,In_543);
and U449 (N_449,In_1694,In_1691);
nand U450 (N_450,In_1311,In_2652);
xnor U451 (N_451,In_2594,In_2991);
xnor U452 (N_452,In_2986,In_2393);
nor U453 (N_453,In_1151,In_1580);
xnor U454 (N_454,In_2240,In_1215);
nand U455 (N_455,In_689,In_546);
or U456 (N_456,In_1227,In_1452);
xnor U457 (N_457,In_1641,In_165);
or U458 (N_458,In_1235,In_2627);
nor U459 (N_459,In_1610,In_1877);
xor U460 (N_460,In_2479,In_1379);
nor U461 (N_461,In_2470,In_557);
or U462 (N_462,In_2564,In_2334);
nor U463 (N_463,In_1243,In_241);
and U464 (N_464,In_903,In_2891);
nor U465 (N_465,In_1200,In_315);
or U466 (N_466,In_486,In_2323);
and U467 (N_467,In_1572,In_1957);
nand U468 (N_468,In_403,In_1493);
nand U469 (N_469,In_1757,In_340);
nand U470 (N_470,In_2166,In_254);
or U471 (N_471,In_998,In_1206);
or U472 (N_472,In_763,In_413);
and U473 (N_473,In_2705,In_1091);
or U474 (N_474,In_1287,In_2093);
nand U475 (N_475,In_904,In_2006);
xnor U476 (N_476,In_496,In_1778);
nor U477 (N_477,In_1326,In_1123);
xnor U478 (N_478,In_2148,In_66);
and U479 (N_479,In_843,In_605);
or U480 (N_480,In_458,In_1637);
nor U481 (N_481,In_1523,In_1942);
or U482 (N_482,In_464,In_2325);
or U483 (N_483,In_1752,In_2122);
xor U484 (N_484,In_1793,In_1830);
nor U485 (N_485,In_1475,In_2882);
xnor U486 (N_486,In_2090,In_2235);
nor U487 (N_487,In_1889,In_2104);
nand U488 (N_488,In_2308,In_2404);
nor U489 (N_489,In_539,In_1922);
nand U490 (N_490,In_1037,In_361);
and U491 (N_491,In_1876,In_2544);
nor U492 (N_492,In_2607,In_1086);
and U493 (N_493,In_1462,In_345);
or U494 (N_494,In_634,In_2262);
xor U495 (N_495,In_1318,In_1030);
nor U496 (N_496,In_94,In_2812);
nor U497 (N_497,In_1716,In_1661);
nand U498 (N_498,In_367,In_61);
nand U499 (N_499,In_2079,In_109);
xor U500 (N_500,In_618,In_2287);
or U501 (N_501,In_1926,In_362);
nor U502 (N_502,In_173,In_1348);
nor U503 (N_503,In_526,In_304);
xor U504 (N_504,In_2593,In_2483);
and U505 (N_505,In_147,In_2760);
and U506 (N_506,In_210,In_2412);
xnor U507 (N_507,In_1310,In_783);
and U508 (N_508,In_2312,In_637);
or U509 (N_509,In_2232,In_1952);
xor U510 (N_510,In_412,In_1654);
nor U511 (N_511,In_1690,In_716);
nor U512 (N_512,In_1454,In_2442);
nor U513 (N_513,In_432,In_2978);
or U514 (N_514,In_2926,In_1468);
and U515 (N_515,In_1078,In_2992);
and U516 (N_516,In_222,In_953);
and U517 (N_517,In_1006,In_1261);
and U518 (N_518,In_2380,In_435);
nor U519 (N_519,In_1194,In_2906);
and U520 (N_520,In_2123,In_576);
nor U521 (N_521,In_1777,In_171);
nand U522 (N_522,In_857,In_706);
or U523 (N_523,In_1849,In_2245);
and U524 (N_524,In_1932,In_1679);
and U525 (N_525,In_2497,In_2860);
xnor U526 (N_526,In_2309,In_2588);
xnor U527 (N_527,In_1034,In_2076);
xor U528 (N_528,In_565,In_2840);
or U529 (N_529,In_2694,In_77);
or U530 (N_530,In_500,In_2603);
xor U531 (N_531,In_2848,In_1625);
or U532 (N_532,In_1812,In_63);
nor U533 (N_533,In_1798,In_1801);
nor U534 (N_534,In_1327,In_1133);
or U535 (N_535,In_1712,In_416);
nor U536 (N_536,In_2642,In_2328);
nor U537 (N_537,In_2746,In_297);
nand U538 (N_538,In_1359,In_2153);
or U539 (N_539,In_1834,In_227);
and U540 (N_540,In_867,In_1856);
xor U541 (N_541,In_2226,In_1535);
or U542 (N_542,In_2919,In_2880);
xnor U543 (N_543,In_2655,In_2912);
nor U544 (N_544,In_461,In_906);
and U545 (N_545,In_680,In_330);
xnor U546 (N_546,In_1790,In_1496);
nand U547 (N_547,In_2795,In_1197);
or U548 (N_548,In_767,In_1417);
xor U549 (N_549,In_156,In_2337);
or U550 (N_550,In_1902,In_2241);
or U551 (N_551,In_1682,In_2033);
nand U552 (N_552,In_1874,In_2725);
and U553 (N_553,In_2558,In_2397);
or U554 (N_554,In_2894,In_2963);
or U555 (N_555,In_1878,In_971);
or U556 (N_556,In_1968,In_2805);
and U557 (N_557,In_2676,In_2942);
nand U558 (N_558,In_1153,In_1534);
nand U559 (N_559,In_2939,In_1255);
nand U560 (N_560,In_1858,In_25);
xnor U561 (N_561,In_1802,In_2902);
xnor U562 (N_562,In_385,In_2684);
nand U563 (N_563,In_1619,In_2819);
nand U564 (N_564,In_2265,In_2273);
nand U565 (N_565,In_2062,In_488);
or U566 (N_566,In_2168,In_2787);
or U567 (N_567,In_2307,In_1628);
nand U568 (N_568,In_1782,In_1060);
nor U569 (N_569,In_1524,In_721);
xnor U570 (N_570,In_1601,In_2227);
xor U571 (N_571,In_600,In_1264);
and U572 (N_572,In_2639,In_2151);
nor U573 (N_573,In_1250,In_456);
and U574 (N_574,In_2706,In_1442);
or U575 (N_575,In_124,In_2960);
and U576 (N_576,In_2274,In_1381);
xor U577 (N_577,In_909,In_1322);
nand U578 (N_578,In_1416,In_1081);
nand U579 (N_579,In_913,In_260);
xor U580 (N_580,In_1915,In_41);
nor U581 (N_581,In_1936,In_2040);
nand U582 (N_582,In_1617,In_776);
nor U583 (N_583,In_1244,In_151);
or U584 (N_584,In_184,In_1516);
nor U585 (N_585,In_2482,In_10);
and U586 (N_586,In_2590,In_2341);
nor U587 (N_587,In_218,In_389);
and U588 (N_588,In_163,In_424);
and U589 (N_589,In_2504,In_522);
and U590 (N_590,In_2331,In_353);
and U591 (N_591,In_443,In_356);
nor U592 (N_592,In_1835,In_2455);
and U593 (N_593,In_84,In_2897);
or U594 (N_594,In_335,In_209);
xnor U595 (N_595,In_1829,In_2764);
nor U596 (N_596,In_167,In_292);
or U597 (N_597,In_1281,In_2211);
and U598 (N_598,In_107,In_2458);
or U599 (N_599,In_2197,In_1141);
xnor U600 (N_600,In_1019,In_2362);
or U601 (N_601,In_2378,In_1884);
or U602 (N_602,In_85,In_1090);
nor U603 (N_603,In_951,In_1566);
nand U604 (N_604,In_386,In_34);
xor U605 (N_605,In_2528,In_2105);
xnor U606 (N_606,In_2599,In_1096);
or U607 (N_607,In_2765,In_2127);
and U608 (N_608,In_1980,In_2946);
and U609 (N_609,In_2051,In_1987);
nand U610 (N_610,In_2070,In_2849);
nand U611 (N_611,In_1996,In_229);
or U612 (N_612,In_1228,In_948);
nand U613 (N_613,In_2841,In_2900);
nor U614 (N_614,In_1738,In_276);
or U615 (N_615,In_624,In_1371);
nand U616 (N_616,In_1823,In_2562);
nor U617 (N_617,In_1461,In_106);
xnor U618 (N_618,In_755,In_1160);
or U619 (N_619,In_2838,In_295);
xnor U620 (N_620,In_1914,In_1841);
or U621 (N_621,In_1015,In_512);
and U622 (N_622,In_482,In_1008);
or U623 (N_623,In_2390,In_1861);
xnor U624 (N_624,In_504,In_1762);
nand U625 (N_625,In_591,In_2899);
and U626 (N_626,In_2082,In_900);
and U627 (N_627,In_191,In_2723);
xor U628 (N_628,In_1527,In_2847);
or U629 (N_629,In_445,In_914);
xor U630 (N_630,In_71,In_236);
or U631 (N_631,In_2125,In_56);
nand U632 (N_632,In_1786,In_118);
xor U633 (N_633,In_2310,In_1248);
nand U634 (N_634,In_1814,In_131);
and U635 (N_635,In_2247,In_1872);
nor U636 (N_636,In_1607,In_249);
nor U637 (N_637,In_2128,In_1029);
nor U638 (N_638,In_2224,In_296);
and U639 (N_639,In_1582,In_357);
nor U640 (N_640,In_1943,In_1007);
and U641 (N_641,In_2567,In_970);
nor U642 (N_642,In_1791,In_1479);
nor U643 (N_643,In_2716,In_2320);
nor U644 (N_644,In_286,In_1279);
nand U645 (N_645,In_1189,In_1526);
or U646 (N_646,In_2835,In_2580);
or U647 (N_647,In_2524,In_732);
nor U648 (N_648,In_774,In_2961);
and U649 (N_649,In_2097,In_1220);
and U650 (N_650,In_545,In_1620);
xor U651 (N_651,In_1446,In_1262);
and U652 (N_652,In_2692,In_2498);
nand U653 (N_653,In_290,In_711);
nand U654 (N_654,In_2579,In_1647);
and U655 (N_655,In_2386,In_1102);
or U656 (N_656,In_1956,In_1766);
nor U657 (N_657,In_402,In_977);
or U658 (N_658,In_269,In_833);
nand U659 (N_659,In_2886,In_457);
nand U660 (N_660,In_2654,In_1323);
xnor U661 (N_661,In_1831,In_2997);
nor U662 (N_662,In_508,In_2525);
xor U663 (N_663,In_1280,In_687);
or U664 (N_664,In_2817,In_2004);
and U665 (N_665,In_1335,In_425);
nor U666 (N_666,In_1329,In_2286);
nor U667 (N_667,In_1130,In_2437);
or U668 (N_668,In_388,In_2000);
xnor U669 (N_669,In_1612,In_2871);
or U670 (N_670,In_2408,In_1372);
nand U671 (N_671,In_2222,In_1003);
or U672 (N_672,In_771,In_1508);
and U673 (N_673,In_2210,In_963);
or U674 (N_674,In_178,In_2698);
or U675 (N_675,In_347,In_794);
and U676 (N_676,In_1207,In_11);
nor U677 (N_677,In_1688,In_804);
or U678 (N_678,In_1509,In_2107);
or U679 (N_679,In_44,In_2719);
and U680 (N_680,In_921,In_1579);
and U681 (N_681,In_1890,In_652);
nor U682 (N_682,In_2585,In_1935);
nand U683 (N_683,In_262,In_733);
and U684 (N_684,In_578,In_2129);
nand U685 (N_685,In_1714,In_326);
xor U686 (N_686,In_2219,In_552);
xnor U687 (N_687,In_257,In_68);
or U688 (N_688,In_2300,In_677);
nor U689 (N_689,In_1054,In_2363);
xnor U690 (N_690,In_2704,In_2881);
xor U691 (N_691,In_1751,In_1923);
or U692 (N_692,In_1950,In_1404);
or U693 (N_693,In_841,In_1651);
nand U694 (N_694,In_2533,In_1402);
nor U695 (N_695,In_2641,In_828);
nor U696 (N_696,In_594,In_2369);
nor U697 (N_697,In_2110,In_2753);
and U698 (N_698,In_679,In_501);
nor U699 (N_699,In_1885,In_36);
nand U700 (N_700,In_2751,In_2876);
and U701 (N_701,In_1558,In_79);
nor U702 (N_702,In_2626,In_2249);
xnor U703 (N_703,In_2370,In_1014);
or U704 (N_704,In_683,In_2454);
or U705 (N_705,In_1826,In_92);
nand U706 (N_706,In_1999,In_2042);
nor U707 (N_707,In_1410,In_2500);
xnor U708 (N_708,In_650,In_2475);
nor U709 (N_709,In_1552,In_1275);
xnor U710 (N_710,In_2914,In_1085);
nor U711 (N_711,In_2869,In_617);
or U712 (N_712,In_1517,In_761);
nor U713 (N_713,In_2085,In_1557);
nand U714 (N_714,In_1109,In_430);
or U715 (N_715,In_2322,In_1570);
nand U716 (N_716,In_325,In_2460);
and U717 (N_717,In_2994,In_1597);
nand U718 (N_718,In_657,In_507);
nor U719 (N_719,In_960,In_487);
nand U720 (N_720,In_1633,In_1678);
nand U721 (N_721,In_1234,In_174);
nand U722 (N_722,In_2709,In_2152);
nor U723 (N_723,In_834,In_1139);
nand U724 (N_724,In_1606,In_251);
or U725 (N_725,In_2535,In_2002);
or U726 (N_726,In_1482,In_938);
or U727 (N_727,In_426,In_1009);
and U728 (N_728,In_481,In_1640);
and U729 (N_729,In_1405,In_1111);
and U730 (N_730,In_2710,In_2964);
nand U731 (N_731,In_2796,In_2382);
xor U732 (N_732,In_2248,In_691);
nand U733 (N_733,In_1809,In_1167);
and U734 (N_734,In_2836,In_2674);
or U735 (N_735,In_162,In_2502);
nor U736 (N_736,In_59,In_101);
or U737 (N_737,In_1772,In_317);
nor U738 (N_738,In_2083,In_1595);
nor U739 (N_739,In_2697,In_2212);
nand U740 (N_740,In_2101,In_1306);
or U741 (N_741,In_2646,In_1700);
and U742 (N_742,In_2496,In_2383);
nor U743 (N_743,In_2527,In_1897);
or U744 (N_744,In_2223,In_704);
and U745 (N_745,In_2321,In_2291);
or U746 (N_746,In_2532,In_155);
and U747 (N_747,In_2471,In_2884);
xnor U748 (N_748,In_2336,In_768);
or U749 (N_749,In_2581,In_284);
or U750 (N_750,In_1380,In_50);
nand U751 (N_751,In_1224,In_1297);
and U752 (N_752,In_2409,In_312);
nor U753 (N_753,In_626,In_1471);
nor U754 (N_754,In_2044,In_1157);
or U755 (N_755,In_2169,In_1346);
or U756 (N_756,In_419,In_2301);
nor U757 (N_757,In_2604,In_2682);
nor U758 (N_758,In_1813,In_1976);
nand U759 (N_759,In_2727,In_1434);
or U760 (N_760,In_609,In_2752);
nor U761 (N_761,In_55,In_2561);
nand U762 (N_762,In_1602,In_1480);
xor U763 (N_763,In_629,In_2139);
or U764 (N_764,In_1401,In_1374);
or U765 (N_765,In_2447,In_1330);
nand U766 (N_766,In_1292,In_1951);
or U767 (N_767,In_1695,In_433);
nor U768 (N_768,In_1565,In_2778);
nor U769 (N_769,In_602,In_376);
or U770 (N_770,In_1542,In_1196);
nand U771 (N_771,In_351,In_836);
nand U772 (N_772,In_1860,In_2766);
nor U773 (N_773,In_415,In_1246);
or U774 (N_774,In_82,In_2574);
nor U775 (N_775,In_2284,In_186);
nand U776 (N_776,In_889,In_2696);
and U777 (N_777,In_1425,In_392);
nor U778 (N_778,In_477,In_2918);
xor U779 (N_779,In_1340,In_517);
nor U780 (N_780,In_1668,In_873);
nand U781 (N_781,In_2218,In_1541);
and U782 (N_782,In_612,In_2634);
or U783 (N_783,In_556,In_941);
nor U784 (N_784,In_847,In_2357);
nor U785 (N_785,In_607,In_614);
and U786 (N_786,In_2459,In_1285);
and U787 (N_787,In_16,In_2413);
or U788 (N_788,In_1815,In_1639);
xnor U789 (N_789,In_2650,In_1663);
and U790 (N_790,In_2637,In_1073);
and U791 (N_791,In_285,In_2141);
nand U792 (N_792,In_120,In_729);
xor U793 (N_793,In_2053,In_2944);
nor U794 (N_794,In_2411,In_1150);
xor U795 (N_795,In_2575,In_2797);
or U796 (N_796,In_2071,In_2132);
or U797 (N_797,In_346,In_320);
nor U798 (N_798,In_2126,In_1403);
nand U799 (N_799,In_2826,In_434);
xor U800 (N_800,In_791,In_37);
nor U801 (N_801,In_2680,In_1028);
nor U802 (N_802,In_911,In_1724);
and U803 (N_803,In_140,In_2276);
or U804 (N_804,In_1916,In_1589);
xor U805 (N_805,In_1760,In_568);
xor U806 (N_806,In_2172,In_8);
nand U807 (N_807,In_1780,In_1135);
nand U808 (N_808,In_1515,In_2181);
xor U809 (N_809,In_2657,In_563);
nor U810 (N_810,In_852,In_1677);
nand U811 (N_811,In_2347,In_1203);
or U812 (N_812,In_2631,In_1013);
xnor U813 (N_813,In_2001,In_1362);
nor U814 (N_814,In_2280,In_2266);
nor U815 (N_815,In_483,In_339);
xnor U816 (N_816,In_1875,In_80);
and U817 (N_817,In_723,In_982);
and U818 (N_818,In_2722,In_746);
xor U819 (N_819,In_1180,In_394);
and U820 (N_820,In_2632,In_2950);
or U821 (N_821,In_103,In_1646);
nand U822 (N_822,In_1126,In_2118);
xor U823 (N_823,In_2799,In_2067);
or U824 (N_824,In_1657,In_1087);
or U825 (N_825,In_1486,In_1719);
xor U826 (N_826,In_2508,In_1567);
xnor U827 (N_827,In_1494,In_1364);
xor U828 (N_828,In_692,In_166);
nor U829 (N_829,In_2589,In_562);
or U830 (N_830,In_255,In_1818);
nand U831 (N_831,In_168,In_1673);
nor U832 (N_832,In_1803,In_1775);
or U833 (N_833,In_2529,In_1779);
and U834 (N_834,In_558,In_190);
nand U835 (N_835,In_1128,In_22);
or U836 (N_836,In_722,In_1232);
or U837 (N_837,In_2669,In_122);
nand U838 (N_838,In_1082,In_72);
nor U839 (N_839,In_2663,In_1370);
nand U840 (N_840,In_404,In_2516);
or U841 (N_841,In_1590,In_259);
nor U842 (N_842,In_727,In_935);
or U843 (N_843,In_250,In_2565);
or U844 (N_844,In_1384,In_708);
nor U845 (N_845,In_2270,In_2446);
nand U846 (N_846,In_705,In_1978);
nor U847 (N_847,In_494,In_813);
or U848 (N_848,In_1276,In_2425);
nor U849 (N_849,In_474,In_1221);
and U850 (N_850,In_1529,In_1931);
nand U851 (N_851,In_2667,In_959);
xor U852 (N_852,In_1018,In_407);
xnor U853 (N_853,In_2788,In_1339);
nand U854 (N_854,In_2728,In_715);
xnor U855 (N_855,In_669,In_2885);
or U856 (N_856,In_2469,In_2536);
and U857 (N_857,In_2664,In_939);
nand U858 (N_858,In_1506,In_2844);
nand U859 (N_859,In_2491,In_2350);
and U860 (N_860,In_1343,In_2505);
xor U861 (N_861,In_1533,In_1547);
and U862 (N_862,In_2731,In_1377);
nand U863 (N_863,In_2932,In_554);
nor U864 (N_864,In_15,In_891);
nor U865 (N_865,In_159,In_1995);
and U866 (N_866,In_753,In_2621);
xor U867 (N_867,In_1518,In_319);
or U868 (N_868,In_1611,In_628);
or U869 (N_869,In_228,In_1270);
xor U870 (N_870,In_309,In_283);
nand U871 (N_871,In_1511,In_2518);
nand U872 (N_872,In_1156,In_1569);
and U873 (N_873,In_170,In_898);
and U874 (N_874,In_516,In_2335);
xnor U875 (N_875,In_1764,In_820);
or U876 (N_876,In_1001,In_2927);
and U877 (N_877,In_1106,In_2450);
nor U878 (N_878,In_1537,In_2714);
nor U879 (N_879,In_164,In_350);
xor U880 (N_880,In_1155,In_2645);
and U881 (N_881,In_2073,In_2106);
or U882 (N_882,In_630,In_1472);
or U883 (N_883,In_397,In_599);
xnor U884 (N_884,In_830,In_842);
xnor U885 (N_885,In_64,In_1840);
nand U886 (N_886,In_1412,In_2416);
and U887 (N_887,In_2054,In_1747);
nand U888 (N_888,In_1164,In_955);
nand U889 (N_889,In_2957,In_2679);
or U890 (N_890,In_2673,In_2855);
and U891 (N_891,In_2385,In_2292);
or U892 (N_892,In_1990,In_752);
nand U893 (N_893,In_1351,In_2087);
nand U894 (N_894,In_1792,In_2288);
and U895 (N_895,In_143,In_2405);
xnor U896 (N_896,In_537,In_2027);
or U897 (N_897,In_450,In_52);
nand U898 (N_898,In_968,In_2099);
nor U899 (N_899,In_1077,In_787);
nor U900 (N_900,In_2021,In_2658);
or U901 (N_901,In_2173,In_2759);
nand U902 (N_902,In_2512,In_2121);
nand U903 (N_903,In_1588,In_365);
xor U904 (N_904,In_2879,In_1910);
or U905 (N_905,In_1148,In_1249);
or U906 (N_906,In_1820,In_1726);
nor U907 (N_907,In_879,In_1460);
nand U908 (N_908,In_221,In_965);
nor U909 (N_909,In_940,In_1784);
and U910 (N_910,In_950,In_1929);
or U911 (N_911,In_1312,In_712);
xnor U912 (N_912,In_1299,In_1658);
nor U913 (N_913,In_1962,In_2354);
nor U914 (N_914,In_645,In_447);
xor U915 (N_915,In_1811,In_743);
and U916 (N_916,In_1512,In_97);
nand U917 (N_917,In_2608,In_1711);
nor U918 (N_918,In_1355,In_1721);
xor U919 (N_919,In_754,In_2733);
or U920 (N_920,In_2171,In_2792);
and U921 (N_921,In_2250,In_1247);
xnor U922 (N_922,In_1718,In_2229);
xnor U923 (N_923,In_440,In_2015);
or U924 (N_924,In_1556,In_916);
and U925 (N_925,In_1072,In_639);
xor U926 (N_926,In_570,In_2779);
nand U927 (N_927,In_878,In_2768);
nand U928 (N_928,In_337,In_2155);
nor U929 (N_929,In_1618,In_1998);
nor U930 (N_930,In_1345,In_2440);
nand U931 (N_931,In_391,In_1879);
nor U932 (N_932,In_1076,In_1470);
or U933 (N_933,In_670,In_747);
nand U934 (N_934,In_2602,In_1769);
nor U935 (N_935,In_2762,In_2570);
and U936 (N_936,In_1549,In_2269);
and U937 (N_937,In_1891,In_121);
nand U938 (N_938,In_2456,In_2344);
nand U939 (N_939,In_1210,In_2772);
nand U940 (N_940,In_431,In_364);
nor U941 (N_941,In_21,In_1948);
and U942 (N_942,In_2800,In_1555);
and U943 (N_943,In_244,In_2970);
nor U944 (N_944,In_1069,In_1465);
nor U945 (N_945,In_2971,In_1159);
and U946 (N_946,In_1457,In_1847);
nor U947 (N_947,In_2553,In_1894);
and U948 (N_948,In_1868,In_2761);
nor U949 (N_949,In_651,In_1584);
nor U950 (N_950,In_2931,In_1017);
nand U951 (N_951,In_2487,In_2857);
nor U952 (N_952,In_2809,In_2261);
and U953 (N_953,In_1510,In_2853);
or U954 (N_954,In_870,In_368);
and U955 (N_955,In_1608,In_1848);
or U956 (N_956,In_2419,In_2018);
or U957 (N_957,In_2332,In_1047);
and U958 (N_958,In_2145,In_1774);
nand U959 (N_959,In_2046,In_1328);
and U960 (N_960,In_2670,In_2583);
xnor U961 (N_961,In_2494,In_2823);
nand U962 (N_962,In_2691,In_817);
or U963 (N_963,In_1649,In_1116);
xnor U964 (N_964,In_548,In_2387);
and U965 (N_965,In_2551,In_371);
nor U966 (N_966,In_2422,In_1543);
and U967 (N_967,In_936,In_29);
and U968 (N_968,In_208,In_1053);
or U969 (N_969,In_1846,In_2984);
nand U970 (N_970,In_216,In_436);
and U971 (N_971,In_2271,In_193);
nand U972 (N_972,In_2406,In_897);
and U973 (N_973,In_2867,In_2989);
and U974 (N_974,In_831,In_2204);
nand U975 (N_975,In_2777,In_976);
or U976 (N_976,In_2011,In_2052);
nor U977 (N_977,In_1505,In_2771);
and U978 (N_978,In_1440,In_2490);
and U979 (N_979,In_606,In_2724);
nand U980 (N_980,In_1208,In_2559);
xor U981 (N_981,In_1382,In_1414);
nand U982 (N_982,In_316,In_2770);
or U983 (N_983,In_2789,In_476);
or U984 (N_984,In_1559,In_2133);
xnor U985 (N_985,In_95,In_749);
nand U986 (N_986,In_993,In_579);
and U987 (N_987,In_2878,In_2666);
and U988 (N_988,In_1985,In_995);
or U989 (N_989,In_1061,In_2783);
nand U990 (N_990,In_1930,In_1918);
xnor U991 (N_991,In_2625,In_784);
or U992 (N_992,In_1048,In_2595);
and U993 (N_993,In_17,In_633);
and U994 (N_994,In_42,In_67);
nand U995 (N_995,In_564,In_2966);
nand U996 (N_996,In_2605,In_1819);
nand U997 (N_997,In_328,In_2242);
nand U998 (N_998,In_1864,In_709);
xnor U999 (N_999,In_176,In_1202);
or U1000 (N_1000,In_2568,In_2556);
xnor U1001 (N_1001,In_2453,In_308);
xor U1002 (N_1002,In_528,In_112);
or U1003 (N_1003,In_595,In_1576);
nor U1004 (N_1004,In_588,In_521);
xor U1005 (N_1005,In_123,In_2872);
and U1006 (N_1006,In_2820,In_2825);
nor U1007 (N_1007,In_2501,In_1870);
or U1008 (N_1008,In_803,In_379);
nor U1009 (N_1009,In_273,In_60);
xnor U1010 (N_1010,In_1981,In_2032);
nor U1011 (N_1011,In_1722,In_2973);
or U1012 (N_1012,In_1975,In_2810);
and U1013 (N_1013,In_2683,In_1333);
and U1014 (N_1014,In_550,In_966);
xnor U1015 (N_1015,In_991,In_1398);
or U1016 (N_1016,In_2142,In_1680);
and U1017 (N_1017,In_2131,In_2217);
or U1018 (N_1018,In_1911,In_2596);
nor U1019 (N_1019,In_187,In_1307);
and U1020 (N_1020,In_785,In_584);
nor U1021 (N_1021,In_789,In_947);
nand U1022 (N_1022,In_1038,In_2672);
nor U1023 (N_1023,In_2993,In_1067);
or U1024 (N_1024,In_293,In_2514);
nor U1025 (N_1025,In_2277,In_802);
or U1026 (N_1026,In_821,In_1174);
or U1027 (N_1027,In_2948,In_2177);
nor U1028 (N_1028,In_375,In_819);
or U1029 (N_1029,In_2426,In_918);
xor U1030 (N_1030,In_175,In_2068);
xor U1031 (N_1031,In_2868,In_266);
nor U1032 (N_1032,In_1585,In_2619);
xnor U1033 (N_1033,In_2358,In_622);
and U1034 (N_1034,In_398,In_1023);
nor U1035 (N_1035,In_510,In_2846);
xor U1036 (N_1036,In_1488,In_2255);
and U1037 (N_1037,In_1578,In_459);
xnor U1038 (N_1038,In_1925,In_702);
xor U1039 (N_1039,In_1871,In_2781);
nand U1040 (N_1040,In_806,In_2084);
nor U1041 (N_1041,In_393,In_1970);
nor U1042 (N_1042,In_323,In_1920);
nor U1043 (N_1043,In_1886,In_822);
and U1044 (N_1044,In_1953,In_826);
nand U1045 (N_1045,In_1225,In_2546);
or U1046 (N_1046,In_2024,In_75);
and U1047 (N_1047,In_1055,In_54);
and U1048 (N_1048,In_1423,In_1630);
xor U1049 (N_1049,In_2384,In_1080);
xnor U1050 (N_1050,In_1286,In_2050);
nor U1051 (N_1051,In_2506,In_1319);
nor U1052 (N_1052,In_627,In_2162);
or U1053 (N_1053,In_894,In_2114);
xnor U1054 (N_1054,In_1733,In_2975);
nor U1055 (N_1055,In_2793,In_2244);
xnor U1056 (N_1056,In_2430,In_1692);
and U1057 (N_1057,In_2859,In_1940);
xor U1058 (N_1058,In_2031,In_70);
nor U1059 (N_1059,In_646,In_2808);
nor U1060 (N_1060,In_1002,In_240);
or U1061 (N_1061,In_2213,In_523);
xnor U1062 (N_1062,In_1032,In_2253);
nor U1063 (N_1063,In_139,In_1421);
nand U1064 (N_1064,In_667,In_2489);
nor U1065 (N_1065,In_2304,In_1360);
nand U1066 (N_1066,In_1687,In_2921);
and U1067 (N_1067,In_2999,In_520);
and U1068 (N_1068,In_1253,In_45);
nand U1069 (N_1069,In_1756,In_2943);
xor U1070 (N_1070,In_932,In_2275);
xnor U1071 (N_1071,In_2695,In_1946);
or U1072 (N_1072,In_2982,In_2088);
xnor U1073 (N_1073,In_1763,In_1426);
or U1074 (N_1074,In_1768,In_816);
nor U1075 (N_1075,In_1463,In_1707);
nor U1076 (N_1076,In_547,In_2609);
or U1077 (N_1077,In_1308,In_2466);
and U1078 (N_1078,In_1622,In_2348);
xor U1079 (N_1079,In_489,In_1237);
nand U1080 (N_1080,In_2049,In_1866);
or U1081 (N_1081,In_1575,In_1742);
nor U1082 (N_1082,In_1881,In_1670);
nor U1083 (N_1083,In_2734,In_2116);
nor U1084 (N_1084,In_1044,In_713);
and U1085 (N_1085,In_2395,In_2555);
or U1086 (N_1086,In_1938,In_2576);
nand U1087 (N_1087,In_952,In_860);
nand U1088 (N_1088,In_2758,In_1383);
nand U1089 (N_1089,In_2418,In_700);
or U1090 (N_1090,In_611,In_849);
nor U1091 (N_1091,In_2191,In_926);
nand U1092 (N_1092,In_2345,In_467);
or U1093 (N_1093,In_2047,In_2510);
nor U1094 (N_1094,In_2965,In_1269);
or U1095 (N_1095,In_1485,In_1010);
or U1096 (N_1096,In_12,In_751);
nand U1097 (N_1097,In_2165,In_2195);
nor U1098 (N_1098,In_923,In_65);
xnor U1099 (N_1099,In_1603,In_231);
and U1100 (N_1100,In_2041,In_2282);
xor U1101 (N_1101,In_1737,In_1144);
nand U1102 (N_1102,In_1912,In_2862);
or U1103 (N_1103,In_1259,In_805);
or U1104 (N_1104,In_2463,In_2225);
xor U1105 (N_1105,In_949,In_615);
or U1106 (N_1106,In_725,In_272);
or U1107 (N_1107,In_1761,In_152);
and U1108 (N_1108,In_104,In_659);
nand U1109 (N_1109,In_1005,In_1448);
xor U1110 (N_1110,In_1059,In_2207);
nor U1111 (N_1111,In_1507,In_2701);
or U1112 (N_1112,In_1124,In_1568);
nor U1113 (N_1113,In_3,In_35);
nor U1114 (N_1114,In_219,In_825);
and U1115 (N_1115,In_1788,In_2693);
nor U1116 (N_1116,In_1185,In_43);
nand U1117 (N_1117,In_1832,In_1163);
and U1118 (N_1118,In_2023,In_2617);
and U1119 (N_1119,In_1033,In_581);
or U1120 (N_1120,In_1363,In_1851);
xnor U1121 (N_1121,In_38,In_1909);
nand U1122 (N_1122,In_1070,In_2638);
nand U1123 (N_1123,In_1825,In_2164);
or U1124 (N_1124,In_1357,In_2077);
and U1125 (N_1125,In_2061,In_1636);
or U1126 (N_1126,In_2656,In_1052);
nor U1127 (N_1127,In_1594,In_2058);
and U1128 (N_1128,In_908,In_2394);
nand U1129 (N_1129,In_2030,In_96);
xor U1130 (N_1130,In_571,In_1497);
xnor U1131 (N_1131,In_2221,In_2929);
nor U1132 (N_1132,In_2449,In_1046);
or U1133 (N_1133,In_1954,In_884);
or U1134 (N_1134,In_2102,In_138);
and U1135 (N_1135,In_1973,In_126);
xor U1136 (N_1136,In_694,In_1079);
nor U1137 (N_1137,In_2296,In_773);
or U1138 (N_1138,In_1118,In_1344);
nor U1139 (N_1139,In_2112,In_2298);
or U1140 (N_1140,In_2120,In_872);
xor U1141 (N_1141,In_1896,In_1908);
and U1142 (N_1142,In_1458,In_359);
nor U1143 (N_1143,In_247,In_1499);
nor U1144 (N_1144,In_676,In_2316);
xnor U1145 (N_1145,In_1000,In_18);
or U1146 (N_1146,In_2822,In_2196);
nand U1147 (N_1147,In_760,In_1476);
and U1148 (N_1148,In_696,In_324);
nor U1149 (N_1149,In_2730,In_2952);
xor U1150 (N_1150,In_261,In_1334);
nand U1151 (N_1151,In_2009,In_381);
nor U1152 (N_1152,In_896,In_252);
and U1153 (N_1153,In_720,In_1191);
nor U1154 (N_1154,In_2231,In_2557);
nor U1155 (N_1155,In_631,In_778);
nor U1156 (N_1156,In_2717,In_134);
and U1157 (N_1157,In_2721,In_890);
or U1158 (N_1158,In_1321,In_1624);
and U1159 (N_1159,In_2969,In_1845);
or U1160 (N_1160,In_1314,In_2423);
xor U1161 (N_1161,In_2089,In_2095);
nand U1162 (N_1162,In_540,In_1844);
and U1163 (N_1163,In_1605,In_782);
nand U1164 (N_1164,In_2330,In_2014);
nand U1165 (N_1165,In_2690,In_2767);
and U1166 (N_1166,In_1583,In_1697);
nor U1167 (N_1167,In_2687,In_541);
nand U1168 (N_1168,In_1702,In_684);
nor U1169 (N_1169,In_1903,In_2850);
or U1170 (N_1170,In_4,In_1278);
nor U1171 (N_1171,In_177,In_185);
and U1172 (N_1172,In_2842,In_1450);
or U1173 (N_1173,In_2339,In_1);
xnor U1174 (N_1174,In_1614,In_1759);
nand U1175 (N_1175,In_2201,In_1361);
xnor U1176 (N_1176,In_2192,In_2094);
nor U1177 (N_1177,In_2283,In_83);
nor U1178 (N_1178,In_1395,In_933);
and U1179 (N_1179,In_2624,In_1149);
or U1180 (N_1180,In_681,In_2432);
xor U1181 (N_1181,In_2530,In_780);
or U1182 (N_1182,In_2974,In_2678);
nor U1183 (N_1183,In_2711,In_306);
and U1184 (N_1184,In_2313,In_846);
or U1185 (N_1185,In_2937,In_1216);
or U1186 (N_1186,In_2549,In_2713);
and U1187 (N_1187,In_1113,In_7);
nor U1188 (N_1188,In_2119,In_382);
nand U1189 (N_1189,In_2586,In_854);
nand U1190 (N_1190,In_1674,In_1186);
nand U1191 (N_1191,In_133,In_1613);
nand U1192 (N_1192,In_1353,In_572);
nor U1193 (N_1193,In_688,In_49);
xor U1194 (N_1194,In_2349,In_1098);
nand U1195 (N_1195,In_1842,In_1177);
nand U1196 (N_1196,In_2012,In_957);
or U1197 (N_1197,In_207,In_1941);
nand U1198 (N_1198,In_2573,In_279);
xor U1199 (N_1199,In_1495,In_1272);
nand U1200 (N_1200,In_2538,In_454);
or U1201 (N_1201,In_2543,In_291);
xnor U1202 (N_1202,In_198,In_1433);
and U1203 (N_1203,In_823,In_1088);
nor U1204 (N_1204,In_2305,In_1012);
nor U1205 (N_1205,In_1806,In_573);
nor U1206 (N_1206,In_2055,In_1439);
and U1207 (N_1207,In_1805,In_238);
or U1208 (N_1208,In_766,In_2268);
or U1209 (N_1209,In_829,In_807);
and U1210 (N_1210,In_179,In_2520);
xor U1211 (N_1211,In_472,In_654);
or U1212 (N_1212,In_2592,In_160);
xor U1213 (N_1213,In_2289,In_2584);
xor U1214 (N_1214,In_405,In_824);
and U1215 (N_1215,In_1522,In_2035);
and U1216 (N_1216,In_1254,In_2134);
nand U1217 (N_1217,In_1701,In_1623);
xnor U1218 (N_1218,In_427,In_421);
nand U1219 (N_1219,In_2436,In_1066);
and U1220 (N_1220,In_585,In_2774);
or U1221 (N_1221,In_2776,In_1937);
nor U1222 (N_1222,In_1004,In_2175);
or U1223 (N_1223,In_2653,In_2279);
or U1224 (N_1224,In_480,In_158);
and U1225 (N_1225,In_2156,In_2303);
nand U1226 (N_1226,In_2063,In_1025);
nor U1227 (N_1227,In_212,In_739);
nor U1228 (N_1228,In_1103,In_2550);
and U1229 (N_1229,In_790,In_2410);
xnor U1230 (N_1230,In_99,In_2324);
xor U1231 (N_1231,In_406,In_2933);
nor U1232 (N_1232,In_81,In_1239);
and U1233 (N_1233,In_587,In_1561);
or U1234 (N_1234,In_2499,In_853);
nand U1235 (N_1235,In_848,In_1114);
xor U1236 (N_1236,In_2548,In_2465);
or U1237 (N_1237,In_1161,In_580);
nand U1238 (N_1238,In_2917,In_1504);
and U1239 (N_1239,In_2317,In_453);
xnor U1240 (N_1240,In_401,In_2916);
or U1241 (N_1241,In_1715,In_2202);
or U1242 (N_1242,In_1852,In_2170);
xnor U1243 (N_1243,In_110,In_1944);
nor U1244 (N_1244,In_13,In_839);
nor U1245 (N_1245,In_2143,In_2361);
and U1246 (N_1246,In_1147,In_1119);
and U1247 (N_1247,In_1171,In_577);
xor U1248 (N_1248,In_2367,In_307);
or U1249 (N_1249,In_2620,In_183);
xnor U1250 (N_1250,In_302,In_268);
nand U1251 (N_1251,In_1313,In_1571);
xor U1252 (N_1252,In_1924,In_756);
nand U1253 (N_1253,In_714,In_943);
nor U1254 (N_1254,In_811,In_2542);
nor U1255 (N_1255,In_125,In_329);
and U1256 (N_1256,In_1456,In_1949);
nor U1257 (N_1257,In_181,In_1181);
and U1258 (N_1258,In_2435,In_2372);
and U1259 (N_1259,In_2839,In_446);
nand U1260 (N_1260,In_321,In_1064);
xnor U1261 (N_1261,In_2889,In_975);
nor U1262 (N_1262,In_1289,In_672);
or U1263 (N_1263,In_2922,In_827);
xnor U1264 (N_1264,In_2258,In_875);
or U1265 (N_1265,In_1487,In_1095);
or U1266 (N_1266,In_2600,In_1703);
and U1267 (N_1267,In_1771,In_1854);
or U1268 (N_1268,In_2628,In_2473);
or U1269 (N_1269,In_1705,In_1429);
nor U1270 (N_1270,In_2415,In_2977);
nand U1271 (N_1271,In_1305,In_2343);
xnor U1272 (N_1272,In_275,In_1776);
or U1273 (N_1273,In_2115,In_439);
and U1274 (N_1274,In_2290,In_845);
or U1275 (N_1275,In_2414,In_1901);
xnor U1276 (N_1276,In_378,In_485);
nor U1277 (N_1277,In_2831,In_2039);
xnor U1278 (N_1278,In_1388,In_1166);
nand U1279 (N_1279,In_682,In_2998);
nor U1280 (N_1280,In_2146,In_332);
and U1281 (N_1281,In_2254,In_946);
nor U1282 (N_1282,In_586,In_2791);
xor U1283 (N_1283,In_2726,In_87);
xnor U1284 (N_1284,In_2740,In_1043);
and U1285 (N_1285,In_1667,In_560);
xnor U1286 (N_1286,In_1453,In_2495);
xnor U1287 (N_1287,In_1997,In_1188);
or U1288 (N_1288,In_915,In_2521);
and U1289 (N_1289,In_1131,In_2451);
nor U1290 (N_1290,In_2481,In_2890);
and U1291 (N_1291,In_2865,In_2988);
xor U1292 (N_1292,In_372,In_1097);
nand U1293 (N_1293,In_417,In_294);
or U1294 (N_1294,In_1201,In_1795);
xor U1295 (N_1295,In_2801,In_1169);
nand U1296 (N_1296,In_2863,In_2208);
xor U1297 (N_1297,In_1530,In_399);
xnor U1298 (N_1298,In_1888,In_772);
and U1299 (N_1299,In_934,In_354);
and U1300 (N_1300,In_1626,In_2485);
nand U1301 (N_1301,In_2074,In_738);
nand U1302 (N_1302,In_1063,In_1979);
xor U1303 (N_1303,In_300,In_1554);
or U1304 (N_1304,In_2554,In_374);
nand U1305 (N_1305,In_2636,In_2909);
nor U1306 (N_1306,In_197,In_1443);
nor U1307 (N_1307,In_27,In_2541);
xor U1308 (N_1308,In_1437,In_1427);
xnor U1309 (N_1309,In_2342,In_2147);
nor U1310 (N_1310,In_182,In_2920);
nor U1311 (N_1311,In_2441,In_1799);
nor U1312 (N_1312,In_815,In_2492);
and U1313 (N_1313,In_148,In_2756);
nand U1314 (N_1314,In_2623,In_1341);
nand U1315 (N_1315,In_310,In_899);
nor U1316 (N_1316,In_1293,In_2388);
or U1317 (N_1317,In_1190,In_658);
nor U1318 (N_1318,In_233,In_1531);
nand U1319 (N_1319,In_1024,In_1655);
and U1320 (N_1320,In_2066,In_925);
and U1321 (N_1321,In_1992,In_1892);
nand U1322 (N_1322,In_748,In_2346);
and U1323 (N_1323,In_647,In_2022);
nand U1324 (N_1324,In_2472,In_395);
nor U1325 (N_1325,In_2729,In_786);
or U1326 (N_1326,In_2786,In_2901);
nand U1327 (N_1327,In_620,In_538);
nor U1328 (N_1328,In_194,In_707);
nand U1329 (N_1329,In_536,In_518);
nor U1330 (N_1330,In_1538,In_837);
xor U1331 (N_1331,In_1438,In_598);
xor U1332 (N_1332,In_438,In_1444);
nand U1333 (N_1333,In_1581,In_1748);
and U1334 (N_1334,In_2230,In_1548);
nand U1335 (N_1335,In_2754,In_2640);
xor U1336 (N_1336,In_214,In_984);
nand U1337 (N_1337,In_2407,In_2522);
nand U1338 (N_1338,In_1631,In_980);
and U1339 (N_1339,In_2743,In_1316);
or U1340 (N_1340,In_2953,In_98);
and U1341 (N_1341,In_1158,In_2389);
and U1342 (N_1342,In_2852,In_2560);
or U1343 (N_1343,In_1212,In_204);
nand U1344 (N_1344,In_2911,In_1553);
nand U1345 (N_1345,In_1502,In_452);
xor U1346 (N_1346,In_492,In_640);
or U1347 (N_1347,In_1294,In_2036);
nor U1348 (N_1348,In_1132,In_1859);
xnor U1349 (N_1349,In_601,In_2098);
xnor U1350 (N_1350,In_2503,In_1827);
nor U1351 (N_1351,In_278,In_1288);
xnor U1352 (N_1352,In_2478,In_1939);
nor U1353 (N_1353,In_265,In_2013);
nor U1354 (N_1354,In_1551,In_996);
xor U1355 (N_1355,In_2928,In_1332);
xor U1356 (N_1356,In_1955,In_1309);
or U1357 (N_1357,In_5,In_2260);
and U1358 (N_1358,In_53,In_1873);
and U1359 (N_1359,In_1026,In_1291);
nor U1360 (N_1360,In_801,In_2028);
nor U1361 (N_1361,In_1521,In_1648);
nor U1362 (N_1362,In_423,In_1397);
xnor U1363 (N_1363,In_1689,In_2081);
and U1364 (N_1364,In_1219,In_2895);
xnor U1365 (N_1365,In_1833,In_1474);
or U1366 (N_1366,In_1600,In_2295);
and U1367 (N_1367,In_527,In_2572);
or U1368 (N_1368,In_974,In_1743);
and U1369 (N_1369,In_223,In_172);
xnor U1370 (N_1370,In_2457,In_1693);
xor U1371 (N_1371,In_1198,In_161);
nor U1372 (N_1372,In_2905,In_90);
xor U1373 (N_1373,In_1899,In_2782);
and U1374 (N_1374,In_2299,In_1125);
nor U1375 (N_1375,In_116,In_1734);
nor U1376 (N_1376,In_1127,In_2117);
nand U1377 (N_1377,In_2157,In_2737);
or U1378 (N_1378,In_632,In_387);
and U1379 (N_1379,In_1117,In_471);
nand U1380 (N_1380,In_2486,In_2515);
or U1381 (N_1381,In_1609,In_1406);
xnor U1382 (N_1382,In_1179,In_1152);
nand U1383 (N_1383,In_1965,In_2748);
xnor U1384 (N_1384,In_1162,In_1199);
or U1385 (N_1385,In_1176,In_2371);
xor U1386 (N_1386,In_1282,In_1120);
nor U1387 (N_1387,In_1390,In_1183);
and U1388 (N_1388,In_1240,In_625);
or U1389 (N_1389,In_1615,In_922);
nand U1390 (N_1390,In_1666,In_662);
nor U1391 (N_1391,In_1843,In_1170);
nand U1392 (N_1392,In_2488,In_1642);
xnor U1393 (N_1393,In_1986,In_142);
and U1394 (N_1394,In_1266,In_2236);
or U1395 (N_1395,In_2396,In_876);
nand U1396 (N_1396,In_2200,In_770);
xor U1397 (N_1397,In_239,In_1389);
nand U1398 (N_1398,In_196,In_2443);
xnor U1399 (N_1399,In_2037,In_1110);
or U1400 (N_1400,In_666,In_2816);
xnor U1401 (N_1401,In_380,In_2167);
nor U1402 (N_1402,In_1824,In_2511);
or U1403 (N_1403,In_2707,In_1074);
or U1404 (N_1404,In_892,In_373);
and U1405 (N_1405,In_226,In_1717);
or U1406 (N_1406,In_866,In_2108);
xnor U1407 (N_1407,In_258,In_1710);
nand U1408 (N_1408,In_2591,In_859);
nand U1409 (N_1409,In_2391,In_812);
or U1410 (N_1410,In_1974,In_1350);
and U1411 (N_1411,In_73,In_569);
and U1412 (N_1412,In_1084,In_1855);
xnor U1413 (N_1413,In_2159,In_2381);
nor U1414 (N_1414,In_1296,In_597);
nor U1415 (N_1415,In_1698,In_341);
nor U1416 (N_1416,In_1366,In_2720);
nand U1417 (N_1417,In_1342,In_1921);
or U1418 (N_1418,In_2215,In_62);
xor U1419 (N_1419,In_2477,In_1184);
and U1420 (N_1420,In_2995,In_444);
nor U1421 (N_1421,In_808,In_2199);
xnor U1422 (N_1422,In_2065,In_2945);
nand U1423 (N_1423,In_1393,In_2981);
and U1424 (N_1424,In_698,In_1927);
or U1425 (N_1425,In_1134,In_2183);
and U1426 (N_1426,In_119,In_1900);
and U1427 (N_1427,In_999,In_931);
or U1428 (N_1428,In_479,In_858);
nand U1429 (N_1429,In_2189,In_1664);
xnor U1430 (N_1430,In_1675,In_1520);
or U1431 (N_1431,In_2246,In_1187);
nand U1432 (N_1432,In_2379,In_1241);
and U1433 (N_1433,In_1804,In_979);
or U1434 (N_1434,In_2629,In_912);
or U1435 (N_1435,In_905,In_2366);
and U1436 (N_1436,In_697,In_665);
xnor U1437 (N_1437,In_1863,In_1947);
nand U1438 (N_1438,In_2749,In_1883);
nand U1439 (N_1439,In_1797,In_643);
or U1440 (N_1440,In_224,In_1528);
and U1441 (N_1441,In_31,In_988);
nor U1442 (N_1442,In_271,In_929);
nand U1443 (N_1443,In_741,In_277);
nand U1444 (N_1444,In_2744,In_810);
or U1445 (N_1445,In_2747,In_2019);
or U1446 (N_1446,In_1129,In_535);
or U1447 (N_1447,In_2587,In_305);
nor U1448 (N_1448,In_2233,In_1503);
and U1449 (N_1449,In_1750,In_1466);
and U1450 (N_1450,In_132,In_1665);
nor U1451 (N_1451,In_945,In_1175);
or U1452 (N_1452,In_2959,In_154);
and U1453 (N_1453,In_901,In_129);
or U1454 (N_1454,In_1713,In_880);
and U1455 (N_1455,In_1056,In_2182);
xnor U1456 (N_1456,In_551,In_1386);
or U1457 (N_1457,In_2571,In_1422);
nand U1458 (N_1458,In_994,In_2688);
and U1459 (N_1459,In_202,In_814);
nand U1460 (N_1460,In_2837,In_2474);
or U1461 (N_1461,In_668,In_1573);
or U1462 (N_1462,In_1656,In_1635);
or U1463 (N_1463,In_1574,In_2517);
nand U1464 (N_1464,In_1787,In_954);
and U1465 (N_1465,In_1376,In_1596);
nor U1466 (N_1466,In_2924,In_2940);
nor U1467 (N_1467,In_1991,In_1563);
or U1468 (N_1468,In_1242,In_1040);
xnor U1469 (N_1469,In_1807,In_636);
and U1470 (N_1470,In_473,In_2091);
nor U1471 (N_1471,In_349,In_2356);
and U1472 (N_1472,In_1519,In_1545);
xor U1473 (N_1473,In_1913,In_298);
nand U1474 (N_1474,In_513,In_1101);
xnor U1475 (N_1475,In_225,In_863);
nor U1476 (N_1476,In_2399,In_1436);
or U1477 (N_1477,In_856,In_1338);
and U1478 (N_1478,In_1075,In_2187);
nor U1479 (N_1479,In_1317,In_574);
and U1480 (N_1480,In_1905,In_2184);
xor U1481 (N_1481,In_1226,In_2263);
xnor U1482 (N_1482,In_930,In_2972);
nand U1483 (N_1483,In_519,In_2402);
nor U1484 (N_1484,In_2537,In_201);
or U1485 (N_1485,In_515,In_1265);
nor U1486 (N_1486,In_2392,In_2566);
xnor U1487 (N_1487,In_2368,In_2214);
or U1488 (N_1488,In_33,In_734);
nand U1489 (N_1489,In_1765,In_1356);
nand U1490 (N_1490,In_1165,In_130);
or U1491 (N_1491,In_1300,In_2908);
xnor U1492 (N_1492,In_511,In_2874);
or U1493 (N_1493,In_23,In_469);
xor U1494 (N_1494,In_1513,In_1413);
xor U1495 (N_1495,In_2534,In_1304);
and U1496 (N_1496,In_1730,In_157);
nand U1497 (N_1497,In_499,In_1022);
nand U1498 (N_1498,In_2821,In_1728);
nor U1499 (N_1499,In_997,In_2633);
xnor U1500 (N_1500,N_499,N_800);
or U1501 (N_1501,N_518,N_1332);
and U1502 (N_1502,N_35,N_1444);
xnor U1503 (N_1503,N_1291,N_798);
or U1504 (N_1504,N_1247,N_866);
and U1505 (N_1505,N_911,N_318);
nor U1506 (N_1506,N_2,N_981);
and U1507 (N_1507,N_1145,N_925);
or U1508 (N_1508,N_1077,N_1290);
and U1509 (N_1509,N_838,N_643);
nand U1510 (N_1510,N_10,N_246);
or U1511 (N_1511,N_11,N_27);
and U1512 (N_1512,N_679,N_658);
or U1513 (N_1513,N_1347,N_1167);
or U1514 (N_1514,N_1335,N_718);
and U1515 (N_1515,N_855,N_285);
nand U1516 (N_1516,N_1386,N_900);
and U1517 (N_1517,N_358,N_948);
nor U1518 (N_1518,N_1397,N_527);
nand U1519 (N_1519,N_775,N_1231);
or U1520 (N_1520,N_29,N_753);
or U1521 (N_1521,N_1334,N_858);
and U1522 (N_1522,N_1030,N_168);
nor U1523 (N_1523,N_553,N_854);
nor U1524 (N_1524,N_1163,N_409);
xnor U1525 (N_1525,N_535,N_145);
nand U1526 (N_1526,N_1243,N_249);
and U1527 (N_1527,N_110,N_44);
xnor U1528 (N_1528,N_173,N_1306);
xor U1529 (N_1529,N_395,N_22);
nor U1530 (N_1530,N_1365,N_1311);
nand U1531 (N_1531,N_376,N_675);
nor U1532 (N_1532,N_75,N_1426);
nand U1533 (N_1533,N_219,N_845);
nand U1534 (N_1534,N_259,N_808);
xor U1535 (N_1535,N_266,N_1092);
xor U1536 (N_1536,N_708,N_677);
or U1537 (N_1537,N_993,N_1049);
nor U1538 (N_1538,N_412,N_136);
xnor U1539 (N_1539,N_1399,N_1435);
or U1540 (N_1540,N_242,N_1074);
and U1541 (N_1541,N_279,N_966);
nor U1542 (N_1542,N_108,N_768);
nor U1543 (N_1543,N_156,N_1417);
nor U1544 (N_1544,N_1010,N_1225);
xor U1545 (N_1545,N_760,N_441);
xor U1546 (N_1546,N_1430,N_443);
or U1547 (N_1547,N_1498,N_1428);
and U1548 (N_1548,N_404,N_1439);
xnor U1549 (N_1549,N_1375,N_55);
nand U1550 (N_1550,N_484,N_359);
or U1551 (N_1551,N_23,N_1127);
xnor U1552 (N_1552,N_1124,N_324);
and U1553 (N_1553,N_148,N_670);
and U1554 (N_1554,N_388,N_352);
or U1555 (N_1555,N_142,N_86);
and U1556 (N_1556,N_1041,N_232);
nand U1557 (N_1557,N_275,N_298);
nand U1558 (N_1558,N_868,N_998);
xor U1559 (N_1559,N_68,N_1034);
and U1560 (N_1560,N_899,N_574);
or U1561 (N_1561,N_398,N_140);
nor U1562 (N_1562,N_1004,N_1045);
nand U1563 (N_1563,N_117,N_1009);
xnor U1564 (N_1564,N_1304,N_365);
xnor U1565 (N_1565,N_1340,N_78);
xnor U1566 (N_1566,N_756,N_505);
nor U1567 (N_1567,N_69,N_573);
xnor U1568 (N_1568,N_1138,N_620);
nand U1569 (N_1569,N_24,N_551);
nor U1570 (N_1570,N_691,N_1204);
nand U1571 (N_1571,N_70,N_1227);
nor U1572 (N_1572,N_65,N_1436);
nand U1573 (N_1573,N_881,N_1473);
nor U1574 (N_1574,N_992,N_1275);
or U1575 (N_1575,N_1406,N_486);
nand U1576 (N_1576,N_373,N_150);
nor U1577 (N_1577,N_678,N_896);
or U1578 (N_1578,N_1285,N_1058);
or U1579 (N_1579,N_1210,N_880);
and U1580 (N_1580,N_585,N_1300);
xnor U1581 (N_1581,N_623,N_436);
xnor U1582 (N_1582,N_419,N_872);
nor U1583 (N_1583,N_652,N_805);
xnor U1584 (N_1584,N_81,N_516);
and U1585 (N_1585,N_433,N_466);
nand U1586 (N_1586,N_1410,N_294);
xor U1587 (N_1587,N_537,N_1273);
and U1588 (N_1588,N_781,N_1368);
nand U1589 (N_1589,N_875,N_1173);
xor U1590 (N_1590,N_685,N_405);
nor U1591 (N_1591,N_1431,N_179);
xnor U1592 (N_1592,N_1061,N_133);
or U1593 (N_1593,N_837,N_299);
xor U1594 (N_1594,N_920,N_1251);
nand U1595 (N_1595,N_1202,N_1080);
nand U1596 (N_1596,N_943,N_622);
nor U1597 (N_1597,N_84,N_542);
nor U1598 (N_1598,N_305,N_751);
nor U1599 (N_1599,N_661,N_515);
nand U1600 (N_1600,N_833,N_1160);
nor U1601 (N_1601,N_238,N_719);
xnor U1602 (N_1602,N_132,N_306);
or U1603 (N_1603,N_733,N_1188);
nor U1604 (N_1604,N_391,N_1494);
nor U1605 (N_1605,N_1423,N_169);
nand U1606 (N_1606,N_774,N_743);
and U1607 (N_1607,N_525,N_171);
nand U1608 (N_1608,N_471,N_1109);
nor U1609 (N_1609,N_859,N_269);
xnor U1610 (N_1610,N_1170,N_188);
and U1611 (N_1611,N_186,N_288);
nor U1612 (N_1612,N_368,N_762);
nand U1613 (N_1613,N_651,N_876);
or U1614 (N_1614,N_1242,N_139);
or U1615 (N_1615,N_1280,N_983);
and U1616 (N_1616,N_1168,N_1257);
nand U1617 (N_1617,N_834,N_625);
and U1618 (N_1618,N_940,N_1027);
or U1619 (N_1619,N_1469,N_45);
and U1620 (N_1620,N_461,N_742);
or U1621 (N_1621,N_1238,N_335);
nor U1622 (N_1622,N_990,N_913);
or U1623 (N_1623,N_767,N_163);
xor U1624 (N_1624,N_1000,N_1298);
or U1625 (N_1625,N_814,N_822);
xnor U1626 (N_1626,N_97,N_206);
nor U1627 (N_1627,N_331,N_271);
nand U1628 (N_1628,N_1040,N_410);
and U1629 (N_1629,N_105,N_343);
nor U1630 (N_1630,N_1294,N_144);
and U1631 (N_1631,N_252,N_1342);
xor U1632 (N_1632,N_502,N_349);
nor U1633 (N_1633,N_1106,N_146);
xor U1634 (N_1634,N_53,N_423);
xnor U1635 (N_1635,N_1310,N_923);
nor U1636 (N_1636,N_350,N_772);
xnor U1637 (N_1637,N_149,N_1020);
and U1638 (N_1638,N_348,N_465);
nand U1639 (N_1639,N_1371,N_1354);
nor U1640 (N_1640,N_453,N_495);
or U1641 (N_1641,N_185,N_548);
nand U1642 (N_1642,N_362,N_96);
and U1643 (N_1643,N_1464,N_209);
or U1644 (N_1644,N_653,N_101);
nand U1645 (N_1645,N_1333,N_501);
nor U1646 (N_1646,N_204,N_690);
and U1647 (N_1647,N_236,N_1266);
nand U1648 (N_1648,N_955,N_668);
xor U1649 (N_1649,N_706,N_892);
and U1650 (N_1650,N_245,N_1068);
nor U1651 (N_1651,N_1383,N_1296);
nand U1652 (N_1652,N_716,N_1262);
xor U1653 (N_1653,N_635,N_1403);
nand U1654 (N_1654,N_48,N_260);
and U1655 (N_1655,N_17,N_1116);
and U1656 (N_1656,N_1054,N_283);
and U1657 (N_1657,N_492,N_965);
nand U1658 (N_1658,N_648,N_1451);
and U1659 (N_1659,N_612,N_284);
nor U1660 (N_1660,N_1203,N_457);
or U1661 (N_1661,N_1098,N_1197);
or U1662 (N_1662,N_1139,N_823);
nand U1663 (N_1663,N_1321,N_222);
nand U1664 (N_1664,N_1302,N_939);
and U1665 (N_1665,N_1478,N_1424);
or U1666 (N_1666,N_182,N_1412);
nand U1667 (N_1667,N_1018,N_1015);
xnor U1668 (N_1668,N_1187,N_208);
and U1669 (N_1669,N_255,N_1355);
nand U1670 (N_1670,N_1212,N_750);
xor U1671 (N_1671,N_1105,N_248);
nand U1672 (N_1672,N_510,N_601);
nor U1673 (N_1673,N_201,N_887);
nor U1674 (N_1674,N_1317,N_570);
xor U1675 (N_1675,N_119,N_50);
nor U1676 (N_1676,N_780,N_309);
xor U1677 (N_1677,N_893,N_942);
xor U1678 (N_1678,N_166,N_212);
nand U1679 (N_1679,N_203,N_910);
or U1680 (N_1680,N_1026,N_104);
xnor U1681 (N_1681,N_795,N_1353);
xor U1682 (N_1682,N_287,N_1208);
nor U1683 (N_1683,N_159,N_1241);
nor U1684 (N_1684,N_46,N_421);
or U1685 (N_1685,N_124,N_563);
and U1686 (N_1686,N_824,N_1462);
nor U1687 (N_1687,N_735,N_1148);
nor U1688 (N_1688,N_1263,N_995);
xor U1689 (N_1689,N_438,N_281);
xor U1690 (N_1690,N_1179,N_107);
nor U1691 (N_1691,N_464,N_1044);
nand U1692 (N_1692,N_909,N_320);
and U1693 (N_1693,N_1463,N_1396);
nand U1694 (N_1694,N_1232,N_1282);
or U1695 (N_1695,N_1432,N_401);
xnor U1696 (N_1696,N_1459,N_1352);
nor U1697 (N_1697,N_844,N_1465);
xnor U1698 (N_1698,N_974,N_901);
nor U1699 (N_1699,N_1229,N_366);
nand U1700 (N_1700,N_771,N_637);
and U1701 (N_1701,N_740,N_544);
or U1702 (N_1702,N_1186,N_1073);
nand U1703 (N_1703,N_1065,N_250);
or U1704 (N_1704,N_1453,N_1388);
xor U1705 (N_1705,N_511,N_33);
nor U1706 (N_1706,N_435,N_1096);
xnor U1707 (N_1707,N_1324,N_536);
and U1708 (N_1708,N_996,N_717);
or U1709 (N_1709,N_1401,N_1377);
nor U1710 (N_1710,N_1035,N_1209);
xnor U1711 (N_1711,N_1316,N_314);
and U1712 (N_1712,N_916,N_1192);
nor U1713 (N_1713,N_646,N_216);
nor U1714 (N_1714,N_857,N_121);
nand U1715 (N_1715,N_540,N_313);
xor U1716 (N_1716,N_569,N_1404);
or U1717 (N_1717,N_789,N_235);
nand U1718 (N_1718,N_1499,N_430);
nor U1719 (N_1719,N_547,N_514);
or U1720 (N_1720,N_432,N_748);
xor U1721 (N_1721,N_697,N_175);
nand U1722 (N_1722,N_999,N_172);
or U1723 (N_1723,N_1166,N_956);
nand U1724 (N_1724,N_1177,N_886);
and U1725 (N_1725,N_1095,N_659);
nand U1726 (N_1726,N_333,N_810);
and U1727 (N_1727,N_1346,N_400);
or U1728 (N_1728,N_1066,N_1370);
nand U1729 (N_1729,N_420,N_958);
or U1730 (N_1730,N_602,N_877);
nand U1731 (N_1731,N_657,N_19);
nor U1732 (N_1732,N_427,N_224);
or U1733 (N_1733,N_962,N_337);
xor U1734 (N_1734,N_1440,N_915);
nand U1735 (N_1735,N_1114,N_125);
and U1736 (N_1736,N_462,N_1284);
xor U1737 (N_1737,N_1323,N_533);
nor U1738 (N_1738,N_82,N_89);
nor U1739 (N_1739,N_88,N_1129);
xnor U1740 (N_1740,N_725,N_1385);
or U1741 (N_1741,N_389,N_897);
or U1742 (N_1742,N_727,N_758);
xnor U1743 (N_1743,N_341,N_312);
nand U1744 (N_1744,N_1483,N_60);
nor U1745 (N_1745,N_381,N_1190);
nor U1746 (N_1746,N_1216,N_1201);
xor U1747 (N_1747,N_1407,N_322);
and U1748 (N_1748,N_933,N_21);
nor U1749 (N_1749,N_1090,N_1117);
and U1750 (N_1750,N_61,N_1207);
and U1751 (N_1751,N_989,N_353);
or U1752 (N_1752,N_666,N_566);
nand U1753 (N_1753,N_1137,N_523);
and U1754 (N_1754,N_634,N_663);
xor U1755 (N_1755,N_1445,N_1158);
nand U1756 (N_1756,N_165,N_1477);
or U1757 (N_1757,N_526,N_194);
or U1758 (N_1758,N_494,N_196);
xnor U1759 (N_1759,N_649,N_31);
xnor U1760 (N_1760,N_827,N_356);
nor U1761 (N_1761,N_426,N_512);
nand U1762 (N_1762,N_1394,N_1362);
or U1763 (N_1763,N_572,N_264);
and U1764 (N_1764,N_746,N_1467);
and U1765 (N_1765,N_832,N_1051);
xor U1766 (N_1766,N_1131,N_673);
nand U1767 (N_1767,N_982,N_1021);
nor U1768 (N_1768,N_195,N_906);
nor U1769 (N_1769,N_785,N_787);
nand U1770 (N_1770,N_1153,N_1199);
nor U1771 (N_1771,N_597,N_302);
and U1772 (N_1772,N_25,N_935);
nor U1773 (N_1773,N_1289,N_485);
and U1774 (N_1774,N_579,N_745);
and U1775 (N_1775,N_681,N_586);
and U1776 (N_1776,N_683,N_98);
nand U1777 (N_1777,N_478,N_672);
or U1778 (N_1778,N_617,N_1339);
or U1779 (N_1779,N_1482,N_967);
xnor U1780 (N_1780,N_1380,N_506);
and U1781 (N_1781,N_600,N_1017);
nor U1782 (N_1782,N_447,N_638);
or U1783 (N_1783,N_42,N_230);
nor U1784 (N_1784,N_338,N_330);
nor U1785 (N_1785,N_557,N_1097);
or U1786 (N_1786,N_1455,N_3);
or U1787 (N_1787,N_289,N_1071);
nor U1788 (N_1788,N_1246,N_1067);
nand U1789 (N_1789,N_1249,N_122);
or U1790 (N_1790,N_874,N_629);
nor U1791 (N_1791,N_761,N_828);
and U1792 (N_1792,N_567,N_975);
and U1793 (N_1793,N_472,N_654);
and U1794 (N_1794,N_841,N_550);
nor U1795 (N_1795,N_801,N_1359);
and U1796 (N_1796,N_197,N_1287);
nand U1797 (N_1797,N_254,N_5);
xor U1798 (N_1798,N_813,N_1055);
nand U1799 (N_1799,N_66,N_723);
nand U1800 (N_1800,N_481,N_1172);
nand U1801 (N_1801,N_1140,N_233);
xor U1802 (N_1802,N_1079,N_190);
xor U1803 (N_1803,N_1016,N_1230);
and U1804 (N_1804,N_1029,N_985);
nand U1805 (N_1805,N_739,N_351);
and U1806 (N_1806,N_327,N_1134);
and U1807 (N_1807,N_731,N_522);
and U1808 (N_1808,N_325,N_30);
and U1809 (N_1809,N_267,N_321);
or U1810 (N_1810,N_1292,N_41);
nand U1811 (N_1811,N_1420,N_1367);
and U1812 (N_1812,N_15,N_1413);
and U1813 (N_1813,N_1261,N_198);
and U1814 (N_1814,N_817,N_883);
and U1815 (N_1815,N_62,N_36);
and U1816 (N_1816,N_1155,N_80);
nand U1817 (N_1817,N_103,N_1226);
xnor U1818 (N_1818,N_997,N_1084);
nor U1819 (N_1819,N_12,N_978);
nand U1820 (N_1820,N_234,N_759);
xnor U1821 (N_1821,N_1272,N_766);
nand U1822 (N_1822,N_1120,N_1326);
xor U1823 (N_1823,N_34,N_843);
xnor U1824 (N_1824,N_729,N_580);
or U1825 (N_1825,N_891,N_393);
or U1826 (N_1826,N_1237,N_1064);
xor U1827 (N_1827,N_696,N_747);
xor U1828 (N_1828,N_741,N_434);
nand U1829 (N_1829,N_1094,N_1075);
or U1830 (N_1830,N_1411,N_240);
or U1831 (N_1831,N_1220,N_662);
nand U1832 (N_1832,N_694,N_702);
xor U1833 (N_1833,N_83,N_1288);
nor U1834 (N_1834,N_418,N_831);
xnor U1835 (N_1835,N_1456,N_802);
or U1836 (N_1836,N_528,N_6);
and U1837 (N_1837,N_972,N_630);
xor U1838 (N_1838,N_300,N_310);
and U1839 (N_1839,N_1119,N_1319);
or U1840 (N_1840,N_1037,N_217);
nor U1841 (N_1841,N_703,N_724);
or U1842 (N_1842,N_1108,N_116);
nor U1843 (N_1843,N_268,N_131);
nor U1844 (N_1844,N_1256,N_1384);
nand U1845 (N_1845,N_1043,N_1457);
and U1846 (N_1846,N_1422,N_459);
xor U1847 (N_1847,N_961,N_1366);
or U1848 (N_1848,N_929,N_986);
or U1849 (N_1849,N_755,N_460);
or U1850 (N_1850,N_1265,N_934);
or U1851 (N_1851,N_1062,N_686);
xnor U1852 (N_1852,N_227,N_777);
nor U1853 (N_1853,N_1038,N_1327);
xnor U1854 (N_1854,N_1048,N_1233);
and U1855 (N_1855,N_37,N_77);
or U1856 (N_1856,N_815,N_562);
nor U1857 (N_1857,N_847,N_1104);
xnor U1858 (N_1858,N_183,N_1374);
xnor U1859 (N_1859,N_92,N_1349);
or U1860 (N_1860,N_701,N_1057);
xor U1861 (N_1861,N_39,N_228);
nand U1862 (N_1862,N_912,N_498);
or U1863 (N_1863,N_991,N_257);
nor U1864 (N_1864,N_431,N_769);
and U1865 (N_1865,N_200,N_40);
or U1866 (N_1866,N_1001,N_1376);
nor U1867 (N_1867,N_180,N_1126);
nor U1868 (N_1868,N_469,N_1031);
xor U1869 (N_1869,N_1112,N_296);
xor U1870 (N_1870,N_976,N_1497);
nand U1871 (N_1871,N_1111,N_1466);
nor U1872 (N_1872,N_1214,N_446);
or U1873 (N_1873,N_821,N_754);
and U1874 (N_1874,N_816,N_738);
xor U1875 (N_1875,N_921,N_26);
and U1876 (N_1876,N_1184,N_736);
or U1877 (N_1877,N_850,N_317);
nand U1878 (N_1878,N_263,N_812);
nor U1879 (N_1879,N_440,N_1063);
or U1880 (N_1880,N_1185,N_396);
or U1881 (N_1881,N_803,N_1492);
xor U1882 (N_1882,N_851,N_390);
nand U1883 (N_1883,N_377,N_1046);
xnor U1884 (N_1884,N_1003,N_928);
xor U1885 (N_1885,N_541,N_261);
xnor U1886 (N_1886,N_450,N_804);
and U1887 (N_1887,N_411,N_951);
and U1888 (N_1888,N_123,N_596);
and U1889 (N_1889,N_959,N_636);
nand U1890 (N_1890,N_1305,N_20);
or U1891 (N_1891,N_592,N_370);
nor U1892 (N_1892,N_626,N_790);
xnor U1893 (N_1893,N_1414,N_732);
xnor U1894 (N_1894,N_1490,N_1224);
and U1895 (N_1895,N_907,N_138);
or U1896 (N_1896,N_950,N_59);
and U1897 (N_1897,N_1433,N_734);
xor U1898 (N_1898,N_1052,N_1418);
nor U1899 (N_1899,N_1434,N_1245);
nand U1900 (N_1900,N_1019,N_1244);
and U1901 (N_1901,N_1475,N_922);
and U1902 (N_1902,N_1053,N_546);
and U1903 (N_1903,N_1060,N_442);
nor U1904 (N_1904,N_1299,N_229);
nand U1905 (N_1905,N_1107,N_603);
nand U1906 (N_1906,N_1337,N_1171);
or U1907 (N_1907,N_917,N_1381);
nand U1908 (N_1908,N_737,N_154);
and U1909 (N_1909,N_595,N_1449);
and U1910 (N_1910,N_470,N_0);
and U1911 (N_1911,N_560,N_763);
and U1912 (N_1912,N_1211,N_334);
nand U1913 (N_1913,N_386,N_1147);
and U1914 (N_1914,N_1144,N_1491);
xor U1915 (N_1915,N_757,N_1024);
xnor U1916 (N_1916,N_957,N_193);
nor U1917 (N_1917,N_231,N_1283);
nand U1918 (N_1918,N_307,N_937);
and U1919 (N_1919,N_120,N_784);
xor U1920 (N_1920,N_403,N_1248);
xor U1921 (N_1921,N_521,N_1328);
and U1922 (N_1922,N_712,N_655);
nand U1923 (N_1923,N_825,N_277);
or U1924 (N_1924,N_94,N_1012);
xnor U1925 (N_1925,N_820,N_1461);
nor U1926 (N_1926,N_111,N_1222);
nand U1927 (N_1927,N_1379,N_239);
nand U1928 (N_1928,N_559,N_591);
nand U1929 (N_1929,N_1496,N_964);
or U1930 (N_1930,N_665,N_364);
xor U1931 (N_1931,N_707,N_660);
nor U1932 (N_1932,N_1269,N_1421);
nand U1933 (N_1933,N_994,N_303);
nand U1934 (N_1934,N_95,N_1110);
or U1935 (N_1935,N_914,N_1348);
nand U1936 (N_1936,N_863,N_1358);
xor U1937 (N_1937,N_902,N_7);
or U1938 (N_1938,N_503,N_531);
and U1939 (N_1939,N_474,N_829);
nand U1940 (N_1940,N_176,N_380);
or U1941 (N_1941,N_1442,N_1183);
and U1942 (N_1942,N_693,N_1143);
xor U1943 (N_1943,N_152,N_496);
xor U1944 (N_1944,N_720,N_276);
nand U1945 (N_1945,N_1329,N_424);
xnor U1946 (N_1946,N_157,N_954);
nand U1947 (N_1947,N_1429,N_555);
and U1948 (N_1948,N_1113,N_109);
or U1949 (N_1949,N_127,N_839);
nor U1950 (N_1950,N_1336,N_968);
nand U1951 (N_1951,N_1364,N_1303);
nand U1952 (N_1952,N_243,N_1318);
nand U1953 (N_1953,N_1078,N_1056);
nor U1954 (N_1954,N_270,N_1416);
nor U1955 (N_1955,N_413,N_286);
xnor U1956 (N_1956,N_1125,N_819);
or U1957 (N_1957,N_864,N_604);
or U1958 (N_1958,N_114,N_189);
xor U1959 (N_1959,N_1441,N_882);
nor U1960 (N_1960,N_1205,N_818);
or U1961 (N_1961,N_765,N_641);
and U1962 (N_1962,N_487,N_1286);
nand U1963 (N_1963,N_1471,N_1135);
nor U1964 (N_1964,N_205,N_616);
and U1965 (N_1965,N_141,N_143);
nand U1966 (N_1966,N_379,N_1474);
and U1967 (N_1967,N_609,N_1360);
nor U1968 (N_1968,N_1322,N_339);
nand U1969 (N_1969,N_1175,N_1142);
or U1970 (N_1970,N_64,N_297);
xnor U1971 (N_1971,N_1356,N_137);
or U1972 (N_1972,N_1258,N_1234);
and U1973 (N_1973,N_422,N_463);
nor U1974 (N_1974,N_644,N_710);
and U1975 (N_1975,N_1361,N_794);
nand U1976 (N_1976,N_316,N_392);
xor U1977 (N_1977,N_1351,N_265);
nor U1978 (N_1978,N_687,N_1382);
xor U1979 (N_1979,N_764,N_1191);
nand U1980 (N_1980,N_1314,N_1118);
xor U1981 (N_1981,N_1484,N_927);
or U1982 (N_1982,N_621,N_184);
and U1983 (N_1983,N_272,N_1452);
or U1984 (N_1984,N_1146,N_278);
or U1985 (N_1985,N_842,N_346);
xor U1986 (N_1986,N_375,N_508);
xor U1987 (N_1987,N_530,N_564);
or U1988 (N_1988,N_695,N_1278);
or U1989 (N_1989,N_782,N_354);
nor U1990 (N_1990,N_456,N_387);
nand U1991 (N_1991,N_632,N_1270);
or U1992 (N_1992,N_153,N_1387);
or U1993 (N_1993,N_262,N_607);
nor U1994 (N_1994,N_898,N_1254);
or U1995 (N_1995,N_517,N_473);
nor U1996 (N_1996,N_1193,N_155);
or U1997 (N_1997,N_76,N_1133);
xor U1998 (N_1998,N_164,N_865);
and U1999 (N_1999,N_210,N_1402);
nor U2000 (N_2000,N_878,N_1239);
or U2001 (N_2001,N_223,N_529);
xor U2002 (N_2002,N_214,N_1345);
and U2003 (N_2003,N_319,N_63);
xnor U2004 (N_2004,N_1460,N_1268);
nor U2005 (N_2005,N_308,N_490);
nor U2006 (N_2006,N_888,N_1400);
xnor U2007 (N_2007,N_479,N_1330);
xnor U2008 (N_2008,N_1132,N_1088);
and U2009 (N_2009,N_793,N_889);
xnor U2010 (N_2010,N_1182,N_328);
nand U2011 (N_2011,N_323,N_336);
nor U2012 (N_2012,N_476,N_192);
or U2013 (N_2013,N_449,N_1450);
nand U2014 (N_2014,N_606,N_840);
or U2015 (N_2015,N_581,N_879);
nor U2016 (N_2016,N_588,N_1217);
nand U2017 (N_2017,N_1223,N_99);
xnor U2018 (N_2018,N_1392,N_273);
nand U2019 (N_2019,N_1389,N_941);
and U2020 (N_2020,N_406,N_714);
nand U2021 (N_2021,N_115,N_1255);
nand U2022 (N_2022,N_482,N_360);
xnor U2023 (N_2023,N_1039,N_689);
or U2024 (N_2024,N_1005,N_280);
nand U2025 (N_2025,N_1130,N_1196);
and U2026 (N_2026,N_1028,N_700);
and U2027 (N_2027,N_856,N_1032);
nor U2028 (N_2028,N_181,N_645);
and U2029 (N_2029,N_692,N_1378);
and U2030 (N_2030,N_797,N_539);
nor U2031 (N_2031,N_584,N_984);
and U2032 (N_2032,N_870,N_575);
nor U2033 (N_2033,N_477,N_1150);
nand U2034 (N_2034,N_407,N_1331);
xor U2035 (N_2035,N_258,N_846);
or U2036 (N_2036,N_680,N_1219);
xnor U2037 (N_2037,N_971,N_274);
and U2038 (N_2038,N_1121,N_332);
or U2039 (N_2039,N_1458,N_969);
or U2040 (N_2040,N_633,N_47);
nor U2041 (N_2041,N_1315,N_93);
nand U2042 (N_2042,N_1264,N_129);
and U2043 (N_2043,N_4,N_345);
or U2044 (N_2044,N_699,N_1115);
xnor U2045 (N_2045,N_87,N_1279);
or U2046 (N_2046,N_56,N_904);
nor U2047 (N_2047,N_605,N_650);
or U2048 (N_2048,N_836,N_1487);
xor U2049 (N_2049,N_786,N_1011);
xnor U2050 (N_2050,N_382,N_952);
or U2051 (N_2051,N_647,N_135);
or U2052 (N_2052,N_51,N_1309);
nor U2053 (N_2053,N_1101,N_744);
and U2054 (N_2054,N_326,N_73);
nor U2055 (N_2055,N_556,N_752);
nand U2056 (N_2056,N_1023,N_458);
xnor U2057 (N_2057,N_329,N_1180);
nor U2058 (N_2058,N_253,N_770);
nand U2059 (N_2059,N_16,N_524);
nor U2060 (N_2060,N_1437,N_520);
nand U2061 (N_2061,N_247,N_429);
and U2062 (N_2062,N_594,N_1076);
xor U2063 (N_2063,N_1174,N_344);
nor U2064 (N_2064,N_1398,N_1082);
nand U2065 (N_2065,N_684,N_945);
nand U2066 (N_2066,N_355,N_849);
nor U2067 (N_2067,N_1086,N_295);
and U2068 (N_2068,N_18,N_613);
and U2069 (N_2069,N_451,N_9);
nor U2070 (N_2070,N_439,N_167);
nand U2071 (N_2071,N_397,N_749);
nor U2072 (N_2072,N_779,N_947);
and U2073 (N_2073,N_704,N_1194);
nand U2074 (N_2074,N_28,N_615);
nor U2075 (N_2075,N_642,N_71);
and U2076 (N_2076,N_170,N_918);
and U2077 (N_2077,N_1059,N_931);
xor U2078 (N_2078,N_806,N_587);
nand U2079 (N_2079,N_549,N_1260);
and U2080 (N_2080,N_884,N_688);
or U2081 (N_2081,N_1050,N_113);
or U2082 (N_2082,N_1164,N_852);
and U2083 (N_2083,N_885,N_1025);
and U2084 (N_2084,N_848,N_1425);
xnor U2085 (N_2085,N_1099,N_571);
or U2086 (N_2086,N_14,N_711);
and U2087 (N_2087,N_773,N_669);
nand U2088 (N_2088,N_973,N_713);
xnor U2089 (N_2089,N_378,N_489);
or U2090 (N_2090,N_830,N_618);
nor U2091 (N_2091,N_100,N_853);
nand U2092 (N_2092,N_578,N_960);
nand U2093 (N_2093,N_576,N_631);
or U2094 (N_2094,N_112,N_174);
nor U2095 (N_2095,N_919,N_513);
nor U2096 (N_2096,N_946,N_558);
xnor U2097 (N_2097,N_507,N_408);
xor U2098 (N_2098,N_415,N_1122);
nand U2099 (N_2099,N_130,N_1093);
and U2100 (N_2100,N_304,N_709);
or U2101 (N_2101,N_932,N_1252);
nor U2102 (N_2102,N_311,N_721);
nor U2103 (N_2103,N_1281,N_908);
nand U2104 (N_2104,N_554,N_371);
xnor U2105 (N_2105,N_134,N_1123);
or U2106 (N_2106,N_361,N_147);
nor U2107 (N_2107,N_38,N_807);
and U2108 (N_2108,N_903,N_128);
xor U2109 (N_2109,N_545,N_177);
nand U2110 (N_2110,N_161,N_244);
and U2111 (N_2111,N_1036,N_1372);
and U2112 (N_2112,N_610,N_1259);
or U2113 (N_2113,N_218,N_671);
or U2114 (N_2114,N_577,N_1307);
and U2115 (N_2115,N_256,N_1);
nor U2116 (N_2116,N_926,N_72);
xnor U2117 (N_2117,N_698,N_1320);
nor U2118 (N_2118,N_924,N_52);
nor U2119 (N_2119,N_74,N_102);
or U2120 (N_2120,N_428,N_504);
and U2121 (N_2121,N_1419,N_293);
xnor U2122 (N_2122,N_85,N_1495);
nand U2123 (N_2123,N_1438,N_977);
nand U2124 (N_2124,N_970,N_867);
nand U2125 (N_2125,N_1154,N_938);
xor U2126 (N_2126,N_58,N_160);
xor U2127 (N_2127,N_611,N_715);
nor U2128 (N_2128,N_1218,N_199);
and U2129 (N_2129,N_979,N_930);
xnor U2130 (N_2130,N_1070,N_226);
or U2131 (N_2131,N_1100,N_402);
nand U2132 (N_2132,N_862,N_445);
nor U2133 (N_2133,N_1338,N_614);
or U2134 (N_2134,N_79,N_1325);
or U2135 (N_2135,N_1363,N_1297);
or U2136 (N_2136,N_215,N_225);
xnor U2137 (N_2137,N_1481,N_448);
nand U2138 (N_2138,N_890,N_290);
and U2139 (N_2139,N_342,N_730);
nor U2140 (N_2140,N_1198,N_1151);
xor U2141 (N_2141,N_565,N_1157);
or U2142 (N_2142,N_1128,N_628);
or U2143 (N_2143,N_796,N_656);
xnor U2144 (N_2144,N_497,N_1152);
xor U2145 (N_2145,N_347,N_1008);
and U2146 (N_2146,N_1087,N_67);
or U2147 (N_2147,N_1301,N_534);
and U2148 (N_2148,N_251,N_1405);
nor U2149 (N_2149,N_599,N_674);
or U2150 (N_2150,N_340,N_1470);
and U2151 (N_2151,N_895,N_1083);
xnor U2152 (N_2152,N_1102,N_726);
nor U2153 (N_2153,N_1069,N_374);
nand U2154 (N_2154,N_416,N_394);
and U2155 (N_2155,N_1485,N_1162);
and U2156 (N_2156,N_372,N_1408);
or U2157 (N_2157,N_519,N_953);
nand U2158 (N_2158,N_237,N_1373);
xnor U2159 (N_2159,N_1195,N_1271);
or U2160 (N_2160,N_1267,N_1476);
and U2161 (N_2161,N_91,N_619);
or U2162 (N_2162,N_282,N_1448);
and U2163 (N_2163,N_475,N_452);
nor U2164 (N_2164,N_49,N_627);
nor U2165 (N_2165,N_1369,N_1103);
or U2166 (N_2166,N_1395,N_963);
nor U2167 (N_2167,N_826,N_667);
nand U2168 (N_2168,N_873,N_202);
and U2169 (N_2169,N_8,N_1493);
xnor U2170 (N_2170,N_1343,N_944);
nor U2171 (N_2171,N_538,N_598);
and U2172 (N_2172,N_728,N_1446);
nor U2173 (N_2173,N_126,N_213);
and U2174 (N_2174,N_1344,N_1228);
xor U2175 (N_2175,N_1002,N_383);
nand U2176 (N_2176,N_1479,N_905);
nand U2177 (N_2177,N_118,N_151);
and U2178 (N_2178,N_860,N_57);
and U2179 (N_2179,N_894,N_809);
and U2180 (N_2180,N_187,N_417);
xor U2181 (N_2181,N_292,N_664);
xor U2182 (N_2182,N_500,N_988);
xnor U2183 (N_2183,N_811,N_640);
or U2184 (N_2184,N_90,N_682);
or U2185 (N_2185,N_467,N_1215);
nand U2186 (N_2186,N_568,N_1472);
nor U2187 (N_2187,N_1085,N_791);
nor U2188 (N_2188,N_869,N_1149);
and U2189 (N_2189,N_949,N_1081);
xor U2190 (N_2190,N_871,N_291);
and U2191 (N_2191,N_1454,N_488);
nor U2192 (N_2192,N_385,N_722);
and U2193 (N_2193,N_399,N_1161);
nor U2194 (N_2194,N_1390,N_241);
xnor U2195 (N_2195,N_357,N_455);
nor U2196 (N_2196,N_1313,N_1480);
nand U2197 (N_2197,N_1006,N_437);
nor U2198 (N_2198,N_1013,N_1033);
and U2199 (N_2199,N_1047,N_1072);
nand U2200 (N_2200,N_1200,N_468);
or U2201 (N_2201,N_207,N_158);
nand U2202 (N_2202,N_1213,N_1189);
nor U2203 (N_2203,N_788,N_1014);
nand U2204 (N_2204,N_1141,N_1293);
nand U2205 (N_2205,N_1250,N_1176);
nor U2206 (N_2206,N_54,N_792);
xnor U2207 (N_2207,N_211,N_589);
and U2208 (N_2208,N_43,N_705);
nand U2209 (N_2209,N_191,N_776);
nor U2210 (N_2210,N_1178,N_582);
xnor U2211 (N_2211,N_1221,N_1156);
xnor U2212 (N_2212,N_532,N_980);
or U2213 (N_2213,N_583,N_162);
xor U2214 (N_2214,N_1391,N_480);
nor U2215 (N_2215,N_220,N_1236);
or U2216 (N_2216,N_987,N_1240);
nand U2217 (N_2217,N_32,N_590);
and U2218 (N_2218,N_1427,N_1165);
nor U2219 (N_2219,N_425,N_13);
nor U2220 (N_2220,N_493,N_1341);
or U2221 (N_2221,N_608,N_444);
xor U2222 (N_2222,N_1447,N_1468);
xnor U2223 (N_2223,N_1308,N_1295);
or U2224 (N_2224,N_1022,N_491);
or U2225 (N_2225,N_367,N_106);
xor U2226 (N_2226,N_1277,N_1350);
or U2227 (N_2227,N_1489,N_861);
and U2228 (N_2228,N_1357,N_363);
or U2229 (N_2229,N_1274,N_1169);
nand U2230 (N_2230,N_1089,N_1042);
nor U2231 (N_2231,N_1393,N_1235);
and U2232 (N_2232,N_414,N_178);
xnor U2233 (N_2233,N_1415,N_1136);
nor U2234 (N_2234,N_1276,N_799);
nor U2235 (N_2235,N_639,N_1409);
nand U2236 (N_2236,N_301,N_561);
nor U2237 (N_2237,N_315,N_509);
or U2238 (N_2238,N_593,N_543);
and U2239 (N_2239,N_835,N_778);
xor U2240 (N_2240,N_676,N_1312);
xnor U2241 (N_2241,N_1488,N_1253);
and U2242 (N_2242,N_1159,N_1181);
xnor U2243 (N_2243,N_483,N_369);
and U2244 (N_2244,N_454,N_384);
xor U2245 (N_2245,N_1091,N_1443);
nor U2246 (N_2246,N_936,N_624);
or U2247 (N_2247,N_783,N_1007);
nor U2248 (N_2248,N_221,N_1486);
xor U2249 (N_2249,N_1206,N_552);
nor U2250 (N_2250,N_973,N_440);
and U2251 (N_2251,N_461,N_977);
nand U2252 (N_2252,N_74,N_114);
nor U2253 (N_2253,N_1182,N_713);
or U2254 (N_2254,N_434,N_80);
or U2255 (N_2255,N_656,N_969);
or U2256 (N_2256,N_92,N_181);
nand U2257 (N_2257,N_121,N_860);
nor U2258 (N_2258,N_684,N_380);
nand U2259 (N_2259,N_742,N_1007);
xnor U2260 (N_2260,N_250,N_989);
and U2261 (N_2261,N_785,N_194);
and U2262 (N_2262,N_420,N_886);
or U2263 (N_2263,N_1162,N_479);
nand U2264 (N_2264,N_895,N_1407);
nand U2265 (N_2265,N_904,N_1045);
or U2266 (N_2266,N_897,N_4);
nand U2267 (N_2267,N_266,N_1093);
xnor U2268 (N_2268,N_689,N_1391);
nor U2269 (N_2269,N_640,N_1232);
nor U2270 (N_2270,N_602,N_739);
nand U2271 (N_2271,N_970,N_968);
or U2272 (N_2272,N_869,N_864);
nor U2273 (N_2273,N_889,N_159);
nor U2274 (N_2274,N_1318,N_838);
nor U2275 (N_2275,N_1323,N_1287);
and U2276 (N_2276,N_368,N_754);
and U2277 (N_2277,N_560,N_1488);
nand U2278 (N_2278,N_124,N_405);
nand U2279 (N_2279,N_220,N_362);
xnor U2280 (N_2280,N_30,N_196);
nand U2281 (N_2281,N_1359,N_960);
nor U2282 (N_2282,N_973,N_665);
or U2283 (N_2283,N_1371,N_1281);
nor U2284 (N_2284,N_876,N_654);
nand U2285 (N_2285,N_1484,N_1219);
nor U2286 (N_2286,N_461,N_974);
nand U2287 (N_2287,N_1087,N_1376);
and U2288 (N_2288,N_1474,N_792);
xnor U2289 (N_2289,N_1271,N_451);
or U2290 (N_2290,N_518,N_583);
or U2291 (N_2291,N_678,N_672);
nand U2292 (N_2292,N_324,N_1456);
and U2293 (N_2293,N_319,N_532);
or U2294 (N_2294,N_622,N_1289);
and U2295 (N_2295,N_633,N_381);
nor U2296 (N_2296,N_497,N_1412);
xnor U2297 (N_2297,N_671,N_1131);
nand U2298 (N_2298,N_789,N_614);
and U2299 (N_2299,N_27,N_913);
and U2300 (N_2300,N_393,N_838);
xnor U2301 (N_2301,N_729,N_791);
nand U2302 (N_2302,N_1037,N_184);
or U2303 (N_2303,N_737,N_766);
xnor U2304 (N_2304,N_187,N_356);
and U2305 (N_2305,N_308,N_111);
nor U2306 (N_2306,N_936,N_1325);
and U2307 (N_2307,N_681,N_819);
nor U2308 (N_2308,N_342,N_1448);
nand U2309 (N_2309,N_1246,N_29);
and U2310 (N_2310,N_299,N_678);
nor U2311 (N_2311,N_134,N_254);
and U2312 (N_2312,N_861,N_72);
and U2313 (N_2313,N_1052,N_506);
and U2314 (N_2314,N_460,N_237);
or U2315 (N_2315,N_221,N_197);
nand U2316 (N_2316,N_237,N_580);
nand U2317 (N_2317,N_987,N_353);
or U2318 (N_2318,N_707,N_32);
or U2319 (N_2319,N_560,N_368);
nor U2320 (N_2320,N_272,N_198);
or U2321 (N_2321,N_663,N_1409);
and U2322 (N_2322,N_368,N_195);
xnor U2323 (N_2323,N_481,N_644);
nor U2324 (N_2324,N_1071,N_1058);
or U2325 (N_2325,N_685,N_491);
and U2326 (N_2326,N_1183,N_1085);
and U2327 (N_2327,N_684,N_685);
nand U2328 (N_2328,N_921,N_1466);
xor U2329 (N_2329,N_758,N_913);
nor U2330 (N_2330,N_426,N_453);
and U2331 (N_2331,N_480,N_175);
or U2332 (N_2332,N_390,N_1456);
nand U2333 (N_2333,N_187,N_722);
nand U2334 (N_2334,N_190,N_512);
or U2335 (N_2335,N_539,N_126);
or U2336 (N_2336,N_164,N_1472);
and U2337 (N_2337,N_982,N_701);
nor U2338 (N_2338,N_276,N_845);
nand U2339 (N_2339,N_631,N_926);
xnor U2340 (N_2340,N_1209,N_709);
nor U2341 (N_2341,N_285,N_960);
nand U2342 (N_2342,N_1202,N_630);
nand U2343 (N_2343,N_519,N_123);
nand U2344 (N_2344,N_317,N_332);
xnor U2345 (N_2345,N_318,N_912);
nor U2346 (N_2346,N_602,N_429);
nor U2347 (N_2347,N_263,N_1283);
xor U2348 (N_2348,N_1480,N_1252);
nor U2349 (N_2349,N_185,N_237);
nor U2350 (N_2350,N_104,N_1353);
xnor U2351 (N_2351,N_1385,N_520);
nand U2352 (N_2352,N_923,N_1103);
and U2353 (N_2353,N_819,N_653);
nand U2354 (N_2354,N_691,N_1335);
nor U2355 (N_2355,N_342,N_892);
nand U2356 (N_2356,N_593,N_983);
nand U2357 (N_2357,N_1234,N_1093);
nor U2358 (N_2358,N_828,N_113);
xor U2359 (N_2359,N_1025,N_1447);
and U2360 (N_2360,N_902,N_882);
nand U2361 (N_2361,N_236,N_78);
nor U2362 (N_2362,N_808,N_1213);
xnor U2363 (N_2363,N_1135,N_1064);
and U2364 (N_2364,N_791,N_1063);
or U2365 (N_2365,N_663,N_1420);
and U2366 (N_2366,N_446,N_900);
xor U2367 (N_2367,N_346,N_717);
and U2368 (N_2368,N_1479,N_1411);
and U2369 (N_2369,N_393,N_1117);
or U2370 (N_2370,N_1093,N_327);
or U2371 (N_2371,N_1318,N_405);
xor U2372 (N_2372,N_210,N_153);
or U2373 (N_2373,N_389,N_1006);
nor U2374 (N_2374,N_201,N_220);
or U2375 (N_2375,N_549,N_329);
nand U2376 (N_2376,N_440,N_1081);
nand U2377 (N_2377,N_460,N_509);
and U2378 (N_2378,N_420,N_230);
or U2379 (N_2379,N_349,N_244);
nor U2380 (N_2380,N_70,N_835);
xor U2381 (N_2381,N_1248,N_1162);
or U2382 (N_2382,N_1326,N_223);
nand U2383 (N_2383,N_1429,N_366);
or U2384 (N_2384,N_817,N_1385);
or U2385 (N_2385,N_887,N_245);
or U2386 (N_2386,N_241,N_501);
or U2387 (N_2387,N_821,N_323);
or U2388 (N_2388,N_1358,N_812);
nand U2389 (N_2389,N_718,N_328);
and U2390 (N_2390,N_53,N_1372);
xor U2391 (N_2391,N_647,N_332);
and U2392 (N_2392,N_1377,N_137);
and U2393 (N_2393,N_714,N_542);
and U2394 (N_2394,N_553,N_457);
nor U2395 (N_2395,N_924,N_1119);
or U2396 (N_2396,N_1272,N_1400);
and U2397 (N_2397,N_644,N_1249);
or U2398 (N_2398,N_1137,N_274);
nor U2399 (N_2399,N_992,N_661);
and U2400 (N_2400,N_309,N_606);
nor U2401 (N_2401,N_815,N_441);
nor U2402 (N_2402,N_959,N_1023);
nand U2403 (N_2403,N_864,N_854);
xnor U2404 (N_2404,N_1121,N_411);
xor U2405 (N_2405,N_1053,N_581);
xor U2406 (N_2406,N_467,N_806);
nand U2407 (N_2407,N_1180,N_840);
nand U2408 (N_2408,N_598,N_241);
or U2409 (N_2409,N_746,N_1431);
or U2410 (N_2410,N_982,N_1249);
or U2411 (N_2411,N_1136,N_54);
nor U2412 (N_2412,N_1184,N_917);
xor U2413 (N_2413,N_1437,N_592);
xnor U2414 (N_2414,N_1118,N_336);
and U2415 (N_2415,N_790,N_907);
xor U2416 (N_2416,N_464,N_1482);
xor U2417 (N_2417,N_784,N_1124);
nand U2418 (N_2418,N_508,N_1397);
and U2419 (N_2419,N_405,N_991);
nand U2420 (N_2420,N_699,N_497);
or U2421 (N_2421,N_523,N_316);
xnor U2422 (N_2422,N_1059,N_83);
nand U2423 (N_2423,N_519,N_272);
and U2424 (N_2424,N_1360,N_431);
and U2425 (N_2425,N_1483,N_1443);
or U2426 (N_2426,N_234,N_791);
xnor U2427 (N_2427,N_837,N_407);
xor U2428 (N_2428,N_622,N_1299);
and U2429 (N_2429,N_765,N_245);
or U2430 (N_2430,N_1415,N_425);
or U2431 (N_2431,N_1108,N_24);
or U2432 (N_2432,N_792,N_205);
nand U2433 (N_2433,N_1368,N_392);
nand U2434 (N_2434,N_409,N_73);
nand U2435 (N_2435,N_520,N_957);
or U2436 (N_2436,N_485,N_522);
nor U2437 (N_2437,N_1009,N_1337);
and U2438 (N_2438,N_114,N_1261);
or U2439 (N_2439,N_1457,N_1072);
nand U2440 (N_2440,N_739,N_981);
xor U2441 (N_2441,N_1269,N_573);
nand U2442 (N_2442,N_943,N_28);
xor U2443 (N_2443,N_92,N_1336);
and U2444 (N_2444,N_200,N_780);
nand U2445 (N_2445,N_896,N_1461);
nand U2446 (N_2446,N_284,N_9);
and U2447 (N_2447,N_609,N_492);
nand U2448 (N_2448,N_1444,N_614);
or U2449 (N_2449,N_897,N_268);
nand U2450 (N_2450,N_325,N_23);
nand U2451 (N_2451,N_535,N_134);
xnor U2452 (N_2452,N_676,N_1468);
or U2453 (N_2453,N_1433,N_1076);
and U2454 (N_2454,N_1275,N_356);
nor U2455 (N_2455,N_853,N_626);
nor U2456 (N_2456,N_1068,N_873);
nand U2457 (N_2457,N_832,N_1413);
or U2458 (N_2458,N_105,N_333);
or U2459 (N_2459,N_325,N_795);
or U2460 (N_2460,N_410,N_1456);
and U2461 (N_2461,N_8,N_395);
and U2462 (N_2462,N_954,N_383);
xor U2463 (N_2463,N_1096,N_529);
or U2464 (N_2464,N_1408,N_743);
nand U2465 (N_2465,N_941,N_964);
or U2466 (N_2466,N_855,N_937);
and U2467 (N_2467,N_867,N_512);
nor U2468 (N_2468,N_758,N_428);
or U2469 (N_2469,N_451,N_205);
nand U2470 (N_2470,N_258,N_1030);
nand U2471 (N_2471,N_268,N_1448);
nor U2472 (N_2472,N_798,N_1065);
or U2473 (N_2473,N_907,N_1099);
xnor U2474 (N_2474,N_1125,N_1198);
and U2475 (N_2475,N_899,N_1270);
nor U2476 (N_2476,N_408,N_595);
or U2477 (N_2477,N_608,N_1089);
and U2478 (N_2478,N_231,N_17);
nor U2479 (N_2479,N_422,N_905);
or U2480 (N_2480,N_192,N_1140);
and U2481 (N_2481,N_154,N_222);
nor U2482 (N_2482,N_117,N_706);
xnor U2483 (N_2483,N_130,N_520);
nand U2484 (N_2484,N_371,N_1481);
nor U2485 (N_2485,N_10,N_1211);
nand U2486 (N_2486,N_1148,N_234);
nor U2487 (N_2487,N_24,N_949);
nand U2488 (N_2488,N_951,N_6);
or U2489 (N_2489,N_321,N_93);
or U2490 (N_2490,N_540,N_65);
and U2491 (N_2491,N_335,N_762);
nor U2492 (N_2492,N_609,N_1073);
nand U2493 (N_2493,N_1463,N_746);
nor U2494 (N_2494,N_1171,N_1071);
nor U2495 (N_2495,N_681,N_1341);
nor U2496 (N_2496,N_39,N_615);
nor U2497 (N_2497,N_9,N_317);
nand U2498 (N_2498,N_1160,N_1477);
nor U2499 (N_2499,N_1018,N_517);
and U2500 (N_2500,N_1314,N_234);
nand U2501 (N_2501,N_89,N_272);
or U2502 (N_2502,N_1457,N_1356);
xnor U2503 (N_2503,N_142,N_1310);
nor U2504 (N_2504,N_525,N_1064);
nor U2505 (N_2505,N_1396,N_544);
xnor U2506 (N_2506,N_191,N_116);
xnor U2507 (N_2507,N_809,N_822);
or U2508 (N_2508,N_1137,N_961);
nor U2509 (N_2509,N_307,N_771);
xnor U2510 (N_2510,N_550,N_1089);
and U2511 (N_2511,N_382,N_812);
and U2512 (N_2512,N_685,N_372);
or U2513 (N_2513,N_763,N_187);
nor U2514 (N_2514,N_23,N_461);
nor U2515 (N_2515,N_1014,N_895);
nor U2516 (N_2516,N_873,N_560);
xor U2517 (N_2517,N_66,N_336);
or U2518 (N_2518,N_1060,N_837);
and U2519 (N_2519,N_549,N_1432);
or U2520 (N_2520,N_929,N_961);
nand U2521 (N_2521,N_319,N_1220);
and U2522 (N_2522,N_628,N_391);
xor U2523 (N_2523,N_9,N_1148);
nor U2524 (N_2524,N_743,N_156);
xnor U2525 (N_2525,N_512,N_409);
and U2526 (N_2526,N_1149,N_479);
and U2527 (N_2527,N_1474,N_1296);
and U2528 (N_2528,N_1384,N_480);
xor U2529 (N_2529,N_1128,N_505);
nand U2530 (N_2530,N_32,N_338);
nand U2531 (N_2531,N_1227,N_1091);
nor U2532 (N_2532,N_365,N_350);
or U2533 (N_2533,N_1308,N_1251);
xnor U2534 (N_2534,N_250,N_171);
and U2535 (N_2535,N_944,N_90);
or U2536 (N_2536,N_1409,N_650);
and U2537 (N_2537,N_387,N_584);
nand U2538 (N_2538,N_1360,N_978);
and U2539 (N_2539,N_786,N_200);
or U2540 (N_2540,N_1330,N_1489);
xnor U2541 (N_2541,N_1396,N_389);
nand U2542 (N_2542,N_1372,N_1380);
nand U2543 (N_2543,N_50,N_550);
nand U2544 (N_2544,N_790,N_548);
xnor U2545 (N_2545,N_555,N_112);
xor U2546 (N_2546,N_365,N_556);
and U2547 (N_2547,N_852,N_400);
nor U2548 (N_2548,N_214,N_611);
nand U2549 (N_2549,N_276,N_204);
and U2550 (N_2550,N_414,N_860);
nand U2551 (N_2551,N_1491,N_676);
nor U2552 (N_2552,N_241,N_672);
nand U2553 (N_2553,N_120,N_956);
or U2554 (N_2554,N_596,N_1259);
nor U2555 (N_2555,N_752,N_1048);
or U2556 (N_2556,N_496,N_895);
nor U2557 (N_2557,N_479,N_900);
nand U2558 (N_2558,N_420,N_1258);
nand U2559 (N_2559,N_1334,N_1037);
xnor U2560 (N_2560,N_549,N_673);
nor U2561 (N_2561,N_156,N_1487);
xnor U2562 (N_2562,N_1211,N_797);
and U2563 (N_2563,N_1387,N_855);
nand U2564 (N_2564,N_377,N_423);
nor U2565 (N_2565,N_1344,N_421);
nor U2566 (N_2566,N_421,N_1383);
nand U2567 (N_2567,N_1036,N_972);
or U2568 (N_2568,N_194,N_1221);
or U2569 (N_2569,N_1088,N_367);
or U2570 (N_2570,N_1084,N_10);
xor U2571 (N_2571,N_1041,N_1249);
nand U2572 (N_2572,N_1039,N_361);
or U2573 (N_2573,N_1404,N_273);
and U2574 (N_2574,N_419,N_924);
nor U2575 (N_2575,N_158,N_604);
and U2576 (N_2576,N_1268,N_393);
xnor U2577 (N_2577,N_233,N_1484);
nor U2578 (N_2578,N_344,N_1310);
or U2579 (N_2579,N_1378,N_887);
xnor U2580 (N_2580,N_1097,N_451);
nor U2581 (N_2581,N_599,N_880);
nand U2582 (N_2582,N_1256,N_723);
or U2583 (N_2583,N_347,N_733);
nand U2584 (N_2584,N_1369,N_955);
nor U2585 (N_2585,N_1082,N_1155);
nand U2586 (N_2586,N_139,N_247);
nor U2587 (N_2587,N_1286,N_890);
nand U2588 (N_2588,N_347,N_1452);
and U2589 (N_2589,N_95,N_1480);
nor U2590 (N_2590,N_727,N_418);
nand U2591 (N_2591,N_1219,N_952);
xor U2592 (N_2592,N_1476,N_974);
nor U2593 (N_2593,N_459,N_410);
nand U2594 (N_2594,N_1350,N_488);
nor U2595 (N_2595,N_264,N_726);
and U2596 (N_2596,N_148,N_1193);
and U2597 (N_2597,N_394,N_1234);
nor U2598 (N_2598,N_1313,N_721);
nor U2599 (N_2599,N_1285,N_1023);
nand U2600 (N_2600,N_305,N_843);
nor U2601 (N_2601,N_250,N_735);
and U2602 (N_2602,N_505,N_1283);
xor U2603 (N_2603,N_925,N_977);
and U2604 (N_2604,N_379,N_479);
or U2605 (N_2605,N_1085,N_1495);
nor U2606 (N_2606,N_705,N_1060);
xor U2607 (N_2607,N_377,N_1496);
nand U2608 (N_2608,N_335,N_355);
nand U2609 (N_2609,N_1227,N_1150);
nor U2610 (N_2610,N_1131,N_850);
xor U2611 (N_2611,N_1372,N_114);
and U2612 (N_2612,N_185,N_1437);
nand U2613 (N_2613,N_724,N_1132);
nor U2614 (N_2614,N_655,N_599);
nor U2615 (N_2615,N_201,N_525);
and U2616 (N_2616,N_1069,N_939);
nand U2617 (N_2617,N_812,N_1240);
or U2618 (N_2618,N_1206,N_752);
and U2619 (N_2619,N_258,N_1117);
and U2620 (N_2620,N_421,N_640);
nand U2621 (N_2621,N_978,N_657);
nor U2622 (N_2622,N_1159,N_854);
nand U2623 (N_2623,N_475,N_719);
nor U2624 (N_2624,N_647,N_1376);
xor U2625 (N_2625,N_724,N_660);
nor U2626 (N_2626,N_732,N_591);
nor U2627 (N_2627,N_536,N_277);
nor U2628 (N_2628,N_1415,N_528);
nand U2629 (N_2629,N_424,N_1286);
nor U2630 (N_2630,N_1092,N_660);
nor U2631 (N_2631,N_161,N_798);
xnor U2632 (N_2632,N_972,N_1141);
xnor U2633 (N_2633,N_202,N_1146);
or U2634 (N_2634,N_1334,N_567);
xor U2635 (N_2635,N_357,N_1441);
nor U2636 (N_2636,N_816,N_410);
nand U2637 (N_2637,N_892,N_378);
or U2638 (N_2638,N_617,N_416);
nand U2639 (N_2639,N_367,N_379);
and U2640 (N_2640,N_529,N_928);
xor U2641 (N_2641,N_1113,N_1334);
xnor U2642 (N_2642,N_505,N_523);
nor U2643 (N_2643,N_1210,N_391);
xor U2644 (N_2644,N_133,N_27);
nand U2645 (N_2645,N_185,N_10);
nor U2646 (N_2646,N_363,N_157);
nand U2647 (N_2647,N_1297,N_246);
or U2648 (N_2648,N_838,N_750);
nor U2649 (N_2649,N_1257,N_72);
or U2650 (N_2650,N_143,N_633);
or U2651 (N_2651,N_905,N_1344);
and U2652 (N_2652,N_816,N_187);
or U2653 (N_2653,N_1023,N_199);
and U2654 (N_2654,N_265,N_503);
and U2655 (N_2655,N_612,N_1131);
and U2656 (N_2656,N_646,N_158);
nand U2657 (N_2657,N_472,N_833);
or U2658 (N_2658,N_1273,N_1148);
or U2659 (N_2659,N_371,N_1336);
or U2660 (N_2660,N_1466,N_989);
or U2661 (N_2661,N_704,N_644);
and U2662 (N_2662,N_380,N_1239);
xnor U2663 (N_2663,N_1438,N_698);
nand U2664 (N_2664,N_596,N_285);
nand U2665 (N_2665,N_224,N_1187);
nor U2666 (N_2666,N_1140,N_1342);
or U2667 (N_2667,N_577,N_283);
or U2668 (N_2668,N_959,N_340);
or U2669 (N_2669,N_1105,N_684);
nand U2670 (N_2670,N_1108,N_538);
and U2671 (N_2671,N_491,N_1333);
xnor U2672 (N_2672,N_1432,N_1007);
or U2673 (N_2673,N_183,N_1454);
and U2674 (N_2674,N_687,N_23);
or U2675 (N_2675,N_1181,N_985);
xor U2676 (N_2676,N_1113,N_751);
nor U2677 (N_2677,N_32,N_669);
xor U2678 (N_2678,N_775,N_1058);
or U2679 (N_2679,N_92,N_830);
nand U2680 (N_2680,N_1243,N_1211);
and U2681 (N_2681,N_777,N_303);
nand U2682 (N_2682,N_818,N_1025);
nor U2683 (N_2683,N_1215,N_947);
or U2684 (N_2684,N_768,N_1076);
nor U2685 (N_2685,N_1494,N_152);
and U2686 (N_2686,N_210,N_807);
nor U2687 (N_2687,N_1162,N_438);
nand U2688 (N_2688,N_871,N_341);
and U2689 (N_2689,N_1328,N_576);
and U2690 (N_2690,N_344,N_943);
and U2691 (N_2691,N_1340,N_34);
nand U2692 (N_2692,N_1283,N_224);
nor U2693 (N_2693,N_897,N_895);
nand U2694 (N_2694,N_1,N_775);
and U2695 (N_2695,N_1281,N_1397);
nand U2696 (N_2696,N_189,N_581);
or U2697 (N_2697,N_1462,N_674);
or U2698 (N_2698,N_268,N_1149);
nand U2699 (N_2699,N_1088,N_241);
and U2700 (N_2700,N_754,N_882);
and U2701 (N_2701,N_734,N_1443);
nand U2702 (N_2702,N_1317,N_1124);
or U2703 (N_2703,N_1378,N_187);
or U2704 (N_2704,N_356,N_1265);
and U2705 (N_2705,N_453,N_1189);
nand U2706 (N_2706,N_1353,N_60);
or U2707 (N_2707,N_870,N_421);
xnor U2708 (N_2708,N_1042,N_1408);
nand U2709 (N_2709,N_523,N_368);
or U2710 (N_2710,N_7,N_51);
and U2711 (N_2711,N_180,N_358);
xnor U2712 (N_2712,N_595,N_218);
xnor U2713 (N_2713,N_302,N_1173);
nand U2714 (N_2714,N_1148,N_613);
and U2715 (N_2715,N_710,N_432);
nand U2716 (N_2716,N_401,N_453);
nand U2717 (N_2717,N_1146,N_388);
xnor U2718 (N_2718,N_1430,N_18);
and U2719 (N_2719,N_627,N_79);
or U2720 (N_2720,N_1191,N_1384);
xor U2721 (N_2721,N_1325,N_925);
nand U2722 (N_2722,N_669,N_800);
and U2723 (N_2723,N_1069,N_1477);
or U2724 (N_2724,N_715,N_276);
and U2725 (N_2725,N_905,N_810);
xnor U2726 (N_2726,N_1322,N_634);
nand U2727 (N_2727,N_885,N_556);
or U2728 (N_2728,N_826,N_96);
xor U2729 (N_2729,N_728,N_378);
nand U2730 (N_2730,N_124,N_174);
nor U2731 (N_2731,N_872,N_319);
and U2732 (N_2732,N_1015,N_1052);
nand U2733 (N_2733,N_1170,N_968);
and U2734 (N_2734,N_786,N_908);
nor U2735 (N_2735,N_195,N_993);
or U2736 (N_2736,N_460,N_1013);
or U2737 (N_2737,N_82,N_915);
nand U2738 (N_2738,N_1014,N_1367);
or U2739 (N_2739,N_574,N_848);
and U2740 (N_2740,N_1273,N_172);
nand U2741 (N_2741,N_440,N_1443);
xor U2742 (N_2742,N_1495,N_1250);
nor U2743 (N_2743,N_1135,N_1323);
nand U2744 (N_2744,N_281,N_1006);
nand U2745 (N_2745,N_288,N_27);
nor U2746 (N_2746,N_777,N_341);
nor U2747 (N_2747,N_66,N_45);
nor U2748 (N_2748,N_1325,N_212);
and U2749 (N_2749,N_721,N_216);
xnor U2750 (N_2750,N_1276,N_87);
nand U2751 (N_2751,N_1124,N_1284);
or U2752 (N_2752,N_449,N_566);
or U2753 (N_2753,N_1100,N_631);
nor U2754 (N_2754,N_1096,N_330);
xnor U2755 (N_2755,N_54,N_359);
xnor U2756 (N_2756,N_363,N_64);
nand U2757 (N_2757,N_742,N_190);
xor U2758 (N_2758,N_1288,N_168);
nand U2759 (N_2759,N_714,N_796);
xnor U2760 (N_2760,N_1183,N_22);
xnor U2761 (N_2761,N_1365,N_100);
nor U2762 (N_2762,N_915,N_1302);
nor U2763 (N_2763,N_42,N_1066);
xnor U2764 (N_2764,N_641,N_1361);
xnor U2765 (N_2765,N_266,N_697);
or U2766 (N_2766,N_867,N_252);
nor U2767 (N_2767,N_1324,N_317);
xor U2768 (N_2768,N_623,N_1040);
or U2769 (N_2769,N_191,N_817);
xnor U2770 (N_2770,N_658,N_954);
nand U2771 (N_2771,N_1088,N_1058);
or U2772 (N_2772,N_962,N_238);
or U2773 (N_2773,N_389,N_1167);
nor U2774 (N_2774,N_406,N_1437);
and U2775 (N_2775,N_102,N_964);
xnor U2776 (N_2776,N_930,N_725);
and U2777 (N_2777,N_888,N_82);
nand U2778 (N_2778,N_25,N_1243);
xnor U2779 (N_2779,N_447,N_1029);
and U2780 (N_2780,N_895,N_1137);
and U2781 (N_2781,N_1355,N_1160);
or U2782 (N_2782,N_436,N_421);
nand U2783 (N_2783,N_926,N_91);
or U2784 (N_2784,N_395,N_250);
nand U2785 (N_2785,N_856,N_503);
nand U2786 (N_2786,N_265,N_239);
or U2787 (N_2787,N_1259,N_234);
and U2788 (N_2788,N_931,N_1319);
or U2789 (N_2789,N_796,N_95);
and U2790 (N_2790,N_961,N_1074);
or U2791 (N_2791,N_1104,N_1221);
xor U2792 (N_2792,N_64,N_1280);
or U2793 (N_2793,N_738,N_314);
xor U2794 (N_2794,N_494,N_65);
nand U2795 (N_2795,N_59,N_1055);
and U2796 (N_2796,N_4,N_71);
xor U2797 (N_2797,N_873,N_618);
xnor U2798 (N_2798,N_226,N_568);
xnor U2799 (N_2799,N_347,N_1050);
xor U2800 (N_2800,N_53,N_1045);
xor U2801 (N_2801,N_292,N_803);
nand U2802 (N_2802,N_606,N_538);
nand U2803 (N_2803,N_897,N_1385);
xnor U2804 (N_2804,N_1432,N_428);
and U2805 (N_2805,N_1371,N_259);
and U2806 (N_2806,N_725,N_1399);
nand U2807 (N_2807,N_1012,N_1380);
and U2808 (N_2808,N_660,N_518);
nand U2809 (N_2809,N_491,N_687);
xor U2810 (N_2810,N_667,N_728);
xnor U2811 (N_2811,N_1203,N_850);
nor U2812 (N_2812,N_719,N_1287);
or U2813 (N_2813,N_1173,N_533);
nor U2814 (N_2814,N_842,N_1424);
nor U2815 (N_2815,N_66,N_323);
and U2816 (N_2816,N_108,N_616);
and U2817 (N_2817,N_257,N_448);
xnor U2818 (N_2818,N_174,N_292);
and U2819 (N_2819,N_371,N_313);
or U2820 (N_2820,N_165,N_527);
and U2821 (N_2821,N_315,N_991);
or U2822 (N_2822,N_308,N_307);
xor U2823 (N_2823,N_344,N_785);
or U2824 (N_2824,N_746,N_962);
and U2825 (N_2825,N_848,N_1214);
xor U2826 (N_2826,N_498,N_637);
nand U2827 (N_2827,N_633,N_248);
or U2828 (N_2828,N_1152,N_14);
nor U2829 (N_2829,N_377,N_1435);
and U2830 (N_2830,N_1486,N_409);
nor U2831 (N_2831,N_555,N_103);
nand U2832 (N_2832,N_1085,N_680);
xor U2833 (N_2833,N_909,N_488);
nand U2834 (N_2834,N_598,N_379);
and U2835 (N_2835,N_1371,N_202);
nor U2836 (N_2836,N_415,N_872);
xnor U2837 (N_2837,N_586,N_1309);
nor U2838 (N_2838,N_1202,N_140);
or U2839 (N_2839,N_755,N_738);
nand U2840 (N_2840,N_1161,N_1190);
or U2841 (N_2841,N_1315,N_971);
and U2842 (N_2842,N_731,N_64);
nand U2843 (N_2843,N_295,N_372);
or U2844 (N_2844,N_1171,N_1405);
and U2845 (N_2845,N_1069,N_732);
nand U2846 (N_2846,N_1167,N_965);
nand U2847 (N_2847,N_915,N_882);
nor U2848 (N_2848,N_385,N_263);
nor U2849 (N_2849,N_412,N_406);
and U2850 (N_2850,N_1289,N_950);
or U2851 (N_2851,N_1080,N_785);
xor U2852 (N_2852,N_497,N_507);
nand U2853 (N_2853,N_85,N_350);
nor U2854 (N_2854,N_362,N_520);
and U2855 (N_2855,N_964,N_1051);
or U2856 (N_2856,N_1261,N_155);
nand U2857 (N_2857,N_1313,N_532);
or U2858 (N_2858,N_1404,N_1147);
and U2859 (N_2859,N_1462,N_1);
nor U2860 (N_2860,N_1338,N_1051);
nor U2861 (N_2861,N_599,N_195);
nand U2862 (N_2862,N_1272,N_1119);
nand U2863 (N_2863,N_1065,N_1342);
nor U2864 (N_2864,N_332,N_1185);
xor U2865 (N_2865,N_31,N_1157);
and U2866 (N_2866,N_806,N_197);
or U2867 (N_2867,N_970,N_548);
nand U2868 (N_2868,N_825,N_1023);
xor U2869 (N_2869,N_1345,N_557);
nand U2870 (N_2870,N_700,N_1102);
nor U2871 (N_2871,N_1349,N_695);
or U2872 (N_2872,N_1286,N_100);
nand U2873 (N_2873,N_212,N_1230);
or U2874 (N_2874,N_1023,N_995);
and U2875 (N_2875,N_1420,N_60);
xnor U2876 (N_2876,N_673,N_652);
nand U2877 (N_2877,N_294,N_546);
nor U2878 (N_2878,N_1231,N_59);
and U2879 (N_2879,N_277,N_235);
xnor U2880 (N_2880,N_1105,N_928);
and U2881 (N_2881,N_1492,N_317);
nor U2882 (N_2882,N_1153,N_81);
and U2883 (N_2883,N_266,N_1010);
and U2884 (N_2884,N_1482,N_1121);
and U2885 (N_2885,N_124,N_680);
or U2886 (N_2886,N_1321,N_1147);
xor U2887 (N_2887,N_125,N_1173);
nor U2888 (N_2888,N_1116,N_651);
or U2889 (N_2889,N_90,N_268);
nand U2890 (N_2890,N_1086,N_1456);
nand U2891 (N_2891,N_1082,N_586);
nand U2892 (N_2892,N_474,N_77);
or U2893 (N_2893,N_1005,N_784);
or U2894 (N_2894,N_918,N_755);
nand U2895 (N_2895,N_461,N_365);
nand U2896 (N_2896,N_734,N_857);
or U2897 (N_2897,N_1265,N_1019);
nand U2898 (N_2898,N_139,N_434);
nand U2899 (N_2899,N_442,N_118);
nand U2900 (N_2900,N_42,N_368);
nor U2901 (N_2901,N_328,N_497);
nand U2902 (N_2902,N_254,N_676);
nand U2903 (N_2903,N_1123,N_1068);
or U2904 (N_2904,N_652,N_584);
or U2905 (N_2905,N_397,N_1030);
or U2906 (N_2906,N_446,N_285);
nand U2907 (N_2907,N_1270,N_1152);
nor U2908 (N_2908,N_635,N_211);
nand U2909 (N_2909,N_456,N_958);
xnor U2910 (N_2910,N_1268,N_1122);
and U2911 (N_2911,N_477,N_513);
and U2912 (N_2912,N_203,N_1161);
xor U2913 (N_2913,N_684,N_238);
xnor U2914 (N_2914,N_1466,N_422);
nor U2915 (N_2915,N_254,N_921);
nand U2916 (N_2916,N_12,N_191);
or U2917 (N_2917,N_1345,N_685);
xor U2918 (N_2918,N_1360,N_1398);
nor U2919 (N_2919,N_115,N_969);
nand U2920 (N_2920,N_320,N_367);
and U2921 (N_2921,N_1278,N_227);
xor U2922 (N_2922,N_501,N_1302);
or U2923 (N_2923,N_335,N_1477);
nor U2924 (N_2924,N_601,N_124);
and U2925 (N_2925,N_654,N_42);
xnor U2926 (N_2926,N_581,N_1344);
xnor U2927 (N_2927,N_550,N_1489);
and U2928 (N_2928,N_1230,N_741);
or U2929 (N_2929,N_1371,N_323);
and U2930 (N_2930,N_502,N_1378);
or U2931 (N_2931,N_1204,N_597);
xor U2932 (N_2932,N_362,N_1305);
xor U2933 (N_2933,N_948,N_824);
xor U2934 (N_2934,N_364,N_111);
nand U2935 (N_2935,N_657,N_447);
or U2936 (N_2936,N_382,N_180);
and U2937 (N_2937,N_350,N_103);
xnor U2938 (N_2938,N_781,N_498);
nand U2939 (N_2939,N_78,N_909);
and U2940 (N_2940,N_19,N_503);
xor U2941 (N_2941,N_126,N_258);
and U2942 (N_2942,N_1045,N_1493);
nand U2943 (N_2943,N_1034,N_843);
xor U2944 (N_2944,N_1479,N_922);
xnor U2945 (N_2945,N_42,N_752);
nor U2946 (N_2946,N_1309,N_859);
xor U2947 (N_2947,N_777,N_37);
nand U2948 (N_2948,N_683,N_657);
nand U2949 (N_2949,N_676,N_1286);
and U2950 (N_2950,N_771,N_748);
or U2951 (N_2951,N_1127,N_881);
nor U2952 (N_2952,N_509,N_244);
and U2953 (N_2953,N_1335,N_91);
and U2954 (N_2954,N_1141,N_684);
nor U2955 (N_2955,N_885,N_276);
xor U2956 (N_2956,N_693,N_257);
xnor U2957 (N_2957,N_59,N_1337);
and U2958 (N_2958,N_1312,N_1002);
nand U2959 (N_2959,N_1217,N_1031);
and U2960 (N_2960,N_342,N_764);
or U2961 (N_2961,N_543,N_106);
nand U2962 (N_2962,N_834,N_204);
or U2963 (N_2963,N_860,N_777);
nand U2964 (N_2964,N_293,N_1450);
and U2965 (N_2965,N_538,N_135);
or U2966 (N_2966,N_291,N_522);
xnor U2967 (N_2967,N_534,N_632);
nand U2968 (N_2968,N_865,N_1180);
nand U2969 (N_2969,N_680,N_644);
xor U2970 (N_2970,N_154,N_308);
xor U2971 (N_2971,N_456,N_94);
or U2972 (N_2972,N_1026,N_1203);
nor U2973 (N_2973,N_379,N_834);
nand U2974 (N_2974,N_1396,N_1400);
xnor U2975 (N_2975,N_1184,N_839);
nand U2976 (N_2976,N_416,N_124);
nand U2977 (N_2977,N_1335,N_1002);
or U2978 (N_2978,N_83,N_658);
nor U2979 (N_2979,N_1317,N_742);
nand U2980 (N_2980,N_1278,N_715);
or U2981 (N_2981,N_805,N_894);
xnor U2982 (N_2982,N_674,N_1057);
nor U2983 (N_2983,N_947,N_1043);
xnor U2984 (N_2984,N_721,N_1366);
and U2985 (N_2985,N_720,N_1332);
nor U2986 (N_2986,N_1111,N_468);
xnor U2987 (N_2987,N_995,N_1054);
nor U2988 (N_2988,N_779,N_1305);
xnor U2989 (N_2989,N_472,N_508);
or U2990 (N_2990,N_828,N_152);
xor U2991 (N_2991,N_632,N_295);
xnor U2992 (N_2992,N_639,N_536);
nand U2993 (N_2993,N_139,N_104);
or U2994 (N_2994,N_1005,N_1445);
and U2995 (N_2995,N_67,N_498);
xnor U2996 (N_2996,N_554,N_876);
and U2997 (N_2997,N_1352,N_1442);
nor U2998 (N_2998,N_1195,N_793);
xnor U2999 (N_2999,N_1014,N_1423);
xnor U3000 (N_3000,N_1879,N_2551);
nand U3001 (N_3001,N_1882,N_2255);
and U3002 (N_3002,N_2933,N_2595);
xnor U3003 (N_3003,N_2567,N_1549);
nand U3004 (N_3004,N_2548,N_2001);
nor U3005 (N_3005,N_2151,N_1834);
nand U3006 (N_3006,N_2161,N_2513);
or U3007 (N_3007,N_2679,N_1802);
nor U3008 (N_3008,N_2114,N_2714);
or U3009 (N_3009,N_2423,N_1575);
nor U3010 (N_3010,N_1610,N_1536);
nor U3011 (N_3011,N_2015,N_2352);
nand U3012 (N_3012,N_2484,N_2462);
nand U3013 (N_3013,N_2380,N_2887);
and U3014 (N_3014,N_2691,N_1939);
or U3015 (N_3015,N_2522,N_1772);
and U3016 (N_3016,N_2978,N_2160);
xnor U3017 (N_3017,N_1754,N_1698);
and U3018 (N_3018,N_2018,N_1700);
nand U3019 (N_3019,N_2372,N_2844);
xnor U3020 (N_3020,N_1823,N_2331);
nand U3021 (N_3021,N_1524,N_2743);
and U3022 (N_3022,N_1737,N_2807);
nand U3023 (N_3023,N_2702,N_2362);
xnor U3024 (N_3024,N_1675,N_1613);
nand U3025 (N_3025,N_2623,N_2611);
nor U3026 (N_3026,N_1629,N_2002);
nor U3027 (N_3027,N_2802,N_2070);
or U3028 (N_3028,N_1544,N_1909);
or U3029 (N_3029,N_1605,N_2606);
or U3030 (N_3030,N_2646,N_2040);
nand U3031 (N_3031,N_1692,N_1586);
or U3032 (N_3032,N_2856,N_2428);
and U3033 (N_3033,N_2073,N_2483);
and U3034 (N_3034,N_2539,N_2816);
nor U3035 (N_3035,N_2089,N_1975);
xnor U3036 (N_3036,N_1896,N_2562);
and U3037 (N_3037,N_2569,N_2166);
xor U3038 (N_3038,N_1506,N_2011);
and U3039 (N_3039,N_1827,N_2666);
nor U3040 (N_3040,N_2659,N_2368);
nand U3041 (N_3041,N_1602,N_2045);
and U3042 (N_3042,N_1601,N_1887);
and U3043 (N_3043,N_2808,N_2062);
nor U3044 (N_3044,N_2051,N_1820);
nand U3045 (N_3045,N_2655,N_2261);
or U3046 (N_3046,N_2007,N_2330);
and U3047 (N_3047,N_1580,N_2192);
and U3048 (N_3048,N_2609,N_2396);
nor U3049 (N_3049,N_2535,N_2039);
or U3050 (N_3050,N_1951,N_1910);
xnor U3051 (N_3051,N_1835,N_1952);
nor U3052 (N_3052,N_1640,N_2306);
xor U3053 (N_3053,N_2767,N_2892);
xor U3054 (N_3054,N_2476,N_2030);
nor U3055 (N_3055,N_1664,N_2193);
nand U3056 (N_3056,N_2194,N_2132);
nor U3057 (N_3057,N_1831,N_1670);
and U3058 (N_3058,N_2176,N_2218);
nand U3059 (N_3059,N_2232,N_2208);
nor U3060 (N_3060,N_1574,N_2849);
nand U3061 (N_3061,N_2478,N_2399);
xor U3062 (N_3062,N_2093,N_2204);
nor U3063 (N_3063,N_2515,N_2966);
nor U3064 (N_3064,N_2628,N_1609);
nand U3065 (N_3065,N_1761,N_1563);
nor U3066 (N_3066,N_2601,N_2980);
or U3067 (N_3067,N_1732,N_2867);
xor U3068 (N_3068,N_1866,N_2509);
nor U3069 (N_3069,N_2963,N_1805);
nand U3070 (N_3070,N_2727,N_2458);
nor U3071 (N_3071,N_1983,N_1763);
nand U3072 (N_3072,N_1890,N_2741);
nand U3073 (N_3073,N_2146,N_2185);
xor U3074 (N_3074,N_1936,N_2793);
xor U3075 (N_3075,N_1961,N_2181);
and U3076 (N_3076,N_1571,N_2481);
xor U3077 (N_3077,N_2106,N_1713);
xnor U3078 (N_3078,N_2141,N_2069);
nor U3079 (N_3079,N_1949,N_1541);
or U3080 (N_3080,N_2454,N_1944);
xor U3081 (N_3081,N_2612,N_2416);
xor U3082 (N_3082,N_2775,N_1870);
nor U3083 (N_3083,N_2426,N_1703);
and U3084 (N_3084,N_1976,N_2742);
nand U3085 (N_3085,N_2855,N_2046);
nand U3086 (N_3086,N_1899,N_1766);
nor U3087 (N_3087,N_1616,N_2836);
and U3088 (N_3088,N_2044,N_1567);
or U3089 (N_3089,N_2578,N_1511);
or U3090 (N_3090,N_2709,N_1998);
and U3091 (N_3091,N_2550,N_1717);
nor U3092 (N_3092,N_1893,N_2603);
nor U3093 (N_3093,N_1597,N_2494);
xnor U3094 (N_3094,N_2697,N_2170);
and U3095 (N_3095,N_2957,N_2005);
nor U3096 (N_3096,N_2252,N_1514);
nand U3097 (N_3097,N_2489,N_1735);
nand U3098 (N_3098,N_1897,N_2173);
nor U3099 (N_3099,N_2427,N_2640);
and U3100 (N_3100,N_1674,N_2443);
nand U3101 (N_3101,N_2260,N_1527);
nor U3102 (N_3102,N_2627,N_2302);
and U3103 (N_3103,N_1995,N_1702);
nor U3104 (N_3104,N_2770,N_2209);
nor U3105 (N_3105,N_2439,N_2350);
xor U3106 (N_3106,N_1788,N_2555);
nor U3107 (N_3107,N_2565,N_2199);
xor U3108 (N_3108,N_2298,N_2013);
nor U3109 (N_3109,N_2277,N_2016);
and U3110 (N_3110,N_2868,N_1693);
or U3111 (N_3111,N_1714,N_2035);
or U3112 (N_3112,N_1639,N_2437);
xor U3113 (N_3113,N_1671,N_2156);
or U3114 (N_3114,N_1724,N_2540);
and U3115 (N_3115,N_2644,N_2099);
or U3116 (N_3116,N_2190,N_1917);
nand U3117 (N_3117,N_2187,N_2829);
or U3118 (N_3118,N_1515,N_1787);
nand U3119 (N_3119,N_1523,N_2754);
or U3120 (N_3120,N_1937,N_1875);
nand U3121 (N_3121,N_2955,N_1762);
xor U3122 (N_3122,N_1753,N_2571);
or U3123 (N_3123,N_2270,N_2516);
nor U3124 (N_3124,N_2970,N_2212);
and U3125 (N_3125,N_1577,N_2663);
xnor U3126 (N_3126,N_1720,N_2752);
nor U3127 (N_3127,N_2634,N_2832);
nor U3128 (N_3128,N_2917,N_1836);
xor U3129 (N_3129,N_2859,N_2325);
nor U3130 (N_3130,N_2133,N_2356);
or U3131 (N_3131,N_2490,N_1614);
nand U3132 (N_3132,N_2833,N_1595);
and U3133 (N_3133,N_1993,N_1554);
or U3134 (N_3134,N_2674,N_2874);
xor U3135 (N_3135,N_1956,N_1749);
nand U3136 (N_3136,N_1842,N_1968);
nor U3137 (N_3137,N_2944,N_2282);
or U3138 (N_3138,N_2835,N_2498);
and U3139 (N_3139,N_1758,N_2086);
or U3140 (N_3140,N_1684,N_1815);
xor U3141 (N_3141,N_2739,N_2009);
xor U3142 (N_3142,N_2171,N_2991);
and U3143 (N_3143,N_1695,N_1545);
xnor U3144 (N_3144,N_1740,N_2196);
xor U3145 (N_3145,N_2537,N_1800);
and U3146 (N_3146,N_2758,N_2673);
and U3147 (N_3147,N_1518,N_1980);
xor U3148 (N_3148,N_2650,N_2852);
nor U3149 (N_3149,N_2463,N_2239);
nor U3150 (N_3150,N_1551,N_2400);
or U3151 (N_3151,N_2632,N_2104);
nand U3152 (N_3152,N_2034,N_2492);
xnor U3153 (N_3153,N_1801,N_2896);
and U3154 (N_3154,N_2154,N_1552);
nand U3155 (N_3155,N_2264,N_2953);
or U3156 (N_3156,N_1969,N_1859);
and U3157 (N_3157,N_1739,N_1612);
nand U3158 (N_3158,N_2485,N_2025);
nor U3159 (N_3159,N_2225,N_1964);
xnor U3160 (N_3160,N_2291,N_2435);
or U3161 (N_3161,N_1532,N_2618);
nor U3162 (N_3162,N_2888,N_2732);
or U3163 (N_3163,N_1764,N_2320);
or U3164 (N_3164,N_2783,N_1885);
or U3165 (N_3165,N_2989,N_2406);
and U3166 (N_3166,N_1867,N_2266);
nor U3167 (N_3167,N_2367,N_2715);
nor U3168 (N_3168,N_2726,N_2520);
and U3169 (N_3169,N_1543,N_1843);
nor U3170 (N_3170,N_2097,N_2708);
nand U3171 (N_3171,N_2737,N_1776);
xor U3172 (N_3172,N_2809,N_1987);
xor U3173 (N_3173,N_2233,N_2465);
nor U3174 (N_3174,N_2622,N_2421);
nor U3175 (N_3175,N_2626,N_2357);
nor U3176 (N_3176,N_1521,N_1811);
nand U3177 (N_3177,N_2444,N_1555);
and U3178 (N_3178,N_1665,N_2607);
and U3179 (N_3179,N_2112,N_2949);
or U3180 (N_3180,N_2651,N_2172);
nor U3181 (N_3181,N_1745,N_2788);
and U3182 (N_3182,N_2870,N_1611);
and U3183 (N_3183,N_1810,N_1565);
xor U3184 (N_3184,N_1818,N_2211);
nand U3185 (N_3185,N_2919,N_2864);
and U3186 (N_3186,N_2667,N_2200);
xor U3187 (N_3187,N_2751,N_2554);
nand U3188 (N_3188,N_2182,N_2075);
xor U3189 (N_3189,N_1856,N_1741);
nor U3190 (N_3190,N_2566,N_2598);
nor U3191 (N_3191,N_1970,N_2012);
nor U3192 (N_3192,N_2499,N_1935);
or U3193 (N_3193,N_1561,N_1519);
xnor U3194 (N_3194,N_1744,N_2256);
or U3195 (N_3195,N_1690,N_1905);
nor U3196 (N_3196,N_1930,N_2162);
or U3197 (N_3197,N_2779,N_1904);
nor U3198 (N_3198,N_2747,N_2765);
nand U3199 (N_3199,N_1965,N_2801);
nor U3200 (N_3200,N_2436,N_1507);
and U3201 (N_3201,N_2126,N_2594);
nor U3202 (N_3202,N_2787,N_1650);
and U3203 (N_3203,N_2414,N_2338);
or U3204 (N_3204,N_1932,N_2766);
xnor U3205 (N_3205,N_2060,N_2297);
nor U3206 (N_3206,N_2313,N_2477);
or U3207 (N_3207,N_2531,N_2799);
nand U3208 (N_3208,N_2983,N_1570);
xor U3209 (N_3209,N_1854,N_2534);
nor U3210 (N_3210,N_1777,N_2231);
and U3211 (N_3211,N_2973,N_2735);
nand U3212 (N_3212,N_2636,N_2547);
or U3213 (N_3213,N_1560,N_2932);
nor U3214 (N_3214,N_1933,N_1847);
xnor U3215 (N_3215,N_1615,N_2149);
and U3216 (N_3216,N_2031,N_2037);
xnor U3217 (N_3217,N_1558,N_1689);
and U3218 (N_3218,N_1718,N_2964);
xor U3219 (N_3219,N_2135,N_2994);
and U3220 (N_3220,N_1869,N_2524);
nand U3221 (N_3221,N_2071,N_2420);
nand U3222 (N_3222,N_2226,N_2480);
or U3223 (N_3223,N_2213,N_1947);
nand U3224 (N_3224,N_2412,N_2755);
or U3225 (N_3225,N_1783,N_2900);
and U3226 (N_3226,N_2502,N_2967);
xor U3227 (N_3227,N_2811,N_2413);
and U3228 (N_3228,N_2158,N_1814);
xor U3229 (N_3229,N_2354,N_1568);
nor U3230 (N_3230,N_1756,N_1999);
and U3231 (N_3231,N_2263,N_2139);
nor U3232 (N_3232,N_1649,N_2335);
nor U3233 (N_3233,N_2665,N_2363);
and U3234 (N_3234,N_2794,N_1799);
or U3235 (N_3235,N_1696,N_2608);
xor U3236 (N_3236,N_1926,N_2823);
or U3237 (N_3237,N_2819,N_2262);
nand U3238 (N_3238,N_1967,N_2865);
nand U3239 (N_3239,N_2180,N_2638);
and U3240 (N_3240,N_1877,N_2813);
xnor U3241 (N_3241,N_2336,N_2445);
nor U3242 (N_3242,N_1709,N_2527);
and U3243 (N_3243,N_2381,N_2629);
nand U3244 (N_3244,N_1906,N_2895);
and U3245 (N_3245,N_1517,N_2822);
nand U3246 (N_3246,N_2203,N_2976);
or U3247 (N_3247,N_1858,N_2908);
nand U3248 (N_3248,N_1747,N_2616);
and U3249 (N_3249,N_2664,N_2789);
or U3250 (N_3250,N_1795,N_1755);
nor U3251 (N_3251,N_2221,N_2961);
or U3252 (N_3252,N_1841,N_2543);
or U3253 (N_3253,N_2348,N_2577);
and U3254 (N_3254,N_2021,N_2355);
nand U3255 (N_3255,N_2408,N_2072);
nor U3256 (N_3256,N_1572,N_2219);
xnor U3257 (N_3257,N_1637,N_2619);
xor U3258 (N_3258,N_1587,N_1529);
nor U3259 (N_3259,N_1729,N_2064);
or U3260 (N_3260,N_2269,N_2625);
and U3261 (N_3261,N_1525,N_2573);
or U3262 (N_3262,N_2430,N_1608);
or U3263 (N_3263,N_2164,N_1804);
nor U3264 (N_3264,N_2710,N_2504);
nor U3265 (N_3265,N_1790,N_2344);
or U3266 (N_3266,N_2810,N_1653);
nor U3267 (N_3267,N_2223,N_2059);
nor U3268 (N_3268,N_2304,N_2505);
or U3269 (N_3269,N_2965,N_2772);
nand U3270 (N_3270,N_1668,N_2753);
nor U3271 (N_3271,N_2087,N_1946);
and U3272 (N_3272,N_1710,N_1550);
nor U3273 (N_3273,N_1868,N_2340);
nand U3274 (N_3274,N_2395,N_2063);
nor U3275 (N_3275,N_1844,N_1547);
xnor U3276 (N_3276,N_1686,N_2169);
nand U3277 (N_3277,N_2750,N_2678);
nor U3278 (N_3278,N_2377,N_2292);
and U3279 (N_3279,N_1908,N_1501);
nand U3280 (N_3280,N_2995,N_2288);
and U3281 (N_3281,N_2425,N_2889);
nand U3282 (N_3282,N_2165,N_2725);
or U3283 (N_3283,N_1786,N_2930);
or U3284 (N_3284,N_1642,N_2364);
and U3285 (N_3285,N_1920,N_1925);
nand U3286 (N_3286,N_2918,N_2497);
xor U3287 (N_3287,N_2092,N_2144);
xnor U3288 (N_3288,N_2718,N_2960);
nand U3289 (N_3289,N_2939,N_2906);
and U3290 (N_3290,N_2817,N_1592);
nor U3291 (N_3291,N_1600,N_2471);
nand U3292 (N_3292,N_2130,N_1807);
xor U3293 (N_3293,N_2748,N_1902);
and U3294 (N_3294,N_2538,N_2319);
nor U3295 (N_3295,N_2140,N_2898);
nand U3296 (N_3296,N_2605,N_2259);
xnor U3297 (N_3297,N_2036,N_1603);
nand U3298 (N_3298,N_2959,N_1526);
and U3299 (N_3299,N_1598,N_2713);
nor U3300 (N_3300,N_2379,N_2880);
and U3301 (N_3301,N_2517,N_2511);
or U3302 (N_3302,N_2560,N_2467);
or U3303 (N_3303,N_1825,N_2373);
and U3304 (N_3304,N_1707,N_2342);
nor U3305 (N_3305,N_1934,N_2241);
xor U3306 (N_3306,N_2456,N_1606);
and U3307 (N_3307,N_1751,N_1656);
nor U3308 (N_3308,N_2409,N_1816);
xor U3309 (N_3309,N_2523,N_2096);
nor U3310 (N_3310,N_2387,N_2376);
nor U3311 (N_3311,N_2159,N_2278);
and U3312 (N_3312,N_2179,N_1851);
or U3313 (N_3313,N_2558,N_1894);
and U3314 (N_3314,N_2828,N_2238);
and U3315 (N_3315,N_2941,N_2806);
or U3316 (N_3316,N_2701,N_1646);
xor U3317 (N_3317,N_2838,N_2777);
xor U3318 (N_3318,N_1556,N_1974);
nand U3319 (N_3319,N_2872,N_1782);
nor U3320 (N_3320,N_2774,N_2386);
or U3321 (N_3321,N_2685,N_2840);
or U3322 (N_3322,N_2615,N_2839);
nor U3323 (N_3323,N_1681,N_1878);
and U3324 (N_3324,N_2660,N_1803);
and U3325 (N_3325,N_2952,N_1848);
xor U3326 (N_3326,N_1645,N_1676);
xor U3327 (N_3327,N_2677,N_2198);
and U3328 (N_3328,N_2118,N_2202);
or U3329 (N_3329,N_1578,N_1509);
xor U3330 (N_3330,N_2496,N_1888);
xnor U3331 (N_3331,N_2843,N_2943);
or U3332 (N_3332,N_2617,N_2067);
nand U3333 (N_3333,N_2921,N_2329);
nor U3334 (N_3334,N_2837,N_2275);
and U3335 (N_3335,N_2762,N_2834);
nor U3336 (N_3336,N_2295,N_2521);
nand U3337 (N_3337,N_2653,N_2576);
or U3338 (N_3338,N_2591,N_1838);
or U3339 (N_3339,N_2704,N_1632);
and U3340 (N_3340,N_2988,N_2700);
and U3341 (N_3341,N_2460,N_2041);
nor U3342 (N_3342,N_2620,N_2633);
nand U3343 (N_3343,N_2652,N_1712);
or U3344 (N_3344,N_1711,N_2215);
nand U3345 (N_3345,N_1837,N_2388);
and U3346 (N_3346,N_2257,N_1721);
nor U3347 (N_3347,N_1876,N_1573);
nand U3348 (N_3348,N_1655,N_2242);
xnor U3349 (N_3349,N_2546,N_2125);
or U3350 (N_3350,N_1798,N_2384);
or U3351 (N_3351,N_2711,N_2857);
or U3352 (N_3352,N_2014,N_2984);
and U3353 (N_3353,N_1569,N_1857);
or U3354 (N_3354,N_2455,N_2109);
nor U3355 (N_3355,N_2730,N_1871);
and U3356 (N_3356,N_1778,N_2150);
and U3357 (N_3357,N_1728,N_2450);
and U3358 (N_3358,N_1641,N_2604);
nand U3359 (N_3359,N_2956,N_2115);
nand U3360 (N_3360,N_2570,N_2600);
nor U3361 (N_3361,N_2472,N_2797);
nand U3362 (N_3362,N_1644,N_2938);
nor U3363 (N_3363,N_2175,N_2382);
nor U3364 (N_3364,N_2643,N_2081);
nor U3365 (N_3365,N_2138,N_2120);
nor U3366 (N_3366,N_1940,N_2286);
nand U3367 (N_3367,N_2545,N_2353);
nand U3368 (N_3368,N_2074,N_2935);
xnor U3369 (N_3369,N_1839,N_2575);
nand U3370 (N_3370,N_2433,N_2365);
nor U3371 (N_3371,N_1981,N_1638);
nand U3372 (N_3372,N_2866,N_2999);
or U3373 (N_3373,N_2503,N_2080);
nand U3374 (N_3374,N_2579,N_2068);
or U3375 (N_3375,N_2587,N_1900);
xnor U3376 (N_3376,N_2103,N_1604);
and U3377 (N_3377,N_2056,N_2296);
nor U3378 (N_3378,N_1502,N_2333);
xor U3379 (N_3379,N_2258,N_2197);
or U3380 (N_3380,N_2585,N_2815);
or U3381 (N_3381,N_2552,N_2177);
nand U3382 (N_3382,N_2533,N_2488);
xnor U3383 (N_3383,N_1624,N_1657);
nand U3384 (N_3384,N_1919,N_2785);
nand U3385 (N_3385,N_2987,N_2916);
or U3386 (N_3386,N_2186,N_2393);
or U3387 (N_3387,N_2500,N_2155);
nor U3388 (N_3388,N_2440,N_2648);
nor U3389 (N_3389,N_2131,N_1531);
nor U3390 (N_3390,N_1594,N_1752);
and U3391 (N_3391,N_2327,N_2911);
xnor U3392 (N_3392,N_2090,N_2026);
nor U3393 (N_3393,N_1830,N_1991);
and U3394 (N_3394,N_1860,N_2345);
nand U3395 (N_3395,N_1673,N_1662);
nor U3396 (N_3396,N_2459,N_2512);
nand U3397 (N_3397,N_2404,N_2403);
nand U3398 (N_3398,N_2105,N_2375);
xor U3399 (N_3399,N_2113,N_1997);
or U3400 (N_3400,N_1738,N_1960);
and U3401 (N_3401,N_2907,N_1760);
nor U3402 (N_3402,N_1564,N_2997);
or U3403 (N_3403,N_1667,N_1955);
xor U3404 (N_3404,N_1679,N_2800);
and U3405 (N_3405,N_1510,N_2422);
or U3406 (N_3406,N_1627,N_1546);
nand U3407 (N_3407,N_2613,N_1622);
and U3408 (N_3408,N_2079,N_2167);
xor U3409 (N_3409,N_2360,N_1821);
nand U3410 (N_3410,N_2776,N_2228);
xnor U3411 (N_3411,N_2798,N_2693);
nand U3412 (N_3412,N_2926,N_2240);
and U3413 (N_3413,N_2134,N_2337);
nand U3414 (N_3414,N_1620,N_2028);
xor U3415 (N_3415,N_2267,N_2826);
and U3416 (N_3416,N_2990,N_2448);
nor U3417 (N_3417,N_2438,N_2121);
or U3418 (N_3418,N_2791,N_2058);
xnor U3419 (N_3419,N_2586,N_2315);
xnor U3420 (N_3420,N_2243,N_2532);
xnor U3421 (N_3421,N_2235,N_1596);
nor U3422 (N_3422,N_1978,N_2424);
nand U3423 (N_3423,N_1648,N_2602);
and U3424 (N_3424,N_1661,N_1535);
xor U3425 (N_3425,N_1534,N_1730);
xnor U3426 (N_3426,N_1773,N_2108);
xor U3427 (N_3427,N_1971,N_2441);
xnor U3428 (N_3428,N_2903,N_2284);
nand U3429 (N_3429,N_2614,N_1808);
and U3430 (N_3430,N_2716,N_2740);
xnor U3431 (N_3431,N_2588,N_2854);
nand U3432 (N_3432,N_2893,N_2078);
nor U3433 (N_3433,N_2736,N_2142);
and U3434 (N_3434,N_2544,N_2847);
or U3435 (N_3435,N_2680,N_1941);
and U3436 (N_3436,N_2214,N_2110);
nand U3437 (N_3437,N_2671,N_1701);
xor U3438 (N_3438,N_2347,N_1775);
nor U3439 (N_3439,N_2899,N_2525);
or U3440 (N_3440,N_2091,N_1538);
nor U3441 (N_3441,N_1715,N_2549);
nand U3442 (N_3442,N_2937,N_2328);
nand U3443 (N_3443,N_2929,N_2820);
and U3444 (N_3444,N_2145,N_2574);
xor U3445 (N_3445,N_2098,N_1522);
nor U3446 (N_3446,N_2369,N_2920);
nor U3447 (N_3447,N_1881,N_2580);
or U3448 (N_3448,N_1660,N_2019);
nand U3449 (N_3449,N_2299,N_1793);
nor U3450 (N_3450,N_2095,N_2993);
xnor U3451 (N_3451,N_2936,N_2311);
xnor U3452 (N_3452,N_2756,N_2317);
nand U3453 (N_3453,N_1789,N_2786);
and U3454 (N_3454,N_2969,N_2236);
xor U3455 (N_3455,N_2023,N_2310);
xor U3456 (N_3456,N_2818,N_1759);
nor U3457 (N_3457,N_2862,N_2687);
and U3458 (N_3458,N_2656,N_2621);
xor U3459 (N_3459,N_2473,N_2804);
nand U3460 (N_3460,N_1880,N_1723);
or U3461 (N_3461,N_2216,N_2249);
xnor U3462 (N_3462,N_1996,N_2008);
xor U3463 (N_3463,N_2407,N_1705);
and U3464 (N_3464,N_2123,N_2206);
and U3465 (N_3465,N_2402,N_1779);
nor U3466 (N_3466,N_2449,N_2274);
or U3467 (N_3467,N_2482,N_1672);
or U3468 (N_3468,N_2842,N_2446);
or U3469 (N_3469,N_1562,N_2289);
nand U3470 (N_3470,N_1548,N_2230);
nor U3471 (N_3471,N_2006,N_2780);
xnor U3472 (N_3472,N_2882,N_2318);
and U3473 (N_3473,N_1768,N_2510);
and U3474 (N_3474,N_1982,N_1634);
or U3475 (N_3475,N_2201,N_2814);
or U3476 (N_3476,N_2530,N_2528);
nor U3477 (N_3477,N_1540,N_1898);
nand U3478 (N_3478,N_2979,N_2812);
nor U3479 (N_3479,N_2703,N_2901);
nand U3480 (N_3480,N_1582,N_1722);
and U3481 (N_3481,N_2392,N_1733);
nand U3482 (N_3482,N_2191,N_2334);
xnor U3483 (N_3483,N_1785,N_2645);
and U3484 (N_3484,N_2821,N_2724);
nand U3485 (N_3485,N_1819,N_2698);
nor U3486 (N_3486,N_2514,N_2501);
nand U3487 (N_3487,N_2890,N_1617);
nor U3488 (N_3488,N_2824,N_2998);
or U3489 (N_3489,N_2038,N_1659);
nor U3490 (N_3490,N_2669,N_2452);
or U3491 (N_3491,N_2782,N_2027);
xor U3492 (N_3492,N_2351,N_1623);
or U3493 (N_3493,N_2017,N_2401);
nand U3494 (N_3494,N_2323,N_2879);
nand U3495 (N_3495,N_1520,N_2052);
or U3496 (N_3496,N_2137,N_2361);
nand U3497 (N_3497,N_2719,N_1508);
xnor U3498 (N_3498,N_1663,N_1791);
xor U3499 (N_3499,N_2946,N_1652);
or U3500 (N_3500,N_2119,N_2707);
nand U3501 (N_3501,N_2850,N_1953);
xnor U3502 (N_3502,N_1746,N_1583);
nand U3503 (N_3503,N_2925,N_2909);
xnor U3504 (N_3504,N_2564,N_1505);
nand U3505 (N_3505,N_1736,N_1706);
and U3506 (N_3506,N_2722,N_1883);
or U3507 (N_3507,N_1719,N_1928);
nor U3508 (N_3508,N_2744,N_2635);
and U3509 (N_3509,N_2661,N_2583);
xor U3510 (N_3510,N_2996,N_1958);
nand U3511 (N_3511,N_1750,N_2696);
or U3512 (N_3512,N_2247,N_2695);
xnor U3513 (N_3513,N_2085,N_2541);
nor U3514 (N_3514,N_1621,N_2004);
or U3515 (N_3515,N_1500,N_2792);
or U3516 (N_3516,N_2881,N_2043);
nor U3517 (N_3517,N_1792,N_2088);
or U3518 (N_3518,N_2581,N_1945);
xnor U3519 (N_3519,N_2124,N_2308);
nand U3520 (N_3520,N_2631,N_1774);
nand U3521 (N_3521,N_1699,N_2487);
or U3522 (N_3522,N_2831,N_1607);
xor U3523 (N_3523,N_1929,N_1593);
xor U3524 (N_3524,N_2234,N_2305);
nand U3525 (N_3525,N_2475,N_1584);
nor U3526 (N_3526,N_1865,N_1781);
xor U3527 (N_3527,N_2928,N_1962);
nand U3528 (N_3528,N_2083,N_2738);
nand U3529 (N_3529,N_1683,N_2846);
nor U3530 (N_3530,N_2706,N_2237);
nand U3531 (N_3531,N_1537,N_2848);
nor U3532 (N_3532,N_1687,N_2720);
xor U3533 (N_3533,N_2905,N_1651);
nor U3534 (N_3534,N_2065,N_1957);
nor U3535 (N_3535,N_2519,N_2077);
and U3536 (N_3536,N_2757,N_2883);
nand U3537 (N_3537,N_1895,N_2188);
or U3538 (N_3538,N_2391,N_1767);
or U3539 (N_3539,N_2332,N_2227);
nand U3540 (N_3540,N_2285,N_1688);
nor U3541 (N_3541,N_2279,N_1809);
and U3542 (N_3542,N_2977,N_2869);
xor U3543 (N_3543,N_2860,N_2464);
nor U3544 (N_3544,N_1966,N_1516);
or U3545 (N_3545,N_2972,N_1985);
nand U3546 (N_3546,N_2934,N_2293);
and U3547 (N_3547,N_2599,N_1588);
nand U3548 (N_3548,N_2924,N_1984);
and U3549 (N_3549,N_1824,N_2431);
or U3550 (N_3550,N_2229,N_1635);
and U3551 (N_3551,N_2468,N_2526);
xnor U3552 (N_3552,N_2733,N_1797);
nand U3553 (N_3553,N_1892,N_2457);
nand U3554 (N_3554,N_2553,N_2884);
nor U3555 (N_3555,N_1931,N_2927);
or U3556 (N_3556,N_2102,N_2584);
xnor U3557 (N_3557,N_2010,N_2163);
nor U3558 (N_3558,N_2951,N_2670);
xor U3559 (N_3559,N_2273,N_2429);
nand U3560 (N_3560,N_1682,N_1990);
or U3561 (N_3561,N_2688,N_2136);
or U3562 (N_3562,N_1566,N_1685);
xnor U3563 (N_3563,N_2300,N_1716);
or U3564 (N_3564,N_2690,N_2061);
or U3565 (N_3565,N_2394,N_2931);
xnor U3566 (N_3566,N_2152,N_2020);
and U3567 (N_3567,N_1666,N_2389);
xor U3568 (N_3568,N_2561,N_2195);
nand U3569 (N_3569,N_2222,N_1654);
and U3570 (N_3570,N_2649,N_1972);
xor U3571 (N_3571,N_1731,N_1915);
or U3572 (N_3572,N_2589,N_2324);
nor U3573 (N_3573,N_1658,N_1942);
xnor U3574 (N_3574,N_2749,N_2129);
or U3575 (N_3575,N_2897,N_2265);
nand U3576 (N_3576,N_2117,N_2434);
or U3577 (N_3577,N_2094,N_1886);
xnor U3578 (N_3578,N_2506,N_2557);
nand U3579 (N_3579,N_1539,N_2128);
or U3580 (N_3580,N_2451,N_2371);
or U3581 (N_3581,N_1889,N_1973);
nor U3582 (N_3582,N_1828,N_2003);
nand U3583 (N_3583,N_2729,N_2411);
and U3584 (N_3584,N_2734,N_1918);
nor U3585 (N_3585,N_2268,N_2374);
xnor U3586 (N_3586,N_1647,N_2971);
or U3587 (N_3587,N_2796,N_2845);
nand U3588 (N_3588,N_2950,N_2220);
or U3589 (N_3589,N_1528,N_2244);
nor U3590 (N_3590,N_2415,N_2873);
nor U3591 (N_3591,N_2383,N_2251);
nor U3592 (N_3592,N_2876,N_2657);
nand U3593 (N_3593,N_2307,N_1630);
nor U3594 (N_3594,N_2322,N_2466);
or U3595 (N_3595,N_2947,N_2474);
xor U3596 (N_3596,N_1948,N_1742);
and U3597 (N_3597,N_2461,N_1988);
nand U3598 (N_3598,N_1533,N_2863);
nor U3599 (N_3599,N_2217,N_2316);
and U3600 (N_3600,N_2122,N_2029);
and U3601 (N_3601,N_1855,N_2692);
xor U3602 (N_3602,N_2910,N_2923);
nand U3603 (N_3603,N_2912,N_2781);
or U3604 (N_3604,N_1903,N_1542);
nor U3605 (N_3605,N_2769,N_1669);
nor U3606 (N_3606,N_2271,N_2805);
nor U3607 (N_3607,N_1989,N_1845);
nand U3608 (N_3608,N_2050,N_2624);
nand U3609 (N_3609,N_1938,N_2309);
nor U3610 (N_3610,N_2419,N_1503);
nor U3611 (N_3611,N_1794,N_2280);
or U3612 (N_3612,N_2853,N_2778);
nand U3613 (N_3613,N_1864,N_2962);
nand U3614 (N_3614,N_1913,N_2945);
xnor U3615 (N_3615,N_2321,N_2795);
nor U3616 (N_3616,N_1576,N_2042);
xor U3617 (N_3617,N_2000,N_2495);
nand U3618 (N_3618,N_2287,N_2572);
nor U3619 (N_3619,N_2447,N_2148);
xnor U3620 (N_3620,N_2699,N_1504);
or U3621 (N_3621,N_2858,N_2168);
nor U3622 (N_3622,N_1912,N_1579);
xnor U3623 (N_3623,N_2764,N_2658);
nor U3624 (N_3624,N_2682,N_1590);
nor U3625 (N_3625,N_2827,N_2276);
nor U3626 (N_3626,N_1846,N_2731);
nand U3627 (N_3627,N_1691,N_2101);
xor U3628 (N_3628,N_1694,N_2250);
nand U3629 (N_3629,N_2830,N_2205);
nand U3630 (N_3630,N_2469,N_1770);
or U3631 (N_3631,N_2157,N_1911);
xnor U3632 (N_3632,N_2803,N_1849);
nand U3633 (N_3633,N_2871,N_2891);
nand U3634 (N_3634,N_1725,N_1812);
xor U3635 (N_3635,N_1757,N_2066);
or U3636 (N_3636,N_1727,N_1923);
xnor U3637 (N_3637,N_2948,N_2033);
and U3638 (N_3638,N_1829,N_2851);
nand U3639 (N_3639,N_1784,N_2189);
and U3640 (N_3640,N_2248,N_2370);
nor U3641 (N_3641,N_1852,N_2784);
xnor U3642 (N_3642,N_1914,N_2082);
nand U3643 (N_3643,N_2717,N_2294);
xnor U3644 (N_3644,N_1771,N_2647);
and U3645 (N_3645,N_1959,N_2728);
nor U3646 (N_3646,N_2654,N_1921);
nor U3647 (N_3647,N_1796,N_2326);
or U3648 (N_3648,N_2723,N_1765);
nand U3649 (N_3649,N_2559,N_2398);
and U3650 (N_3650,N_2417,N_1832);
and U3651 (N_3651,N_2721,N_2705);
nand U3652 (N_3652,N_2339,N_2385);
xnor U3653 (N_3653,N_1625,N_2143);
and U3654 (N_3654,N_2048,N_2032);
and U3655 (N_3655,N_1874,N_2184);
or U3656 (N_3656,N_1954,N_2116);
xor U3657 (N_3657,N_2290,N_2301);
nand U3658 (N_3658,N_2746,N_2610);
or U3659 (N_3659,N_1530,N_1826);
and U3660 (N_3660,N_2975,N_2518);
xnor U3661 (N_3661,N_2343,N_2153);
nand U3662 (N_3662,N_2915,N_1643);
xor U3663 (N_3663,N_2359,N_2902);
xnor U3664 (N_3664,N_1631,N_2681);
or U3665 (N_3665,N_2773,N_2974);
nand U3666 (N_3666,N_2245,N_1589);
nand U3667 (N_3667,N_1992,N_2272);
nand U3668 (N_3668,N_1862,N_1950);
nor U3669 (N_3669,N_1884,N_1924);
and U3670 (N_3670,N_2592,N_1863);
or U3671 (N_3671,N_1697,N_1678);
xor U3672 (N_3672,N_2790,N_2084);
or U3673 (N_3673,N_2942,N_2442);
or U3674 (N_3674,N_1977,N_2712);
or U3675 (N_3675,N_1628,N_2432);
or U3676 (N_3676,N_2596,N_2341);
xnor U3677 (N_3677,N_2954,N_1748);
xnor U3678 (N_3678,N_2914,N_2507);
nor U3679 (N_3679,N_2055,N_2418);
nor U3680 (N_3680,N_1585,N_1817);
nor U3681 (N_3681,N_1853,N_2178);
xor U3682 (N_3682,N_2886,N_2841);
and U3683 (N_3683,N_1986,N_2639);
nor U3684 (N_3684,N_2346,N_2281);
nor U3685 (N_3685,N_2397,N_1806);
and U3686 (N_3686,N_1704,N_1901);
or U3687 (N_3687,N_1553,N_2076);
nand U3688 (N_3688,N_2875,N_2210);
and U3689 (N_3689,N_2981,N_2053);
or U3690 (N_3690,N_2563,N_2940);
and U3691 (N_3691,N_2885,N_1559);
nand U3692 (N_3692,N_1581,N_2982);
xnor U3693 (N_3693,N_1734,N_2675);
nand U3694 (N_3694,N_1513,N_1979);
nor U3695 (N_3695,N_2877,N_2568);
nor U3696 (N_3696,N_2913,N_2641);
and U3697 (N_3697,N_2246,N_2878);
nor U3698 (N_3698,N_1677,N_2894);
nand U3699 (N_3699,N_1618,N_1891);
and U3700 (N_3700,N_2642,N_2536);
or U3701 (N_3701,N_2358,N_2759);
or U3702 (N_3702,N_2985,N_2768);
nand U3703 (N_3703,N_2689,N_2107);
or U3704 (N_3704,N_1963,N_1922);
xor U3705 (N_3705,N_1813,N_2771);
and U3706 (N_3706,N_2590,N_2024);
nor U3707 (N_3707,N_1850,N_2453);
or U3708 (N_3708,N_2111,N_2491);
nor U3709 (N_3709,N_2314,N_2054);
xnor U3710 (N_3710,N_2486,N_1626);
or U3711 (N_3711,N_1708,N_2127);
and U3712 (N_3712,N_2825,N_2676);
xnor U3713 (N_3713,N_1591,N_1916);
or U3714 (N_3714,N_2662,N_2968);
or U3715 (N_3715,N_2922,N_2283);
nand U3716 (N_3716,N_1726,N_2378);
nand U3717 (N_3717,N_1769,N_2630);
nor U3718 (N_3718,N_2493,N_2100);
or U3719 (N_3719,N_2390,N_2047);
and U3720 (N_3720,N_2760,N_1840);
nand U3721 (N_3721,N_2147,N_1872);
and U3722 (N_3722,N_2694,N_1833);
and U3723 (N_3723,N_1873,N_2405);
and U3724 (N_3724,N_2761,N_1861);
xnor U3725 (N_3725,N_2745,N_2479);
and U3726 (N_3726,N_2904,N_1907);
nor U3727 (N_3727,N_2366,N_2224);
or U3728 (N_3728,N_2763,N_2861);
nand U3729 (N_3729,N_2470,N_2637);
or U3730 (N_3730,N_2049,N_2174);
nand U3731 (N_3731,N_1927,N_2529);
nand U3732 (N_3732,N_2992,N_2672);
and U3733 (N_3733,N_2508,N_2686);
or U3734 (N_3734,N_2022,N_2582);
and U3735 (N_3735,N_2986,N_2593);
and U3736 (N_3736,N_2410,N_1633);
nand U3737 (N_3737,N_1943,N_2556);
and U3738 (N_3738,N_2542,N_1994);
or U3739 (N_3739,N_2684,N_2668);
nor U3740 (N_3740,N_2303,N_1680);
or U3741 (N_3741,N_2057,N_1636);
and U3742 (N_3742,N_2349,N_2183);
and U3743 (N_3743,N_2312,N_1512);
or U3744 (N_3744,N_2597,N_1599);
and U3745 (N_3745,N_1780,N_1619);
and U3746 (N_3746,N_2958,N_2207);
nor U3747 (N_3747,N_1743,N_2253);
and U3748 (N_3748,N_1557,N_2254);
nand U3749 (N_3749,N_2683,N_1822);
nand U3750 (N_3750,N_1861,N_2011);
nand U3751 (N_3751,N_2059,N_2742);
and U3752 (N_3752,N_2693,N_2773);
nor U3753 (N_3753,N_1859,N_2614);
and U3754 (N_3754,N_2445,N_1687);
or U3755 (N_3755,N_1783,N_2670);
nand U3756 (N_3756,N_2060,N_2274);
xor U3757 (N_3757,N_1626,N_2101);
xnor U3758 (N_3758,N_2658,N_2464);
nor U3759 (N_3759,N_1666,N_1804);
nor U3760 (N_3760,N_2707,N_2296);
and U3761 (N_3761,N_2267,N_2325);
and U3762 (N_3762,N_1574,N_2031);
or U3763 (N_3763,N_1728,N_2713);
nor U3764 (N_3764,N_1659,N_2231);
xnor U3765 (N_3765,N_2779,N_2732);
or U3766 (N_3766,N_2394,N_2099);
or U3767 (N_3767,N_2476,N_2749);
xor U3768 (N_3768,N_1730,N_2109);
and U3769 (N_3769,N_2963,N_2947);
xor U3770 (N_3770,N_1906,N_1763);
xnor U3771 (N_3771,N_2173,N_1646);
or U3772 (N_3772,N_1550,N_2475);
and U3773 (N_3773,N_2936,N_2731);
and U3774 (N_3774,N_1616,N_2868);
nor U3775 (N_3775,N_2340,N_2074);
and U3776 (N_3776,N_2197,N_1941);
xnor U3777 (N_3777,N_1502,N_2092);
or U3778 (N_3778,N_1615,N_2262);
xnor U3779 (N_3779,N_2457,N_2330);
nand U3780 (N_3780,N_1812,N_1574);
nand U3781 (N_3781,N_2806,N_2132);
nor U3782 (N_3782,N_2376,N_2656);
nor U3783 (N_3783,N_2464,N_2123);
or U3784 (N_3784,N_2221,N_2443);
nor U3785 (N_3785,N_2328,N_1559);
and U3786 (N_3786,N_2296,N_2151);
or U3787 (N_3787,N_2566,N_2135);
xor U3788 (N_3788,N_2106,N_1533);
xnor U3789 (N_3789,N_1686,N_1653);
nand U3790 (N_3790,N_2162,N_2288);
nand U3791 (N_3791,N_2677,N_2227);
nand U3792 (N_3792,N_2419,N_1759);
xnor U3793 (N_3793,N_1852,N_1918);
nand U3794 (N_3794,N_1615,N_2601);
and U3795 (N_3795,N_2449,N_2559);
xnor U3796 (N_3796,N_1526,N_2154);
xnor U3797 (N_3797,N_2917,N_2689);
nand U3798 (N_3798,N_1694,N_2861);
xnor U3799 (N_3799,N_2389,N_2931);
nand U3800 (N_3800,N_2967,N_2076);
or U3801 (N_3801,N_2152,N_1510);
nand U3802 (N_3802,N_2075,N_1966);
or U3803 (N_3803,N_2880,N_2674);
and U3804 (N_3804,N_1707,N_1734);
or U3805 (N_3805,N_2186,N_2029);
xnor U3806 (N_3806,N_2806,N_2405);
and U3807 (N_3807,N_2382,N_1757);
nand U3808 (N_3808,N_1530,N_1691);
xor U3809 (N_3809,N_2019,N_2058);
and U3810 (N_3810,N_2566,N_2822);
nand U3811 (N_3811,N_2606,N_2309);
or U3812 (N_3812,N_2196,N_2478);
nor U3813 (N_3813,N_2863,N_2611);
nand U3814 (N_3814,N_1532,N_1933);
nor U3815 (N_3815,N_2473,N_2788);
xnor U3816 (N_3816,N_1931,N_1682);
and U3817 (N_3817,N_2794,N_2686);
nand U3818 (N_3818,N_1722,N_2911);
nor U3819 (N_3819,N_1712,N_2455);
xnor U3820 (N_3820,N_2098,N_2760);
nand U3821 (N_3821,N_2060,N_1912);
or U3822 (N_3822,N_2581,N_2987);
xor U3823 (N_3823,N_1925,N_2618);
or U3824 (N_3824,N_2743,N_1806);
and U3825 (N_3825,N_2813,N_2417);
or U3826 (N_3826,N_2089,N_2967);
and U3827 (N_3827,N_2107,N_1780);
or U3828 (N_3828,N_2526,N_2953);
nor U3829 (N_3829,N_1863,N_1665);
nand U3830 (N_3830,N_2005,N_2246);
and U3831 (N_3831,N_1728,N_2233);
or U3832 (N_3832,N_1721,N_2915);
and U3833 (N_3833,N_2214,N_2411);
nor U3834 (N_3834,N_2694,N_2774);
nand U3835 (N_3835,N_2302,N_2529);
and U3836 (N_3836,N_2248,N_1548);
xor U3837 (N_3837,N_2257,N_2158);
xnor U3838 (N_3838,N_1855,N_2581);
or U3839 (N_3839,N_2476,N_1913);
or U3840 (N_3840,N_2977,N_2053);
nand U3841 (N_3841,N_1868,N_2648);
xor U3842 (N_3842,N_2080,N_2987);
nor U3843 (N_3843,N_2861,N_2764);
nand U3844 (N_3844,N_2533,N_1585);
nor U3845 (N_3845,N_1786,N_2414);
and U3846 (N_3846,N_2212,N_2639);
nor U3847 (N_3847,N_1657,N_2612);
xnor U3848 (N_3848,N_1885,N_2809);
and U3849 (N_3849,N_1928,N_2478);
xor U3850 (N_3850,N_2980,N_2303);
nand U3851 (N_3851,N_2503,N_1730);
or U3852 (N_3852,N_2142,N_2826);
nor U3853 (N_3853,N_2162,N_2783);
xor U3854 (N_3854,N_2929,N_1755);
and U3855 (N_3855,N_2009,N_1621);
xor U3856 (N_3856,N_1577,N_2844);
nand U3857 (N_3857,N_1604,N_1636);
or U3858 (N_3858,N_1515,N_2088);
and U3859 (N_3859,N_2678,N_2024);
xnor U3860 (N_3860,N_2406,N_1581);
or U3861 (N_3861,N_2212,N_2819);
and U3862 (N_3862,N_1653,N_2741);
or U3863 (N_3863,N_1574,N_2527);
and U3864 (N_3864,N_1621,N_1676);
nand U3865 (N_3865,N_2077,N_2535);
xor U3866 (N_3866,N_2616,N_2240);
or U3867 (N_3867,N_2116,N_2007);
and U3868 (N_3868,N_2551,N_1743);
xor U3869 (N_3869,N_1515,N_2478);
nor U3870 (N_3870,N_1988,N_1692);
nand U3871 (N_3871,N_2552,N_2876);
xnor U3872 (N_3872,N_1671,N_1825);
xor U3873 (N_3873,N_2832,N_1774);
xnor U3874 (N_3874,N_1639,N_2884);
nor U3875 (N_3875,N_1708,N_2444);
and U3876 (N_3876,N_2448,N_1605);
and U3877 (N_3877,N_1951,N_2291);
and U3878 (N_3878,N_1654,N_1724);
xnor U3879 (N_3879,N_1627,N_2803);
nor U3880 (N_3880,N_1572,N_2942);
nand U3881 (N_3881,N_1867,N_2029);
and U3882 (N_3882,N_2819,N_1659);
nor U3883 (N_3883,N_2810,N_1643);
and U3884 (N_3884,N_1781,N_2085);
and U3885 (N_3885,N_2693,N_1761);
xnor U3886 (N_3886,N_2760,N_2549);
nand U3887 (N_3887,N_1754,N_1750);
and U3888 (N_3888,N_1813,N_2007);
nand U3889 (N_3889,N_2573,N_1521);
or U3890 (N_3890,N_2080,N_1941);
xnor U3891 (N_3891,N_2202,N_2355);
xor U3892 (N_3892,N_2397,N_2878);
nand U3893 (N_3893,N_1612,N_2513);
or U3894 (N_3894,N_2368,N_1967);
nand U3895 (N_3895,N_1580,N_1741);
xnor U3896 (N_3896,N_1995,N_1934);
nor U3897 (N_3897,N_2230,N_1859);
or U3898 (N_3898,N_2058,N_2371);
nand U3899 (N_3899,N_2453,N_1888);
nor U3900 (N_3900,N_2021,N_1862);
nand U3901 (N_3901,N_1558,N_2204);
nor U3902 (N_3902,N_1839,N_1821);
nor U3903 (N_3903,N_2642,N_2057);
nand U3904 (N_3904,N_2273,N_1787);
nand U3905 (N_3905,N_1711,N_2632);
nand U3906 (N_3906,N_1841,N_1898);
nor U3907 (N_3907,N_2652,N_2018);
xor U3908 (N_3908,N_2947,N_2872);
nand U3909 (N_3909,N_2255,N_2676);
and U3910 (N_3910,N_2690,N_2963);
xor U3911 (N_3911,N_2568,N_2483);
and U3912 (N_3912,N_1919,N_2107);
nor U3913 (N_3913,N_2590,N_1522);
nand U3914 (N_3914,N_1629,N_2509);
xor U3915 (N_3915,N_2027,N_2026);
nand U3916 (N_3916,N_2617,N_1758);
and U3917 (N_3917,N_2070,N_2698);
and U3918 (N_3918,N_1578,N_2773);
or U3919 (N_3919,N_2734,N_1961);
nand U3920 (N_3920,N_2574,N_1780);
or U3921 (N_3921,N_1574,N_2241);
xnor U3922 (N_3922,N_1600,N_1909);
or U3923 (N_3923,N_2807,N_2897);
xnor U3924 (N_3924,N_2811,N_1533);
and U3925 (N_3925,N_2188,N_2588);
and U3926 (N_3926,N_2136,N_2127);
xnor U3927 (N_3927,N_2765,N_2226);
or U3928 (N_3928,N_1615,N_1899);
nand U3929 (N_3929,N_2379,N_2807);
and U3930 (N_3930,N_2845,N_1847);
xor U3931 (N_3931,N_1538,N_2623);
and U3932 (N_3932,N_2743,N_1756);
and U3933 (N_3933,N_1569,N_2042);
and U3934 (N_3934,N_2754,N_2117);
nand U3935 (N_3935,N_1501,N_2877);
or U3936 (N_3936,N_2958,N_1825);
and U3937 (N_3937,N_1501,N_1891);
nor U3938 (N_3938,N_2991,N_2870);
nand U3939 (N_3939,N_2365,N_2423);
or U3940 (N_3940,N_2167,N_1823);
nand U3941 (N_3941,N_1917,N_2081);
xor U3942 (N_3942,N_1681,N_2865);
or U3943 (N_3943,N_2171,N_2519);
nor U3944 (N_3944,N_1983,N_1954);
xnor U3945 (N_3945,N_1722,N_2821);
or U3946 (N_3946,N_2802,N_1756);
or U3947 (N_3947,N_2748,N_2286);
nand U3948 (N_3948,N_2916,N_2221);
and U3949 (N_3949,N_1830,N_2814);
nor U3950 (N_3950,N_1885,N_1708);
nand U3951 (N_3951,N_2020,N_2851);
or U3952 (N_3952,N_1949,N_2653);
and U3953 (N_3953,N_2719,N_2458);
or U3954 (N_3954,N_2812,N_1547);
or U3955 (N_3955,N_1532,N_2799);
and U3956 (N_3956,N_2616,N_2182);
or U3957 (N_3957,N_2171,N_2365);
or U3958 (N_3958,N_2470,N_2406);
nand U3959 (N_3959,N_2575,N_2318);
nor U3960 (N_3960,N_2035,N_1532);
or U3961 (N_3961,N_1796,N_2316);
xnor U3962 (N_3962,N_1674,N_2270);
and U3963 (N_3963,N_2143,N_1905);
nand U3964 (N_3964,N_2777,N_1785);
and U3965 (N_3965,N_2674,N_2998);
or U3966 (N_3966,N_2811,N_1540);
and U3967 (N_3967,N_2287,N_2492);
or U3968 (N_3968,N_2090,N_1899);
xnor U3969 (N_3969,N_1772,N_1833);
nand U3970 (N_3970,N_1755,N_1876);
and U3971 (N_3971,N_1981,N_2135);
nor U3972 (N_3972,N_2871,N_2019);
nor U3973 (N_3973,N_1524,N_1906);
nand U3974 (N_3974,N_1616,N_2033);
and U3975 (N_3975,N_1852,N_1818);
xor U3976 (N_3976,N_2910,N_2066);
nand U3977 (N_3977,N_2561,N_2422);
or U3978 (N_3978,N_1655,N_2722);
xor U3979 (N_3979,N_1770,N_1828);
nor U3980 (N_3980,N_2227,N_2367);
xnor U3981 (N_3981,N_2735,N_1878);
or U3982 (N_3982,N_1828,N_2237);
nor U3983 (N_3983,N_2370,N_1951);
nor U3984 (N_3984,N_1589,N_1992);
xor U3985 (N_3985,N_2937,N_2015);
nand U3986 (N_3986,N_1858,N_2090);
nand U3987 (N_3987,N_2069,N_2705);
nor U3988 (N_3988,N_2044,N_2563);
nor U3989 (N_3989,N_1681,N_2965);
and U3990 (N_3990,N_2255,N_1912);
xor U3991 (N_3991,N_2607,N_2358);
or U3992 (N_3992,N_2840,N_2200);
xnor U3993 (N_3993,N_1617,N_2666);
nand U3994 (N_3994,N_1666,N_2698);
nor U3995 (N_3995,N_2952,N_2503);
nor U3996 (N_3996,N_2965,N_2245);
and U3997 (N_3997,N_2297,N_2604);
or U3998 (N_3998,N_2731,N_2227);
nand U3999 (N_3999,N_2822,N_2185);
nand U4000 (N_4000,N_1767,N_2149);
nand U4001 (N_4001,N_2244,N_1816);
xnor U4002 (N_4002,N_1794,N_2799);
and U4003 (N_4003,N_2639,N_2898);
xnor U4004 (N_4004,N_2478,N_1979);
or U4005 (N_4005,N_2488,N_1716);
nor U4006 (N_4006,N_2857,N_1867);
or U4007 (N_4007,N_2856,N_2218);
nor U4008 (N_4008,N_2139,N_1884);
or U4009 (N_4009,N_2629,N_2207);
and U4010 (N_4010,N_1602,N_2472);
xor U4011 (N_4011,N_2227,N_2546);
and U4012 (N_4012,N_2527,N_2111);
and U4013 (N_4013,N_1628,N_2056);
nand U4014 (N_4014,N_2195,N_2732);
nor U4015 (N_4015,N_1631,N_1991);
or U4016 (N_4016,N_2984,N_2265);
or U4017 (N_4017,N_2206,N_2342);
nor U4018 (N_4018,N_2433,N_2768);
or U4019 (N_4019,N_2319,N_1603);
or U4020 (N_4020,N_2525,N_2103);
and U4021 (N_4021,N_2816,N_1717);
nand U4022 (N_4022,N_1603,N_2575);
xor U4023 (N_4023,N_2247,N_1891);
nor U4024 (N_4024,N_2372,N_2290);
and U4025 (N_4025,N_1959,N_2901);
nor U4026 (N_4026,N_2351,N_1628);
nand U4027 (N_4027,N_2462,N_1938);
nand U4028 (N_4028,N_2931,N_2478);
xnor U4029 (N_4029,N_2506,N_1737);
or U4030 (N_4030,N_1736,N_2888);
and U4031 (N_4031,N_1994,N_1519);
or U4032 (N_4032,N_2406,N_1980);
xnor U4033 (N_4033,N_2487,N_2706);
nand U4034 (N_4034,N_1585,N_2621);
xor U4035 (N_4035,N_2890,N_2459);
and U4036 (N_4036,N_1858,N_2872);
or U4037 (N_4037,N_2017,N_1904);
and U4038 (N_4038,N_1683,N_2465);
xor U4039 (N_4039,N_1994,N_2471);
nand U4040 (N_4040,N_1845,N_2759);
nand U4041 (N_4041,N_2273,N_1701);
or U4042 (N_4042,N_2635,N_2895);
or U4043 (N_4043,N_1602,N_1877);
or U4044 (N_4044,N_2230,N_1896);
or U4045 (N_4045,N_2710,N_2883);
nand U4046 (N_4046,N_2070,N_1692);
nor U4047 (N_4047,N_1926,N_1662);
nor U4048 (N_4048,N_2847,N_1902);
xnor U4049 (N_4049,N_2876,N_1946);
nor U4050 (N_4050,N_2703,N_2714);
and U4051 (N_4051,N_2202,N_1593);
nand U4052 (N_4052,N_2302,N_2140);
and U4053 (N_4053,N_2868,N_1691);
xnor U4054 (N_4054,N_1750,N_2250);
nor U4055 (N_4055,N_2350,N_2269);
xnor U4056 (N_4056,N_2633,N_2294);
xor U4057 (N_4057,N_2613,N_2190);
and U4058 (N_4058,N_2127,N_2201);
nand U4059 (N_4059,N_2621,N_2203);
xnor U4060 (N_4060,N_2875,N_2588);
xnor U4061 (N_4061,N_2612,N_2089);
or U4062 (N_4062,N_2926,N_2485);
xor U4063 (N_4063,N_2554,N_2134);
or U4064 (N_4064,N_1852,N_2435);
and U4065 (N_4065,N_2284,N_2283);
nor U4066 (N_4066,N_1891,N_1795);
and U4067 (N_4067,N_2059,N_2782);
nand U4068 (N_4068,N_2768,N_2267);
nor U4069 (N_4069,N_2713,N_2213);
xnor U4070 (N_4070,N_2740,N_2900);
nand U4071 (N_4071,N_1960,N_1867);
or U4072 (N_4072,N_2233,N_2615);
or U4073 (N_4073,N_2260,N_2976);
and U4074 (N_4074,N_1602,N_2610);
nand U4075 (N_4075,N_1922,N_1759);
and U4076 (N_4076,N_1592,N_1943);
nor U4077 (N_4077,N_2278,N_2698);
or U4078 (N_4078,N_2627,N_1721);
or U4079 (N_4079,N_2939,N_2938);
xnor U4080 (N_4080,N_1745,N_2757);
xor U4081 (N_4081,N_1973,N_1936);
or U4082 (N_4082,N_2295,N_2419);
and U4083 (N_4083,N_2551,N_2781);
xnor U4084 (N_4084,N_1629,N_2400);
nand U4085 (N_4085,N_2631,N_2149);
or U4086 (N_4086,N_2262,N_1903);
xnor U4087 (N_4087,N_1646,N_2136);
and U4088 (N_4088,N_2554,N_2282);
nor U4089 (N_4089,N_1878,N_2570);
xnor U4090 (N_4090,N_1636,N_2904);
nand U4091 (N_4091,N_2530,N_2942);
or U4092 (N_4092,N_1887,N_2900);
and U4093 (N_4093,N_2148,N_1558);
xnor U4094 (N_4094,N_1979,N_1588);
xnor U4095 (N_4095,N_2218,N_1786);
xor U4096 (N_4096,N_1638,N_1582);
and U4097 (N_4097,N_2734,N_2667);
nor U4098 (N_4098,N_2711,N_1960);
nand U4099 (N_4099,N_1702,N_2296);
nor U4100 (N_4100,N_2737,N_1845);
nand U4101 (N_4101,N_1786,N_2069);
or U4102 (N_4102,N_2711,N_2185);
nand U4103 (N_4103,N_1608,N_2279);
xnor U4104 (N_4104,N_1970,N_2806);
or U4105 (N_4105,N_1714,N_2404);
nor U4106 (N_4106,N_2100,N_2102);
or U4107 (N_4107,N_2297,N_1982);
nand U4108 (N_4108,N_2886,N_2338);
and U4109 (N_4109,N_2585,N_2381);
or U4110 (N_4110,N_1650,N_2358);
and U4111 (N_4111,N_1838,N_2602);
nor U4112 (N_4112,N_1585,N_2191);
and U4113 (N_4113,N_2865,N_1897);
or U4114 (N_4114,N_2114,N_2761);
and U4115 (N_4115,N_2012,N_2073);
xnor U4116 (N_4116,N_2218,N_2157);
nand U4117 (N_4117,N_2179,N_1519);
xor U4118 (N_4118,N_2357,N_2642);
nor U4119 (N_4119,N_1735,N_1830);
nor U4120 (N_4120,N_2522,N_2613);
xor U4121 (N_4121,N_2181,N_1747);
nand U4122 (N_4122,N_2252,N_1568);
or U4123 (N_4123,N_2654,N_1641);
nand U4124 (N_4124,N_2075,N_2453);
nor U4125 (N_4125,N_1894,N_1674);
nor U4126 (N_4126,N_2284,N_1547);
xnor U4127 (N_4127,N_2374,N_1826);
nor U4128 (N_4128,N_2218,N_2551);
and U4129 (N_4129,N_1821,N_1830);
nor U4130 (N_4130,N_2130,N_2512);
xnor U4131 (N_4131,N_2964,N_2226);
or U4132 (N_4132,N_2262,N_2088);
nor U4133 (N_4133,N_1889,N_2579);
nand U4134 (N_4134,N_2846,N_2670);
or U4135 (N_4135,N_1531,N_2422);
xnor U4136 (N_4136,N_2940,N_1731);
or U4137 (N_4137,N_2370,N_2000);
nand U4138 (N_4138,N_2676,N_2989);
nor U4139 (N_4139,N_2637,N_2875);
nand U4140 (N_4140,N_1501,N_2609);
xor U4141 (N_4141,N_1900,N_2856);
or U4142 (N_4142,N_1846,N_2655);
nand U4143 (N_4143,N_2521,N_2010);
nand U4144 (N_4144,N_2250,N_1963);
nor U4145 (N_4145,N_1942,N_2643);
and U4146 (N_4146,N_2580,N_2159);
xnor U4147 (N_4147,N_2994,N_1607);
or U4148 (N_4148,N_2237,N_2181);
xor U4149 (N_4149,N_2779,N_1790);
nand U4150 (N_4150,N_2576,N_2732);
or U4151 (N_4151,N_2506,N_2318);
nor U4152 (N_4152,N_2990,N_2924);
nor U4153 (N_4153,N_1553,N_1788);
or U4154 (N_4154,N_2882,N_2339);
nand U4155 (N_4155,N_2842,N_1741);
nand U4156 (N_4156,N_2276,N_2729);
xor U4157 (N_4157,N_2730,N_2215);
nor U4158 (N_4158,N_1859,N_1930);
nor U4159 (N_4159,N_2665,N_2153);
and U4160 (N_4160,N_2774,N_2288);
and U4161 (N_4161,N_1743,N_2442);
xor U4162 (N_4162,N_1724,N_2709);
nor U4163 (N_4163,N_2609,N_2553);
nand U4164 (N_4164,N_2408,N_1504);
or U4165 (N_4165,N_2167,N_2395);
xor U4166 (N_4166,N_2210,N_2257);
nand U4167 (N_4167,N_2602,N_2062);
and U4168 (N_4168,N_2023,N_1789);
or U4169 (N_4169,N_1660,N_1547);
nand U4170 (N_4170,N_2566,N_2555);
and U4171 (N_4171,N_2819,N_2477);
nor U4172 (N_4172,N_2955,N_2075);
xnor U4173 (N_4173,N_2844,N_2881);
or U4174 (N_4174,N_2897,N_1842);
nor U4175 (N_4175,N_2518,N_2717);
or U4176 (N_4176,N_2158,N_1798);
nand U4177 (N_4177,N_2011,N_1760);
xor U4178 (N_4178,N_2970,N_1531);
and U4179 (N_4179,N_1657,N_2425);
xnor U4180 (N_4180,N_2508,N_2605);
or U4181 (N_4181,N_2658,N_1719);
nor U4182 (N_4182,N_1996,N_1938);
nor U4183 (N_4183,N_2769,N_2408);
xor U4184 (N_4184,N_1748,N_2309);
nor U4185 (N_4185,N_1551,N_2716);
or U4186 (N_4186,N_2477,N_2610);
and U4187 (N_4187,N_1602,N_1591);
xnor U4188 (N_4188,N_2046,N_1516);
and U4189 (N_4189,N_2980,N_2780);
or U4190 (N_4190,N_2214,N_2721);
nor U4191 (N_4191,N_2129,N_1527);
nor U4192 (N_4192,N_2057,N_2047);
and U4193 (N_4193,N_2468,N_2309);
or U4194 (N_4194,N_1986,N_1935);
nand U4195 (N_4195,N_2062,N_1912);
nor U4196 (N_4196,N_2211,N_1726);
and U4197 (N_4197,N_2124,N_2026);
nand U4198 (N_4198,N_2248,N_2870);
nand U4199 (N_4199,N_2225,N_2754);
xnor U4200 (N_4200,N_2996,N_2644);
or U4201 (N_4201,N_2491,N_2414);
and U4202 (N_4202,N_2011,N_2365);
xnor U4203 (N_4203,N_2995,N_2599);
nand U4204 (N_4204,N_2556,N_2247);
nand U4205 (N_4205,N_2329,N_2582);
or U4206 (N_4206,N_1540,N_2122);
or U4207 (N_4207,N_2205,N_2636);
or U4208 (N_4208,N_2858,N_2460);
or U4209 (N_4209,N_2025,N_1799);
and U4210 (N_4210,N_1868,N_2547);
or U4211 (N_4211,N_1905,N_1959);
xnor U4212 (N_4212,N_2514,N_1823);
xnor U4213 (N_4213,N_2582,N_2634);
nand U4214 (N_4214,N_2672,N_2318);
or U4215 (N_4215,N_1692,N_2801);
xor U4216 (N_4216,N_1622,N_2639);
and U4217 (N_4217,N_2375,N_1803);
and U4218 (N_4218,N_2151,N_1824);
and U4219 (N_4219,N_2047,N_1962);
and U4220 (N_4220,N_1874,N_2890);
nor U4221 (N_4221,N_1740,N_1657);
and U4222 (N_4222,N_1656,N_1854);
nor U4223 (N_4223,N_1644,N_2572);
nor U4224 (N_4224,N_1513,N_2431);
and U4225 (N_4225,N_1552,N_1964);
nor U4226 (N_4226,N_2503,N_2014);
and U4227 (N_4227,N_2932,N_1924);
and U4228 (N_4228,N_1932,N_2436);
and U4229 (N_4229,N_2776,N_2392);
or U4230 (N_4230,N_1508,N_2032);
nor U4231 (N_4231,N_2278,N_1962);
xnor U4232 (N_4232,N_2765,N_1647);
or U4233 (N_4233,N_2652,N_2431);
xor U4234 (N_4234,N_1929,N_2637);
and U4235 (N_4235,N_1957,N_1831);
nor U4236 (N_4236,N_2085,N_1641);
xor U4237 (N_4237,N_2083,N_2893);
nor U4238 (N_4238,N_2594,N_2953);
or U4239 (N_4239,N_2485,N_2417);
or U4240 (N_4240,N_2808,N_1717);
and U4241 (N_4241,N_2783,N_2518);
and U4242 (N_4242,N_2850,N_1576);
xor U4243 (N_4243,N_1536,N_2384);
nand U4244 (N_4244,N_2496,N_1765);
nand U4245 (N_4245,N_1794,N_2780);
and U4246 (N_4246,N_2472,N_2081);
nor U4247 (N_4247,N_1622,N_2387);
nand U4248 (N_4248,N_1535,N_2533);
and U4249 (N_4249,N_1674,N_1505);
nand U4250 (N_4250,N_1970,N_2792);
and U4251 (N_4251,N_2792,N_2137);
and U4252 (N_4252,N_2895,N_1592);
nor U4253 (N_4253,N_2556,N_2220);
or U4254 (N_4254,N_2816,N_2996);
nand U4255 (N_4255,N_1856,N_2383);
xor U4256 (N_4256,N_2351,N_1835);
nor U4257 (N_4257,N_2641,N_2549);
nor U4258 (N_4258,N_2728,N_2242);
xor U4259 (N_4259,N_1735,N_2003);
or U4260 (N_4260,N_2503,N_2362);
xnor U4261 (N_4261,N_1673,N_1991);
xor U4262 (N_4262,N_2525,N_1738);
and U4263 (N_4263,N_1564,N_1532);
xor U4264 (N_4264,N_1831,N_2880);
nor U4265 (N_4265,N_2966,N_1776);
nor U4266 (N_4266,N_1538,N_2747);
or U4267 (N_4267,N_2595,N_1562);
nor U4268 (N_4268,N_1681,N_2272);
xnor U4269 (N_4269,N_2676,N_2767);
nand U4270 (N_4270,N_2982,N_2612);
nor U4271 (N_4271,N_1896,N_2107);
nand U4272 (N_4272,N_2792,N_1776);
or U4273 (N_4273,N_2378,N_2566);
nand U4274 (N_4274,N_2719,N_2083);
nand U4275 (N_4275,N_2150,N_1596);
xor U4276 (N_4276,N_2333,N_2577);
or U4277 (N_4277,N_2703,N_1595);
or U4278 (N_4278,N_2369,N_1605);
xor U4279 (N_4279,N_2117,N_2150);
xor U4280 (N_4280,N_2628,N_2673);
and U4281 (N_4281,N_2252,N_1788);
and U4282 (N_4282,N_2191,N_2416);
nor U4283 (N_4283,N_2541,N_2797);
nor U4284 (N_4284,N_1726,N_1826);
and U4285 (N_4285,N_2257,N_2196);
xnor U4286 (N_4286,N_1698,N_2288);
nor U4287 (N_4287,N_2209,N_1794);
xnor U4288 (N_4288,N_1971,N_1794);
nor U4289 (N_4289,N_2602,N_1572);
nor U4290 (N_4290,N_1709,N_2070);
and U4291 (N_4291,N_2689,N_2113);
and U4292 (N_4292,N_2936,N_2585);
nand U4293 (N_4293,N_2081,N_1536);
and U4294 (N_4294,N_2161,N_1957);
nand U4295 (N_4295,N_2630,N_1615);
nand U4296 (N_4296,N_1803,N_2695);
and U4297 (N_4297,N_1580,N_1659);
or U4298 (N_4298,N_2965,N_2863);
nand U4299 (N_4299,N_2717,N_2501);
or U4300 (N_4300,N_2437,N_1731);
nand U4301 (N_4301,N_2993,N_2910);
nor U4302 (N_4302,N_2625,N_2238);
or U4303 (N_4303,N_2465,N_1761);
xnor U4304 (N_4304,N_1956,N_2198);
nor U4305 (N_4305,N_2636,N_2404);
and U4306 (N_4306,N_1651,N_2788);
nand U4307 (N_4307,N_2235,N_2594);
nand U4308 (N_4308,N_2663,N_2240);
and U4309 (N_4309,N_2574,N_2266);
or U4310 (N_4310,N_2432,N_1863);
xor U4311 (N_4311,N_2259,N_2708);
nor U4312 (N_4312,N_2502,N_2526);
nor U4313 (N_4313,N_1549,N_1590);
and U4314 (N_4314,N_2597,N_1803);
nor U4315 (N_4315,N_1961,N_2286);
nand U4316 (N_4316,N_1617,N_2384);
and U4317 (N_4317,N_2646,N_1554);
or U4318 (N_4318,N_1559,N_1609);
or U4319 (N_4319,N_1645,N_2292);
nand U4320 (N_4320,N_2805,N_2259);
or U4321 (N_4321,N_2530,N_2869);
nor U4322 (N_4322,N_2988,N_2236);
xnor U4323 (N_4323,N_2685,N_2624);
or U4324 (N_4324,N_2542,N_2694);
and U4325 (N_4325,N_1835,N_2077);
xnor U4326 (N_4326,N_2150,N_2068);
nor U4327 (N_4327,N_1916,N_2208);
nand U4328 (N_4328,N_2832,N_2271);
xor U4329 (N_4329,N_2918,N_2660);
nand U4330 (N_4330,N_2671,N_2330);
nor U4331 (N_4331,N_2504,N_2929);
xnor U4332 (N_4332,N_2979,N_2888);
or U4333 (N_4333,N_2267,N_1924);
nand U4334 (N_4334,N_2021,N_1725);
xor U4335 (N_4335,N_2071,N_2215);
nor U4336 (N_4336,N_2379,N_2751);
nor U4337 (N_4337,N_2682,N_2509);
nor U4338 (N_4338,N_2629,N_2086);
nand U4339 (N_4339,N_2811,N_1766);
nor U4340 (N_4340,N_2113,N_2703);
xor U4341 (N_4341,N_2357,N_2573);
nand U4342 (N_4342,N_1874,N_1718);
xnor U4343 (N_4343,N_2634,N_2814);
nor U4344 (N_4344,N_2248,N_1773);
xnor U4345 (N_4345,N_1902,N_2116);
nor U4346 (N_4346,N_2767,N_2845);
nand U4347 (N_4347,N_2150,N_2848);
or U4348 (N_4348,N_2145,N_2987);
or U4349 (N_4349,N_2280,N_2008);
and U4350 (N_4350,N_2365,N_2122);
nor U4351 (N_4351,N_1932,N_1685);
xor U4352 (N_4352,N_2383,N_2494);
or U4353 (N_4353,N_2276,N_2688);
xor U4354 (N_4354,N_1953,N_2785);
nand U4355 (N_4355,N_2746,N_2231);
or U4356 (N_4356,N_1561,N_2449);
nor U4357 (N_4357,N_2696,N_2019);
nand U4358 (N_4358,N_1561,N_2857);
xnor U4359 (N_4359,N_1940,N_2563);
xnor U4360 (N_4360,N_2981,N_1692);
nor U4361 (N_4361,N_1700,N_2990);
nand U4362 (N_4362,N_1577,N_2049);
nand U4363 (N_4363,N_1547,N_2440);
xnor U4364 (N_4364,N_2863,N_2320);
nor U4365 (N_4365,N_2306,N_1886);
nor U4366 (N_4366,N_2841,N_2139);
or U4367 (N_4367,N_2902,N_2109);
xor U4368 (N_4368,N_2756,N_2153);
nor U4369 (N_4369,N_2375,N_2940);
xor U4370 (N_4370,N_2847,N_2976);
nand U4371 (N_4371,N_2445,N_2395);
and U4372 (N_4372,N_2849,N_2339);
nor U4373 (N_4373,N_1576,N_2326);
nand U4374 (N_4374,N_2427,N_1961);
xnor U4375 (N_4375,N_2890,N_2360);
or U4376 (N_4376,N_1517,N_1967);
nand U4377 (N_4377,N_2244,N_2233);
xnor U4378 (N_4378,N_2728,N_1623);
nor U4379 (N_4379,N_1776,N_2354);
or U4380 (N_4380,N_2219,N_1915);
xnor U4381 (N_4381,N_2677,N_1703);
nand U4382 (N_4382,N_2105,N_1983);
nand U4383 (N_4383,N_1950,N_2292);
xnor U4384 (N_4384,N_2748,N_2425);
xnor U4385 (N_4385,N_2520,N_1782);
xnor U4386 (N_4386,N_2891,N_2138);
and U4387 (N_4387,N_2715,N_2319);
nand U4388 (N_4388,N_2586,N_2226);
or U4389 (N_4389,N_2135,N_2584);
xor U4390 (N_4390,N_2605,N_2246);
xnor U4391 (N_4391,N_1797,N_1668);
and U4392 (N_4392,N_2099,N_2639);
nand U4393 (N_4393,N_2384,N_2824);
nor U4394 (N_4394,N_2912,N_2199);
and U4395 (N_4395,N_2983,N_2873);
nor U4396 (N_4396,N_2728,N_1686);
nand U4397 (N_4397,N_2376,N_2154);
and U4398 (N_4398,N_2984,N_2886);
nor U4399 (N_4399,N_2525,N_1718);
nor U4400 (N_4400,N_1941,N_2853);
and U4401 (N_4401,N_2281,N_2476);
and U4402 (N_4402,N_2603,N_2030);
or U4403 (N_4403,N_1658,N_2309);
or U4404 (N_4404,N_1724,N_2490);
and U4405 (N_4405,N_1567,N_2819);
or U4406 (N_4406,N_1601,N_2824);
and U4407 (N_4407,N_2178,N_2493);
nand U4408 (N_4408,N_2328,N_1506);
xnor U4409 (N_4409,N_2579,N_1596);
nor U4410 (N_4410,N_2763,N_2691);
nand U4411 (N_4411,N_1547,N_2349);
nor U4412 (N_4412,N_1985,N_1675);
nor U4413 (N_4413,N_2728,N_2384);
xor U4414 (N_4414,N_2519,N_2570);
or U4415 (N_4415,N_1506,N_1738);
and U4416 (N_4416,N_1897,N_1518);
and U4417 (N_4417,N_1978,N_2225);
xor U4418 (N_4418,N_1793,N_1744);
and U4419 (N_4419,N_2318,N_2699);
nor U4420 (N_4420,N_2945,N_2898);
xnor U4421 (N_4421,N_2310,N_2657);
or U4422 (N_4422,N_2170,N_2712);
and U4423 (N_4423,N_2815,N_2309);
nor U4424 (N_4424,N_2984,N_1692);
or U4425 (N_4425,N_2092,N_1945);
nand U4426 (N_4426,N_2351,N_1806);
nor U4427 (N_4427,N_2710,N_2441);
or U4428 (N_4428,N_2579,N_2156);
nand U4429 (N_4429,N_2415,N_1746);
and U4430 (N_4430,N_2252,N_2297);
or U4431 (N_4431,N_1706,N_2199);
or U4432 (N_4432,N_1660,N_2329);
or U4433 (N_4433,N_2610,N_1558);
nor U4434 (N_4434,N_2330,N_2378);
nor U4435 (N_4435,N_2450,N_2928);
and U4436 (N_4436,N_2088,N_1965);
xnor U4437 (N_4437,N_1829,N_1835);
nand U4438 (N_4438,N_2434,N_2770);
xnor U4439 (N_4439,N_2464,N_2944);
xnor U4440 (N_4440,N_2208,N_2092);
xnor U4441 (N_4441,N_2060,N_2300);
nand U4442 (N_4442,N_2569,N_2186);
xnor U4443 (N_4443,N_2782,N_2385);
and U4444 (N_4444,N_2337,N_2752);
nand U4445 (N_4445,N_2523,N_1608);
nand U4446 (N_4446,N_2046,N_1703);
xnor U4447 (N_4447,N_2769,N_1685);
nor U4448 (N_4448,N_1782,N_2208);
and U4449 (N_4449,N_2041,N_2015);
or U4450 (N_4450,N_2663,N_2770);
and U4451 (N_4451,N_2670,N_2861);
xor U4452 (N_4452,N_2129,N_2829);
and U4453 (N_4453,N_1806,N_2779);
and U4454 (N_4454,N_2775,N_1573);
nand U4455 (N_4455,N_1928,N_2718);
xnor U4456 (N_4456,N_2482,N_2892);
xor U4457 (N_4457,N_2607,N_1972);
nand U4458 (N_4458,N_2789,N_2363);
nor U4459 (N_4459,N_2503,N_2600);
xnor U4460 (N_4460,N_1866,N_2553);
and U4461 (N_4461,N_1744,N_2038);
xor U4462 (N_4462,N_1984,N_1545);
nor U4463 (N_4463,N_1788,N_2437);
or U4464 (N_4464,N_2899,N_1840);
nand U4465 (N_4465,N_1922,N_2459);
xor U4466 (N_4466,N_2185,N_2808);
nand U4467 (N_4467,N_2319,N_2505);
and U4468 (N_4468,N_1747,N_1636);
nand U4469 (N_4469,N_1670,N_2521);
or U4470 (N_4470,N_2321,N_2075);
xor U4471 (N_4471,N_2577,N_2217);
or U4472 (N_4472,N_2712,N_1561);
and U4473 (N_4473,N_2919,N_2335);
and U4474 (N_4474,N_2176,N_2401);
and U4475 (N_4475,N_1670,N_2125);
nand U4476 (N_4476,N_2526,N_1911);
nor U4477 (N_4477,N_1566,N_2405);
or U4478 (N_4478,N_1529,N_2469);
or U4479 (N_4479,N_2090,N_1722);
xor U4480 (N_4480,N_1890,N_1733);
nor U4481 (N_4481,N_2199,N_1996);
xor U4482 (N_4482,N_2795,N_2174);
or U4483 (N_4483,N_2161,N_2553);
and U4484 (N_4484,N_1953,N_2617);
or U4485 (N_4485,N_1912,N_2980);
nand U4486 (N_4486,N_2037,N_2736);
nand U4487 (N_4487,N_1686,N_2984);
and U4488 (N_4488,N_2383,N_2537);
or U4489 (N_4489,N_1730,N_1619);
nor U4490 (N_4490,N_2031,N_1776);
and U4491 (N_4491,N_2034,N_2648);
or U4492 (N_4492,N_1749,N_1919);
nand U4493 (N_4493,N_2993,N_2677);
xor U4494 (N_4494,N_1723,N_1952);
nor U4495 (N_4495,N_2118,N_2251);
or U4496 (N_4496,N_2656,N_2825);
xnor U4497 (N_4497,N_2755,N_2385);
nor U4498 (N_4498,N_2387,N_2455);
nor U4499 (N_4499,N_1538,N_1754);
and U4500 (N_4500,N_3046,N_3505);
nand U4501 (N_4501,N_4178,N_3243);
and U4502 (N_4502,N_3453,N_3765);
or U4503 (N_4503,N_3360,N_3784);
and U4504 (N_4504,N_3574,N_3860);
and U4505 (N_4505,N_3473,N_4002);
and U4506 (N_4506,N_3682,N_3768);
or U4507 (N_4507,N_4031,N_3281);
nor U4508 (N_4508,N_3304,N_4399);
and U4509 (N_4509,N_4317,N_3322);
or U4510 (N_4510,N_3001,N_3769);
nor U4511 (N_4511,N_4411,N_4400);
nand U4512 (N_4512,N_4352,N_4386);
and U4513 (N_4513,N_3987,N_4013);
nor U4514 (N_4514,N_4493,N_3671);
nand U4515 (N_4515,N_3502,N_4329);
nor U4516 (N_4516,N_3020,N_3255);
nor U4517 (N_4517,N_3704,N_3551);
xnor U4518 (N_4518,N_4026,N_3115);
and U4519 (N_4519,N_4402,N_3374);
xnor U4520 (N_4520,N_3880,N_4180);
nor U4521 (N_4521,N_3073,N_3145);
or U4522 (N_4522,N_3938,N_4005);
nand U4523 (N_4523,N_3324,N_3434);
nand U4524 (N_4524,N_3101,N_3925);
nor U4525 (N_4525,N_4405,N_3107);
or U4526 (N_4526,N_4189,N_3709);
or U4527 (N_4527,N_3189,N_4122);
or U4528 (N_4528,N_3516,N_4255);
and U4529 (N_4529,N_3405,N_3681);
xor U4530 (N_4530,N_3592,N_3290);
xnor U4531 (N_4531,N_3264,N_3526);
nand U4532 (N_4532,N_3731,N_3739);
nand U4533 (N_4533,N_3433,N_3685);
or U4534 (N_4534,N_3150,N_3156);
xnor U4535 (N_4535,N_3792,N_4258);
nor U4536 (N_4536,N_3003,N_4210);
or U4537 (N_4537,N_4024,N_4312);
nand U4538 (N_4538,N_3440,N_3445);
nand U4539 (N_4539,N_4141,N_3665);
or U4540 (N_4540,N_3999,N_3241);
nand U4541 (N_4541,N_4269,N_3287);
and U4542 (N_4542,N_3129,N_4135);
nand U4543 (N_4543,N_3175,N_3836);
nand U4544 (N_4544,N_3154,N_3949);
nor U4545 (N_4545,N_3057,N_3247);
and U4546 (N_4546,N_4191,N_3415);
and U4547 (N_4547,N_3518,N_4345);
nand U4548 (N_4548,N_4254,N_4334);
xnor U4549 (N_4549,N_3767,N_4415);
nor U4550 (N_4550,N_3441,N_3985);
xnor U4551 (N_4551,N_3418,N_3855);
xnor U4552 (N_4552,N_3652,N_3978);
and U4553 (N_4553,N_3967,N_3561);
or U4554 (N_4554,N_3104,N_4357);
nand U4555 (N_4555,N_3818,N_3893);
nand U4556 (N_4556,N_4459,N_4238);
nor U4557 (N_4557,N_3948,N_4052);
or U4558 (N_4558,N_4124,N_3197);
xor U4559 (N_4559,N_4398,N_3598);
nor U4560 (N_4560,N_4030,N_3383);
and U4561 (N_4561,N_3538,N_4051);
nand U4562 (N_4562,N_3071,N_3402);
nand U4563 (N_4563,N_4170,N_3930);
and U4564 (N_4564,N_3299,N_3063);
or U4565 (N_4565,N_3074,N_4097);
and U4566 (N_4566,N_3379,N_4251);
xor U4567 (N_4567,N_4145,N_4166);
and U4568 (N_4568,N_3958,N_3636);
or U4569 (N_4569,N_3781,N_3677);
xor U4570 (N_4570,N_3325,N_3966);
xor U4571 (N_4571,N_3594,N_3075);
nand U4572 (N_4572,N_3267,N_4136);
nor U4573 (N_4573,N_3779,N_4098);
nand U4574 (N_4574,N_4094,N_3376);
or U4575 (N_4575,N_4279,N_3220);
nand U4576 (N_4576,N_3041,N_3599);
nor U4577 (N_4577,N_3435,N_3806);
and U4578 (N_4578,N_3161,N_4343);
xnor U4579 (N_4579,N_3457,N_3712);
xor U4580 (N_4580,N_3149,N_4099);
or U4581 (N_4581,N_3761,N_3400);
nand U4582 (N_4582,N_4483,N_3375);
and U4583 (N_4583,N_3586,N_3790);
and U4584 (N_4584,N_3483,N_4028);
nor U4585 (N_4585,N_3617,N_3625);
xnor U4586 (N_4586,N_3662,N_4445);
nor U4587 (N_4587,N_3979,N_3755);
nand U4588 (N_4588,N_3113,N_3294);
and U4589 (N_4589,N_3633,N_4292);
or U4590 (N_4590,N_4486,N_4425);
nor U4591 (N_4591,N_3648,N_3173);
and U4592 (N_4592,N_4195,N_3248);
nand U4593 (N_4593,N_3621,N_3749);
and U4594 (N_4594,N_3286,N_3968);
xor U4595 (N_4595,N_3766,N_3077);
nand U4596 (N_4596,N_4117,N_4440);
xor U4597 (N_4597,N_4340,N_3803);
nor U4598 (N_4598,N_3411,N_3942);
or U4599 (N_4599,N_3618,N_4139);
or U4600 (N_4600,N_3353,N_4320);
nor U4601 (N_4601,N_3035,N_3345);
nand U4602 (N_4602,N_3794,N_4457);
nand U4603 (N_4603,N_3488,N_3686);
nor U4604 (N_4604,N_3951,N_3996);
nand U4605 (N_4605,N_4046,N_4370);
or U4606 (N_4606,N_3829,N_3280);
xor U4607 (N_4607,N_3461,N_3399);
and U4608 (N_4608,N_3807,N_4385);
nor U4609 (N_4609,N_3357,N_4092);
nor U4610 (N_4610,N_3471,N_3065);
or U4611 (N_4611,N_4042,N_3301);
nor U4612 (N_4612,N_4147,N_3036);
or U4613 (N_4613,N_3438,N_3560);
or U4614 (N_4614,N_3506,N_3995);
and U4615 (N_4615,N_4077,N_3130);
and U4616 (N_4616,N_4430,N_3510);
or U4617 (N_4617,N_3187,N_3827);
or U4618 (N_4618,N_3038,N_3170);
and U4619 (N_4619,N_3311,N_3689);
nand U4620 (N_4620,N_3511,N_3935);
nor U4621 (N_4621,N_4346,N_4218);
and U4622 (N_4622,N_4290,N_3292);
nor U4623 (N_4623,N_3657,N_3832);
xnor U4624 (N_4624,N_4164,N_4194);
or U4625 (N_4625,N_4458,N_4216);
nor U4626 (N_4626,N_3229,N_4333);
and U4627 (N_4627,N_3080,N_3040);
nor U4628 (N_4628,N_4332,N_3437);
or U4629 (N_4629,N_3959,N_3016);
nand U4630 (N_4630,N_3257,N_3915);
nand U4631 (N_4631,N_4416,N_3097);
xor U4632 (N_4632,N_3004,N_3477);
nand U4633 (N_4633,N_3941,N_3205);
or U4634 (N_4634,N_3815,N_3992);
and U4635 (N_4635,N_4066,N_4063);
or U4636 (N_4636,N_3796,N_4132);
xnor U4637 (N_4637,N_4438,N_4184);
xnor U4638 (N_4638,N_3328,N_3495);
and U4639 (N_4639,N_4471,N_4219);
nand U4640 (N_4640,N_3470,N_4101);
or U4641 (N_4641,N_4085,N_4015);
nand U4642 (N_4642,N_3349,N_3939);
and U4643 (N_4643,N_3868,N_3552);
or U4644 (N_4644,N_3913,N_4247);
nor U4645 (N_4645,N_3982,N_3244);
nand U4646 (N_4646,N_4494,N_4225);
xnor U4647 (N_4647,N_3603,N_4050);
or U4648 (N_4648,N_4499,N_3122);
or U4649 (N_4649,N_3578,N_3033);
and U4650 (N_4650,N_3158,N_3607);
nor U4651 (N_4651,N_3427,N_3312);
xnor U4652 (N_4652,N_3953,N_3852);
or U4653 (N_4653,N_3523,N_3678);
or U4654 (N_4654,N_4300,N_3947);
nand U4655 (N_4655,N_3031,N_3697);
nor U4656 (N_4656,N_3023,N_3305);
xor U4657 (N_4657,N_4082,N_4162);
or U4658 (N_4658,N_3624,N_3562);
nor U4659 (N_4659,N_3017,N_4177);
xor U4660 (N_4660,N_4442,N_4153);
nand U4661 (N_4661,N_4463,N_4407);
nor U4662 (N_4662,N_3593,N_4091);
xnor U4663 (N_4663,N_3088,N_4389);
or U4664 (N_4664,N_4263,N_3507);
and U4665 (N_4665,N_3310,N_3135);
and U4666 (N_4666,N_4485,N_4439);
or U4667 (N_4667,N_3112,N_4070);
nor U4668 (N_4668,N_4133,N_3386);
or U4669 (N_4669,N_3645,N_3820);
or U4670 (N_4670,N_3320,N_3791);
xor U4671 (N_4671,N_4409,N_3174);
nor U4672 (N_4672,N_3332,N_3045);
xnor U4673 (N_4673,N_3447,N_3192);
xnor U4674 (N_4674,N_3724,N_4327);
xor U4675 (N_4675,N_3927,N_4404);
and U4676 (N_4676,N_3034,N_3632);
or U4677 (N_4677,N_3185,N_4110);
xnor U4678 (N_4678,N_4296,N_3850);
nand U4679 (N_4679,N_3250,N_4089);
and U4680 (N_4680,N_3917,N_3943);
xnor U4681 (N_4681,N_4281,N_3335);
xnor U4682 (N_4682,N_3690,N_3843);
nand U4683 (N_4683,N_4201,N_4473);
and U4684 (N_4684,N_4237,N_3898);
xnor U4685 (N_4685,N_4149,N_3459);
nor U4686 (N_4686,N_3343,N_3133);
and U4687 (N_4687,N_3078,N_3841);
xnor U4688 (N_4688,N_4016,N_3907);
or U4689 (N_4689,N_3619,N_4331);
and U4690 (N_4690,N_4093,N_3861);
nor U4691 (N_4691,N_4495,N_4420);
or U4692 (N_4692,N_3398,N_4190);
xnor U4693 (N_4693,N_3989,N_4069);
nand U4694 (N_4694,N_4482,N_4088);
xnor U4695 (N_4695,N_4137,N_3816);
xor U4696 (N_4696,N_3740,N_3100);
or U4697 (N_4697,N_3557,N_3647);
nand U4698 (N_4698,N_3475,N_3152);
and U4699 (N_4699,N_3629,N_4062);
xor U4700 (N_4700,N_3472,N_3702);
or U4701 (N_4701,N_4130,N_4007);
nand U4702 (N_4702,N_4232,N_3993);
or U4703 (N_4703,N_3997,N_3454);
nor U4704 (N_4704,N_3567,N_3710);
xnor U4705 (N_4705,N_3916,N_3191);
xnor U4706 (N_4706,N_4221,N_4277);
nor U4707 (N_4707,N_4020,N_3782);
xor U4708 (N_4708,N_3214,N_3971);
or U4709 (N_4709,N_3503,N_3216);
nand U4710 (N_4710,N_4034,N_3872);
or U4711 (N_4711,N_3443,N_3123);
and U4712 (N_4712,N_3222,N_4114);
nor U4713 (N_4713,N_4227,N_3921);
nand U4714 (N_4714,N_4308,N_3810);
nand U4715 (N_4715,N_4150,N_3429);
and U4716 (N_4716,N_4361,N_3641);
and U4717 (N_4717,N_3809,N_3933);
nor U4718 (N_4718,N_3675,N_3487);
or U4719 (N_4719,N_3082,N_3600);
xor U4720 (N_4720,N_3278,N_4228);
nand U4721 (N_4721,N_3556,N_4121);
or U4722 (N_4722,N_3753,N_3414);
nor U4723 (N_4723,N_3478,N_3356);
or U4724 (N_4724,N_3032,N_3109);
nor U4725 (N_4725,N_3079,N_3773);
xnor U4726 (N_4726,N_4033,N_4397);
and U4727 (N_4727,N_3026,N_4017);
nor U4728 (N_4728,N_3204,N_4481);
xnor U4729 (N_4729,N_3742,N_3695);
or U4730 (N_4730,N_3052,N_4090);
and U4731 (N_4731,N_3878,N_3011);
xnor U4732 (N_4732,N_4429,N_3751);
and U4733 (N_4733,N_3849,N_4037);
and U4734 (N_4734,N_4073,N_3616);
nand U4735 (N_4735,N_4220,N_4450);
nor U4736 (N_4736,N_4396,N_3393);
nor U4737 (N_4737,N_4342,N_3548);
and U4738 (N_4738,N_3984,N_3591);
xnor U4739 (N_4739,N_3352,N_3143);
nand U4740 (N_4740,N_4165,N_4198);
nand U4741 (N_4741,N_3846,N_3659);
nor U4742 (N_4742,N_4043,N_4079);
nor U4743 (N_4743,N_3698,N_4241);
nand U4744 (N_4744,N_3851,N_4422);
and U4745 (N_4745,N_3354,N_4128);
nor U4746 (N_4746,N_4154,N_3262);
or U4747 (N_4747,N_3347,N_3330);
nand U4748 (N_4748,N_3277,N_3595);
nor U4749 (N_4749,N_3362,N_3805);
xor U4750 (N_4750,N_3568,N_3608);
nor U4751 (N_4751,N_4120,N_3468);
or U4752 (N_4752,N_4266,N_3159);
and U4753 (N_4753,N_4175,N_3514);
nand U4754 (N_4754,N_3489,N_3882);
or U4755 (N_4755,N_4182,N_4435);
nor U4756 (N_4756,N_3303,N_4081);
or U4757 (N_4757,N_3295,N_3142);
nand U4758 (N_4758,N_3823,N_3572);
nand U4759 (N_4759,N_3327,N_4437);
nand U4760 (N_4760,N_4209,N_3750);
nand U4761 (N_4761,N_3417,N_3355);
xnor U4762 (N_4762,N_3431,N_3000);
xnor U4763 (N_4763,N_4148,N_3723);
and U4764 (N_4764,N_3172,N_3676);
and U4765 (N_4765,N_3237,N_4095);
nor U4766 (N_4766,N_3181,N_3064);
xnor U4767 (N_4767,N_3436,N_4027);
nor U4768 (N_4768,N_4466,N_3008);
and U4769 (N_4769,N_3165,N_3039);
nor U4770 (N_4770,N_4179,N_3961);
or U4771 (N_4771,N_3348,N_3134);
xor U4772 (N_4772,N_4061,N_3654);
and U4773 (N_4773,N_3711,N_4348);
xnor U4774 (N_4774,N_3169,N_3132);
nor U4775 (N_4775,N_3331,N_3946);
xor U4776 (N_4776,N_3637,N_3370);
nor U4777 (N_4777,N_4116,N_4003);
and U4778 (N_4778,N_3642,N_3479);
xor U4779 (N_4779,N_3367,N_3908);
xor U4780 (N_4780,N_4211,N_3455);
xor U4781 (N_4781,N_3825,N_3350);
xnor U4782 (N_4782,N_3053,N_3821);
or U4783 (N_4783,N_3344,N_3308);
nand U4784 (N_4784,N_4284,N_3558);
nand U4785 (N_4785,N_3125,N_3070);
nor U4786 (N_4786,N_3924,N_3426);
and U4787 (N_4787,N_4354,N_4444);
xnor U4788 (N_4788,N_3384,N_3559);
or U4789 (N_4789,N_3474,N_4115);
xor U4790 (N_4790,N_3804,N_3883);
nor U4791 (N_4791,N_3777,N_3911);
nor U4792 (N_4792,N_4204,N_3407);
xnor U4793 (N_4793,N_4246,N_3589);
or U4794 (N_4794,N_4252,N_4140);
or U4795 (N_4795,N_4100,N_4108);
and U4796 (N_4796,N_4183,N_4371);
xnor U4797 (N_4797,N_3144,N_4205);
nor U4798 (N_4798,N_4109,N_3178);
nand U4799 (N_4799,N_4186,N_4375);
or U4800 (N_4800,N_4274,N_3565);
nand U4801 (N_4801,N_4072,N_4282);
nand U4802 (N_4802,N_3381,N_4142);
xor U4803 (N_4803,N_4199,N_4474);
xor U4804 (N_4804,N_3746,N_4301);
nand U4805 (N_4805,N_3148,N_4270);
nand U4806 (N_4806,N_3059,N_4309);
and U4807 (N_4807,N_3266,N_3060);
nand U4808 (N_4808,N_3635,N_3176);
nor U4809 (N_4809,N_3668,N_4229);
or U4810 (N_4810,N_4103,N_3168);
xor U4811 (N_4811,N_4288,N_4169);
nor U4812 (N_4812,N_3166,N_3926);
or U4813 (N_4813,N_4382,N_4298);
nor U4814 (N_4814,N_4000,N_3102);
nor U4815 (N_4815,N_3465,N_3091);
or U4816 (N_4816,N_3021,N_3009);
xnor U4817 (N_4817,N_4259,N_3658);
and U4818 (N_4818,N_4350,N_3279);
and U4819 (N_4819,N_3541,N_3700);
and U4820 (N_4820,N_4452,N_3014);
nor U4821 (N_4821,N_4068,N_3451);
xnor U4822 (N_4822,N_3812,N_3801);
nand U4823 (N_4823,N_3745,N_3814);
and U4824 (N_4824,N_3316,N_3136);
nand U4825 (N_4825,N_3138,N_3201);
nor U4826 (N_4826,N_3061,N_3274);
or U4827 (N_4827,N_3687,N_3094);
nand U4828 (N_4828,N_3177,N_4240);
nor U4829 (N_4829,N_4264,N_4224);
and U4830 (N_4830,N_4231,N_3272);
and U4831 (N_4831,N_4021,N_3265);
nor U4832 (N_4832,N_4161,N_3620);
or U4833 (N_4833,N_4022,N_3162);
xnor U4834 (N_4834,N_4275,N_4160);
xor U4835 (N_4835,N_3164,N_4353);
nor U4836 (N_4836,N_3903,N_3232);
nor U4837 (N_4837,N_4260,N_4470);
xnor U4838 (N_4838,N_4469,N_3242);
or U4839 (N_4839,N_4322,N_3095);
and U4840 (N_4840,N_3936,N_3638);
and U4841 (N_4841,N_4087,N_3691);
xor U4842 (N_4842,N_4086,N_3307);
and U4843 (N_4843,N_4048,N_4324);
or U4844 (N_4844,N_3692,N_4377);
or U4845 (N_4845,N_3547,N_3121);
and U4846 (N_4846,N_3420,N_3391);
nor U4847 (N_4847,N_4223,N_3378);
xor U4848 (N_4848,N_3321,N_3037);
xor U4849 (N_4849,N_3737,N_3928);
nand U4850 (N_4850,N_4498,N_3337);
nor U4851 (N_4851,N_3536,N_4436);
nand U4852 (N_4852,N_4143,N_3890);
and U4853 (N_4853,N_3644,N_4014);
nor U4854 (N_4854,N_3892,N_4384);
xor U4855 (N_4855,N_3452,N_4480);
nand U4856 (N_4856,N_4055,N_3501);
and U4857 (N_4857,N_4291,N_3213);
or U4858 (N_4858,N_3655,N_4339);
nor U4859 (N_4859,N_4200,N_3865);
nand U4860 (N_4860,N_3584,N_3221);
xor U4861 (N_4861,N_3885,N_3854);
nand U4862 (N_4862,N_4302,N_4112);
xnor U4863 (N_4863,N_4041,N_3858);
xor U4864 (N_4864,N_4394,N_3285);
nor U4865 (N_4865,N_4202,N_4239);
nand U4866 (N_4866,N_3628,N_3802);
xor U4867 (N_4867,N_3528,N_3934);
xor U4868 (N_4868,N_4059,N_4113);
nand U4869 (N_4869,N_3464,N_4047);
xnor U4870 (N_4870,N_4158,N_3550);
or U4871 (N_4871,N_3194,N_3537);
nor U4872 (N_4872,N_3298,N_3351);
and U4873 (N_4873,N_4187,N_3891);
and U4874 (N_4874,N_3527,N_4214);
or U4875 (N_4875,N_3975,N_3763);
and U4876 (N_4876,N_3627,N_4387);
or U4877 (N_4877,N_4208,N_3297);
nand U4878 (N_4878,N_4257,N_3534);
xor U4879 (N_4879,N_3207,N_3424);
nor U4880 (N_4880,N_3976,N_3828);
nor U4881 (N_4881,N_4249,N_3602);
and U4882 (N_4882,N_4383,N_3795);
nand U4883 (N_4883,N_3186,N_4197);
or U4884 (N_4884,N_3604,N_3615);
or U4885 (N_4885,N_3529,N_3833);
and U4886 (N_4886,N_4039,N_4476);
nor U4887 (N_4887,N_3482,N_3270);
and U4888 (N_4888,N_4146,N_4134);
and U4889 (N_4889,N_3124,N_4456);
or U4890 (N_4890,N_3099,N_3233);
and U4891 (N_4891,N_4464,N_3910);
and U4892 (N_4892,N_4390,N_4454);
nor U4893 (N_4893,N_3542,N_3899);
and U4894 (N_4894,N_3713,N_4323);
and U4895 (N_4895,N_3896,N_3844);
nand U4896 (N_4896,N_4376,N_4212);
or U4897 (N_4897,N_3089,N_3258);
nand U4898 (N_4898,N_3653,N_3845);
xor U4899 (N_4899,N_3252,N_4360);
and U4900 (N_4900,N_3840,N_3056);
nor U4901 (N_4901,N_3126,N_4076);
xor U4902 (N_4902,N_4156,N_3722);
and U4903 (N_4903,N_4465,N_3081);
or U4904 (N_4904,N_4372,N_3334);
nor U4905 (N_4905,N_3983,N_3043);
nand U4906 (N_4906,N_3022,N_4467);
nand U4907 (N_4907,N_3432,N_4451);
and U4908 (N_4908,N_3359,N_3208);
or U4909 (N_4909,N_3206,N_3006);
nor U4910 (N_4910,N_3778,N_4152);
or U4911 (N_4911,N_3775,N_4049);
and U4912 (N_4912,N_3005,N_3498);
or U4913 (N_4913,N_3042,N_4268);
or U4914 (N_4914,N_4379,N_4267);
nor U4915 (N_4915,N_4431,N_4064);
nand U4916 (N_4916,N_3717,N_4126);
nand U4917 (N_4917,N_3571,N_3634);
xnor U4918 (N_4918,N_3863,N_3922);
nand U4919 (N_4919,N_3480,N_3403);
or U4920 (N_4920,N_4419,N_3314);
nor U4921 (N_4921,N_3067,N_4276);
nor U4922 (N_4922,N_3679,N_4188);
and U4923 (N_4923,N_3952,N_3085);
and U4924 (N_4924,N_3813,N_3062);
nor U4925 (N_4925,N_3111,N_3981);
xor U4926 (N_4926,N_3371,N_3072);
nor U4927 (N_4927,N_3293,N_3396);
nand U4928 (N_4928,N_4297,N_4421);
and U4929 (N_4929,N_3449,N_3630);
and U4930 (N_4930,N_4316,N_3980);
and U4931 (N_4931,N_3467,N_3923);
nand U4932 (N_4932,N_3817,N_3988);
nand U4933 (N_4933,N_4029,N_3365);
or U4934 (N_4934,N_4391,N_3945);
nor U4935 (N_4935,N_4138,N_3881);
nor U4936 (N_4936,N_3199,N_4185);
or U4937 (N_4937,N_3614,N_3597);
or U4938 (N_4938,N_4347,N_3273);
nor U4939 (N_4939,N_3870,N_3289);
or U4940 (N_4940,N_3730,N_3117);
nand U4941 (N_4941,N_3797,N_3228);
and U4942 (N_4942,N_3573,N_4356);
or U4943 (N_4943,N_3302,N_3323);
and U4944 (N_4944,N_3086,N_4172);
nor U4945 (N_4945,N_3744,N_3613);
xor U4946 (N_4946,N_4127,N_4044);
nor U4947 (N_4947,N_4374,N_3030);
and U4948 (N_4948,N_3772,N_4058);
nor U4949 (N_4949,N_3309,N_4412);
and U4950 (N_4950,N_3412,N_4111);
or U4951 (N_4951,N_3512,N_3994);
nor U4952 (N_4952,N_4432,N_3051);
nor U4953 (N_4953,N_3340,N_4299);
or U4954 (N_4954,N_3847,N_4171);
xor U4955 (N_4955,N_4233,N_3196);
nand U4956 (N_4956,N_3463,N_4446);
and U4957 (N_4957,N_3157,N_3069);
and U4958 (N_4958,N_3932,N_3410);
and U4959 (N_4959,N_3533,N_4025);
and U4960 (N_4960,N_3842,N_3387);
nand U4961 (N_4961,N_4181,N_3364);
nor U4962 (N_4962,N_4355,N_3066);
xnor U4963 (N_4963,N_4491,N_3622);
xor U4964 (N_4964,N_3962,N_3377);
or U4965 (N_4965,N_3875,N_4330);
nor U4966 (N_4966,N_3392,N_3105);
nor U4967 (N_4967,N_4380,N_4203);
xnor U4968 (N_4968,N_3050,N_4083);
xor U4969 (N_4969,N_4176,N_3515);
nand U4970 (N_4970,N_4071,N_3239);
nor U4971 (N_4971,N_3920,N_3422);
nor U4972 (N_4972,N_3912,N_4018);
xnor U4973 (N_4973,N_3611,N_3862);
xnor U4974 (N_4974,N_3227,N_3734);
nand U4975 (N_4975,N_3848,N_3888);
nor U4976 (N_4976,N_3098,N_3596);
or U4977 (N_4977,N_3103,N_3373);
nor U4978 (N_4978,N_4448,N_3831);
xnor U4979 (N_4979,N_4487,N_4406);
nor U4980 (N_4980,N_3905,N_3397);
xnor U4981 (N_4981,N_3128,N_4032);
and U4982 (N_4982,N_4490,N_3493);
and U4983 (N_4983,N_3577,N_3580);
xnor U4984 (N_4984,N_3448,N_4373);
and U4985 (N_4985,N_3834,N_4011);
nor U4986 (N_4986,N_3643,N_4023);
nand U4987 (N_4987,N_4107,N_4362);
xor U4988 (N_4988,N_3372,N_3756);
and U4989 (N_4989,N_4057,N_3822);
and U4990 (N_4990,N_3808,N_3120);
xor U4991 (N_4991,N_3783,N_3492);
or U4992 (N_4992,N_3669,N_4265);
nor U4993 (N_4993,N_3137,N_3956);
and U4994 (N_4994,N_4193,N_4060);
nand U4995 (N_4995,N_4294,N_3857);
and U4996 (N_4996,N_3369,N_4215);
xnor U4997 (N_4997,N_4311,N_4256);
or U4998 (N_4998,N_3874,N_3546);
or U4999 (N_4999,N_4341,N_4102);
nor U5000 (N_5000,N_3076,N_3444);
and U5001 (N_5001,N_3743,N_3703);
nand U5002 (N_5002,N_4307,N_3184);
nor U5003 (N_5003,N_3793,N_3696);
nor U5004 (N_5004,N_3762,N_3466);
xnor U5005 (N_5005,N_3900,N_3182);
xor U5006 (N_5006,N_3339,N_4242);
nor U5007 (N_5007,N_3884,N_3879);
nand U5008 (N_5008,N_3263,N_4235);
and U5009 (N_5009,N_4477,N_4244);
xnor U5010 (N_5010,N_4196,N_3859);
xor U5011 (N_5011,N_3486,N_3450);
nor U5012 (N_5012,N_4009,N_4335);
and U5013 (N_5013,N_4250,N_4496);
nand U5014 (N_5014,N_3549,N_4078);
nor U5015 (N_5015,N_3771,N_4125);
nand U5016 (N_5016,N_3606,N_4222);
nand U5017 (N_5017,N_3748,N_4295);
nor U5018 (N_5018,N_4318,N_4447);
and U5019 (N_5019,N_4105,N_3028);
nand U5020 (N_5020,N_3570,N_3238);
and U5021 (N_5021,N_3715,N_4056);
nor U5022 (N_5022,N_4038,N_3090);
or U5023 (N_5023,N_3271,N_3918);
nor U5024 (N_5024,N_4012,N_3283);
nand U5025 (N_5025,N_4403,N_3760);
or U5026 (N_5026,N_3439,N_4074);
nor U5027 (N_5027,N_4349,N_3876);
or U5028 (N_5028,N_4129,N_3093);
nand U5029 (N_5029,N_4326,N_3336);
nor U5030 (N_5030,N_3973,N_4413);
or U5031 (N_5031,N_3545,N_3705);
nand U5032 (N_5032,N_3522,N_4319);
xor U5033 (N_5033,N_3735,N_3179);
nand U5034 (N_5034,N_3146,N_4433);
xor U5035 (N_5035,N_4271,N_3666);
and U5036 (N_5036,N_3284,N_3612);
or U5037 (N_5037,N_3147,N_3720);
xor U5038 (N_5038,N_4230,N_3719);
xor U5039 (N_5039,N_3931,N_3048);
nor U5040 (N_5040,N_3901,N_4151);
and U5041 (N_5041,N_3346,N_3333);
and U5042 (N_5042,N_3757,N_3096);
and U5043 (N_5043,N_3998,N_4378);
nand U5044 (N_5044,N_4336,N_3664);
nor U5045 (N_5045,N_3764,N_3867);
nor U5046 (N_5046,N_3315,N_3087);
and U5047 (N_5047,N_4453,N_4065);
nor U5048 (N_5048,N_3555,N_3889);
nand U5049 (N_5049,N_4344,N_4443);
nor U5050 (N_5050,N_3253,N_3590);
xor U5051 (N_5051,N_3716,N_4314);
xnor U5052 (N_5052,N_3579,N_3219);
nand U5053 (N_5053,N_4278,N_3306);
nor U5054 (N_5054,N_3871,N_3225);
xnor U5055 (N_5055,N_3496,N_4262);
xnor U5056 (N_5056,N_4475,N_3012);
nor U5057 (N_5057,N_3151,N_3131);
or U5058 (N_5058,N_3358,N_4414);
or U5059 (N_5059,N_4163,N_3902);
and U5060 (N_5060,N_3212,N_3230);
nand U5061 (N_5061,N_3799,N_4305);
xor U5062 (N_5062,N_4119,N_3726);
or U5063 (N_5063,N_3811,N_4304);
or U5064 (N_5064,N_4417,N_3395);
nand U5065 (N_5065,N_3787,N_3010);
nor U5066 (N_5066,N_3167,N_3068);
nand U5067 (N_5067,N_4460,N_4489);
and U5068 (N_5068,N_3183,N_4462);
xnor U5069 (N_5069,N_3127,N_3338);
xnor U5070 (N_5070,N_4337,N_3819);
or U5071 (N_5071,N_3963,N_3249);
xor U5072 (N_5072,N_3366,N_3563);
nand U5073 (N_5073,N_3955,N_4168);
and U5074 (N_5074,N_3240,N_3291);
and U5075 (N_5075,N_3195,N_3202);
xnor U5076 (N_5076,N_3401,N_4053);
or U5077 (N_5077,N_3626,N_3409);
xor U5078 (N_5078,N_4303,N_3200);
and U5079 (N_5079,N_3895,N_4313);
and U5080 (N_5080,N_3141,N_3774);
xor U5081 (N_5081,N_4217,N_4434);
nor U5082 (N_5082,N_3027,N_3203);
and U5083 (N_5083,N_3342,N_3914);
xnor U5084 (N_5084,N_4106,N_3517);
nor U5085 (N_5085,N_3776,N_3428);
nand U5086 (N_5086,N_3521,N_3582);
nor U5087 (N_5087,N_3389,N_3838);
nor U5088 (N_5088,N_4131,N_3631);
and U5089 (N_5089,N_3013,N_3217);
nand U5090 (N_5090,N_3673,N_3708);
xor U5091 (N_5091,N_3919,N_3211);
or U5092 (N_5092,N_3084,N_3873);
and U5093 (N_5093,N_3160,N_3944);
and U5094 (N_5094,N_3830,N_4364);
nand U5095 (N_5095,N_4328,N_4306);
or U5096 (N_5096,N_3210,N_3583);
nor U5097 (N_5097,N_4424,N_3856);
or U5098 (N_5098,N_4253,N_3276);
nor U5099 (N_5099,N_3694,N_3543);
nand U5100 (N_5100,N_3909,N_3758);
xnor U5101 (N_5101,N_4468,N_4449);
or U5102 (N_5102,N_3268,N_3937);
nor U5103 (N_5103,N_4401,N_3540);
nor U5104 (N_5104,N_4035,N_3725);
nor U5105 (N_5105,N_4157,N_4472);
nor U5106 (N_5106,N_3960,N_3251);
and U5107 (N_5107,N_3904,N_4441);
nor U5108 (N_5108,N_3623,N_3974);
nor U5109 (N_5109,N_4358,N_3002);
nor U5110 (N_5110,N_3118,N_3044);
and U5111 (N_5111,N_3853,N_4365);
or U5112 (N_5112,N_3198,N_3341);
nand U5113 (N_5113,N_4226,N_3119);
or U5114 (N_5114,N_3800,N_4293);
and U5115 (N_5115,N_3733,N_3564);
or U5116 (N_5116,N_3886,N_3015);
and U5117 (N_5117,N_3539,N_3231);
xor U5118 (N_5118,N_3954,N_3260);
or U5119 (N_5119,N_3484,N_4488);
and U5120 (N_5120,N_3786,N_3382);
xnor U5121 (N_5121,N_3180,N_3269);
nor U5122 (N_5122,N_3513,N_4428);
nor U5123 (N_5123,N_4096,N_3707);
or U5124 (N_5124,N_4236,N_3499);
xnor U5125 (N_5125,N_4287,N_3798);
nand U5126 (N_5126,N_3458,N_4192);
or U5127 (N_5127,N_4381,N_3929);
or U5128 (N_5128,N_3581,N_3683);
and U5129 (N_5129,N_3991,N_3296);
and U5130 (N_5130,N_3714,N_3494);
nor U5131 (N_5131,N_4159,N_3609);
nand U5132 (N_5132,N_3727,N_3535);
nand U5133 (N_5133,N_4008,N_3576);
nor U5134 (N_5134,N_3058,N_3532);
xor U5135 (N_5135,N_4426,N_3055);
nand U5136 (N_5136,N_3940,N_3588);
and U5137 (N_5137,N_3701,N_3245);
xnor U5138 (N_5138,N_3363,N_4067);
xor U5139 (N_5139,N_3110,N_3234);
or U5140 (N_5140,N_3866,N_3729);
and U5141 (N_5141,N_3326,N_4004);
nand U5142 (N_5142,N_3163,N_4272);
or U5143 (N_5143,N_3824,N_4118);
or U5144 (N_5144,N_4144,N_3047);
or U5145 (N_5145,N_3780,N_3569);
and U5146 (N_5146,N_3977,N_4040);
xor U5147 (N_5147,N_3261,N_3462);
nor U5148 (N_5148,N_3684,N_3736);
or U5149 (N_5149,N_3114,N_3759);
nand U5150 (N_5150,N_3663,N_3670);
nor U5151 (N_5151,N_3282,N_3728);
or U5152 (N_5152,N_4283,N_4243);
or U5153 (N_5153,N_3752,N_4359);
and U5154 (N_5154,N_3394,N_3408);
or U5155 (N_5155,N_3361,N_3788);
nor U5156 (N_5156,N_3656,N_3688);
nand U5157 (N_5157,N_3423,N_4084);
and U5158 (N_5158,N_3869,N_3485);
or U5159 (N_5159,N_3246,N_3413);
xor U5160 (N_5160,N_3877,N_4497);
and U5161 (N_5161,N_3585,N_3442);
nor U5162 (N_5162,N_3388,N_4325);
or U5163 (N_5163,N_3639,N_3610);
nor U5164 (N_5164,N_3406,N_3218);
and U5165 (N_5165,N_4285,N_3481);
nand U5166 (N_5166,N_3837,N_4427);
nor U5167 (N_5167,N_4174,N_3380);
nor U5168 (N_5168,N_3965,N_3193);
or U5169 (N_5169,N_4104,N_3721);
xnor U5170 (N_5170,N_4261,N_3508);
xor U5171 (N_5171,N_4388,N_3519);
nand U5172 (N_5172,N_3531,N_3236);
nor U5173 (N_5173,N_3500,N_4080);
and U5174 (N_5174,N_3706,N_3025);
nor U5175 (N_5175,N_3430,N_3171);
nor U5176 (N_5176,N_3969,N_3839);
xor U5177 (N_5177,N_3425,N_4280);
and U5178 (N_5178,N_4363,N_3153);
xor U5179 (N_5179,N_3007,N_4395);
or U5180 (N_5180,N_3319,N_4351);
xor U5181 (N_5181,N_3826,N_4245);
xor U5182 (N_5182,N_3476,N_3209);
xor U5183 (N_5183,N_3190,N_4054);
or U5184 (N_5184,N_3223,N_3575);
xnor U5185 (N_5185,N_4001,N_3530);
or U5186 (N_5186,N_3256,N_4173);
nand U5187 (N_5187,N_3385,N_3950);
nor U5188 (N_5188,N_4273,N_3544);
or U5189 (N_5189,N_3421,N_3108);
nand U5190 (N_5190,N_4366,N_3018);
or U5191 (N_5191,N_3416,N_3254);
or U5192 (N_5192,N_3680,N_4484);
nor U5193 (N_5193,N_3235,N_3674);
nor U5194 (N_5194,N_3054,N_4075);
nand U5195 (N_5195,N_3970,N_3738);
or U5196 (N_5196,N_3446,N_3651);
or U5197 (N_5197,N_4393,N_3024);
xnor U5198 (N_5198,N_3019,N_3864);
nand U5199 (N_5199,N_3672,N_4123);
and U5200 (N_5200,N_3509,N_3140);
nand U5201 (N_5201,N_4045,N_4455);
xnor U5202 (N_5202,N_3275,N_3313);
or U5203 (N_5203,N_3504,N_4367);
or U5204 (N_5204,N_4207,N_3390);
nor U5205 (N_5205,N_3329,N_4006);
nand U5206 (N_5206,N_3520,N_3906);
and U5207 (N_5207,N_4492,N_3226);
xnor U5208 (N_5208,N_3491,N_3460);
and U5209 (N_5209,N_4248,N_3964);
nand U5210 (N_5210,N_4461,N_4423);
and U5211 (N_5211,N_3667,N_4010);
or U5212 (N_5212,N_4338,N_3640);
nor U5213 (N_5213,N_4286,N_3990);
xor U5214 (N_5214,N_4410,N_3660);
or U5215 (N_5215,N_3601,N_3288);
or U5216 (N_5216,N_3083,N_3887);
xor U5217 (N_5217,N_3566,N_3215);
nand U5218 (N_5218,N_4368,N_3419);
or U5219 (N_5219,N_4206,N_3029);
nand U5220 (N_5220,N_3587,N_3497);
nand U5221 (N_5221,N_3718,N_4479);
xor U5222 (N_5222,N_3368,N_4369);
nor U5223 (N_5223,N_3490,N_4234);
xnor U5224 (N_5224,N_3224,N_3789);
and U5225 (N_5225,N_3770,N_3554);
nand U5226 (N_5226,N_3957,N_3404);
nand U5227 (N_5227,N_3835,N_3553);
xnor U5228 (N_5228,N_4155,N_3785);
or U5229 (N_5229,N_3155,N_3741);
nor U5230 (N_5230,N_4310,N_3106);
nor U5231 (N_5231,N_3092,N_4036);
nor U5232 (N_5232,N_3747,N_3300);
xor U5233 (N_5233,N_3139,N_4167);
or U5234 (N_5234,N_3525,N_3318);
or U5235 (N_5235,N_3986,N_3524);
xor U5236 (N_5236,N_3649,N_3699);
xor U5237 (N_5237,N_4392,N_3897);
nand U5238 (N_5238,N_3646,N_3661);
and U5239 (N_5239,N_3754,N_3116);
or U5240 (N_5240,N_3650,N_4418);
nor U5241 (N_5241,N_3469,N_3049);
or U5242 (N_5242,N_4408,N_4478);
nand U5243 (N_5243,N_4315,N_4019);
or U5244 (N_5244,N_4321,N_3188);
and U5245 (N_5245,N_4213,N_3259);
xnor U5246 (N_5246,N_3693,N_4289);
and U5247 (N_5247,N_3317,N_3456);
or U5248 (N_5248,N_3894,N_3732);
xor U5249 (N_5249,N_3972,N_3605);
nand U5250 (N_5250,N_3327,N_4223);
xor U5251 (N_5251,N_4451,N_3137);
and U5252 (N_5252,N_3950,N_3378);
nor U5253 (N_5253,N_3191,N_3757);
and U5254 (N_5254,N_3370,N_3997);
nand U5255 (N_5255,N_3397,N_3199);
and U5256 (N_5256,N_3183,N_3898);
nand U5257 (N_5257,N_3747,N_3633);
and U5258 (N_5258,N_4303,N_4434);
xor U5259 (N_5259,N_4051,N_4409);
and U5260 (N_5260,N_3331,N_3631);
or U5261 (N_5261,N_3927,N_3178);
or U5262 (N_5262,N_3298,N_3087);
nand U5263 (N_5263,N_3393,N_3021);
nor U5264 (N_5264,N_3113,N_4101);
xnor U5265 (N_5265,N_3104,N_3128);
or U5266 (N_5266,N_4164,N_4404);
nor U5267 (N_5267,N_3343,N_3215);
nand U5268 (N_5268,N_3723,N_3818);
xnor U5269 (N_5269,N_3754,N_4346);
and U5270 (N_5270,N_3834,N_3414);
nand U5271 (N_5271,N_4011,N_3145);
nand U5272 (N_5272,N_4134,N_3281);
nand U5273 (N_5273,N_3203,N_4435);
or U5274 (N_5274,N_3895,N_4024);
nand U5275 (N_5275,N_3456,N_3354);
nor U5276 (N_5276,N_3439,N_3339);
xor U5277 (N_5277,N_4476,N_4494);
nand U5278 (N_5278,N_3496,N_4092);
or U5279 (N_5279,N_3361,N_3329);
or U5280 (N_5280,N_4017,N_4326);
nor U5281 (N_5281,N_3949,N_3818);
and U5282 (N_5282,N_4178,N_4264);
or U5283 (N_5283,N_3898,N_3255);
nor U5284 (N_5284,N_3739,N_3201);
xnor U5285 (N_5285,N_4380,N_3414);
and U5286 (N_5286,N_4299,N_3483);
and U5287 (N_5287,N_4090,N_3952);
nor U5288 (N_5288,N_4423,N_3230);
and U5289 (N_5289,N_3391,N_3188);
nor U5290 (N_5290,N_3992,N_3073);
and U5291 (N_5291,N_3375,N_3433);
nor U5292 (N_5292,N_3916,N_4288);
and U5293 (N_5293,N_4045,N_3357);
xnor U5294 (N_5294,N_4181,N_3315);
xor U5295 (N_5295,N_3227,N_4159);
xnor U5296 (N_5296,N_3588,N_4045);
or U5297 (N_5297,N_3022,N_4109);
nor U5298 (N_5298,N_3758,N_3707);
or U5299 (N_5299,N_3316,N_4339);
nor U5300 (N_5300,N_3584,N_3730);
xor U5301 (N_5301,N_4072,N_4445);
and U5302 (N_5302,N_4295,N_4157);
xnor U5303 (N_5303,N_3424,N_4026);
xnor U5304 (N_5304,N_3578,N_3979);
nor U5305 (N_5305,N_4416,N_3860);
xnor U5306 (N_5306,N_3846,N_4173);
nor U5307 (N_5307,N_4079,N_3993);
nand U5308 (N_5308,N_4328,N_3880);
nor U5309 (N_5309,N_3034,N_3479);
nand U5310 (N_5310,N_3154,N_4119);
nand U5311 (N_5311,N_3539,N_3885);
and U5312 (N_5312,N_3802,N_3805);
nand U5313 (N_5313,N_3572,N_4334);
or U5314 (N_5314,N_3163,N_3269);
or U5315 (N_5315,N_4243,N_3092);
xnor U5316 (N_5316,N_4118,N_4297);
nand U5317 (N_5317,N_3035,N_3601);
xnor U5318 (N_5318,N_4141,N_3457);
and U5319 (N_5319,N_3249,N_4126);
nand U5320 (N_5320,N_3115,N_4157);
or U5321 (N_5321,N_3839,N_3764);
nand U5322 (N_5322,N_3208,N_3172);
xnor U5323 (N_5323,N_3287,N_3805);
or U5324 (N_5324,N_3737,N_3521);
nor U5325 (N_5325,N_3899,N_4488);
nand U5326 (N_5326,N_4414,N_4463);
xor U5327 (N_5327,N_3241,N_3119);
nor U5328 (N_5328,N_3708,N_3066);
and U5329 (N_5329,N_3859,N_3273);
xor U5330 (N_5330,N_3934,N_3947);
nor U5331 (N_5331,N_3801,N_3954);
or U5332 (N_5332,N_3457,N_3424);
nand U5333 (N_5333,N_4490,N_3367);
and U5334 (N_5334,N_3755,N_3662);
xor U5335 (N_5335,N_4270,N_4335);
nor U5336 (N_5336,N_3248,N_3000);
nand U5337 (N_5337,N_3997,N_4198);
or U5338 (N_5338,N_4458,N_3056);
nand U5339 (N_5339,N_4257,N_3948);
nor U5340 (N_5340,N_3482,N_3227);
and U5341 (N_5341,N_3278,N_4210);
nor U5342 (N_5342,N_4340,N_3661);
or U5343 (N_5343,N_3380,N_4346);
and U5344 (N_5344,N_3026,N_3928);
nor U5345 (N_5345,N_3239,N_3299);
xor U5346 (N_5346,N_3456,N_4358);
nand U5347 (N_5347,N_4142,N_3385);
xor U5348 (N_5348,N_3335,N_3050);
nor U5349 (N_5349,N_3069,N_3852);
xnor U5350 (N_5350,N_3887,N_3090);
xnor U5351 (N_5351,N_3024,N_3343);
nor U5352 (N_5352,N_4222,N_4438);
nand U5353 (N_5353,N_3260,N_3477);
and U5354 (N_5354,N_4271,N_4100);
nor U5355 (N_5355,N_3960,N_4411);
xor U5356 (N_5356,N_3512,N_3553);
nor U5357 (N_5357,N_3875,N_3395);
nor U5358 (N_5358,N_3973,N_4360);
nand U5359 (N_5359,N_3086,N_3695);
nor U5360 (N_5360,N_3018,N_4406);
nand U5361 (N_5361,N_3474,N_3040);
or U5362 (N_5362,N_3019,N_3998);
nor U5363 (N_5363,N_4432,N_3898);
and U5364 (N_5364,N_3096,N_4406);
nor U5365 (N_5365,N_3246,N_3804);
and U5366 (N_5366,N_4397,N_3012);
or U5367 (N_5367,N_4125,N_4302);
nand U5368 (N_5368,N_3026,N_3775);
nor U5369 (N_5369,N_3909,N_4217);
nor U5370 (N_5370,N_3918,N_4290);
nand U5371 (N_5371,N_3069,N_4054);
and U5372 (N_5372,N_3760,N_3332);
nand U5373 (N_5373,N_3479,N_3876);
nor U5374 (N_5374,N_4044,N_3214);
or U5375 (N_5375,N_3920,N_3646);
nor U5376 (N_5376,N_3249,N_3104);
or U5377 (N_5377,N_3903,N_4211);
or U5378 (N_5378,N_3284,N_3971);
xor U5379 (N_5379,N_3693,N_3117);
or U5380 (N_5380,N_3946,N_3467);
and U5381 (N_5381,N_4077,N_3498);
xor U5382 (N_5382,N_3556,N_3818);
or U5383 (N_5383,N_4256,N_4214);
nand U5384 (N_5384,N_4272,N_3762);
xnor U5385 (N_5385,N_3315,N_3369);
nand U5386 (N_5386,N_3648,N_3256);
xor U5387 (N_5387,N_4368,N_3484);
xnor U5388 (N_5388,N_3449,N_4385);
nand U5389 (N_5389,N_3087,N_4345);
or U5390 (N_5390,N_3858,N_3395);
nand U5391 (N_5391,N_3754,N_3506);
nand U5392 (N_5392,N_3261,N_3782);
and U5393 (N_5393,N_3097,N_4495);
xnor U5394 (N_5394,N_4091,N_4393);
xor U5395 (N_5395,N_3396,N_4084);
nand U5396 (N_5396,N_3614,N_4185);
nor U5397 (N_5397,N_3281,N_4151);
xor U5398 (N_5398,N_4222,N_3215);
or U5399 (N_5399,N_3958,N_4469);
xor U5400 (N_5400,N_3813,N_3112);
nor U5401 (N_5401,N_4230,N_4236);
and U5402 (N_5402,N_3400,N_3063);
nor U5403 (N_5403,N_3241,N_4121);
xnor U5404 (N_5404,N_3842,N_3384);
nor U5405 (N_5405,N_4151,N_3797);
nor U5406 (N_5406,N_4322,N_3266);
xnor U5407 (N_5407,N_3677,N_3679);
nor U5408 (N_5408,N_4167,N_4407);
and U5409 (N_5409,N_3757,N_3994);
nand U5410 (N_5410,N_3225,N_3083);
or U5411 (N_5411,N_3198,N_4157);
nand U5412 (N_5412,N_3050,N_4363);
nor U5413 (N_5413,N_3294,N_4349);
xnor U5414 (N_5414,N_4133,N_3795);
xor U5415 (N_5415,N_4055,N_3342);
nor U5416 (N_5416,N_3313,N_3889);
xor U5417 (N_5417,N_3834,N_4206);
or U5418 (N_5418,N_3136,N_3007);
xnor U5419 (N_5419,N_4101,N_3125);
nor U5420 (N_5420,N_3702,N_4494);
nor U5421 (N_5421,N_4160,N_3817);
or U5422 (N_5422,N_4396,N_3327);
nor U5423 (N_5423,N_3816,N_4181);
nand U5424 (N_5424,N_4487,N_4380);
and U5425 (N_5425,N_3092,N_3854);
and U5426 (N_5426,N_3672,N_3390);
nand U5427 (N_5427,N_3937,N_3575);
or U5428 (N_5428,N_4040,N_4107);
nand U5429 (N_5429,N_4397,N_3332);
nand U5430 (N_5430,N_4216,N_4024);
nand U5431 (N_5431,N_3792,N_3977);
or U5432 (N_5432,N_3570,N_3596);
nand U5433 (N_5433,N_3383,N_3096);
nor U5434 (N_5434,N_4382,N_3233);
xor U5435 (N_5435,N_3937,N_4275);
nand U5436 (N_5436,N_4098,N_3687);
xnor U5437 (N_5437,N_4457,N_3657);
xnor U5438 (N_5438,N_3693,N_3310);
or U5439 (N_5439,N_3600,N_3700);
nand U5440 (N_5440,N_3916,N_4079);
and U5441 (N_5441,N_3710,N_4057);
nor U5442 (N_5442,N_4437,N_3823);
nor U5443 (N_5443,N_3192,N_4208);
xor U5444 (N_5444,N_4013,N_4195);
nand U5445 (N_5445,N_4056,N_3322);
and U5446 (N_5446,N_3271,N_3105);
or U5447 (N_5447,N_3235,N_3572);
nor U5448 (N_5448,N_4141,N_4128);
and U5449 (N_5449,N_4097,N_3965);
nor U5450 (N_5450,N_3675,N_4487);
and U5451 (N_5451,N_3768,N_3252);
nor U5452 (N_5452,N_4266,N_3118);
and U5453 (N_5453,N_3085,N_3955);
nor U5454 (N_5454,N_3865,N_4104);
nand U5455 (N_5455,N_3387,N_3047);
and U5456 (N_5456,N_3612,N_4472);
nor U5457 (N_5457,N_4043,N_3739);
xnor U5458 (N_5458,N_4196,N_4284);
nor U5459 (N_5459,N_3715,N_3672);
nor U5460 (N_5460,N_3677,N_3141);
nor U5461 (N_5461,N_3837,N_4322);
or U5462 (N_5462,N_3465,N_3889);
nor U5463 (N_5463,N_3687,N_4485);
xor U5464 (N_5464,N_3708,N_3070);
or U5465 (N_5465,N_3675,N_3995);
nor U5466 (N_5466,N_3954,N_4427);
and U5467 (N_5467,N_4450,N_3787);
or U5468 (N_5468,N_4031,N_3079);
or U5469 (N_5469,N_3164,N_3824);
and U5470 (N_5470,N_3968,N_3723);
nor U5471 (N_5471,N_3494,N_3445);
or U5472 (N_5472,N_3387,N_4209);
or U5473 (N_5473,N_4211,N_3526);
nand U5474 (N_5474,N_3755,N_4154);
nand U5475 (N_5475,N_3499,N_4437);
nor U5476 (N_5476,N_3114,N_3705);
xnor U5477 (N_5477,N_3442,N_3048);
or U5478 (N_5478,N_3723,N_3742);
nor U5479 (N_5479,N_3523,N_4378);
xnor U5480 (N_5480,N_3803,N_4206);
or U5481 (N_5481,N_4034,N_3843);
nand U5482 (N_5482,N_4436,N_3542);
nor U5483 (N_5483,N_3263,N_4218);
and U5484 (N_5484,N_3292,N_4186);
xor U5485 (N_5485,N_3077,N_3337);
xor U5486 (N_5486,N_3894,N_4274);
and U5487 (N_5487,N_3980,N_3926);
nand U5488 (N_5488,N_3153,N_3112);
or U5489 (N_5489,N_3970,N_4138);
xor U5490 (N_5490,N_3583,N_3570);
nor U5491 (N_5491,N_3293,N_4006);
xnor U5492 (N_5492,N_3402,N_3401);
and U5493 (N_5493,N_3890,N_4216);
nand U5494 (N_5494,N_4485,N_3963);
nor U5495 (N_5495,N_3621,N_4047);
nor U5496 (N_5496,N_3018,N_4303);
nand U5497 (N_5497,N_3058,N_3934);
and U5498 (N_5498,N_4083,N_4270);
nand U5499 (N_5499,N_4125,N_4135);
xnor U5500 (N_5500,N_4445,N_3855);
nor U5501 (N_5501,N_3723,N_3792);
xor U5502 (N_5502,N_3075,N_4207);
and U5503 (N_5503,N_3410,N_3648);
nor U5504 (N_5504,N_4229,N_3240);
nand U5505 (N_5505,N_4470,N_3750);
nand U5506 (N_5506,N_3625,N_4305);
and U5507 (N_5507,N_3084,N_4472);
or U5508 (N_5508,N_4292,N_3404);
and U5509 (N_5509,N_3871,N_3779);
nor U5510 (N_5510,N_4207,N_3796);
and U5511 (N_5511,N_3048,N_3748);
or U5512 (N_5512,N_4016,N_3092);
and U5513 (N_5513,N_3149,N_3755);
and U5514 (N_5514,N_4367,N_3819);
and U5515 (N_5515,N_4270,N_3614);
xnor U5516 (N_5516,N_3072,N_4460);
nand U5517 (N_5517,N_4157,N_4179);
nor U5518 (N_5518,N_3118,N_3074);
xnor U5519 (N_5519,N_3413,N_4097);
xor U5520 (N_5520,N_4051,N_3404);
and U5521 (N_5521,N_3565,N_3876);
xor U5522 (N_5522,N_3739,N_4099);
nor U5523 (N_5523,N_3922,N_4279);
or U5524 (N_5524,N_3259,N_3922);
nand U5525 (N_5525,N_4377,N_3409);
nand U5526 (N_5526,N_4488,N_3510);
or U5527 (N_5527,N_3940,N_3854);
and U5528 (N_5528,N_3251,N_3784);
and U5529 (N_5529,N_3094,N_3961);
nor U5530 (N_5530,N_4326,N_3190);
or U5531 (N_5531,N_3798,N_3003);
and U5532 (N_5532,N_3856,N_3321);
nor U5533 (N_5533,N_4084,N_3411);
or U5534 (N_5534,N_3686,N_3312);
or U5535 (N_5535,N_3428,N_4240);
xnor U5536 (N_5536,N_3966,N_4031);
xnor U5537 (N_5537,N_4160,N_3639);
and U5538 (N_5538,N_3804,N_4237);
xnor U5539 (N_5539,N_3530,N_4377);
or U5540 (N_5540,N_4283,N_3794);
xor U5541 (N_5541,N_3105,N_3575);
nand U5542 (N_5542,N_3341,N_3474);
and U5543 (N_5543,N_3773,N_4438);
or U5544 (N_5544,N_3447,N_3634);
nand U5545 (N_5545,N_4322,N_3535);
nor U5546 (N_5546,N_3757,N_3843);
nand U5547 (N_5547,N_4397,N_3847);
or U5548 (N_5548,N_3801,N_3311);
or U5549 (N_5549,N_3503,N_4459);
nand U5550 (N_5550,N_3409,N_4208);
xor U5551 (N_5551,N_4127,N_3743);
or U5552 (N_5552,N_3562,N_3532);
and U5553 (N_5553,N_3208,N_3952);
nand U5554 (N_5554,N_3600,N_3629);
or U5555 (N_5555,N_3584,N_3366);
nand U5556 (N_5556,N_4199,N_3261);
or U5557 (N_5557,N_4347,N_3434);
nand U5558 (N_5558,N_4051,N_4010);
and U5559 (N_5559,N_3058,N_4113);
nand U5560 (N_5560,N_4476,N_4498);
xor U5561 (N_5561,N_3825,N_3643);
and U5562 (N_5562,N_3322,N_3937);
or U5563 (N_5563,N_3966,N_3071);
nor U5564 (N_5564,N_3595,N_3874);
and U5565 (N_5565,N_3348,N_3334);
and U5566 (N_5566,N_3030,N_4236);
and U5567 (N_5567,N_3366,N_3623);
and U5568 (N_5568,N_3574,N_3722);
or U5569 (N_5569,N_3992,N_3261);
nor U5570 (N_5570,N_3450,N_3564);
and U5571 (N_5571,N_3786,N_3886);
or U5572 (N_5572,N_4467,N_3781);
or U5573 (N_5573,N_4250,N_3128);
or U5574 (N_5574,N_4385,N_3174);
nand U5575 (N_5575,N_4246,N_4399);
nor U5576 (N_5576,N_3224,N_3250);
and U5577 (N_5577,N_3627,N_3544);
nand U5578 (N_5578,N_3934,N_3428);
and U5579 (N_5579,N_3023,N_3419);
nand U5580 (N_5580,N_3793,N_3742);
xor U5581 (N_5581,N_3756,N_4440);
nor U5582 (N_5582,N_3150,N_4295);
xnor U5583 (N_5583,N_4191,N_3073);
nor U5584 (N_5584,N_4400,N_3657);
or U5585 (N_5585,N_4454,N_4391);
and U5586 (N_5586,N_3954,N_3956);
nor U5587 (N_5587,N_3210,N_3393);
or U5588 (N_5588,N_4407,N_3934);
or U5589 (N_5589,N_3333,N_3825);
xor U5590 (N_5590,N_3027,N_3495);
nor U5591 (N_5591,N_3177,N_3907);
and U5592 (N_5592,N_3120,N_4119);
and U5593 (N_5593,N_3271,N_3565);
nor U5594 (N_5594,N_3388,N_3631);
or U5595 (N_5595,N_4116,N_4308);
and U5596 (N_5596,N_3924,N_3991);
nand U5597 (N_5597,N_3837,N_3591);
nand U5598 (N_5598,N_4172,N_3579);
nor U5599 (N_5599,N_3823,N_3328);
nor U5600 (N_5600,N_3660,N_3828);
nor U5601 (N_5601,N_3513,N_3486);
nor U5602 (N_5602,N_3479,N_3617);
and U5603 (N_5603,N_4124,N_3132);
and U5604 (N_5604,N_3340,N_3897);
nand U5605 (N_5605,N_3773,N_3861);
xnor U5606 (N_5606,N_4397,N_3094);
nor U5607 (N_5607,N_3310,N_4241);
xor U5608 (N_5608,N_4466,N_3488);
xnor U5609 (N_5609,N_3153,N_3874);
nor U5610 (N_5610,N_3981,N_4442);
xnor U5611 (N_5611,N_3181,N_3475);
nand U5612 (N_5612,N_4217,N_3421);
nand U5613 (N_5613,N_4233,N_3336);
nor U5614 (N_5614,N_3167,N_3318);
and U5615 (N_5615,N_3285,N_3549);
nor U5616 (N_5616,N_3882,N_3528);
or U5617 (N_5617,N_4224,N_3589);
nand U5618 (N_5618,N_3052,N_3263);
nor U5619 (N_5619,N_4125,N_3722);
nand U5620 (N_5620,N_3531,N_3984);
nand U5621 (N_5621,N_3071,N_3109);
xnor U5622 (N_5622,N_3400,N_3768);
nand U5623 (N_5623,N_3828,N_3961);
and U5624 (N_5624,N_3517,N_4382);
xnor U5625 (N_5625,N_4051,N_3427);
or U5626 (N_5626,N_4438,N_3538);
nand U5627 (N_5627,N_4084,N_4028);
or U5628 (N_5628,N_3164,N_3114);
or U5629 (N_5629,N_3754,N_4490);
or U5630 (N_5630,N_4428,N_3296);
or U5631 (N_5631,N_3124,N_3251);
xnor U5632 (N_5632,N_3322,N_3386);
or U5633 (N_5633,N_4066,N_4258);
nand U5634 (N_5634,N_3543,N_3426);
and U5635 (N_5635,N_3590,N_3939);
and U5636 (N_5636,N_4202,N_3360);
nand U5637 (N_5637,N_3011,N_3143);
nor U5638 (N_5638,N_3607,N_4089);
nor U5639 (N_5639,N_4334,N_3607);
and U5640 (N_5640,N_3816,N_4102);
nor U5641 (N_5641,N_3720,N_4144);
xor U5642 (N_5642,N_4204,N_4080);
and U5643 (N_5643,N_3262,N_3282);
and U5644 (N_5644,N_4278,N_4467);
xor U5645 (N_5645,N_4315,N_4400);
and U5646 (N_5646,N_3731,N_4434);
and U5647 (N_5647,N_4372,N_3253);
nand U5648 (N_5648,N_3029,N_3210);
or U5649 (N_5649,N_3845,N_3990);
xor U5650 (N_5650,N_4105,N_4076);
nand U5651 (N_5651,N_3077,N_4237);
nand U5652 (N_5652,N_4349,N_3698);
nor U5653 (N_5653,N_3844,N_3837);
nor U5654 (N_5654,N_3734,N_3969);
nor U5655 (N_5655,N_4276,N_4348);
nor U5656 (N_5656,N_3047,N_3395);
nor U5657 (N_5657,N_3643,N_3452);
xor U5658 (N_5658,N_4337,N_3929);
nor U5659 (N_5659,N_3678,N_4376);
nor U5660 (N_5660,N_3089,N_3995);
nand U5661 (N_5661,N_3370,N_3091);
nand U5662 (N_5662,N_3798,N_4321);
nand U5663 (N_5663,N_3282,N_4031);
nand U5664 (N_5664,N_3190,N_4286);
and U5665 (N_5665,N_3999,N_4089);
nor U5666 (N_5666,N_4218,N_3261);
xnor U5667 (N_5667,N_3980,N_3119);
or U5668 (N_5668,N_3619,N_3127);
nor U5669 (N_5669,N_4123,N_3368);
nor U5670 (N_5670,N_3428,N_4471);
nor U5671 (N_5671,N_3704,N_3347);
and U5672 (N_5672,N_4349,N_4441);
nor U5673 (N_5673,N_3731,N_4128);
nand U5674 (N_5674,N_3981,N_3221);
xnor U5675 (N_5675,N_3450,N_3312);
and U5676 (N_5676,N_4248,N_3350);
and U5677 (N_5677,N_4473,N_4315);
nand U5678 (N_5678,N_3882,N_3954);
nand U5679 (N_5679,N_3745,N_3413);
xor U5680 (N_5680,N_4376,N_4229);
xor U5681 (N_5681,N_3054,N_3402);
nand U5682 (N_5682,N_4127,N_3870);
nor U5683 (N_5683,N_4360,N_4155);
and U5684 (N_5684,N_3202,N_4389);
and U5685 (N_5685,N_4246,N_3892);
or U5686 (N_5686,N_3383,N_3218);
nand U5687 (N_5687,N_3197,N_3403);
or U5688 (N_5688,N_4254,N_3723);
and U5689 (N_5689,N_3132,N_3512);
nor U5690 (N_5690,N_3304,N_3491);
nor U5691 (N_5691,N_4093,N_4069);
and U5692 (N_5692,N_3911,N_4214);
xor U5693 (N_5693,N_3405,N_4051);
and U5694 (N_5694,N_3439,N_3370);
xor U5695 (N_5695,N_3947,N_3907);
and U5696 (N_5696,N_4488,N_3126);
or U5697 (N_5697,N_4176,N_3452);
nor U5698 (N_5698,N_4298,N_3891);
nor U5699 (N_5699,N_3560,N_3993);
and U5700 (N_5700,N_3737,N_3725);
or U5701 (N_5701,N_3544,N_3681);
nand U5702 (N_5702,N_3243,N_3713);
or U5703 (N_5703,N_4159,N_3006);
or U5704 (N_5704,N_3929,N_3935);
xor U5705 (N_5705,N_3505,N_3807);
nor U5706 (N_5706,N_4442,N_3076);
or U5707 (N_5707,N_4398,N_3182);
and U5708 (N_5708,N_4312,N_4353);
nand U5709 (N_5709,N_3458,N_3615);
xor U5710 (N_5710,N_3403,N_3957);
nor U5711 (N_5711,N_4078,N_4490);
xnor U5712 (N_5712,N_3551,N_4293);
and U5713 (N_5713,N_3490,N_3340);
and U5714 (N_5714,N_4319,N_3863);
xnor U5715 (N_5715,N_4051,N_4241);
or U5716 (N_5716,N_4119,N_3832);
nand U5717 (N_5717,N_4410,N_4289);
nand U5718 (N_5718,N_3683,N_3562);
nor U5719 (N_5719,N_3602,N_3424);
xor U5720 (N_5720,N_3496,N_3953);
nand U5721 (N_5721,N_3090,N_3151);
or U5722 (N_5722,N_3725,N_3917);
nand U5723 (N_5723,N_3518,N_4051);
nand U5724 (N_5724,N_3369,N_4471);
nand U5725 (N_5725,N_3177,N_3362);
and U5726 (N_5726,N_4046,N_3167);
nor U5727 (N_5727,N_4306,N_4287);
nand U5728 (N_5728,N_4271,N_3534);
xnor U5729 (N_5729,N_4164,N_3502);
xnor U5730 (N_5730,N_3604,N_3586);
or U5731 (N_5731,N_3667,N_3562);
nor U5732 (N_5732,N_3717,N_3627);
and U5733 (N_5733,N_4135,N_4074);
nor U5734 (N_5734,N_3863,N_3772);
xnor U5735 (N_5735,N_3105,N_4340);
nand U5736 (N_5736,N_3505,N_4222);
or U5737 (N_5737,N_3830,N_3239);
and U5738 (N_5738,N_3979,N_4482);
nor U5739 (N_5739,N_3562,N_3059);
and U5740 (N_5740,N_4148,N_4174);
and U5741 (N_5741,N_4468,N_4219);
and U5742 (N_5742,N_3324,N_3481);
xnor U5743 (N_5743,N_3408,N_3091);
and U5744 (N_5744,N_3407,N_3313);
and U5745 (N_5745,N_3366,N_3715);
and U5746 (N_5746,N_3307,N_4205);
nand U5747 (N_5747,N_4385,N_4353);
nor U5748 (N_5748,N_4193,N_3169);
and U5749 (N_5749,N_3117,N_4371);
and U5750 (N_5750,N_4464,N_3237);
nor U5751 (N_5751,N_3399,N_4226);
or U5752 (N_5752,N_3929,N_3465);
xnor U5753 (N_5753,N_3178,N_3455);
or U5754 (N_5754,N_4457,N_4086);
nand U5755 (N_5755,N_3102,N_3416);
or U5756 (N_5756,N_4191,N_3973);
and U5757 (N_5757,N_3428,N_3244);
and U5758 (N_5758,N_3008,N_4316);
or U5759 (N_5759,N_3510,N_3187);
nand U5760 (N_5760,N_4003,N_3687);
nor U5761 (N_5761,N_4040,N_3878);
nand U5762 (N_5762,N_3694,N_3348);
or U5763 (N_5763,N_4042,N_3277);
or U5764 (N_5764,N_3404,N_3895);
or U5765 (N_5765,N_3710,N_4405);
or U5766 (N_5766,N_3793,N_3247);
and U5767 (N_5767,N_3701,N_4362);
nor U5768 (N_5768,N_4243,N_3773);
nand U5769 (N_5769,N_3517,N_3079);
nor U5770 (N_5770,N_3008,N_3850);
and U5771 (N_5771,N_3834,N_4471);
and U5772 (N_5772,N_3068,N_4363);
nand U5773 (N_5773,N_3172,N_4496);
xor U5774 (N_5774,N_4005,N_3705);
xnor U5775 (N_5775,N_4321,N_3092);
or U5776 (N_5776,N_4461,N_3116);
nand U5777 (N_5777,N_4212,N_3680);
and U5778 (N_5778,N_4282,N_3134);
nand U5779 (N_5779,N_4073,N_3226);
xor U5780 (N_5780,N_4486,N_3546);
xor U5781 (N_5781,N_4087,N_3102);
nor U5782 (N_5782,N_3126,N_4421);
or U5783 (N_5783,N_3481,N_3476);
xor U5784 (N_5784,N_3518,N_3282);
and U5785 (N_5785,N_3474,N_3328);
or U5786 (N_5786,N_4010,N_3154);
or U5787 (N_5787,N_3357,N_3875);
nand U5788 (N_5788,N_3757,N_3300);
or U5789 (N_5789,N_4461,N_3885);
or U5790 (N_5790,N_3598,N_3838);
nor U5791 (N_5791,N_3268,N_4106);
nor U5792 (N_5792,N_3785,N_3392);
or U5793 (N_5793,N_3485,N_3856);
nand U5794 (N_5794,N_3983,N_4346);
and U5795 (N_5795,N_3066,N_4171);
and U5796 (N_5796,N_4170,N_3231);
nand U5797 (N_5797,N_3955,N_4054);
xor U5798 (N_5798,N_4172,N_3177);
nor U5799 (N_5799,N_3807,N_4211);
nand U5800 (N_5800,N_3397,N_3163);
nand U5801 (N_5801,N_3127,N_3446);
and U5802 (N_5802,N_3903,N_3919);
and U5803 (N_5803,N_4257,N_3638);
and U5804 (N_5804,N_3779,N_4345);
and U5805 (N_5805,N_4181,N_3102);
and U5806 (N_5806,N_3437,N_3759);
nor U5807 (N_5807,N_3094,N_4329);
xnor U5808 (N_5808,N_3133,N_3660);
and U5809 (N_5809,N_4037,N_3256);
nor U5810 (N_5810,N_3399,N_3726);
nand U5811 (N_5811,N_3745,N_3001);
or U5812 (N_5812,N_4304,N_3050);
and U5813 (N_5813,N_3813,N_3862);
nand U5814 (N_5814,N_3713,N_3640);
or U5815 (N_5815,N_4157,N_4456);
or U5816 (N_5816,N_3321,N_3133);
or U5817 (N_5817,N_4001,N_3414);
or U5818 (N_5818,N_3484,N_4147);
xnor U5819 (N_5819,N_3138,N_4012);
nor U5820 (N_5820,N_3922,N_4263);
nor U5821 (N_5821,N_3390,N_3483);
or U5822 (N_5822,N_3150,N_3694);
xnor U5823 (N_5823,N_3055,N_3425);
and U5824 (N_5824,N_4118,N_4103);
and U5825 (N_5825,N_3823,N_4469);
and U5826 (N_5826,N_3424,N_4061);
or U5827 (N_5827,N_3335,N_4146);
or U5828 (N_5828,N_3373,N_4476);
nor U5829 (N_5829,N_3728,N_4134);
or U5830 (N_5830,N_3367,N_4199);
or U5831 (N_5831,N_4281,N_3128);
or U5832 (N_5832,N_4325,N_3473);
nand U5833 (N_5833,N_3794,N_4035);
or U5834 (N_5834,N_4433,N_3023);
xnor U5835 (N_5835,N_3568,N_3178);
nand U5836 (N_5836,N_3762,N_4408);
nor U5837 (N_5837,N_4461,N_3251);
xnor U5838 (N_5838,N_3982,N_4234);
and U5839 (N_5839,N_4427,N_3073);
nor U5840 (N_5840,N_3836,N_3575);
nor U5841 (N_5841,N_3470,N_3910);
nand U5842 (N_5842,N_3535,N_4019);
nand U5843 (N_5843,N_4379,N_4158);
or U5844 (N_5844,N_3511,N_3616);
and U5845 (N_5845,N_4304,N_3747);
xor U5846 (N_5846,N_4339,N_3872);
nor U5847 (N_5847,N_3308,N_3120);
nand U5848 (N_5848,N_4347,N_3098);
xnor U5849 (N_5849,N_3721,N_3988);
nor U5850 (N_5850,N_3203,N_3535);
nor U5851 (N_5851,N_3347,N_4153);
xnor U5852 (N_5852,N_4204,N_3246);
or U5853 (N_5853,N_3410,N_3171);
xor U5854 (N_5854,N_3967,N_3399);
nand U5855 (N_5855,N_3048,N_3381);
and U5856 (N_5856,N_3208,N_3040);
xor U5857 (N_5857,N_4149,N_3055);
and U5858 (N_5858,N_3117,N_3860);
nor U5859 (N_5859,N_3119,N_4264);
nor U5860 (N_5860,N_3347,N_4040);
nor U5861 (N_5861,N_3125,N_4358);
or U5862 (N_5862,N_4253,N_3788);
nor U5863 (N_5863,N_4109,N_4191);
or U5864 (N_5864,N_3288,N_3031);
and U5865 (N_5865,N_3764,N_4377);
xor U5866 (N_5866,N_3720,N_3784);
or U5867 (N_5867,N_3133,N_3179);
and U5868 (N_5868,N_3375,N_3423);
and U5869 (N_5869,N_3793,N_4189);
and U5870 (N_5870,N_3995,N_3150);
nand U5871 (N_5871,N_4432,N_3924);
nor U5872 (N_5872,N_3950,N_3643);
nor U5873 (N_5873,N_4043,N_3214);
and U5874 (N_5874,N_4372,N_3521);
and U5875 (N_5875,N_3787,N_3209);
nor U5876 (N_5876,N_3125,N_3335);
nand U5877 (N_5877,N_4122,N_3810);
xor U5878 (N_5878,N_4049,N_3610);
xnor U5879 (N_5879,N_3507,N_3370);
or U5880 (N_5880,N_3952,N_4347);
or U5881 (N_5881,N_4019,N_3584);
or U5882 (N_5882,N_3231,N_4393);
xor U5883 (N_5883,N_4004,N_3656);
nand U5884 (N_5884,N_3362,N_3646);
and U5885 (N_5885,N_3472,N_3292);
nor U5886 (N_5886,N_3732,N_3107);
nand U5887 (N_5887,N_3832,N_3567);
and U5888 (N_5888,N_3282,N_3577);
xor U5889 (N_5889,N_4217,N_4106);
nor U5890 (N_5890,N_3875,N_3955);
or U5891 (N_5891,N_3682,N_3758);
nor U5892 (N_5892,N_3351,N_3368);
nand U5893 (N_5893,N_4059,N_4102);
and U5894 (N_5894,N_3832,N_3472);
or U5895 (N_5895,N_3924,N_3460);
nor U5896 (N_5896,N_3813,N_3349);
nand U5897 (N_5897,N_4307,N_3285);
and U5898 (N_5898,N_4115,N_4218);
and U5899 (N_5899,N_4238,N_3667);
and U5900 (N_5900,N_3537,N_4439);
or U5901 (N_5901,N_4046,N_3923);
or U5902 (N_5902,N_4228,N_4450);
xnor U5903 (N_5903,N_3056,N_3003);
nand U5904 (N_5904,N_4149,N_3800);
or U5905 (N_5905,N_3066,N_4443);
and U5906 (N_5906,N_3934,N_4488);
nor U5907 (N_5907,N_3689,N_4449);
or U5908 (N_5908,N_3866,N_3070);
and U5909 (N_5909,N_4058,N_3781);
nand U5910 (N_5910,N_3557,N_3767);
nand U5911 (N_5911,N_3954,N_3562);
and U5912 (N_5912,N_3201,N_4369);
nor U5913 (N_5913,N_3192,N_3320);
and U5914 (N_5914,N_3969,N_4123);
nor U5915 (N_5915,N_3439,N_4048);
and U5916 (N_5916,N_4189,N_4460);
and U5917 (N_5917,N_4484,N_3796);
xnor U5918 (N_5918,N_3429,N_3449);
nand U5919 (N_5919,N_3504,N_3034);
or U5920 (N_5920,N_3405,N_4389);
xnor U5921 (N_5921,N_3108,N_3105);
or U5922 (N_5922,N_3641,N_4044);
or U5923 (N_5923,N_3213,N_3879);
nand U5924 (N_5924,N_3222,N_3023);
nand U5925 (N_5925,N_3538,N_3768);
or U5926 (N_5926,N_4243,N_4443);
nand U5927 (N_5927,N_4437,N_3364);
and U5928 (N_5928,N_3540,N_3959);
nor U5929 (N_5929,N_3059,N_4254);
and U5930 (N_5930,N_3756,N_3574);
xnor U5931 (N_5931,N_4198,N_3417);
xor U5932 (N_5932,N_4303,N_4274);
nand U5933 (N_5933,N_3440,N_4135);
nand U5934 (N_5934,N_4143,N_3992);
nand U5935 (N_5935,N_3284,N_4029);
or U5936 (N_5936,N_4278,N_4394);
nand U5937 (N_5937,N_4292,N_3707);
xnor U5938 (N_5938,N_4479,N_4247);
nand U5939 (N_5939,N_4244,N_3911);
or U5940 (N_5940,N_3579,N_4456);
nor U5941 (N_5941,N_3519,N_4161);
xor U5942 (N_5942,N_3053,N_3647);
or U5943 (N_5943,N_3064,N_3736);
nand U5944 (N_5944,N_3025,N_3453);
xnor U5945 (N_5945,N_3790,N_4263);
or U5946 (N_5946,N_4410,N_3230);
nor U5947 (N_5947,N_4070,N_3996);
or U5948 (N_5948,N_4273,N_3888);
nor U5949 (N_5949,N_3787,N_3772);
nor U5950 (N_5950,N_3797,N_3139);
and U5951 (N_5951,N_3007,N_4491);
and U5952 (N_5952,N_4488,N_4199);
or U5953 (N_5953,N_3239,N_3388);
or U5954 (N_5954,N_3740,N_4147);
or U5955 (N_5955,N_3066,N_4281);
nand U5956 (N_5956,N_4055,N_3826);
or U5957 (N_5957,N_4429,N_3860);
xnor U5958 (N_5958,N_3589,N_4204);
xor U5959 (N_5959,N_4400,N_3447);
and U5960 (N_5960,N_4246,N_3666);
xnor U5961 (N_5961,N_4238,N_3281);
xnor U5962 (N_5962,N_3358,N_3940);
xor U5963 (N_5963,N_3984,N_3140);
xnor U5964 (N_5964,N_3779,N_4454);
or U5965 (N_5965,N_4207,N_3666);
and U5966 (N_5966,N_4011,N_4459);
nor U5967 (N_5967,N_3960,N_3039);
nand U5968 (N_5968,N_3440,N_3877);
and U5969 (N_5969,N_4240,N_3069);
and U5970 (N_5970,N_4492,N_4450);
nand U5971 (N_5971,N_3228,N_4314);
nand U5972 (N_5972,N_3785,N_3027);
nand U5973 (N_5973,N_3311,N_3481);
nor U5974 (N_5974,N_3393,N_3614);
nor U5975 (N_5975,N_3301,N_3120);
xnor U5976 (N_5976,N_3146,N_4434);
or U5977 (N_5977,N_4254,N_4117);
and U5978 (N_5978,N_3891,N_3094);
and U5979 (N_5979,N_4048,N_3372);
xnor U5980 (N_5980,N_4418,N_3202);
nor U5981 (N_5981,N_3732,N_3643);
xor U5982 (N_5982,N_3886,N_3873);
nand U5983 (N_5983,N_3911,N_3570);
xnor U5984 (N_5984,N_4166,N_3856);
xnor U5985 (N_5985,N_3047,N_3879);
nand U5986 (N_5986,N_4284,N_3855);
nand U5987 (N_5987,N_3411,N_4107);
xor U5988 (N_5988,N_4456,N_4324);
xor U5989 (N_5989,N_4084,N_3507);
and U5990 (N_5990,N_3897,N_4434);
or U5991 (N_5991,N_3559,N_3400);
nand U5992 (N_5992,N_3153,N_4173);
or U5993 (N_5993,N_4366,N_3096);
xnor U5994 (N_5994,N_4371,N_3472);
nand U5995 (N_5995,N_3525,N_3221);
nor U5996 (N_5996,N_4306,N_4423);
and U5997 (N_5997,N_4483,N_3935);
and U5998 (N_5998,N_3247,N_3927);
or U5999 (N_5999,N_3427,N_3115);
and U6000 (N_6000,N_5798,N_4594);
or U6001 (N_6001,N_4565,N_5501);
xor U6002 (N_6002,N_5267,N_4866);
and U6003 (N_6003,N_4836,N_5371);
nor U6004 (N_6004,N_5236,N_4981);
nand U6005 (N_6005,N_5198,N_4642);
xor U6006 (N_6006,N_5781,N_4831);
nor U6007 (N_6007,N_5191,N_4598);
nand U6008 (N_6008,N_5780,N_5278);
or U6009 (N_6009,N_5681,N_4504);
and U6010 (N_6010,N_4509,N_5183);
xor U6011 (N_6011,N_5987,N_5468);
or U6012 (N_6012,N_5339,N_4973);
or U6013 (N_6013,N_4741,N_4891);
nor U6014 (N_6014,N_5435,N_4714);
nor U6015 (N_6015,N_5715,N_4809);
and U6016 (N_6016,N_5767,N_4898);
xor U6017 (N_6017,N_5441,N_5054);
xor U6018 (N_6018,N_4656,N_4721);
nand U6019 (N_6019,N_5481,N_4757);
nand U6020 (N_6020,N_5050,N_5231);
or U6021 (N_6021,N_5943,N_5437);
or U6022 (N_6022,N_4750,N_5793);
nor U6023 (N_6023,N_5997,N_5756);
or U6024 (N_6024,N_4747,N_5065);
or U6025 (N_6025,N_5123,N_5012);
nor U6026 (N_6026,N_5227,N_4906);
or U6027 (N_6027,N_5776,N_5952);
nand U6028 (N_6028,N_5521,N_5740);
nand U6029 (N_6029,N_5090,N_5659);
nand U6030 (N_6030,N_5008,N_4698);
and U6031 (N_6031,N_5888,N_4863);
nand U6032 (N_6032,N_5608,N_5390);
xnor U6033 (N_6033,N_5306,N_5823);
nand U6034 (N_6034,N_4845,N_4812);
or U6035 (N_6035,N_5792,N_5380);
and U6036 (N_6036,N_4848,N_4502);
xnor U6037 (N_6037,N_5140,N_5408);
and U6038 (N_6038,N_4790,N_5185);
nand U6039 (N_6039,N_5735,N_5653);
nor U6040 (N_6040,N_5247,N_5121);
nor U6041 (N_6041,N_5930,N_4955);
nand U6042 (N_6042,N_5354,N_5310);
and U6043 (N_6043,N_5496,N_5901);
or U6044 (N_6044,N_5852,N_5387);
nor U6045 (N_6045,N_5162,N_4666);
nand U6046 (N_6046,N_5456,N_5016);
xnor U6047 (N_6047,N_4529,N_4507);
nor U6048 (N_6048,N_5960,N_4984);
nand U6049 (N_6049,N_5986,N_5899);
nand U6050 (N_6050,N_5818,N_5137);
and U6051 (N_6051,N_5266,N_5438);
and U6052 (N_6052,N_4618,N_5051);
xnor U6053 (N_6053,N_4725,N_4897);
xor U6054 (N_6054,N_5141,N_4534);
xnor U6055 (N_6055,N_4907,N_5196);
and U6056 (N_6056,N_4644,N_5924);
xnor U6057 (N_6057,N_5142,N_4885);
or U6058 (N_6058,N_5839,N_4899);
nor U6059 (N_6059,N_4752,N_5144);
and U6060 (N_6060,N_5499,N_4886);
and U6061 (N_6061,N_5938,N_5955);
nor U6062 (N_6062,N_4811,N_4988);
and U6063 (N_6063,N_5203,N_5993);
nor U6064 (N_6064,N_5741,N_5648);
nand U6065 (N_6065,N_5230,N_5136);
nand U6066 (N_6066,N_5394,N_5447);
nand U6067 (N_6067,N_5417,N_4832);
xor U6068 (N_6068,N_5294,N_4537);
nand U6069 (N_6069,N_5432,N_4646);
or U6070 (N_6070,N_5816,N_5106);
and U6071 (N_6071,N_5634,N_4568);
xor U6072 (N_6072,N_5353,N_5598);
xnor U6073 (N_6073,N_5133,N_4779);
or U6074 (N_6074,N_5277,N_4879);
or U6075 (N_6075,N_5836,N_4890);
or U6076 (N_6076,N_5926,N_4634);
nand U6077 (N_6077,N_5918,N_5486);
nand U6078 (N_6078,N_5972,N_5199);
and U6079 (N_6079,N_5484,N_5817);
nor U6080 (N_6080,N_5866,N_4737);
nand U6081 (N_6081,N_4630,N_5061);
or U6082 (N_6082,N_5876,N_5859);
nor U6083 (N_6083,N_5094,N_5083);
and U6084 (N_6084,N_4573,N_5594);
and U6085 (N_6085,N_5385,N_4754);
or U6086 (N_6086,N_4655,N_5596);
or U6087 (N_6087,N_5743,N_4658);
nor U6088 (N_6088,N_4579,N_5957);
xor U6089 (N_6089,N_4830,N_5244);
xor U6090 (N_6090,N_5341,N_5936);
xor U6091 (N_6091,N_5245,N_5873);
xnor U6092 (N_6092,N_5082,N_4728);
and U6093 (N_6093,N_5639,N_5105);
nand U6094 (N_6094,N_4603,N_5810);
xor U6095 (N_6095,N_5584,N_5988);
xor U6096 (N_6096,N_5014,N_4970);
nor U6097 (N_6097,N_5188,N_5098);
nor U6098 (N_6098,N_4956,N_5223);
nor U6099 (N_6099,N_4787,N_5066);
nand U6100 (N_6100,N_5386,N_5512);
or U6101 (N_6101,N_4690,N_5580);
nor U6102 (N_6102,N_5265,N_5835);
nor U6103 (N_6103,N_5604,N_5612);
nand U6104 (N_6104,N_5044,N_5749);
or U6105 (N_6105,N_5329,N_5643);
nand U6106 (N_6106,N_5931,N_5379);
nor U6107 (N_6107,N_4510,N_5115);
and U6108 (N_6108,N_4678,N_4635);
nor U6109 (N_6109,N_4806,N_5109);
or U6110 (N_6110,N_4540,N_4519);
nand U6111 (N_6111,N_5312,N_4841);
nand U6112 (N_6112,N_5732,N_4616);
nor U6113 (N_6113,N_5449,N_4993);
or U6114 (N_6114,N_5164,N_5268);
nor U6115 (N_6115,N_5007,N_5728);
nand U6116 (N_6116,N_5346,N_4872);
and U6117 (N_6117,N_5998,N_5440);
nor U6118 (N_6118,N_5210,N_5791);
and U6119 (N_6119,N_5625,N_4976);
nor U6120 (N_6120,N_5976,N_5959);
or U6121 (N_6121,N_5912,N_4539);
xor U6122 (N_6122,N_5962,N_4778);
or U6123 (N_6123,N_5610,N_4992);
and U6124 (N_6124,N_5577,N_4566);
or U6125 (N_6125,N_5365,N_4758);
and U6126 (N_6126,N_4919,N_5886);
nand U6127 (N_6127,N_5645,N_5261);
xor U6128 (N_6128,N_5779,N_4917);
nor U6129 (N_6129,N_5338,N_4876);
xnor U6130 (N_6130,N_5434,N_5360);
nor U6131 (N_6131,N_5614,N_5323);
or U6132 (N_6132,N_5139,N_5273);
or U6133 (N_6133,N_5337,N_4915);
and U6134 (N_6134,N_5286,N_4952);
xnor U6135 (N_6135,N_5946,N_5799);
or U6136 (N_6136,N_5590,N_5970);
nand U6137 (N_6137,N_4523,N_5472);
or U6138 (N_6138,N_5631,N_5152);
nor U6139 (N_6139,N_5678,N_5842);
and U6140 (N_6140,N_4705,N_5975);
or U6141 (N_6141,N_4559,N_4774);
or U6142 (N_6142,N_5856,N_5797);
nand U6143 (N_6143,N_5118,N_5522);
nor U6144 (N_6144,N_5724,N_5455);
and U6145 (N_6145,N_4798,N_5956);
nor U6146 (N_6146,N_5321,N_5126);
or U6147 (N_6147,N_5689,N_5576);
nor U6148 (N_6148,N_4718,N_4662);
nand U6149 (N_6149,N_5308,N_5197);
xnor U6150 (N_6150,N_4934,N_5655);
nand U6151 (N_6151,N_5696,N_5705);
or U6152 (N_6152,N_5361,N_5350);
nand U6153 (N_6153,N_5285,N_5507);
and U6154 (N_6154,N_5815,N_5745);
or U6155 (N_6155,N_4985,N_4800);
nor U6156 (N_6156,N_5863,N_5181);
nand U6157 (N_6157,N_5347,N_5651);
nor U6158 (N_6158,N_4726,N_5738);
nor U6159 (N_6159,N_4614,N_5914);
or U6160 (N_6160,N_5463,N_4517);
nor U6161 (N_6161,N_5465,N_5964);
nor U6162 (N_6162,N_5257,N_4914);
xor U6163 (N_6163,N_5910,N_5155);
nor U6164 (N_6164,N_5695,N_5896);
xnor U6165 (N_6165,N_4556,N_5707);
or U6166 (N_6166,N_5450,N_4949);
and U6167 (N_6167,N_5958,N_4749);
xnor U6168 (N_6168,N_5733,N_4677);
nor U6169 (N_6169,N_4768,N_4802);
and U6170 (N_6170,N_5567,N_4561);
nand U6171 (N_6171,N_5748,N_4609);
or U6172 (N_6172,N_5649,N_4613);
nand U6173 (N_6173,N_5771,N_5553);
and U6174 (N_6174,N_5058,N_5420);
and U6175 (N_6175,N_5328,N_5027);
nand U6176 (N_6176,N_5990,N_5628);
xnor U6177 (N_6177,N_5404,N_5263);
nor U6178 (N_6178,N_5744,N_5889);
nand U6179 (N_6179,N_5364,N_5550);
xor U6180 (N_6180,N_5828,N_5428);
xnor U6181 (N_6181,N_5934,N_5063);
or U6182 (N_6182,N_4834,N_5949);
xnor U6183 (N_6183,N_4659,N_5047);
and U6184 (N_6184,N_5848,N_5737);
nand U6185 (N_6185,N_5518,N_5693);
nand U6186 (N_6186,N_4815,N_5974);
xnor U6187 (N_6187,N_4982,N_5951);
or U6188 (N_6188,N_5723,N_4818);
nand U6189 (N_6189,N_4829,N_5304);
nand U6190 (N_6190,N_4796,N_5963);
or U6191 (N_6191,N_5813,N_5478);
and U6192 (N_6192,N_4505,N_5332);
nor U6193 (N_6193,N_5857,N_4626);
or U6194 (N_6194,N_5146,N_5297);
and U6195 (N_6195,N_5769,N_4580);
xor U6196 (N_6196,N_4944,N_5929);
nor U6197 (N_6197,N_5362,N_4680);
and U6198 (N_6198,N_4777,N_5143);
nor U6199 (N_6199,N_5887,N_5103);
nand U6200 (N_6200,N_5851,N_5671);
and U6201 (N_6201,N_4954,N_4637);
nand U6202 (N_6202,N_4974,N_5709);
and U6203 (N_6203,N_4686,N_5833);
xor U6204 (N_6204,N_4627,N_5497);
or U6205 (N_6205,N_5629,N_5225);
or U6206 (N_6206,N_5582,N_4661);
and U6207 (N_6207,N_5333,N_5630);
xnor U6208 (N_6208,N_5205,N_5099);
xor U6209 (N_6209,N_5416,N_5461);
nor U6210 (N_6210,N_5270,N_4625);
and U6211 (N_6211,N_5831,N_5832);
xor U6212 (N_6212,N_5402,N_5241);
nand U6213 (N_6213,N_5274,N_5454);
nor U6214 (N_6214,N_4695,N_4895);
nor U6215 (N_6215,N_5878,N_5057);
nor U6216 (N_6216,N_5091,N_5357);
or U6217 (N_6217,N_4512,N_5754);
nand U6218 (N_6218,N_5819,N_5571);
or U6219 (N_6219,N_5664,N_5683);
nor U6220 (N_6220,N_4732,N_5513);
or U6221 (N_6221,N_5822,N_4582);
nand U6222 (N_6222,N_4665,N_5947);
nand U6223 (N_6223,N_4918,N_5840);
or U6224 (N_6224,N_5165,N_5814);
xnor U6225 (N_6225,N_5107,N_5445);
nand U6226 (N_6226,N_4583,N_5037);
nor U6227 (N_6227,N_5690,N_4847);
nand U6228 (N_6228,N_4735,N_4927);
nor U6229 (N_6229,N_4912,N_5812);
or U6230 (N_6230,N_4590,N_5657);
and U6231 (N_6231,N_5429,N_5159);
and U6232 (N_6232,N_5158,N_5838);
xor U6233 (N_6233,N_4986,N_5149);
nor U6234 (N_6234,N_5564,N_5971);
nor U6235 (N_6235,N_4727,N_5384);
or U6236 (N_6236,N_5853,N_4837);
and U6237 (N_6237,N_4654,N_4544);
or U6238 (N_6238,N_4854,N_4513);
nor U6239 (N_6239,N_4522,N_5932);
nand U6240 (N_6240,N_4615,N_5560);
xor U6241 (N_6241,N_4980,N_5234);
or U6242 (N_6242,N_5295,N_4861);
or U6243 (N_6243,N_5593,N_5556);
nand U6244 (N_6244,N_5829,N_4780);
and U6245 (N_6245,N_5427,N_5194);
and U6246 (N_6246,N_4803,N_4763);
nor U6247 (N_6247,N_5633,N_4596);
and U6248 (N_6248,N_4549,N_5334);
nor U6249 (N_6249,N_5568,N_4547);
and U6250 (N_6250,N_4821,N_4884);
and U6251 (N_6251,N_5232,N_4610);
xor U6252 (N_6252,N_5006,N_5296);
xor U6253 (N_6253,N_5130,N_5498);
xnor U6254 (N_6254,N_5868,N_5788);
and U6255 (N_6255,N_5279,N_5087);
and U6256 (N_6256,N_4515,N_4572);
or U6257 (N_6257,N_4853,N_4764);
nand U6258 (N_6258,N_4524,N_5336);
or U6259 (N_6259,N_4586,N_5423);
nand U6260 (N_6260,N_4875,N_5011);
and U6261 (N_6261,N_5999,N_4971);
nand U6262 (N_6262,N_4520,N_5714);
or U6263 (N_6263,N_4676,N_4870);
nand U6264 (N_6264,N_4570,N_5457);
nor U6265 (N_6265,N_5311,N_5370);
nand U6266 (N_6266,N_5401,N_5944);
nor U6267 (N_6267,N_4553,N_5881);
and U6268 (N_6268,N_5022,N_4855);
nor U6269 (N_6269,N_4647,N_5026);
xnor U6270 (N_6270,N_5249,N_5563);
nor U6271 (N_6271,N_5376,N_5581);
xor U6272 (N_6272,N_5706,N_5076);
or U6273 (N_6273,N_4894,N_5674);
and U6274 (N_6274,N_4938,N_4604);
and U6275 (N_6275,N_5056,N_4704);
nand U6276 (N_6276,N_5613,N_4643);
and U6277 (N_6277,N_4781,N_5509);
nand U6278 (N_6278,N_4801,N_5699);
xor U6279 (N_6279,N_5623,N_5064);
xor U6280 (N_6280,N_5669,N_5355);
and U6281 (N_6281,N_5351,N_5684);
xor U6282 (N_6282,N_5204,N_5504);
xor U6283 (N_6283,N_5945,N_5915);
nor U6284 (N_6284,N_5757,N_5182);
xnor U6285 (N_6285,N_5795,N_5908);
xnor U6286 (N_6286,N_5948,N_5460);
or U6287 (N_6287,N_4692,N_5555);
and U6288 (N_6288,N_5212,N_5487);
nand U6289 (N_6289,N_5451,N_5073);
nand U6290 (N_6290,N_4833,N_4810);
or U6291 (N_6291,N_4587,N_5403);
nor U6292 (N_6292,N_5395,N_4900);
nand U6293 (N_6293,N_4733,N_5624);
and U6294 (N_6294,N_5692,N_4593);
and U6295 (N_6295,N_5117,N_5597);
xor U6296 (N_6296,N_5092,N_5535);
xnor U6297 (N_6297,N_5900,N_5884);
xnor U6298 (N_6298,N_5045,N_5586);
and U6299 (N_6299,N_5532,N_5890);
xnor U6300 (N_6300,N_5825,N_5519);
xnor U6301 (N_6301,N_5869,N_5175);
nor U6302 (N_6302,N_5939,N_4925);
nor U6303 (N_6303,N_5207,N_4827);
xnor U6304 (N_6304,N_4709,N_4712);
and U6305 (N_6305,N_5129,N_5281);
xnor U6306 (N_6306,N_4964,N_4959);
and U6307 (N_6307,N_5178,N_5009);
nand U6308 (N_6308,N_4730,N_5222);
nor U6309 (N_6309,N_4857,N_5324);
and U6310 (N_6310,N_4632,N_4702);
and U6311 (N_6311,N_5790,N_4995);
nor U6312 (N_6312,N_5870,N_5415);
and U6313 (N_6313,N_4877,N_5067);
or U6314 (N_6314,N_5242,N_4935);
nand U6315 (N_6315,N_4669,N_5966);
or U6316 (N_6316,N_4904,N_4710);
xor U6317 (N_6317,N_5722,N_5545);
or U6318 (N_6318,N_5768,N_5761);
or U6319 (N_6319,N_4922,N_5994);
nand U6320 (N_6320,N_5661,N_5516);
nor U6321 (N_6321,N_5784,N_4706);
nand U6322 (N_6322,N_4667,N_5941);
nand U6323 (N_6323,N_5485,N_4765);
xnor U6324 (N_6324,N_5475,N_5985);
nand U6325 (N_6325,N_5796,N_5293);
nand U6326 (N_6326,N_4849,N_5736);
nand U6327 (N_6327,N_5902,N_5200);
nor U6328 (N_6328,N_4628,N_5700);
nor U6329 (N_6329,N_5820,N_5770);
xnor U6330 (N_6330,N_5031,N_5954);
and U6331 (N_6331,N_4941,N_5824);
and U6332 (N_6332,N_5766,N_5138);
nand U6333 (N_6333,N_5837,N_4672);
or U6334 (N_6334,N_5538,N_5973);
nand U6335 (N_6335,N_5500,N_4543);
nand U6336 (N_6336,N_5157,N_5359);
nor U6337 (N_6337,N_5883,N_5526);
and U6338 (N_6338,N_5760,N_5844);
nand U6339 (N_6339,N_5208,N_4951);
and U6340 (N_6340,N_5601,N_4612);
nor U6341 (N_6341,N_5302,N_5179);
and U6342 (N_6342,N_5697,N_4567);
and U6343 (N_6343,N_5148,N_4864);
xnor U6344 (N_6344,N_4932,N_5569);
nor U6345 (N_6345,N_5081,N_5453);
or U6346 (N_6346,N_5119,N_5032);
and U6347 (N_6347,N_5272,N_5524);
and U6348 (N_6348,N_5885,N_5980);
and U6349 (N_6349,N_5043,N_4557);
and U6350 (N_6350,N_5309,N_5239);
or U6351 (N_6351,N_5366,N_5575);
and U6352 (N_6352,N_4681,N_4761);
nor U6353 (N_6353,N_4550,N_4916);
nor U6354 (N_6354,N_5174,N_4697);
nor U6355 (N_6355,N_5235,N_5573);
xnor U6356 (N_6356,N_5611,N_5599);
or U6357 (N_6357,N_5950,N_5762);
or U6358 (N_6358,N_5953,N_5382);
nor U6359 (N_6359,N_5187,N_5214);
and U6360 (N_6360,N_5551,N_4622);
xnor U6361 (N_6361,N_5080,N_4893);
nor U6362 (N_6362,N_5202,N_5284);
nor U6363 (N_6363,N_5635,N_4953);
or U6364 (N_6364,N_5477,N_4688);
and U6365 (N_6365,N_5619,N_5292);
xnor U6366 (N_6366,N_5656,N_4511);
and U6367 (N_6367,N_5493,N_4624);
and U6368 (N_6368,N_4660,N_4648);
or U6369 (N_6369,N_5755,N_4571);
or U6370 (N_6370,N_5246,N_5372);
nor U6371 (N_6371,N_5120,N_5746);
xor U6372 (N_6372,N_5846,N_5414);
and U6373 (N_6373,N_5991,N_5112);
and U6374 (N_6374,N_5774,N_5909);
and U6375 (N_6375,N_5411,N_4723);
xor U6376 (N_6376,N_4668,N_4651);
and U6377 (N_6377,N_4736,N_5882);
or U6378 (N_6378,N_5880,N_5226);
or U6379 (N_6379,N_4751,N_5340);
and U6380 (N_6380,N_4923,N_4880);
nor U6381 (N_6381,N_4942,N_5548);
or U6382 (N_6382,N_5010,N_5928);
xnor U6383 (N_6383,N_4564,N_4850);
and U6384 (N_6384,N_5794,N_5036);
or U6385 (N_6385,N_5969,N_5430);
nor U6386 (N_6386,N_4928,N_4860);
xor U6387 (N_6387,N_5125,N_5271);
and U6388 (N_6388,N_5872,N_5255);
nor U6389 (N_6389,N_4687,N_4773);
xnor U6390 (N_6390,N_4595,N_4805);
nand U6391 (N_6391,N_5343,N_5905);
nor U6392 (N_6392,N_5084,N_5666);
and U6393 (N_6393,N_4584,N_4972);
and U6394 (N_6394,N_5543,N_4722);
nor U6395 (N_6395,N_5480,N_5326);
nand U6396 (N_6396,N_5269,N_4936);
nand U6397 (N_6397,N_5074,N_5708);
nor U6398 (N_6398,N_5436,N_4776);
xnor U6399 (N_6399,N_5618,N_5570);
nand U6400 (N_6400,N_4852,N_5458);
nand U6401 (N_6401,N_4783,N_4913);
xor U6402 (N_6402,N_5685,N_5217);
or U6403 (N_6403,N_5965,N_5248);
or U6404 (N_6404,N_5718,N_5483);
xor U6405 (N_6405,N_5237,N_5055);
and U6406 (N_6406,N_4978,N_4620);
nand U6407 (N_6407,N_4611,N_5879);
or U6408 (N_6408,N_4716,N_4910);
xnor U6409 (N_6409,N_5342,N_4530);
xnor U6410 (N_6410,N_4943,N_5153);
nand U6411 (N_6411,N_5005,N_5919);
and U6412 (N_6412,N_5114,N_5062);
xor U6413 (N_6413,N_5785,N_4623);
xor U6414 (N_6414,N_5029,N_5373);
nand U6415 (N_6415,N_5001,N_4926);
nand U6416 (N_6416,N_4558,N_5989);
or U6417 (N_6417,N_5804,N_5190);
nand U6418 (N_6418,N_5800,N_4858);
nor U6419 (N_6419,N_4674,N_5775);
nand U6420 (N_6420,N_4889,N_4696);
or U6421 (N_6421,N_4629,N_4711);
xor U6422 (N_6422,N_5168,N_5156);
or U6423 (N_6423,N_4742,N_4619);
xnor U6424 (N_6424,N_5982,N_5020);
and U6425 (N_6425,N_5942,N_5034);
xnor U6426 (N_6426,N_4921,N_5917);
xnor U6427 (N_6427,N_5452,N_5977);
nor U6428 (N_6428,N_4794,N_5579);
and U6429 (N_6429,N_4685,N_4621);
xnor U6430 (N_6430,N_4767,N_5801);
xor U6431 (N_6431,N_4844,N_5777);
nor U6432 (N_6432,N_5617,N_5508);
or U6433 (N_6433,N_4948,N_5894);
or U6434 (N_6434,N_4961,N_5712);
nand U6435 (N_6435,N_5327,N_5898);
nor U6436 (N_6436,N_5320,N_5469);
nand U6437 (N_6437,N_5996,N_4684);
and U6438 (N_6438,N_5542,N_4693);
xnor U6439 (N_6439,N_4592,N_5782);
nand U6440 (N_6440,N_4528,N_4631);
nand U6441 (N_6441,N_5251,N_4527);
and U6442 (N_6442,N_4975,N_5252);
or U6443 (N_6443,N_4939,N_4552);
nand U6444 (N_6444,N_5565,N_4526);
or U6445 (N_6445,N_5368,N_5363);
xnor U6446 (N_6446,N_5215,N_4835);
or U6447 (N_6447,N_5116,N_5462);
xor U6448 (N_6448,N_4645,N_5253);
or U6449 (N_6449,N_5721,N_5688);
nand U6450 (N_6450,N_4786,N_5393);
nor U6451 (N_6451,N_5053,N_5135);
and U6452 (N_6452,N_5730,N_5433);
and U6453 (N_6453,N_5670,N_5559);
nand U6454 (N_6454,N_4569,N_5161);
and U6455 (N_6455,N_4892,N_4541);
nand U6456 (N_6456,N_5444,N_5169);
xor U6457 (N_6457,N_5515,N_5626);
and U6458 (N_6458,N_5672,N_4599);
and U6459 (N_6459,N_5425,N_4820);
nand U6460 (N_6460,N_5547,N_5392);
or U6461 (N_6461,N_5218,N_4968);
nor U6462 (N_6462,N_5086,N_4508);
xnor U6463 (N_6463,N_4881,N_5163);
nand U6464 (N_6464,N_4775,N_5046);
nor U6465 (N_6465,N_5419,N_4597);
or U6466 (N_6466,N_5821,N_5038);
or U6467 (N_6467,N_4856,N_5102);
nor U6468 (N_6468,N_4760,N_5520);
or U6469 (N_6469,N_4542,N_5002);
nand U6470 (N_6470,N_5124,N_4503);
nand U6471 (N_6471,N_5319,N_4514);
and U6472 (N_6472,N_4911,N_5422);
xnor U6473 (N_6473,N_5206,N_5077);
nor U6474 (N_6474,N_5752,N_5984);
nor U6475 (N_6475,N_5510,N_5763);
and U6476 (N_6476,N_5147,N_5479);
xnor U6477 (N_6477,N_5529,N_5834);
nand U6478 (N_6478,N_4882,N_5916);
nand U6479 (N_6479,N_5622,N_5476);
or U6480 (N_6480,N_5827,N_5621);
xnor U6481 (N_6481,N_4675,N_5154);
and U6482 (N_6482,N_5644,N_5561);
xnor U6483 (N_6483,N_5867,N_5330);
xor U6484 (N_6484,N_5167,N_4538);
or U6485 (N_6485,N_5258,N_5111);
and U6486 (N_6486,N_4873,N_5861);
xnor U6487 (N_6487,N_5687,N_4762);
nand U6488 (N_6488,N_5727,N_5276);
nor U6489 (N_6489,N_5742,N_5747);
and U6490 (N_6490,N_5667,N_5467);
nor U6491 (N_6491,N_4924,N_5676);
xnor U6492 (N_6492,N_4772,N_5325);
nor U6493 (N_6493,N_5374,N_5021);
nor U6494 (N_6494,N_5132,N_5787);
and U6495 (N_6495,N_4851,N_4753);
nor U6496 (N_6496,N_5189,N_4724);
and U6497 (N_6497,N_5603,N_5017);
nand U6498 (N_6498,N_5783,N_5826);
xnor U6499 (N_6499,N_5716,N_5079);
nor U6500 (N_6500,N_4983,N_5530);
nor U6501 (N_6501,N_5717,N_4962);
and U6502 (N_6502,N_5446,N_5961);
nand U6503 (N_6503,N_4525,N_5862);
nor U6504 (N_6504,N_5220,N_5940);
or U6505 (N_6505,N_5317,N_4846);
and U6506 (N_6506,N_4531,N_5698);
nor U6507 (N_6507,N_4591,N_5367);
nor U6508 (N_6508,N_5398,N_5151);
nor U6509 (N_6509,N_5874,N_5041);
nand U6510 (N_6510,N_5410,N_4825);
nor U6511 (N_6511,N_4969,N_5171);
nor U6512 (N_6512,N_5809,N_5595);
nand U6513 (N_6513,N_5421,N_4990);
nor U6514 (N_6514,N_4769,N_5211);
xnor U6515 (N_6515,N_4713,N_5316);
or U6516 (N_6516,N_5280,N_5806);
or U6517 (N_6517,N_4694,N_4766);
or U6518 (N_6518,N_4554,N_5383);
nand U6519 (N_6519,N_5647,N_5283);
nand U6520 (N_6520,N_5654,N_5170);
and U6521 (N_6521,N_5979,N_5525);
nand U6522 (N_6522,N_5701,N_5391);
nand U6523 (N_6523,N_5734,N_5558);
or U6524 (N_6524,N_4731,N_5589);
or U6525 (N_6525,N_4920,N_5843);
or U6526 (N_6526,N_4791,N_5301);
or U6527 (N_6527,N_4828,N_4516);
xor U6528 (N_6528,N_4822,N_4867);
xor U6529 (N_6529,N_4608,N_5591);
nor U6530 (N_6530,N_4967,N_5907);
nor U6531 (N_6531,N_5702,N_4789);
nand U6532 (N_6532,N_5290,N_5620);
nor U6533 (N_6533,N_5131,N_5865);
nor U6534 (N_6534,N_4548,N_5933);
nor U6535 (N_6535,N_5369,N_5850);
nand U6536 (N_6536,N_5682,N_4797);
nor U6537 (N_6537,N_5491,N_5668);
and U6538 (N_6538,N_5042,N_5562);
nor U6539 (N_6539,N_4602,N_5331);
nor U6540 (N_6540,N_5243,N_5895);
xor U6541 (N_6541,N_5920,N_5075);
and U6542 (N_6542,N_5259,N_4551);
nor U6543 (N_6543,N_5642,N_5413);
nand U6544 (N_6544,N_5640,N_4808);
nand U6545 (N_6545,N_4689,N_5922);
or U6546 (N_6546,N_4720,N_5068);
nand U6547 (N_6547,N_5514,N_5786);
nand U6548 (N_6548,N_5023,N_5602);
xnor U6549 (N_6549,N_5015,N_5470);
xnor U6550 (N_6550,N_5399,N_4997);
nor U6551 (N_6551,N_5765,N_4795);
and U6552 (N_6552,N_5572,N_4719);
and U6553 (N_6553,N_4999,N_4909);
xnor U6554 (N_6554,N_5240,N_5720);
and U6555 (N_6555,N_5228,N_5679);
and U6556 (N_6556,N_4649,N_5096);
nand U6557 (N_6557,N_5172,N_4929);
nor U6558 (N_6558,N_5632,N_5592);
and U6559 (N_6559,N_5811,N_5110);
and U6560 (N_6560,N_5505,N_5400);
xor U6561 (N_6561,N_5923,N_5305);
nor U6562 (N_6562,N_5160,N_5566);
nor U6563 (N_6563,N_4826,N_5059);
xor U6564 (N_6564,N_5303,N_5442);
or U6565 (N_6565,N_4729,N_4843);
nand U6566 (N_6566,N_4759,N_5726);
and U6567 (N_6567,N_5300,N_4842);
nand U6568 (N_6568,N_4940,N_5650);
or U6569 (N_6569,N_5322,N_4883);
or U6570 (N_6570,N_5877,N_5431);
and U6571 (N_6571,N_4500,N_5967);
nor U6572 (N_6572,N_4606,N_5534);
nand U6573 (N_6573,N_5638,N_5180);
nor U6574 (N_6574,N_5019,N_4521);
xnor U6575 (N_6575,N_5049,N_4600);
nand U6576 (N_6576,N_4585,N_5615);
nor U6577 (N_6577,N_5256,N_5546);
nand U6578 (N_6578,N_5855,N_5318);
nor U6579 (N_6579,N_5927,N_4601);
xnor U6580 (N_6580,N_5492,N_4535);
xor U6581 (N_6581,N_5348,N_4588);
and U6582 (N_6582,N_5177,N_4862);
and U6583 (N_6583,N_4734,N_4717);
nand U6584 (N_6584,N_5983,N_4977);
or U6585 (N_6585,N_5443,N_4744);
nor U6586 (N_6586,N_4533,N_5166);
or U6587 (N_6587,N_5195,N_4638);
nor U6588 (N_6588,N_5201,N_5751);
xor U6589 (N_6589,N_5527,N_5627);
or U6590 (N_6590,N_4931,N_4640);
xor U6591 (N_6591,N_5471,N_5725);
or U6592 (N_6592,N_5407,N_4998);
and U6593 (N_6593,N_4743,N_4819);
nand U6594 (N_6594,N_4578,N_4868);
xnor U6595 (N_6595,N_4958,N_4657);
or U6596 (N_6596,N_4589,N_5101);
xor U6597 (N_6597,N_4946,N_4902);
xnor U6598 (N_6598,N_5352,N_4546);
nand U6599 (N_6599,N_4560,N_5052);
xnor U6600 (N_6600,N_5803,N_5464);
and U6601 (N_6601,N_5636,N_5375);
nor U6602 (N_6602,N_4930,N_4671);
or U6603 (N_6603,N_4740,N_5511);
or U6604 (N_6604,N_5925,N_5652);
or U6605 (N_6605,N_5864,N_5490);
nand U6606 (N_6606,N_4605,N_5097);
and U6607 (N_6607,N_5426,N_4607);
nand U6608 (N_6608,N_5719,N_5104);
nand U6609 (N_6609,N_5313,N_5221);
nand U6610 (N_6610,N_4903,N_5291);
nand U6611 (N_6611,N_4545,N_4908);
nand U6612 (N_6612,N_4838,N_5128);
xnor U6613 (N_6613,N_4699,N_4670);
and U6614 (N_6614,N_5531,N_5607);
xor U6615 (N_6615,N_5127,N_4673);
nand U6616 (N_6616,N_5078,N_4788);
and U6617 (N_6617,N_5184,N_5517);
nand U6618 (N_6618,N_5897,N_5409);
nand U6619 (N_6619,N_5854,N_4865);
or U6620 (N_6620,N_4784,N_5466);
xnor U6621 (N_6621,N_4664,N_5287);
xor U6622 (N_6622,N_4577,N_5663);
xor U6623 (N_6623,N_5921,N_5802);
or U6624 (N_6624,N_4633,N_4816);
xnor U6625 (N_6625,N_5298,N_5254);
nor U6626 (N_6626,N_4707,N_5024);
xnor U6627 (N_6627,N_5913,N_4701);
nor U6628 (N_6628,N_5000,N_5229);
or U6629 (N_6629,N_4869,N_4799);
and U6630 (N_6630,N_4663,N_5003);
nor U6631 (N_6631,N_4979,N_4653);
nand U6632 (N_6632,N_5750,N_5040);
nor U6633 (N_6633,N_4965,N_4814);
nand U6634 (N_6634,N_5871,N_4874);
nand U6635 (N_6635,N_5892,N_5315);
or U6636 (N_6636,N_5377,N_5694);
or U6637 (N_6637,N_4682,N_5176);
and U6638 (N_6638,N_5388,N_4896);
nand U6639 (N_6639,N_5405,N_5544);
and U6640 (N_6640,N_5753,N_4945);
xnor U6641 (N_6641,N_5406,N_4991);
nand U6642 (N_6642,N_5397,N_4650);
or U6643 (N_6643,N_4994,N_5418);
nand U6644 (N_6644,N_5713,N_5122);
nand U6645 (N_6645,N_4840,N_5906);
nand U6646 (N_6646,N_5903,N_4888);
or U6647 (N_6647,N_5739,N_5841);
and U6648 (N_6648,N_4782,N_5904);
and U6649 (N_6649,N_5540,N_5070);
and U6650 (N_6650,N_5473,N_5968);
and U6651 (N_6651,N_5554,N_5396);
xor U6652 (N_6652,N_5665,N_5072);
or U6653 (N_6653,N_5609,N_5299);
and U6654 (N_6654,N_5808,N_5060);
nor U6655 (N_6655,N_5759,N_4745);
nand U6656 (N_6656,N_4950,N_5646);
nor U6657 (N_6657,N_4617,N_5549);
nor U6658 (N_6658,N_5209,N_4804);
nor U6659 (N_6659,N_5893,N_4807);
and U6660 (N_6660,N_5587,N_4989);
nor U6661 (N_6661,N_4996,N_4963);
nand U6662 (N_6662,N_5028,N_5219);
or U6663 (N_6663,N_5710,N_4652);
or U6664 (N_6664,N_5093,N_5807);
xnor U6665 (N_6665,N_5704,N_5606);
xnor U6666 (N_6666,N_5100,N_4933);
and U6667 (N_6667,N_5088,N_5213);
nand U6668 (N_6668,N_4823,N_4746);
or U6669 (N_6669,N_5145,N_4839);
or U6670 (N_6670,N_4756,N_5013);
and U6671 (N_6671,N_4793,N_4871);
and U6672 (N_6672,N_5494,N_5605);
xnor U6673 (N_6673,N_5389,N_5691);
nand U6674 (N_6674,N_5875,N_5089);
or U6675 (N_6675,N_5173,N_5711);
nor U6676 (N_6676,N_5585,N_5528);
and U6677 (N_6677,N_5541,N_5578);
nor U6678 (N_6678,N_4937,N_5314);
and U6679 (N_6679,N_5764,N_5085);
nor U6680 (N_6680,N_4563,N_5250);
nor U6681 (N_6681,N_5069,N_5660);
and U6682 (N_6682,N_5039,N_4536);
or U6683 (N_6683,N_4957,N_4792);
xnor U6684 (N_6684,N_4748,N_5356);
xor U6685 (N_6685,N_5275,N_4501);
nor U6686 (N_6686,N_5537,N_4703);
nand U6687 (N_6687,N_4562,N_5004);
xnor U6688 (N_6688,N_5035,N_5658);
and U6689 (N_6689,N_5459,N_5482);
or U6690 (N_6690,N_5345,N_5539);
or U6691 (N_6691,N_5439,N_5071);
xnor U6692 (N_6692,N_5616,N_5772);
nor U6693 (N_6693,N_4905,N_4966);
xnor U6694 (N_6694,N_5502,N_4708);
and U6695 (N_6695,N_4683,N_5978);
nor U6696 (N_6696,N_5533,N_5686);
or U6697 (N_6697,N_5489,N_5193);
nand U6698 (N_6698,N_4817,N_4771);
or U6699 (N_6699,N_4555,N_5680);
or U6700 (N_6700,N_5381,N_5778);
nand U6701 (N_6701,N_5307,N_5731);
nand U6702 (N_6702,N_5860,N_5673);
and U6703 (N_6703,N_5995,N_5424);
xnor U6704 (N_6704,N_5216,N_5574);
nand U6705 (N_6705,N_5503,N_5911);
or U6706 (N_6706,N_5335,N_5289);
or U6707 (N_6707,N_5048,N_5758);
nor U6708 (N_6708,N_5845,N_4639);
and U6709 (N_6709,N_5858,N_4715);
and U6710 (N_6710,N_4506,N_4576);
nand U6711 (N_6711,N_5830,N_5224);
nor U6712 (N_6712,N_5588,N_5033);
nand U6713 (N_6713,N_4574,N_5773);
nand U6714 (N_6714,N_4785,N_4700);
xnor U6715 (N_6715,N_5030,N_5378);
xor U6716 (N_6716,N_5150,N_4901);
nand U6717 (N_6717,N_5552,N_5358);
nor U6718 (N_6718,N_5805,N_4770);
nand U6719 (N_6719,N_5891,N_5536);
xnor U6720 (N_6720,N_5637,N_5729);
nor U6721 (N_6721,N_5233,N_5849);
xor U6722 (N_6722,N_4532,N_5238);
nor U6723 (N_6723,N_5641,N_5108);
nand U6724 (N_6724,N_5264,N_4575);
and U6725 (N_6725,N_5935,N_5018);
nand U6726 (N_6726,N_5937,N_5677);
xor U6727 (N_6727,N_5600,N_5789);
or U6728 (N_6728,N_4691,N_5523);
xnor U6729 (N_6729,N_4947,N_5488);
nor U6730 (N_6730,N_4878,N_5506);
nand U6731 (N_6731,N_5349,N_4679);
and U6732 (N_6732,N_4581,N_5344);
nor U6733 (N_6733,N_5448,N_5981);
nor U6734 (N_6734,N_5113,N_4987);
nor U6735 (N_6735,N_4641,N_4636);
nand U6736 (N_6736,N_4738,N_4859);
or U6737 (N_6737,N_5474,N_4824);
and U6738 (N_6738,N_4813,N_5186);
xor U6739 (N_6739,N_5992,N_5134);
nor U6740 (N_6740,N_5412,N_4518);
nor U6741 (N_6741,N_5262,N_4887);
or U6742 (N_6742,N_5557,N_5282);
and U6743 (N_6743,N_5847,N_5662);
xnor U6744 (N_6744,N_5192,N_5703);
nand U6745 (N_6745,N_5583,N_5025);
xnor U6746 (N_6746,N_5095,N_5288);
nand U6747 (N_6747,N_4755,N_5675);
nor U6748 (N_6748,N_4960,N_5260);
or U6749 (N_6749,N_5495,N_4739);
xor U6750 (N_6750,N_5964,N_5233);
or U6751 (N_6751,N_5831,N_5533);
xnor U6752 (N_6752,N_5299,N_5990);
and U6753 (N_6753,N_5231,N_5101);
nor U6754 (N_6754,N_4582,N_4939);
nor U6755 (N_6755,N_4777,N_5542);
and U6756 (N_6756,N_5863,N_5822);
nand U6757 (N_6757,N_4761,N_4649);
and U6758 (N_6758,N_4855,N_4675);
or U6759 (N_6759,N_5323,N_5424);
or U6760 (N_6760,N_5073,N_5745);
xor U6761 (N_6761,N_5668,N_5746);
or U6762 (N_6762,N_5839,N_5390);
xnor U6763 (N_6763,N_4996,N_4667);
xor U6764 (N_6764,N_5750,N_4854);
nor U6765 (N_6765,N_4509,N_5655);
or U6766 (N_6766,N_5152,N_4665);
nand U6767 (N_6767,N_5439,N_5909);
xnor U6768 (N_6768,N_5294,N_5079);
nand U6769 (N_6769,N_4974,N_5640);
nand U6770 (N_6770,N_5102,N_5177);
or U6771 (N_6771,N_5195,N_5399);
nor U6772 (N_6772,N_4923,N_4639);
xor U6773 (N_6773,N_4689,N_5186);
nand U6774 (N_6774,N_5335,N_5699);
xnor U6775 (N_6775,N_5312,N_5122);
nand U6776 (N_6776,N_4955,N_4522);
nor U6777 (N_6777,N_4790,N_4979);
or U6778 (N_6778,N_5834,N_4811);
and U6779 (N_6779,N_4691,N_5734);
and U6780 (N_6780,N_5166,N_4975);
and U6781 (N_6781,N_5995,N_5774);
nor U6782 (N_6782,N_4664,N_5810);
or U6783 (N_6783,N_5668,N_5808);
and U6784 (N_6784,N_5501,N_4529);
xor U6785 (N_6785,N_4871,N_5284);
or U6786 (N_6786,N_4689,N_4877);
and U6787 (N_6787,N_4994,N_5827);
and U6788 (N_6788,N_4996,N_4886);
xnor U6789 (N_6789,N_5816,N_5352);
or U6790 (N_6790,N_5710,N_5426);
xnor U6791 (N_6791,N_4972,N_5862);
nand U6792 (N_6792,N_4716,N_5944);
or U6793 (N_6793,N_5131,N_5039);
and U6794 (N_6794,N_5820,N_5881);
and U6795 (N_6795,N_4700,N_4637);
xor U6796 (N_6796,N_4968,N_5967);
or U6797 (N_6797,N_5412,N_4680);
xor U6798 (N_6798,N_5106,N_4600);
nand U6799 (N_6799,N_5350,N_4806);
nor U6800 (N_6800,N_5845,N_5888);
nand U6801 (N_6801,N_4919,N_4958);
nand U6802 (N_6802,N_5575,N_5425);
xnor U6803 (N_6803,N_4569,N_4836);
xnor U6804 (N_6804,N_5289,N_5488);
nor U6805 (N_6805,N_5253,N_5939);
or U6806 (N_6806,N_5012,N_5842);
or U6807 (N_6807,N_4646,N_5857);
and U6808 (N_6808,N_5231,N_4897);
nand U6809 (N_6809,N_5495,N_4844);
and U6810 (N_6810,N_4657,N_4765);
or U6811 (N_6811,N_5750,N_4983);
nand U6812 (N_6812,N_5652,N_5734);
nor U6813 (N_6813,N_4667,N_4912);
xnor U6814 (N_6814,N_4924,N_4911);
xor U6815 (N_6815,N_5741,N_5193);
or U6816 (N_6816,N_5588,N_5274);
and U6817 (N_6817,N_5882,N_5141);
or U6818 (N_6818,N_5680,N_4618);
and U6819 (N_6819,N_4545,N_5929);
nand U6820 (N_6820,N_4665,N_5283);
or U6821 (N_6821,N_4521,N_5515);
and U6822 (N_6822,N_4722,N_5860);
nor U6823 (N_6823,N_4574,N_5513);
and U6824 (N_6824,N_5421,N_4549);
or U6825 (N_6825,N_5953,N_5639);
nand U6826 (N_6826,N_5512,N_5749);
and U6827 (N_6827,N_5068,N_4767);
nand U6828 (N_6828,N_5754,N_5107);
nor U6829 (N_6829,N_5349,N_5120);
and U6830 (N_6830,N_5136,N_5840);
nand U6831 (N_6831,N_4892,N_5847);
and U6832 (N_6832,N_5653,N_5081);
or U6833 (N_6833,N_5567,N_4724);
nand U6834 (N_6834,N_4636,N_5783);
or U6835 (N_6835,N_5942,N_4529);
or U6836 (N_6836,N_4862,N_5627);
or U6837 (N_6837,N_5757,N_5185);
and U6838 (N_6838,N_5124,N_5456);
and U6839 (N_6839,N_5328,N_4768);
and U6840 (N_6840,N_5558,N_5281);
and U6841 (N_6841,N_5449,N_5861);
and U6842 (N_6842,N_4981,N_5385);
or U6843 (N_6843,N_5895,N_5103);
nor U6844 (N_6844,N_5710,N_5200);
or U6845 (N_6845,N_4942,N_4714);
xnor U6846 (N_6846,N_5777,N_4740);
nand U6847 (N_6847,N_4905,N_4731);
and U6848 (N_6848,N_4685,N_5779);
or U6849 (N_6849,N_4689,N_5834);
nor U6850 (N_6850,N_4880,N_4865);
and U6851 (N_6851,N_5603,N_4588);
or U6852 (N_6852,N_5127,N_4786);
xor U6853 (N_6853,N_5870,N_5444);
nor U6854 (N_6854,N_4501,N_5870);
nor U6855 (N_6855,N_5821,N_4639);
and U6856 (N_6856,N_5525,N_4593);
and U6857 (N_6857,N_4567,N_5365);
and U6858 (N_6858,N_4786,N_4840);
xor U6859 (N_6859,N_5304,N_4510);
or U6860 (N_6860,N_5251,N_5401);
and U6861 (N_6861,N_5616,N_5026);
nand U6862 (N_6862,N_4997,N_5698);
nand U6863 (N_6863,N_4678,N_5850);
and U6864 (N_6864,N_4710,N_5446);
or U6865 (N_6865,N_4707,N_5469);
nand U6866 (N_6866,N_5212,N_5499);
nand U6867 (N_6867,N_4592,N_5349);
nor U6868 (N_6868,N_4962,N_5070);
or U6869 (N_6869,N_5915,N_5356);
nand U6870 (N_6870,N_4614,N_5205);
nor U6871 (N_6871,N_4584,N_5385);
and U6872 (N_6872,N_5922,N_4829);
and U6873 (N_6873,N_5751,N_5155);
and U6874 (N_6874,N_4586,N_5704);
nand U6875 (N_6875,N_5056,N_4873);
or U6876 (N_6876,N_4858,N_4595);
nand U6877 (N_6877,N_4596,N_5310);
and U6878 (N_6878,N_5054,N_5940);
or U6879 (N_6879,N_4546,N_4623);
and U6880 (N_6880,N_5255,N_5102);
nand U6881 (N_6881,N_5809,N_4797);
nor U6882 (N_6882,N_5267,N_5765);
or U6883 (N_6883,N_5102,N_4564);
nand U6884 (N_6884,N_5206,N_5124);
or U6885 (N_6885,N_5588,N_5786);
nand U6886 (N_6886,N_5796,N_5791);
nand U6887 (N_6887,N_4816,N_5721);
nand U6888 (N_6888,N_5858,N_5980);
xnor U6889 (N_6889,N_5367,N_5319);
or U6890 (N_6890,N_5363,N_4652);
xor U6891 (N_6891,N_5616,N_5110);
nand U6892 (N_6892,N_5494,N_5764);
xnor U6893 (N_6893,N_5229,N_5048);
nor U6894 (N_6894,N_5000,N_4947);
nor U6895 (N_6895,N_5523,N_5924);
or U6896 (N_6896,N_5738,N_4652);
and U6897 (N_6897,N_4999,N_5384);
nand U6898 (N_6898,N_5907,N_4907);
and U6899 (N_6899,N_4601,N_4816);
xor U6900 (N_6900,N_5794,N_5557);
xor U6901 (N_6901,N_4833,N_5692);
or U6902 (N_6902,N_5138,N_4657);
nand U6903 (N_6903,N_5594,N_4849);
xor U6904 (N_6904,N_5616,N_4802);
or U6905 (N_6905,N_5721,N_5444);
nand U6906 (N_6906,N_4702,N_5637);
or U6907 (N_6907,N_5670,N_5113);
nor U6908 (N_6908,N_5319,N_5389);
xnor U6909 (N_6909,N_5714,N_4883);
or U6910 (N_6910,N_4703,N_5840);
and U6911 (N_6911,N_5152,N_5532);
and U6912 (N_6912,N_4744,N_5613);
nand U6913 (N_6913,N_5960,N_5622);
nand U6914 (N_6914,N_5490,N_5370);
nor U6915 (N_6915,N_4937,N_5221);
or U6916 (N_6916,N_5159,N_4886);
xor U6917 (N_6917,N_5248,N_5675);
xor U6918 (N_6918,N_4754,N_5154);
nand U6919 (N_6919,N_5458,N_4896);
and U6920 (N_6920,N_4926,N_5029);
nand U6921 (N_6921,N_4859,N_4526);
nor U6922 (N_6922,N_5508,N_4611);
xor U6923 (N_6923,N_5915,N_5885);
xor U6924 (N_6924,N_5874,N_4574);
nor U6925 (N_6925,N_5410,N_4547);
nand U6926 (N_6926,N_4830,N_5441);
xnor U6927 (N_6927,N_5390,N_4604);
and U6928 (N_6928,N_4705,N_5972);
and U6929 (N_6929,N_5138,N_5695);
nand U6930 (N_6930,N_5160,N_5581);
or U6931 (N_6931,N_5100,N_5098);
nor U6932 (N_6932,N_4977,N_4731);
nand U6933 (N_6933,N_4599,N_5537);
and U6934 (N_6934,N_5082,N_5640);
xnor U6935 (N_6935,N_4747,N_5313);
and U6936 (N_6936,N_5431,N_5034);
nand U6937 (N_6937,N_4581,N_5844);
and U6938 (N_6938,N_4740,N_5092);
xor U6939 (N_6939,N_4907,N_5455);
nand U6940 (N_6940,N_5165,N_5428);
xor U6941 (N_6941,N_5113,N_5698);
xnor U6942 (N_6942,N_4748,N_5823);
or U6943 (N_6943,N_4816,N_4959);
or U6944 (N_6944,N_5324,N_5497);
and U6945 (N_6945,N_5913,N_5655);
nand U6946 (N_6946,N_4946,N_5254);
or U6947 (N_6947,N_5999,N_5324);
nor U6948 (N_6948,N_4678,N_5936);
xor U6949 (N_6949,N_5840,N_4839);
nor U6950 (N_6950,N_5420,N_4736);
and U6951 (N_6951,N_5402,N_5032);
or U6952 (N_6952,N_5263,N_5699);
nand U6953 (N_6953,N_4892,N_5401);
xnor U6954 (N_6954,N_5296,N_5070);
nand U6955 (N_6955,N_5500,N_5101);
xor U6956 (N_6956,N_4974,N_5292);
nor U6957 (N_6957,N_5869,N_4708);
nor U6958 (N_6958,N_4511,N_5762);
nor U6959 (N_6959,N_5209,N_5785);
nor U6960 (N_6960,N_4547,N_5738);
nor U6961 (N_6961,N_4804,N_5266);
xnor U6962 (N_6962,N_5470,N_5159);
or U6963 (N_6963,N_5317,N_5920);
xor U6964 (N_6964,N_5917,N_5811);
or U6965 (N_6965,N_5808,N_5262);
and U6966 (N_6966,N_4561,N_5729);
nor U6967 (N_6967,N_4845,N_5885);
nor U6968 (N_6968,N_5279,N_5826);
and U6969 (N_6969,N_5448,N_5189);
and U6970 (N_6970,N_5088,N_5191);
nand U6971 (N_6971,N_4669,N_5601);
xnor U6972 (N_6972,N_5546,N_5732);
xor U6973 (N_6973,N_4537,N_5049);
xnor U6974 (N_6974,N_5450,N_4593);
nor U6975 (N_6975,N_5582,N_5800);
nand U6976 (N_6976,N_5225,N_5395);
nand U6977 (N_6977,N_4996,N_5487);
nand U6978 (N_6978,N_5086,N_4761);
or U6979 (N_6979,N_5640,N_5738);
xor U6980 (N_6980,N_5201,N_5258);
or U6981 (N_6981,N_5140,N_4534);
nor U6982 (N_6982,N_5675,N_5315);
nand U6983 (N_6983,N_5182,N_4997);
nor U6984 (N_6984,N_4530,N_4528);
nand U6985 (N_6985,N_5987,N_5940);
or U6986 (N_6986,N_5099,N_5988);
nand U6987 (N_6987,N_5253,N_4634);
xor U6988 (N_6988,N_5542,N_5507);
and U6989 (N_6989,N_5255,N_5585);
nand U6990 (N_6990,N_5492,N_4933);
and U6991 (N_6991,N_5126,N_5144);
xnor U6992 (N_6992,N_5515,N_5533);
and U6993 (N_6993,N_4952,N_4985);
nand U6994 (N_6994,N_4724,N_5889);
xor U6995 (N_6995,N_4741,N_5505);
and U6996 (N_6996,N_5989,N_4554);
nand U6997 (N_6997,N_5693,N_5981);
nor U6998 (N_6998,N_5222,N_5057);
nor U6999 (N_6999,N_4962,N_4528);
nand U7000 (N_7000,N_4874,N_5568);
and U7001 (N_7001,N_4943,N_5007);
or U7002 (N_7002,N_4554,N_4504);
nand U7003 (N_7003,N_5734,N_5584);
and U7004 (N_7004,N_5065,N_4503);
and U7005 (N_7005,N_4648,N_5004);
or U7006 (N_7006,N_5084,N_5317);
xnor U7007 (N_7007,N_4620,N_5712);
or U7008 (N_7008,N_5826,N_5488);
xnor U7009 (N_7009,N_5045,N_5196);
and U7010 (N_7010,N_5348,N_5587);
nor U7011 (N_7011,N_5881,N_4534);
and U7012 (N_7012,N_5304,N_5038);
nor U7013 (N_7013,N_4597,N_5580);
and U7014 (N_7014,N_5163,N_5719);
xnor U7015 (N_7015,N_5958,N_5137);
and U7016 (N_7016,N_5734,N_5825);
nand U7017 (N_7017,N_5488,N_4641);
nor U7018 (N_7018,N_5940,N_5974);
xor U7019 (N_7019,N_4798,N_5183);
or U7020 (N_7020,N_5946,N_4967);
or U7021 (N_7021,N_5191,N_4981);
or U7022 (N_7022,N_5232,N_4536);
nand U7023 (N_7023,N_5326,N_4824);
nand U7024 (N_7024,N_5357,N_5883);
xor U7025 (N_7025,N_5464,N_5635);
nor U7026 (N_7026,N_5159,N_5769);
xnor U7027 (N_7027,N_4610,N_5832);
or U7028 (N_7028,N_5460,N_5370);
and U7029 (N_7029,N_4502,N_5575);
nand U7030 (N_7030,N_4932,N_5303);
nand U7031 (N_7031,N_5115,N_4601);
or U7032 (N_7032,N_4745,N_4698);
nor U7033 (N_7033,N_4509,N_5756);
nand U7034 (N_7034,N_5443,N_4822);
xor U7035 (N_7035,N_5775,N_5103);
nand U7036 (N_7036,N_5742,N_5690);
nor U7037 (N_7037,N_4724,N_5873);
and U7038 (N_7038,N_5370,N_5036);
nand U7039 (N_7039,N_4805,N_5618);
and U7040 (N_7040,N_5570,N_5985);
and U7041 (N_7041,N_4674,N_5454);
or U7042 (N_7042,N_5599,N_5182);
or U7043 (N_7043,N_4706,N_4977);
and U7044 (N_7044,N_5321,N_4802);
nand U7045 (N_7045,N_5933,N_4503);
and U7046 (N_7046,N_4738,N_5296);
or U7047 (N_7047,N_5100,N_5788);
or U7048 (N_7048,N_5296,N_5728);
nand U7049 (N_7049,N_5092,N_5246);
or U7050 (N_7050,N_5108,N_5788);
and U7051 (N_7051,N_5107,N_5146);
xnor U7052 (N_7052,N_4731,N_4539);
nand U7053 (N_7053,N_4657,N_4611);
nand U7054 (N_7054,N_5010,N_4593);
or U7055 (N_7055,N_4798,N_5608);
xor U7056 (N_7056,N_5564,N_5686);
xnor U7057 (N_7057,N_5037,N_5742);
nor U7058 (N_7058,N_5147,N_5609);
or U7059 (N_7059,N_5027,N_5605);
nor U7060 (N_7060,N_5203,N_5941);
xnor U7061 (N_7061,N_5219,N_5036);
and U7062 (N_7062,N_4612,N_5021);
xnor U7063 (N_7063,N_5838,N_5974);
and U7064 (N_7064,N_5515,N_5501);
nor U7065 (N_7065,N_4832,N_5980);
nor U7066 (N_7066,N_5203,N_4806);
nor U7067 (N_7067,N_5714,N_4614);
or U7068 (N_7068,N_5053,N_5068);
nor U7069 (N_7069,N_4781,N_5502);
or U7070 (N_7070,N_5943,N_5851);
nand U7071 (N_7071,N_4929,N_5657);
xnor U7072 (N_7072,N_4729,N_4694);
and U7073 (N_7073,N_5648,N_5980);
or U7074 (N_7074,N_5506,N_5557);
and U7075 (N_7075,N_5656,N_5691);
nor U7076 (N_7076,N_5759,N_5781);
and U7077 (N_7077,N_5302,N_5935);
xnor U7078 (N_7078,N_5727,N_5075);
xor U7079 (N_7079,N_5867,N_4807);
and U7080 (N_7080,N_4866,N_4754);
nor U7081 (N_7081,N_5975,N_4879);
nor U7082 (N_7082,N_5936,N_5108);
and U7083 (N_7083,N_5026,N_5906);
xnor U7084 (N_7084,N_5540,N_4834);
xnor U7085 (N_7085,N_5838,N_5352);
nor U7086 (N_7086,N_5255,N_4504);
and U7087 (N_7087,N_4691,N_5968);
nand U7088 (N_7088,N_4802,N_4766);
nor U7089 (N_7089,N_4936,N_4555);
nor U7090 (N_7090,N_4934,N_4677);
xor U7091 (N_7091,N_4711,N_5707);
nand U7092 (N_7092,N_4834,N_5985);
xor U7093 (N_7093,N_5477,N_5589);
nand U7094 (N_7094,N_4855,N_4770);
xor U7095 (N_7095,N_4920,N_5464);
and U7096 (N_7096,N_5914,N_4688);
nor U7097 (N_7097,N_5669,N_4940);
and U7098 (N_7098,N_5923,N_5888);
nand U7099 (N_7099,N_5210,N_4763);
and U7100 (N_7100,N_5832,N_4697);
and U7101 (N_7101,N_5363,N_5633);
xnor U7102 (N_7102,N_5885,N_5146);
xnor U7103 (N_7103,N_5708,N_5487);
nand U7104 (N_7104,N_5513,N_5371);
and U7105 (N_7105,N_5985,N_5033);
nor U7106 (N_7106,N_5353,N_5030);
or U7107 (N_7107,N_5494,N_5241);
nand U7108 (N_7108,N_5804,N_5483);
or U7109 (N_7109,N_5858,N_4878);
xor U7110 (N_7110,N_5343,N_4593);
nand U7111 (N_7111,N_4720,N_4947);
nor U7112 (N_7112,N_5472,N_5422);
nand U7113 (N_7113,N_5169,N_5781);
nor U7114 (N_7114,N_5780,N_5973);
xor U7115 (N_7115,N_5363,N_5001);
nand U7116 (N_7116,N_5524,N_5980);
and U7117 (N_7117,N_5141,N_5271);
or U7118 (N_7118,N_4893,N_5837);
or U7119 (N_7119,N_5626,N_4935);
and U7120 (N_7120,N_5534,N_5424);
nor U7121 (N_7121,N_4502,N_4628);
or U7122 (N_7122,N_5394,N_5050);
and U7123 (N_7123,N_4767,N_5255);
nand U7124 (N_7124,N_5914,N_4643);
xor U7125 (N_7125,N_5096,N_4947);
nor U7126 (N_7126,N_5986,N_5797);
and U7127 (N_7127,N_4833,N_5778);
nor U7128 (N_7128,N_5684,N_5275);
nand U7129 (N_7129,N_5393,N_5396);
and U7130 (N_7130,N_4602,N_4680);
nor U7131 (N_7131,N_5739,N_5211);
or U7132 (N_7132,N_5662,N_4826);
xnor U7133 (N_7133,N_4528,N_5892);
and U7134 (N_7134,N_5861,N_4729);
nor U7135 (N_7135,N_5650,N_5386);
nor U7136 (N_7136,N_5107,N_5780);
nor U7137 (N_7137,N_5789,N_4992);
and U7138 (N_7138,N_4887,N_4851);
xor U7139 (N_7139,N_5611,N_5011);
and U7140 (N_7140,N_5842,N_5343);
xor U7141 (N_7141,N_4798,N_4556);
xnor U7142 (N_7142,N_5351,N_4741);
and U7143 (N_7143,N_5962,N_5782);
nand U7144 (N_7144,N_4614,N_5422);
xor U7145 (N_7145,N_5470,N_4694);
and U7146 (N_7146,N_5684,N_5230);
and U7147 (N_7147,N_4990,N_5533);
or U7148 (N_7148,N_5216,N_4561);
nand U7149 (N_7149,N_5292,N_5666);
and U7150 (N_7150,N_5434,N_5756);
nand U7151 (N_7151,N_4623,N_5310);
and U7152 (N_7152,N_5370,N_5259);
xor U7153 (N_7153,N_4766,N_5977);
nand U7154 (N_7154,N_5367,N_4765);
or U7155 (N_7155,N_5578,N_4994);
nand U7156 (N_7156,N_4605,N_5528);
and U7157 (N_7157,N_5749,N_4938);
nor U7158 (N_7158,N_5873,N_5256);
nor U7159 (N_7159,N_5867,N_5132);
and U7160 (N_7160,N_5778,N_5755);
nor U7161 (N_7161,N_5026,N_5622);
or U7162 (N_7162,N_5987,N_5626);
and U7163 (N_7163,N_5823,N_5968);
and U7164 (N_7164,N_5674,N_5051);
or U7165 (N_7165,N_5669,N_4580);
nor U7166 (N_7166,N_5280,N_5676);
nor U7167 (N_7167,N_4789,N_5760);
and U7168 (N_7168,N_5328,N_4938);
and U7169 (N_7169,N_4664,N_4642);
nor U7170 (N_7170,N_4923,N_5903);
or U7171 (N_7171,N_5263,N_4623);
xor U7172 (N_7172,N_5034,N_5850);
and U7173 (N_7173,N_5782,N_5321);
nor U7174 (N_7174,N_4618,N_5586);
and U7175 (N_7175,N_4545,N_4683);
xor U7176 (N_7176,N_4513,N_4745);
nand U7177 (N_7177,N_5350,N_5127);
and U7178 (N_7178,N_4795,N_5146);
nor U7179 (N_7179,N_5123,N_5356);
nor U7180 (N_7180,N_5850,N_5692);
and U7181 (N_7181,N_4596,N_4892);
and U7182 (N_7182,N_4785,N_5271);
nor U7183 (N_7183,N_5831,N_5241);
and U7184 (N_7184,N_5427,N_5759);
nor U7185 (N_7185,N_4583,N_5327);
nor U7186 (N_7186,N_4730,N_4885);
and U7187 (N_7187,N_5439,N_4608);
and U7188 (N_7188,N_5830,N_4563);
nor U7189 (N_7189,N_5710,N_5005);
and U7190 (N_7190,N_5378,N_5026);
xnor U7191 (N_7191,N_5073,N_4743);
nand U7192 (N_7192,N_4527,N_5069);
nor U7193 (N_7193,N_5080,N_4968);
nand U7194 (N_7194,N_5567,N_5893);
nand U7195 (N_7195,N_5788,N_4933);
nand U7196 (N_7196,N_5526,N_5058);
nand U7197 (N_7197,N_5812,N_5588);
xnor U7198 (N_7198,N_5224,N_4628);
nor U7199 (N_7199,N_4664,N_5807);
nor U7200 (N_7200,N_5611,N_4660);
nor U7201 (N_7201,N_5400,N_4908);
and U7202 (N_7202,N_5416,N_4569);
xor U7203 (N_7203,N_5651,N_5777);
nor U7204 (N_7204,N_5420,N_5381);
nand U7205 (N_7205,N_4586,N_5138);
and U7206 (N_7206,N_5450,N_4970);
or U7207 (N_7207,N_4664,N_4764);
nand U7208 (N_7208,N_4773,N_4965);
and U7209 (N_7209,N_5764,N_5289);
nor U7210 (N_7210,N_4674,N_5999);
xor U7211 (N_7211,N_5617,N_5278);
or U7212 (N_7212,N_5172,N_5280);
or U7213 (N_7213,N_4952,N_4768);
nand U7214 (N_7214,N_4931,N_5223);
or U7215 (N_7215,N_5602,N_5261);
or U7216 (N_7216,N_4976,N_5572);
nor U7217 (N_7217,N_5581,N_4508);
and U7218 (N_7218,N_5557,N_4873);
nand U7219 (N_7219,N_5971,N_5338);
and U7220 (N_7220,N_4906,N_4958);
and U7221 (N_7221,N_5253,N_5422);
and U7222 (N_7222,N_5472,N_5093);
nand U7223 (N_7223,N_4629,N_4743);
and U7224 (N_7224,N_5313,N_5995);
and U7225 (N_7225,N_5335,N_5191);
and U7226 (N_7226,N_5320,N_5034);
nand U7227 (N_7227,N_4987,N_5137);
nor U7228 (N_7228,N_5521,N_5675);
and U7229 (N_7229,N_5595,N_5142);
nor U7230 (N_7230,N_5758,N_5415);
nor U7231 (N_7231,N_5125,N_4764);
and U7232 (N_7232,N_5070,N_4879);
nand U7233 (N_7233,N_5380,N_4557);
and U7234 (N_7234,N_5233,N_5487);
and U7235 (N_7235,N_4990,N_5713);
or U7236 (N_7236,N_5826,N_5281);
xor U7237 (N_7237,N_5392,N_5524);
nor U7238 (N_7238,N_5392,N_4552);
or U7239 (N_7239,N_4836,N_4979);
xor U7240 (N_7240,N_5887,N_4778);
nand U7241 (N_7241,N_4937,N_5749);
nor U7242 (N_7242,N_5786,N_5077);
nor U7243 (N_7243,N_5552,N_5714);
and U7244 (N_7244,N_5593,N_4655);
nor U7245 (N_7245,N_4635,N_5368);
xnor U7246 (N_7246,N_5735,N_5613);
nand U7247 (N_7247,N_4772,N_4843);
xnor U7248 (N_7248,N_5848,N_5672);
nor U7249 (N_7249,N_5027,N_5497);
or U7250 (N_7250,N_5870,N_5064);
xor U7251 (N_7251,N_5141,N_5974);
and U7252 (N_7252,N_5835,N_5152);
nor U7253 (N_7253,N_5274,N_5500);
nor U7254 (N_7254,N_5605,N_5585);
or U7255 (N_7255,N_5744,N_5931);
and U7256 (N_7256,N_4834,N_5017);
nor U7257 (N_7257,N_5023,N_4974);
or U7258 (N_7258,N_5506,N_5754);
xor U7259 (N_7259,N_5275,N_4815);
or U7260 (N_7260,N_5443,N_4965);
xnor U7261 (N_7261,N_5825,N_5395);
and U7262 (N_7262,N_5982,N_4830);
nand U7263 (N_7263,N_5677,N_5576);
and U7264 (N_7264,N_5692,N_4789);
or U7265 (N_7265,N_4705,N_5039);
nand U7266 (N_7266,N_5006,N_5521);
nor U7267 (N_7267,N_5047,N_4747);
nand U7268 (N_7268,N_5974,N_5458);
and U7269 (N_7269,N_5870,N_5026);
nor U7270 (N_7270,N_5746,N_5869);
nor U7271 (N_7271,N_4687,N_4527);
nand U7272 (N_7272,N_5769,N_4966);
or U7273 (N_7273,N_4587,N_5915);
nor U7274 (N_7274,N_5932,N_4780);
nor U7275 (N_7275,N_5034,N_5159);
nor U7276 (N_7276,N_5084,N_5343);
nand U7277 (N_7277,N_5712,N_4583);
nor U7278 (N_7278,N_5930,N_5441);
and U7279 (N_7279,N_5682,N_5859);
or U7280 (N_7280,N_4761,N_4723);
or U7281 (N_7281,N_4878,N_5701);
or U7282 (N_7282,N_5210,N_5753);
nor U7283 (N_7283,N_5580,N_5760);
and U7284 (N_7284,N_5576,N_5314);
and U7285 (N_7285,N_5791,N_4509);
nand U7286 (N_7286,N_5476,N_5238);
nor U7287 (N_7287,N_5231,N_4636);
xor U7288 (N_7288,N_5737,N_5356);
and U7289 (N_7289,N_5705,N_5451);
nor U7290 (N_7290,N_5686,N_5167);
xnor U7291 (N_7291,N_5401,N_5023);
and U7292 (N_7292,N_5620,N_5455);
xor U7293 (N_7293,N_5981,N_5628);
nand U7294 (N_7294,N_5600,N_5408);
xor U7295 (N_7295,N_5298,N_5970);
or U7296 (N_7296,N_5487,N_5151);
nor U7297 (N_7297,N_4739,N_5474);
nor U7298 (N_7298,N_5821,N_5658);
and U7299 (N_7299,N_5664,N_4854);
or U7300 (N_7300,N_4726,N_4891);
nor U7301 (N_7301,N_5240,N_5825);
and U7302 (N_7302,N_4680,N_5481);
xor U7303 (N_7303,N_5299,N_4947);
or U7304 (N_7304,N_4968,N_5564);
or U7305 (N_7305,N_5542,N_4797);
and U7306 (N_7306,N_5986,N_4612);
or U7307 (N_7307,N_5741,N_5960);
and U7308 (N_7308,N_5881,N_4558);
nand U7309 (N_7309,N_5310,N_4975);
nand U7310 (N_7310,N_5741,N_4883);
xor U7311 (N_7311,N_5436,N_5617);
nand U7312 (N_7312,N_5616,N_5282);
xor U7313 (N_7313,N_5055,N_5003);
or U7314 (N_7314,N_4960,N_5947);
and U7315 (N_7315,N_5830,N_4874);
and U7316 (N_7316,N_5292,N_5925);
xnor U7317 (N_7317,N_5698,N_4775);
or U7318 (N_7318,N_4802,N_5856);
nand U7319 (N_7319,N_5697,N_5541);
nor U7320 (N_7320,N_4675,N_5559);
xnor U7321 (N_7321,N_5529,N_4887);
xnor U7322 (N_7322,N_5122,N_5391);
xor U7323 (N_7323,N_5119,N_5474);
and U7324 (N_7324,N_5408,N_4853);
or U7325 (N_7325,N_5810,N_4897);
and U7326 (N_7326,N_4945,N_5657);
nor U7327 (N_7327,N_5643,N_4597);
or U7328 (N_7328,N_5833,N_5346);
xnor U7329 (N_7329,N_5377,N_5213);
or U7330 (N_7330,N_5885,N_5280);
nor U7331 (N_7331,N_5697,N_4842);
nand U7332 (N_7332,N_5216,N_5516);
and U7333 (N_7333,N_5959,N_4898);
and U7334 (N_7334,N_4548,N_5653);
or U7335 (N_7335,N_4706,N_4580);
nand U7336 (N_7336,N_5582,N_4835);
nor U7337 (N_7337,N_5469,N_5679);
nand U7338 (N_7338,N_5880,N_4563);
nand U7339 (N_7339,N_5430,N_4526);
xnor U7340 (N_7340,N_5602,N_5367);
xnor U7341 (N_7341,N_5987,N_4520);
and U7342 (N_7342,N_5575,N_4967);
or U7343 (N_7343,N_5956,N_5125);
or U7344 (N_7344,N_5556,N_5198);
xnor U7345 (N_7345,N_5315,N_5457);
nor U7346 (N_7346,N_5312,N_5323);
xor U7347 (N_7347,N_5430,N_4827);
nor U7348 (N_7348,N_5648,N_5545);
nand U7349 (N_7349,N_4885,N_5619);
and U7350 (N_7350,N_5003,N_5103);
xnor U7351 (N_7351,N_5841,N_5086);
and U7352 (N_7352,N_5314,N_5131);
xor U7353 (N_7353,N_4898,N_5160);
and U7354 (N_7354,N_4792,N_5689);
or U7355 (N_7355,N_5676,N_5988);
xnor U7356 (N_7356,N_5829,N_5169);
or U7357 (N_7357,N_5601,N_4980);
xor U7358 (N_7358,N_4960,N_4745);
xnor U7359 (N_7359,N_5983,N_5703);
or U7360 (N_7360,N_5400,N_5724);
xor U7361 (N_7361,N_5273,N_4849);
nor U7362 (N_7362,N_4706,N_4826);
nor U7363 (N_7363,N_4568,N_4502);
nor U7364 (N_7364,N_5051,N_5668);
and U7365 (N_7365,N_4991,N_5526);
and U7366 (N_7366,N_5754,N_5563);
nand U7367 (N_7367,N_4801,N_4735);
nor U7368 (N_7368,N_5437,N_4988);
and U7369 (N_7369,N_5859,N_4690);
and U7370 (N_7370,N_5187,N_5357);
and U7371 (N_7371,N_5504,N_5990);
nand U7372 (N_7372,N_5017,N_4592);
nor U7373 (N_7373,N_5343,N_4857);
nand U7374 (N_7374,N_5502,N_5956);
xnor U7375 (N_7375,N_4768,N_4608);
nand U7376 (N_7376,N_5908,N_5556);
or U7377 (N_7377,N_4816,N_5633);
or U7378 (N_7378,N_4924,N_4887);
nand U7379 (N_7379,N_5842,N_4687);
and U7380 (N_7380,N_5636,N_4874);
xor U7381 (N_7381,N_4893,N_4685);
and U7382 (N_7382,N_5626,N_5836);
or U7383 (N_7383,N_4545,N_5840);
or U7384 (N_7384,N_5203,N_5023);
nor U7385 (N_7385,N_4578,N_5694);
and U7386 (N_7386,N_5373,N_4721);
and U7387 (N_7387,N_4746,N_5781);
xor U7388 (N_7388,N_5315,N_5568);
or U7389 (N_7389,N_5616,N_4724);
nand U7390 (N_7390,N_5390,N_5693);
nand U7391 (N_7391,N_5721,N_4755);
and U7392 (N_7392,N_5888,N_5952);
or U7393 (N_7393,N_5604,N_5773);
nor U7394 (N_7394,N_5963,N_5384);
nand U7395 (N_7395,N_4541,N_5912);
xor U7396 (N_7396,N_4843,N_5774);
and U7397 (N_7397,N_4653,N_5468);
nor U7398 (N_7398,N_5017,N_5777);
xnor U7399 (N_7399,N_5506,N_5398);
or U7400 (N_7400,N_5727,N_5268);
xnor U7401 (N_7401,N_5420,N_4580);
or U7402 (N_7402,N_5204,N_5608);
xnor U7403 (N_7403,N_5732,N_5666);
or U7404 (N_7404,N_4586,N_5449);
nand U7405 (N_7405,N_5685,N_4734);
nand U7406 (N_7406,N_5285,N_4595);
nand U7407 (N_7407,N_4810,N_4633);
or U7408 (N_7408,N_5355,N_5348);
and U7409 (N_7409,N_5648,N_5651);
nand U7410 (N_7410,N_4567,N_5423);
xnor U7411 (N_7411,N_5216,N_5958);
and U7412 (N_7412,N_5977,N_5372);
and U7413 (N_7413,N_5947,N_4547);
nand U7414 (N_7414,N_4851,N_5949);
xnor U7415 (N_7415,N_5702,N_5264);
xnor U7416 (N_7416,N_5588,N_5105);
xnor U7417 (N_7417,N_5517,N_5734);
xnor U7418 (N_7418,N_5499,N_4925);
or U7419 (N_7419,N_5066,N_5267);
or U7420 (N_7420,N_5962,N_4568);
xor U7421 (N_7421,N_5065,N_5076);
and U7422 (N_7422,N_4617,N_5984);
and U7423 (N_7423,N_4800,N_5028);
nor U7424 (N_7424,N_5909,N_4890);
nor U7425 (N_7425,N_5530,N_5041);
xnor U7426 (N_7426,N_5233,N_5738);
nand U7427 (N_7427,N_5908,N_5942);
nor U7428 (N_7428,N_5307,N_5902);
nand U7429 (N_7429,N_5041,N_5759);
xor U7430 (N_7430,N_4742,N_5893);
nor U7431 (N_7431,N_5605,N_5163);
xor U7432 (N_7432,N_4980,N_4865);
or U7433 (N_7433,N_5583,N_5829);
nor U7434 (N_7434,N_4679,N_4570);
and U7435 (N_7435,N_5519,N_4674);
nor U7436 (N_7436,N_5881,N_4901);
and U7437 (N_7437,N_5547,N_4794);
and U7438 (N_7438,N_5787,N_5760);
and U7439 (N_7439,N_5695,N_5537);
or U7440 (N_7440,N_5000,N_5816);
or U7441 (N_7441,N_4725,N_4645);
and U7442 (N_7442,N_5873,N_5106);
xor U7443 (N_7443,N_5541,N_5512);
and U7444 (N_7444,N_4778,N_5674);
nand U7445 (N_7445,N_4757,N_5757);
xnor U7446 (N_7446,N_4993,N_5910);
or U7447 (N_7447,N_5908,N_5339);
and U7448 (N_7448,N_4874,N_4846);
or U7449 (N_7449,N_4841,N_5892);
and U7450 (N_7450,N_5492,N_4512);
xnor U7451 (N_7451,N_5262,N_5479);
nand U7452 (N_7452,N_4851,N_5248);
and U7453 (N_7453,N_4767,N_4596);
nand U7454 (N_7454,N_5048,N_5799);
or U7455 (N_7455,N_4714,N_4802);
nand U7456 (N_7456,N_5094,N_4916);
and U7457 (N_7457,N_4761,N_5933);
nand U7458 (N_7458,N_5338,N_5056);
and U7459 (N_7459,N_5542,N_5069);
nand U7460 (N_7460,N_5653,N_5316);
and U7461 (N_7461,N_5570,N_5313);
nor U7462 (N_7462,N_5037,N_5547);
and U7463 (N_7463,N_4990,N_5020);
nand U7464 (N_7464,N_4994,N_4881);
nand U7465 (N_7465,N_4735,N_5325);
nand U7466 (N_7466,N_5493,N_5722);
and U7467 (N_7467,N_4638,N_5540);
xnor U7468 (N_7468,N_5483,N_5065);
and U7469 (N_7469,N_5720,N_4586);
xor U7470 (N_7470,N_5142,N_4518);
and U7471 (N_7471,N_5607,N_5486);
nor U7472 (N_7472,N_5899,N_4814);
or U7473 (N_7473,N_5418,N_4709);
nand U7474 (N_7474,N_5972,N_5675);
or U7475 (N_7475,N_4984,N_5813);
nor U7476 (N_7476,N_4503,N_5351);
nand U7477 (N_7477,N_4798,N_4791);
nand U7478 (N_7478,N_5913,N_5169);
nor U7479 (N_7479,N_4684,N_5719);
xnor U7480 (N_7480,N_5121,N_5408);
xor U7481 (N_7481,N_5532,N_5141);
nand U7482 (N_7482,N_4963,N_4910);
nand U7483 (N_7483,N_4961,N_5284);
nor U7484 (N_7484,N_5807,N_4567);
nand U7485 (N_7485,N_5525,N_5896);
xor U7486 (N_7486,N_4679,N_5239);
nand U7487 (N_7487,N_5645,N_5333);
xnor U7488 (N_7488,N_4826,N_5035);
and U7489 (N_7489,N_5489,N_5151);
nor U7490 (N_7490,N_5137,N_5884);
nor U7491 (N_7491,N_5375,N_5291);
nand U7492 (N_7492,N_4920,N_5021);
nor U7493 (N_7493,N_4924,N_4938);
xor U7494 (N_7494,N_5133,N_4592);
nand U7495 (N_7495,N_5859,N_4769);
nor U7496 (N_7496,N_5085,N_4722);
or U7497 (N_7497,N_5366,N_4784);
xnor U7498 (N_7498,N_4552,N_5167);
or U7499 (N_7499,N_5871,N_5937);
xor U7500 (N_7500,N_6129,N_7139);
nand U7501 (N_7501,N_6868,N_6412);
nor U7502 (N_7502,N_6712,N_6741);
xnor U7503 (N_7503,N_6484,N_6462);
nand U7504 (N_7504,N_6704,N_6325);
xor U7505 (N_7505,N_6249,N_7494);
nand U7506 (N_7506,N_6326,N_6611);
and U7507 (N_7507,N_6901,N_7267);
nor U7508 (N_7508,N_6347,N_7155);
and U7509 (N_7509,N_7362,N_7048);
xnor U7510 (N_7510,N_6582,N_6851);
nand U7511 (N_7511,N_6236,N_7392);
nor U7512 (N_7512,N_7261,N_6899);
or U7513 (N_7513,N_6620,N_7061);
nand U7514 (N_7514,N_6389,N_7219);
nor U7515 (N_7515,N_6109,N_6319);
nor U7516 (N_7516,N_6787,N_6452);
nand U7517 (N_7517,N_7352,N_6059);
nand U7518 (N_7518,N_7310,N_6497);
xnor U7519 (N_7519,N_7264,N_7197);
and U7520 (N_7520,N_6967,N_6124);
xnor U7521 (N_7521,N_7427,N_6070);
nand U7522 (N_7522,N_7449,N_6626);
nand U7523 (N_7523,N_6323,N_7314);
or U7524 (N_7524,N_6309,N_6625);
or U7525 (N_7525,N_6943,N_6633);
xor U7526 (N_7526,N_6227,N_6313);
xnor U7527 (N_7527,N_6371,N_7172);
xnor U7528 (N_7528,N_6890,N_6913);
or U7529 (N_7529,N_6618,N_7320);
xor U7530 (N_7530,N_6599,N_6072);
xor U7531 (N_7531,N_6420,N_6503);
and U7532 (N_7532,N_7017,N_6948);
xnor U7533 (N_7533,N_6841,N_6796);
nor U7534 (N_7534,N_6519,N_6446);
and U7535 (N_7535,N_7159,N_6286);
and U7536 (N_7536,N_6266,N_6487);
or U7537 (N_7537,N_6336,N_6111);
and U7538 (N_7538,N_6630,N_7082);
and U7539 (N_7539,N_7445,N_6729);
nor U7540 (N_7540,N_7063,N_6905);
or U7541 (N_7541,N_6646,N_6264);
and U7542 (N_7542,N_6235,N_6566);
xor U7543 (N_7543,N_6030,N_6894);
nand U7544 (N_7544,N_6064,N_7015);
nand U7545 (N_7545,N_7185,N_6833);
xnor U7546 (N_7546,N_6298,N_6364);
xnor U7547 (N_7547,N_6613,N_6937);
xnor U7548 (N_7548,N_7242,N_6270);
or U7549 (N_7549,N_6492,N_6548);
and U7550 (N_7550,N_6971,N_7198);
nand U7551 (N_7551,N_7254,N_6136);
or U7552 (N_7552,N_6306,N_6550);
nand U7553 (N_7553,N_7128,N_7122);
and U7554 (N_7554,N_6588,N_6220);
nand U7555 (N_7555,N_7078,N_7035);
xor U7556 (N_7556,N_6414,N_7377);
xnor U7557 (N_7557,N_6234,N_6255);
xnor U7558 (N_7558,N_6567,N_7216);
nor U7559 (N_7559,N_6005,N_6048);
or U7560 (N_7560,N_6593,N_7292);
or U7561 (N_7561,N_6038,N_6650);
and U7562 (N_7562,N_7464,N_7084);
and U7563 (N_7563,N_7107,N_7079);
xnor U7564 (N_7564,N_7145,N_6490);
nand U7565 (N_7565,N_6099,N_6056);
and U7566 (N_7566,N_7057,N_6361);
xor U7567 (N_7567,N_6568,N_6804);
nor U7568 (N_7568,N_6277,N_6822);
nor U7569 (N_7569,N_6746,N_6055);
or U7570 (N_7570,N_7325,N_6053);
nand U7571 (N_7571,N_6574,N_6384);
or U7572 (N_7572,N_6366,N_6311);
xnor U7573 (N_7573,N_6376,N_7337);
nor U7574 (N_7574,N_6663,N_6466);
nor U7575 (N_7575,N_6532,N_7273);
and U7576 (N_7576,N_6797,N_6239);
xor U7577 (N_7577,N_6816,N_6421);
and U7578 (N_7578,N_6196,N_7201);
nand U7579 (N_7579,N_6495,N_6541);
nand U7580 (N_7580,N_6597,N_7199);
and U7581 (N_7581,N_6085,N_6723);
nor U7582 (N_7582,N_6839,N_7054);
nor U7583 (N_7583,N_6500,N_6314);
xnor U7584 (N_7584,N_7074,N_6821);
nand U7585 (N_7585,N_6911,N_6138);
nor U7586 (N_7586,N_6223,N_7420);
and U7587 (N_7587,N_6684,N_6212);
or U7588 (N_7588,N_6150,N_6991);
nor U7589 (N_7589,N_6681,N_6502);
nor U7590 (N_7590,N_7289,N_6610);
nand U7591 (N_7591,N_7455,N_6169);
and U7592 (N_7592,N_6986,N_6510);
nor U7593 (N_7593,N_6455,N_6225);
or U7594 (N_7594,N_6962,N_7448);
xor U7595 (N_7595,N_6125,N_6592);
xor U7596 (N_7596,N_6965,N_6852);
or U7597 (N_7597,N_6450,N_7226);
and U7598 (N_7598,N_6357,N_6291);
nand U7599 (N_7599,N_6984,N_6934);
or U7600 (N_7600,N_6843,N_6637);
nand U7601 (N_7601,N_6065,N_6781);
nor U7602 (N_7602,N_6793,N_7453);
and U7603 (N_7603,N_6281,N_6692);
nor U7604 (N_7604,N_6496,N_6387);
nand U7605 (N_7605,N_7348,N_6857);
and U7606 (N_7606,N_6200,N_6020);
or U7607 (N_7607,N_6246,N_6278);
nand U7608 (N_7608,N_6823,N_6101);
nor U7609 (N_7609,N_6267,N_7120);
or U7610 (N_7610,N_6263,N_6832);
nand U7611 (N_7611,N_6044,N_6132);
or U7612 (N_7612,N_6434,N_6602);
nand U7613 (N_7613,N_7477,N_7402);
and U7614 (N_7614,N_6182,N_6732);
nor U7615 (N_7615,N_6092,N_6858);
or U7616 (N_7616,N_6506,N_7460);
nor U7617 (N_7617,N_7333,N_7075);
xnor U7618 (N_7618,N_6390,N_6794);
or U7619 (N_7619,N_6722,N_7398);
nand U7620 (N_7620,N_7425,N_6062);
nor U7621 (N_7621,N_7132,N_7279);
nand U7622 (N_7622,N_6657,N_7415);
xnor U7623 (N_7623,N_6190,N_7255);
xor U7624 (N_7624,N_7375,N_6244);
nor U7625 (N_7625,N_6449,N_6697);
nor U7626 (N_7626,N_6120,N_6607);
and U7627 (N_7627,N_6022,N_7376);
nand U7628 (N_7628,N_6185,N_6825);
nor U7629 (N_7629,N_7131,N_6558);
or U7630 (N_7630,N_6454,N_7134);
nor U7631 (N_7631,N_6711,N_7330);
nor U7632 (N_7632,N_6942,N_6703);
xor U7633 (N_7633,N_6511,N_7496);
xnor U7634 (N_7634,N_6140,N_7150);
nand U7635 (N_7635,N_6609,N_6354);
nor U7636 (N_7636,N_6779,N_6769);
or U7637 (N_7637,N_6456,N_6393);
or U7638 (N_7638,N_6702,N_6583);
nand U7639 (N_7639,N_7162,N_7277);
nand U7640 (N_7640,N_7336,N_7469);
nand U7641 (N_7641,N_6594,N_7104);
and U7642 (N_7642,N_6363,N_7056);
xor U7643 (N_7643,N_7036,N_7157);
nor U7644 (N_7644,N_6501,N_6912);
xor U7645 (N_7645,N_6829,N_6964);
nor U7646 (N_7646,N_7234,N_6772);
nand U7647 (N_7647,N_6049,N_6238);
and U7648 (N_7648,N_6666,N_6745);
and U7649 (N_7649,N_6014,N_7437);
nand U7650 (N_7650,N_7382,N_7108);
or U7651 (N_7651,N_6878,N_7374);
or U7652 (N_7652,N_7285,N_6985);
xor U7653 (N_7653,N_6312,N_7360);
nor U7654 (N_7654,N_6766,N_7443);
xnor U7655 (N_7655,N_6751,N_6262);
and U7656 (N_7656,N_6584,N_6218);
and U7657 (N_7657,N_7149,N_6980);
xnor U7658 (N_7658,N_6369,N_6814);
nor U7659 (N_7659,N_7097,N_6435);
and U7660 (N_7660,N_7462,N_6844);
or U7661 (N_7661,N_6189,N_7371);
xnor U7662 (N_7662,N_7182,N_7429);
nor U7663 (N_7663,N_7004,N_6867);
nand U7664 (N_7664,N_7418,N_7112);
or U7665 (N_7665,N_6368,N_6755);
xnor U7666 (N_7666,N_7235,N_6648);
nor U7667 (N_7667,N_7065,N_7301);
or U7668 (N_7668,N_6727,N_6747);
nand U7669 (N_7669,N_7147,N_7327);
and U7670 (N_7670,N_6860,N_6675);
xnor U7671 (N_7671,N_7372,N_6443);
nor U7672 (N_7672,N_6670,N_7032);
nand U7673 (N_7673,N_6790,N_6830);
and U7674 (N_7674,N_6876,N_6404);
xnor U7675 (N_7675,N_6687,N_6343);
nand U7676 (N_7676,N_7384,N_7091);
xor U7677 (N_7677,N_7302,N_6904);
nand U7678 (N_7678,N_7355,N_6162);
xnor U7679 (N_7679,N_7380,N_7148);
or U7680 (N_7680,N_6688,N_7321);
or U7681 (N_7681,N_6674,N_6098);
xnor U7682 (N_7682,N_6331,N_7208);
nand U7683 (N_7683,N_7110,N_6957);
and U7684 (N_7684,N_6931,N_6505);
and U7685 (N_7685,N_7368,N_7002);
or U7686 (N_7686,N_6335,N_6569);
or U7687 (N_7687,N_6175,N_6093);
and U7688 (N_7688,N_7111,N_6696);
or U7689 (N_7689,N_6103,N_6184);
nor U7690 (N_7690,N_7458,N_7184);
nand U7691 (N_7691,N_6115,N_6046);
nand U7692 (N_7692,N_6021,N_6591);
nand U7693 (N_7693,N_6536,N_7123);
nor U7694 (N_7694,N_7269,N_6820);
or U7695 (N_7695,N_7169,N_6976);
or U7696 (N_7696,N_7188,N_7013);
nor U7697 (N_7697,N_6203,N_6627);
nor U7698 (N_7698,N_6534,N_7158);
xor U7699 (N_7699,N_6889,N_6071);
nand U7700 (N_7700,N_6273,N_6174);
xor U7701 (N_7701,N_6564,N_6595);
or U7702 (N_7702,N_6873,N_6771);
nand U7703 (N_7703,N_7164,N_7117);
and U7704 (N_7704,N_6641,N_7266);
or U7705 (N_7705,N_7177,N_6514);
nand U7706 (N_7706,N_7391,N_6951);
and U7707 (N_7707,N_7105,N_6284);
nor U7708 (N_7708,N_7040,N_6693);
and U7709 (N_7709,N_6661,N_6803);
and U7710 (N_7710,N_7262,N_6458);
nor U7711 (N_7711,N_6679,N_6764);
nor U7712 (N_7712,N_6440,N_7451);
and U7713 (N_7713,N_6955,N_6758);
and U7714 (N_7714,N_6301,N_7282);
and U7715 (N_7715,N_6515,N_6073);
nor U7716 (N_7716,N_6252,N_6612);
nor U7717 (N_7717,N_6016,N_6467);
or U7718 (N_7718,N_7023,N_6815);
nor U7719 (N_7719,N_6530,N_7142);
nor U7720 (N_7720,N_6840,N_6474);
nor U7721 (N_7721,N_6600,N_7435);
or U7722 (N_7722,N_6345,N_7334);
xnor U7723 (N_7723,N_6348,N_7341);
xor U7724 (N_7724,N_7176,N_7479);
nor U7725 (N_7725,N_6141,N_6892);
or U7726 (N_7726,N_6094,N_6122);
xor U7727 (N_7727,N_6516,N_7011);
nor U7728 (N_7728,N_7088,N_6081);
and U7729 (N_7729,N_6686,N_6292);
nand U7730 (N_7730,N_6026,N_6050);
or U7731 (N_7731,N_6527,N_6042);
nand U7732 (N_7732,N_6339,N_6280);
nor U7733 (N_7733,N_6398,N_7179);
nand U7734 (N_7734,N_6139,N_6854);
and U7735 (N_7735,N_6216,N_6116);
and U7736 (N_7736,N_7001,N_7119);
and U7737 (N_7737,N_7335,N_6211);
nor U7738 (N_7738,N_7474,N_6573);
or U7739 (N_7739,N_6812,N_6575);
or U7740 (N_7740,N_6748,N_6917);
xor U7741 (N_7741,N_6149,N_7161);
nor U7742 (N_7742,N_7346,N_7007);
xor U7743 (N_7743,N_6134,N_7370);
nand U7744 (N_7744,N_6918,N_6349);
nor U7745 (N_7745,N_7353,N_6039);
or U7746 (N_7746,N_7010,N_6682);
or U7747 (N_7747,N_7483,N_6112);
or U7748 (N_7748,N_6981,N_6513);
xnor U7749 (N_7749,N_6145,N_6035);
xor U7750 (N_7750,N_6906,N_7433);
and U7751 (N_7751,N_7138,N_6842);
nand U7752 (N_7752,N_7359,N_7031);
nand U7753 (N_7753,N_6240,N_6721);
nand U7754 (N_7754,N_7005,N_7049);
nor U7755 (N_7755,N_6517,N_6483);
nand U7756 (N_7756,N_6327,N_7135);
nor U7757 (N_7757,N_6874,N_7365);
nand U7758 (N_7758,N_6895,N_6767);
nor U7759 (N_7759,N_6153,N_6818);
nor U7760 (N_7760,N_6872,N_6552);
or U7761 (N_7761,N_6002,N_6828);
xnor U7762 (N_7762,N_6233,N_6925);
nand U7763 (N_7763,N_6468,N_7072);
nor U7764 (N_7764,N_6864,N_7080);
and U7765 (N_7765,N_6250,N_7356);
nand U7766 (N_7766,N_7101,N_6855);
or U7767 (N_7767,N_7196,N_6941);
nor U7768 (N_7768,N_7407,N_6378);
nor U7769 (N_7769,N_6032,N_7026);
nor U7770 (N_7770,N_6921,N_7440);
nand U7771 (N_7771,N_7339,N_7307);
and U7772 (N_7772,N_6034,N_6598);
or U7773 (N_7773,N_7432,N_6067);
xor U7774 (N_7774,N_6596,N_6316);
or U7775 (N_7775,N_6863,N_6628);
nand U7776 (N_7776,N_6375,N_6219);
nor U7777 (N_7777,N_6845,N_6655);
nor U7778 (N_7778,N_6528,N_6315);
nor U7779 (N_7779,N_6866,N_6608);
xor U7780 (N_7780,N_6037,N_6498);
or U7781 (N_7781,N_6756,N_6358);
and U7782 (N_7782,N_6318,N_6113);
nor U7783 (N_7783,N_6425,N_6271);
and U7784 (N_7784,N_6341,N_7073);
and U7785 (N_7785,N_6105,N_7058);
or U7786 (N_7786,N_7423,N_7442);
nand U7787 (N_7787,N_6481,N_7489);
and U7788 (N_7788,N_7373,N_6441);
or U7789 (N_7789,N_7038,N_7484);
nand U7790 (N_7790,N_7083,N_7042);
or U7791 (N_7791,N_7250,N_6401);
xor U7792 (N_7792,N_6869,N_6813);
or U7793 (N_7793,N_6388,N_6248);
and U7794 (N_7794,N_6806,N_6181);
and U7795 (N_7795,N_7465,N_6953);
and U7796 (N_7796,N_6915,N_6296);
nand U7797 (N_7797,N_6213,N_6229);
and U7798 (N_7798,N_7168,N_6760);
xnor U7799 (N_7799,N_6352,N_7475);
nand U7800 (N_7800,N_6410,N_7397);
xnor U7801 (N_7801,N_7152,N_7284);
nand U7802 (N_7802,N_6619,N_7309);
nor U7803 (N_7803,N_6151,N_6805);
and U7804 (N_7804,N_6750,N_6902);
or U7805 (N_7805,N_7280,N_6846);
nand U7806 (N_7806,N_6547,N_7143);
or U7807 (N_7807,N_6432,N_7270);
xor U7808 (N_7808,N_7175,N_7288);
and U7809 (N_7809,N_6529,N_6260);
xor U7810 (N_7810,N_6691,N_6636);
or U7811 (N_7811,N_6893,N_6765);
or U7812 (N_7812,N_6537,N_6587);
or U7813 (N_7813,N_7410,N_7102);
nor U7814 (N_7814,N_6254,N_6165);
and U7815 (N_7815,N_6954,N_6275);
and U7816 (N_7816,N_7227,N_7220);
and U7817 (N_7817,N_7204,N_7470);
and U7818 (N_7818,N_6551,N_7069);
nand U7819 (N_7819,N_7064,N_6265);
nor U7820 (N_7820,N_6685,N_7251);
xnor U7821 (N_7821,N_6572,N_6399);
nor U7822 (N_7822,N_7447,N_6819);
nand U7823 (N_7823,N_6195,N_7043);
nor U7824 (N_7824,N_7467,N_6012);
nand U7825 (N_7825,N_7385,N_7441);
nand U7826 (N_7826,N_6850,N_6473);
and U7827 (N_7827,N_6423,N_6783);
nand U7828 (N_7828,N_7236,N_6733);
xnor U7829 (N_7829,N_7303,N_6777);
nor U7830 (N_7830,N_6966,N_7488);
nor U7831 (N_7831,N_6290,N_6983);
xor U7832 (N_7832,N_7490,N_6770);
nand U7833 (N_7833,N_6647,N_7154);
xnor U7834 (N_7834,N_7430,N_7369);
xor U7835 (N_7835,N_7178,N_6835);
nor U7836 (N_7836,N_7332,N_6713);
xnor U7837 (N_7837,N_7311,N_6159);
nand U7838 (N_7838,N_7312,N_6643);
nor U7839 (N_7839,N_7252,N_6903);
nor U7840 (N_7840,N_6540,N_7287);
and U7841 (N_7841,N_7318,N_7140);
or U7842 (N_7842,N_6063,N_7019);
or U7843 (N_7843,N_6694,N_6415);
and U7844 (N_7844,N_6973,N_7194);
and U7845 (N_7845,N_7103,N_7225);
xnor U7846 (N_7846,N_6782,N_7106);
xnor U7847 (N_7847,N_6909,N_6146);
and U7848 (N_7848,N_6875,N_6933);
and U7849 (N_7849,N_7231,N_6871);
or U7850 (N_7850,N_6019,N_6993);
and U7851 (N_7851,N_6945,N_6272);
and U7852 (N_7852,N_6757,N_6104);
and U7853 (N_7853,N_6987,N_6776);
nand U7854 (N_7854,N_7009,N_6877);
and U7855 (N_7855,N_6308,N_6431);
and U7856 (N_7856,N_7067,N_6914);
and U7857 (N_7857,N_7446,N_6952);
and U7858 (N_7858,N_7482,N_6972);
nor U7859 (N_7859,N_6471,N_6654);
nor U7860 (N_7860,N_7491,N_6442);
nor U7861 (N_7861,N_6958,N_6381);
or U7862 (N_7862,N_6762,N_6898);
xnor U7863 (N_7863,N_6743,N_6166);
nand U7864 (N_7864,N_7315,N_7444);
xnor U7865 (N_7865,N_6365,N_6144);
nor U7866 (N_7866,N_6025,N_6380);
and U7867 (N_7867,N_7317,N_6383);
nand U7868 (N_7868,N_6332,N_6482);
nor U7869 (N_7869,N_6659,N_6011);
nor U7870 (N_7870,N_6095,N_7223);
or U7871 (N_7871,N_7381,N_7338);
or U7872 (N_7872,N_7481,N_7221);
nand U7873 (N_7873,N_6413,N_6653);
and U7874 (N_7874,N_6744,N_6058);
nand U7875 (N_7875,N_6087,N_6924);
xor U7876 (N_7876,N_6640,N_6257);
xnor U7877 (N_7877,N_6464,N_7020);
xor U7878 (N_7878,N_6089,N_6553);
and U7879 (N_7879,N_7025,N_6695);
xor U7880 (N_7880,N_6489,N_6559);
or U7881 (N_7881,N_6960,N_7077);
nand U7882 (N_7882,N_7224,N_6884);
nand U7883 (N_7883,N_6405,N_6448);
or U7884 (N_7884,N_6461,N_7322);
nand U7885 (N_7885,N_6810,N_7003);
and U7886 (N_7886,N_6997,N_7434);
xnor U7887 (N_7887,N_7187,N_6809);
and U7888 (N_7888,N_6717,N_6652);
and U7889 (N_7889,N_6604,N_7478);
nor U7890 (N_7890,N_7272,N_7008);
and U7891 (N_7891,N_7492,N_6060);
nor U7892 (N_7892,N_7345,N_6992);
xor U7893 (N_7893,N_7343,N_6157);
xnor U7894 (N_7894,N_6963,N_6671);
and U7895 (N_7895,N_7401,N_6199);
and U7896 (N_7896,N_7253,N_6831);
nand U7897 (N_7897,N_7411,N_6673);
xor U7898 (N_7898,N_7240,N_6672);
nor U7899 (N_7899,N_6268,N_7361);
and U7900 (N_7900,N_6560,N_6579);
or U7901 (N_7901,N_6775,N_6436);
nand U7902 (N_7902,N_7241,N_7275);
xnor U7903 (N_7903,N_7495,N_6725);
or U7904 (N_7904,N_6662,N_6076);
or U7905 (N_7905,N_6397,N_7342);
and U7906 (N_7906,N_7459,N_7153);
and U7907 (N_7907,N_7471,N_6539);
and U7908 (N_7908,N_6133,N_7055);
nand U7909 (N_7909,N_7166,N_7093);
nand U7910 (N_7910,N_6276,N_6407);
nor U7911 (N_7911,N_7296,N_6754);
or U7912 (N_7912,N_6131,N_6930);
and U7913 (N_7913,N_6826,N_7463);
xnor U7914 (N_7914,N_6377,N_6526);
nand U7915 (N_7915,N_7278,N_7405);
nand U7916 (N_7916,N_6848,N_7213);
and U7917 (N_7917,N_7476,N_6834);
xnor U7918 (N_7918,N_6355,N_7367);
nor U7919 (N_7919,N_6251,N_7214);
nor U7920 (N_7920,N_7222,N_6521);
nand U7921 (N_7921,N_6041,N_6439);
or U7922 (N_7922,N_6180,N_7039);
or U7923 (N_7923,N_7232,N_6043);
xor U7924 (N_7924,N_6799,N_6130);
nand U7925 (N_7925,N_6261,N_6974);
and U7926 (N_7926,N_7243,N_6601);
nand U7927 (N_7927,N_6561,N_6677);
nor U7928 (N_7928,N_7328,N_7233);
and U7929 (N_7929,N_6245,N_6198);
or U7930 (N_7930,N_6665,N_6690);
and U7931 (N_7931,N_7129,N_6668);
or U7932 (N_7932,N_6338,N_6989);
nor U7933 (N_7933,N_6800,N_6028);
and U7934 (N_7934,N_6545,N_6475);
xnor U7935 (N_7935,N_7121,N_6716);
xor U7936 (N_7936,N_7066,N_6302);
nand U7937 (N_7937,N_6645,N_7095);
or U7938 (N_7938,N_6753,N_6667);
nor U7939 (N_7939,N_6001,N_6617);
nor U7940 (N_7940,N_6183,N_7414);
nor U7941 (N_7941,N_6644,N_6900);
or U7942 (N_7942,N_6207,N_6571);
nand U7943 (N_7943,N_6269,N_6699);
nor U7944 (N_7944,N_6961,N_6763);
xnor U7945 (N_7945,N_7136,N_6170);
xor U7946 (N_7946,N_6386,N_6350);
or U7947 (N_7947,N_6137,N_6533);
nor U7948 (N_7948,N_6907,N_7183);
xor U7949 (N_7949,N_7404,N_7412);
and U7950 (N_7950,N_6724,N_6555);
and U7951 (N_7951,N_6356,N_7294);
nor U7952 (N_7952,N_6847,N_6304);
xor U7953 (N_7953,N_6052,N_7499);
and U7954 (N_7954,N_6340,N_7281);
nand U7955 (N_7955,N_6156,N_7389);
xor U7956 (N_7956,N_6947,N_6920);
or U7957 (N_7957,N_7388,N_6215);
xor U7958 (N_7958,N_6908,N_6886);
and U7959 (N_7959,N_7081,N_7305);
or U7960 (N_7960,N_6990,N_6047);
xnor U7961 (N_7961,N_7190,N_6752);
xnor U7962 (N_7962,N_6202,N_7260);
or U7963 (N_7963,N_6808,N_6922);
and U7964 (N_7964,N_6520,N_7028);
and U7965 (N_7965,N_6445,N_7417);
nand U7966 (N_7966,N_7092,N_6698);
or U7967 (N_7967,N_6135,N_6798);
nor U7968 (N_7968,N_6710,N_6231);
xor U7969 (N_7969,N_6451,N_6715);
xor U7970 (N_7970,N_6683,N_7012);
and U7971 (N_7971,N_6299,N_6074);
and U7972 (N_7972,N_7274,N_6512);
or U7973 (N_7973,N_6719,N_6285);
and U7974 (N_7974,N_6658,N_7256);
or U7975 (N_7975,N_6581,N_6117);
xnor U7976 (N_7976,N_6224,N_6367);
nand U7977 (N_7977,N_6549,N_6168);
xor U7978 (N_7978,N_7357,N_6968);
nand U7979 (N_7979,N_6472,N_6485);
and U7980 (N_7980,N_6253,N_7466);
nor U7981 (N_7981,N_7000,N_6478);
and U7982 (N_7982,N_6576,N_7394);
and U7983 (N_7983,N_7052,N_6538);
and U7984 (N_7984,N_6031,N_6488);
nand U7985 (N_7985,N_7228,N_7379);
and U7986 (N_7986,N_6546,N_6228);
nor U7987 (N_7987,N_6396,N_7126);
nor U7988 (N_7988,N_7298,N_6051);
or U7989 (N_7989,N_7165,N_6194);
nor U7990 (N_7990,N_7306,N_6241);
and U7991 (N_7991,N_6554,N_6297);
xnor U7992 (N_7992,N_6362,N_7099);
xor U7993 (N_7993,N_6373,N_6346);
or U7994 (N_7994,N_6258,N_6631);
and U7995 (N_7995,N_6294,N_6230);
and U7996 (N_7996,N_7351,N_6940);
nand U7997 (N_7997,N_6676,N_7291);
xor U7998 (N_7998,N_6114,N_6023);
and U7999 (N_7999,N_7383,N_6204);
nand U8000 (N_8000,N_7059,N_6084);
and U8001 (N_8001,N_7034,N_6802);
and U8002 (N_8002,N_6328,N_7244);
nor U8003 (N_8003,N_7452,N_6603);
xnor U8004 (N_8004,N_7205,N_7195);
nor U8005 (N_8005,N_7191,N_7498);
xor U8006 (N_8006,N_6896,N_7413);
or U8007 (N_8007,N_6861,N_6544);
xor U8008 (N_8008,N_6995,N_7124);
and U8009 (N_8009,N_6580,N_7340);
nand U8010 (N_8010,N_7217,N_7046);
nor U8011 (N_8011,N_6469,N_6243);
or U8012 (N_8012,N_6242,N_6161);
or U8013 (N_8013,N_6656,N_6996);
nand U8014 (N_8014,N_6881,N_6008);
and U8015 (N_8015,N_7246,N_6179);
or U8016 (N_8016,N_6509,N_6792);
nand U8017 (N_8017,N_6780,N_6978);
and U8018 (N_8018,N_6279,N_7308);
nand U8019 (N_8019,N_7146,N_7144);
nand U8020 (N_8020,N_6639,N_6556);
nor U8021 (N_8021,N_7044,N_7493);
and U8022 (N_8022,N_7050,N_6811);
or U8023 (N_8023,N_7115,N_6077);
and U8024 (N_8024,N_7419,N_7167);
or U8025 (N_8025,N_6817,N_6994);
nor U8026 (N_8026,N_7118,N_7130);
nor U8027 (N_8027,N_6635,N_7047);
and U8028 (N_8028,N_7211,N_6624);
nor U8029 (N_8029,N_7424,N_6623);
or U8030 (N_8030,N_6192,N_6862);
nand U8031 (N_8031,N_6735,N_7203);
and U8032 (N_8032,N_6045,N_6107);
and U8033 (N_8033,N_6057,N_6344);
and U8034 (N_8034,N_7487,N_6206);
and U8035 (N_8035,N_7090,N_6928);
xnor U8036 (N_8036,N_6621,N_6226);
nand U8037 (N_8037,N_7358,N_6409);
or U8038 (N_8038,N_6438,N_6370);
xnor U8039 (N_8039,N_7457,N_6946);
and U8040 (N_8040,N_6788,N_7386);
nor U8041 (N_8041,N_6880,N_6742);
nand U8042 (N_8042,N_7408,N_6324);
xnor U8043 (N_8043,N_7127,N_6360);
or U8044 (N_8044,N_6177,N_6395);
nor U8045 (N_8045,N_6988,N_7006);
and U8046 (N_8046,N_7087,N_7114);
nand U8047 (N_8047,N_6416,N_6123);
and U8048 (N_8048,N_7300,N_7209);
nand U8049 (N_8049,N_6259,N_7387);
or U8050 (N_8050,N_7156,N_6320);
and U8051 (N_8051,N_6849,N_7436);
nor U8052 (N_8052,N_6761,N_6121);
or U8053 (N_8053,N_6480,N_7045);
nor U8054 (N_8054,N_6463,N_7094);
nand U8055 (N_8055,N_7431,N_7238);
or U8056 (N_8056,N_6205,N_6882);
nor U8057 (N_8057,N_6033,N_7473);
or U8058 (N_8058,N_6209,N_6689);
nand U8059 (N_8059,N_6171,N_6883);
nand U8060 (N_8060,N_6838,N_6148);
xnor U8061 (N_8061,N_6916,N_7125);
or U8062 (N_8062,N_7258,N_6078);
or U8063 (N_8063,N_7259,N_7409);
and U8064 (N_8064,N_6522,N_6565);
xor U8065 (N_8065,N_6678,N_6079);
nor U8066 (N_8066,N_7071,N_7468);
nand U8067 (N_8067,N_6036,N_6091);
xnor U8068 (N_8068,N_6428,N_7076);
nand U8069 (N_8069,N_6570,N_6614);
and U8070 (N_8070,N_7016,N_6402);
and U8071 (N_8071,N_6163,N_6669);
nor U8072 (N_8072,N_6563,N_7189);
or U8073 (N_8073,N_6232,N_6429);
nor U8074 (N_8074,N_7033,N_6126);
nor U8075 (N_8075,N_7393,N_7014);
and U8076 (N_8076,N_6066,N_6629);
and U8077 (N_8077,N_6615,N_7276);
nand U8078 (N_8078,N_7024,N_7344);
and U8079 (N_8079,N_7041,N_6333);
xor U8080 (N_8080,N_6082,N_6295);
nand U8081 (N_8081,N_7450,N_6300);
nor U8082 (N_8082,N_7486,N_6586);
nor U8083 (N_8083,N_6330,N_7237);
nand U8084 (N_8084,N_6680,N_6382);
nor U8085 (N_8085,N_6307,N_6086);
nor U8086 (N_8086,N_6859,N_6068);
or U8087 (N_8087,N_7133,N_7173);
xnor U8088 (N_8088,N_7174,N_6499);
nor U8089 (N_8089,N_6193,N_7363);
and U8090 (N_8090,N_7053,N_6317);
or U8091 (N_8091,N_7319,N_7200);
nor U8092 (N_8092,N_6759,N_7113);
nand U8093 (N_8093,N_6731,N_6329);
or U8094 (N_8094,N_7037,N_6939);
nor U8095 (N_8095,N_6929,N_6969);
or U8096 (N_8096,N_6837,N_7390);
and U8097 (N_8097,N_6923,N_7206);
nand U8098 (N_8098,N_7268,N_7263);
nand U8099 (N_8099,N_6949,N_6176);
and U8100 (N_8100,N_6562,N_6004);
nor U8101 (N_8101,N_6097,N_7439);
nand U8102 (N_8102,N_7428,N_7068);
and U8103 (N_8103,N_6102,N_7329);
and U8104 (N_8104,N_6827,N_7290);
xnor U8105 (N_8105,N_6418,N_6470);
nor U8106 (N_8106,N_7060,N_6768);
nand U8107 (N_8107,N_6664,N_6392);
nand U8108 (N_8108,N_6789,N_6557);
xnor U8109 (N_8109,N_6444,N_7070);
xnor U8110 (N_8110,N_6288,N_6247);
or U8111 (N_8111,N_7472,N_6160);
or U8112 (N_8112,N_6524,N_7349);
nor U8113 (N_8113,N_6891,N_6433);
and U8114 (N_8114,N_6143,N_6795);
and U8115 (N_8115,N_7202,N_6870);
nand U8116 (N_8116,N_6426,N_6998);
nand U8117 (N_8117,N_6740,N_6453);
and U8118 (N_8118,N_7207,N_6406);
nand U8119 (N_8119,N_7180,N_6734);
or U8120 (N_8120,N_7497,N_6027);
nand U8121 (N_8121,N_6508,N_7364);
xnor U8122 (N_8122,N_7304,N_7027);
nor U8123 (N_8123,N_6459,N_6956);
nand U8124 (N_8124,N_6289,N_7378);
or U8125 (N_8125,N_7085,N_7193);
nor U8126 (N_8126,N_6638,N_7350);
xor U8127 (N_8127,N_6642,N_7215);
xor U8128 (N_8128,N_6885,N_7416);
nand U8129 (N_8129,N_6730,N_6164);
nor U8130 (N_8130,N_6391,N_6801);
nand U8131 (N_8131,N_7151,N_6525);
or U8132 (N_8132,N_6590,N_6634);
nor U8133 (N_8133,N_6372,N_7239);
xnor U8134 (N_8134,N_6749,N_7299);
xor U8135 (N_8135,N_6003,N_7354);
nand U8136 (N_8136,N_6950,N_6379);
and U8137 (N_8137,N_7163,N_7403);
nand U8138 (N_8138,N_7245,N_6208);
and U8139 (N_8139,N_7248,N_7286);
and U8140 (N_8140,N_6411,N_6106);
and U8141 (N_8141,N_6128,N_7171);
or U8142 (N_8142,N_6494,N_7212);
and U8143 (N_8143,N_6221,N_7426);
nand U8144 (N_8144,N_6424,N_6447);
xor U8145 (N_8145,N_6853,N_6507);
or U8146 (N_8146,N_6493,N_6147);
or U8147 (N_8147,N_6778,N_6222);
nor U8148 (N_8148,N_6310,N_6061);
nand U8149 (N_8149,N_7480,N_6606);
nand U8150 (N_8150,N_6010,N_6486);
nor U8151 (N_8151,N_6351,N_6660);
or U8152 (N_8152,N_7170,N_7096);
xor U8153 (N_8153,N_7295,N_6651);
xor U8154 (N_8154,N_6427,N_6394);
xnor U8155 (N_8155,N_6999,N_7265);
nor U8156 (N_8156,N_6616,N_7485);
xor U8157 (N_8157,N_6403,N_6359);
or U8158 (N_8158,N_7316,N_6979);
nor U8159 (N_8159,N_6017,N_6523);
and U8160 (N_8160,N_7022,N_6430);
and U8161 (N_8161,N_6707,N_7454);
or U8162 (N_8162,N_6585,N_7021);
nand U8163 (N_8163,N_6706,N_6807);
xor U8164 (N_8164,N_6408,N_6938);
and U8165 (N_8165,N_6936,N_6040);
nand U8166 (N_8166,N_7181,N_6975);
nand U8167 (N_8167,N_6736,N_7029);
xnor U8168 (N_8168,N_7422,N_6944);
nand U8169 (N_8169,N_6784,N_6342);
xor U8170 (N_8170,N_6632,N_6910);
nor U8171 (N_8171,N_7229,N_6256);
or U8172 (N_8172,N_6718,N_6927);
or U8173 (N_8173,N_6321,N_6007);
and U8174 (N_8174,N_6305,N_6006);
or U8175 (N_8175,N_6142,N_7347);
xnor U8176 (N_8176,N_6622,N_6088);
xnor U8177 (N_8177,N_7109,N_6080);
or U8178 (N_8178,N_6535,N_6108);
nor U8179 (N_8179,N_6024,N_7399);
xor U8180 (N_8180,N_7086,N_6353);
nor U8181 (N_8181,N_6926,N_7271);
xor U8182 (N_8182,N_6385,N_6479);
or U8183 (N_8183,N_6303,N_6856);
and U8184 (N_8184,N_6738,N_7324);
nor U8185 (N_8185,N_6460,N_6069);
nor U8186 (N_8186,N_6865,N_6274);
nor U8187 (N_8187,N_6700,N_6477);
and U8188 (N_8188,N_6720,N_6054);
and U8189 (N_8189,N_7293,N_6774);
nand U8190 (N_8190,N_6543,N_6118);
or U8191 (N_8191,N_7366,N_6457);
nand U8192 (N_8192,N_6465,N_6127);
or U8193 (N_8193,N_7247,N_6322);
nand U8194 (N_8194,N_7331,N_6013);
and U8195 (N_8195,N_6491,N_6110);
nand U8196 (N_8196,N_6000,N_6577);
xor U8197 (N_8197,N_7141,N_6029);
or U8198 (N_8198,N_7297,N_6178);
nand U8199 (N_8199,N_6705,N_6701);
and U8200 (N_8200,N_6714,N_6935);
and U8201 (N_8201,N_7210,N_6919);
xor U8202 (N_8202,N_6186,N_6791);
or U8203 (N_8203,N_6167,N_6649);
nor U8204 (N_8204,N_6083,N_6009);
xnor U8205 (N_8205,N_6158,N_6476);
or U8206 (N_8206,N_7030,N_6786);
nor U8207 (N_8207,N_6897,N_7089);
xnor U8208 (N_8208,N_6191,N_7018);
and U8209 (N_8209,N_7218,N_7100);
xor U8210 (N_8210,N_7249,N_7062);
nand U8211 (N_8211,N_6737,N_7313);
or U8212 (N_8212,N_6879,N_6187);
nand U8213 (N_8213,N_6293,N_7400);
or U8214 (N_8214,N_7396,N_6400);
nand U8215 (N_8215,N_6518,N_6709);
nor U8216 (N_8216,N_6100,N_6739);
xnor U8217 (N_8217,N_6982,N_6075);
and U8218 (N_8218,N_6728,N_6287);
nor U8219 (N_8219,N_6531,N_7160);
xnor U8220 (N_8220,N_7461,N_6172);
xnor U8221 (N_8221,N_6337,N_6589);
and U8222 (N_8222,N_6578,N_6173);
nor U8223 (N_8223,N_6773,N_7186);
or U8224 (N_8224,N_6201,N_6090);
or U8225 (N_8225,N_7230,N_6217);
nor U8226 (N_8226,N_6959,N_6334);
or U8227 (N_8227,N_6888,N_6542);
nor U8228 (N_8228,N_6210,N_6015);
or U8229 (N_8229,N_6197,N_6726);
nor U8230 (N_8230,N_6237,N_6977);
nor U8231 (N_8231,N_7098,N_6282);
nand U8232 (N_8232,N_6824,N_7421);
nand U8233 (N_8233,N_6970,N_7116);
and U8234 (N_8234,N_7192,N_7283);
nand U8235 (N_8235,N_6708,N_7395);
xnor U8236 (N_8236,N_7137,N_6152);
nand U8237 (N_8237,N_7323,N_6437);
nand U8238 (N_8238,N_6836,N_6887);
nand U8239 (N_8239,N_6214,N_6417);
nor U8240 (N_8240,N_7438,N_7326);
nor U8241 (N_8241,N_6155,N_6422);
nand U8242 (N_8242,N_7257,N_7406);
nand U8243 (N_8243,N_6504,N_6154);
nor U8244 (N_8244,N_6096,N_6374);
nand U8245 (N_8245,N_6188,N_6119);
or U8246 (N_8246,N_7456,N_6785);
nor U8247 (N_8247,N_7051,N_6605);
nor U8248 (N_8248,N_6932,N_6018);
xor U8249 (N_8249,N_6283,N_6419);
nor U8250 (N_8250,N_6183,N_6505);
and U8251 (N_8251,N_6340,N_6627);
or U8252 (N_8252,N_7138,N_7210);
and U8253 (N_8253,N_6738,N_7410);
nor U8254 (N_8254,N_6287,N_7085);
xnor U8255 (N_8255,N_6901,N_6425);
and U8256 (N_8256,N_6717,N_6207);
and U8257 (N_8257,N_6393,N_7437);
xnor U8258 (N_8258,N_6599,N_6054);
xor U8259 (N_8259,N_7004,N_7037);
xor U8260 (N_8260,N_6774,N_7235);
nor U8261 (N_8261,N_6861,N_6532);
or U8262 (N_8262,N_6194,N_7437);
nand U8263 (N_8263,N_6582,N_6323);
nand U8264 (N_8264,N_7108,N_6977);
or U8265 (N_8265,N_7466,N_6216);
nand U8266 (N_8266,N_7180,N_7086);
and U8267 (N_8267,N_6921,N_6924);
and U8268 (N_8268,N_6291,N_6224);
and U8269 (N_8269,N_6543,N_7203);
or U8270 (N_8270,N_6889,N_6178);
xor U8271 (N_8271,N_6538,N_6360);
and U8272 (N_8272,N_7102,N_6931);
xor U8273 (N_8273,N_6937,N_6093);
nand U8274 (N_8274,N_6787,N_6858);
or U8275 (N_8275,N_6655,N_7259);
nand U8276 (N_8276,N_6365,N_6765);
and U8277 (N_8277,N_6660,N_6790);
or U8278 (N_8278,N_6041,N_7361);
nand U8279 (N_8279,N_7172,N_7343);
or U8280 (N_8280,N_6969,N_6109);
nor U8281 (N_8281,N_6557,N_6172);
xor U8282 (N_8282,N_6688,N_6106);
or U8283 (N_8283,N_6903,N_6139);
or U8284 (N_8284,N_6806,N_6150);
nand U8285 (N_8285,N_6355,N_6690);
nand U8286 (N_8286,N_7315,N_6644);
and U8287 (N_8287,N_6302,N_6742);
or U8288 (N_8288,N_6730,N_7408);
and U8289 (N_8289,N_6831,N_6718);
nand U8290 (N_8290,N_6606,N_6705);
nor U8291 (N_8291,N_6790,N_7110);
and U8292 (N_8292,N_6521,N_6041);
nand U8293 (N_8293,N_6445,N_6322);
xnor U8294 (N_8294,N_7483,N_6366);
nand U8295 (N_8295,N_6528,N_6614);
nand U8296 (N_8296,N_6125,N_7213);
nor U8297 (N_8297,N_6801,N_6404);
or U8298 (N_8298,N_6930,N_7317);
xnor U8299 (N_8299,N_7026,N_6845);
nand U8300 (N_8300,N_6223,N_6464);
nand U8301 (N_8301,N_6257,N_7268);
nand U8302 (N_8302,N_6930,N_7219);
nand U8303 (N_8303,N_7383,N_6269);
xor U8304 (N_8304,N_6955,N_7238);
and U8305 (N_8305,N_6014,N_6897);
xor U8306 (N_8306,N_6823,N_6046);
xnor U8307 (N_8307,N_6004,N_7393);
nand U8308 (N_8308,N_6883,N_7457);
and U8309 (N_8309,N_6644,N_7433);
nand U8310 (N_8310,N_7393,N_7305);
or U8311 (N_8311,N_7284,N_6430);
and U8312 (N_8312,N_6184,N_6895);
and U8313 (N_8313,N_6487,N_6326);
or U8314 (N_8314,N_7178,N_6040);
nand U8315 (N_8315,N_6368,N_7279);
nand U8316 (N_8316,N_6728,N_7232);
or U8317 (N_8317,N_7156,N_6599);
and U8318 (N_8318,N_6725,N_6146);
and U8319 (N_8319,N_7480,N_7433);
xnor U8320 (N_8320,N_7191,N_7192);
or U8321 (N_8321,N_6721,N_6541);
nor U8322 (N_8322,N_6182,N_7011);
nor U8323 (N_8323,N_6328,N_7373);
nor U8324 (N_8324,N_6270,N_6736);
or U8325 (N_8325,N_6571,N_6099);
or U8326 (N_8326,N_6052,N_7239);
and U8327 (N_8327,N_7028,N_6333);
xor U8328 (N_8328,N_7352,N_7440);
nor U8329 (N_8329,N_6522,N_7160);
xor U8330 (N_8330,N_7259,N_6847);
and U8331 (N_8331,N_7098,N_6913);
nand U8332 (N_8332,N_6244,N_6924);
nor U8333 (N_8333,N_6761,N_7421);
nor U8334 (N_8334,N_6643,N_6328);
and U8335 (N_8335,N_7207,N_7423);
xnor U8336 (N_8336,N_6770,N_7095);
nor U8337 (N_8337,N_6956,N_6550);
nor U8338 (N_8338,N_6631,N_7300);
nor U8339 (N_8339,N_7414,N_6940);
and U8340 (N_8340,N_6996,N_6915);
nand U8341 (N_8341,N_6792,N_7284);
or U8342 (N_8342,N_6589,N_6366);
and U8343 (N_8343,N_6752,N_7224);
and U8344 (N_8344,N_6408,N_7073);
nor U8345 (N_8345,N_6422,N_7284);
nand U8346 (N_8346,N_6324,N_6569);
or U8347 (N_8347,N_6384,N_7497);
xnor U8348 (N_8348,N_7110,N_6366);
or U8349 (N_8349,N_7277,N_6732);
xnor U8350 (N_8350,N_6574,N_6275);
and U8351 (N_8351,N_7467,N_6385);
and U8352 (N_8352,N_6300,N_6856);
nor U8353 (N_8353,N_6654,N_6975);
xor U8354 (N_8354,N_6121,N_6472);
and U8355 (N_8355,N_6235,N_6176);
nor U8356 (N_8356,N_6640,N_6700);
and U8357 (N_8357,N_6270,N_6677);
or U8358 (N_8358,N_6675,N_6301);
nand U8359 (N_8359,N_6112,N_6146);
nor U8360 (N_8360,N_6349,N_7362);
nand U8361 (N_8361,N_7310,N_7048);
xor U8362 (N_8362,N_6641,N_6609);
nor U8363 (N_8363,N_7185,N_6671);
nor U8364 (N_8364,N_7365,N_6634);
xnor U8365 (N_8365,N_6043,N_6051);
and U8366 (N_8366,N_6603,N_7364);
xor U8367 (N_8367,N_6540,N_6989);
nor U8368 (N_8368,N_6013,N_6682);
nand U8369 (N_8369,N_7227,N_6218);
or U8370 (N_8370,N_6130,N_6892);
nor U8371 (N_8371,N_7355,N_7479);
or U8372 (N_8372,N_6139,N_6727);
nand U8373 (N_8373,N_7128,N_6798);
nand U8374 (N_8374,N_6611,N_6605);
xor U8375 (N_8375,N_6849,N_7489);
nor U8376 (N_8376,N_6172,N_6185);
xnor U8377 (N_8377,N_6330,N_7482);
and U8378 (N_8378,N_6575,N_6600);
nor U8379 (N_8379,N_6512,N_6345);
nor U8380 (N_8380,N_6760,N_6694);
nand U8381 (N_8381,N_6233,N_6491);
nor U8382 (N_8382,N_6530,N_7273);
nor U8383 (N_8383,N_6551,N_6539);
and U8384 (N_8384,N_6426,N_7073);
nand U8385 (N_8385,N_6302,N_7478);
or U8386 (N_8386,N_7347,N_6138);
and U8387 (N_8387,N_6581,N_7217);
nor U8388 (N_8388,N_7499,N_6237);
nor U8389 (N_8389,N_6802,N_6318);
nand U8390 (N_8390,N_6379,N_6916);
or U8391 (N_8391,N_7267,N_6001);
xor U8392 (N_8392,N_7192,N_6353);
xor U8393 (N_8393,N_6336,N_6755);
or U8394 (N_8394,N_6513,N_6047);
nand U8395 (N_8395,N_6018,N_6965);
xnor U8396 (N_8396,N_6181,N_7451);
nor U8397 (N_8397,N_6003,N_6910);
nor U8398 (N_8398,N_7495,N_6091);
or U8399 (N_8399,N_6676,N_6819);
or U8400 (N_8400,N_6827,N_7137);
and U8401 (N_8401,N_7050,N_6667);
or U8402 (N_8402,N_6227,N_7284);
xnor U8403 (N_8403,N_7376,N_6607);
or U8404 (N_8404,N_6852,N_6514);
xnor U8405 (N_8405,N_6250,N_6903);
nand U8406 (N_8406,N_6793,N_6133);
nand U8407 (N_8407,N_7301,N_7211);
and U8408 (N_8408,N_6301,N_6618);
xnor U8409 (N_8409,N_7406,N_7385);
and U8410 (N_8410,N_6190,N_6084);
nand U8411 (N_8411,N_6007,N_6851);
or U8412 (N_8412,N_7022,N_6303);
or U8413 (N_8413,N_7055,N_6980);
nor U8414 (N_8414,N_7153,N_7225);
nor U8415 (N_8415,N_7196,N_6344);
or U8416 (N_8416,N_7183,N_6232);
and U8417 (N_8417,N_7169,N_6162);
and U8418 (N_8418,N_6561,N_7276);
nor U8419 (N_8419,N_6228,N_6165);
and U8420 (N_8420,N_6297,N_6408);
or U8421 (N_8421,N_6983,N_7246);
nor U8422 (N_8422,N_7136,N_7086);
nand U8423 (N_8423,N_7183,N_6705);
or U8424 (N_8424,N_6807,N_6367);
xnor U8425 (N_8425,N_6015,N_6126);
nor U8426 (N_8426,N_7372,N_7075);
and U8427 (N_8427,N_6445,N_6520);
and U8428 (N_8428,N_7133,N_7213);
nand U8429 (N_8429,N_6211,N_7223);
nand U8430 (N_8430,N_7495,N_7290);
and U8431 (N_8431,N_6006,N_6623);
and U8432 (N_8432,N_6647,N_6088);
or U8433 (N_8433,N_6396,N_6779);
nand U8434 (N_8434,N_6414,N_6251);
xnor U8435 (N_8435,N_7425,N_6548);
xor U8436 (N_8436,N_6422,N_6195);
or U8437 (N_8437,N_6255,N_7049);
xnor U8438 (N_8438,N_7179,N_6273);
and U8439 (N_8439,N_6148,N_6687);
and U8440 (N_8440,N_6157,N_7057);
xor U8441 (N_8441,N_6257,N_6759);
or U8442 (N_8442,N_6728,N_7472);
and U8443 (N_8443,N_6291,N_6960);
nand U8444 (N_8444,N_6253,N_6086);
or U8445 (N_8445,N_7391,N_6481);
xor U8446 (N_8446,N_6750,N_7117);
xor U8447 (N_8447,N_6110,N_7184);
or U8448 (N_8448,N_6245,N_6421);
nor U8449 (N_8449,N_7078,N_6537);
xor U8450 (N_8450,N_7449,N_6613);
or U8451 (N_8451,N_7372,N_6994);
nand U8452 (N_8452,N_7252,N_6019);
nor U8453 (N_8453,N_6522,N_6402);
or U8454 (N_8454,N_7061,N_7318);
nand U8455 (N_8455,N_6915,N_6687);
and U8456 (N_8456,N_6148,N_7089);
and U8457 (N_8457,N_6945,N_6282);
and U8458 (N_8458,N_7233,N_6158);
or U8459 (N_8459,N_7065,N_7191);
nand U8460 (N_8460,N_6572,N_7139);
or U8461 (N_8461,N_6582,N_7297);
nand U8462 (N_8462,N_6709,N_6584);
nor U8463 (N_8463,N_6407,N_6221);
or U8464 (N_8464,N_6466,N_6166);
nor U8465 (N_8465,N_6120,N_6376);
nand U8466 (N_8466,N_7003,N_6769);
nor U8467 (N_8467,N_7417,N_6814);
nor U8468 (N_8468,N_6274,N_7009);
or U8469 (N_8469,N_6429,N_6750);
nand U8470 (N_8470,N_6875,N_7181);
nor U8471 (N_8471,N_6271,N_6054);
or U8472 (N_8472,N_6503,N_7255);
xnor U8473 (N_8473,N_6293,N_6683);
or U8474 (N_8474,N_7224,N_6324);
xor U8475 (N_8475,N_6610,N_6044);
nor U8476 (N_8476,N_6255,N_7109);
and U8477 (N_8477,N_7203,N_6824);
xnor U8478 (N_8478,N_6531,N_6701);
nor U8479 (N_8479,N_6162,N_6398);
and U8480 (N_8480,N_6083,N_7191);
and U8481 (N_8481,N_6585,N_7301);
nand U8482 (N_8482,N_6004,N_6113);
nand U8483 (N_8483,N_6236,N_6774);
nor U8484 (N_8484,N_6973,N_6265);
xor U8485 (N_8485,N_7296,N_7002);
or U8486 (N_8486,N_7409,N_6364);
and U8487 (N_8487,N_6505,N_6467);
and U8488 (N_8488,N_6707,N_7015);
nor U8489 (N_8489,N_7122,N_6703);
or U8490 (N_8490,N_6691,N_7266);
nor U8491 (N_8491,N_7187,N_6061);
xnor U8492 (N_8492,N_7202,N_6607);
xnor U8493 (N_8493,N_7104,N_6964);
and U8494 (N_8494,N_6491,N_7270);
nor U8495 (N_8495,N_6981,N_6822);
and U8496 (N_8496,N_6076,N_7328);
xor U8497 (N_8497,N_7272,N_6877);
or U8498 (N_8498,N_6758,N_6433);
nand U8499 (N_8499,N_6539,N_7115);
nor U8500 (N_8500,N_6368,N_7261);
or U8501 (N_8501,N_6832,N_7255);
nand U8502 (N_8502,N_6532,N_6996);
nor U8503 (N_8503,N_6521,N_6893);
nor U8504 (N_8504,N_7145,N_6453);
nand U8505 (N_8505,N_6294,N_6244);
nand U8506 (N_8506,N_6497,N_6293);
or U8507 (N_8507,N_7286,N_6003);
xor U8508 (N_8508,N_6591,N_6941);
nor U8509 (N_8509,N_6743,N_6578);
or U8510 (N_8510,N_6824,N_6959);
nor U8511 (N_8511,N_7377,N_6936);
nor U8512 (N_8512,N_7132,N_7369);
xnor U8513 (N_8513,N_6851,N_6354);
nand U8514 (N_8514,N_6563,N_6987);
nor U8515 (N_8515,N_6893,N_6675);
nor U8516 (N_8516,N_6615,N_7222);
and U8517 (N_8517,N_6781,N_6032);
nor U8518 (N_8518,N_6665,N_7026);
nand U8519 (N_8519,N_7046,N_6322);
nand U8520 (N_8520,N_6447,N_6367);
nor U8521 (N_8521,N_7402,N_6569);
nor U8522 (N_8522,N_6788,N_6471);
nand U8523 (N_8523,N_7499,N_7472);
and U8524 (N_8524,N_7110,N_6750);
and U8525 (N_8525,N_7252,N_6581);
nor U8526 (N_8526,N_6886,N_7105);
xnor U8527 (N_8527,N_7104,N_6666);
nor U8528 (N_8528,N_6163,N_7136);
xor U8529 (N_8529,N_7043,N_6316);
and U8530 (N_8530,N_6074,N_6304);
and U8531 (N_8531,N_7479,N_6222);
nor U8532 (N_8532,N_6991,N_7142);
nand U8533 (N_8533,N_6782,N_6458);
and U8534 (N_8534,N_6578,N_7495);
or U8535 (N_8535,N_6266,N_6522);
nor U8536 (N_8536,N_7268,N_6555);
and U8537 (N_8537,N_6700,N_6588);
and U8538 (N_8538,N_7355,N_6661);
nand U8539 (N_8539,N_6575,N_6015);
nand U8540 (N_8540,N_7350,N_6660);
and U8541 (N_8541,N_6521,N_6647);
nand U8542 (N_8542,N_6141,N_7377);
xor U8543 (N_8543,N_6787,N_6888);
nor U8544 (N_8544,N_7087,N_6171);
and U8545 (N_8545,N_6134,N_6379);
xor U8546 (N_8546,N_6035,N_6046);
xor U8547 (N_8547,N_7124,N_6109);
nor U8548 (N_8548,N_7123,N_7368);
or U8549 (N_8549,N_6969,N_7143);
xnor U8550 (N_8550,N_6548,N_6376);
or U8551 (N_8551,N_6911,N_6786);
and U8552 (N_8552,N_6606,N_6146);
nor U8553 (N_8553,N_7184,N_7136);
xor U8554 (N_8554,N_6563,N_6799);
and U8555 (N_8555,N_6425,N_7485);
and U8556 (N_8556,N_7046,N_6000);
or U8557 (N_8557,N_7060,N_6952);
nand U8558 (N_8558,N_7259,N_7339);
xnor U8559 (N_8559,N_6649,N_6495);
xnor U8560 (N_8560,N_6610,N_6705);
or U8561 (N_8561,N_6198,N_6913);
or U8562 (N_8562,N_6010,N_6882);
nand U8563 (N_8563,N_6423,N_7017);
and U8564 (N_8564,N_6059,N_7475);
or U8565 (N_8565,N_6048,N_7039);
or U8566 (N_8566,N_6517,N_6535);
nor U8567 (N_8567,N_6909,N_6839);
or U8568 (N_8568,N_7131,N_7321);
nor U8569 (N_8569,N_6987,N_6384);
xor U8570 (N_8570,N_6664,N_6292);
and U8571 (N_8571,N_6841,N_6144);
or U8572 (N_8572,N_6935,N_6432);
xnor U8573 (N_8573,N_6552,N_7408);
nor U8574 (N_8574,N_6450,N_6532);
and U8575 (N_8575,N_6222,N_7259);
nand U8576 (N_8576,N_6772,N_7420);
or U8577 (N_8577,N_6604,N_6863);
nor U8578 (N_8578,N_7056,N_7235);
and U8579 (N_8579,N_7375,N_6687);
nand U8580 (N_8580,N_6108,N_7290);
or U8581 (N_8581,N_7137,N_6382);
nor U8582 (N_8582,N_6752,N_6175);
and U8583 (N_8583,N_6780,N_6273);
and U8584 (N_8584,N_6780,N_6104);
nand U8585 (N_8585,N_6546,N_6199);
and U8586 (N_8586,N_6026,N_6943);
xor U8587 (N_8587,N_6964,N_6017);
and U8588 (N_8588,N_7460,N_6797);
and U8589 (N_8589,N_6729,N_6177);
nor U8590 (N_8590,N_7240,N_7054);
xnor U8591 (N_8591,N_6544,N_7046);
xnor U8592 (N_8592,N_6959,N_7384);
or U8593 (N_8593,N_7034,N_6416);
or U8594 (N_8594,N_6107,N_6389);
or U8595 (N_8595,N_6830,N_6494);
xnor U8596 (N_8596,N_7070,N_6215);
nor U8597 (N_8597,N_7159,N_6359);
nand U8598 (N_8598,N_7072,N_6209);
xnor U8599 (N_8599,N_6119,N_7071);
xor U8600 (N_8600,N_6533,N_7418);
and U8601 (N_8601,N_7210,N_7302);
or U8602 (N_8602,N_6054,N_6644);
nand U8603 (N_8603,N_7307,N_6353);
xor U8604 (N_8604,N_6704,N_6850);
xnor U8605 (N_8605,N_7057,N_6112);
nor U8606 (N_8606,N_7010,N_6125);
or U8607 (N_8607,N_7102,N_7078);
and U8608 (N_8608,N_6308,N_6480);
or U8609 (N_8609,N_6323,N_6811);
xnor U8610 (N_8610,N_6640,N_7003);
or U8611 (N_8611,N_6895,N_6341);
nor U8612 (N_8612,N_7325,N_6587);
or U8613 (N_8613,N_7141,N_6428);
nor U8614 (N_8614,N_6988,N_6865);
nor U8615 (N_8615,N_7137,N_7200);
or U8616 (N_8616,N_7465,N_7105);
xnor U8617 (N_8617,N_6869,N_6754);
nor U8618 (N_8618,N_7484,N_7314);
or U8619 (N_8619,N_6952,N_7463);
xor U8620 (N_8620,N_6116,N_6035);
nor U8621 (N_8621,N_6214,N_6522);
nand U8622 (N_8622,N_6381,N_7048);
xnor U8623 (N_8623,N_6717,N_7486);
nor U8624 (N_8624,N_7152,N_6433);
xnor U8625 (N_8625,N_7101,N_6496);
and U8626 (N_8626,N_6168,N_6856);
or U8627 (N_8627,N_7189,N_7437);
or U8628 (N_8628,N_6229,N_7493);
nand U8629 (N_8629,N_6582,N_6957);
nor U8630 (N_8630,N_6599,N_7306);
and U8631 (N_8631,N_7016,N_6040);
and U8632 (N_8632,N_6365,N_6120);
xnor U8633 (N_8633,N_6224,N_6241);
nor U8634 (N_8634,N_7108,N_7340);
xor U8635 (N_8635,N_6898,N_7372);
nor U8636 (N_8636,N_7365,N_6343);
or U8637 (N_8637,N_6751,N_6036);
or U8638 (N_8638,N_7018,N_7164);
nand U8639 (N_8639,N_7266,N_6702);
nor U8640 (N_8640,N_7244,N_6195);
and U8641 (N_8641,N_6514,N_6008);
or U8642 (N_8642,N_7392,N_7477);
or U8643 (N_8643,N_6799,N_7226);
nand U8644 (N_8644,N_7170,N_7077);
nand U8645 (N_8645,N_6553,N_6477);
xor U8646 (N_8646,N_6251,N_6605);
nand U8647 (N_8647,N_7142,N_6482);
xnor U8648 (N_8648,N_6625,N_7280);
and U8649 (N_8649,N_7200,N_6086);
or U8650 (N_8650,N_7379,N_7030);
nor U8651 (N_8651,N_6171,N_7114);
and U8652 (N_8652,N_7191,N_6266);
nand U8653 (N_8653,N_6755,N_6635);
xor U8654 (N_8654,N_7043,N_6783);
nor U8655 (N_8655,N_7169,N_7133);
nand U8656 (N_8656,N_7074,N_7007);
or U8657 (N_8657,N_6926,N_6847);
or U8658 (N_8658,N_6210,N_6055);
nor U8659 (N_8659,N_6079,N_7228);
or U8660 (N_8660,N_6467,N_7331);
or U8661 (N_8661,N_6738,N_7097);
nor U8662 (N_8662,N_7469,N_7383);
nand U8663 (N_8663,N_6790,N_7101);
xor U8664 (N_8664,N_7131,N_7035);
and U8665 (N_8665,N_6830,N_7098);
and U8666 (N_8666,N_7219,N_7193);
nand U8667 (N_8667,N_6741,N_6185);
nor U8668 (N_8668,N_6220,N_6571);
nor U8669 (N_8669,N_7390,N_7047);
xor U8670 (N_8670,N_7234,N_7469);
nand U8671 (N_8671,N_6145,N_6802);
nand U8672 (N_8672,N_6902,N_7422);
nor U8673 (N_8673,N_6575,N_6383);
nor U8674 (N_8674,N_7130,N_7440);
nor U8675 (N_8675,N_6579,N_7344);
nor U8676 (N_8676,N_7280,N_6931);
nor U8677 (N_8677,N_6804,N_6271);
or U8678 (N_8678,N_7287,N_6749);
and U8679 (N_8679,N_7294,N_7003);
or U8680 (N_8680,N_6361,N_6201);
nor U8681 (N_8681,N_7212,N_6746);
nor U8682 (N_8682,N_6368,N_6568);
nor U8683 (N_8683,N_6680,N_6507);
and U8684 (N_8684,N_6645,N_6079);
and U8685 (N_8685,N_6266,N_6452);
nor U8686 (N_8686,N_7479,N_6163);
and U8687 (N_8687,N_6853,N_7254);
or U8688 (N_8688,N_6401,N_6665);
and U8689 (N_8689,N_6936,N_6818);
nand U8690 (N_8690,N_7458,N_6285);
nand U8691 (N_8691,N_6450,N_6920);
nand U8692 (N_8692,N_6438,N_7377);
and U8693 (N_8693,N_6160,N_6418);
nor U8694 (N_8694,N_7459,N_7109);
nand U8695 (N_8695,N_7482,N_6481);
nand U8696 (N_8696,N_7334,N_6612);
xnor U8697 (N_8697,N_7091,N_6321);
and U8698 (N_8698,N_7075,N_6394);
nand U8699 (N_8699,N_7412,N_7018);
xnor U8700 (N_8700,N_6576,N_6339);
and U8701 (N_8701,N_6776,N_6880);
nor U8702 (N_8702,N_6513,N_6048);
xor U8703 (N_8703,N_6289,N_6485);
xor U8704 (N_8704,N_7229,N_7210);
xor U8705 (N_8705,N_7194,N_6885);
or U8706 (N_8706,N_7245,N_7030);
nor U8707 (N_8707,N_6002,N_6623);
or U8708 (N_8708,N_6009,N_7391);
xnor U8709 (N_8709,N_7397,N_7369);
or U8710 (N_8710,N_6247,N_6516);
or U8711 (N_8711,N_6853,N_6081);
nand U8712 (N_8712,N_6287,N_6468);
and U8713 (N_8713,N_6646,N_6017);
and U8714 (N_8714,N_6912,N_7163);
and U8715 (N_8715,N_6933,N_7250);
and U8716 (N_8716,N_7314,N_6055);
nor U8717 (N_8717,N_6513,N_6390);
xnor U8718 (N_8718,N_6705,N_6981);
xor U8719 (N_8719,N_6682,N_6494);
nor U8720 (N_8720,N_6161,N_7108);
xor U8721 (N_8721,N_7399,N_6498);
nor U8722 (N_8722,N_7214,N_6918);
nor U8723 (N_8723,N_6123,N_6771);
xor U8724 (N_8724,N_6317,N_6286);
nand U8725 (N_8725,N_6607,N_6362);
nand U8726 (N_8726,N_6213,N_7349);
xor U8727 (N_8727,N_6326,N_6552);
nor U8728 (N_8728,N_7448,N_6963);
or U8729 (N_8729,N_6503,N_6128);
and U8730 (N_8730,N_6574,N_6656);
nor U8731 (N_8731,N_6179,N_7173);
nand U8732 (N_8732,N_7015,N_6561);
or U8733 (N_8733,N_6714,N_6009);
nor U8734 (N_8734,N_7338,N_6907);
or U8735 (N_8735,N_6337,N_7267);
or U8736 (N_8736,N_7261,N_6836);
nor U8737 (N_8737,N_7298,N_6317);
nand U8738 (N_8738,N_7182,N_6058);
and U8739 (N_8739,N_7108,N_6291);
and U8740 (N_8740,N_6190,N_6531);
and U8741 (N_8741,N_6339,N_7204);
or U8742 (N_8742,N_6933,N_6865);
or U8743 (N_8743,N_6072,N_6248);
or U8744 (N_8744,N_7444,N_6114);
nand U8745 (N_8745,N_7322,N_6378);
nor U8746 (N_8746,N_6228,N_6915);
or U8747 (N_8747,N_6121,N_6853);
or U8748 (N_8748,N_7460,N_6073);
and U8749 (N_8749,N_6080,N_6655);
xor U8750 (N_8750,N_6825,N_6568);
or U8751 (N_8751,N_7400,N_6856);
or U8752 (N_8752,N_6102,N_7105);
and U8753 (N_8753,N_6061,N_6130);
nand U8754 (N_8754,N_6662,N_7082);
xor U8755 (N_8755,N_6148,N_7431);
nand U8756 (N_8756,N_6464,N_6749);
nor U8757 (N_8757,N_6137,N_6747);
and U8758 (N_8758,N_6469,N_6267);
or U8759 (N_8759,N_6509,N_6249);
nor U8760 (N_8760,N_6313,N_6838);
xor U8761 (N_8761,N_6470,N_6489);
and U8762 (N_8762,N_6376,N_7352);
nand U8763 (N_8763,N_7149,N_6488);
and U8764 (N_8764,N_6384,N_7125);
xnor U8765 (N_8765,N_6820,N_7097);
nor U8766 (N_8766,N_6016,N_6238);
and U8767 (N_8767,N_6542,N_6739);
nor U8768 (N_8768,N_7288,N_7256);
xnor U8769 (N_8769,N_7297,N_6092);
nand U8770 (N_8770,N_7028,N_7014);
or U8771 (N_8771,N_6233,N_6530);
and U8772 (N_8772,N_7263,N_6417);
nand U8773 (N_8773,N_7140,N_7106);
nand U8774 (N_8774,N_7464,N_7174);
or U8775 (N_8775,N_7448,N_6130);
xor U8776 (N_8776,N_6380,N_6484);
xor U8777 (N_8777,N_6014,N_7202);
or U8778 (N_8778,N_6329,N_6311);
xor U8779 (N_8779,N_7122,N_6393);
nand U8780 (N_8780,N_7286,N_6887);
and U8781 (N_8781,N_6335,N_6405);
nand U8782 (N_8782,N_7371,N_6782);
xor U8783 (N_8783,N_6177,N_7142);
nand U8784 (N_8784,N_7062,N_6817);
and U8785 (N_8785,N_6189,N_6790);
nor U8786 (N_8786,N_6166,N_7428);
nand U8787 (N_8787,N_6078,N_6818);
xnor U8788 (N_8788,N_7440,N_6171);
or U8789 (N_8789,N_6644,N_6434);
nor U8790 (N_8790,N_6313,N_7210);
and U8791 (N_8791,N_6419,N_6438);
and U8792 (N_8792,N_6363,N_6851);
or U8793 (N_8793,N_7369,N_6505);
or U8794 (N_8794,N_6876,N_6784);
nand U8795 (N_8795,N_6814,N_6967);
and U8796 (N_8796,N_6893,N_6608);
or U8797 (N_8797,N_6886,N_6904);
nand U8798 (N_8798,N_6600,N_6176);
nand U8799 (N_8799,N_7478,N_7289);
or U8800 (N_8800,N_6633,N_6219);
or U8801 (N_8801,N_7246,N_6926);
nand U8802 (N_8802,N_6518,N_7299);
or U8803 (N_8803,N_6182,N_6343);
xor U8804 (N_8804,N_6101,N_6780);
and U8805 (N_8805,N_7378,N_6143);
nor U8806 (N_8806,N_6175,N_6680);
or U8807 (N_8807,N_6675,N_6850);
nand U8808 (N_8808,N_6211,N_6210);
nor U8809 (N_8809,N_7330,N_6760);
nand U8810 (N_8810,N_7322,N_7203);
nand U8811 (N_8811,N_6053,N_6740);
nor U8812 (N_8812,N_6880,N_6947);
nor U8813 (N_8813,N_7393,N_7135);
nand U8814 (N_8814,N_6505,N_6495);
and U8815 (N_8815,N_7266,N_6881);
and U8816 (N_8816,N_6671,N_6882);
or U8817 (N_8817,N_6170,N_6952);
or U8818 (N_8818,N_6022,N_6144);
nand U8819 (N_8819,N_7465,N_6153);
nand U8820 (N_8820,N_7152,N_7140);
nor U8821 (N_8821,N_6745,N_6990);
nor U8822 (N_8822,N_7015,N_6139);
nor U8823 (N_8823,N_7311,N_7106);
or U8824 (N_8824,N_6748,N_7425);
nor U8825 (N_8825,N_6637,N_7257);
nand U8826 (N_8826,N_7174,N_6427);
nor U8827 (N_8827,N_6952,N_6969);
and U8828 (N_8828,N_6255,N_6450);
and U8829 (N_8829,N_6697,N_6462);
and U8830 (N_8830,N_6900,N_7348);
nor U8831 (N_8831,N_6633,N_7483);
xor U8832 (N_8832,N_6338,N_7205);
and U8833 (N_8833,N_6336,N_6351);
nand U8834 (N_8834,N_6495,N_6257);
nor U8835 (N_8835,N_6903,N_6799);
nand U8836 (N_8836,N_6233,N_6183);
xnor U8837 (N_8837,N_6828,N_6730);
and U8838 (N_8838,N_7479,N_6042);
and U8839 (N_8839,N_7042,N_7268);
nand U8840 (N_8840,N_6267,N_6802);
nand U8841 (N_8841,N_7448,N_7018);
nand U8842 (N_8842,N_6773,N_6713);
or U8843 (N_8843,N_6604,N_6575);
and U8844 (N_8844,N_6086,N_7397);
nand U8845 (N_8845,N_6375,N_7425);
or U8846 (N_8846,N_7068,N_6567);
and U8847 (N_8847,N_6048,N_6591);
or U8848 (N_8848,N_6678,N_7292);
and U8849 (N_8849,N_6144,N_6531);
nor U8850 (N_8850,N_6018,N_6327);
or U8851 (N_8851,N_6337,N_6708);
and U8852 (N_8852,N_6935,N_6686);
nand U8853 (N_8853,N_7177,N_7117);
or U8854 (N_8854,N_7474,N_7259);
nand U8855 (N_8855,N_7428,N_7213);
or U8856 (N_8856,N_7424,N_6542);
or U8857 (N_8857,N_6399,N_6895);
xor U8858 (N_8858,N_7305,N_6017);
nand U8859 (N_8859,N_6579,N_6233);
nor U8860 (N_8860,N_6422,N_6006);
nand U8861 (N_8861,N_7257,N_6856);
xor U8862 (N_8862,N_7353,N_6385);
nand U8863 (N_8863,N_6966,N_6364);
xor U8864 (N_8864,N_6673,N_6860);
nand U8865 (N_8865,N_7440,N_7370);
or U8866 (N_8866,N_7168,N_7328);
and U8867 (N_8867,N_6715,N_6287);
and U8868 (N_8868,N_6509,N_6657);
nand U8869 (N_8869,N_7018,N_6110);
nand U8870 (N_8870,N_7363,N_7069);
and U8871 (N_8871,N_6404,N_6625);
or U8872 (N_8872,N_7160,N_7197);
nor U8873 (N_8873,N_6009,N_6732);
nand U8874 (N_8874,N_6745,N_6607);
or U8875 (N_8875,N_7189,N_6492);
nand U8876 (N_8876,N_6835,N_7202);
nor U8877 (N_8877,N_6098,N_7091);
xor U8878 (N_8878,N_6294,N_7376);
and U8879 (N_8879,N_6446,N_7353);
and U8880 (N_8880,N_7213,N_7356);
nand U8881 (N_8881,N_7387,N_7323);
xor U8882 (N_8882,N_6734,N_6820);
and U8883 (N_8883,N_6081,N_6637);
nand U8884 (N_8884,N_6363,N_6779);
or U8885 (N_8885,N_7452,N_7182);
and U8886 (N_8886,N_7255,N_6422);
nor U8887 (N_8887,N_6257,N_7016);
nand U8888 (N_8888,N_6518,N_6195);
xor U8889 (N_8889,N_6876,N_6924);
nand U8890 (N_8890,N_7408,N_6145);
nor U8891 (N_8891,N_7197,N_6030);
and U8892 (N_8892,N_6498,N_6597);
or U8893 (N_8893,N_7318,N_6245);
nand U8894 (N_8894,N_6201,N_6989);
xnor U8895 (N_8895,N_6602,N_6408);
nand U8896 (N_8896,N_7347,N_7018);
or U8897 (N_8897,N_6962,N_7233);
or U8898 (N_8898,N_6942,N_7039);
nand U8899 (N_8899,N_6765,N_6278);
or U8900 (N_8900,N_6004,N_6190);
nand U8901 (N_8901,N_6460,N_6755);
nor U8902 (N_8902,N_6573,N_6198);
nor U8903 (N_8903,N_7353,N_6233);
and U8904 (N_8904,N_6775,N_6631);
nand U8905 (N_8905,N_7456,N_6221);
or U8906 (N_8906,N_7131,N_6957);
and U8907 (N_8907,N_7307,N_6808);
and U8908 (N_8908,N_7469,N_7392);
and U8909 (N_8909,N_6130,N_6089);
nand U8910 (N_8910,N_7346,N_6825);
xor U8911 (N_8911,N_6598,N_7411);
nand U8912 (N_8912,N_7388,N_6811);
and U8913 (N_8913,N_7371,N_6850);
xor U8914 (N_8914,N_7243,N_7239);
or U8915 (N_8915,N_7292,N_7062);
nand U8916 (N_8916,N_7014,N_6576);
or U8917 (N_8917,N_6127,N_6019);
nand U8918 (N_8918,N_6022,N_7087);
or U8919 (N_8919,N_6344,N_7130);
and U8920 (N_8920,N_6257,N_6656);
and U8921 (N_8921,N_6094,N_6950);
nand U8922 (N_8922,N_6772,N_6337);
nor U8923 (N_8923,N_6178,N_6187);
nand U8924 (N_8924,N_7291,N_7121);
nor U8925 (N_8925,N_6964,N_6747);
nor U8926 (N_8926,N_6088,N_7486);
nand U8927 (N_8927,N_6938,N_7083);
xnor U8928 (N_8928,N_7354,N_7234);
xor U8929 (N_8929,N_6684,N_6028);
nand U8930 (N_8930,N_6843,N_6779);
or U8931 (N_8931,N_6460,N_6485);
and U8932 (N_8932,N_6071,N_7196);
nor U8933 (N_8933,N_7255,N_6742);
xnor U8934 (N_8934,N_7489,N_7447);
or U8935 (N_8935,N_6771,N_6818);
nand U8936 (N_8936,N_6857,N_6051);
nand U8937 (N_8937,N_7055,N_6080);
and U8938 (N_8938,N_6418,N_7371);
or U8939 (N_8939,N_6123,N_6227);
xor U8940 (N_8940,N_6241,N_7272);
xor U8941 (N_8941,N_6508,N_6927);
and U8942 (N_8942,N_6752,N_7127);
nor U8943 (N_8943,N_7219,N_6823);
and U8944 (N_8944,N_7111,N_6828);
and U8945 (N_8945,N_6377,N_6896);
nand U8946 (N_8946,N_6395,N_6499);
and U8947 (N_8947,N_6237,N_6603);
and U8948 (N_8948,N_7406,N_7315);
xnor U8949 (N_8949,N_7031,N_6734);
and U8950 (N_8950,N_7338,N_6353);
nor U8951 (N_8951,N_7189,N_6819);
nand U8952 (N_8952,N_6776,N_6186);
nand U8953 (N_8953,N_6912,N_7417);
xnor U8954 (N_8954,N_6191,N_6206);
nand U8955 (N_8955,N_6727,N_7431);
nor U8956 (N_8956,N_6595,N_7293);
nand U8957 (N_8957,N_7256,N_6164);
and U8958 (N_8958,N_7017,N_7415);
xnor U8959 (N_8959,N_6277,N_6891);
and U8960 (N_8960,N_6557,N_6050);
nor U8961 (N_8961,N_6645,N_6021);
nand U8962 (N_8962,N_7497,N_6099);
or U8963 (N_8963,N_6699,N_7188);
nor U8964 (N_8964,N_7157,N_7031);
or U8965 (N_8965,N_6667,N_6159);
or U8966 (N_8966,N_6081,N_6782);
xnor U8967 (N_8967,N_6180,N_6667);
nand U8968 (N_8968,N_6855,N_6808);
nand U8969 (N_8969,N_6485,N_7450);
nand U8970 (N_8970,N_6051,N_6359);
xnor U8971 (N_8971,N_7334,N_7287);
nor U8972 (N_8972,N_6399,N_6485);
nand U8973 (N_8973,N_6560,N_6168);
xnor U8974 (N_8974,N_6529,N_6321);
nand U8975 (N_8975,N_7269,N_6854);
or U8976 (N_8976,N_7386,N_6770);
or U8977 (N_8977,N_6492,N_6448);
and U8978 (N_8978,N_6249,N_7329);
nand U8979 (N_8979,N_6167,N_7132);
xor U8980 (N_8980,N_6053,N_6439);
xor U8981 (N_8981,N_6717,N_6999);
nor U8982 (N_8982,N_7341,N_6408);
xnor U8983 (N_8983,N_6169,N_7462);
xnor U8984 (N_8984,N_6257,N_6777);
and U8985 (N_8985,N_7379,N_6211);
or U8986 (N_8986,N_6355,N_6289);
xnor U8987 (N_8987,N_6508,N_7491);
and U8988 (N_8988,N_6276,N_6317);
nor U8989 (N_8989,N_7475,N_6366);
nand U8990 (N_8990,N_6074,N_7427);
nor U8991 (N_8991,N_6859,N_7041);
or U8992 (N_8992,N_6504,N_6280);
xor U8993 (N_8993,N_7399,N_6154);
nor U8994 (N_8994,N_7448,N_6559);
and U8995 (N_8995,N_6580,N_6085);
nand U8996 (N_8996,N_6608,N_6680);
and U8997 (N_8997,N_7412,N_7212);
and U8998 (N_8998,N_7035,N_6588);
or U8999 (N_8999,N_7024,N_6816);
nand U9000 (N_9000,N_7666,N_8626);
xnor U9001 (N_9001,N_8182,N_8557);
or U9002 (N_9002,N_7534,N_8648);
xnor U9003 (N_9003,N_8365,N_8984);
or U9004 (N_9004,N_8128,N_7912);
nand U9005 (N_9005,N_8653,N_8979);
nor U9006 (N_9006,N_8733,N_8873);
or U9007 (N_9007,N_8125,N_8506);
nor U9008 (N_9008,N_8574,N_7807);
nor U9009 (N_9009,N_8722,N_7724);
or U9010 (N_9010,N_8679,N_8613);
or U9011 (N_9011,N_8573,N_7767);
xor U9012 (N_9012,N_8167,N_8638);
nor U9013 (N_9013,N_8185,N_8316);
nand U9014 (N_9014,N_8717,N_8224);
and U9015 (N_9015,N_8403,N_8452);
nand U9016 (N_9016,N_7952,N_7799);
or U9017 (N_9017,N_8639,N_8404);
xnor U9018 (N_9018,N_8269,N_8333);
nand U9019 (N_9019,N_8256,N_8086);
nor U9020 (N_9020,N_7926,N_8650);
and U9021 (N_9021,N_8659,N_8533);
nand U9022 (N_9022,N_7521,N_8723);
xor U9023 (N_9023,N_8521,N_8575);
or U9024 (N_9024,N_8137,N_8629);
nand U9025 (N_9025,N_7833,N_8692);
xor U9026 (N_9026,N_8524,N_8024);
nand U9027 (N_9027,N_8395,N_7838);
and U9028 (N_9028,N_7786,N_7658);
and U9029 (N_9029,N_7585,N_7847);
or U9030 (N_9030,N_7955,N_7975);
nand U9031 (N_9031,N_8095,N_8487);
xnor U9032 (N_9032,N_8989,N_8541);
nand U9033 (N_9033,N_8078,N_7871);
or U9034 (N_9034,N_7698,N_8826);
and U9035 (N_9035,N_8448,N_7587);
or U9036 (N_9036,N_8587,N_7715);
and U9037 (N_9037,N_7738,N_8177);
xor U9038 (N_9038,N_7832,N_8703);
or U9039 (N_9039,N_8774,N_8340);
nor U9040 (N_9040,N_8975,N_7553);
nand U9041 (N_9041,N_8896,N_8415);
nor U9042 (N_9042,N_8329,N_8569);
xor U9043 (N_9043,N_8258,N_7879);
xnor U9044 (N_9044,N_8772,N_8549);
nor U9045 (N_9045,N_7999,N_7728);
nand U9046 (N_9046,N_8065,N_8740);
and U9047 (N_9047,N_8370,N_8903);
and U9048 (N_9048,N_7776,N_7577);
nand U9049 (N_9049,N_8938,N_7506);
nor U9050 (N_9050,N_8165,N_8335);
nand U9051 (N_9051,N_7761,N_8787);
or U9052 (N_9052,N_7522,N_8062);
and U9053 (N_9053,N_8363,N_7866);
nor U9054 (N_9054,N_7524,N_8806);
and U9055 (N_9055,N_8630,N_8614);
nor U9056 (N_9056,N_7629,N_8360);
nand U9057 (N_9057,N_7665,N_8241);
nor U9058 (N_9058,N_8059,N_7951);
nor U9059 (N_9059,N_7798,N_8757);
or U9060 (N_9060,N_8930,N_8718);
nand U9061 (N_9061,N_8645,N_8243);
and U9062 (N_9062,N_8282,N_7993);
xor U9063 (N_9063,N_8788,N_7523);
xor U9064 (N_9064,N_8479,N_8127);
and U9065 (N_9065,N_7809,N_8738);
nor U9066 (N_9066,N_8496,N_7802);
and U9067 (N_9067,N_8001,N_8838);
nand U9068 (N_9068,N_7875,N_8463);
nor U9069 (N_9069,N_8298,N_8249);
xnor U9070 (N_9070,N_8158,N_7707);
nand U9071 (N_9071,N_7920,N_7624);
and U9072 (N_9072,N_7970,N_8015);
xor U9073 (N_9073,N_7749,N_8414);
nor U9074 (N_9074,N_8144,N_7998);
or U9075 (N_9075,N_7708,N_8622);
nand U9076 (N_9076,N_8719,N_8002);
xnor U9077 (N_9077,N_7566,N_8747);
nand U9078 (N_9078,N_8545,N_7742);
nand U9079 (N_9079,N_8210,N_8766);
nor U9080 (N_9080,N_8320,N_8209);
and U9081 (N_9081,N_8584,N_8368);
nor U9082 (N_9082,N_8123,N_8477);
nand U9083 (N_9083,N_8773,N_7796);
nor U9084 (N_9084,N_8832,N_8369);
or U9085 (N_9085,N_7601,N_7922);
nor U9086 (N_9086,N_7830,N_7514);
nor U9087 (N_9087,N_7891,N_8051);
or U9088 (N_9088,N_7722,N_8789);
xnor U9089 (N_9089,N_8735,N_8874);
and U9090 (N_9090,N_7909,N_8279);
nand U9091 (N_9091,N_8830,N_8852);
and U9092 (N_9092,N_7840,N_8563);
nand U9093 (N_9093,N_8118,N_8461);
nor U9094 (N_9094,N_7633,N_8802);
and U9095 (N_9095,N_8032,N_7932);
nor U9096 (N_9096,N_8712,N_8381);
xnor U9097 (N_9097,N_8000,N_7701);
and U9098 (N_9098,N_8306,N_7801);
or U9099 (N_9099,N_7588,N_7874);
or U9100 (N_9100,N_8536,N_8726);
nand U9101 (N_9101,N_7509,N_8163);
and U9102 (N_9102,N_7712,N_8605);
or U9103 (N_9103,N_7500,N_7923);
nor U9104 (N_9104,N_8300,N_7659);
and U9105 (N_9105,N_7681,N_8528);
nand U9106 (N_9106,N_7815,N_8084);
nor U9107 (N_9107,N_8834,N_8516);
or U9108 (N_9108,N_8089,N_7649);
nand U9109 (N_9109,N_7925,N_8121);
nand U9110 (N_9110,N_8221,N_8152);
nand U9111 (N_9111,N_8073,N_8105);
nor U9112 (N_9112,N_8963,N_8715);
xnor U9113 (N_9113,N_7619,N_7638);
or U9114 (N_9114,N_8977,N_7532);
xor U9115 (N_9115,N_7605,N_8254);
nor U9116 (N_9116,N_7579,N_7705);
or U9117 (N_9117,N_8186,N_8696);
or U9118 (N_9118,N_8429,N_8753);
or U9119 (N_9119,N_7949,N_8571);
nor U9120 (N_9120,N_7667,N_8960);
or U9121 (N_9121,N_8503,N_8055);
or U9122 (N_9122,N_8804,N_8421);
nor U9123 (N_9123,N_8619,N_8231);
or U9124 (N_9124,N_8682,N_7824);
nand U9125 (N_9125,N_8156,N_7727);
and U9126 (N_9126,N_8449,N_7508);
nor U9127 (N_9127,N_8771,N_8262);
nand U9128 (N_9128,N_7657,N_8932);
nand U9129 (N_9129,N_8920,N_8029);
nor U9130 (N_9130,N_8546,N_8512);
nand U9131 (N_9131,N_8099,N_7897);
xnor U9132 (N_9132,N_7716,N_8887);
and U9133 (N_9133,N_8017,N_8828);
and U9134 (N_9134,N_8367,N_8651);
or U9135 (N_9135,N_7812,N_8204);
and U9136 (N_9136,N_7687,N_8390);
nor U9137 (N_9137,N_7621,N_8762);
nor U9138 (N_9138,N_7614,N_7718);
and U9139 (N_9139,N_7511,N_8981);
and U9140 (N_9140,N_8969,N_8933);
and U9141 (N_9141,N_7694,N_8854);
or U9142 (N_9142,N_8219,N_8862);
nand U9143 (N_9143,N_7976,N_7714);
xor U9144 (N_9144,N_8202,N_7792);
nand U9145 (N_9145,N_7977,N_8674);
or U9146 (N_9146,N_8867,N_8866);
and U9147 (N_9147,N_7930,N_8748);
nor U9148 (N_9148,N_8225,N_8223);
nor U9149 (N_9149,N_8926,N_8778);
xor U9150 (N_9150,N_8423,N_8750);
xor U9151 (N_9151,N_8120,N_8011);
nor U9152 (N_9152,N_7573,N_7651);
nor U9153 (N_9153,N_8042,N_8678);
and U9154 (N_9154,N_7725,N_7545);
or U9155 (N_9155,N_8013,N_8267);
and U9156 (N_9156,N_7870,N_8326);
nand U9157 (N_9157,N_8285,N_7544);
nor U9158 (N_9158,N_7820,N_7917);
nand U9159 (N_9159,N_7984,N_8473);
or U9160 (N_9160,N_8428,N_8990);
nand U9161 (N_9161,N_7726,N_8208);
and U9162 (N_9162,N_8673,N_8978);
nand U9163 (N_9163,N_8490,N_8507);
xnor U9164 (N_9164,N_8129,N_8610);
or U9165 (N_9165,N_8686,N_8486);
xnor U9166 (N_9166,N_8627,N_7885);
and U9167 (N_9167,N_7757,N_8705);
nand U9168 (N_9168,N_7965,N_7916);
xor U9169 (N_9169,N_8378,N_8822);
xor U9170 (N_9170,N_8841,N_8080);
and U9171 (N_9171,N_8038,N_8550);
or U9172 (N_9172,N_8230,N_7581);
and U9173 (N_9173,N_8965,N_8359);
nor U9174 (N_9174,N_7873,N_8636);
or U9175 (N_9175,N_8211,N_8139);
nor U9176 (N_9176,N_8661,N_8079);
nor U9177 (N_9177,N_7555,N_7668);
nor U9178 (N_9178,N_8149,N_8576);
nand U9179 (N_9179,N_8777,N_8554);
xnor U9180 (N_9180,N_8034,N_7859);
nor U9181 (N_9181,N_8025,N_8336);
nor U9182 (N_9182,N_8364,N_8294);
nor U9183 (N_9183,N_7700,N_8160);
xor U9184 (N_9184,N_8611,N_7857);
and U9185 (N_9185,N_8019,N_7630);
xnor U9186 (N_9186,N_8312,N_8842);
nor U9187 (N_9187,N_7967,N_8976);
nor U9188 (N_9188,N_7743,N_8052);
or U9189 (N_9189,N_8594,N_7759);
nor U9190 (N_9190,N_8330,N_7887);
xor U9191 (N_9191,N_7686,N_8270);
and U9192 (N_9192,N_8746,N_8586);
and U9193 (N_9193,N_7836,N_7663);
nor U9194 (N_9194,N_8143,N_8472);
nor U9195 (N_9195,N_8592,N_8839);
nor U9196 (N_9196,N_8244,N_8328);
nor U9197 (N_9197,N_8663,N_7852);
nand U9198 (N_9198,N_7939,N_7986);
and U9199 (N_9199,N_8341,N_7919);
nand U9200 (N_9200,N_8606,N_8483);
and U9201 (N_9201,N_8642,N_8155);
nand U9202 (N_9202,N_8094,N_8140);
xor U9203 (N_9203,N_8603,N_8445);
and U9204 (N_9204,N_8814,N_8407);
nor U9205 (N_9205,N_7782,N_8810);
xor U9206 (N_9206,N_7530,N_7888);
or U9207 (N_9207,N_8667,N_7893);
or U9208 (N_9208,N_8646,N_7773);
xnor U9209 (N_9209,N_8173,N_8767);
or U9210 (N_9210,N_8598,N_8222);
nor U9211 (N_9211,N_7631,N_7613);
and U9212 (N_9212,N_8096,N_8676);
or U9213 (N_9213,N_8565,N_8302);
or U9214 (N_9214,N_8184,N_8878);
xnor U9215 (N_9215,N_8540,N_8985);
nand U9216 (N_9216,N_8464,N_8572);
nor U9217 (N_9217,N_8205,N_7642);
nand U9218 (N_9218,N_7981,N_8044);
and U9219 (N_9219,N_8396,N_8092);
xor U9220 (N_9220,N_7770,N_8652);
nor U9221 (N_9221,N_7565,N_8426);
xor U9222 (N_9222,N_8315,N_8836);
and U9223 (N_9223,N_7823,N_8314);
nand U9224 (N_9224,N_8162,N_8088);
xor U9225 (N_9225,N_8510,N_8945);
nand U9226 (N_9226,N_7685,N_7933);
and U9227 (N_9227,N_8688,N_8580);
xnor U9228 (N_9228,N_8453,N_7813);
or U9229 (N_9229,N_8045,N_7793);
xnor U9230 (N_9230,N_7961,N_7768);
nand U9231 (N_9231,N_8220,N_8730);
nand U9232 (N_9232,N_8954,N_7515);
nor U9233 (N_9233,N_7853,N_8462);
xnor U9234 (N_9234,N_8431,N_7869);
or U9235 (N_9235,N_7570,N_7695);
or U9236 (N_9236,N_8133,N_8508);
nor U9237 (N_9237,N_7906,N_8885);
xnor U9238 (N_9238,N_8548,N_8928);
nand U9239 (N_9239,N_7914,N_8194);
nand U9240 (N_9240,N_8801,N_8523);
nand U9241 (N_9241,N_8958,N_7626);
nand U9242 (N_9242,N_8552,N_8704);
and U9243 (N_9243,N_7697,N_7525);
or U9244 (N_9244,N_7542,N_8699);
xnor U9245 (N_9245,N_8591,N_7778);
or U9246 (N_9246,N_8175,N_8391);
nand U9247 (N_9247,N_8456,N_8710);
xor U9248 (N_9248,N_8869,N_8897);
and U9249 (N_9249,N_8737,N_8408);
nor U9250 (N_9250,N_8698,N_8103);
or U9251 (N_9251,N_7635,N_8317);
nor U9252 (N_9252,N_8337,N_7600);
nand U9253 (N_9253,N_8147,N_7683);
nor U9254 (N_9254,N_8641,N_7568);
and U9255 (N_9255,N_7872,N_8784);
xnor U9256 (N_9256,N_7602,N_8207);
nand U9257 (N_9257,N_8402,N_8539);
or U9258 (N_9258,N_7516,N_8693);
nor U9259 (N_9259,N_7856,N_8036);
xnor U9260 (N_9260,N_7652,N_8366);
xor U9261 (N_9261,N_8690,N_8716);
and U9262 (N_9262,N_8906,N_7719);
or U9263 (N_9263,N_7901,N_8634);
xor U9264 (N_9264,N_8427,N_8388);
nand U9265 (N_9265,N_8988,N_8919);
nor U9266 (N_9266,N_8325,N_8174);
or U9267 (N_9267,N_8235,N_7898);
and U9268 (N_9268,N_7609,N_8176);
and U9269 (N_9269,N_7862,N_8198);
xnor U9270 (N_9270,N_8560,N_8239);
nor U9271 (N_9271,N_7746,N_7550);
and U9272 (N_9272,N_8022,N_8600);
nor U9273 (N_9273,N_7662,N_8820);
and U9274 (N_9274,N_7945,N_8907);
xnor U9275 (N_9275,N_7504,N_7547);
xnor U9276 (N_9276,N_7858,N_8082);
nor U9277 (N_9277,N_7561,N_7758);
and U9278 (N_9278,N_7953,N_7501);
nor U9279 (N_9279,N_8203,N_8070);
and U9280 (N_9280,N_8765,N_8392);
nand U9281 (N_9281,N_8706,N_8769);
or U9282 (N_9282,N_7894,N_7639);
nor U9283 (N_9283,N_7988,N_8941);
or U9284 (N_9284,N_8432,N_7689);
nand U9285 (N_9285,N_8009,N_8383);
xnor U9286 (N_9286,N_8293,N_8434);
xnor U9287 (N_9287,N_8498,N_8242);
and U9288 (N_9288,N_7591,N_8962);
nand U9289 (N_9289,N_8201,N_8405);
nand U9290 (N_9290,N_7507,N_8470);
and U9291 (N_9291,N_7985,N_8342);
and U9292 (N_9292,N_8216,N_8899);
and U9293 (N_9293,N_8680,N_8687);
xor U9294 (N_9294,N_8343,N_8786);
xor U9295 (N_9295,N_7983,N_8491);
nor U9296 (N_9296,N_7829,N_7740);
nor U9297 (N_9297,N_7541,N_8465);
and U9298 (N_9298,N_8732,N_7637);
nor U9299 (N_9299,N_8284,N_7822);
nor U9300 (N_9300,N_7854,N_8884);
and U9301 (N_9301,N_8280,N_8997);
nand U9302 (N_9302,N_7526,N_7849);
or U9303 (N_9303,N_8106,N_8247);
nand U9304 (N_9304,N_8871,N_7603);
and U9305 (N_9305,N_8311,N_8063);
or U9306 (N_9306,N_8373,N_7878);
and U9307 (N_9307,N_8555,N_7850);
and U9308 (N_9308,N_8098,N_8334);
xor U9309 (N_9309,N_7938,N_8588);
or U9310 (N_9310,N_8911,N_8713);
or U9311 (N_9311,N_8640,N_7537);
and U9312 (N_9312,N_8910,N_7966);
and U9313 (N_9313,N_7911,N_7596);
and U9314 (N_9314,N_7992,N_7831);
and U9315 (N_9315,N_7628,N_7785);
or U9316 (N_9316,N_8877,N_8662);
xor U9317 (N_9317,N_8664,N_8188);
nand U9318 (N_9318,N_8595,N_8308);
or U9319 (N_9319,N_8898,N_8803);
xnor U9320 (N_9320,N_8108,N_7580);
xnor U9321 (N_9321,N_8081,N_7764);
nor U9322 (N_9322,N_7676,N_7554);
and U9323 (N_9323,N_8991,N_7623);
and U9324 (N_9324,N_7861,N_7944);
xor U9325 (N_9325,N_7680,N_8087);
nor U9326 (N_9326,N_8245,N_7702);
xnor U9327 (N_9327,N_8425,N_8271);
nand U9328 (N_9328,N_7766,N_8827);
or U9329 (N_9329,N_8050,N_7641);
nor U9330 (N_9330,N_7502,N_8913);
xor U9331 (N_9331,N_8649,N_8831);
or U9332 (N_9332,N_7654,N_8957);
nor U9333 (N_9333,N_8509,N_8179);
nand U9334 (N_9334,N_8353,N_7814);
or U9335 (N_9335,N_7670,N_8891);
nand U9336 (N_9336,N_7994,N_8457);
nand U9337 (N_9337,N_7540,N_7943);
xor U9338 (N_9338,N_8362,N_8657);
xnor U9339 (N_9339,N_8272,N_7996);
nand U9340 (N_9340,N_8049,N_7611);
and U9341 (N_9341,N_8537,N_8864);
or U9342 (N_9342,N_8754,N_7784);
nand U9343 (N_9343,N_8593,N_8134);
and U9344 (N_9344,N_8357,N_7851);
xor U9345 (N_9345,N_7599,N_7972);
xor U9346 (N_9346,N_8348,N_8468);
or U9347 (N_9347,N_8808,N_8596);
or U9348 (N_9348,N_7929,N_8450);
nand U9349 (N_9349,N_8812,N_8518);
or U9350 (N_9350,N_8665,N_8422);
nand U9351 (N_9351,N_8499,N_8060);
and U9352 (N_9352,N_8263,N_8601);
nand U9353 (N_9353,N_7675,N_8455);
xnor U9354 (N_9354,N_8475,N_7989);
and U9355 (N_9355,N_7699,N_8039);
xnor U9356 (N_9356,N_8781,N_8237);
and U9357 (N_9357,N_8529,N_8908);
or U9358 (N_9358,N_7868,N_8743);
or U9359 (N_9359,N_8206,N_8790);
nand U9360 (N_9360,N_7720,N_7552);
nand U9361 (N_9361,N_8213,N_7618);
xnor U9362 (N_9362,N_8807,N_7634);
nand U9363 (N_9363,N_7513,N_7771);
nand U9364 (N_9364,N_8775,N_8872);
nand U9365 (N_9365,N_8138,N_7648);
and U9366 (N_9366,N_7732,N_8685);
xor U9367 (N_9367,N_7877,N_7558);
nand U9368 (N_9368,N_8809,N_7997);
xnor U9369 (N_9369,N_7576,N_7549);
or U9370 (N_9370,N_7598,N_8145);
and U9371 (N_9371,N_8351,N_8542);
xor U9372 (N_9372,N_7733,N_7647);
nand U9373 (N_9373,N_7512,N_7693);
and U9374 (N_9374,N_8354,N_7661);
and U9375 (N_9375,N_8522,N_7803);
nand U9376 (N_9376,N_7797,N_8924);
nand U9377 (N_9377,N_7848,N_8292);
or U9378 (N_9378,N_7760,N_8701);
nand U9379 (N_9379,N_8447,N_8443);
nor U9380 (N_9380,N_8929,N_8811);
or U9381 (N_9381,N_8534,N_8582);
nor U9382 (N_9382,N_8371,N_8894);
or U9383 (N_9383,N_8115,N_7846);
and U9384 (N_9384,N_7765,N_7736);
xnor U9385 (N_9385,N_8067,N_7671);
and U9386 (N_9386,N_8943,N_8238);
xor U9387 (N_9387,N_8322,N_7627);
or U9388 (N_9388,N_8525,N_8905);
xor U9389 (N_9389,N_8240,N_8181);
nand U9390 (N_9390,N_7571,N_7789);
or U9391 (N_9391,N_7557,N_8346);
xnor U9392 (N_9392,N_8734,N_8577);
and U9393 (N_9393,N_7937,N_8633);
nand U9394 (N_9394,N_8006,N_8519);
or U9395 (N_9395,N_8916,N_8482);
and U9396 (N_9396,N_7546,N_8966);
nand U9397 (N_9397,N_8376,N_7737);
nor U9398 (N_9398,N_8953,N_8794);
nand U9399 (N_9399,N_8150,N_8901);
and U9400 (N_9400,N_8377,N_7503);
xnor U9401 (N_9401,N_8892,N_8492);
nor U9402 (N_9402,N_7845,N_8909);
or U9403 (N_9403,N_8180,N_8578);
or U9404 (N_9404,N_8999,N_8077);
nand U9405 (N_9405,N_8355,N_8250);
or U9406 (N_9406,N_8252,N_7610);
nor U9407 (N_9407,N_8375,N_8356);
nand U9408 (N_9408,N_7584,N_8097);
nand U9409 (N_9409,N_8998,N_7721);
nor U9410 (N_9410,N_8947,N_7548);
xor U9411 (N_9411,N_8670,N_7918);
nand U9412 (N_9412,N_8489,N_7655);
xnor U9413 (N_9413,N_8004,N_8028);
or U9414 (N_9414,N_8585,N_8526);
nand U9415 (N_9415,N_7517,N_8914);
xnor U9416 (N_9416,N_8110,N_8513);
and U9417 (N_9417,N_8433,N_8972);
or U9418 (N_9418,N_8331,N_7543);
or U9419 (N_9419,N_8783,N_8564);
and U9420 (N_9420,N_7867,N_7934);
or U9421 (N_9421,N_8865,N_8967);
nand U9422 (N_9422,N_8142,N_8021);
nand U9423 (N_9423,N_8344,N_7908);
xnor U9424 (N_9424,N_8792,N_7775);
and U9425 (N_9425,N_8727,N_8752);
xnor U9426 (N_9426,N_8949,N_8782);
nor U9427 (N_9427,N_7959,N_8399);
and U9428 (N_9428,N_7781,N_7617);
nand U9429 (N_9429,N_7706,N_8218);
xnor U9430 (N_9430,N_8131,N_8530);
nand U9431 (N_9431,N_7987,N_7653);
xnor U9432 (N_9432,N_8227,N_8112);
xnor U9433 (N_9433,N_8301,N_8883);
nor U9434 (N_9434,N_7597,N_7974);
nor U9435 (N_9435,N_8956,N_7622);
xor U9436 (N_9436,N_8829,N_8466);
xnor U9437 (N_9437,N_8511,N_7834);
nor U9438 (N_9438,N_8915,N_8946);
xnor U9439 (N_9439,N_8818,N_8855);
xor U9440 (N_9440,N_7954,N_8621);
and U9441 (N_9441,N_7620,N_7713);
nand U9442 (N_9442,N_8857,N_8758);
and U9443 (N_9443,N_7674,N_8993);
and U9444 (N_9444,N_7656,N_8845);
or U9445 (N_9445,N_7817,N_7835);
and U9446 (N_9446,N_7744,N_8602);
xor U9447 (N_9447,N_8056,N_8955);
or U9448 (N_9448,N_8853,N_8460);
xor U9449 (N_9449,N_8259,N_7971);
nand U9450 (N_9450,N_7794,N_8725);
xnor U9451 (N_9451,N_7536,N_7692);
nand U9452 (N_9452,N_8851,N_8451);
nor U9453 (N_9453,N_8844,N_8964);
and U9454 (N_9454,N_8389,N_8961);
and U9455 (N_9455,N_8944,N_7969);
xnor U9456 (N_9456,N_8440,N_8823);
or U9457 (N_9457,N_8100,N_8037);
and U9458 (N_9458,N_8164,N_7753);
nand U9459 (N_9459,N_8339,N_8467);
nor U9460 (N_9460,N_7762,N_8514);
or U9461 (N_9461,N_8553,N_8912);
or U9462 (N_9462,N_8323,N_8313);
nor U9463 (N_9463,N_7886,N_8739);
and U9464 (N_9464,N_7673,N_8076);
nand U9465 (N_9465,N_8870,N_8361);
xnor U9466 (N_9466,N_8072,N_7505);
nor U9467 (N_9467,N_7941,N_8628);
or U9468 (N_9468,N_7569,N_8816);
and U9469 (N_9469,N_8058,N_7973);
xor U9470 (N_9470,N_7677,N_8620);
nor U9471 (N_9471,N_8132,N_8776);
xnor U9472 (N_9472,N_8114,N_8994);
nand U9473 (N_9473,N_7644,N_8068);
nor U9474 (N_9474,N_7519,N_7783);
and U9475 (N_9475,N_8900,N_7556);
nand U9476 (N_9476,N_7608,N_7902);
or U9477 (N_9477,N_8085,N_8793);
xnor U9478 (N_9478,N_8876,N_8623);
xnor U9479 (N_9479,N_8295,N_8141);
and U9480 (N_9480,N_8691,N_8304);
or U9481 (N_9481,N_8531,N_8234);
nand U9482 (N_9482,N_8625,N_7946);
or U9483 (N_9483,N_7593,N_8441);
nor U9484 (N_9484,N_8590,N_8454);
xor U9485 (N_9485,N_8583,N_8570);
nor U9486 (N_9486,N_8309,N_8760);
nand U9487 (N_9487,N_8435,N_8805);
nand U9488 (N_9488,N_8658,N_8566);
xnor U9489 (N_9489,N_8817,N_8023);
xnor U9490 (N_9490,N_8412,N_8255);
or U9491 (N_9491,N_7865,N_8959);
xor U9492 (N_9492,N_7964,N_8502);
xor U9493 (N_9493,N_8305,N_8277);
nand U9494 (N_9494,N_8161,N_7560);
xor U9495 (N_9495,N_7769,N_8939);
or U9496 (N_9496,N_8821,N_8410);
and U9497 (N_9497,N_8090,N_8151);
and U9498 (N_9498,N_8289,N_7690);
nand U9499 (N_9499,N_7883,N_8260);
and U9500 (N_9500,N_8178,N_8515);
or U9501 (N_9501,N_8951,N_8195);
or U9502 (N_9502,N_8035,N_8971);
nand U9503 (N_9503,N_8996,N_7559);
xor U9504 (N_9504,N_8824,N_7696);
xnor U9505 (N_9505,N_8196,N_7723);
nor U9506 (N_9506,N_8200,N_7889);
nor U9507 (N_9507,N_7863,N_8494);
and U9508 (N_9508,N_8278,N_8952);
and U9509 (N_9509,N_8439,N_7788);
nand U9510 (N_9510,N_7913,N_8122);
nor U9511 (N_9511,N_8091,N_8631);
nand U9512 (N_9512,N_7595,N_8481);
or U9513 (N_9513,N_8856,N_7684);
nor U9514 (N_9514,N_8655,N_7590);
and U9515 (N_9515,N_7819,N_7935);
xor U9516 (N_9516,N_8567,N_8597);
nor U9517 (N_9517,N_7772,N_8755);
or U9518 (N_9518,N_8868,N_7960);
and U9519 (N_9519,N_8689,N_8543);
and U9520 (N_9520,N_7607,N_8493);
nand U9521 (N_9521,N_8902,N_8744);
xnor U9522 (N_9522,N_8697,N_8970);
nor U9523 (N_9523,N_8191,N_8071);
or U9524 (N_9524,N_7777,N_8318);
xor U9525 (N_9525,N_7927,N_8992);
nor U9526 (N_9526,N_8768,N_8400);
xor U9527 (N_9527,N_8925,N_8074);
nand U9528 (N_9528,N_7586,N_8624);
and U9529 (N_9529,N_8707,N_8815);
or U9530 (N_9530,N_8236,N_8764);
nand U9531 (N_9531,N_7825,N_7895);
or U9532 (N_9532,N_8274,N_8437);
or U9533 (N_9533,N_8709,N_8647);
xor U9534 (N_9534,N_8014,N_7660);
nand U9535 (N_9535,N_8974,N_8504);
nor U9536 (N_9536,N_8417,N_8796);
and U9537 (N_9537,N_7664,N_8413);
or U9538 (N_9538,N_8172,N_8109);
and U9539 (N_9539,N_7646,N_8257);
or U9540 (N_9540,N_7669,N_8229);
nor U9541 (N_9541,N_7703,N_8632);
and U9542 (N_9542,N_8579,N_7709);
or U9543 (N_9543,N_7968,N_8107);
nor U9544 (N_9544,N_8860,N_8940);
or U9545 (N_9545,N_8299,N_8027);
xor U9546 (N_9546,N_8995,N_8731);
nor U9547 (N_9547,N_8551,N_7616);
or U9548 (N_9548,N_8183,N_8478);
nor U9549 (N_9549,N_7957,N_8736);
nand U9550 (N_9550,N_7890,N_7739);
xnor U9551 (N_9551,N_8759,N_7527);
xor U9552 (N_9552,N_7564,N_8918);
or U9553 (N_9553,N_8166,N_8922);
nor U9554 (N_9554,N_8189,N_7589);
and U9555 (N_9555,N_8005,N_8350);
and U9556 (N_9556,N_8168,N_8048);
nand U9557 (N_9557,N_7583,N_7843);
nand U9558 (N_9558,N_8283,N_8116);
or U9559 (N_9559,N_8980,N_7790);
and U9560 (N_9560,N_8199,N_8656);
xnor U9561 (N_9561,N_8668,N_7958);
nor U9562 (N_9562,N_8948,N_8040);
nor U9563 (N_9563,N_7828,N_7899);
nor U9564 (N_9564,N_8046,N_7717);
nand U9565 (N_9565,N_8745,N_7691);
xor U9566 (N_9566,N_7884,N_7734);
xnor U9567 (N_9567,N_7921,N_8386);
or U9568 (N_9568,N_8660,N_8927);
nand U9569 (N_9569,N_7962,N_7811);
nand U9570 (N_9570,N_8193,N_8875);
and U9571 (N_9571,N_8119,N_7567);
xor U9572 (N_9572,N_8791,N_8275);
nor U9573 (N_9573,N_8458,N_7751);
nand U9574 (N_9574,N_8380,N_8474);
and U9575 (N_9575,N_8785,N_8556);
xor U9576 (N_9576,N_8031,N_8558);
and U9577 (N_9577,N_8030,N_8616);
nor U9578 (N_9578,N_8819,N_8281);
xor U9579 (N_9579,N_8547,N_8986);
nor U9580 (N_9580,N_8171,N_8635);
xor U9581 (N_9581,N_8136,N_8589);
and U9582 (N_9582,N_8170,N_8837);
xor U9583 (N_9583,N_8780,N_8982);
or U9584 (N_9584,N_8111,N_8290);
and U9585 (N_9585,N_8497,N_7748);
or U9586 (N_9586,N_7940,N_8264);
xnor U9587 (N_9587,N_7827,N_8212);
or U9588 (N_9588,N_8987,N_8485);
xor U9589 (N_9589,N_8469,N_8517);
and U9590 (N_9590,N_7990,N_8886);
or U9591 (N_9591,N_8532,N_8833);
xnor U9592 (N_9592,N_8406,N_7808);
nand U9593 (N_9593,N_8148,N_7821);
and U9594 (N_9594,N_7592,N_8273);
nand U9595 (N_9595,N_8020,N_8276);
and U9596 (N_9596,N_8480,N_8847);
nor U9597 (N_9597,N_8047,N_8287);
or U9598 (N_9598,N_7936,N_8057);
or U9599 (N_9599,N_8983,N_7779);
nor U9600 (N_9600,N_8026,N_8288);
nor U9601 (N_9601,N_7991,N_8500);
and U9602 (N_9602,N_8848,N_7956);
and U9603 (N_9603,N_7729,N_8612);
xor U9604 (N_9604,N_7950,N_7910);
nor U9605 (N_9605,N_8416,N_7982);
or U9606 (N_9606,N_8253,N_7855);
nor U9607 (N_9607,N_7679,N_7826);
nor U9608 (N_9608,N_7963,N_8398);
nand U9609 (N_9609,N_8675,N_7562);
or U9610 (N_9610,N_8544,N_8319);
or U9611 (N_9611,N_8617,N_8895);
and U9612 (N_9612,N_8728,N_8214);
xnor U9613 (N_9613,N_8153,N_8419);
xor U9614 (N_9614,N_8527,N_7640);
xnor U9615 (N_9615,N_8104,N_8197);
nor U9616 (N_9616,N_7805,N_8850);
or U9617 (N_9617,N_8968,N_8003);
xor U9618 (N_9618,N_8379,N_8352);
and U9619 (N_9619,N_8154,N_8169);
nand U9620 (N_9620,N_8714,N_8677);
nor U9621 (N_9621,N_8384,N_8372);
nor U9622 (N_9622,N_7606,N_8721);
nor U9623 (N_9623,N_7800,N_8307);
nand U9624 (N_9624,N_8618,N_7810);
nand U9625 (N_9625,N_7907,N_8157);
or U9626 (N_9626,N_8232,N_8385);
nor U9627 (N_9627,N_8888,N_8538);
and U9628 (N_9628,N_7704,N_8724);
and U9629 (N_9629,N_8799,N_8495);
or U9630 (N_9630,N_8146,N_8066);
nand U9631 (N_9631,N_7844,N_8904);
nand U9632 (N_9632,N_7763,N_7741);
and U9633 (N_9633,N_7735,N_8438);
nand U9634 (N_9634,N_8124,N_8840);
nand U9635 (N_9635,N_7645,N_8672);
or U9636 (N_9636,N_8931,N_8061);
and U9637 (N_9637,N_8889,N_8459);
xor U9638 (N_9638,N_8268,N_8942);
xnor U9639 (N_9639,N_8858,N_8347);
and U9640 (N_9640,N_8520,N_8615);
and U9641 (N_9641,N_7904,N_7731);
xor U9642 (N_9642,N_7755,N_8007);
or U9643 (N_9643,N_8797,N_7612);
or U9644 (N_9644,N_8358,N_7594);
xnor U9645 (N_9645,N_8568,N_8893);
and U9646 (N_9646,N_7578,N_8266);
xnor U9647 (N_9647,N_8190,N_8751);
nand U9648 (N_9648,N_7791,N_8881);
nand U9649 (N_9649,N_8251,N_8702);
or U9650 (N_9650,N_8921,N_7650);
xnor U9651 (N_9651,N_8561,N_8973);
or U9652 (N_9652,N_7864,N_8684);
nor U9653 (N_9653,N_7615,N_7979);
nand U9654 (N_9654,N_8296,N_7625);
and U9655 (N_9655,N_7643,N_8033);
xor U9656 (N_9656,N_7900,N_8644);
nor U9657 (N_9657,N_8863,N_8708);
xnor U9658 (N_9658,N_8770,N_8756);
and U9659 (N_9659,N_8761,N_8397);
and U9660 (N_9660,N_8711,N_8671);
or U9661 (N_9661,N_7947,N_8297);
or U9662 (N_9662,N_8700,N_7572);
nor U9663 (N_9663,N_7876,N_8505);
nor U9664 (N_9664,N_8637,N_8950);
xnor U9665 (N_9665,N_7531,N_7551);
nand U9666 (N_9666,N_8835,N_8393);
and U9667 (N_9667,N_8599,N_8430);
and U9668 (N_9668,N_7839,N_8321);
nor U9669 (N_9669,N_7905,N_8064);
nor U9670 (N_9670,N_8101,N_7604);
xor U9671 (N_9671,N_7520,N_7774);
and U9672 (N_9672,N_7582,N_7795);
nand U9673 (N_9673,N_8923,N_7980);
xor U9674 (N_9674,N_8303,N_8695);
and U9675 (N_9675,N_7529,N_7804);
or U9676 (N_9676,N_8217,N_7942);
nand U9677 (N_9677,N_7978,N_8117);
nor U9678 (N_9678,N_8795,N_8215);
or U9679 (N_9679,N_7780,N_8859);
and U9680 (N_9680,N_7632,N_8562);
nor U9681 (N_9681,N_8394,N_8742);
nor U9682 (N_9682,N_7528,N_7710);
or U9683 (N_9683,N_8135,N_8043);
xor U9684 (N_9684,N_8825,N_8324);
or U9685 (N_9685,N_8436,N_8779);
nand U9686 (N_9686,N_8694,N_7787);
or U9687 (N_9687,N_8882,N_8917);
and U9688 (N_9688,N_8581,N_7711);
xnor U9689 (N_9689,N_7880,N_8374);
or U9690 (N_9690,N_8401,N_8126);
or U9691 (N_9691,N_8669,N_8763);
and U9692 (N_9692,N_8666,N_8501);
or U9693 (N_9693,N_8261,N_8880);
xor U9694 (N_9694,N_8609,N_7948);
nand U9695 (N_9695,N_8332,N_7754);
or U9696 (N_9696,N_8741,N_7841);
nand U9697 (N_9697,N_7688,N_8349);
nand U9698 (N_9698,N_7881,N_7896);
and U9699 (N_9699,N_8535,N_8053);
nor U9700 (N_9700,N_8411,N_7816);
and U9701 (N_9701,N_8069,N_7682);
or U9702 (N_9702,N_8075,N_8798);
or U9703 (N_9703,N_7575,N_8813);
or U9704 (N_9704,N_8012,N_8749);
xor U9705 (N_9705,N_8936,N_8607);
xnor U9706 (N_9706,N_8446,N_8192);
and U9707 (N_9707,N_8484,N_8338);
nor U9708 (N_9708,N_7837,N_7747);
nand U9709 (N_9709,N_7745,N_7510);
and U9710 (N_9710,N_8113,N_8681);
nor U9711 (N_9711,N_8418,N_8937);
xor U9712 (N_9712,N_8409,N_7818);
nor U9713 (N_9713,N_8849,N_8248);
nand U9714 (N_9714,N_8720,N_7924);
nor U9715 (N_9715,N_7928,N_8729);
or U9716 (N_9716,N_8228,N_8233);
nand U9717 (N_9717,N_8159,N_7882);
or U9718 (N_9718,N_8010,N_8187);
xnor U9719 (N_9719,N_7539,N_7533);
nand U9720 (N_9720,N_8683,N_7892);
xor U9721 (N_9721,N_8420,N_8130);
and U9722 (N_9722,N_8083,N_8291);
nand U9723 (N_9723,N_7574,N_8444);
nor U9724 (N_9724,N_8861,N_8041);
and U9725 (N_9725,N_7756,N_8102);
or U9726 (N_9726,N_8018,N_8286);
nor U9727 (N_9727,N_7518,N_8843);
or U9728 (N_9728,N_8890,N_7538);
nand U9729 (N_9729,N_7563,N_7750);
nor U9730 (N_9730,N_7995,N_8846);
xnor U9731 (N_9731,N_8643,N_8442);
nand U9732 (N_9732,N_8935,N_8265);
nor U9733 (N_9733,N_8800,N_8559);
xnor U9734 (N_9734,N_7730,N_8226);
xnor U9735 (N_9735,N_8604,N_8093);
and U9736 (N_9736,N_8608,N_7752);
and U9737 (N_9737,N_8424,N_8016);
nand U9738 (N_9738,N_8934,N_8008);
nand U9739 (N_9739,N_8654,N_8382);
nand U9740 (N_9740,N_8310,N_8471);
or U9741 (N_9741,N_7535,N_7860);
nor U9742 (N_9742,N_8345,N_7915);
nor U9743 (N_9743,N_8054,N_8476);
and U9744 (N_9744,N_7931,N_7672);
nand U9745 (N_9745,N_8246,N_8488);
nor U9746 (N_9746,N_7678,N_8879);
nor U9747 (N_9747,N_7806,N_8387);
xnor U9748 (N_9748,N_7903,N_7636);
and U9749 (N_9749,N_8327,N_7842);
and U9750 (N_9750,N_8512,N_8045);
xor U9751 (N_9751,N_7724,N_8077);
or U9752 (N_9752,N_8630,N_7573);
and U9753 (N_9753,N_7715,N_7782);
and U9754 (N_9754,N_7610,N_8104);
xor U9755 (N_9755,N_7978,N_8852);
or U9756 (N_9756,N_7918,N_8393);
xor U9757 (N_9757,N_7782,N_8925);
nor U9758 (N_9758,N_8680,N_8762);
or U9759 (N_9759,N_8081,N_8146);
nand U9760 (N_9760,N_7676,N_7612);
or U9761 (N_9761,N_8997,N_7830);
xor U9762 (N_9762,N_8787,N_8558);
or U9763 (N_9763,N_7983,N_8998);
nor U9764 (N_9764,N_7566,N_8196);
or U9765 (N_9765,N_7779,N_8389);
nor U9766 (N_9766,N_7629,N_7981);
and U9767 (N_9767,N_8542,N_7959);
nor U9768 (N_9768,N_7648,N_8153);
xnor U9769 (N_9769,N_8268,N_7641);
xnor U9770 (N_9770,N_7515,N_8047);
xnor U9771 (N_9771,N_8500,N_7660);
and U9772 (N_9772,N_7821,N_7697);
xor U9773 (N_9773,N_8390,N_8322);
xor U9774 (N_9774,N_8487,N_8591);
nand U9775 (N_9775,N_7617,N_8599);
xnor U9776 (N_9776,N_8551,N_8305);
and U9777 (N_9777,N_7914,N_8940);
or U9778 (N_9778,N_8468,N_7651);
or U9779 (N_9779,N_8610,N_7844);
and U9780 (N_9780,N_7981,N_8656);
nand U9781 (N_9781,N_8934,N_8268);
xnor U9782 (N_9782,N_8611,N_8695);
xnor U9783 (N_9783,N_8957,N_8938);
and U9784 (N_9784,N_8354,N_8001);
or U9785 (N_9785,N_8582,N_7798);
xor U9786 (N_9786,N_8440,N_8268);
nand U9787 (N_9787,N_7661,N_8391);
nor U9788 (N_9788,N_8163,N_8470);
nor U9789 (N_9789,N_8508,N_8693);
or U9790 (N_9790,N_7588,N_8442);
nand U9791 (N_9791,N_7807,N_8704);
nor U9792 (N_9792,N_8206,N_7993);
nor U9793 (N_9793,N_7859,N_7947);
or U9794 (N_9794,N_8277,N_7671);
nand U9795 (N_9795,N_8985,N_8717);
or U9796 (N_9796,N_8544,N_8043);
and U9797 (N_9797,N_7957,N_8823);
nor U9798 (N_9798,N_7574,N_8792);
or U9799 (N_9799,N_8280,N_7981);
and U9800 (N_9800,N_8257,N_8164);
nor U9801 (N_9801,N_8529,N_8808);
and U9802 (N_9802,N_8928,N_8887);
nand U9803 (N_9803,N_8960,N_7826);
nand U9804 (N_9804,N_8807,N_7958);
xnor U9805 (N_9805,N_7807,N_8718);
and U9806 (N_9806,N_8610,N_8978);
xor U9807 (N_9807,N_8454,N_7669);
and U9808 (N_9808,N_8711,N_7633);
or U9809 (N_9809,N_8537,N_8289);
or U9810 (N_9810,N_8473,N_7723);
nor U9811 (N_9811,N_7865,N_7916);
or U9812 (N_9812,N_8764,N_8727);
nand U9813 (N_9813,N_7635,N_8510);
nor U9814 (N_9814,N_8437,N_8822);
nand U9815 (N_9815,N_7598,N_8445);
nor U9816 (N_9816,N_7802,N_7716);
and U9817 (N_9817,N_8456,N_8930);
and U9818 (N_9818,N_8379,N_8430);
and U9819 (N_9819,N_8288,N_8598);
and U9820 (N_9820,N_7567,N_8137);
nor U9821 (N_9821,N_8375,N_7748);
or U9822 (N_9822,N_7959,N_8825);
and U9823 (N_9823,N_8622,N_7818);
nor U9824 (N_9824,N_7511,N_8819);
nor U9825 (N_9825,N_8237,N_8117);
and U9826 (N_9826,N_7599,N_7738);
xor U9827 (N_9827,N_8038,N_8110);
nand U9828 (N_9828,N_8596,N_7629);
xor U9829 (N_9829,N_8532,N_8058);
xnor U9830 (N_9830,N_8624,N_8057);
nand U9831 (N_9831,N_8622,N_8352);
or U9832 (N_9832,N_8189,N_8024);
xor U9833 (N_9833,N_7675,N_7828);
or U9834 (N_9834,N_7960,N_8241);
nor U9835 (N_9835,N_8999,N_7852);
or U9836 (N_9836,N_7901,N_7534);
nand U9837 (N_9837,N_8365,N_7666);
xor U9838 (N_9838,N_7581,N_7670);
xnor U9839 (N_9839,N_8036,N_8676);
nor U9840 (N_9840,N_8389,N_8745);
xnor U9841 (N_9841,N_8866,N_8539);
or U9842 (N_9842,N_8662,N_8529);
nor U9843 (N_9843,N_8130,N_8809);
xnor U9844 (N_9844,N_7830,N_8802);
nor U9845 (N_9845,N_8651,N_8543);
xnor U9846 (N_9846,N_7641,N_8480);
nor U9847 (N_9847,N_8526,N_7956);
or U9848 (N_9848,N_7758,N_8019);
xnor U9849 (N_9849,N_7713,N_7848);
nor U9850 (N_9850,N_8843,N_8489);
nor U9851 (N_9851,N_8351,N_7604);
and U9852 (N_9852,N_7851,N_8083);
or U9853 (N_9853,N_8125,N_8184);
xor U9854 (N_9854,N_8156,N_8981);
nor U9855 (N_9855,N_8500,N_8145);
and U9856 (N_9856,N_8866,N_8183);
xnor U9857 (N_9857,N_8764,N_7633);
and U9858 (N_9858,N_8013,N_8607);
or U9859 (N_9859,N_8349,N_8640);
nor U9860 (N_9860,N_7978,N_8713);
nand U9861 (N_9861,N_7863,N_8559);
xnor U9862 (N_9862,N_7972,N_8134);
and U9863 (N_9863,N_8611,N_8364);
xnor U9864 (N_9864,N_8331,N_7714);
nor U9865 (N_9865,N_8276,N_8283);
or U9866 (N_9866,N_8410,N_7727);
nor U9867 (N_9867,N_8404,N_8861);
or U9868 (N_9868,N_7506,N_8694);
xnor U9869 (N_9869,N_7594,N_8964);
nand U9870 (N_9870,N_8638,N_7641);
nor U9871 (N_9871,N_8459,N_8213);
or U9872 (N_9872,N_7974,N_8668);
and U9873 (N_9873,N_8610,N_7657);
nand U9874 (N_9874,N_8009,N_7852);
or U9875 (N_9875,N_7633,N_8281);
xnor U9876 (N_9876,N_8326,N_8555);
and U9877 (N_9877,N_8607,N_8782);
nand U9878 (N_9878,N_7799,N_7868);
xnor U9879 (N_9879,N_8679,N_7723);
xnor U9880 (N_9880,N_8675,N_8265);
or U9881 (N_9881,N_8980,N_7641);
or U9882 (N_9882,N_8061,N_8740);
nand U9883 (N_9883,N_8836,N_7569);
xor U9884 (N_9884,N_7948,N_8737);
xnor U9885 (N_9885,N_8222,N_8989);
and U9886 (N_9886,N_8698,N_8080);
xnor U9887 (N_9887,N_8505,N_7983);
or U9888 (N_9888,N_8088,N_8472);
or U9889 (N_9889,N_8473,N_8131);
nand U9890 (N_9890,N_7614,N_7647);
xor U9891 (N_9891,N_8438,N_7888);
and U9892 (N_9892,N_7692,N_8219);
nand U9893 (N_9893,N_7910,N_7717);
xor U9894 (N_9894,N_8309,N_8669);
or U9895 (N_9895,N_8200,N_8987);
and U9896 (N_9896,N_8171,N_7989);
or U9897 (N_9897,N_8583,N_7932);
or U9898 (N_9898,N_8708,N_8453);
nor U9899 (N_9899,N_8108,N_8558);
xor U9900 (N_9900,N_8626,N_8764);
nor U9901 (N_9901,N_8140,N_7564);
and U9902 (N_9902,N_8936,N_8514);
xnor U9903 (N_9903,N_8110,N_8588);
and U9904 (N_9904,N_8891,N_8949);
or U9905 (N_9905,N_8104,N_8173);
and U9906 (N_9906,N_7608,N_8714);
nor U9907 (N_9907,N_8344,N_8470);
nand U9908 (N_9908,N_8305,N_8743);
nor U9909 (N_9909,N_7627,N_8538);
nor U9910 (N_9910,N_7675,N_8630);
and U9911 (N_9911,N_7728,N_8302);
and U9912 (N_9912,N_7709,N_8504);
nand U9913 (N_9913,N_8483,N_8601);
and U9914 (N_9914,N_8016,N_8954);
and U9915 (N_9915,N_8820,N_7844);
nor U9916 (N_9916,N_7660,N_8883);
or U9917 (N_9917,N_8048,N_7576);
xor U9918 (N_9918,N_8614,N_7732);
xor U9919 (N_9919,N_8481,N_7571);
nand U9920 (N_9920,N_8973,N_7880);
nor U9921 (N_9921,N_8466,N_8941);
or U9922 (N_9922,N_8839,N_8821);
nand U9923 (N_9923,N_8868,N_8317);
nor U9924 (N_9924,N_7696,N_8130);
and U9925 (N_9925,N_8411,N_7885);
and U9926 (N_9926,N_8244,N_8180);
and U9927 (N_9927,N_7606,N_8596);
nand U9928 (N_9928,N_7965,N_8820);
or U9929 (N_9929,N_8125,N_8588);
and U9930 (N_9930,N_8564,N_8829);
or U9931 (N_9931,N_8098,N_7905);
xnor U9932 (N_9932,N_7559,N_7531);
and U9933 (N_9933,N_8028,N_8309);
and U9934 (N_9934,N_7898,N_8334);
and U9935 (N_9935,N_8941,N_7635);
or U9936 (N_9936,N_8907,N_8988);
nand U9937 (N_9937,N_7767,N_8225);
nand U9938 (N_9938,N_8865,N_8603);
nand U9939 (N_9939,N_8924,N_8765);
xnor U9940 (N_9940,N_8679,N_8689);
nand U9941 (N_9941,N_8237,N_7840);
or U9942 (N_9942,N_7601,N_8479);
and U9943 (N_9943,N_7957,N_8652);
and U9944 (N_9944,N_8554,N_7725);
and U9945 (N_9945,N_8541,N_8161);
xnor U9946 (N_9946,N_8323,N_7949);
nor U9947 (N_9947,N_8960,N_8761);
xnor U9948 (N_9948,N_8290,N_8856);
and U9949 (N_9949,N_8172,N_8211);
and U9950 (N_9950,N_7861,N_8646);
nand U9951 (N_9951,N_8331,N_8403);
xor U9952 (N_9952,N_7631,N_8863);
and U9953 (N_9953,N_8220,N_8243);
nor U9954 (N_9954,N_8010,N_8990);
and U9955 (N_9955,N_8805,N_8725);
and U9956 (N_9956,N_8090,N_7582);
nand U9957 (N_9957,N_8175,N_8153);
xnor U9958 (N_9958,N_8343,N_7839);
and U9959 (N_9959,N_8528,N_8178);
or U9960 (N_9960,N_7857,N_7786);
nor U9961 (N_9961,N_8219,N_8904);
xnor U9962 (N_9962,N_8471,N_7798);
or U9963 (N_9963,N_7730,N_7806);
nor U9964 (N_9964,N_7539,N_8634);
xnor U9965 (N_9965,N_8477,N_8575);
or U9966 (N_9966,N_8551,N_7664);
nor U9967 (N_9967,N_8537,N_7701);
or U9968 (N_9968,N_8212,N_7836);
and U9969 (N_9969,N_8055,N_8889);
and U9970 (N_9970,N_7682,N_8762);
and U9971 (N_9971,N_8273,N_7975);
xor U9972 (N_9972,N_7834,N_8386);
nor U9973 (N_9973,N_8824,N_8386);
and U9974 (N_9974,N_8109,N_8876);
xnor U9975 (N_9975,N_8820,N_7770);
or U9976 (N_9976,N_7579,N_7652);
nand U9977 (N_9977,N_8679,N_7579);
nor U9978 (N_9978,N_8199,N_8672);
or U9979 (N_9979,N_7877,N_8662);
nor U9980 (N_9980,N_8217,N_8278);
and U9981 (N_9981,N_8039,N_7587);
or U9982 (N_9982,N_7620,N_7621);
and U9983 (N_9983,N_8239,N_8917);
xor U9984 (N_9984,N_7771,N_7895);
or U9985 (N_9985,N_8885,N_8815);
xnor U9986 (N_9986,N_8681,N_8400);
xor U9987 (N_9987,N_8028,N_8612);
xnor U9988 (N_9988,N_8241,N_8586);
nor U9989 (N_9989,N_8041,N_8664);
nand U9990 (N_9990,N_8098,N_8778);
xnor U9991 (N_9991,N_8118,N_7728);
or U9992 (N_9992,N_8230,N_8635);
or U9993 (N_9993,N_8676,N_7956);
and U9994 (N_9994,N_8614,N_8965);
nand U9995 (N_9995,N_8621,N_8171);
and U9996 (N_9996,N_7500,N_8571);
xnor U9997 (N_9997,N_7832,N_8079);
and U9998 (N_9998,N_7743,N_8576);
and U9999 (N_9999,N_8024,N_8273);
and U10000 (N_10000,N_8997,N_8284);
and U10001 (N_10001,N_7607,N_7569);
xor U10002 (N_10002,N_8764,N_7833);
or U10003 (N_10003,N_8474,N_8457);
nor U10004 (N_10004,N_7792,N_8584);
nor U10005 (N_10005,N_8378,N_8323);
and U10006 (N_10006,N_8542,N_7549);
nand U10007 (N_10007,N_8356,N_8116);
and U10008 (N_10008,N_7568,N_7832);
and U10009 (N_10009,N_8134,N_8587);
or U10010 (N_10010,N_8303,N_8523);
and U10011 (N_10011,N_7500,N_7746);
xor U10012 (N_10012,N_8351,N_8333);
nand U10013 (N_10013,N_8291,N_7613);
nor U10014 (N_10014,N_8234,N_8436);
or U10015 (N_10015,N_8955,N_8240);
or U10016 (N_10016,N_8294,N_8725);
or U10017 (N_10017,N_8088,N_8007);
and U10018 (N_10018,N_8327,N_8834);
nand U10019 (N_10019,N_8581,N_7684);
nand U10020 (N_10020,N_8531,N_8697);
nor U10021 (N_10021,N_7877,N_7549);
nor U10022 (N_10022,N_8905,N_8163);
nand U10023 (N_10023,N_8046,N_7623);
xor U10024 (N_10024,N_7916,N_8612);
or U10025 (N_10025,N_8564,N_7532);
xor U10026 (N_10026,N_8924,N_7994);
nor U10027 (N_10027,N_8604,N_7506);
nand U10028 (N_10028,N_8054,N_7543);
nor U10029 (N_10029,N_7500,N_8787);
nand U10030 (N_10030,N_8723,N_8115);
or U10031 (N_10031,N_7828,N_8776);
nand U10032 (N_10032,N_7934,N_8466);
or U10033 (N_10033,N_7642,N_8463);
or U10034 (N_10034,N_7981,N_8031);
or U10035 (N_10035,N_8620,N_7537);
and U10036 (N_10036,N_8054,N_8336);
xnor U10037 (N_10037,N_8187,N_8022);
and U10038 (N_10038,N_8639,N_8173);
nor U10039 (N_10039,N_8001,N_7753);
nand U10040 (N_10040,N_8406,N_8825);
nand U10041 (N_10041,N_7957,N_7649);
nand U10042 (N_10042,N_7863,N_8805);
nor U10043 (N_10043,N_8444,N_8731);
nand U10044 (N_10044,N_8189,N_8943);
nand U10045 (N_10045,N_8186,N_7959);
and U10046 (N_10046,N_7520,N_8048);
nor U10047 (N_10047,N_7691,N_7988);
nor U10048 (N_10048,N_8426,N_7746);
and U10049 (N_10049,N_7510,N_7797);
or U10050 (N_10050,N_8307,N_7883);
xnor U10051 (N_10051,N_8473,N_8015);
xor U10052 (N_10052,N_8335,N_8299);
or U10053 (N_10053,N_8432,N_8759);
or U10054 (N_10054,N_8747,N_8839);
and U10055 (N_10055,N_8040,N_8173);
xor U10056 (N_10056,N_8772,N_8765);
and U10057 (N_10057,N_7973,N_8043);
nor U10058 (N_10058,N_8445,N_8053);
nand U10059 (N_10059,N_8021,N_8965);
or U10060 (N_10060,N_8911,N_7588);
nor U10061 (N_10061,N_8387,N_7604);
and U10062 (N_10062,N_7896,N_8631);
nand U10063 (N_10063,N_8533,N_7763);
or U10064 (N_10064,N_8483,N_8136);
xnor U10065 (N_10065,N_7983,N_7900);
nand U10066 (N_10066,N_7971,N_8409);
and U10067 (N_10067,N_8101,N_8589);
xor U10068 (N_10068,N_8761,N_7752);
nand U10069 (N_10069,N_7894,N_8997);
nand U10070 (N_10070,N_8352,N_7842);
and U10071 (N_10071,N_8380,N_8319);
xor U10072 (N_10072,N_8563,N_8763);
xor U10073 (N_10073,N_8887,N_8468);
and U10074 (N_10074,N_8234,N_8994);
nor U10075 (N_10075,N_8905,N_7528);
nand U10076 (N_10076,N_8673,N_7656);
and U10077 (N_10077,N_8395,N_8562);
xnor U10078 (N_10078,N_8875,N_8349);
xnor U10079 (N_10079,N_8097,N_7825);
xor U10080 (N_10080,N_7712,N_7611);
and U10081 (N_10081,N_8011,N_7965);
and U10082 (N_10082,N_7580,N_8001);
or U10083 (N_10083,N_8393,N_7605);
nor U10084 (N_10084,N_7733,N_8437);
xnor U10085 (N_10085,N_8098,N_8699);
nand U10086 (N_10086,N_7612,N_7682);
xnor U10087 (N_10087,N_8087,N_7562);
nor U10088 (N_10088,N_8331,N_8660);
nor U10089 (N_10089,N_8376,N_8292);
or U10090 (N_10090,N_7844,N_8947);
xor U10091 (N_10091,N_8912,N_8677);
nand U10092 (N_10092,N_8968,N_8874);
or U10093 (N_10093,N_8263,N_8138);
and U10094 (N_10094,N_8718,N_7840);
xor U10095 (N_10095,N_7619,N_8005);
or U10096 (N_10096,N_7973,N_8537);
xnor U10097 (N_10097,N_8077,N_8203);
xor U10098 (N_10098,N_7821,N_8898);
or U10099 (N_10099,N_8823,N_8419);
xor U10100 (N_10100,N_8474,N_8349);
nand U10101 (N_10101,N_7857,N_7866);
and U10102 (N_10102,N_8548,N_8793);
nor U10103 (N_10103,N_8591,N_7566);
or U10104 (N_10104,N_8260,N_8105);
or U10105 (N_10105,N_8926,N_8591);
and U10106 (N_10106,N_8449,N_8404);
nor U10107 (N_10107,N_7627,N_8581);
nand U10108 (N_10108,N_8155,N_8540);
xnor U10109 (N_10109,N_7740,N_8206);
xor U10110 (N_10110,N_8937,N_8057);
or U10111 (N_10111,N_7792,N_7939);
nor U10112 (N_10112,N_8013,N_8966);
and U10113 (N_10113,N_8578,N_7535);
and U10114 (N_10114,N_7613,N_7780);
or U10115 (N_10115,N_7876,N_8641);
and U10116 (N_10116,N_7511,N_8784);
nor U10117 (N_10117,N_7935,N_8660);
xor U10118 (N_10118,N_8339,N_8086);
nor U10119 (N_10119,N_7804,N_8999);
and U10120 (N_10120,N_7665,N_8691);
or U10121 (N_10121,N_8249,N_8009);
and U10122 (N_10122,N_8269,N_8272);
nand U10123 (N_10123,N_8181,N_7705);
xnor U10124 (N_10124,N_8871,N_8860);
xor U10125 (N_10125,N_8524,N_8764);
and U10126 (N_10126,N_8571,N_8805);
xnor U10127 (N_10127,N_8985,N_7994);
and U10128 (N_10128,N_7607,N_8500);
or U10129 (N_10129,N_7541,N_8512);
xor U10130 (N_10130,N_7675,N_8429);
nor U10131 (N_10131,N_7883,N_8031);
or U10132 (N_10132,N_8291,N_7742);
or U10133 (N_10133,N_8597,N_7796);
nor U10134 (N_10134,N_7708,N_7669);
nand U10135 (N_10135,N_8099,N_7889);
xor U10136 (N_10136,N_8458,N_8581);
xor U10137 (N_10137,N_8541,N_8481);
xor U10138 (N_10138,N_8120,N_8294);
or U10139 (N_10139,N_7579,N_7868);
and U10140 (N_10140,N_8927,N_8433);
and U10141 (N_10141,N_8475,N_8467);
nand U10142 (N_10142,N_8077,N_8760);
xor U10143 (N_10143,N_7560,N_8787);
nand U10144 (N_10144,N_7960,N_7850);
and U10145 (N_10145,N_8762,N_7929);
or U10146 (N_10146,N_7517,N_8703);
nand U10147 (N_10147,N_7948,N_7566);
nand U10148 (N_10148,N_8367,N_8350);
nand U10149 (N_10149,N_8904,N_8206);
or U10150 (N_10150,N_7864,N_8685);
xnor U10151 (N_10151,N_8112,N_8704);
and U10152 (N_10152,N_8716,N_8037);
xor U10153 (N_10153,N_8438,N_8542);
nand U10154 (N_10154,N_7787,N_8844);
and U10155 (N_10155,N_8501,N_8643);
nor U10156 (N_10156,N_8429,N_8285);
xnor U10157 (N_10157,N_7823,N_7834);
and U10158 (N_10158,N_8916,N_7931);
nand U10159 (N_10159,N_8987,N_8094);
nor U10160 (N_10160,N_8873,N_7860);
or U10161 (N_10161,N_8834,N_8065);
xnor U10162 (N_10162,N_8003,N_8301);
nand U10163 (N_10163,N_8858,N_8248);
xnor U10164 (N_10164,N_8565,N_8658);
and U10165 (N_10165,N_8696,N_8959);
xnor U10166 (N_10166,N_8595,N_8549);
and U10167 (N_10167,N_8777,N_8983);
nor U10168 (N_10168,N_8083,N_8977);
xor U10169 (N_10169,N_8238,N_7617);
or U10170 (N_10170,N_7775,N_8189);
xnor U10171 (N_10171,N_8682,N_7821);
or U10172 (N_10172,N_8158,N_8573);
or U10173 (N_10173,N_8672,N_7595);
xor U10174 (N_10174,N_8486,N_8575);
xor U10175 (N_10175,N_8433,N_7675);
nand U10176 (N_10176,N_8982,N_8381);
or U10177 (N_10177,N_8376,N_7979);
nor U10178 (N_10178,N_8469,N_7823);
or U10179 (N_10179,N_7781,N_8691);
and U10180 (N_10180,N_7701,N_7725);
and U10181 (N_10181,N_8424,N_8191);
or U10182 (N_10182,N_8610,N_8201);
xnor U10183 (N_10183,N_7832,N_8191);
xnor U10184 (N_10184,N_8956,N_7795);
or U10185 (N_10185,N_8778,N_8193);
nand U10186 (N_10186,N_8179,N_7704);
or U10187 (N_10187,N_8308,N_7852);
and U10188 (N_10188,N_7940,N_8806);
nor U10189 (N_10189,N_8742,N_8834);
and U10190 (N_10190,N_8819,N_7853);
or U10191 (N_10191,N_7827,N_8841);
and U10192 (N_10192,N_8815,N_8989);
nand U10193 (N_10193,N_8715,N_7989);
and U10194 (N_10194,N_7827,N_8514);
and U10195 (N_10195,N_8712,N_8350);
xor U10196 (N_10196,N_8174,N_8537);
xnor U10197 (N_10197,N_8723,N_7611);
xnor U10198 (N_10198,N_8373,N_8892);
xor U10199 (N_10199,N_8504,N_8797);
nand U10200 (N_10200,N_8661,N_7632);
or U10201 (N_10201,N_8845,N_7792);
nand U10202 (N_10202,N_8204,N_8472);
nand U10203 (N_10203,N_8586,N_8545);
and U10204 (N_10204,N_8391,N_8914);
or U10205 (N_10205,N_7992,N_8080);
xor U10206 (N_10206,N_8617,N_7693);
or U10207 (N_10207,N_7653,N_8420);
and U10208 (N_10208,N_8393,N_7950);
xor U10209 (N_10209,N_8082,N_8508);
xnor U10210 (N_10210,N_8416,N_8540);
nor U10211 (N_10211,N_8080,N_8344);
nor U10212 (N_10212,N_8303,N_8716);
xor U10213 (N_10213,N_8301,N_8532);
nand U10214 (N_10214,N_8158,N_8530);
or U10215 (N_10215,N_8742,N_8599);
nand U10216 (N_10216,N_7996,N_8147);
nand U10217 (N_10217,N_8240,N_7521);
nand U10218 (N_10218,N_7997,N_8714);
nand U10219 (N_10219,N_7982,N_8049);
nand U10220 (N_10220,N_7671,N_8020);
or U10221 (N_10221,N_8141,N_8937);
or U10222 (N_10222,N_8632,N_7660);
and U10223 (N_10223,N_8617,N_8667);
or U10224 (N_10224,N_7667,N_7640);
or U10225 (N_10225,N_7768,N_8676);
nor U10226 (N_10226,N_8654,N_8869);
nand U10227 (N_10227,N_7694,N_7754);
and U10228 (N_10228,N_7697,N_8438);
and U10229 (N_10229,N_8082,N_8887);
and U10230 (N_10230,N_8475,N_8298);
or U10231 (N_10231,N_8223,N_8850);
nor U10232 (N_10232,N_8914,N_7562);
nor U10233 (N_10233,N_8772,N_8127);
and U10234 (N_10234,N_8779,N_8923);
or U10235 (N_10235,N_7963,N_8188);
nand U10236 (N_10236,N_8171,N_8074);
or U10237 (N_10237,N_7906,N_7644);
and U10238 (N_10238,N_8764,N_8456);
or U10239 (N_10239,N_7722,N_7942);
or U10240 (N_10240,N_7995,N_8505);
nor U10241 (N_10241,N_8777,N_8544);
or U10242 (N_10242,N_8390,N_8991);
xor U10243 (N_10243,N_8516,N_8504);
nand U10244 (N_10244,N_8619,N_7770);
nor U10245 (N_10245,N_7649,N_7882);
or U10246 (N_10246,N_8536,N_7515);
and U10247 (N_10247,N_7592,N_8683);
xor U10248 (N_10248,N_8529,N_8213);
and U10249 (N_10249,N_8417,N_8060);
nor U10250 (N_10250,N_8874,N_7556);
xnor U10251 (N_10251,N_8620,N_8720);
and U10252 (N_10252,N_7829,N_7915);
xor U10253 (N_10253,N_8330,N_7700);
or U10254 (N_10254,N_8989,N_7693);
or U10255 (N_10255,N_8520,N_8183);
nor U10256 (N_10256,N_8001,N_8190);
nand U10257 (N_10257,N_8677,N_7863);
nand U10258 (N_10258,N_8660,N_8382);
or U10259 (N_10259,N_8924,N_8305);
or U10260 (N_10260,N_7794,N_7798);
nor U10261 (N_10261,N_8540,N_8300);
xor U10262 (N_10262,N_7525,N_8175);
nand U10263 (N_10263,N_8043,N_7604);
nor U10264 (N_10264,N_8815,N_7827);
xor U10265 (N_10265,N_8061,N_8934);
and U10266 (N_10266,N_8910,N_7912);
or U10267 (N_10267,N_8305,N_8690);
and U10268 (N_10268,N_8590,N_8183);
nor U10269 (N_10269,N_8417,N_8811);
and U10270 (N_10270,N_8925,N_7536);
or U10271 (N_10271,N_8411,N_7795);
nor U10272 (N_10272,N_7949,N_8005);
xnor U10273 (N_10273,N_8438,N_8867);
or U10274 (N_10274,N_8855,N_8622);
or U10275 (N_10275,N_7956,N_7824);
nor U10276 (N_10276,N_8515,N_8026);
nor U10277 (N_10277,N_8037,N_8592);
or U10278 (N_10278,N_8760,N_7793);
and U10279 (N_10279,N_8163,N_8349);
nand U10280 (N_10280,N_8551,N_8751);
nand U10281 (N_10281,N_8697,N_7805);
nor U10282 (N_10282,N_7604,N_8293);
nand U10283 (N_10283,N_7862,N_8088);
and U10284 (N_10284,N_8308,N_7756);
and U10285 (N_10285,N_8179,N_7949);
xnor U10286 (N_10286,N_7654,N_7662);
nand U10287 (N_10287,N_8300,N_8571);
and U10288 (N_10288,N_8705,N_8913);
nand U10289 (N_10289,N_7978,N_8569);
nor U10290 (N_10290,N_8989,N_8138);
nand U10291 (N_10291,N_8891,N_8083);
or U10292 (N_10292,N_8845,N_8691);
nor U10293 (N_10293,N_8203,N_8288);
nor U10294 (N_10294,N_8377,N_7532);
or U10295 (N_10295,N_7991,N_7612);
nor U10296 (N_10296,N_8631,N_8230);
or U10297 (N_10297,N_8854,N_8670);
xor U10298 (N_10298,N_7827,N_8627);
xor U10299 (N_10299,N_8394,N_7578);
nor U10300 (N_10300,N_8563,N_8719);
and U10301 (N_10301,N_8487,N_7516);
nor U10302 (N_10302,N_8730,N_8343);
xnor U10303 (N_10303,N_8443,N_7647);
nor U10304 (N_10304,N_7684,N_8264);
or U10305 (N_10305,N_8362,N_7838);
xor U10306 (N_10306,N_7506,N_7878);
or U10307 (N_10307,N_7579,N_8534);
or U10308 (N_10308,N_7541,N_8073);
and U10309 (N_10309,N_7895,N_7598);
and U10310 (N_10310,N_8184,N_8584);
xor U10311 (N_10311,N_8569,N_8340);
or U10312 (N_10312,N_7579,N_8022);
and U10313 (N_10313,N_8863,N_8574);
or U10314 (N_10314,N_7800,N_8352);
nand U10315 (N_10315,N_8883,N_7868);
and U10316 (N_10316,N_7687,N_8964);
and U10317 (N_10317,N_8299,N_7674);
xnor U10318 (N_10318,N_7855,N_8373);
or U10319 (N_10319,N_8031,N_7551);
nand U10320 (N_10320,N_8309,N_8903);
nand U10321 (N_10321,N_7565,N_8415);
xor U10322 (N_10322,N_7833,N_8746);
xor U10323 (N_10323,N_8888,N_7991);
xnor U10324 (N_10324,N_8976,N_8663);
or U10325 (N_10325,N_8741,N_8780);
nand U10326 (N_10326,N_7760,N_8515);
xnor U10327 (N_10327,N_8962,N_8693);
nor U10328 (N_10328,N_8531,N_8821);
and U10329 (N_10329,N_8941,N_7586);
nor U10330 (N_10330,N_8405,N_7540);
xnor U10331 (N_10331,N_8401,N_7809);
or U10332 (N_10332,N_8625,N_8917);
nor U10333 (N_10333,N_8477,N_7744);
xnor U10334 (N_10334,N_8248,N_7919);
nor U10335 (N_10335,N_8585,N_8622);
nand U10336 (N_10336,N_8459,N_8882);
nand U10337 (N_10337,N_8912,N_8544);
nor U10338 (N_10338,N_8629,N_7815);
nor U10339 (N_10339,N_8576,N_8378);
nand U10340 (N_10340,N_7836,N_8925);
nor U10341 (N_10341,N_7935,N_8561);
xor U10342 (N_10342,N_8432,N_7596);
and U10343 (N_10343,N_8398,N_8926);
xor U10344 (N_10344,N_8929,N_8988);
or U10345 (N_10345,N_8388,N_7535);
and U10346 (N_10346,N_8498,N_8390);
nand U10347 (N_10347,N_7792,N_7871);
or U10348 (N_10348,N_8229,N_8152);
nor U10349 (N_10349,N_8439,N_8958);
or U10350 (N_10350,N_8476,N_8993);
and U10351 (N_10351,N_8282,N_8463);
or U10352 (N_10352,N_8062,N_7527);
nor U10353 (N_10353,N_8512,N_8108);
or U10354 (N_10354,N_7528,N_7875);
and U10355 (N_10355,N_8304,N_8821);
nand U10356 (N_10356,N_8127,N_7752);
nand U10357 (N_10357,N_7545,N_8360);
xor U10358 (N_10358,N_7668,N_8945);
and U10359 (N_10359,N_8847,N_7838);
or U10360 (N_10360,N_8749,N_8879);
nor U10361 (N_10361,N_8075,N_8350);
or U10362 (N_10362,N_7848,N_8142);
or U10363 (N_10363,N_8247,N_8796);
xnor U10364 (N_10364,N_7643,N_8745);
nor U10365 (N_10365,N_8080,N_7911);
nand U10366 (N_10366,N_8994,N_8439);
nand U10367 (N_10367,N_7589,N_7723);
nor U10368 (N_10368,N_7930,N_8425);
xor U10369 (N_10369,N_8461,N_8740);
or U10370 (N_10370,N_8284,N_8613);
xnor U10371 (N_10371,N_7882,N_8085);
and U10372 (N_10372,N_8103,N_8801);
or U10373 (N_10373,N_7854,N_8222);
nand U10374 (N_10374,N_8513,N_8984);
or U10375 (N_10375,N_8786,N_8949);
nand U10376 (N_10376,N_7953,N_8502);
or U10377 (N_10377,N_8109,N_8907);
or U10378 (N_10378,N_7721,N_8761);
xnor U10379 (N_10379,N_8480,N_8096);
nand U10380 (N_10380,N_8770,N_8737);
or U10381 (N_10381,N_8147,N_8887);
nor U10382 (N_10382,N_8451,N_8622);
and U10383 (N_10383,N_8313,N_8245);
nand U10384 (N_10384,N_8688,N_8321);
or U10385 (N_10385,N_8601,N_8014);
and U10386 (N_10386,N_8058,N_7823);
xnor U10387 (N_10387,N_7837,N_7898);
nor U10388 (N_10388,N_8663,N_7694);
xor U10389 (N_10389,N_8882,N_7526);
nor U10390 (N_10390,N_8846,N_7915);
xor U10391 (N_10391,N_8905,N_7753);
and U10392 (N_10392,N_8180,N_7914);
xor U10393 (N_10393,N_7558,N_8929);
nand U10394 (N_10394,N_7620,N_8466);
nor U10395 (N_10395,N_8700,N_7709);
nand U10396 (N_10396,N_8826,N_7966);
or U10397 (N_10397,N_8209,N_8362);
nor U10398 (N_10398,N_8310,N_7796);
nor U10399 (N_10399,N_8886,N_8847);
xor U10400 (N_10400,N_7593,N_7881);
nor U10401 (N_10401,N_7577,N_8412);
xnor U10402 (N_10402,N_8018,N_8044);
and U10403 (N_10403,N_8793,N_8724);
or U10404 (N_10404,N_8873,N_8785);
nand U10405 (N_10405,N_7516,N_7661);
or U10406 (N_10406,N_8974,N_7729);
and U10407 (N_10407,N_8972,N_7975);
and U10408 (N_10408,N_8749,N_8287);
and U10409 (N_10409,N_7771,N_8694);
and U10410 (N_10410,N_8863,N_7687);
or U10411 (N_10411,N_8877,N_7882);
and U10412 (N_10412,N_8469,N_7564);
nand U10413 (N_10413,N_8113,N_8588);
nor U10414 (N_10414,N_8512,N_8347);
or U10415 (N_10415,N_8903,N_8436);
nand U10416 (N_10416,N_8944,N_8982);
and U10417 (N_10417,N_7595,N_7965);
and U10418 (N_10418,N_7691,N_8404);
nor U10419 (N_10419,N_8357,N_8119);
or U10420 (N_10420,N_8446,N_7774);
xor U10421 (N_10421,N_8501,N_8071);
xor U10422 (N_10422,N_7845,N_8961);
and U10423 (N_10423,N_7736,N_7741);
and U10424 (N_10424,N_8537,N_8010);
xnor U10425 (N_10425,N_8579,N_8344);
nand U10426 (N_10426,N_8004,N_7842);
and U10427 (N_10427,N_7809,N_8002);
xor U10428 (N_10428,N_7763,N_7575);
and U10429 (N_10429,N_8865,N_8430);
nand U10430 (N_10430,N_8540,N_8973);
and U10431 (N_10431,N_8282,N_8869);
or U10432 (N_10432,N_8166,N_8018);
nand U10433 (N_10433,N_8621,N_8414);
or U10434 (N_10434,N_7810,N_8200);
and U10435 (N_10435,N_7928,N_7717);
or U10436 (N_10436,N_7798,N_8783);
nor U10437 (N_10437,N_7567,N_8227);
nand U10438 (N_10438,N_8364,N_8110);
or U10439 (N_10439,N_8866,N_7773);
and U10440 (N_10440,N_8010,N_7651);
xor U10441 (N_10441,N_8452,N_7756);
nor U10442 (N_10442,N_7845,N_8065);
and U10443 (N_10443,N_7947,N_8139);
and U10444 (N_10444,N_7825,N_7663);
nor U10445 (N_10445,N_8625,N_8794);
or U10446 (N_10446,N_8948,N_8529);
or U10447 (N_10447,N_8424,N_8020);
nand U10448 (N_10448,N_8990,N_7634);
xnor U10449 (N_10449,N_8501,N_7804);
and U10450 (N_10450,N_8959,N_8579);
nor U10451 (N_10451,N_8910,N_8357);
or U10452 (N_10452,N_8855,N_7951);
or U10453 (N_10453,N_8574,N_8705);
or U10454 (N_10454,N_8231,N_7723);
and U10455 (N_10455,N_7915,N_8921);
nand U10456 (N_10456,N_8546,N_8463);
nand U10457 (N_10457,N_8677,N_8956);
nand U10458 (N_10458,N_8005,N_8322);
xnor U10459 (N_10459,N_8412,N_7987);
nor U10460 (N_10460,N_8998,N_8406);
and U10461 (N_10461,N_8525,N_7507);
nor U10462 (N_10462,N_8995,N_8327);
nor U10463 (N_10463,N_8349,N_8523);
nand U10464 (N_10464,N_8850,N_7736);
nor U10465 (N_10465,N_8158,N_8602);
xor U10466 (N_10466,N_8967,N_8546);
nand U10467 (N_10467,N_8131,N_8480);
xnor U10468 (N_10468,N_8485,N_8472);
xnor U10469 (N_10469,N_7680,N_8155);
nor U10470 (N_10470,N_8616,N_7876);
nand U10471 (N_10471,N_8813,N_7844);
nor U10472 (N_10472,N_8629,N_7977);
xor U10473 (N_10473,N_7866,N_8985);
nand U10474 (N_10474,N_8612,N_7646);
or U10475 (N_10475,N_8578,N_8584);
nand U10476 (N_10476,N_8774,N_7733);
nand U10477 (N_10477,N_7657,N_8284);
nand U10478 (N_10478,N_7805,N_8970);
and U10479 (N_10479,N_7741,N_7969);
xnor U10480 (N_10480,N_8897,N_8381);
xor U10481 (N_10481,N_8260,N_8122);
or U10482 (N_10482,N_7626,N_8920);
xor U10483 (N_10483,N_8261,N_8661);
nand U10484 (N_10484,N_8934,N_8986);
and U10485 (N_10485,N_8193,N_7692);
nor U10486 (N_10486,N_8301,N_8861);
xor U10487 (N_10487,N_7950,N_7966);
nand U10488 (N_10488,N_8547,N_8687);
and U10489 (N_10489,N_8751,N_7823);
nor U10490 (N_10490,N_8983,N_8316);
and U10491 (N_10491,N_7780,N_7966);
and U10492 (N_10492,N_8367,N_7999);
xnor U10493 (N_10493,N_8250,N_7728);
and U10494 (N_10494,N_8221,N_7813);
or U10495 (N_10495,N_8428,N_8796);
nor U10496 (N_10496,N_8020,N_7553);
or U10497 (N_10497,N_7793,N_8465);
nor U10498 (N_10498,N_8165,N_7560);
xnor U10499 (N_10499,N_8531,N_8176);
or U10500 (N_10500,N_10008,N_9806);
xor U10501 (N_10501,N_9556,N_9099);
and U10502 (N_10502,N_9329,N_9561);
nand U10503 (N_10503,N_9490,N_9448);
or U10504 (N_10504,N_10430,N_9557);
or U10505 (N_10505,N_9343,N_9546);
and U10506 (N_10506,N_10344,N_9920);
nand U10507 (N_10507,N_10465,N_10437);
nor U10508 (N_10508,N_10161,N_9152);
nand U10509 (N_10509,N_10179,N_9446);
or U10510 (N_10510,N_10387,N_9381);
or U10511 (N_10511,N_10115,N_10258);
nor U10512 (N_10512,N_9312,N_9819);
and U10513 (N_10513,N_9271,N_10325);
or U10514 (N_10514,N_10025,N_9229);
xnor U10515 (N_10515,N_9307,N_9670);
or U10516 (N_10516,N_9379,N_10353);
and U10517 (N_10517,N_10201,N_9209);
and U10518 (N_10518,N_10034,N_10094);
nand U10519 (N_10519,N_9757,N_10475);
or U10520 (N_10520,N_9019,N_9413);
nor U10521 (N_10521,N_9097,N_9979);
nor U10522 (N_10522,N_9440,N_9130);
nor U10523 (N_10523,N_9380,N_9762);
nor U10524 (N_10524,N_9200,N_9435);
or U10525 (N_10525,N_9080,N_9974);
xor U10526 (N_10526,N_9710,N_9746);
or U10527 (N_10527,N_10333,N_9215);
nand U10528 (N_10528,N_9189,N_9374);
or U10529 (N_10529,N_10020,N_9454);
xnor U10530 (N_10530,N_9277,N_10436);
and U10531 (N_10531,N_10454,N_9754);
nor U10532 (N_10532,N_9989,N_9947);
xor U10533 (N_10533,N_10260,N_10379);
xnor U10534 (N_10534,N_10184,N_10269);
or U10535 (N_10535,N_10375,N_9980);
nand U10536 (N_10536,N_9079,N_9709);
and U10537 (N_10537,N_10164,N_9437);
or U10538 (N_10538,N_10399,N_9639);
and U10539 (N_10539,N_9694,N_9999);
or U10540 (N_10540,N_10239,N_10048);
xor U10541 (N_10541,N_9664,N_10172);
nor U10542 (N_10542,N_9933,N_9216);
xor U10543 (N_10543,N_9264,N_9081);
xor U10544 (N_10544,N_10187,N_9239);
and U10545 (N_10545,N_9993,N_10147);
and U10546 (N_10546,N_9958,N_10204);
nand U10547 (N_10547,N_9011,N_9839);
nor U10548 (N_10548,N_9513,N_9112);
and U10549 (N_10549,N_9320,N_10494);
nor U10550 (N_10550,N_9175,N_10460);
xnor U10551 (N_10551,N_9100,N_9850);
and U10552 (N_10552,N_10037,N_9953);
nand U10553 (N_10553,N_9549,N_9500);
nor U10554 (N_10554,N_9082,N_9544);
nand U10555 (N_10555,N_9732,N_10116);
or U10556 (N_10556,N_10195,N_10484);
nand U10557 (N_10557,N_10336,N_10256);
nand U10558 (N_10558,N_10095,N_9375);
or U10559 (N_10559,N_9316,N_9144);
nor U10560 (N_10560,N_10284,N_10050);
xnor U10561 (N_10561,N_9140,N_9049);
and U10562 (N_10562,N_10045,N_10408);
xor U10563 (N_10563,N_10428,N_10485);
nand U10564 (N_10564,N_10107,N_9624);
xor U10565 (N_10565,N_10087,N_9625);
or U10566 (N_10566,N_10042,N_9337);
and U10567 (N_10567,N_10218,N_9627);
xor U10568 (N_10568,N_10234,N_10137);
nor U10569 (N_10569,N_9891,N_9445);
and U10570 (N_10570,N_9161,N_9588);
nand U10571 (N_10571,N_9397,N_9996);
or U10572 (N_10572,N_9185,N_10056);
nand U10573 (N_10573,N_9341,N_9118);
or U10574 (N_10574,N_9395,N_9474);
nand U10575 (N_10575,N_9160,N_9038);
nor U10576 (N_10576,N_9815,N_10426);
nand U10577 (N_10577,N_9838,N_9632);
and U10578 (N_10578,N_9062,N_9016);
nand U10579 (N_10579,N_9228,N_9602);
xor U10580 (N_10580,N_10074,N_9044);
nor U10581 (N_10581,N_10182,N_10401);
xor U10582 (N_10582,N_10285,N_9836);
or U10583 (N_10583,N_10031,N_10362);
and U10584 (N_10584,N_9050,N_10466);
and U10585 (N_10585,N_10313,N_9310);
and U10586 (N_10586,N_9998,N_9163);
nor U10587 (N_10587,N_9230,N_9033);
and U10588 (N_10588,N_9027,N_10103);
nand U10589 (N_10589,N_9008,N_10223);
nor U10590 (N_10590,N_9706,N_9467);
or U10591 (N_10591,N_9692,N_9243);
and U10592 (N_10592,N_9906,N_10104);
or U10593 (N_10593,N_9294,N_9018);
nand U10594 (N_10594,N_10470,N_9350);
and U10595 (N_10595,N_10007,N_10487);
or U10596 (N_10596,N_10089,N_10294);
and U10597 (N_10597,N_10091,N_9262);
nor U10598 (N_10598,N_9333,N_10365);
and U10599 (N_10599,N_10127,N_9852);
or U10600 (N_10600,N_9418,N_9897);
and U10601 (N_10601,N_9031,N_10073);
nor U10602 (N_10602,N_9862,N_9761);
nand U10603 (N_10603,N_9325,N_9197);
or U10604 (N_10604,N_9269,N_9314);
nand U10605 (N_10605,N_9499,N_9524);
nor U10606 (N_10606,N_9916,N_10114);
and U10607 (N_10607,N_9505,N_9677);
nand U10608 (N_10608,N_10281,N_9973);
or U10609 (N_10609,N_9537,N_10129);
xnor U10610 (N_10610,N_10273,N_10270);
nor U10611 (N_10611,N_9292,N_9508);
nor U10612 (N_10612,N_10146,N_9076);
xor U10613 (N_10613,N_9957,N_9476);
nand U10614 (N_10614,N_9599,N_9604);
nor U10615 (N_10615,N_9928,N_9988);
xor U10616 (N_10616,N_9948,N_9491);
xor U10617 (N_10617,N_10446,N_9313);
or U10618 (N_10618,N_10210,N_9198);
xor U10619 (N_10619,N_9219,N_10392);
and U10620 (N_10620,N_9309,N_9338);
and U10621 (N_10621,N_10349,N_9117);
xnor U10622 (N_10622,N_10021,N_9914);
or U10623 (N_10623,N_10158,N_9274);
xnor U10624 (N_10624,N_9799,N_9004);
or U10625 (N_10625,N_9816,N_9032);
or U10626 (N_10626,N_10332,N_10493);
or U10627 (N_10627,N_9638,N_9378);
and U10628 (N_10628,N_9558,N_10311);
nand U10629 (N_10629,N_9825,N_9072);
or U10630 (N_10630,N_9360,N_9302);
xnor U10631 (N_10631,N_9103,N_10002);
nand U10632 (N_10632,N_9407,N_9786);
xnor U10633 (N_10633,N_9766,N_10018);
xnor U10634 (N_10634,N_9859,N_10228);
nand U10635 (N_10635,N_10154,N_10183);
or U10636 (N_10636,N_9978,N_9181);
and U10637 (N_10637,N_10192,N_9055);
or U10638 (N_10638,N_9934,N_9365);
nor U10639 (N_10639,N_10383,N_9559);
nand U10640 (N_10640,N_9647,N_9344);
nor U10641 (N_10641,N_9751,N_10326);
or U10642 (N_10642,N_10283,N_9869);
nand U10643 (N_10643,N_9362,N_10377);
and U10644 (N_10644,N_9529,N_9452);
or U10645 (N_10645,N_9811,N_9770);
nand U10646 (N_10646,N_9636,N_9293);
xnor U10647 (N_10647,N_10439,N_9182);
xor U10648 (N_10648,N_9865,N_9719);
and U10649 (N_10649,N_9217,N_9172);
or U10650 (N_10650,N_9077,N_9483);
nand U10651 (N_10651,N_9394,N_9405);
nor U10652 (N_10652,N_10272,N_10355);
xnor U10653 (N_10653,N_9201,N_10105);
nand U10654 (N_10654,N_9183,N_9104);
xnor U10655 (N_10655,N_10134,N_9875);
nor U10656 (N_10656,N_9039,N_9731);
or U10657 (N_10657,N_9823,N_10163);
and U10658 (N_10658,N_9115,N_9346);
and U10659 (N_10659,N_10225,N_10293);
nor U10660 (N_10660,N_9860,N_9401);
xnor U10661 (N_10661,N_9656,N_10479);
nor U10662 (N_10662,N_9439,N_9794);
nor U10663 (N_10663,N_9792,N_9330);
nor U10664 (N_10664,N_10111,N_10345);
xor U10665 (N_10665,N_9901,N_10176);
nor U10666 (N_10666,N_10188,N_9713);
xor U10667 (N_10667,N_9389,N_9841);
nor U10668 (N_10668,N_9699,N_9569);
nand U10669 (N_10669,N_9233,N_9252);
nor U10670 (N_10670,N_9772,N_10099);
xor U10671 (N_10671,N_9940,N_9048);
xnor U10672 (N_10672,N_9258,N_9393);
xnor U10673 (N_10673,N_10062,N_9662);
or U10674 (N_10674,N_10309,N_9619);
or U10675 (N_10675,N_9598,N_10419);
and U10676 (N_10676,N_9937,N_9015);
nor U10677 (N_10677,N_9961,N_9242);
nor U10678 (N_10678,N_9273,N_9773);
xnor U10679 (N_10679,N_10409,N_10429);
nand U10680 (N_10680,N_10122,N_9574);
or U10681 (N_10681,N_9881,N_9226);
or U10682 (N_10682,N_10030,N_10203);
xnor U10683 (N_10683,N_9681,N_9223);
xor U10684 (N_10684,N_10206,N_10453);
and U10685 (N_10685,N_9560,N_9105);
nand U10686 (N_10686,N_9603,N_9297);
nor U10687 (N_10687,N_9725,N_10330);
nand U10688 (N_10688,N_9580,N_9246);
or U10689 (N_10689,N_9923,N_9613);
nor U10690 (N_10690,N_9517,N_10486);
or U10691 (N_10691,N_10120,N_9040);
nand U10692 (N_10692,N_9388,N_10382);
nor U10693 (N_10693,N_10124,N_9892);
and U10694 (N_10694,N_10462,N_9386);
xnor U10695 (N_10695,N_9621,N_10098);
and U10696 (N_10696,N_9615,N_9538);
or U10697 (N_10697,N_9323,N_9495);
nor U10698 (N_10698,N_10075,N_9530);
and U10699 (N_10699,N_9628,N_10067);
and U10700 (N_10700,N_9668,N_10472);
or U10701 (N_10701,N_9275,N_10391);
nand U10702 (N_10702,N_9760,N_9912);
and U10703 (N_10703,N_9506,N_10194);
or U10704 (N_10704,N_9884,N_9340);
nor U10705 (N_10705,N_9141,N_10335);
nand U10706 (N_10706,N_9813,N_9193);
nand U10707 (N_10707,N_9489,N_9856);
nor U10708 (N_10708,N_9543,N_9122);
or U10709 (N_10709,N_9426,N_9114);
nor U10710 (N_10710,N_9473,N_9562);
nor U10711 (N_10711,N_9564,N_10352);
xor U10712 (N_10712,N_9903,N_9465);
xnor U10713 (N_10713,N_10110,N_9113);
xnor U10714 (N_10714,N_9202,N_10354);
or U10715 (N_10715,N_9255,N_9878);
nand U10716 (N_10716,N_9410,N_9449);
nor U10717 (N_10717,N_10029,N_10235);
nand U10718 (N_10718,N_9917,N_10059);
or U10719 (N_10719,N_9600,N_10009);
and U10720 (N_10720,N_9504,N_9204);
or U10721 (N_10721,N_10035,N_9391);
or U10722 (N_10722,N_9463,N_10338);
nand U10723 (N_10723,N_9353,N_9409);
nand U10724 (N_10724,N_9646,N_9817);
nand U10725 (N_10725,N_9643,N_10458);
nand U10726 (N_10726,N_9167,N_9003);
nand U10727 (N_10727,N_10036,N_9990);
nor U10728 (N_10728,N_9190,N_9907);
or U10729 (N_10729,N_10010,N_9651);
or U10730 (N_10730,N_9400,N_10128);
xor U10731 (N_10731,N_9089,N_9475);
nand U10732 (N_10732,N_9868,N_9419);
and U10733 (N_10733,N_10320,N_9013);
or U10734 (N_10734,N_9304,N_9671);
xor U10735 (N_10735,N_9212,N_10144);
or U10736 (N_10736,N_9522,N_9985);
nand U10737 (N_10737,N_9433,N_10226);
nor U10738 (N_10738,N_9567,N_10214);
nand U10739 (N_10739,N_9908,N_9581);
nor U10740 (N_10740,N_10277,N_10019);
or U10741 (N_10741,N_9471,N_10085);
or U10742 (N_10742,N_9095,N_9351);
and U10743 (N_10743,N_9828,N_9359);
nor U10744 (N_10744,N_9047,N_9256);
or U10745 (N_10745,N_10054,N_9837);
nor U10746 (N_10746,N_9871,N_9888);
or U10747 (N_10747,N_9752,N_10456);
and U10748 (N_10748,N_9683,N_10496);
xnor U10749 (N_10749,N_9436,N_9220);
nor U10750 (N_10750,N_10440,N_10003);
nor U10751 (N_10751,N_10431,N_9800);
nor U10752 (N_10752,N_9168,N_10083);
and U10753 (N_10753,N_9139,N_10395);
xor U10754 (N_10754,N_10473,N_9430);
nand U10755 (N_10755,N_9222,N_9371);
nand U10756 (N_10756,N_10425,N_9586);
nand U10757 (N_10757,N_9146,N_9592);
nand U10758 (N_10758,N_10152,N_10422);
or U10759 (N_10759,N_9626,N_9195);
xor U10760 (N_10760,N_9180,N_10334);
nor U10761 (N_10761,N_9834,N_9245);
nand U10762 (N_10762,N_10298,N_10027);
or U10763 (N_10763,N_9648,N_10464);
nor U10764 (N_10764,N_9142,N_9963);
xor U10765 (N_10765,N_9363,N_9879);
and U10766 (N_10766,N_10369,N_10014);
and U10767 (N_10767,N_9976,N_10141);
or U10768 (N_10768,N_10407,N_9824);
nand U10769 (N_10769,N_9518,N_9136);
xor U10770 (N_10770,N_10477,N_9432);
nor U10771 (N_10771,N_9318,N_9131);
or U10772 (N_10772,N_9915,N_9956);
nor U10773 (N_10773,N_9631,N_9753);
and U10774 (N_10774,N_9416,N_9158);
nand U10775 (N_10775,N_9798,N_9895);
nand U10776 (N_10776,N_9864,N_10243);
or U10777 (N_10777,N_10167,N_9241);
and U10778 (N_10778,N_9480,N_9820);
nand U10779 (N_10779,N_10498,N_10230);
and U10780 (N_10780,N_9326,N_10288);
xnor U10781 (N_10781,N_10400,N_9539);
or U10782 (N_10782,N_9286,N_10237);
or U10783 (N_10783,N_9555,N_9411);
nor U10784 (N_10784,N_9120,N_9171);
nand U10785 (N_10785,N_9065,N_9470);
xor U10786 (N_10786,N_9654,N_10471);
nor U10787 (N_10787,N_10046,N_9166);
and U10788 (N_10788,N_9263,N_9675);
or U10789 (N_10789,N_9462,N_9342);
nand U10790 (N_10790,N_9285,N_9116);
nor U10791 (N_10791,N_10271,N_9810);
xor U10792 (N_10792,N_9296,N_9455);
and U10793 (N_10793,N_10079,N_9279);
nor U10794 (N_10794,N_9165,N_9650);
xnor U10795 (N_10795,N_9857,N_10165);
and U10796 (N_10796,N_9431,N_10121);
nor U10797 (N_10797,N_9087,N_9074);
or U10798 (N_10798,N_9578,N_9265);
or U10799 (N_10799,N_9938,N_9069);
and U10800 (N_10800,N_9899,N_10255);
xnor U10801 (N_10801,N_10451,N_9855);
xor U10802 (N_10802,N_9403,N_10199);
xnor U10803 (N_10803,N_9024,N_9300);
nand U10804 (N_10804,N_10337,N_9067);
and U10805 (N_10805,N_9637,N_10489);
nor U10806 (N_10806,N_9020,N_10312);
nor U10807 (N_10807,N_10457,N_9696);
xnor U10808 (N_10808,N_9162,N_10495);
xnor U10809 (N_10809,N_9644,N_9744);
and U10810 (N_10810,N_9579,N_9488);
nor U10811 (N_10811,N_9147,N_10308);
or U10812 (N_10812,N_9485,N_9248);
nor U10813 (N_10813,N_9234,N_9053);
and U10814 (N_10814,N_10213,N_9102);
or U10815 (N_10815,N_10178,N_9657);
or U10816 (N_10816,N_9601,N_9034);
nor U10817 (N_10817,N_10300,N_9494);
xnor U10818 (N_10818,N_9932,N_9863);
and U10819 (N_10819,N_9306,N_10236);
or U10820 (N_10820,N_9968,N_10278);
xor U10821 (N_10821,N_10295,N_9383);
xnor U10822 (N_10822,N_9807,N_10343);
nor U10823 (N_10823,N_9390,N_10424);
xor U10824 (N_10824,N_10219,N_9714);
or U10825 (N_10825,N_9704,N_10126);
xnor U10826 (N_10826,N_10394,N_9225);
nor U10827 (N_10827,N_9686,N_10467);
or U10828 (N_10828,N_9666,N_10434);
or U10829 (N_10829,N_9966,N_9553);
and U10830 (N_10830,N_9291,N_9481);
nor U10831 (N_10831,N_9459,N_9127);
and U10832 (N_10832,N_10069,N_10497);
and U10833 (N_10833,N_9712,N_9482);
nor U10834 (N_10834,N_9697,N_9520);
and U10835 (N_10835,N_9640,N_10038);
nand U10836 (N_10836,N_10197,N_9918);
or U10837 (N_10837,N_9691,N_9213);
and U10838 (N_10838,N_9612,N_10314);
nor U10839 (N_10839,N_9620,N_10372);
nand U10840 (N_10840,N_9420,N_10291);
xnor U10841 (N_10841,N_9883,N_9573);
nand U10842 (N_10842,N_10322,N_9781);
xnor U10843 (N_10843,N_9121,N_10052);
and U10844 (N_10844,N_10060,N_9597);
and U10845 (N_10845,N_9428,N_10414);
or U10846 (N_10846,N_10367,N_10044);
nand U10847 (N_10847,N_9835,N_9594);
or U10848 (N_10848,N_9023,N_9108);
xor U10849 (N_10849,N_10357,N_9874);
and U10850 (N_10850,N_9649,N_10043);
nor U10851 (N_10851,N_9808,N_9177);
xnor U10852 (N_10852,N_9005,N_9098);
xnor U10853 (N_10853,N_10371,N_10171);
and U10854 (N_10854,N_9443,N_9355);
and U10855 (N_10855,N_10156,N_9926);
nor U10856 (N_10856,N_9398,N_10403);
or U10857 (N_10857,N_9715,N_10202);
nor U10858 (N_10858,N_10101,N_9231);
nand U10859 (N_10859,N_9844,N_9126);
or U10860 (N_10860,N_9521,N_9610);
xnor U10861 (N_10861,N_10323,N_9060);
and U10862 (N_10862,N_9042,N_9930);
xnor U10863 (N_10863,N_10358,N_9145);
and U10864 (N_10864,N_10246,N_10024);
nand U10865 (N_10865,N_9965,N_9669);
nor U10866 (N_10866,N_9893,N_9111);
and U10867 (N_10867,N_10339,N_9991);
nor U10868 (N_10868,N_9373,N_9073);
or U10869 (N_10869,N_9137,N_9345);
and U10870 (N_10870,N_9913,N_9191);
xor U10871 (N_10871,N_9187,N_9516);
xnor U10872 (N_10872,N_10445,N_10132);
xnor U10873 (N_10873,N_9756,N_10315);
nor U10874 (N_10874,N_9154,N_10212);
and U10875 (N_10875,N_10096,N_9605);
xnor U10876 (N_10876,N_9995,N_10448);
or U10877 (N_10877,N_9030,N_9526);
nor U10878 (N_10878,N_9818,N_9469);
xor U10879 (N_10879,N_9525,N_10398);
and U10880 (N_10880,N_10118,N_10265);
nor U10881 (N_10881,N_9339,N_9791);
nand U10882 (N_10882,N_9421,N_9583);
and U10883 (N_10883,N_9925,N_9290);
and U10884 (N_10884,N_10274,N_9955);
and U10885 (N_10885,N_9509,N_10380);
nand U10886 (N_10886,N_9944,N_9203);
nor U10887 (N_10887,N_9498,N_10415);
or U10888 (N_10888,N_9025,N_10081);
and U10889 (N_10889,N_9960,N_10469);
nand U10890 (N_10890,N_9571,N_9106);
nor U10891 (N_10891,N_9540,N_10148);
nand U10892 (N_10892,N_9964,N_9851);
xnor U10893 (N_10893,N_9422,N_9853);
or U10894 (N_10894,N_10181,N_10480);
xor U10895 (N_10895,N_10254,N_10209);
nand U10896 (N_10896,N_9550,N_10193);
nand U10897 (N_10897,N_9251,N_9678);
nor U10898 (N_10898,N_9829,N_9214);
nor U10899 (N_10899,N_9037,N_9970);
xnor U10900 (N_10900,N_9737,N_9478);
nand U10901 (N_10901,N_9684,N_9584);
or U10902 (N_10902,N_9890,N_9000);
nor U10903 (N_10903,N_10488,N_10447);
or U10904 (N_10904,N_10262,N_9809);
xor U10905 (N_10905,N_9867,N_9332);
nor U10906 (N_10906,N_10138,N_10061);
nor U10907 (N_10907,N_9858,N_10442);
and U10908 (N_10908,N_9797,N_10376);
nand U10909 (N_10909,N_9924,N_10013);
and U10910 (N_10910,N_9493,N_9542);
or U10911 (N_10911,N_9563,N_9028);
xor U10912 (N_10912,N_9789,N_9009);
and U10913 (N_10913,N_10175,N_10396);
or U10914 (N_10914,N_10109,N_10170);
or U10915 (N_10915,N_10249,N_9845);
and U10916 (N_10916,N_9250,N_9464);
nand U10917 (N_10917,N_10282,N_9184);
and U10918 (N_10918,N_9589,N_9492);
xor U10919 (N_10919,N_9240,N_9268);
and U10920 (N_10920,N_10160,N_9922);
nor U10921 (N_10921,N_9457,N_9460);
or U10922 (N_10922,N_9477,N_10289);
nor U10923 (N_10923,N_9259,N_10402);
xor U10924 (N_10924,N_10065,N_9745);
and U10925 (N_10925,N_9660,N_9658);
xnor U10926 (N_10926,N_9655,N_9554);
or U10927 (N_10927,N_9758,N_10275);
and U10928 (N_10928,N_10386,N_9535);
or U10929 (N_10929,N_9723,N_9527);
nand U10930 (N_10930,N_10301,N_9531);
nand U10931 (N_10931,N_10420,N_9902);
and U10932 (N_10932,N_9739,N_10198);
and U10933 (N_10933,N_9833,N_9324);
nor U10934 (N_10934,N_9730,N_9790);
or U10935 (N_10935,N_9054,N_9534);
xnor U10936 (N_10936,N_10299,N_9911);
nor U10937 (N_10937,N_10039,N_9425);
nand U10938 (N_10938,N_9528,N_10321);
nor U10939 (N_10939,N_10499,N_10032);
nand U10940 (N_10940,N_9261,N_9063);
nand U10941 (N_10941,N_9919,N_9311);
or U10942 (N_10942,N_10168,N_10017);
nor U10943 (N_10943,N_9986,N_9179);
nor U10944 (N_10944,N_10208,N_9847);
and U10945 (N_10945,N_9969,N_10072);
nor U10946 (N_10946,N_9629,N_10151);
and U10947 (N_10947,N_10055,N_9587);
nand U10948 (N_10948,N_9134,N_9877);
nor U10949 (N_10949,N_10329,N_9734);
nand U10950 (N_10950,N_9576,N_9450);
nor U10951 (N_10951,N_9803,N_9061);
and U10952 (N_10952,N_9497,N_10404);
nor U10953 (N_10953,N_9148,N_9224);
and U10954 (N_10954,N_9981,N_10232);
xnor U10955 (N_10955,N_10106,N_9109);
or U10956 (N_10956,N_9427,N_9910);
nor U10957 (N_10957,N_10304,N_9793);
xor U10958 (N_10958,N_9093,N_9512);
nor U10959 (N_10959,N_9848,N_10241);
or U10960 (N_10960,N_9764,N_9357);
nor U10961 (N_10961,N_9396,N_9367);
and U10962 (N_10962,N_9315,N_9249);
xnor U10963 (N_10963,N_10051,N_9617);
nand U10964 (N_10964,N_9257,N_9994);
and U10965 (N_10965,N_10341,N_9846);
nor U10966 (N_10966,N_10342,N_9633);
or U10967 (N_10967,N_10324,N_9085);
xnor U10968 (N_10968,N_9736,N_10307);
nor U10969 (N_10969,N_9043,N_9523);
nand U10970 (N_10970,N_10443,N_9232);
xor U10971 (N_10971,N_10047,N_9652);
nor U10972 (N_10972,N_9768,N_10108);
nor U10973 (N_10973,N_9741,N_10026);
or U10974 (N_10974,N_9429,N_9412);
and U10975 (N_10975,N_10346,N_10080);
nand U10976 (N_10976,N_9805,N_9444);
and U10977 (N_10977,N_9630,N_10340);
or U10978 (N_10978,N_9110,N_9123);
xor U10979 (N_10979,N_10247,N_10251);
and U10980 (N_10980,N_9987,N_9949);
nor U10981 (N_10981,N_9972,N_9227);
and U10982 (N_10982,N_10427,N_10433);
or U10983 (N_10983,N_10360,N_9236);
nor U10984 (N_10984,N_9690,N_9254);
and U10985 (N_10985,N_9441,N_9173);
nor U10986 (N_10986,N_9176,N_9174);
or U10987 (N_10987,N_9046,N_9585);
or U10988 (N_10988,N_9366,N_10461);
nand U10989 (N_10989,N_9006,N_10410);
nand U10990 (N_10990,N_9788,N_9541);
or U10991 (N_10991,N_9188,N_10390);
nand U10992 (N_10992,N_9515,N_9356);
nand U10993 (N_10993,N_9728,N_9399);
or U10994 (N_10994,N_9572,N_9942);
nand U10995 (N_10995,N_9205,N_9634);
or U10996 (N_10996,N_9207,N_9208);
or U10997 (N_10997,N_9842,N_9336);
nand U10998 (N_10998,N_10476,N_9321);
and U10999 (N_10999,N_9931,N_10366);
xor U11000 (N_11000,N_9186,N_10397);
or U11001 (N_11001,N_9486,N_9308);
xor U11002 (N_11002,N_9361,N_10068);
and U11003 (N_11003,N_9453,N_10016);
or U11004 (N_11004,N_10296,N_9665);
or U11005 (N_11005,N_9716,N_9088);
or U11006 (N_11006,N_9423,N_9950);
xor U11007 (N_11007,N_9107,N_9606);
or U11008 (N_11008,N_9281,N_9078);
or U11009 (N_11009,N_9577,N_9702);
xnor U11010 (N_11010,N_9369,N_10153);
nor U11011 (N_11011,N_9921,N_9717);
xor U11012 (N_11012,N_9724,N_9645);
or U11013 (N_11013,N_10131,N_9056);
or U11014 (N_11014,N_10305,N_9661);
xnor U11015 (N_11015,N_10064,N_9952);
nand U11016 (N_11016,N_10370,N_9849);
and U11017 (N_11017,N_9778,N_10205);
xor U11018 (N_11018,N_10292,N_10250);
nor U11019 (N_11019,N_9083,N_10066);
nor U11020 (N_11020,N_10438,N_10240);
and U11021 (N_11021,N_9726,N_10455);
or U11022 (N_11022,N_9936,N_9503);
nor U11023 (N_11023,N_10173,N_9802);
or U11024 (N_11024,N_9551,N_10364);
xnor U11025 (N_11025,N_9155,N_10418);
and U11026 (N_11026,N_10432,N_9763);
nor U11027 (N_11027,N_10139,N_9663);
nor U11028 (N_11028,N_9532,N_10331);
or U11029 (N_11029,N_10280,N_10006);
xnor U11030 (N_11030,N_10088,N_9347);
or U11031 (N_11031,N_9507,N_10155);
nand U11032 (N_11032,N_9997,N_10263);
xnor U11033 (N_11033,N_10090,N_9830);
and U11034 (N_11034,N_10351,N_9780);
nor U11035 (N_11035,N_9278,N_10190);
xnor U11036 (N_11036,N_9672,N_9718);
or U11037 (N_11037,N_10058,N_10159);
nand U11038 (N_11038,N_10049,N_10022);
and U11039 (N_11039,N_9566,N_9237);
or U11040 (N_11040,N_10452,N_9235);
xor U11041 (N_11041,N_9616,N_9682);
nand U11042 (N_11042,N_10224,N_9461);
xnor U11043 (N_11043,N_10216,N_9959);
nor U11044 (N_11044,N_9607,N_9889);
nor U11045 (N_11045,N_9951,N_9376);
nand U11046 (N_11046,N_10350,N_10186);
and U11047 (N_11047,N_10450,N_10076);
and U11048 (N_11048,N_9064,N_9280);
nor U11049 (N_11049,N_9689,N_9096);
nand U11050 (N_11050,N_9068,N_10449);
nand U11051 (N_11051,N_10416,N_9092);
or U11052 (N_11052,N_10004,N_10063);
or U11053 (N_11053,N_10264,N_9267);
and U11054 (N_11054,N_9880,N_9698);
nand U11055 (N_11055,N_9547,N_9317);
xor U11056 (N_11056,N_10356,N_9748);
or U11057 (N_11057,N_9769,N_9622);
and U11058 (N_11058,N_9707,N_9750);
nand U11059 (N_11059,N_9349,N_10384);
and U11060 (N_11060,N_9733,N_9284);
nand U11061 (N_11061,N_10196,N_9570);
nand U11062 (N_11062,N_9484,N_9687);
or U11063 (N_11063,N_9667,N_9036);
or U11064 (N_11064,N_9001,N_10150);
xor U11065 (N_11065,N_9283,N_9735);
and U11066 (N_11066,N_9017,N_9693);
nor U11067 (N_11067,N_9090,N_9358);
and U11068 (N_11068,N_9084,N_9133);
or U11069 (N_11069,N_10117,N_9676);
and U11070 (N_11070,N_9447,N_9608);
nor U11071 (N_11071,N_10077,N_9695);
nor U11072 (N_11072,N_9623,N_9674);
xnor U11073 (N_11073,N_10421,N_10015);
xor U11074 (N_11074,N_9618,N_10097);
xnor U11075 (N_11075,N_9774,N_10227);
xor U11076 (N_11076,N_9331,N_9295);
nand U11077 (N_11077,N_10220,N_9468);
nor U11078 (N_11078,N_9288,N_9086);
or U11079 (N_11079,N_9272,N_9548);
nand U11080 (N_11080,N_9372,N_9035);
xnor U11081 (N_11081,N_9466,N_9787);
or U11082 (N_11082,N_10347,N_10136);
xor U11083 (N_11083,N_9392,N_9727);
xnor U11084 (N_11084,N_10119,N_10459);
nor U11085 (N_11085,N_10478,N_9635);
xor U11086 (N_11086,N_9496,N_9352);
or U11087 (N_11087,N_9138,N_9124);
nand U11088 (N_11088,N_10406,N_9299);
or U11089 (N_11089,N_9159,N_9832);
nor U11090 (N_11090,N_10238,N_10242);
nor U11091 (N_11091,N_9992,N_9533);
and U11092 (N_11092,N_9238,N_10481);
nand U11093 (N_11093,N_10267,N_9382);
or U11094 (N_11094,N_10200,N_9876);
nand U11095 (N_11095,N_9012,N_10040);
or U11096 (N_11096,N_10435,N_9568);
nor U11097 (N_11097,N_9404,N_9536);
nand U11098 (N_11098,N_9045,N_10302);
nor U11099 (N_11099,N_9010,N_9022);
nand U11100 (N_11100,N_9218,N_10279);
or U11101 (N_11101,N_9059,N_9157);
xor U11102 (N_11102,N_10005,N_9742);
nor U11103 (N_11103,N_10231,N_9552);
or U11104 (N_11104,N_10468,N_9385);
and U11105 (N_11105,N_10215,N_10244);
xor U11106 (N_11106,N_9402,N_9840);
nand U11107 (N_11107,N_10417,N_10229);
xnor U11108 (N_11108,N_9377,N_9821);
xnor U11109 (N_11109,N_9327,N_9886);
nand U11110 (N_11110,N_10303,N_10413);
and U11111 (N_11111,N_9370,N_9711);
nand U11112 (N_11112,N_9775,N_10423);
and U11113 (N_11113,N_10207,N_9927);
nand U11114 (N_11114,N_9861,N_10130);
and U11115 (N_11115,N_9673,N_9747);
nand U11116 (N_11116,N_9685,N_10125);
or U11117 (N_11117,N_10483,N_9070);
and U11118 (N_11118,N_9870,N_9014);
nand U11119 (N_11119,N_10162,N_10185);
nor U11120 (N_11120,N_9354,N_9708);
nand U11121 (N_11121,N_9091,N_9935);
xor U11122 (N_11122,N_10001,N_10028);
nor U11123 (N_11123,N_10222,N_10113);
or U11124 (N_11124,N_9565,N_9156);
xor U11125 (N_11125,N_9143,N_10259);
and U11126 (N_11126,N_9211,N_9782);
and U11127 (N_11127,N_9729,N_9796);
and U11128 (N_11128,N_9700,N_10286);
nor U11129 (N_11129,N_10374,N_9221);
nor U11130 (N_11130,N_10135,N_9680);
nand U11131 (N_11131,N_9983,N_10378);
or U11132 (N_11132,N_10123,N_9058);
xnor U11133 (N_11133,N_9334,N_10180);
nand U11134 (N_11134,N_9743,N_10297);
and U11135 (N_11135,N_9101,N_10492);
xnor U11136 (N_11136,N_9149,N_10253);
nor U11137 (N_11137,N_9384,N_9150);
or U11138 (N_11138,N_10388,N_10140);
and U11139 (N_11139,N_10306,N_9276);
and U11140 (N_11140,N_10041,N_9954);
nand U11141 (N_11141,N_9442,N_9749);
nand U11142 (N_11142,N_10057,N_9287);
xor U11143 (N_11143,N_10405,N_10441);
xnor U11144 (N_11144,N_9872,N_9002);
xor U11145 (N_11145,N_9328,N_9804);
nand U11146 (N_11146,N_10287,N_9812);
nand U11147 (N_11147,N_9831,N_9210);
nand U11148 (N_11148,N_9298,N_9415);
nand U11149 (N_11149,N_10318,N_9151);
nand U11150 (N_11150,N_9282,N_9135);
nand U11151 (N_11151,N_9909,N_10169);
xnor U11152 (N_11152,N_9206,N_9487);
nor U11153 (N_11153,N_9801,N_9822);
or U11154 (N_11154,N_9514,N_9946);
and U11155 (N_11155,N_9896,N_9319);
nand U11156 (N_11156,N_9472,N_9501);
nand U11157 (N_11157,N_9705,N_9289);
nand U11158 (N_11158,N_10189,N_9458);
or U11159 (N_11159,N_9784,N_10133);
nand U11160 (N_11160,N_10310,N_9885);
and U11161 (N_11161,N_10368,N_10261);
and U11162 (N_11162,N_9335,N_9779);
or U11163 (N_11163,N_9945,N_10221);
nor U11164 (N_11164,N_9939,N_10328);
nand U11165 (N_11165,N_9814,N_9301);
nor U11166 (N_11166,N_9740,N_9943);
nor U11167 (N_11167,N_10233,N_10071);
nand U11168 (N_11168,N_9322,N_10053);
xor U11169 (N_11169,N_9075,N_9071);
nand U11170 (N_11170,N_9755,N_9244);
nor U11171 (N_11171,N_9776,N_9129);
nor U11172 (N_11172,N_10363,N_9738);
xor U11173 (N_11173,N_9192,N_9066);
and U11174 (N_11174,N_9434,N_9456);
nand U11175 (N_11175,N_9196,N_10268);
nand U11176 (N_11176,N_10086,N_10482);
xnor U11177 (N_11177,N_9785,N_9898);
and U11178 (N_11178,N_9679,N_9866);
nor U11179 (N_11179,N_10078,N_10361);
xor U11180 (N_11180,N_9051,N_10252);
nor U11181 (N_11181,N_10389,N_10070);
or U11182 (N_11182,N_9826,N_9642);
nand U11183 (N_11183,N_9029,N_10033);
and U11184 (N_11184,N_9194,N_10217);
and U11185 (N_11185,N_9511,N_9007);
and U11186 (N_11186,N_9882,N_9591);
nand U11187 (N_11187,N_9424,N_10191);
nand U11188 (N_11188,N_9387,N_9519);
or U11189 (N_11189,N_9873,N_9722);
xor U11190 (N_11190,N_9266,N_10092);
or U11191 (N_11191,N_9348,N_9904);
or U11192 (N_11192,N_10149,N_9967);
nor U11193 (N_11193,N_10100,N_10257);
and U11194 (N_11194,N_10444,N_10319);
or U11195 (N_11195,N_9905,N_9982);
xor U11196 (N_11196,N_10012,N_10082);
or U11197 (N_11197,N_9247,N_9026);
or U11198 (N_11198,N_9887,N_9783);
xor U11199 (N_11199,N_10381,N_9169);
nand U11200 (N_11200,N_10145,N_9270);
nand U11201 (N_11201,N_9720,N_10112);
xnor U11202 (N_11202,N_10290,N_10157);
xnor U11203 (N_11203,N_9479,N_10011);
xor U11204 (N_11204,N_10143,N_9596);
xnor U11205 (N_11205,N_9759,N_10385);
and U11206 (N_11206,N_9178,N_9502);
or U11207 (N_11207,N_10211,N_10166);
and U11208 (N_11208,N_10142,N_9929);
or U11209 (N_11209,N_9021,N_10102);
xnor U11210 (N_11210,N_10412,N_9414);
and U11211 (N_11211,N_10490,N_9593);
and U11212 (N_11212,N_9119,N_10317);
xnor U11213 (N_11213,N_10474,N_9827);
xnor U11214 (N_11214,N_9854,N_9941);
and U11215 (N_11215,N_9575,N_9590);
nor U11216 (N_11216,N_10393,N_9771);
and U11217 (N_11217,N_9364,N_9894);
nand U11218 (N_11218,N_9094,N_9408);
nand U11219 (N_11219,N_9132,N_9052);
or U11220 (N_11220,N_9406,N_10348);
and U11221 (N_11221,N_9701,N_9199);
and U11222 (N_11222,N_9611,N_9984);
xor U11223 (N_11223,N_9614,N_9368);
xor U11224 (N_11224,N_9170,N_10491);
or U11225 (N_11225,N_10359,N_9975);
nand U11226 (N_11226,N_9125,N_9545);
or U11227 (N_11227,N_9303,N_10093);
nor U11228 (N_11228,N_9777,N_10276);
or U11229 (N_11229,N_9609,N_9305);
xor U11230 (N_11230,N_10174,N_9971);
or U11231 (N_11231,N_10463,N_9438);
nand U11232 (N_11232,N_9582,N_9900);
xor U11233 (N_11233,N_9451,N_10084);
nand U11234 (N_11234,N_9843,N_9260);
nand U11235 (N_11235,N_9417,N_9510);
nand U11236 (N_11236,N_10373,N_9767);
nand U11237 (N_11237,N_9688,N_10411);
nor U11238 (N_11238,N_9153,N_10023);
xnor U11239 (N_11239,N_9977,N_10245);
nor U11240 (N_11240,N_9765,N_9962);
xnor U11241 (N_11241,N_9703,N_10000);
and U11242 (N_11242,N_9659,N_9595);
nand U11243 (N_11243,N_10266,N_9128);
nand U11244 (N_11244,N_9164,N_10248);
or U11245 (N_11245,N_10327,N_10177);
and U11246 (N_11246,N_9057,N_10316);
nor U11247 (N_11247,N_9795,N_9721);
nor U11248 (N_11248,N_9253,N_9041);
nand U11249 (N_11249,N_9641,N_9653);
nand U11250 (N_11250,N_10187,N_10381);
and U11251 (N_11251,N_9292,N_10260);
nor U11252 (N_11252,N_9537,N_10479);
nor U11253 (N_11253,N_9449,N_10465);
nor U11254 (N_11254,N_10186,N_9977);
nor U11255 (N_11255,N_10005,N_9360);
or U11256 (N_11256,N_9015,N_9956);
xor U11257 (N_11257,N_9644,N_10387);
nor U11258 (N_11258,N_10017,N_9762);
or U11259 (N_11259,N_10111,N_10246);
nand U11260 (N_11260,N_10195,N_10448);
nand U11261 (N_11261,N_9438,N_10343);
nor U11262 (N_11262,N_9795,N_9382);
xnor U11263 (N_11263,N_10365,N_9814);
and U11264 (N_11264,N_10285,N_9876);
xor U11265 (N_11265,N_10334,N_10338);
nor U11266 (N_11266,N_9106,N_9740);
xor U11267 (N_11267,N_9511,N_9676);
nand U11268 (N_11268,N_9445,N_9984);
nor U11269 (N_11269,N_10089,N_9103);
and U11270 (N_11270,N_10168,N_9975);
and U11271 (N_11271,N_9728,N_9597);
xnor U11272 (N_11272,N_9154,N_10113);
xnor U11273 (N_11273,N_10285,N_9213);
nand U11274 (N_11274,N_9094,N_9564);
nand U11275 (N_11275,N_9164,N_10143);
xor U11276 (N_11276,N_9084,N_9890);
and U11277 (N_11277,N_9843,N_10114);
xnor U11278 (N_11278,N_9928,N_9941);
xor U11279 (N_11279,N_10475,N_9170);
and U11280 (N_11280,N_10206,N_10171);
xnor U11281 (N_11281,N_10140,N_10360);
or U11282 (N_11282,N_9534,N_9632);
nand U11283 (N_11283,N_9490,N_9140);
nor U11284 (N_11284,N_10443,N_9530);
xor U11285 (N_11285,N_10174,N_9890);
nand U11286 (N_11286,N_9967,N_9225);
nor U11287 (N_11287,N_10336,N_9913);
xnor U11288 (N_11288,N_9579,N_9805);
xor U11289 (N_11289,N_9453,N_10354);
xor U11290 (N_11290,N_10360,N_9647);
nand U11291 (N_11291,N_9476,N_9667);
and U11292 (N_11292,N_10462,N_9667);
xnor U11293 (N_11293,N_9745,N_9177);
nand U11294 (N_11294,N_9600,N_10281);
nor U11295 (N_11295,N_9716,N_10070);
and U11296 (N_11296,N_9022,N_9808);
xor U11297 (N_11297,N_9406,N_9982);
or U11298 (N_11298,N_10082,N_9233);
xor U11299 (N_11299,N_9696,N_9992);
nor U11300 (N_11300,N_10328,N_9886);
or U11301 (N_11301,N_10265,N_9097);
or U11302 (N_11302,N_10063,N_10375);
nor U11303 (N_11303,N_9011,N_9891);
nand U11304 (N_11304,N_9303,N_9492);
nor U11305 (N_11305,N_9611,N_9917);
and U11306 (N_11306,N_9785,N_10092);
or U11307 (N_11307,N_9445,N_9845);
xnor U11308 (N_11308,N_10346,N_9355);
and U11309 (N_11309,N_9387,N_10342);
or U11310 (N_11310,N_9338,N_9328);
nor U11311 (N_11311,N_9767,N_9673);
or U11312 (N_11312,N_9493,N_9874);
nand U11313 (N_11313,N_9009,N_10457);
xnor U11314 (N_11314,N_10112,N_9044);
and U11315 (N_11315,N_10125,N_10137);
nand U11316 (N_11316,N_9769,N_9033);
nor U11317 (N_11317,N_9389,N_9369);
nor U11318 (N_11318,N_10402,N_10199);
or U11319 (N_11319,N_10204,N_10393);
nand U11320 (N_11320,N_9332,N_9616);
nor U11321 (N_11321,N_10050,N_9905);
or U11322 (N_11322,N_9213,N_9724);
or U11323 (N_11323,N_9027,N_10137);
and U11324 (N_11324,N_9397,N_9078);
nor U11325 (N_11325,N_9764,N_10485);
nor U11326 (N_11326,N_10265,N_9208);
xnor U11327 (N_11327,N_9929,N_10318);
and U11328 (N_11328,N_9538,N_9574);
or U11329 (N_11329,N_9828,N_10032);
and U11330 (N_11330,N_9385,N_9257);
or U11331 (N_11331,N_10349,N_9738);
or U11332 (N_11332,N_9289,N_9652);
xor U11333 (N_11333,N_9022,N_9299);
and U11334 (N_11334,N_9288,N_10077);
xnor U11335 (N_11335,N_10440,N_9272);
nor U11336 (N_11336,N_9753,N_9763);
nand U11337 (N_11337,N_9884,N_10327);
and U11338 (N_11338,N_9312,N_10430);
and U11339 (N_11339,N_10126,N_9616);
and U11340 (N_11340,N_10183,N_10470);
or U11341 (N_11341,N_10001,N_9983);
xor U11342 (N_11342,N_10224,N_9846);
or U11343 (N_11343,N_9230,N_9260);
and U11344 (N_11344,N_9372,N_10273);
or U11345 (N_11345,N_9417,N_10100);
and U11346 (N_11346,N_9717,N_9782);
nor U11347 (N_11347,N_9579,N_9058);
xor U11348 (N_11348,N_10093,N_9948);
xnor U11349 (N_11349,N_9854,N_10304);
or U11350 (N_11350,N_10261,N_9122);
and U11351 (N_11351,N_9174,N_10273);
nor U11352 (N_11352,N_10447,N_10095);
and U11353 (N_11353,N_10112,N_9100);
and U11354 (N_11354,N_9625,N_9726);
or U11355 (N_11355,N_9809,N_9135);
xnor U11356 (N_11356,N_10405,N_9071);
or U11357 (N_11357,N_9165,N_9508);
or U11358 (N_11358,N_9602,N_9664);
xnor U11359 (N_11359,N_10188,N_9565);
nand U11360 (N_11360,N_9850,N_9525);
xnor U11361 (N_11361,N_9867,N_10268);
nor U11362 (N_11362,N_9565,N_10217);
and U11363 (N_11363,N_9660,N_9698);
nor U11364 (N_11364,N_10075,N_9483);
xnor U11365 (N_11365,N_10108,N_10105);
xor U11366 (N_11366,N_9616,N_9697);
xor U11367 (N_11367,N_10127,N_9180);
nand U11368 (N_11368,N_9132,N_9116);
nand U11369 (N_11369,N_10264,N_10060);
or U11370 (N_11370,N_9849,N_9857);
nand U11371 (N_11371,N_9689,N_9889);
nor U11372 (N_11372,N_9404,N_9688);
and U11373 (N_11373,N_9224,N_9877);
xnor U11374 (N_11374,N_10004,N_10080);
nor U11375 (N_11375,N_9756,N_10424);
nand U11376 (N_11376,N_9031,N_9411);
xor U11377 (N_11377,N_10018,N_10379);
or U11378 (N_11378,N_9213,N_9560);
or U11379 (N_11379,N_10303,N_9823);
xor U11380 (N_11380,N_9260,N_9922);
or U11381 (N_11381,N_10481,N_9297);
and U11382 (N_11382,N_9670,N_10291);
nor U11383 (N_11383,N_9166,N_9948);
or U11384 (N_11384,N_10442,N_10145);
and U11385 (N_11385,N_10084,N_9370);
xnor U11386 (N_11386,N_10353,N_10220);
and U11387 (N_11387,N_10401,N_9938);
and U11388 (N_11388,N_9204,N_10399);
xnor U11389 (N_11389,N_9096,N_9264);
and U11390 (N_11390,N_9877,N_10109);
or U11391 (N_11391,N_9312,N_9880);
nor U11392 (N_11392,N_10291,N_9309);
or U11393 (N_11393,N_9554,N_9009);
and U11394 (N_11394,N_10194,N_9662);
or U11395 (N_11395,N_9570,N_9574);
and U11396 (N_11396,N_9398,N_9409);
and U11397 (N_11397,N_9968,N_10289);
nor U11398 (N_11398,N_9319,N_9042);
or U11399 (N_11399,N_9184,N_10092);
nor U11400 (N_11400,N_9721,N_10048);
xnor U11401 (N_11401,N_9469,N_9834);
xor U11402 (N_11402,N_10400,N_10386);
or U11403 (N_11403,N_10286,N_9893);
and U11404 (N_11404,N_9513,N_9520);
nand U11405 (N_11405,N_9156,N_9587);
and U11406 (N_11406,N_10114,N_10307);
or U11407 (N_11407,N_10239,N_9638);
xor U11408 (N_11408,N_9622,N_10296);
and U11409 (N_11409,N_10199,N_10119);
nor U11410 (N_11410,N_9670,N_9928);
nand U11411 (N_11411,N_9492,N_9263);
and U11412 (N_11412,N_9807,N_9834);
and U11413 (N_11413,N_9119,N_9093);
or U11414 (N_11414,N_9796,N_9061);
and U11415 (N_11415,N_10057,N_9433);
xnor U11416 (N_11416,N_10027,N_10411);
and U11417 (N_11417,N_9923,N_10021);
and U11418 (N_11418,N_9089,N_9572);
xor U11419 (N_11419,N_10493,N_9194);
and U11420 (N_11420,N_9527,N_9482);
nor U11421 (N_11421,N_9766,N_10436);
nor U11422 (N_11422,N_10021,N_9755);
or U11423 (N_11423,N_9334,N_9843);
nand U11424 (N_11424,N_9358,N_9170);
or U11425 (N_11425,N_10154,N_10184);
xor U11426 (N_11426,N_9533,N_9933);
nor U11427 (N_11427,N_9806,N_10082);
nand U11428 (N_11428,N_9521,N_9574);
nor U11429 (N_11429,N_10437,N_9578);
nand U11430 (N_11430,N_10392,N_9887);
or U11431 (N_11431,N_9546,N_10006);
nand U11432 (N_11432,N_9712,N_10008);
nand U11433 (N_11433,N_9932,N_9444);
nor U11434 (N_11434,N_9193,N_9078);
and U11435 (N_11435,N_9803,N_10139);
xor U11436 (N_11436,N_10029,N_9890);
and U11437 (N_11437,N_9365,N_9892);
nor U11438 (N_11438,N_9478,N_9157);
nor U11439 (N_11439,N_9223,N_9540);
nand U11440 (N_11440,N_9187,N_9471);
or U11441 (N_11441,N_9999,N_9681);
nand U11442 (N_11442,N_10352,N_9543);
or U11443 (N_11443,N_9513,N_9276);
and U11444 (N_11444,N_9120,N_9573);
or U11445 (N_11445,N_9485,N_10229);
nand U11446 (N_11446,N_9320,N_9493);
xnor U11447 (N_11447,N_9271,N_9211);
nand U11448 (N_11448,N_9880,N_10086);
nor U11449 (N_11449,N_9312,N_9268);
nand U11450 (N_11450,N_9002,N_9407);
nor U11451 (N_11451,N_10423,N_9684);
and U11452 (N_11452,N_9293,N_9553);
xnor U11453 (N_11453,N_10272,N_9908);
xor U11454 (N_11454,N_9388,N_10274);
nand U11455 (N_11455,N_9750,N_10200);
and U11456 (N_11456,N_9535,N_9334);
xor U11457 (N_11457,N_9092,N_10485);
or U11458 (N_11458,N_9014,N_9600);
xor U11459 (N_11459,N_9822,N_9569);
or U11460 (N_11460,N_10036,N_10311);
and U11461 (N_11461,N_10098,N_9601);
nand U11462 (N_11462,N_9005,N_10120);
and U11463 (N_11463,N_9556,N_9996);
nor U11464 (N_11464,N_10198,N_9155);
xnor U11465 (N_11465,N_9919,N_9129);
xnor U11466 (N_11466,N_9521,N_10420);
and U11467 (N_11467,N_9543,N_9683);
xor U11468 (N_11468,N_9525,N_9714);
xor U11469 (N_11469,N_10349,N_10190);
and U11470 (N_11470,N_9141,N_10128);
nor U11471 (N_11471,N_10353,N_9087);
nand U11472 (N_11472,N_9886,N_10056);
or U11473 (N_11473,N_9113,N_10397);
or U11474 (N_11474,N_9508,N_9640);
nand U11475 (N_11475,N_9843,N_10070);
or U11476 (N_11476,N_10340,N_9022);
nor U11477 (N_11477,N_9011,N_9096);
nor U11478 (N_11478,N_9629,N_10193);
xnor U11479 (N_11479,N_10384,N_9834);
nand U11480 (N_11480,N_10294,N_9971);
nor U11481 (N_11481,N_9541,N_9117);
xor U11482 (N_11482,N_9392,N_10419);
and U11483 (N_11483,N_9148,N_9584);
and U11484 (N_11484,N_10344,N_9948);
nand U11485 (N_11485,N_9782,N_9530);
nor U11486 (N_11486,N_9032,N_9313);
nor U11487 (N_11487,N_9056,N_9447);
nor U11488 (N_11488,N_10238,N_9352);
nand U11489 (N_11489,N_10382,N_9583);
nor U11490 (N_11490,N_9967,N_9580);
or U11491 (N_11491,N_9182,N_10235);
or U11492 (N_11492,N_9298,N_9583);
nor U11493 (N_11493,N_9782,N_10189);
xnor U11494 (N_11494,N_10420,N_10231);
or U11495 (N_11495,N_10339,N_10437);
and U11496 (N_11496,N_9954,N_9105);
xnor U11497 (N_11497,N_9103,N_9389);
xor U11498 (N_11498,N_10140,N_9443);
or U11499 (N_11499,N_10128,N_10215);
nor U11500 (N_11500,N_9679,N_9250);
nand U11501 (N_11501,N_9102,N_9563);
xnor U11502 (N_11502,N_9252,N_10110);
xor U11503 (N_11503,N_9081,N_9787);
nand U11504 (N_11504,N_9246,N_10312);
nand U11505 (N_11505,N_10121,N_9733);
and U11506 (N_11506,N_9224,N_9696);
xor U11507 (N_11507,N_10477,N_9387);
xnor U11508 (N_11508,N_9310,N_9777);
nor U11509 (N_11509,N_9168,N_9665);
xnor U11510 (N_11510,N_10488,N_9316);
nor U11511 (N_11511,N_10057,N_9370);
nor U11512 (N_11512,N_10219,N_10310);
or U11513 (N_11513,N_9192,N_9323);
xnor U11514 (N_11514,N_10204,N_9618);
xnor U11515 (N_11515,N_9788,N_10410);
nand U11516 (N_11516,N_9845,N_10194);
and U11517 (N_11517,N_10470,N_9151);
nor U11518 (N_11518,N_9096,N_10046);
nand U11519 (N_11519,N_10072,N_10230);
nor U11520 (N_11520,N_10491,N_9703);
nor U11521 (N_11521,N_9690,N_10070);
xor U11522 (N_11522,N_10009,N_10297);
or U11523 (N_11523,N_9316,N_9952);
nor U11524 (N_11524,N_9336,N_10142);
or U11525 (N_11525,N_9922,N_10375);
nor U11526 (N_11526,N_10365,N_9519);
nand U11527 (N_11527,N_10251,N_9384);
xor U11528 (N_11528,N_9919,N_9909);
or U11529 (N_11529,N_9528,N_10341);
nand U11530 (N_11530,N_9343,N_10328);
and U11531 (N_11531,N_10225,N_9376);
or U11532 (N_11532,N_9032,N_10348);
xor U11533 (N_11533,N_10047,N_9619);
xnor U11534 (N_11534,N_9365,N_9430);
nand U11535 (N_11535,N_10217,N_9937);
and U11536 (N_11536,N_10004,N_9061);
nor U11537 (N_11537,N_9701,N_9207);
and U11538 (N_11538,N_9716,N_10307);
nand U11539 (N_11539,N_10459,N_9032);
and U11540 (N_11540,N_9018,N_9271);
nand U11541 (N_11541,N_9101,N_9434);
or U11542 (N_11542,N_9332,N_9435);
nand U11543 (N_11543,N_9029,N_9093);
nand U11544 (N_11544,N_9787,N_9403);
or U11545 (N_11545,N_9723,N_10472);
xnor U11546 (N_11546,N_10343,N_10047);
xnor U11547 (N_11547,N_9483,N_10119);
nand U11548 (N_11548,N_9460,N_10181);
nand U11549 (N_11549,N_9762,N_9923);
xnor U11550 (N_11550,N_9293,N_9058);
xnor U11551 (N_11551,N_9132,N_9509);
xor U11552 (N_11552,N_10479,N_9378);
xnor U11553 (N_11553,N_9742,N_9147);
nor U11554 (N_11554,N_9190,N_9298);
and U11555 (N_11555,N_9627,N_9065);
nand U11556 (N_11556,N_9339,N_10218);
or U11557 (N_11557,N_9895,N_10394);
xor U11558 (N_11558,N_9708,N_10484);
xnor U11559 (N_11559,N_9776,N_10337);
nor U11560 (N_11560,N_10363,N_9518);
nand U11561 (N_11561,N_9384,N_9746);
or U11562 (N_11562,N_10482,N_9954);
or U11563 (N_11563,N_10398,N_9438);
or U11564 (N_11564,N_10211,N_9992);
nand U11565 (N_11565,N_9563,N_9307);
or U11566 (N_11566,N_9972,N_9850);
and U11567 (N_11567,N_10041,N_9339);
xor U11568 (N_11568,N_10160,N_10029);
xnor U11569 (N_11569,N_9337,N_10256);
or U11570 (N_11570,N_9595,N_9680);
xnor U11571 (N_11571,N_9518,N_9369);
or U11572 (N_11572,N_9583,N_9109);
nand U11573 (N_11573,N_9859,N_10406);
xor U11574 (N_11574,N_9869,N_9192);
or U11575 (N_11575,N_9841,N_9943);
or U11576 (N_11576,N_9944,N_10465);
nor U11577 (N_11577,N_9764,N_10159);
nor U11578 (N_11578,N_10130,N_9007);
xor U11579 (N_11579,N_9453,N_10439);
xor U11580 (N_11580,N_10217,N_10434);
nand U11581 (N_11581,N_10400,N_9814);
xor U11582 (N_11582,N_9683,N_9112);
and U11583 (N_11583,N_9131,N_10341);
xor U11584 (N_11584,N_9547,N_9144);
and U11585 (N_11585,N_10058,N_10342);
and U11586 (N_11586,N_10387,N_9789);
nand U11587 (N_11587,N_9906,N_9072);
or U11588 (N_11588,N_10459,N_9890);
and U11589 (N_11589,N_9854,N_10465);
nand U11590 (N_11590,N_10360,N_9766);
or U11591 (N_11591,N_10144,N_9368);
nand U11592 (N_11592,N_9441,N_10204);
xnor U11593 (N_11593,N_9831,N_10282);
nor U11594 (N_11594,N_10079,N_9967);
nor U11595 (N_11595,N_9363,N_10217);
or U11596 (N_11596,N_9202,N_9632);
nor U11597 (N_11597,N_10061,N_10327);
or U11598 (N_11598,N_9661,N_9796);
nor U11599 (N_11599,N_10395,N_9515);
nor U11600 (N_11600,N_9775,N_9304);
and U11601 (N_11601,N_9518,N_10282);
xor U11602 (N_11602,N_10062,N_9519);
nor U11603 (N_11603,N_9909,N_10016);
xnor U11604 (N_11604,N_9025,N_9030);
and U11605 (N_11605,N_10252,N_10439);
nor U11606 (N_11606,N_10213,N_9515);
nand U11607 (N_11607,N_10104,N_9313);
xnor U11608 (N_11608,N_9098,N_9008);
and U11609 (N_11609,N_9901,N_9641);
xor U11610 (N_11610,N_9201,N_10152);
nand U11611 (N_11611,N_10106,N_10013);
and U11612 (N_11612,N_9934,N_10296);
xnor U11613 (N_11613,N_10358,N_10156);
and U11614 (N_11614,N_9090,N_10436);
nor U11615 (N_11615,N_10391,N_10291);
nand U11616 (N_11616,N_9321,N_9726);
nor U11617 (N_11617,N_10265,N_9079);
nor U11618 (N_11618,N_9742,N_9827);
or U11619 (N_11619,N_10245,N_9286);
xnor U11620 (N_11620,N_10347,N_9998);
xnor U11621 (N_11621,N_9006,N_10140);
xor U11622 (N_11622,N_9249,N_9411);
or U11623 (N_11623,N_9232,N_9160);
xor U11624 (N_11624,N_10331,N_9763);
xnor U11625 (N_11625,N_9466,N_10343);
xnor U11626 (N_11626,N_10036,N_9683);
xor U11627 (N_11627,N_9114,N_10024);
or U11628 (N_11628,N_9876,N_9095);
nor U11629 (N_11629,N_10019,N_10410);
xnor U11630 (N_11630,N_10214,N_10257);
and U11631 (N_11631,N_9991,N_9278);
or U11632 (N_11632,N_9270,N_9806);
nor U11633 (N_11633,N_9124,N_9458);
nand U11634 (N_11634,N_9776,N_10002);
nor U11635 (N_11635,N_9756,N_10004);
nor U11636 (N_11636,N_10219,N_9728);
xnor U11637 (N_11637,N_9203,N_9128);
xnor U11638 (N_11638,N_9607,N_9318);
and U11639 (N_11639,N_9653,N_9960);
or U11640 (N_11640,N_9854,N_9202);
nor U11641 (N_11641,N_9360,N_9618);
or U11642 (N_11642,N_10219,N_9596);
and U11643 (N_11643,N_9837,N_9811);
nand U11644 (N_11644,N_10472,N_9358);
and U11645 (N_11645,N_10433,N_9537);
nor U11646 (N_11646,N_9249,N_10087);
nand U11647 (N_11647,N_9328,N_9839);
and U11648 (N_11648,N_9613,N_10353);
xnor U11649 (N_11649,N_9858,N_9409);
or U11650 (N_11650,N_9352,N_9735);
nor U11651 (N_11651,N_10113,N_9641);
nor U11652 (N_11652,N_9247,N_9479);
and U11653 (N_11653,N_9162,N_10119);
or U11654 (N_11654,N_9458,N_9371);
and U11655 (N_11655,N_9732,N_9500);
xor U11656 (N_11656,N_9020,N_9113);
and U11657 (N_11657,N_9761,N_9370);
or U11658 (N_11658,N_10136,N_10046);
and U11659 (N_11659,N_10210,N_9358);
or U11660 (N_11660,N_9481,N_9415);
and U11661 (N_11661,N_10252,N_9951);
and U11662 (N_11662,N_10048,N_9802);
xor U11663 (N_11663,N_10216,N_9021);
nand U11664 (N_11664,N_9949,N_9716);
and U11665 (N_11665,N_9251,N_9601);
or U11666 (N_11666,N_9166,N_10197);
nand U11667 (N_11667,N_10090,N_9970);
or U11668 (N_11668,N_10378,N_9528);
or U11669 (N_11669,N_10167,N_9586);
and U11670 (N_11670,N_9930,N_9727);
nand U11671 (N_11671,N_10212,N_10487);
nand U11672 (N_11672,N_9233,N_9208);
xor U11673 (N_11673,N_9877,N_10215);
nand U11674 (N_11674,N_10117,N_9496);
and U11675 (N_11675,N_9846,N_10106);
xor U11676 (N_11676,N_9267,N_9503);
and U11677 (N_11677,N_10297,N_9560);
nor U11678 (N_11678,N_10271,N_9931);
and U11679 (N_11679,N_10212,N_9545);
and U11680 (N_11680,N_10433,N_9128);
and U11681 (N_11681,N_9269,N_9622);
or U11682 (N_11682,N_10112,N_9281);
xnor U11683 (N_11683,N_9860,N_9153);
xor U11684 (N_11684,N_9136,N_9300);
nand U11685 (N_11685,N_9440,N_10337);
or U11686 (N_11686,N_9025,N_9389);
nand U11687 (N_11687,N_9504,N_9097);
and U11688 (N_11688,N_9171,N_9660);
nand U11689 (N_11689,N_9816,N_10255);
nor U11690 (N_11690,N_10163,N_9124);
and U11691 (N_11691,N_10297,N_9138);
xnor U11692 (N_11692,N_9038,N_9497);
xor U11693 (N_11693,N_10495,N_9885);
xnor U11694 (N_11694,N_9568,N_9003);
xor U11695 (N_11695,N_9543,N_9117);
nand U11696 (N_11696,N_10372,N_9435);
xnor U11697 (N_11697,N_9977,N_9641);
xor U11698 (N_11698,N_9054,N_10288);
xnor U11699 (N_11699,N_10430,N_10374);
and U11700 (N_11700,N_10298,N_9452);
xor U11701 (N_11701,N_10366,N_9583);
and U11702 (N_11702,N_9554,N_10099);
and U11703 (N_11703,N_9811,N_9676);
nand U11704 (N_11704,N_10025,N_10201);
and U11705 (N_11705,N_10054,N_10334);
nor U11706 (N_11706,N_10305,N_9496);
nand U11707 (N_11707,N_10159,N_10443);
nor U11708 (N_11708,N_9721,N_10293);
or U11709 (N_11709,N_10185,N_9301);
and U11710 (N_11710,N_9172,N_9105);
nand U11711 (N_11711,N_9871,N_10471);
xor U11712 (N_11712,N_9248,N_9345);
xnor U11713 (N_11713,N_10434,N_9823);
nand U11714 (N_11714,N_9335,N_9359);
or U11715 (N_11715,N_9235,N_10379);
nor U11716 (N_11716,N_10228,N_10298);
and U11717 (N_11717,N_9024,N_9636);
xnor U11718 (N_11718,N_9410,N_9375);
or U11719 (N_11719,N_10330,N_9102);
or U11720 (N_11720,N_9430,N_9651);
nor U11721 (N_11721,N_9199,N_9404);
xnor U11722 (N_11722,N_9847,N_10346);
nor U11723 (N_11723,N_9971,N_9519);
xor U11724 (N_11724,N_9440,N_9142);
nor U11725 (N_11725,N_9180,N_9459);
xor U11726 (N_11726,N_9126,N_9785);
nand U11727 (N_11727,N_9555,N_9209);
nor U11728 (N_11728,N_9762,N_10418);
nor U11729 (N_11729,N_9293,N_10317);
xor U11730 (N_11730,N_9701,N_9640);
nor U11731 (N_11731,N_9243,N_9851);
nand U11732 (N_11732,N_10199,N_9623);
nor U11733 (N_11733,N_10410,N_10118);
and U11734 (N_11734,N_10464,N_9844);
nand U11735 (N_11735,N_10088,N_9513);
and U11736 (N_11736,N_10443,N_9466);
and U11737 (N_11737,N_10206,N_9191);
or U11738 (N_11738,N_10282,N_9769);
and U11739 (N_11739,N_10065,N_9579);
nand U11740 (N_11740,N_10327,N_9937);
xnor U11741 (N_11741,N_9518,N_9835);
or U11742 (N_11742,N_9069,N_10285);
nand U11743 (N_11743,N_9605,N_9076);
xnor U11744 (N_11744,N_9643,N_10486);
and U11745 (N_11745,N_9719,N_9462);
or U11746 (N_11746,N_9818,N_9659);
nand U11747 (N_11747,N_9024,N_9772);
xor U11748 (N_11748,N_10251,N_10496);
xnor U11749 (N_11749,N_10227,N_9496);
nand U11750 (N_11750,N_10430,N_10339);
and U11751 (N_11751,N_9812,N_9109);
nor U11752 (N_11752,N_9863,N_9389);
nand U11753 (N_11753,N_10492,N_9886);
xor U11754 (N_11754,N_9046,N_9697);
nor U11755 (N_11755,N_10061,N_9191);
or U11756 (N_11756,N_10480,N_10447);
and U11757 (N_11757,N_9044,N_9751);
nand U11758 (N_11758,N_9979,N_9447);
nand U11759 (N_11759,N_10339,N_10377);
or U11760 (N_11760,N_9875,N_9184);
and U11761 (N_11761,N_9433,N_10146);
or U11762 (N_11762,N_9662,N_10085);
nand U11763 (N_11763,N_10333,N_9929);
and U11764 (N_11764,N_9190,N_9671);
xor U11765 (N_11765,N_9363,N_9207);
nor U11766 (N_11766,N_9801,N_9133);
nand U11767 (N_11767,N_9059,N_9946);
nand U11768 (N_11768,N_9027,N_9931);
or U11769 (N_11769,N_9705,N_9806);
nand U11770 (N_11770,N_9875,N_9456);
nor U11771 (N_11771,N_9493,N_10416);
and U11772 (N_11772,N_9826,N_9870);
nand U11773 (N_11773,N_9421,N_9851);
and U11774 (N_11774,N_9730,N_10243);
and U11775 (N_11775,N_9957,N_9035);
nor U11776 (N_11776,N_10192,N_9435);
nand U11777 (N_11777,N_10195,N_9170);
xor U11778 (N_11778,N_9475,N_9446);
xnor U11779 (N_11779,N_10193,N_10049);
and U11780 (N_11780,N_9583,N_9851);
and U11781 (N_11781,N_9520,N_10208);
nand U11782 (N_11782,N_9987,N_10454);
nand U11783 (N_11783,N_9106,N_9274);
and U11784 (N_11784,N_9089,N_10273);
or U11785 (N_11785,N_9164,N_9301);
or U11786 (N_11786,N_9033,N_10011);
xor U11787 (N_11787,N_10088,N_10337);
or U11788 (N_11788,N_9059,N_9691);
and U11789 (N_11789,N_9841,N_9883);
nor U11790 (N_11790,N_9976,N_10108);
nor U11791 (N_11791,N_10464,N_10168);
or U11792 (N_11792,N_9706,N_9582);
nand U11793 (N_11793,N_9927,N_9008);
and U11794 (N_11794,N_9106,N_9825);
nor U11795 (N_11795,N_9899,N_10298);
or U11796 (N_11796,N_9260,N_9302);
xor U11797 (N_11797,N_9498,N_10114);
and U11798 (N_11798,N_9932,N_9767);
or U11799 (N_11799,N_9623,N_9260);
nor U11800 (N_11800,N_9327,N_10185);
xnor U11801 (N_11801,N_10423,N_10209);
nand U11802 (N_11802,N_9495,N_9969);
nand U11803 (N_11803,N_9318,N_9804);
nand U11804 (N_11804,N_10267,N_9885);
xor U11805 (N_11805,N_10205,N_10223);
or U11806 (N_11806,N_10042,N_10072);
nand U11807 (N_11807,N_9608,N_10328);
or U11808 (N_11808,N_10191,N_9419);
xor U11809 (N_11809,N_9110,N_9601);
xnor U11810 (N_11810,N_10275,N_10400);
xnor U11811 (N_11811,N_10032,N_9205);
or U11812 (N_11812,N_10092,N_9151);
nor U11813 (N_11813,N_10440,N_9157);
xnor U11814 (N_11814,N_9797,N_9677);
nand U11815 (N_11815,N_10167,N_9301);
and U11816 (N_11816,N_9277,N_10490);
or U11817 (N_11817,N_10102,N_9274);
or U11818 (N_11818,N_9533,N_10307);
and U11819 (N_11819,N_9145,N_9912);
nor U11820 (N_11820,N_9127,N_9706);
xor U11821 (N_11821,N_9163,N_9400);
or U11822 (N_11822,N_10490,N_9562);
nor U11823 (N_11823,N_9483,N_10216);
and U11824 (N_11824,N_9223,N_9399);
and U11825 (N_11825,N_9754,N_9452);
nand U11826 (N_11826,N_9130,N_9506);
nand U11827 (N_11827,N_9963,N_10113);
nand U11828 (N_11828,N_9416,N_9257);
and U11829 (N_11829,N_9166,N_10064);
xnor U11830 (N_11830,N_9298,N_9147);
nor U11831 (N_11831,N_10311,N_9206);
or U11832 (N_11832,N_9787,N_9922);
or U11833 (N_11833,N_10481,N_10131);
nor U11834 (N_11834,N_9442,N_9087);
xor U11835 (N_11835,N_9886,N_10121);
xor U11836 (N_11836,N_9893,N_10275);
nor U11837 (N_11837,N_10282,N_9843);
nand U11838 (N_11838,N_10048,N_10141);
and U11839 (N_11839,N_9326,N_10294);
xnor U11840 (N_11840,N_10317,N_9875);
xor U11841 (N_11841,N_9962,N_9423);
or U11842 (N_11842,N_9881,N_9371);
nor U11843 (N_11843,N_9009,N_9283);
nand U11844 (N_11844,N_10379,N_10120);
nand U11845 (N_11845,N_9338,N_9500);
or U11846 (N_11846,N_10180,N_9174);
and U11847 (N_11847,N_9761,N_10469);
xor U11848 (N_11848,N_9017,N_9353);
nand U11849 (N_11849,N_10461,N_10419);
xor U11850 (N_11850,N_9437,N_10389);
xor U11851 (N_11851,N_10067,N_9744);
nor U11852 (N_11852,N_9432,N_9272);
xor U11853 (N_11853,N_10238,N_9126);
or U11854 (N_11854,N_9393,N_10380);
nand U11855 (N_11855,N_9886,N_9242);
xor U11856 (N_11856,N_10360,N_10045);
and U11857 (N_11857,N_10466,N_10487);
xor U11858 (N_11858,N_9211,N_9537);
or U11859 (N_11859,N_9804,N_9529);
nand U11860 (N_11860,N_9664,N_9451);
and U11861 (N_11861,N_9273,N_9834);
and U11862 (N_11862,N_10314,N_10172);
nand U11863 (N_11863,N_9062,N_9855);
nor U11864 (N_11864,N_9123,N_10376);
or U11865 (N_11865,N_9780,N_10164);
nor U11866 (N_11866,N_10023,N_9794);
nor U11867 (N_11867,N_10437,N_9990);
and U11868 (N_11868,N_9018,N_9468);
nand U11869 (N_11869,N_9419,N_10202);
and U11870 (N_11870,N_9063,N_9108);
nor U11871 (N_11871,N_9718,N_9320);
nor U11872 (N_11872,N_9810,N_10153);
nand U11873 (N_11873,N_10097,N_9667);
xnor U11874 (N_11874,N_9752,N_9492);
and U11875 (N_11875,N_10145,N_10290);
or U11876 (N_11876,N_9235,N_9962);
nor U11877 (N_11877,N_9239,N_10055);
and U11878 (N_11878,N_9093,N_9237);
nor U11879 (N_11879,N_9494,N_9352);
xor U11880 (N_11880,N_9415,N_9965);
or U11881 (N_11881,N_9408,N_9881);
and U11882 (N_11882,N_9735,N_9676);
nand U11883 (N_11883,N_10454,N_9160);
nor U11884 (N_11884,N_9011,N_9030);
nor U11885 (N_11885,N_9110,N_9668);
nor U11886 (N_11886,N_9552,N_10011);
or U11887 (N_11887,N_10005,N_9411);
or U11888 (N_11888,N_10449,N_10284);
and U11889 (N_11889,N_9364,N_9040);
or U11890 (N_11890,N_9365,N_9574);
nor U11891 (N_11891,N_10262,N_9062);
or U11892 (N_11892,N_10157,N_10244);
and U11893 (N_11893,N_9174,N_10100);
xor U11894 (N_11894,N_9749,N_10471);
xor U11895 (N_11895,N_9157,N_9951);
nor U11896 (N_11896,N_9421,N_9637);
or U11897 (N_11897,N_9067,N_9121);
xor U11898 (N_11898,N_9510,N_9522);
and U11899 (N_11899,N_9405,N_9548);
nand U11900 (N_11900,N_9152,N_9189);
or U11901 (N_11901,N_9236,N_10306);
nand U11902 (N_11902,N_9040,N_9915);
and U11903 (N_11903,N_10162,N_9989);
or U11904 (N_11904,N_9660,N_10292);
nor U11905 (N_11905,N_10273,N_9969);
and U11906 (N_11906,N_9247,N_9345);
nor U11907 (N_11907,N_10267,N_10054);
and U11908 (N_11908,N_10486,N_10436);
or U11909 (N_11909,N_10203,N_9879);
xnor U11910 (N_11910,N_9004,N_9828);
nand U11911 (N_11911,N_9722,N_9610);
nand U11912 (N_11912,N_9063,N_10386);
nor U11913 (N_11913,N_9992,N_9873);
or U11914 (N_11914,N_10498,N_9076);
nand U11915 (N_11915,N_9860,N_9275);
nand U11916 (N_11916,N_10186,N_10205);
or U11917 (N_11917,N_9376,N_10241);
xor U11918 (N_11918,N_9010,N_9856);
nand U11919 (N_11919,N_9833,N_10023);
nor U11920 (N_11920,N_9924,N_9488);
nand U11921 (N_11921,N_9163,N_9152);
and U11922 (N_11922,N_9509,N_10180);
xor U11923 (N_11923,N_10382,N_9762);
nor U11924 (N_11924,N_9756,N_10358);
xor U11925 (N_11925,N_9044,N_9195);
and U11926 (N_11926,N_9475,N_9507);
nor U11927 (N_11927,N_9520,N_9665);
xnor U11928 (N_11928,N_9923,N_10218);
or U11929 (N_11929,N_9453,N_9217);
or U11930 (N_11930,N_9311,N_9601);
and U11931 (N_11931,N_9475,N_9255);
xor U11932 (N_11932,N_10426,N_9588);
xor U11933 (N_11933,N_9985,N_9005);
nand U11934 (N_11934,N_10466,N_9693);
nand U11935 (N_11935,N_9452,N_9807);
or U11936 (N_11936,N_10182,N_10388);
nand U11937 (N_11937,N_9902,N_9686);
and U11938 (N_11938,N_9650,N_9156);
nand U11939 (N_11939,N_9671,N_10046);
nor U11940 (N_11940,N_9639,N_9312);
xor U11941 (N_11941,N_9187,N_10428);
or U11942 (N_11942,N_9326,N_9955);
xor U11943 (N_11943,N_10302,N_10257);
nor U11944 (N_11944,N_9015,N_9794);
nor U11945 (N_11945,N_9065,N_9926);
nor U11946 (N_11946,N_10078,N_9713);
nand U11947 (N_11947,N_9534,N_9727);
and U11948 (N_11948,N_10213,N_10388);
or U11949 (N_11949,N_10033,N_10225);
nand U11950 (N_11950,N_10388,N_10323);
xor U11951 (N_11951,N_10066,N_9261);
nor U11952 (N_11952,N_10276,N_9192);
or U11953 (N_11953,N_9630,N_9584);
and U11954 (N_11954,N_10272,N_10032);
and U11955 (N_11955,N_10361,N_9353);
or U11956 (N_11956,N_10189,N_9078);
or U11957 (N_11957,N_10434,N_10196);
xor U11958 (N_11958,N_9055,N_9866);
xnor U11959 (N_11959,N_10494,N_9403);
or U11960 (N_11960,N_9503,N_9790);
nand U11961 (N_11961,N_10224,N_10296);
or U11962 (N_11962,N_9060,N_10183);
or U11963 (N_11963,N_9933,N_9434);
nor U11964 (N_11964,N_10026,N_9071);
and U11965 (N_11965,N_10158,N_9758);
and U11966 (N_11966,N_9243,N_9803);
and U11967 (N_11967,N_10480,N_10392);
and U11968 (N_11968,N_10402,N_10335);
or U11969 (N_11969,N_9041,N_10458);
xor U11970 (N_11970,N_9532,N_10062);
nand U11971 (N_11971,N_10136,N_9208);
xor U11972 (N_11972,N_9015,N_9592);
nand U11973 (N_11973,N_9546,N_9641);
or U11974 (N_11974,N_9378,N_10051);
and U11975 (N_11975,N_9677,N_9980);
and U11976 (N_11976,N_9567,N_9635);
nor U11977 (N_11977,N_9994,N_9502);
nor U11978 (N_11978,N_9907,N_9545);
nand U11979 (N_11979,N_10302,N_9485);
nand U11980 (N_11980,N_9251,N_9077);
or U11981 (N_11981,N_9080,N_9301);
nand U11982 (N_11982,N_9347,N_9672);
xor U11983 (N_11983,N_9340,N_10358);
nor U11984 (N_11984,N_9846,N_9106);
nand U11985 (N_11985,N_9985,N_9315);
and U11986 (N_11986,N_9966,N_10466);
or U11987 (N_11987,N_9961,N_9863);
xnor U11988 (N_11988,N_9453,N_9264);
nand U11989 (N_11989,N_9251,N_9612);
nand U11990 (N_11990,N_10295,N_9938);
nand U11991 (N_11991,N_9833,N_9760);
and U11992 (N_11992,N_9893,N_9602);
nor U11993 (N_11993,N_10279,N_9222);
nor U11994 (N_11994,N_9291,N_9139);
xor U11995 (N_11995,N_9288,N_9404);
nor U11996 (N_11996,N_10211,N_9442);
or U11997 (N_11997,N_10178,N_10372);
and U11998 (N_11998,N_10434,N_9670);
nor U11999 (N_11999,N_9446,N_10036);
nand U12000 (N_12000,N_10865,N_11287);
and U12001 (N_12001,N_11255,N_10885);
or U12002 (N_12002,N_11436,N_10712);
and U12003 (N_12003,N_10754,N_10632);
xor U12004 (N_12004,N_10923,N_10912);
and U12005 (N_12005,N_10718,N_11268);
nor U12006 (N_12006,N_10975,N_11306);
nand U12007 (N_12007,N_11189,N_11216);
and U12008 (N_12008,N_10594,N_11199);
nor U12009 (N_12009,N_10612,N_11186);
nand U12010 (N_12010,N_10661,N_10650);
or U12011 (N_12011,N_11825,N_11024);
or U12012 (N_12012,N_10515,N_11442);
and U12013 (N_12013,N_10777,N_11129);
and U12014 (N_12014,N_11307,N_11979);
nor U12015 (N_12015,N_10895,N_11217);
and U12016 (N_12016,N_10868,N_11848);
nand U12017 (N_12017,N_11691,N_11385);
nand U12018 (N_12018,N_11430,N_10817);
xor U12019 (N_12019,N_10607,N_11159);
or U12020 (N_12020,N_11044,N_11944);
xor U12021 (N_12021,N_11459,N_10557);
nor U12022 (N_12022,N_11135,N_11651);
nor U12023 (N_12023,N_11987,N_10966);
and U12024 (N_12024,N_11886,N_11816);
and U12025 (N_12025,N_10507,N_11184);
xnor U12026 (N_12026,N_11820,N_11210);
nand U12027 (N_12027,N_10506,N_10510);
and U12028 (N_12028,N_11512,N_10910);
xnor U12029 (N_12029,N_10555,N_11959);
and U12030 (N_12030,N_11851,N_11293);
xnor U12031 (N_12031,N_11000,N_10630);
or U12032 (N_12032,N_11371,N_11971);
nand U12033 (N_12033,N_11212,N_11443);
and U12034 (N_12034,N_10784,N_11516);
or U12035 (N_12035,N_11058,N_10853);
xor U12036 (N_12036,N_10531,N_11069);
and U12037 (N_12037,N_10806,N_11552);
and U12038 (N_12038,N_10989,N_11859);
xor U12039 (N_12039,N_10883,N_10929);
and U12040 (N_12040,N_11940,N_11741);
nor U12041 (N_12041,N_11116,N_11327);
xnor U12042 (N_12042,N_10711,N_10695);
nor U12043 (N_12043,N_11049,N_10964);
nand U12044 (N_12044,N_11869,N_11203);
and U12045 (N_12045,N_11348,N_11304);
nand U12046 (N_12046,N_11624,N_11679);
and U12047 (N_12047,N_11141,N_10578);
and U12048 (N_12048,N_11014,N_11879);
or U12049 (N_12049,N_11949,N_11487);
and U12050 (N_12050,N_11294,N_10542);
nand U12051 (N_12051,N_11994,N_11642);
nand U12052 (N_12052,N_10748,N_11975);
xnor U12053 (N_12053,N_11126,N_11154);
nand U12054 (N_12054,N_10702,N_11751);
nor U12055 (N_12055,N_11220,N_10887);
xor U12056 (N_12056,N_10856,N_11079);
or U12057 (N_12057,N_11308,N_11221);
and U12058 (N_12058,N_10591,N_11331);
nor U12059 (N_12059,N_10898,N_10862);
nor U12060 (N_12060,N_11004,N_11062);
nor U12061 (N_12061,N_10790,N_11781);
xor U12062 (N_12062,N_11561,N_10680);
or U12063 (N_12063,N_10823,N_11547);
nor U12064 (N_12064,N_11928,N_10717);
xnor U12065 (N_12065,N_10775,N_11709);
xor U12066 (N_12066,N_10819,N_11657);
xnor U12067 (N_12067,N_11701,N_10888);
nand U12068 (N_12068,N_10974,N_11322);
and U12069 (N_12069,N_10689,N_10602);
nor U12070 (N_12070,N_11284,N_11907);
nor U12071 (N_12071,N_10592,N_11314);
nor U12072 (N_12072,N_11380,N_10734);
and U12073 (N_12073,N_10771,N_10921);
and U12074 (N_12074,N_11121,N_10938);
or U12075 (N_12075,N_10681,N_10664);
nor U12076 (N_12076,N_10770,N_11952);
xor U12077 (N_12077,N_11565,N_11965);
or U12078 (N_12078,N_11066,N_11763);
nor U12079 (N_12079,N_11310,N_11463);
and U12080 (N_12080,N_11855,N_11895);
nand U12081 (N_12081,N_11048,N_11418);
xor U12082 (N_12082,N_10861,N_10967);
xor U12083 (N_12083,N_10992,N_11392);
or U12084 (N_12084,N_11860,N_10631);
and U12085 (N_12085,N_11911,N_11457);
nor U12086 (N_12086,N_10659,N_10932);
and U12087 (N_12087,N_11586,N_11060);
xor U12088 (N_12088,N_11146,N_11970);
nand U12089 (N_12089,N_11540,N_11168);
xor U12090 (N_12090,N_11724,N_10629);
nand U12091 (N_12091,N_10697,N_10520);
and U12092 (N_12092,N_10687,N_10572);
nand U12093 (N_12093,N_11027,N_10599);
xnor U12094 (N_12094,N_11341,N_11983);
xnor U12095 (N_12095,N_11645,N_11767);
nand U12096 (N_12096,N_10658,N_11889);
and U12097 (N_12097,N_11630,N_10956);
or U12098 (N_12098,N_10778,N_11431);
or U12099 (N_12099,N_11156,N_11275);
xor U12100 (N_12100,N_10696,N_11039);
xor U12101 (N_12101,N_11521,N_11881);
nand U12102 (N_12102,N_11511,N_11299);
or U12103 (N_12103,N_11517,N_10601);
xnor U12104 (N_12104,N_11927,N_11400);
nor U12105 (N_12105,N_11241,N_11787);
nand U12106 (N_12106,N_11384,N_11622);
nand U12107 (N_12107,N_11102,N_11976);
nand U12108 (N_12108,N_11765,N_11080);
xor U12109 (N_12109,N_11695,N_11481);
xnor U12110 (N_12110,N_11742,N_11967);
and U12111 (N_12111,N_11095,N_11803);
xnor U12112 (N_12112,N_10803,N_11346);
xnor U12113 (N_12113,N_11974,N_11366);
nor U12114 (N_12114,N_11799,N_11351);
nor U12115 (N_12115,N_11167,N_11887);
nor U12116 (N_12116,N_11728,N_11599);
nand U12117 (N_12117,N_11582,N_11961);
or U12118 (N_12118,N_10634,N_11251);
nor U12119 (N_12119,N_11098,N_11835);
and U12120 (N_12120,N_11417,N_11922);
nand U12121 (N_12121,N_11295,N_10651);
nor U12122 (N_12122,N_11437,N_11575);
nand U12123 (N_12123,N_10675,N_11405);
or U12124 (N_12124,N_11899,N_11668);
nand U12125 (N_12125,N_10527,N_11812);
or U12126 (N_12126,N_11573,N_11553);
xor U12127 (N_12127,N_11413,N_11420);
xor U12128 (N_12128,N_11254,N_10788);
nor U12129 (N_12129,N_11929,N_11421);
nor U12130 (N_12130,N_10627,N_11091);
nor U12131 (N_12131,N_11412,N_10677);
nor U12132 (N_12132,N_10571,N_10831);
and U12133 (N_12133,N_10722,N_10762);
nor U12134 (N_12134,N_11106,N_10869);
and U12135 (N_12135,N_10657,N_11529);
nand U12136 (N_12136,N_11682,N_11791);
xnor U12137 (N_12137,N_10809,N_10955);
and U12138 (N_12138,N_10562,N_10866);
and U12139 (N_12139,N_10528,N_11277);
nand U12140 (N_12140,N_11097,N_10625);
or U12141 (N_12141,N_11477,N_11035);
xnor U12142 (N_12142,N_11636,N_11667);
or U12143 (N_12143,N_10808,N_10952);
or U12144 (N_12144,N_10894,N_10615);
nand U12145 (N_12145,N_11725,N_11219);
and U12146 (N_12146,N_10846,N_10600);
and U12147 (N_12147,N_10774,N_11905);
and U12148 (N_12148,N_11760,N_10833);
nor U12149 (N_12149,N_11289,N_11061);
and U12150 (N_12150,N_10716,N_11491);
nand U12151 (N_12151,N_11347,N_10783);
xor U12152 (N_12152,N_10751,N_11263);
xor U12153 (N_12153,N_10636,N_11894);
or U12154 (N_12154,N_11828,N_11654);
nor U12155 (N_12155,N_11797,N_10842);
and U12156 (N_12156,N_11073,N_11447);
nor U12157 (N_12157,N_10699,N_10559);
and U12158 (N_12158,N_10972,N_11950);
nand U12159 (N_12159,N_11356,N_10667);
xnor U12160 (N_12160,N_11114,N_10517);
and U12161 (N_12161,N_11977,N_11954);
nor U12162 (N_12162,N_11604,N_10947);
or U12163 (N_12163,N_11015,N_11696);
xnor U12164 (N_12164,N_11833,N_11017);
nor U12165 (N_12165,N_10776,N_11958);
nor U12166 (N_12166,N_10649,N_11666);
and U12167 (N_12167,N_11943,N_11629);
and U12168 (N_12168,N_11509,N_11993);
or U12169 (N_12169,N_10715,N_11224);
nor U12170 (N_12170,N_11856,N_11500);
nor U12171 (N_12171,N_10577,N_10884);
and U12172 (N_12172,N_11598,N_11662);
nor U12173 (N_12173,N_11689,N_11182);
and U12174 (N_12174,N_10737,N_10647);
and U12175 (N_12175,N_10849,N_11147);
xor U12176 (N_12176,N_11603,N_10540);
nor U12177 (N_12177,N_11486,N_10549);
or U12178 (N_12178,N_11096,N_11478);
xnor U12179 (N_12179,N_11090,N_11433);
and U12180 (N_12180,N_11882,N_11962);
and U12181 (N_12181,N_10903,N_11467);
nor U12182 (N_12182,N_11580,N_11948);
nand U12183 (N_12183,N_11452,N_11115);
nand U12184 (N_12184,N_11085,N_11874);
xnor U12185 (N_12185,N_11370,N_11271);
nand U12186 (N_12186,N_11536,N_10997);
and U12187 (N_12187,N_11609,N_11204);
xor U12188 (N_12188,N_11533,N_11546);
and U12189 (N_12189,N_10946,N_11558);
nor U12190 (N_12190,N_11631,N_11699);
nand U12191 (N_12191,N_10935,N_10976);
and U12192 (N_12192,N_11716,N_11532);
xor U12193 (N_12193,N_11045,N_11610);
and U12194 (N_12194,N_11910,N_11422);
and U12195 (N_12195,N_10991,N_10851);
nand U12196 (N_12196,N_11041,N_10613);
nand U12197 (N_12197,N_10605,N_11785);
xnor U12198 (N_12198,N_11206,N_11735);
xnor U12199 (N_12199,N_11995,N_10503);
xnor U12200 (N_12200,N_11902,N_11822);
or U12201 (N_12201,N_11504,N_10710);
or U12202 (N_12202,N_10530,N_11262);
nor U12203 (N_12203,N_11278,N_11214);
or U12204 (N_12204,N_11719,N_11108);
and U12205 (N_12205,N_10901,N_11817);
xnor U12206 (N_12206,N_11826,N_11570);
and U12207 (N_12207,N_11151,N_11576);
nand U12208 (N_12208,N_10951,N_11737);
xnor U12209 (N_12209,N_11143,N_11615);
or U12210 (N_12210,N_11480,N_11906);
nand U12211 (N_12211,N_10792,N_11530);
nor U12212 (N_12212,N_11485,N_11296);
or U12213 (N_12213,N_11426,N_11072);
nor U12214 (N_12214,N_11428,N_11900);
nor U12215 (N_12215,N_11475,N_11534);
and U12216 (N_12216,N_11231,N_11769);
and U12217 (N_12217,N_11164,N_11434);
nor U12218 (N_12218,N_11786,N_10509);
nor U12219 (N_12219,N_11321,N_11846);
nor U12220 (N_12220,N_11871,N_10837);
and U12221 (N_12221,N_11955,N_11568);
xnor U12222 (N_12222,N_10983,N_10535);
nor U12223 (N_12223,N_11708,N_10977);
nor U12224 (N_12224,N_10684,N_11409);
nand U12225 (N_12225,N_10598,N_11827);
or U12226 (N_12226,N_11814,N_10532);
and U12227 (N_12227,N_11508,N_10642);
or U12228 (N_12228,N_11921,N_10899);
xor U12229 (N_12229,N_11885,N_11734);
or U12230 (N_12230,N_11474,N_10606);
nor U12231 (N_12231,N_11957,N_10682);
nand U12232 (N_12232,N_10906,N_11753);
or U12233 (N_12233,N_11614,N_10871);
nor U12234 (N_12234,N_10720,N_11557);
nand U12235 (N_12235,N_11276,N_10628);
nand U12236 (N_12236,N_10739,N_11258);
and U12237 (N_12237,N_11989,N_10781);
nand U12238 (N_12238,N_10798,N_11286);
nor U12239 (N_12239,N_10860,N_10545);
nand U12240 (N_12240,N_10824,N_11292);
or U12241 (N_12241,N_11363,N_11242);
or U12242 (N_12242,N_11768,N_10999);
and U12243 (N_12243,N_11118,N_11495);
nor U12244 (N_12244,N_11152,N_11402);
and U12245 (N_12245,N_11325,N_11564);
nor U12246 (N_12246,N_11766,N_11253);
xor U12247 (N_12247,N_11665,N_10981);
nor U12248 (N_12248,N_11483,N_11729);
nand U12249 (N_12249,N_10950,N_11718);
and U12250 (N_12250,N_11055,N_11686);
xor U12251 (N_12251,N_11194,N_11174);
nand U12252 (N_12252,N_11963,N_11171);
and U12253 (N_12253,N_11824,N_11594);
xor U12254 (N_12254,N_11243,N_11290);
nor U12255 (N_12255,N_10750,N_11070);
xor U12256 (N_12256,N_10922,N_10738);
and U12257 (N_12257,N_11208,N_11240);
and U12258 (N_12258,N_10890,N_11040);
nand U12259 (N_12259,N_10889,N_10990);
nor U12260 (N_12260,N_10841,N_11344);
nand U12261 (N_12261,N_11100,N_11230);
nor U12262 (N_12262,N_11756,N_11775);
nand U12263 (N_12263,N_11128,N_11446);
xnor U12264 (N_12264,N_11369,N_11225);
or U12265 (N_12265,N_11301,N_10586);
xnor U12266 (N_12266,N_10988,N_11169);
and U12267 (N_12267,N_11809,N_11790);
nand U12268 (N_12268,N_10789,N_11499);
and U12269 (N_12269,N_11201,N_10513);
nand U12270 (N_12270,N_10700,N_11687);
and U12271 (N_12271,N_11757,N_11064);
nand U12272 (N_12272,N_11780,N_11632);
nor U12273 (N_12273,N_10914,N_11444);
and U12274 (N_12274,N_10834,N_10585);
nor U12275 (N_12275,N_11406,N_11541);
or U12276 (N_12276,N_11266,N_10508);
nand U12277 (N_12277,N_11640,N_11663);
xor U12278 (N_12278,N_10996,N_11454);
nand U12279 (N_12279,N_10822,N_10931);
nand U12280 (N_12280,N_10646,N_10985);
or U12281 (N_12281,N_10969,N_11228);
and U12282 (N_12282,N_11273,N_11706);
and U12283 (N_12283,N_11138,N_11005);
and U12284 (N_12284,N_10550,N_11367);
and U12285 (N_12285,N_11320,N_11345);
or U12286 (N_12286,N_10656,N_11795);
or U12287 (N_12287,N_11986,N_11776);
and U12288 (N_12288,N_10624,N_10958);
and U12289 (N_12289,N_11641,N_10730);
xnor U12290 (N_12290,N_10679,N_11783);
or U12291 (N_12291,N_11606,N_11111);
or U12292 (N_12292,N_11403,N_11990);
and U12293 (N_12293,N_11032,N_10795);
nand U12294 (N_12294,N_10690,N_10588);
and U12295 (N_12295,N_11960,N_11711);
nand U12296 (N_12296,N_11601,N_10937);
xnor U12297 (N_12297,N_11488,N_11572);
xor U12298 (N_12298,N_11120,N_11647);
and U12299 (N_12299,N_11365,N_10876);
xnor U12300 (N_12300,N_10668,N_11870);
nor U12301 (N_12301,N_11818,N_11019);
xor U12302 (N_12302,N_11053,N_11323);
or U12303 (N_12303,N_11238,N_10812);
nor U12304 (N_12304,N_10835,N_10797);
nor U12305 (N_12305,N_10863,N_10925);
nor U12306 (N_12306,N_11257,N_11655);
or U12307 (N_12307,N_11195,N_10949);
nor U12308 (N_12308,N_11052,N_10643);
xor U12309 (N_12309,N_11806,N_10911);
nand U12310 (N_12310,N_10576,N_11893);
nand U12311 (N_12311,N_10526,N_11567);
nand U12312 (N_12312,N_11288,N_11337);
nand U12313 (N_12313,N_11834,N_10852);
and U12314 (N_12314,N_11867,N_11730);
or U12315 (N_12315,N_11700,N_10941);
nand U12316 (N_12316,N_11831,N_11969);
xnor U12317 (N_12317,N_11901,N_11597);
and U12318 (N_12318,N_10701,N_11209);
xor U12319 (N_12319,N_11891,N_10534);
and U12320 (N_12320,N_11311,N_11917);
nand U12321 (N_12321,N_11819,N_10580);
or U12322 (N_12322,N_11162,N_10728);
nor U12323 (N_12323,N_11992,N_11334);
nand U12324 (N_12324,N_10704,N_11236);
xor U12325 (N_12325,N_11036,N_11461);
and U12326 (N_12326,N_11643,N_11233);
or U12327 (N_12327,N_11416,N_10500);
xor U12328 (N_12328,N_10896,N_11999);
or U12329 (N_12329,N_11688,N_10794);
or U12330 (N_12330,N_11713,N_10785);
nor U12331 (N_12331,N_10971,N_11110);
nor U12332 (N_12332,N_10595,N_11823);
nor U12333 (N_12333,N_10832,N_11249);
and U12334 (N_12334,N_10799,N_10916);
nand U12335 (N_12335,N_10619,N_11291);
or U12336 (N_12336,N_11166,N_11252);
xnor U12337 (N_12337,N_10622,N_10512);
nor U12338 (N_12338,N_10959,N_11023);
nand U12339 (N_12339,N_11744,N_11043);
and U12340 (N_12340,N_10544,N_10870);
and U12341 (N_12341,N_11551,N_10940);
or U12342 (N_12342,N_10787,N_10676);
xor U12343 (N_12343,N_11223,N_11669);
nor U12344 (N_12344,N_11281,N_11218);
nor U12345 (N_12345,N_11340,N_11165);
xnor U12346 (N_12346,N_11411,N_11089);
and U12347 (N_12347,N_10654,N_11067);
and U12348 (N_12348,N_10829,N_10740);
nand U12349 (N_12349,N_11777,N_10674);
xor U12350 (N_12350,N_10546,N_11896);
or U12351 (N_12351,N_11229,N_11947);
and U12352 (N_12352,N_11578,N_10825);
xnor U12353 (N_12353,N_11717,N_11361);
xnor U12354 (N_12354,N_10752,N_11782);
xnor U12355 (N_12355,N_11051,N_10918);
nand U12356 (N_12356,N_11261,N_10987);
nor U12357 (N_12357,N_10780,N_11747);
xor U12358 (N_12358,N_11131,N_11710);
or U12359 (N_12359,N_11071,N_10742);
xnor U12360 (N_12360,N_10928,N_11620);
or U12361 (N_12361,N_11427,N_11602);
nand U12362 (N_12362,N_11857,N_11432);
xnor U12363 (N_12363,N_11868,N_10779);
and U12364 (N_12364,N_11938,N_10805);
or U12365 (N_12365,N_11681,N_11639);
and U12366 (N_12366,N_10924,N_11383);
nand U12367 (N_12367,N_10984,N_11560);
or U12368 (N_12368,N_10980,N_11661);
xnor U12369 (N_12369,N_11376,N_11796);
and U12370 (N_12370,N_10804,N_10683);
nand U12371 (N_12371,N_10583,N_11646);
and U12372 (N_12372,N_10706,N_11458);
or U12373 (N_12373,N_11503,N_11324);
or U12374 (N_12374,N_11247,N_11117);
and U12375 (N_12375,N_11811,N_11836);
or U12376 (N_12376,N_11664,N_10843);
nand U12377 (N_12377,N_10982,N_10693);
nor U12378 (N_12378,N_11941,N_11650);
or U12379 (N_12379,N_10685,N_11909);
or U12380 (N_12380,N_11456,N_10936);
and U12381 (N_12381,N_10886,N_11013);
nor U12382 (N_12382,N_11211,N_10960);
nand U12383 (N_12383,N_10786,N_11876);
nor U12384 (N_12384,N_10574,N_11007);
nor U12385 (N_12385,N_11685,N_11722);
xnor U12386 (N_12386,N_11991,N_10694);
or U12387 (N_12387,N_11192,N_11502);
nand U12388 (N_12388,N_11083,N_10719);
and U12389 (N_12389,N_11137,N_10858);
nand U12390 (N_12390,N_11399,N_11462);
or U12391 (N_12391,N_10566,N_11155);
nor U12392 (N_12392,N_10857,N_11333);
and U12393 (N_12393,N_10645,N_11269);
xnor U12394 (N_12394,N_10855,N_10705);
or U12395 (N_12395,N_11723,N_11123);
or U12396 (N_12396,N_10590,N_11094);
or U12397 (N_12397,N_11774,N_10801);
xor U12398 (N_12398,N_10660,N_11801);
and U12399 (N_12399,N_11496,N_11778);
xor U12400 (N_12400,N_11414,N_11621);
nand U12401 (N_12401,N_11946,N_10961);
nor U12402 (N_12402,N_11997,N_11903);
and U12403 (N_12403,N_10848,N_11634);
nor U12404 (N_12404,N_10617,N_11644);
nand U12405 (N_12405,N_11671,N_10671);
nand U12406 (N_12406,N_11305,N_11397);
nand U12407 (N_12407,N_11523,N_10908);
or U12408 (N_12408,N_11638,N_10864);
xor U12409 (N_12409,N_10733,N_10558);
nor U12410 (N_12410,N_11972,N_11526);
and U12411 (N_12411,N_11942,N_11538);
nand U12412 (N_12412,N_10648,N_11232);
and U12413 (N_12413,N_11357,N_11600);
nand U12414 (N_12414,N_11956,N_11933);
nor U12415 (N_12415,N_11173,N_11338);
and U12416 (N_12416,N_11732,N_11497);
xnor U12417 (N_12417,N_10807,N_11676);
xnor U12418 (N_12418,N_11528,N_11248);
and U12419 (N_12419,N_10678,N_11771);
or U12420 (N_12420,N_11720,N_11313);
nor U12421 (N_12421,N_10814,N_11755);
and U12422 (N_12422,N_11157,N_11840);
nand U12423 (N_12423,N_11673,N_11520);
nor U12424 (N_12424,N_11592,N_11009);
nor U12425 (N_12425,N_10611,N_10623);
and U12426 (N_12426,N_11105,N_11754);
and U12427 (N_12427,N_11193,N_11800);
nor U12428 (N_12428,N_11473,N_10713);
and U12429 (N_12429,N_10943,N_11133);
and U12430 (N_12430,N_11339,N_10907);
xnor U12431 (N_12431,N_11318,N_10547);
nor U12432 (N_12432,N_11556,N_10995);
nand U12433 (N_12433,N_10939,N_11852);
nor U12434 (N_12434,N_10703,N_11239);
nand U12435 (N_12435,N_11270,N_11740);
and U12436 (N_12436,N_10663,N_11845);
and U12437 (N_12437,N_10597,N_10548);
or U12438 (N_12438,N_11466,N_11677);
xnor U12439 (N_12439,N_10859,N_11559);
nand U12440 (N_12440,N_10973,N_11030);
nor U12441 (N_12441,N_11059,N_11020);
or U12442 (N_12442,N_11425,N_11998);
nor U12443 (N_12443,N_10948,N_11374);
xnor U12444 (N_12444,N_11581,N_11429);
xor U12445 (N_12445,N_10793,N_11435);
nand U12446 (N_12446,N_11591,N_11279);
nor U12447 (N_12447,N_11448,N_11761);
nand U12448 (N_12448,N_11616,N_10723);
or U12449 (N_12449,N_11054,N_10618);
nand U12450 (N_12450,N_11011,N_11404);
nor U12451 (N_12451,N_11142,N_11476);
nand U12452 (N_12452,N_10934,N_10891);
xor U12453 (N_12453,N_11507,N_10570);
nor U12454 (N_12454,N_10641,N_10756);
and U12455 (N_12455,N_10818,N_11381);
xor U12456 (N_12456,N_10963,N_10993);
nor U12457 (N_12457,N_11075,N_11342);
nand U12458 (N_12458,N_11635,N_10729);
nand U12459 (N_12459,N_10769,N_11838);
or U12460 (N_12460,N_10920,N_11460);
nor U12461 (N_12461,N_11764,N_11675);
nand U12462 (N_12462,N_11583,N_11649);
nand U12463 (N_12463,N_11489,N_11316);
nand U12464 (N_12464,N_11596,N_11861);
and U12465 (N_12465,N_11136,N_11798);
and U12466 (N_12466,N_10554,N_10708);
nand U12467 (N_12467,N_10881,N_11197);
nor U12468 (N_12468,N_11884,N_11163);
or U12469 (N_12469,N_10998,N_11862);
nand U12470 (N_12470,N_11554,N_11309);
and U12471 (N_12471,N_11183,N_11518);
nand U12472 (N_12472,N_11770,N_11789);
and U12473 (N_12473,N_10744,N_11608);
nand U12474 (N_12474,N_11139,N_11637);
nand U12475 (N_12475,N_11315,N_10877);
or U12476 (N_12476,N_11731,N_11721);
nor U12477 (N_12477,N_10945,N_11864);
or U12478 (N_12478,N_11916,N_11234);
or U12479 (N_12479,N_10915,N_11660);
nand U12480 (N_12480,N_10757,N_11056);
xnor U12481 (N_12481,N_10800,N_10662);
and U12482 (N_12482,N_11805,N_11577);
or U12483 (N_12483,N_11527,N_11034);
xnor U12484 (N_12484,N_10511,N_10875);
and U12485 (N_12485,N_11841,N_11693);
and U12486 (N_12486,N_11585,N_11104);
or U12487 (N_12487,N_11658,N_10874);
xor U12488 (N_12488,N_11829,N_11379);
xnor U12489 (N_12489,N_11362,N_10968);
and U12490 (N_12490,N_10686,N_11464);
xor U12491 (N_12491,N_10669,N_11865);
nor U12492 (N_12492,N_10626,N_11196);
nor U12493 (N_12493,N_11150,N_11022);
nand U12494 (N_12494,N_11934,N_10782);
nor U12495 (N_12495,N_10575,N_10826);
and U12496 (N_12496,N_11752,N_10610);
or U12497 (N_12497,N_10569,N_11283);
and U12498 (N_12498,N_11648,N_11388);
and U12499 (N_12499,N_10673,N_11285);
xnor U12500 (N_12500,N_11830,N_11127);
nor U12501 (N_12501,N_11419,N_11904);
xor U12502 (N_12502,N_11914,N_11953);
and U12503 (N_12503,N_10767,N_11025);
xor U12504 (N_12504,N_10844,N_11545);
or U12505 (N_12505,N_11794,N_11659);
xor U12506 (N_12506,N_10603,N_11440);
and U12507 (N_12507,N_10536,N_11264);
nor U12508 (N_12508,N_10965,N_11683);
or U12509 (N_12509,N_10732,N_11569);
xnor U12510 (N_12510,N_10529,N_10791);
or U12511 (N_12511,N_10909,N_11873);
nand U12512 (N_12512,N_10614,N_11618);
and U12513 (N_12513,N_10638,N_11498);
and U12514 (N_12514,N_10753,N_11449);
nor U12515 (N_12515,N_11026,N_11395);
and U12516 (N_12516,N_10581,N_10525);
nor U12517 (N_12517,N_11843,N_11101);
nand U12518 (N_12518,N_11890,N_11784);
and U12519 (N_12519,N_11063,N_10593);
nor U12520 (N_12520,N_11057,N_11298);
and U12521 (N_12521,N_11172,N_11018);
nand U12522 (N_12522,N_11074,N_11613);
and U12523 (N_12523,N_10878,N_11892);
nor U12524 (N_12524,N_11762,N_11390);
xnor U12525 (N_12525,N_11302,N_11368);
xor U12526 (N_12526,N_10802,N_10560);
xor U12527 (N_12527,N_10553,N_11748);
or U12528 (N_12528,N_10505,N_11303);
xnor U12529 (N_12529,N_11490,N_10893);
or U12530 (N_12530,N_11082,N_11445);
or U12531 (N_12531,N_11003,N_10653);
xnor U12532 (N_12532,N_10747,N_11535);
nor U12533 (N_12533,N_11181,N_11544);
nor U12534 (N_12534,N_10979,N_11988);
or U12535 (N_12535,N_11758,N_11617);
xor U12536 (N_12536,N_11349,N_10589);
nor U12537 (N_12537,N_10880,N_11130);
and U12538 (N_12538,N_11562,N_11537);
xor U12539 (N_12539,N_11215,N_11712);
xnor U12540 (N_12540,N_11850,N_10587);
or U12541 (N_12541,N_11566,N_11908);
and U12542 (N_12542,N_11028,N_11424);
nand U12543 (N_12543,N_10522,N_11513);
nor U12544 (N_12544,N_11919,N_11046);
nand U12545 (N_12545,N_11398,N_11707);
or U12546 (N_12546,N_11555,N_11531);
nand U12547 (N_12547,N_11633,N_11698);
xnor U12548 (N_12548,N_10827,N_10524);
and U12549 (N_12549,N_10635,N_11759);
or U12550 (N_12550,N_11140,N_10930);
nand U12551 (N_12551,N_10727,N_11332);
xor U12552 (N_12552,N_10927,N_11012);
and U12553 (N_12553,N_11574,N_11945);
and U12554 (N_12554,N_11470,N_11875);
nand U12555 (N_12555,N_10672,N_10773);
nor U12556 (N_12556,N_11068,N_10761);
or U12557 (N_12557,N_11703,N_10746);
xor U12558 (N_12558,N_10552,N_11524);
nor U12559 (N_12559,N_11590,N_11149);
nand U12560 (N_12560,N_11493,N_11265);
xnor U12561 (N_12561,N_11389,N_11226);
or U12562 (N_12562,N_11612,N_11280);
xnor U12563 (N_12563,N_11579,N_10573);
nand U12564 (N_12564,N_10759,N_11042);
and U12565 (N_12565,N_11179,N_11652);
and U12566 (N_12566,N_11951,N_11328);
or U12567 (N_12567,N_11372,N_11694);
or U12568 (N_12568,N_11897,N_10944);
and U12569 (N_12569,N_11350,N_11235);
nor U12570 (N_12570,N_10637,N_11936);
or U12571 (N_12571,N_10905,N_11702);
or U12572 (N_12572,N_11849,N_10582);
nor U12573 (N_12573,N_11122,N_11092);
nand U12574 (N_12574,N_11872,N_11360);
nor U12575 (N_12575,N_11119,N_10913);
or U12576 (N_12576,N_11866,N_10691);
xnor U12577 (N_12577,N_10900,N_11382);
or U12578 (N_12578,N_10564,N_11514);
or U12579 (N_12579,N_11656,N_10741);
nor U12580 (N_12580,N_11746,N_11282);
xor U12581 (N_12581,N_11912,N_11627);
and U12582 (N_12582,N_10726,N_11743);
nand U12583 (N_12583,N_10954,N_11494);
xor U12584 (N_12584,N_11563,N_11387);
nor U12585 (N_12585,N_11029,N_10745);
and U12586 (N_12586,N_11807,N_11571);
nor U12587 (N_12587,N_10902,N_11001);
nand U12588 (N_12588,N_10725,N_11964);
nor U12589 (N_12589,N_11373,N_10533);
or U12590 (N_12590,N_11037,N_11359);
and U12591 (N_12591,N_10854,N_10584);
nand U12592 (N_12592,N_11125,N_10766);
and U12593 (N_12593,N_10688,N_10840);
and U12594 (N_12594,N_11336,N_11482);
and U12595 (N_12595,N_11006,N_11396);
and U12596 (N_12596,N_10551,N_10882);
xnor U12597 (N_12597,N_11438,N_11898);
xnor U12598 (N_12598,N_11343,N_11021);
nor U12599 (N_12599,N_10519,N_11016);
or U12600 (N_12600,N_11050,N_11918);
or U12601 (N_12601,N_11185,N_10709);
and U12602 (N_12602,N_11472,N_10714);
nand U12603 (N_12603,N_11134,N_11047);
or U12604 (N_12604,N_11198,N_10665);
nor U12605 (N_12605,N_10616,N_10609);
or U12606 (N_12606,N_11355,N_11736);
nand U12607 (N_12607,N_11705,N_11358);
nand U12608 (N_12608,N_11930,N_11858);
or U12609 (N_12609,N_11492,N_11844);
nand U12610 (N_12610,N_11297,N_11619);
nand U12611 (N_12611,N_11628,N_11525);
nor U12612 (N_12612,N_10640,N_11501);
or U12613 (N_12613,N_11739,N_10892);
nor U12614 (N_12614,N_11160,N_11260);
nand U12615 (N_12615,N_11804,N_10813);
or U12616 (N_12616,N_10755,N_11441);
nand U12617 (N_12617,N_11837,N_11996);
xor U12618 (N_12618,N_11832,N_10579);
and U12619 (N_12619,N_11772,N_11109);
and U12620 (N_12620,N_10567,N_11926);
or U12621 (N_12621,N_11415,N_11439);
xor U12622 (N_12622,N_11300,N_10758);
nor U12623 (N_12623,N_11968,N_11888);
nand U12624 (N_12624,N_11113,N_11479);
xor U12625 (N_12625,N_11202,N_10707);
nand U12626 (N_12626,N_11272,N_11733);
and U12627 (N_12627,N_10724,N_11329);
xor U12628 (N_12628,N_11839,N_11593);
nor U12629 (N_12629,N_11227,N_11738);
xor U12630 (N_12630,N_11915,N_10828);
and U12631 (N_12631,N_10538,N_11810);
nor U12632 (N_12632,N_11222,N_10518);
nor U12633 (N_12633,N_11808,N_11191);
xor U12634 (N_12634,N_11727,N_11170);
nand U12635 (N_12635,N_11468,N_11465);
xnor U12636 (N_12636,N_11522,N_10820);
or U12637 (N_12637,N_11543,N_10897);
and U12638 (N_12638,N_10867,N_11190);
nor U12639 (N_12639,N_11245,N_10721);
xor U12640 (N_12640,N_11773,N_11176);
nand U12641 (N_12641,N_10816,N_10768);
nand U12642 (N_12642,N_10743,N_10633);
and U12643 (N_12643,N_11065,N_11450);
nand U12644 (N_12644,N_11453,N_11588);
xor U12645 (N_12645,N_10760,N_11692);
and U12646 (N_12646,N_11312,N_11144);
nand U12647 (N_12647,N_11966,N_10523);
and U12648 (N_12648,N_11423,N_11853);
nor U12649 (N_12649,N_11407,N_10698);
nor U12650 (N_12650,N_11935,N_11352);
xor U12651 (N_12651,N_11931,N_11484);
nand U12652 (N_12652,N_10620,N_11330);
nor U12653 (N_12653,N_11161,N_11033);
xor U12654 (N_12654,N_11103,N_11175);
nand U12655 (N_12655,N_11924,N_11244);
xor U12656 (N_12656,N_10811,N_10873);
nor U12657 (N_12657,N_11010,N_11726);
or U12658 (N_12658,N_10772,N_11584);
or U12659 (N_12659,N_11672,N_10970);
nand U12660 (N_12660,N_10608,N_11749);
xnor U12661 (N_12661,N_11158,N_10563);
or U12662 (N_12662,N_11112,N_10919);
and U12663 (N_12663,N_10514,N_11792);
and U12664 (N_12664,N_11145,N_11883);
or U12665 (N_12665,N_11200,N_10621);
or U12666 (N_12666,N_11410,N_11877);
nor U12667 (N_12667,N_11549,N_11802);
and U12668 (N_12668,N_10504,N_11821);
xor U12669 (N_12669,N_11854,N_11471);
nor U12670 (N_12670,N_10735,N_11506);
or U12671 (N_12671,N_10692,N_11878);
nor U12672 (N_12672,N_11205,N_11880);
and U12673 (N_12673,N_11038,N_10764);
nor U12674 (N_12674,N_10838,N_11093);
and U12675 (N_12675,N_11246,N_11925);
xor U12676 (N_12676,N_11256,N_11187);
nor U12677 (N_12677,N_11539,N_11326);
nand U12678 (N_12678,N_11813,N_11354);
nor U12679 (N_12679,N_11088,N_11077);
xor U12680 (N_12680,N_11335,N_11267);
nand U12681 (N_12681,N_10994,N_11680);
and U12682 (N_12682,N_11981,N_10904);
and U12683 (N_12683,N_11401,N_10933);
xnor U12684 (N_12684,N_11542,N_10596);
nand U12685 (N_12685,N_10543,N_11750);
nand U12686 (N_12686,N_11678,N_10986);
xnor U12687 (N_12687,N_10872,N_10556);
and U12688 (N_12688,N_11515,N_10516);
or U12689 (N_12689,N_11595,N_10501);
nand U12690 (N_12690,N_11607,N_10749);
and U12691 (N_12691,N_11086,N_10847);
and U12692 (N_12692,N_11611,N_11469);
nor U12693 (N_12693,N_10670,N_11319);
and U12694 (N_12694,N_11148,N_10655);
and U12695 (N_12695,N_11937,N_11375);
xor U12696 (N_12696,N_10539,N_11378);
xor U12697 (N_12697,N_10731,N_10644);
or U12698 (N_12698,N_10879,N_11589);
nor U12699 (N_12699,N_11081,N_10568);
nor U12700 (N_12700,N_11394,N_11084);
xnor U12701 (N_12701,N_11745,N_11982);
and U12702 (N_12702,N_11623,N_11008);
xor U12703 (N_12703,N_10796,N_10962);
nand U12704 (N_12704,N_11788,N_10815);
nand U12705 (N_12705,N_11714,N_11076);
and U12706 (N_12706,N_11386,N_11391);
nand U12707 (N_12707,N_11177,N_11548);
nor U12708 (N_12708,N_11984,N_11519);
nor U12709 (N_12709,N_11259,N_11099);
and U12710 (N_12710,N_10942,N_11107);
nor U12711 (N_12711,N_10917,N_10850);
or U12712 (N_12712,N_11353,N_11132);
or U12713 (N_12713,N_11863,N_11078);
xor U12714 (N_12714,N_11913,N_11815);
nand U12715 (N_12715,N_11985,N_11124);
nand U12716 (N_12716,N_11697,N_11455);
nand U12717 (N_12717,N_11510,N_11920);
or U12718 (N_12718,N_11250,N_11213);
nor U12719 (N_12719,N_10836,N_11178);
nor U12720 (N_12720,N_11847,N_10830);
nor U12721 (N_12721,N_10521,N_11377);
and U12722 (N_12722,N_10957,N_10652);
and U12723 (N_12723,N_11923,N_11704);
xnor U12724 (N_12724,N_11408,N_11684);
xnor U12725 (N_12725,N_11939,N_10561);
nand U12726 (N_12726,N_11779,N_11587);
nand U12727 (N_12727,N_10810,N_11653);
and U12728 (N_12728,N_11451,N_10978);
nor U12729 (N_12729,N_11207,N_11505);
and U12730 (N_12730,N_11670,N_10953);
and U12731 (N_12731,N_11550,N_10926);
or U12732 (N_12732,N_11364,N_11188);
and U12733 (N_12733,N_10639,N_11980);
and U12734 (N_12734,N_11031,N_11674);
and U12735 (N_12735,N_11625,N_10502);
nand U12736 (N_12736,N_10821,N_11153);
nand U12737 (N_12737,N_10839,N_11715);
or U12738 (N_12738,N_10845,N_10537);
nand U12739 (N_12739,N_11087,N_11932);
nor U12740 (N_12740,N_11237,N_10736);
and U12741 (N_12741,N_10565,N_11793);
or U12742 (N_12742,N_10763,N_11317);
xnor U12743 (N_12743,N_10604,N_11978);
or U12744 (N_12744,N_11690,N_11842);
and U12745 (N_12745,N_10765,N_11626);
nand U12746 (N_12746,N_11180,N_10666);
xnor U12747 (N_12747,N_11002,N_10541);
nor U12748 (N_12748,N_11393,N_11973);
nand U12749 (N_12749,N_11605,N_11274);
and U12750 (N_12750,N_11888,N_11016);
nand U12751 (N_12751,N_11584,N_11950);
and U12752 (N_12752,N_11421,N_11622);
or U12753 (N_12753,N_11290,N_11369);
and U12754 (N_12754,N_11232,N_11933);
and U12755 (N_12755,N_10777,N_10668);
and U12756 (N_12756,N_10541,N_11580);
nor U12757 (N_12757,N_10694,N_10563);
xnor U12758 (N_12758,N_11882,N_11652);
or U12759 (N_12759,N_11115,N_11916);
nor U12760 (N_12760,N_11167,N_11703);
xor U12761 (N_12761,N_11257,N_11065);
and U12762 (N_12762,N_10922,N_10527);
or U12763 (N_12763,N_11355,N_10538);
xnor U12764 (N_12764,N_10505,N_11786);
xor U12765 (N_12765,N_11857,N_10673);
nand U12766 (N_12766,N_10706,N_10840);
or U12767 (N_12767,N_11594,N_10804);
nand U12768 (N_12768,N_11786,N_11179);
nand U12769 (N_12769,N_10977,N_10857);
xor U12770 (N_12770,N_10955,N_11430);
or U12771 (N_12771,N_11083,N_11969);
and U12772 (N_12772,N_11335,N_11673);
nand U12773 (N_12773,N_11243,N_11763);
or U12774 (N_12774,N_11081,N_11015);
and U12775 (N_12775,N_10666,N_11007);
or U12776 (N_12776,N_11367,N_11067);
and U12777 (N_12777,N_10952,N_10905);
xnor U12778 (N_12778,N_10622,N_11289);
xnor U12779 (N_12779,N_11207,N_10994);
or U12780 (N_12780,N_11383,N_11862);
nor U12781 (N_12781,N_11230,N_11633);
nor U12782 (N_12782,N_10651,N_10800);
and U12783 (N_12783,N_11107,N_11092);
xnor U12784 (N_12784,N_11192,N_10535);
nor U12785 (N_12785,N_11887,N_10639);
xor U12786 (N_12786,N_11888,N_10933);
nand U12787 (N_12787,N_10657,N_11865);
nand U12788 (N_12788,N_11204,N_11318);
nor U12789 (N_12789,N_10696,N_10802);
or U12790 (N_12790,N_10917,N_11212);
nand U12791 (N_12791,N_10969,N_11442);
xor U12792 (N_12792,N_10969,N_11444);
nand U12793 (N_12793,N_11900,N_11759);
and U12794 (N_12794,N_11762,N_11973);
or U12795 (N_12795,N_10990,N_11481);
and U12796 (N_12796,N_11155,N_11460);
nor U12797 (N_12797,N_11852,N_10734);
and U12798 (N_12798,N_11598,N_11557);
or U12799 (N_12799,N_10735,N_11674);
or U12800 (N_12800,N_11293,N_10977);
nor U12801 (N_12801,N_11664,N_11427);
nor U12802 (N_12802,N_10576,N_10686);
or U12803 (N_12803,N_10832,N_11312);
nand U12804 (N_12804,N_11227,N_10951);
and U12805 (N_12805,N_11441,N_10655);
xor U12806 (N_12806,N_11598,N_10872);
nand U12807 (N_12807,N_11897,N_10690);
nor U12808 (N_12808,N_10820,N_11545);
and U12809 (N_12809,N_11056,N_10530);
and U12810 (N_12810,N_10505,N_11907);
nand U12811 (N_12811,N_11713,N_11122);
nor U12812 (N_12812,N_11109,N_10817);
or U12813 (N_12813,N_11090,N_11385);
xor U12814 (N_12814,N_11170,N_10573);
xnor U12815 (N_12815,N_10767,N_10540);
nor U12816 (N_12816,N_11791,N_11185);
nand U12817 (N_12817,N_11372,N_11288);
or U12818 (N_12818,N_11964,N_10569);
nand U12819 (N_12819,N_11494,N_11678);
or U12820 (N_12820,N_10689,N_11286);
nand U12821 (N_12821,N_11139,N_10678);
or U12822 (N_12822,N_11177,N_11920);
or U12823 (N_12823,N_11847,N_11592);
nand U12824 (N_12824,N_10900,N_11598);
xor U12825 (N_12825,N_11451,N_10930);
nor U12826 (N_12826,N_10765,N_11337);
and U12827 (N_12827,N_11156,N_11414);
nand U12828 (N_12828,N_11065,N_11490);
and U12829 (N_12829,N_10744,N_11504);
nand U12830 (N_12830,N_11456,N_11695);
nand U12831 (N_12831,N_11359,N_11702);
nand U12832 (N_12832,N_11954,N_11865);
nand U12833 (N_12833,N_11284,N_10730);
or U12834 (N_12834,N_10532,N_11392);
xnor U12835 (N_12835,N_11968,N_10966);
and U12836 (N_12836,N_11326,N_11469);
or U12837 (N_12837,N_10604,N_10501);
xnor U12838 (N_12838,N_11966,N_11747);
and U12839 (N_12839,N_11953,N_11813);
and U12840 (N_12840,N_11027,N_11588);
or U12841 (N_12841,N_11198,N_10732);
nand U12842 (N_12842,N_10571,N_11252);
nor U12843 (N_12843,N_11229,N_11668);
xnor U12844 (N_12844,N_11522,N_10610);
and U12845 (N_12845,N_11901,N_11814);
nor U12846 (N_12846,N_11163,N_11764);
or U12847 (N_12847,N_11165,N_11299);
or U12848 (N_12848,N_10901,N_11432);
and U12849 (N_12849,N_11761,N_10896);
and U12850 (N_12850,N_10768,N_10672);
or U12851 (N_12851,N_11019,N_11736);
nand U12852 (N_12852,N_10670,N_11694);
nand U12853 (N_12853,N_11385,N_10999);
or U12854 (N_12854,N_11447,N_10665);
and U12855 (N_12855,N_11423,N_11602);
nor U12856 (N_12856,N_10928,N_10713);
or U12857 (N_12857,N_10882,N_11175);
nand U12858 (N_12858,N_11081,N_11715);
or U12859 (N_12859,N_10732,N_11359);
or U12860 (N_12860,N_11600,N_11133);
xnor U12861 (N_12861,N_10580,N_11944);
and U12862 (N_12862,N_11819,N_11399);
nor U12863 (N_12863,N_11604,N_11140);
nor U12864 (N_12864,N_11377,N_10962);
xnor U12865 (N_12865,N_11382,N_11183);
nor U12866 (N_12866,N_11688,N_10938);
nor U12867 (N_12867,N_10551,N_11182);
and U12868 (N_12868,N_11796,N_11406);
and U12869 (N_12869,N_11537,N_11647);
nand U12870 (N_12870,N_11065,N_11902);
or U12871 (N_12871,N_11164,N_11989);
xnor U12872 (N_12872,N_10786,N_11605);
nor U12873 (N_12873,N_10659,N_11179);
nor U12874 (N_12874,N_11750,N_11973);
and U12875 (N_12875,N_10815,N_11814);
nor U12876 (N_12876,N_10781,N_10645);
xnor U12877 (N_12877,N_11568,N_11290);
and U12878 (N_12878,N_11586,N_10843);
and U12879 (N_12879,N_11291,N_11282);
xnor U12880 (N_12880,N_10632,N_10915);
nand U12881 (N_12881,N_11671,N_10514);
or U12882 (N_12882,N_10727,N_11526);
nor U12883 (N_12883,N_10527,N_11577);
nand U12884 (N_12884,N_11710,N_11196);
xor U12885 (N_12885,N_11795,N_11854);
nor U12886 (N_12886,N_10978,N_11708);
or U12887 (N_12887,N_10926,N_11190);
nor U12888 (N_12888,N_10802,N_10684);
or U12889 (N_12889,N_11676,N_11948);
xnor U12890 (N_12890,N_11115,N_11864);
nand U12891 (N_12891,N_10742,N_11992);
or U12892 (N_12892,N_10601,N_11572);
and U12893 (N_12893,N_11307,N_10874);
nand U12894 (N_12894,N_11866,N_10541);
or U12895 (N_12895,N_11673,N_11142);
nor U12896 (N_12896,N_11223,N_10826);
and U12897 (N_12897,N_10854,N_11335);
nor U12898 (N_12898,N_11832,N_11011);
nand U12899 (N_12899,N_10974,N_11151);
xor U12900 (N_12900,N_11093,N_10905);
xor U12901 (N_12901,N_11002,N_11659);
nor U12902 (N_12902,N_10711,N_10516);
or U12903 (N_12903,N_11909,N_11753);
and U12904 (N_12904,N_11793,N_11441);
xor U12905 (N_12905,N_11048,N_10969);
nand U12906 (N_12906,N_11995,N_11457);
xnor U12907 (N_12907,N_11203,N_11154);
or U12908 (N_12908,N_11777,N_11351);
nor U12909 (N_12909,N_11839,N_11098);
nor U12910 (N_12910,N_11659,N_10768);
xor U12911 (N_12911,N_11007,N_11827);
and U12912 (N_12912,N_11078,N_10629);
nor U12913 (N_12913,N_11017,N_11831);
and U12914 (N_12914,N_11757,N_11233);
and U12915 (N_12915,N_10906,N_11033);
xor U12916 (N_12916,N_11315,N_11795);
xor U12917 (N_12917,N_11599,N_11104);
or U12918 (N_12918,N_11291,N_11913);
nand U12919 (N_12919,N_11010,N_11163);
nand U12920 (N_12920,N_10567,N_11217);
or U12921 (N_12921,N_10968,N_11009);
nand U12922 (N_12922,N_11351,N_11093);
or U12923 (N_12923,N_11687,N_10523);
and U12924 (N_12924,N_11474,N_11526);
or U12925 (N_12925,N_11412,N_11468);
or U12926 (N_12926,N_11167,N_11900);
and U12927 (N_12927,N_11288,N_11205);
and U12928 (N_12928,N_11636,N_11605);
xnor U12929 (N_12929,N_11381,N_10752);
or U12930 (N_12930,N_11779,N_10744);
nand U12931 (N_12931,N_11067,N_11022);
nor U12932 (N_12932,N_10751,N_10913);
and U12933 (N_12933,N_11791,N_11464);
nand U12934 (N_12934,N_11054,N_11724);
xnor U12935 (N_12935,N_10747,N_11390);
or U12936 (N_12936,N_10931,N_10951);
nand U12937 (N_12937,N_11613,N_11878);
nor U12938 (N_12938,N_10674,N_11504);
xor U12939 (N_12939,N_11571,N_10843);
nand U12940 (N_12940,N_11058,N_11491);
nor U12941 (N_12941,N_10809,N_11593);
xnor U12942 (N_12942,N_11817,N_10598);
nand U12943 (N_12943,N_11184,N_11361);
nand U12944 (N_12944,N_10888,N_11608);
nand U12945 (N_12945,N_11232,N_11010);
and U12946 (N_12946,N_11645,N_11929);
nor U12947 (N_12947,N_10962,N_10591);
and U12948 (N_12948,N_11120,N_11114);
nor U12949 (N_12949,N_10600,N_11528);
nor U12950 (N_12950,N_11230,N_11457);
and U12951 (N_12951,N_10821,N_10550);
and U12952 (N_12952,N_10629,N_11687);
nand U12953 (N_12953,N_11333,N_11907);
xor U12954 (N_12954,N_11646,N_10793);
nand U12955 (N_12955,N_10961,N_10831);
or U12956 (N_12956,N_11819,N_11083);
xor U12957 (N_12957,N_10965,N_10735);
xnor U12958 (N_12958,N_11610,N_11359);
or U12959 (N_12959,N_10727,N_10946);
or U12960 (N_12960,N_11183,N_11168);
and U12961 (N_12961,N_11357,N_11954);
nor U12962 (N_12962,N_11469,N_10773);
xor U12963 (N_12963,N_11492,N_11173);
and U12964 (N_12964,N_10933,N_11198);
nand U12965 (N_12965,N_10962,N_11549);
nand U12966 (N_12966,N_10553,N_10794);
and U12967 (N_12967,N_11569,N_11373);
nand U12968 (N_12968,N_11124,N_11406);
or U12969 (N_12969,N_11432,N_11405);
or U12970 (N_12970,N_10659,N_10987);
or U12971 (N_12971,N_11573,N_11008);
and U12972 (N_12972,N_10833,N_10623);
and U12973 (N_12973,N_10938,N_11922);
nor U12974 (N_12974,N_11116,N_11346);
and U12975 (N_12975,N_11103,N_11598);
nand U12976 (N_12976,N_11643,N_10727);
nor U12977 (N_12977,N_11845,N_11468);
nor U12978 (N_12978,N_11127,N_10816);
nand U12979 (N_12979,N_10795,N_11846);
xnor U12980 (N_12980,N_11305,N_10825);
or U12981 (N_12981,N_10855,N_10661);
nand U12982 (N_12982,N_11145,N_10926);
or U12983 (N_12983,N_11839,N_10904);
xor U12984 (N_12984,N_10600,N_11944);
nand U12985 (N_12985,N_10726,N_11578);
xor U12986 (N_12986,N_11615,N_10580);
xor U12987 (N_12987,N_10680,N_11932);
and U12988 (N_12988,N_10864,N_11526);
and U12989 (N_12989,N_10990,N_11257);
or U12990 (N_12990,N_11205,N_11047);
nor U12991 (N_12991,N_11200,N_10928);
nor U12992 (N_12992,N_11318,N_10566);
xnor U12993 (N_12993,N_11520,N_10923);
and U12994 (N_12994,N_11691,N_11585);
xnor U12995 (N_12995,N_11681,N_11267);
nand U12996 (N_12996,N_11501,N_10868);
and U12997 (N_12997,N_11844,N_11831);
nor U12998 (N_12998,N_11466,N_10688);
nand U12999 (N_12999,N_10580,N_11304);
nor U13000 (N_13000,N_10884,N_11979);
xnor U13001 (N_13001,N_11634,N_11559);
or U13002 (N_13002,N_11122,N_11939);
xor U13003 (N_13003,N_11512,N_11545);
xnor U13004 (N_13004,N_10825,N_11156);
nand U13005 (N_13005,N_10806,N_10578);
or U13006 (N_13006,N_11638,N_11744);
or U13007 (N_13007,N_11799,N_10871);
or U13008 (N_13008,N_11462,N_11665);
nor U13009 (N_13009,N_11717,N_11740);
or U13010 (N_13010,N_10926,N_11303);
or U13011 (N_13011,N_11690,N_11907);
nand U13012 (N_13012,N_10692,N_11989);
nor U13013 (N_13013,N_11178,N_11551);
nor U13014 (N_13014,N_10809,N_11462);
nand U13015 (N_13015,N_11718,N_10904);
nor U13016 (N_13016,N_11455,N_10936);
nor U13017 (N_13017,N_11657,N_10994);
nand U13018 (N_13018,N_11160,N_11033);
xor U13019 (N_13019,N_11653,N_11404);
and U13020 (N_13020,N_11247,N_11550);
or U13021 (N_13021,N_11046,N_11849);
nand U13022 (N_13022,N_10838,N_11115);
nor U13023 (N_13023,N_11807,N_10940);
or U13024 (N_13024,N_11679,N_10604);
xnor U13025 (N_13025,N_11883,N_11653);
nor U13026 (N_13026,N_10746,N_10604);
and U13027 (N_13027,N_10618,N_11504);
nor U13028 (N_13028,N_11179,N_11886);
nor U13029 (N_13029,N_11917,N_11042);
and U13030 (N_13030,N_10921,N_11707);
xor U13031 (N_13031,N_11731,N_10820);
and U13032 (N_13032,N_11873,N_11188);
nand U13033 (N_13033,N_11290,N_11215);
and U13034 (N_13034,N_10885,N_11900);
and U13035 (N_13035,N_10718,N_10739);
nor U13036 (N_13036,N_11089,N_11577);
or U13037 (N_13037,N_11012,N_11697);
and U13038 (N_13038,N_10512,N_11412);
nand U13039 (N_13039,N_10673,N_11255);
or U13040 (N_13040,N_11048,N_11129);
nand U13041 (N_13041,N_11938,N_11474);
nor U13042 (N_13042,N_11589,N_11688);
or U13043 (N_13043,N_11514,N_11489);
nor U13044 (N_13044,N_10943,N_10640);
and U13045 (N_13045,N_10586,N_11381);
nand U13046 (N_13046,N_10702,N_11367);
nand U13047 (N_13047,N_10966,N_10584);
nand U13048 (N_13048,N_11053,N_10744);
or U13049 (N_13049,N_10761,N_11444);
or U13050 (N_13050,N_11964,N_11954);
xnor U13051 (N_13051,N_11507,N_11725);
nor U13052 (N_13052,N_11952,N_10756);
nor U13053 (N_13053,N_10792,N_11932);
xor U13054 (N_13054,N_10811,N_11218);
nand U13055 (N_13055,N_11806,N_10546);
nor U13056 (N_13056,N_11771,N_10761);
and U13057 (N_13057,N_10636,N_11764);
and U13058 (N_13058,N_11035,N_11609);
nand U13059 (N_13059,N_10952,N_10540);
or U13060 (N_13060,N_11724,N_11835);
and U13061 (N_13061,N_11859,N_11911);
or U13062 (N_13062,N_11162,N_11575);
nor U13063 (N_13063,N_11103,N_10860);
nand U13064 (N_13064,N_11661,N_10710);
xor U13065 (N_13065,N_10781,N_11444);
xnor U13066 (N_13066,N_11335,N_11474);
nand U13067 (N_13067,N_11656,N_11726);
nand U13068 (N_13068,N_11187,N_10721);
or U13069 (N_13069,N_11931,N_11515);
or U13070 (N_13070,N_11119,N_11698);
nor U13071 (N_13071,N_11347,N_10516);
or U13072 (N_13072,N_10840,N_11408);
and U13073 (N_13073,N_11096,N_10713);
nand U13074 (N_13074,N_11756,N_11345);
and U13075 (N_13075,N_11675,N_11601);
and U13076 (N_13076,N_11047,N_10568);
xnor U13077 (N_13077,N_10971,N_10754);
nand U13078 (N_13078,N_10581,N_11867);
and U13079 (N_13079,N_10527,N_11041);
and U13080 (N_13080,N_11602,N_11004);
nand U13081 (N_13081,N_10987,N_11581);
xnor U13082 (N_13082,N_10543,N_11640);
and U13083 (N_13083,N_11720,N_11682);
and U13084 (N_13084,N_11520,N_10691);
xor U13085 (N_13085,N_11268,N_11929);
nand U13086 (N_13086,N_10696,N_10504);
or U13087 (N_13087,N_11680,N_11825);
nor U13088 (N_13088,N_10569,N_10898);
nand U13089 (N_13089,N_11425,N_10864);
xnor U13090 (N_13090,N_10521,N_11886);
or U13091 (N_13091,N_11574,N_11081);
or U13092 (N_13092,N_11049,N_11462);
nand U13093 (N_13093,N_11286,N_11499);
or U13094 (N_13094,N_11963,N_11275);
nand U13095 (N_13095,N_11604,N_11667);
xor U13096 (N_13096,N_11491,N_11409);
nand U13097 (N_13097,N_11094,N_11879);
and U13098 (N_13098,N_11481,N_11709);
or U13099 (N_13099,N_10822,N_10901);
or U13100 (N_13100,N_11049,N_11499);
nor U13101 (N_13101,N_11231,N_10985);
nor U13102 (N_13102,N_10538,N_10535);
xnor U13103 (N_13103,N_11460,N_11363);
nor U13104 (N_13104,N_10767,N_11377);
or U13105 (N_13105,N_10845,N_11665);
and U13106 (N_13106,N_11781,N_11140);
nand U13107 (N_13107,N_10693,N_10913);
and U13108 (N_13108,N_11746,N_10518);
and U13109 (N_13109,N_11800,N_11351);
nor U13110 (N_13110,N_11126,N_10686);
nor U13111 (N_13111,N_11359,N_11000);
and U13112 (N_13112,N_11913,N_11222);
or U13113 (N_13113,N_11354,N_11447);
and U13114 (N_13114,N_11073,N_11302);
or U13115 (N_13115,N_10758,N_11826);
or U13116 (N_13116,N_10910,N_10827);
or U13117 (N_13117,N_11736,N_10685);
or U13118 (N_13118,N_10647,N_11751);
nand U13119 (N_13119,N_11470,N_11406);
nand U13120 (N_13120,N_10904,N_11979);
and U13121 (N_13121,N_11367,N_11667);
nand U13122 (N_13122,N_11953,N_10682);
nand U13123 (N_13123,N_10556,N_11716);
xnor U13124 (N_13124,N_11427,N_11952);
or U13125 (N_13125,N_11723,N_11095);
nor U13126 (N_13126,N_11273,N_10937);
and U13127 (N_13127,N_11232,N_11572);
nor U13128 (N_13128,N_11168,N_11665);
xnor U13129 (N_13129,N_10683,N_11532);
nor U13130 (N_13130,N_10944,N_10765);
and U13131 (N_13131,N_10914,N_11046);
nand U13132 (N_13132,N_11637,N_11184);
nand U13133 (N_13133,N_10952,N_10669);
or U13134 (N_13134,N_10620,N_10538);
xor U13135 (N_13135,N_11456,N_11750);
xor U13136 (N_13136,N_11946,N_11523);
nand U13137 (N_13137,N_11070,N_11663);
and U13138 (N_13138,N_10913,N_11132);
nor U13139 (N_13139,N_10922,N_11871);
nor U13140 (N_13140,N_11719,N_10869);
and U13141 (N_13141,N_11805,N_11761);
nor U13142 (N_13142,N_11038,N_11150);
xnor U13143 (N_13143,N_11955,N_10508);
and U13144 (N_13144,N_11263,N_11030);
or U13145 (N_13145,N_10852,N_11308);
and U13146 (N_13146,N_11614,N_10554);
nor U13147 (N_13147,N_11767,N_10969);
nor U13148 (N_13148,N_10985,N_11978);
nand U13149 (N_13149,N_10668,N_10719);
nor U13150 (N_13150,N_11289,N_11573);
nand U13151 (N_13151,N_11735,N_11156);
nand U13152 (N_13152,N_11226,N_11507);
xnor U13153 (N_13153,N_11669,N_10914);
and U13154 (N_13154,N_10961,N_10983);
and U13155 (N_13155,N_11886,N_10806);
nand U13156 (N_13156,N_11809,N_11430);
or U13157 (N_13157,N_10664,N_11365);
nor U13158 (N_13158,N_11992,N_10736);
nand U13159 (N_13159,N_11677,N_11183);
or U13160 (N_13160,N_11894,N_11097);
nand U13161 (N_13161,N_11119,N_11180);
nor U13162 (N_13162,N_11254,N_10981);
nand U13163 (N_13163,N_11953,N_11786);
and U13164 (N_13164,N_11614,N_11424);
nor U13165 (N_13165,N_11054,N_10555);
nor U13166 (N_13166,N_11952,N_10846);
nor U13167 (N_13167,N_11400,N_11509);
and U13168 (N_13168,N_10887,N_10520);
xor U13169 (N_13169,N_10666,N_10569);
xor U13170 (N_13170,N_11370,N_11194);
nor U13171 (N_13171,N_10738,N_11565);
nand U13172 (N_13172,N_11716,N_11352);
nand U13173 (N_13173,N_10953,N_11950);
or U13174 (N_13174,N_11405,N_10869);
and U13175 (N_13175,N_11253,N_11573);
and U13176 (N_13176,N_10746,N_10580);
and U13177 (N_13177,N_10958,N_11476);
xnor U13178 (N_13178,N_10659,N_10712);
nor U13179 (N_13179,N_11727,N_11070);
nand U13180 (N_13180,N_11454,N_11150);
xor U13181 (N_13181,N_10747,N_10726);
nand U13182 (N_13182,N_11357,N_11410);
nand U13183 (N_13183,N_10511,N_11586);
or U13184 (N_13184,N_10533,N_11357);
xor U13185 (N_13185,N_10995,N_11215);
and U13186 (N_13186,N_11026,N_11014);
nor U13187 (N_13187,N_11601,N_11810);
nor U13188 (N_13188,N_10962,N_11413);
nor U13189 (N_13189,N_11477,N_10761);
xnor U13190 (N_13190,N_10538,N_10523);
nand U13191 (N_13191,N_10533,N_11868);
or U13192 (N_13192,N_10801,N_11695);
nand U13193 (N_13193,N_10830,N_11277);
nor U13194 (N_13194,N_11090,N_11320);
and U13195 (N_13195,N_10519,N_11628);
nor U13196 (N_13196,N_11220,N_11589);
or U13197 (N_13197,N_10880,N_11687);
nand U13198 (N_13198,N_11089,N_10652);
or U13199 (N_13199,N_10560,N_11530);
nand U13200 (N_13200,N_11847,N_11644);
and U13201 (N_13201,N_11494,N_11457);
nand U13202 (N_13202,N_10878,N_11394);
nand U13203 (N_13203,N_11388,N_11167);
or U13204 (N_13204,N_11370,N_11369);
nor U13205 (N_13205,N_11270,N_11359);
nor U13206 (N_13206,N_11646,N_10734);
and U13207 (N_13207,N_11528,N_10801);
nand U13208 (N_13208,N_11746,N_10944);
or U13209 (N_13209,N_10688,N_11838);
and U13210 (N_13210,N_10584,N_10853);
and U13211 (N_13211,N_11291,N_11660);
nor U13212 (N_13212,N_11328,N_11197);
or U13213 (N_13213,N_11098,N_11924);
and U13214 (N_13214,N_10920,N_11939);
and U13215 (N_13215,N_11099,N_11058);
or U13216 (N_13216,N_11951,N_11513);
or U13217 (N_13217,N_11448,N_10891);
nand U13218 (N_13218,N_11757,N_11291);
or U13219 (N_13219,N_11857,N_11441);
xor U13220 (N_13220,N_11437,N_11117);
nand U13221 (N_13221,N_10748,N_11582);
xnor U13222 (N_13222,N_11117,N_11114);
or U13223 (N_13223,N_11593,N_11509);
nand U13224 (N_13224,N_11496,N_11101);
nor U13225 (N_13225,N_10955,N_10802);
and U13226 (N_13226,N_11672,N_10522);
and U13227 (N_13227,N_10742,N_10801);
and U13228 (N_13228,N_11501,N_10739);
or U13229 (N_13229,N_11919,N_11198);
nand U13230 (N_13230,N_11222,N_11889);
or U13231 (N_13231,N_11342,N_10941);
or U13232 (N_13232,N_11019,N_11039);
and U13233 (N_13233,N_11018,N_11767);
and U13234 (N_13234,N_11641,N_10501);
nor U13235 (N_13235,N_10737,N_10989);
nor U13236 (N_13236,N_11798,N_11164);
or U13237 (N_13237,N_11875,N_11130);
or U13238 (N_13238,N_11505,N_11927);
or U13239 (N_13239,N_10939,N_11019);
and U13240 (N_13240,N_10771,N_11620);
nor U13241 (N_13241,N_11402,N_10594);
or U13242 (N_13242,N_11333,N_10503);
nor U13243 (N_13243,N_11417,N_11149);
and U13244 (N_13244,N_11555,N_11365);
or U13245 (N_13245,N_11324,N_10653);
xnor U13246 (N_13246,N_11951,N_11598);
or U13247 (N_13247,N_11162,N_11753);
xor U13248 (N_13248,N_11040,N_11199);
nor U13249 (N_13249,N_11584,N_10626);
nor U13250 (N_13250,N_11233,N_10936);
nor U13251 (N_13251,N_11100,N_11999);
xnor U13252 (N_13252,N_11866,N_11177);
and U13253 (N_13253,N_11648,N_11995);
and U13254 (N_13254,N_11887,N_11121);
xnor U13255 (N_13255,N_11571,N_11843);
nor U13256 (N_13256,N_11375,N_11870);
nor U13257 (N_13257,N_11630,N_10939);
nor U13258 (N_13258,N_11578,N_10661);
nor U13259 (N_13259,N_10607,N_11771);
xor U13260 (N_13260,N_10806,N_10834);
xor U13261 (N_13261,N_10695,N_10910);
xor U13262 (N_13262,N_10641,N_10700);
or U13263 (N_13263,N_10605,N_10850);
or U13264 (N_13264,N_11810,N_11028);
or U13265 (N_13265,N_11268,N_11469);
or U13266 (N_13266,N_11980,N_10709);
xnor U13267 (N_13267,N_11439,N_10888);
nor U13268 (N_13268,N_11046,N_11898);
or U13269 (N_13269,N_10732,N_10570);
nor U13270 (N_13270,N_11846,N_10796);
nor U13271 (N_13271,N_10868,N_11228);
and U13272 (N_13272,N_11222,N_11377);
or U13273 (N_13273,N_11185,N_10630);
xor U13274 (N_13274,N_11419,N_10591);
nand U13275 (N_13275,N_11394,N_10526);
nand U13276 (N_13276,N_11314,N_11270);
nand U13277 (N_13277,N_10659,N_11404);
and U13278 (N_13278,N_10925,N_10874);
and U13279 (N_13279,N_11281,N_10704);
xor U13280 (N_13280,N_11981,N_11439);
nor U13281 (N_13281,N_11103,N_11755);
and U13282 (N_13282,N_11990,N_11443);
xnor U13283 (N_13283,N_11009,N_11612);
or U13284 (N_13284,N_11794,N_11064);
and U13285 (N_13285,N_11158,N_10982);
or U13286 (N_13286,N_11037,N_11353);
and U13287 (N_13287,N_11703,N_11738);
xor U13288 (N_13288,N_11603,N_11073);
xor U13289 (N_13289,N_11381,N_10972);
xor U13290 (N_13290,N_11838,N_10919);
nand U13291 (N_13291,N_11394,N_10749);
or U13292 (N_13292,N_11310,N_11682);
xnor U13293 (N_13293,N_11865,N_11630);
nor U13294 (N_13294,N_11464,N_10928);
or U13295 (N_13295,N_11516,N_11451);
and U13296 (N_13296,N_11056,N_11000);
and U13297 (N_13297,N_11546,N_10732);
or U13298 (N_13298,N_10877,N_10710);
nand U13299 (N_13299,N_10967,N_10853);
or U13300 (N_13300,N_11891,N_11929);
xor U13301 (N_13301,N_10850,N_10620);
nor U13302 (N_13302,N_10510,N_11893);
nor U13303 (N_13303,N_11814,N_10884);
nor U13304 (N_13304,N_11360,N_11334);
or U13305 (N_13305,N_11030,N_10898);
xnor U13306 (N_13306,N_10906,N_11478);
nor U13307 (N_13307,N_11485,N_10934);
or U13308 (N_13308,N_11602,N_10872);
or U13309 (N_13309,N_10657,N_10722);
and U13310 (N_13310,N_11211,N_10728);
nor U13311 (N_13311,N_11422,N_10735);
nand U13312 (N_13312,N_11450,N_11430);
or U13313 (N_13313,N_11306,N_11567);
nand U13314 (N_13314,N_11246,N_10521);
nor U13315 (N_13315,N_11440,N_10541);
xor U13316 (N_13316,N_10906,N_11908);
nand U13317 (N_13317,N_11440,N_11007);
xnor U13318 (N_13318,N_10703,N_11361);
and U13319 (N_13319,N_11198,N_11717);
or U13320 (N_13320,N_10528,N_11706);
or U13321 (N_13321,N_10534,N_11344);
nor U13322 (N_13322,N_11489,N_11684);
or U13323 (N_13323,N_11855,N_11087);
xor U13324 (N_13324,N_11445,N_10953);
and U13325 (N_13325,N_11715,N_11377);
nand U13326 (N_13326,N_11708,N_11230);
and U13327 (N_13327,N_10512,N_11423);
xor U13328 (N_13328,N_11575,N_11210);
xor U13329 (N_13329,N_11435,N_11068);
or U13330 (N_13330,N_11833,N_11504);
nand U13331 (N_13331,N_11086,N_11089);
nor U13332 (N_13332,N_10603,N_10574);
nor U13333 (N_13333,N_11398,N_11590);
xnor U13334 (N_13334,N_11208,N_11144);
and U13335 (N_13335,N_11423,N_11392);
nand U13336 (N_13336,N_11425,N_11469);
and U13337 (N_13337,N_11192,N_10563);
nor U13338 (N_13338,N_11426,N_10823);
or U13339 (N_13339,N_11314,N_11931);
nor U13340 (N_13340,N_11227,N_11813);
and U13341 (N_13341,N_10805,N_10626);
xnor U13342 (N_13342,N_10738,N_10822);
xor U13343 (N_13343,N_11743,N_10757);
xor U13344 (N_13344,N_11131,N_10555);
nor U13345 (N_13345,N_11205,N_11766);
xor U13346 (N_13346,N_11346,N_11122);
or U13347 (N_13347,N_11412,N_10757);
xnor U13348 (N_13348,N_10554,N_11660);
nand U13349 (N_13349,N_11454,N_11892);
nor U13350 (N_13350,N_10670,N_10975);
xor U13351 (N_13351,N_10705,N_10592);
nand U13352 (N_13352,N_11878,N_10719);
xor U13353 (N_13353,N_10847,N_11305);
and U13354 (N_13354,N_11781,N_10774);
nor U13355 (N_13355,N_10649,N_10681);
and U13356 (N_13356,N_10984,N_10945);
or U13357 (N_13357,N_11367,N_11738);
and U13358 (N_13358,N_11611,N_11912);
and U13359 (N_13359,N_11038,N_11751);
and U13360 (N_13360,N_10943,N_10875);
and U13361 (N_13361,N_10826,N_11179);
or U13362 (N_13362,N_11205,N_11214);
nor U13363 (N_13363,N_11969,N_10631);
and U13364 (N_13364,N_11282,N_11550);
nor U13365 (N_13365,N_11180,N_11139);
nor U13366 (N_13366,N_10868,N_11835);
nor U13367 (N_13367,N_11664,N_10857);
nand U13368 (N_13368,N_10840,N_11548);
nand U13369 (N_13369,N_10658,N_11014);
or U13370 (N_13370,N_11316,N_11425);
and U13371 (N_13371,N_11088,N_10612);
xnor U13372 (N_13372,N_11371,N_11158);
nor U13373 (N_13373,N_11909,N_11292);
or U13374 (N_13374,N_10808,N_10618);
and U13375 (N_13375,N_10981,N_11633);
nand U13376 (N_13376,N_10972,N_10892);
or U13377 (N_13377,N_11880,N_11662);
nor U13378 (N_13378,N_11442,N_11081);
or U13379 (N_13379,N_10553,N_10533);
xor U13380 (N_13380,N_11214,N_11620);
nand U13381 (N_13381,N_11640,N_11184);
and U13382 (N_13382,N_11018,N_10854);
or U13383 (N_13383,N_11703,N_11423);
nor U13384 (N_13384,N_11395,N_10824);
nand U13385 (N_13385,N_10791,N_10967);
or U13386 (N_13386,N_11052,N_10649);
or U13387 (N_13387,N_10774,N_11737);
or U13388 (N_13388,N_11704,N_10946);
and U13389 (N_13389,N_11818,N_11354);
nand U13390 (N_13390,N_11190,N_11018);
nor U13391 (N_13391,N_10750,N_11433);
nand U13392 (N_13392,N_11900,N_10863);
xnor U13393 (N_13393,N_11323,N_10675);
nor U13394 (N_13394,N_10678,N_11710);
nor U13395 (N_13395,N_10987,N_11739);
nor U13396 (N_13396,N_11642,N_11864);
xor U13397 (N_13397,N_11227,N_11798);
xnor U13398 (N_13398,N_10821,N_10973);
or U13399 (N_13399,N_11439,N_11899);
xnor U13400 (N_13400,N_10755,N_10726);
xnor U13401 (N_13401,N_11365,N_11320);
nor U13402 (N_13402,N_11098,N_10903);
nor U13403 (N_13403,N_10992,N_11772);
or U13404 (N_13404,N_11201,N_11447);
or U13405 (N_13405,N_10825,N_11718);
and U13406 (N_13406,N_11342,N_11319);
nand U13407 (N_13407,N_11823,N_10564);
xor U13408 (N_13408,N_11201,N_11582);
or U13409 (N_13409,N_11068,N_10900);
nor U13410 (N_13410,N_10880,N_10762);
and U13411 (N_13411,N_11362,N_11373);
xor U13412 (N_13412,N_10969,N_11652);
or U13413 (N_13413,N_11667,N_11871);
nand U13414 (N_13414,N_11612,N_11918);
and U13415 (N_13415,N_11839,N_11217);
xor U13416 (N_13416,N_10957,N_11412);
or U13417 (N_13417,N_10566,N_10666);
and U13418 (N_13418,N_11342,N_10919);
nand U13419 (N_13419,N_10738,N_10715);
nand U13420 (N_13420,N_11339,N_10658);
xor U13421 (N_13421,N_11606,N_11133);
xor U13422 (N_13422,N_11304,N_11676);
or U13423 (N_13423,N_10500,N_10992);
and U13424 (N_13424,N_11322,N_11275);
or U13425 (N_13425,N_11512,N_11413);
and U13426 (N_13426,N_10538,N_11568);
nand U13427 (N_13427,N_11446,N_11722);
or U13428 (N_13428,N_10993,N_11954);
or U13429 (N_13429,N_11582,N_10893);
and U13430 (N_13430,N_11023,N_11132);
nand U13431 (N_13431,N_11617,N_11547);
nand U13432 (N_13432,N_11522,N_11213);
nor U13433 (N_13433,N_11191,N_10581);
xnor U13434 (N_13434,N_11201,N_11655);
nand U13435 (N_13435,N_10649,N_10586);
nand U13436 (N_13436,N_10843,N_11063);
nor U13437 (N_13437,N_11187,N_11201);
nand U13438 (N_13438,N_11761,N_11525);
nand U13439 (N_13439,N_10656,N_10632);
nand U13440 (N_13440,N_10533,N_11737);
xnor U13441 (N_13441,N_11515,N_11733);
and U13442 (N_13442,N_11100,N_11479);
nor U13443 (N_13443,N_11330,N_10992);
and U13444 (N_13444,N_10884,N_10844);
nor U13445 (N_13445,N_11435,N_10506);
and U13446 (N_13446,N_11077,N_10512);
and U13447 (N_13447,N_11000,N_11652);
nor U13448 (N_13448,N_11699,N_11122);
nor U13449 (N_13449,N_11865,N_10553);
nand U13450 (N_13450,N_11765,N_11145);
nand U13451 (N_13451,N_11697,N_11514);
nor U13452 (N_13452,N_11937,N_10523);
and U13453 (N_13453,N_11196,N_11935);
xnor U13454 (N_13454,N_11504,N_11614);
xnor U13455 (N_13455,N_11368,N_11906);
nand U13456 (N_13456,N_11902,N_10670);
and U13457 (N_13457,N_11151,N_10630);
nor U13458 (N_13458,N_11461,N_10618);
and U13459 (N_13459,N_11340,N_10862);
nand U13460 (N_13460,N_11660,N_11779);
or U13461 (N_13461,N_11708,N_11977);
and U13462 (N_13462,N_10990,N_11850);
nor U13463 (N_13463,N_11938,N_11063);
nor U13464 (N_13464,N_11492,N_11264);
and U13465 (N_13465,N_11118,N_10984);
xnor U13466 (N_13466,N_11249,N_10592);
nand U13467 (N_13467,N_10999,N_11362);
xor U13468 (N_13468,N_10688,N_11270);
or U13469 (N_13469,N_11307,N_11861);
and U13470 (N_13470,N_10734,N_11337);
and U13471 (N_13471,N_10665,N_11724);
and U13472 (N_13472,N_11085,N_10782);
or U13473 (N_13473,N_10514,N_11782);
nor U13474 (N_13474,N_11107,N_11585);
or U13475 (N_13475,N_10750,N_10682);
xnor U13476 (N_13476,N_11730,N_11243);
or U13477 (N_13477,N_10795,N_11796);
nor U13478 (N_13478,N_10937,N_11387);
and U13479 (N_13479,N_11083,N_11196);
nand U13480 (N_13480,N_10959,N_11596);
or U13481 (N_13481,N_10963,N_11447);
nand U13482 (N_13482,N_10506,N_11553);
xnor U13483 (N_13483,N_11192,N_11103);
xnor U13484 (N_13484,N_10773,N_10837);
nand U13485 (N_13485,N_11479,N_10504);
nand U13486 (N_13486,N_10748,N_10523);
or U13487 (N_13487,N_10534,N_11067);
and U13488 (N_13488,N_10998,N_11304);
nand U13489 (N_13489,N_10541,N_10630);
nand U13490 (N_13490,N_11055,N_10867);
xor U13491 (N_13491,N_11746,N_11501);
and U13492 (N_13492,N_11105,N_11359);
or U13493 (N_13493,N_11573,N_11966);
nand U13494 (N_13494,N_10882,N_10648);
nand U13495 (N_13495,N_11053,N_11870);
nor U13496 (N_13496,N_11600,N_11097);
nand U13497 (N_13497,N_11879,N_11318);
or U13498 (N_13498,N_11693,N_10895);
xor U13499 (N_13499,N_10517,N_10871);
and U13500 (N_13500,N_12568,N_13112);
or U13501 (N_13501,N_12349,N_12981);
xnor U13502 (N_13502,N_13238,N_12551);
xor U13503 (N_13503,N_13225,N_12446);
or U13504 (N_13504,N_13377,N_12254);
xnor U13505 (N_13505,N_13263,N_12619);
nor U13506 (N_13506,N_12351,N_13142);
or U13507 (N_13507,N_13228,N_12628);
nor U13508 (N_13508,N_12313,N_13386);
nor U13509 (N_13509,N_12958,N_12176);
xnor U13510 (N_13510,N_13281,N_12122);
nand U13511 (N_13511,N_13250,N_13064);
and U13512 (N_13512,N_12260,N_13163);
or U13513 (N_13513,N_12144,N_12462);
xor U13514 (N_13514,N_13130,N_12866);
nor U13515 (N_13515,N_12851,N_13196);
xnor U13516 (N_13516,N_12782,N_13192);
and U13517 (N_13517,N_12787,N_13469);
nor U13518 (N_13518,N_12068,N_12956);
nand U13519 (N_13519,N_13014,N_12973);
nand U13520 (N_13520,N_12165,N_12448);
nor U13521 (N_13521,N_13448,N_13447);
nand U13522 (N_13522,N_13237,N_13091);
or U13523 (N_13523,N_13158,N_12198);
or U13524 (N_13524,N_13331,N_13017);
and U13525 (N_13525,N_12649,N_12560);
xnor U13526 (N_13526,N_12783,N_12997);
and U13527 (N_13527,N_12069,N_13026);
nor U13528 (N_13528,N_13231,N_13421);
nor U13529 (N_13529,N_12710,N_13495);
or U13530 (N_13530,N_12749,N_12250);
nor U13531 (N_13531,N_12368,N_12652);
xor U13532 (N_13532,N_12917,N_13122);
xnor U13533 (N_13533,N_13370,N_12631);
xnor U13534 (N_13534,N_12561,N_13292);
and U13535 (N_13535,N_12900,N_13369);
xor U13536 (N_13536,N_12110,N_13162);
nand U13537 (N_13537,N_12142,N_12959);
nand U13538 (N_13538,N_12440,N_12449);
nand U13539 (N_13539,N_12643,N_13305);
or U13540 (N_13540,N_12663,N_13407);
xor U13541 (N_13541,N_13352,N_13120);
xnor U13542 (N_13542,N_13145,N_12856);
and U13543 (N_13543,N_12739,N_12849);
and U13544 (N_13544,N_12056,N_12416);
xor U13545 (N_13545,N_12614,N_12211);
nor U13546 (N_13546,N_13279,N_12918);
xnor U13547 (N_13547,N_13126,N_13392);
and U13548 (N_13548,N_12057,N_12813);
nand U13549 (N_13549,N_12228,N_13188);
or U13550 (N_13550,N_12433,N_12341);
nand U13551 (N_13551,N_13310,N_13136);
nand U13552 (N_13552,N_12669,N_12378);
xor U13553 (N_13553,N_13390,N_12027);
or U13554 (N_13554,N_12659,N_12302);
and U13555 (N_13555,N_12232,N_12279);
xnor U13556 (N_13556,N_13182,N_13143);
or U13557 (N_13557,N_13243,N_12156);
or U13558 (N_13558,N_12885,N_12894);
nand U13559 (N_13559,N_12764,N_13488);
nand U13560 (N_13560,N_12342,N_13037);
or U13561 (N_13561,N_13436,N_12740);
or U13562 (N_13562,N_12453,N_13170);
or U13563 (N_13563,N_13131,N_12795);
xnor U13564 (N_13564,N_12274,N_12840);
nor U13565 (N_13565,N_13315,N_12486);
nand U13566 (N_13566,N_13052,N_12640);
or U13567 (N_13567,N_12184,N_12296);
nand U13568 (N_13568,N_13465,N_13150);
nand U13569 (N_13569,N_12412,N_12475);
or U13570 (N_13570,N_12968,N_12319);
xnor U13571 (N_13571,N_12479,N_12802);
nor U13572 (N_13572,N_12267,N_12678);
nor U13573 (N_13573,N_12510,N_12245);
or U13574 (N_13574,N_12213,N_12012);
or U13575 (N_13575,N_12294,N_12452);
xnor U13576 (N_13576,N_12556,N_12109);
nor U13577 (N_13577,N_12391,N_12707);
or U13578 (N_13578,N_13001,N_13341);
nand U13579 (N_13579,N_12099,N_13351);
xor U13580 (N_13580,N_12686,N_12424);
nand U13581 (N_13581,N_13372,N_12219);
xor U13582 (N_13582,N_12162,N_12426);
nand U13583 (N_13583,N_12158,N_13374);
xnor U13584 (N_13584,N_12089,N_12778);
or U13585 (N_13585,N_12550,N_12819);
xor U13586 (N_13586,N_12251,N_12916);
xnor U13587 (N_13587,N_13391,N_13245);
or U13588 (N_13588,N_13235,N_12687);
or U13589 (N_13589,N_12902,N_12011);
nand U13590 (N_13590,N_12494,N_13476);
and U13591 (N_13591,N_12932,N_12114);
or U13592 (N_13592,N_12582,N_12344);
and U13593 (N_13593,N_12645,N_12079);
and U13594 (N_13594,N_13334,N_13124);
nor U13595 (N_13595,N_12573,N_13173);
xor U13596 (N_13596,N_13206,N_12334);
xor U13597 (N_13597,N_12388,N_12415);
or U13598 (N_13598,N_12082,N_12854);
nor U13599 (N_13599,N_13306,N_13220);
nor U13600 (N_13600,N_12712,N_12464);
or U13601 (N_13601,N_13480,N_12681);
nor U13602 (N_13602,N_12199,N_13103);
nor U13603 (N_13603,N_12946,N_12549);
nand U13604 (N_13604,N_12193,N_12352);
nand U13605 (N_13605,N_12493,N_13467);
or U13606 (N_13606,N_12673,N_13239);
nand U13607 (N_13607,N_12656,N_12704);
nor U13608 (N_13608,N_13035,N_12421);
nand U13609 (N_13609,N_13267,N_12218);
and U13610 (N_13610,N_12090,N_13254);
xnor U13611 (N_13611,N_13345,N_12806);
and U13612 (N_13612,N_12272,N_12411);
nand U13613 (N_13613,N_12076,N_12935);
nor U13614 (N_13614,N_12390,N_12459);
or U13615 (N_13615,N_13474,N_13113);
nand U13616 (N_13616,N_13160,N_12034);
or U13617 (N_13617,N_12048,N_12238);
and U13618 (N_13618,N_12996,N_12280);
xnor U13619 (N_13619,N_12516,N_12719);
xor U13620 (N_13620,N_12197,N_12468);
and U13621 (N_13621,N_12519,N_13159);
or U13622 (N_13622,N_12853,N_12376);
or U13623 (N_13623,N_12419,N_12395);
nor U13624 (N_13624,N_13078,N_12485);
nor U13625 (N_13625,N_12999,N_12389);
nor U13626 (N_13626,N_12128,N_13289);
nand U13627 (N_13627,N_13384,N_12123);
xnor U13628 (N_13628,N_13032,N_13025);
or U13629 (N_13629,N_12767,N_13168);
or U13630 (N_13630,N_12898,N_12949);
nor U13631 (N_13631,N_12796,N_13083);
nand U13632 (N_13632,N_12742,N_13294);
and U13633 (N_13633,N_12666,N_12625);
or U13634 (N_13634,N_12350,N_12270);
nand U13635 (N_13635,N_13319,N_12192);
and U13636 (N_13636,N_13388,N_12558);
nand U13637 (N_13637,N_12063,N_13381);
and U13638 (N_13638,N_12658,N_13455);
or U13639 (N_13639,N_12538,N_12733);
or U13640 (N_13640,N_12758,N_12569);
nand U13641 (N_13641,N_12978,N_13011);
nand U13642 (N_13642,N_13435,N_12769);
nand U13643 (N_13643,N_12492,N_13401);
or U13644 (N_13644,N_12784,N_13146);
or U13645 (N_13645,N_12072,N_12848);
and U13646 (N_13646,N_12970,N_12400);
nor U13647 (N_13647,N_13321,N_12629);
and U13648 (N_13648,N_12869,N_12327);
nor U13649 (N_13649,N_13361,N_12566);
nand U13650 (N_13650,N_12333,N_12505);
and U13651 (N_13651,N_12682,N_13434);
and U13652 (N_13652,N_12330,N_13073);
or U13653 (N_13653,N_12170,N_12044);
or U13654 (N_13654,N_12471,N_13060);
and U13655 (N_13655,N_12445,N_12256);
xnor U13656 (N_13656,N_12525,N_12283);
nor U13657 (N_13657,N_13403,N_12222);
or U13658 (N_13658,N_12950,N_13333);
nand U13659 (N_13659,N_12896,N_12797);
nor U13660 (N_13660,N_13348,N_13007);
nor U13661 (N_13661,N_12358,N_12129);
xor U13662 (N_13662,N_12496,N_12096);
nand U13663 (N_13663,N_12227,N_12458);
or U13664 (N_13664,N_13338,N_12537);
or U13665 (N_13665,N_12071,N_13497);
nand U13666 (N_13666,N_13087,N_13471);
and U13667 (N_13667,N_12842,N_12820);
xnor U13668 (N_13668,N_13117,N_13302);
or U13669 (N_13669,N_12960,N_12595);
or U13670 (N_13670,N_12367,N_12974);
xor U13671 (N_13671,N_13227,N_13412);
or U13672 (N_13672,N_12600,N_13127);
xor U13673 (N_13673,N_13320,N_12230);
or U13674 (N_13674,N_12952,N_13489);
and U13675 (N_13675,N_12246,N_12859);
or U13676 (N_13676,N_12627,N_12506);
and U13677 (N_13677,N_13499,N_12661);
or U13678 (N_13678,N_13065,N_12321);
nand U13679 (N_13679,N_12613,N_12305);
nor U13680 (N_13680,N_13340,N_13493);
and U13681 (N_13681,N_12926,N_12530);
nand U13682 (N_13682,N_12830,N_12945);
nand U13683 (N_13683,N_13058,N_12407);
or U13684 (N_13684,N_12405,N_12861);
xnor U13685 (N_13685,N_13140,N_12638);
nor U13686 (N_13686,N_12857,N_12779);
nand U13687 (N_13687,N_13428,N_12382);
nor U13688 (N_13688,N_12759,N_12845);
or U13689 (N_13689,N_12356,N_12570);
xor U13690 (N_13690,N_12451,N_13194);
and U13691 (N_13691,N_12091,N_12683);
or U13692 (N_13692,N_12513,N_13347);
nor U13693 (N_13693,N_12244,N_13008);
and U13694 (N_13694,N_12284,N_12650);
or U13695 (N_13695,N_12237,N_12632);
or U13696 (N_13696,N_12157,N_12654);
xor U13697 (N_13697,N_13462,N_13062);
nand U13698 (N_13698,N_13230,N_12798);
nor U13699 (N_13699,N_12042,N_12689);
nor U13700 (N_13700,N_13234,N_12013);
xor U13701 (N_13701,N_13128,N_12312);
xnor U13702 (N_13702,N_12860,N_13191);
or U13703 (N_13703,N_12025,N_12140);
xnor U13704 (N_13704,N_13241,N_12488);
nor U13705 (N_13705,N_12756,N_12206);
and U13706 (N_13706,N_12065,N_13149);
nor U13707 (N_13707,N_13393,N_12169);
xor U13708 (N_13708,N_13287,N_12107);
nand U13709 (N_13709,N_12817,N_12024);
or U13710 (N_13710,N_12533,N_12168);
nor U13711 (N_13711,N_12092,N_13222);
xor U13712 (N_13712,N_12980,N_12924);
nor U13713 (N_13713,N_12546,N_12331);
nand U13714 (N_13714,N_12276,N_13077);
nand U13715 (N_13715,N_13186,N_12553);
and U13716 (N_13716,N_12088,N_12726);
nand U13717 (N_13717,N_12768,N_12810);
and U13718 (N_13718,N_12786,N_12508);
nand U13719 (N_13719,N_12354,N_13108);
nor U13720 (N_13720,N_12927,N_13203);
nor U13721 (N_13721,N_12723,N_13209);
or U13722 (N_13722,N_13045,N_12130);
nand U13723 (N_13723,N_12423,N_12383);
nand U13724 (N_13724,N_12921,N_13072);
nand U13725 (N_13725,N_12990,N_12290);
xor U13726 (N_13726,N_13041,N_13012);
nand U13727 (N_13727,N_12131,N_12816);
and U13728 (N_13728,N_12967,N_12149);
nand U13729 (N_13729,N_13270,N_12911);
nor U13730 (N_13730,N_12685,N_13244);
and U13731 (N_13731,N_12404,N_13354);
xor U13732 (N_13732,N_12439,N_12708);
nor U13733 (N_13733,N_12171,N_13490);
and U13734 (N_13734,N_12392,N_12146);
and U13735 (N_13735,N_12172,N_13094);
xor U13736 (N_13736,N_13223,N_12234);
nor U13737 (N_13737,N_12657,N_12429);
xor U13738 (N_13738,N_12035,N_12535);
nand U13739 (N_13739,N_12583,N_13387);
nor U13740 (N_13740,N_13139,N_13483);
nor U13741 (N_13741,N_13275,N_12434);
nor U13742 (N_13742,N_13180,N_12626);
nand U13743 (N_13743,N_12223,N_13208);
xor U13744 (N_13744,N_12040,N_13445);
xor U13745 (N_13745,N_12252,N_12067);
nor U13746 (N_13746,N_12509,N_12991);
nand U13747 (N_13747,N_12695,N_12907);
and U13748 (N_13748,N_13024,N_12744);
or U13749 (N_13749,N_13380,N_13290);
or U13750 (N_13750,N_12913,N_13213);
xnor U13751 (N_13751,N_12731,N_12037);
nor U13752 (N_13752,N_13383,N_13336);
nor U13753 (N_13753,N_12930,N_12258);
nand U13754 (N_13754,N_12292,N_12807);
or U13755 (N_13755,N_12752,N_12257);
and U13756 (N_13756,N_13265,N_12966);
nor U13757 (N_13757,N_12151,N_12671);
xnor U13758 (N_13758,N_12616,N_12147);
xnor U13759 (N_13759,N_12692,N_12381);
xnor U13760 (N_13760,N_12541,N_12502);
xor U13761 (N_13761,N_12191,N_12763);
or U13762 (N_13762,N_12125,N_12175);
and U13763 (N_13763,N_12112,N_13079);
nor U13764 (N_13764,N_12837,N_12348);
or U13765 (N_13765,N_13394,N_12922);
nand U13766 (N_13766,N_12877,N_12221);
or U13767 (N_13767,N_12635,N_12047);
nand U13768 (N_13768,N_12791,N_12548);
nor U13769 (N_13769,N_12514,N_12487);
and U13770 (N_13770,N_12982,N_12014);
or U13771 (N_13771,N_13258,N_12736);
xnor U13772 (N_13772,N_12021,N_12906);
nand U13773 (N_13773,N_12753,N_12004);
or U13774 (N_13774,N_13107,N_12755);
nand U13775 (N_13775,N_13408,N_12873);
nand U13776 (N_13776,N_12329,N_13324);
nor U13777 (N_13777,N_13433,N_12772);
or U13778 (N_13778,N_12827,N_13019);
nor U13779 (N_13779,N_12241,N_12714);
xnor U13780 (N_13780,N_12379,N_13304);
or U13781 (N_13781,N_12380,N_13458);
and U13782 (N_13782,N_13076,N_12512);
and U13783 (N_13783,N_12585,N_12402);
nand U13784 (N_13784,N_12983,N_12608);
xnor U13785 (N_13785,N_12346,N_12372);
nor U13786 (N_13786,N_12467,N_13397);
nor U13787 (N_13787,N_12792,N_12651);
xor U13788 (N_13788,N_12119,N_12361);
nand U13789 (N_13789,N_12594,N_12336);
or U13790 (N_13790,N_13312,N_13262);
nor U13791 (N_13791,N_12466,N_13111);
nor U13792 (N_13792,N_12846,N_12427);
or U13793 (N_13793,N_12443,N_13185);
nand U13794 (N_13794,N_12567,N_13311);
nand U13795 (N_13795,N_12882,N_13028);
nand U13796 (N_13796,N_12141,N_12915);
nand U13797 (N_13797,N_13473,N_12134);
or U13798 (N_13798,N_12403,N_12217);
and U13799 (N_13799,N_12364,N_13424);
nor U13800 (N_13800,N_13400,N_13399);
nand U13801 (N_13801,N_12442,N_13257);
and U13802 (N_13802,N_12291,N_12410);
xnor U13803 (N_13803,N_12912,N_12944);
nor U13804 (N_13804,N_13438,N_12295);
nand U13805 (N_13805,N_13382,N_12087);
nor U13806 (N_13806,N_12563,N_12043);
and U13807 (N_13807,N_13328,N_12006);
nand U13808 (N_13808,N_12064,N_12000);
and U13809 (N_13809,N_13410,N_13482);
and U13810 (N_13810,N_13085,N_12239);
or U13811 (N_13811,N_13439,N_12102);
nand U13812 (N_13812,N_12003,N_13043);
nand U13813 (N_13813,N_13119,N_12843);
xnor U13814 (N_13814,N_12660,N_12622);
nor U13815 (N_13815,N_12318,N_12463);
nor U13816 (N_13816,N_12016,N_13385);
nor U13817 (N_13817,N_12653,N_12053);
xnor U13818 (N_13818,N_13349,N_12871);
and U13819 (N_13819,N_13316,N_12889);
nor U13820 (N_13820,N_12891,N_12677);
nor U13821 (N_13821,N_12428,N_13088);
nor U13822 (N_13822,N_12397,N_13313);
or U13823 (N_13823,N_12437,N_12979);
and U13824 (N_13824,N_12115,N_13406);
nor U13825 (N_13825,N_12706,N_13039);
nor U13826 (N_13826,N_12822,N_12590);
nor U13827 (N_13827,N_12507,N_12201);
nor U13828 (N_13828,N_12621,N_12910);
and U13829 (N_13829,N_12240,N_12722);
or U13830 (N_13830,N_13441,N_12992);
nand U13831 (N_13831,N_12818,N_12435);
nand U13832 (N_13832,N_13066,N_12461);
nor U13833 (N_13833,N_13280,N_12059);
nor U13834 (N_13834,N_13189,N_12300);
xnor U13835 (N_13835,N_12738,N_12504);
xor U13836 (N_13836,N_12316,N_12668);
nor U13837 (N_13837,N_13426,N_12580);
or U13838 (N_13838,N_12143,N_12998);
nor U13839 (N_13839,N_12518,N_13100);
nor U13840 (N_13840,N_12282,N_12324);
nor U13841 (N_13841,N_13190,N_12465);
xnor U13842 (N_13842,N_12394,N_12278);
xnor U13843 (N_13843,N_12940,N_13022);
and U13844 (N_13844,N_12103,N_12699);
xor U13845 (N_13845,N_12852,N_12441);
nor U13846 (N_13846,N_12498,N_12747);
and U13847 (N_13847,N_12941,N_12696);
nor U13848 (N_13848,N_12483,N_13283);
or U13849 (N_13849,N_12094,N_12263);
nand U13850 (N_13850,N_13346,N_13456);
nand U13851 (N_13851,N_13200,N_12205);
nor U13852 (N_13852,N_12803,N_12994);
or U13853 (N_13853,N_12060,N_12371);
xnor U13854 (N_13854,N_12844,N_12760);
xnor U13855 (N_13855,N_12357,N_12933);
and U13856 (N_13856,N_12224,N_12478);
xor U13857 (N_13857,N_13004,N_13027);
and U13858 (N_13858,N_12167,N_12775);
nor U13859 (N_13859,N_12148,N_13003);
xnor U13860 (N_13860,N_12152,N_13307);
xor U13861 (N_13861,N_12189,N_12247);
and U13862 (N_13862,N_13260,N_12444);
xor U13863 (N_13863,N_13224,N_13494);
or U13864 (N_13864,N_13362,N_13296);
xor U13865 (N_13865,N_13102,N_12804);
and U13866 (N_13866,N_13266,N_12401);
nor U13867 (N_13867,N_12320,N_12592);
xor U13868 (N_13868,N_12317,N_12373);
or U13869 (N_13869,N_13242,N_12809);
xor U13870 (N_13870,N_12539,N_12709);
xnor U13871 (N_13871,N_13444,N_13031);
nand U13872 (N_13872,N_12482,N_12266);
or U13873 (N_13873,N_12249,N_12794);
nand U13874 (N_13874,N_13081,N_12269);
xnor U13875 (N_13875,N_12178,N_13147);
nand U13876 (N_13876,N_13365,N_13118);
and U13877 (N_13877,N_12557,N_12194);
nor U13878 (N_13878,N_13459,N_12919);
and U13879 (N_13879,N_13156,N_12049);
or U13880 (N_13880,N_12620,N_12624);
nor U13881 (N_13881,N_12363,N_12001);
nor U13882 (N_13882,N_12095,N_13057);
and U13883 (N_13883,N_13151,N_13165);
and U13884 (N_13884,N_12497,N_12936);
xnor U13885 (N_13885,N_12961,N_12957);
or U13886 (N_13886,N_12116,N_12417);
nor U13887 (N_13887,N_13212,N_13452);
nor U13888 (N_13888,N_12431,N_13472);
nor U13889 (N_13889,N_13099,N_12477);
or U13890 (N_13890,N_12185,N_12914);
nor U13891 (N_13891,N_13121,N_12879);
xnor U13892 (N_13892,N_12264,N_12026);
or U13893 (N_13893,N_12934,N_12552);
xor U13894 (N_13894,N_12457,N_13366);
nor U13895 (N_13895,N_12603,N_13233);
and U13896 (N_13896,N_12038,N_12534);
nor U13897 (N_13897,N_12664,N_12200);
and U13898 (N_13898,N_12823,N_12008);
xnor U13899 (N_13899,N_12186,N_12338);
and U13900 (N_13900,N_13277,N_13274);
nor U13901 (N_13901,N_12587,N_12559);
nor U13902 (N_13902,N_12489,N_13442);
and U13903 (N_13903,N_12301,N_12062);
xor U13904 (N_13904,N_13272,N_13269);
nand U13905 (N_13905,N_13398,N_13468);
xnor U13906 (N_13906,N_13067,N_12288);
nor U13907 (N_13907,N_13084,N_12623);
xor U13908 (N_13908,N_13479,N_12078);
nand U13909 (N_13909,N_13323,N_13418);
or U13910 (N_13910,N_13055,N_13429);
or U13911 (N_13911,N_12527,N_12811);
or U13912 (N_13912,N_12637,N_13049);
or U13913 (N_13913,N_13171,N_13175);
xnor U13914 (N_13914,N_12748,N_12897);
and U13915 (N_13915,N_12501,N_12225);
or U13916 (N_13916,N_12460,N_13236);
xor U13917 (N_13917,N_12883,N_13061);
and U13918 (N_13918,N_13309,N_13046);
xnor U13919 (N_13919,N_12515,N_12903);
or U13920 (N_13920,N_12299,N_12571);
nand U13921 (N_13921,N_12762,N_12310);
and U13922 (N_13922,N_12780,N_12536);
or U13923 (N_13923,N_12577,N_12886);
nand U13924 (N_13924,N_13042,N_12277);
xor U13925 (N_13925,N_12542,N_12868);
and U13926 (N_13926,N_13299,N_12727);
xor U13927 (N_13927,N_13148,N_13461);
or U13928 (N_13928,N_13216,N_12183);
and U13929 (N_13929,N_13261,N_12480);
xor U13930 (N_13930,N_12925,N_13367);
or U13931 (N_13931,N_13379,N_13376);
xor U13932 (N_13932,N_13314,N_12343);
nand U13933 (N_13933,N_12177,N_12304);
and U13934 (N_13934,N_13295,N_12135);
or U13935 (N_13935,N_13018,N_13110);
nand U13936 (N_13936,N_12523,N_12215);
nand U13937 (N_13937,N_12899,N_12281);
or U13938 (N_13938,N_12863,N_13359);
and U13939 (N_13939,N_13086,N_12589);
nand U13940 (N_13940,N_13104,N_12872);
xor U13941 (N_13941,N_12084,N_12406);
or U13942 (N_13942,N_12725,N_12540);
and U13943 (N_13943,N_12500,N_13353);
or U13944 (N_13944,N_13184,N_13330);
or U13945 (N_13945,N_12229,N_13034);
nand U13946 (N_13946,N_12097,N_12137);
nand U13947 (N_13947,N_13044,N_12297);
or U13948 (N_13948,N_13132,N_12839);
nand U13949 (N_13949,N_12881,N_12604);
xnor U13950 (N_13950,N_12605,N_12432);
nor U13951 (N_13951,N_13423,N_13286);
nor U13952 (N_13952,N_12473,N_12328);
and U13953 (N_13953,N_13422,N_12154);
or U13954 (N_13954,N_12150,N_12610);
and U13955 (N_13955,N_13470,N_12901);
or U13956 (N_13956,N_12161,N_13326);
nor U13957 (N_13957,N_12015,N_12120);
nand U13958 (N_13958,N_12684,N_13202);
and U13959 (N_13959,N_12989,N_12323);
or U13960 (N_13960,N_12133,N_12855);
nand U13961 (N_13961,N_13339,N_13069);
xnor U13962 (N_13962,N_12741,N_12781);
and U13963 (N_13963,N_13373,N_12833);
xnor U13964 (N_13964,N_12495,N_12572);
or U13965 (N_13965,N_12220,N_13443);
nor U13966 (N_13966,N_12750,N_12771);
xor U13967 (N_13967,N_13082,N_12208);
xor U13968 (N_13968,N_12598,N_13251);
nand U13969 (N_13969,N_12033,N_12895);
nor U13970 (N_13970,N_12963,N_12028);
or U13971 (N_13971,N_13360,N_13317);
and U13972 (N_13972,N_13015,N_13040);
or U13973 (N_13973,N_12720,N_13252);
nor U13974 (N_13974,N_13009,N_13463);
and U13975 (N_13975,N_13453,N_13288);
or U13976 (N_13976,N_12374,N_13451);
nand U13977 (N_13977,N_13181,N_13335);
or U13978 (N_13978,N_12179,N_12010);
and U13979 (N_13979,N_13054,N_13350);
and U13980 (N_13980,N_12526,N_13217);
nand U13981 (N_13981,N_12735,N_12667);
nor U13982 (N_13982,N_13343,N_12075);
nor U13983 (N_13983,N_12905,N_12607);
and U13984 (N_13984,N_13389,N_13464);
xnor U13985 (N_13985,N_12564,N_12884);
and U13986 (N_13986,N_13101,N_13106);
nor U13987 (N_13987,N_12522,N_13329);
and U13988 (N_13988,N_12204,N_13276);
and U13989 (N_13989,N_12606,N_12588);
xor U13990 (N_13990,N_13167,N_12369);
xor U13991 (N_13991,N_12335,N_12314);
or U13992 (N_13992,N_12009,N_12209);
and U13993 (N_13993,N_13172,N_12387);
nor U13994 (N_13994,N_13090,N_13415);
or U13995 (N_13995,N_12159,N_12073);
and U13996 (N_13996,N_13282,N_13249);
xor U13997 (N_13997,N_12155,N_12022);
xnor U13998 (N_13998,N_13116,N_12019);
nand U13999 (N_13999,N_12481,N_12639);
xnor U14000 (N_14000,N_12644,N_12948);
or U14001 (N_14001,N_13430,N_12132);
nand U14002 (N_14002,N_13268,N_12977);
nand U14003 (N_14003,N_12212,N_12825);
nand U14004 (N_14004,N_12986,N_12521);
or U14005 (N_14005,N_12100,N_12841);
or U14006 (N_14006,N_12337,N_12988);
xor U14007 (N_14007,N_12511,N_13138);
nor U14008 (N_14008,N_12174,N_12698);
and U14009 (N_14009,N_13300,N_12718);
or U14010 (N_14010,N_13070,N_12694);
and U14011 (N_14011,N_13195,N_13137);
nand U14012 (N_14012,N_12955,N_12824);
xor U14013 (N_14013,N_12243,N_13178);
or U14014 (N_14014,N_13036,N_12793);
or U14015 (N_14015,N_12020,N_12052);
xor U14016 (N_14016,N_12262,N_12565);
nor U14017 (N_14017,N_12746,N_12655);
nand U14018 (N_14018,N_12418,N_12216);
xnor U14019 (N_14019,N_12231,N_12145);
xor U14020 (N_14020,N_12413,N_12360);
xor U14021 (N_14021,N_13240,N_12286);
and U14022 (N_14022,N_12061,N_12826);
xor U14023 (N_14023,N_12838,N_13219);
and U14024 (N_14024,N_12705,N_12751);
xnor U14025 (N_14025,N_12408,N_12113);
or U14026 (N_14026,N_12578,N_12734);
and U14027 (N_14027,N_12581,N_13486);
xnor U14028 (N_14028,N_13485,N_12051);
nor U14029 (N_14029,N_13416,N_12646);
xor U14030 (N_14030,N_12636,N_13109);
or U14031 (N_14031,N_12285,N_12160);
nor U14032 (N_14032,N_12181,N_13183);
or U14033 (N_14033,N_12259,N_12951);
xor U14034 (N_14034,N_13030,N_13246);
or U14035 (N_14035,N_13154,N_12377);
nor U14036 (N_14036,N_13404,N_12969);
nand U14037 (N_14037,N_13000,N_12612);
nor U14038 (N_14038,N_12555,N_13141);
xor U14039 (N_14039,N_13431,N_12384);
or U14040 (N_14040,N_12287,N_12207);
and U14041 (N_14041,N_13068,N_12821);
and U14042 (N_14042,N_12831,N_13297);
nor U14043 (N_14043,N_12765,N_12662);
nor U14044 (N_14044,N_12080,N_12648);
nor U14045 (N_14045,N_12814,N_12834);
and U14046 (N_14046,N_12713,N_12942);
nor U14047 (N_14047,N_12688,N_12340);
and U14048 (N_14048,N_12964,N_13419);
or U14049 (N_14049,N_13050,N_12365);
or U14050 (N_14050,N_12490,N_13356);
nor U14051 (N_14051,N_12308,N_13358);
or U14052 (N_14052,N_12203,N_13023);
nor U14053 (N_14053,N_13215,N_12046);
nand U14054 (N_14054,N_13047,N_13092);
nor U14055 (N_14055,N_12469,N_12339);
xnor U14056 (N_14056,N_12503,N_12306);
or U14057 (N_14057,N_12584,N_13214);
nand U14058 (N_14058,N_13063,N_13002);
xor U14059 (N_14059,N_12325,N_12743);
and U14060 (N_14060,N_12943,N_12928);
or U14061 (N_14061,N_13013,N_12630);
and U14062 (N_14062,N_12430,N_13484);
xnor U14063 (N_14063,N_12332,N_12265);
nand U14064 (N_14064,N_12562,N_12456);
nand U14065 (N_14065,N_13293,N_13477);
or U14066 (N_14066,N_12665,N_12790);
nand U14067 (N_14067,N_12828,N_12393);
or U14068 (N_14068,N_12976,N_13135);
nor U14069 (N_14069,N_13021,N_12138);
nand U14070 (N_14070,N_13048,N_13395);
xnor U14071 (N_14071,N_12018,N_12529);
nor U14072 (N_14072,N_13020,N_12773);
and U14073 (N_14073,N_12633,N_13440);
nand U14074 (N_14074,N_13198,N_12680);
and U14075 (N_14075,N_12732,N_13371);
nor U14076 (N_14076,N_12770,N_12691);
and U14077 (N_14077,N_12058,N_12180);
and U14078 (N_14078,N_13177,N_13357);
xnor U14079 (N_14079,N_13375,N_12436);
nand U14080 (N_14080,N_12386,N_13327);
xor U14081 (N_14081,N_12472,N_12615);
nor U14082 (N_14082,N_13207,N_12920);
and U14083 (N_14083,N_13278,N_12908);
xnor U14084 (N_14084,N_13457,N_13475);
and U14085 (N_14085,N_12359,N_12531);
nand U14086 (N_14086,N_13285,N_12850);
nor U14087 (N_14087,N_13187,N_12066);
or U14088 (N_14088,N_12166,N_12326);
xnor U14089 (N_14089,N_12106,N_12375);
or U14090 (N_14090,N_12596,N_12353);
and U14091 (N_14091,N_13402,N_12788);
nor U14092 (N_14092,N_12880,N_12450);
and U14093 (N_14093,N_13125,N_12962);
nor U14094 (N_14094,N_12757,N_12422);
or U14095 (N_14095,N_12345,N_12878);
xnor U14096 (N_14096,N_13204,N_12586);
or U14097 (N_14097,N_13318,N_12030);
and U14098 (N_14098,N_12904,N_13332);
nand U14099 (N_14099,N_13115,N_12995);
nand U14100 (N_14100,N_12947,N_12799);
nand U14101 (N_14101,N_13256,N_13096);
xnor U14102 (N_14102,N_13420,N_13449);
xor U14103 (N_14103,N_12690,N_12108);
or U14104 (N_14104,N_12124,N_12055);
nand U14105 (N_14105,N_12214,N_12355);
or U14106 (N_14106,N_12937,N_12528);
or U14107 (N_14107,N_12591,N_12647);
xor U14108 (N_14108,N_12093,N_12864);
xor U14109 (N_14109,N_13291,N_12847);
nor U14110 (N_14110,N_12036,N_12697);
and U14111 (N_14111,N_12987,N_12261);
or U14112 (N_14112,N_13271,N_12023);
or U14113 (N_14113,N_12579,N_12425);
nor U14114 (N_14114,N_13425,N_12307);
nor U14115 (N_14115,N_12777,N_12985);
or U14116 (N_14116,N_12311,N_13259);
and U14117 (N_14117,N_13437,N_12597);
nand U14118 (N_14118,N_12737,N_13221);
xnor U14119 (N_14119,N_13364,N_12104);
nand U14120 (N_14120,N_12273,N_12599);
nor U14121 (N_14121,N_12729,N_12776);
xor U14122 (N_14122,N_12724,N_12275);
nor U14123 (N_14123,N_12474,N_13450);
xnor U14124 (N_14124,N_12255,N_13264);
and U14125 (N_14125,N_13414,N_12785);
or U14126 (N_14126,N_12870,N_12164);
or U14127 (N_14127,N_13089,N_12153);
nor U14128 (N_14128,N_13161,N_13129);
or U14129 (N_14129,N_12532,N_12975);
xor U14130 (N_14130,N_13226,N_12173);
and U14131 (N_14131,N_12953,N_12118);
nand U14132 (N_14132,N_13051,N_12865);
or U14133 (N_14133,N_12196,N_12017);
nor U14134 (N_14134,N_13409,N_13355);
or U14135 (N_14135,N_12370,N_12032);
or U14136 (N_14136,N_12543,N_13201);
nand U14137 (N_14137,N_13053,N_13255);
nor U14138 (N_14138,N_12309,N_13303);
and U14139 (N_14139,N_12805,N_12676);
or U14140 (N_14140,N_12235,N_12139);
or U14141 (N_14141,N_12182,N_12575);
or U14142 (N_14142,N_13133,N_12576);
and U14143 (N_14143,N_13193,N_12298);
or U14144 (N_14144,N_12002,N_12163);
or U14145 (N_14145,N_13174,N_13197);
xnor U14146 (N_14146,N_13413,N_13460);
nand U14147 (N_14147,N_12126,N_12909);
nor U14148 (N_14148,N_13247,N_12693);
or U14149 (N_14149,N_12385,N_12835);
or U14150 (N_14150,N_12862,N_13157);
nor U14151 (N_14151,N_13166,N_12874);
nand U14152 (N_14152,N_13169,N_12923);
nor U14153 (N_14153,N_13071,N_12438);
nand U14154 (N_14154,N_12041,N_13095);
nor U14155 (N_14155,N_12700,N_12618);
and U14156 (N_14156,N_12081,N_12812);
nand U14157 (N_14157,N_12702,N_13498);
xor U14158 (N_14158,N_12892,N_12289);
nor U14159 (N_14159,N_12858,N_12031);
and U14160 (N_14160,N_13337,N_13308);
xnor U14161 (N_14161,N_13097,N_13033);
or U14162 (N_14162,N_12054,N_12226);
and U14163 (N_14163,N_13016,N_12554);
and U14164 (N_14164,N_12679,N_12045);
nand U14165 (N_14165,N_12674,N_13164);
nor U14166 (N_14166,N_12602,N_12520);
or U14167 (N_14167,N_12236,N_12611);
and U14168 (N_14168,N_13005,N_12398);
nor U14169 (N_14169,N_13378,N_12268);
or U14170 (N_14170,N_13273,N_13123);
nor U14171 (N_14171,N_13481,N_12761);
nand U14172 (N_14172,N_13176,N_12829);
nand U14173 (N_14173,N_12233,N_12347);
nand U14174 (N_14174,N_12366,N_12085);
xnor U14175 (N_14175,N_12789,N_12101);
and U14176 (N_14176,N_13229,N_12086);
and U14177 (N_14177,N_12188,N_12029);
and U14178 (N_14178,N_12454,N_12938);
or U14179 (N_14179,N_13152,N_13487);
or U14180 (N_14180,N_12074,N_12253);
and U14181 (N_14181,N_12717,N_12491);
nor U14182 (N_14182,N_12642,N_13080);
xor U14183 (N_14183,N_12774,N_12547);
and U14184 (N_14184,N_13074,N_13284);
and U14185 (N_14185,N_13363,N_12005);
nor U14186 (N_14186,N_12574,N_12832);
xnor U14187 (N_14187,N_13478,N_12121);
xnor U14188 (N_14188,N_12721,N_12815);
nor U14189 (N_14189,N_12271,N_13417);
or U14190 (N_14190,N_12609,N_12715);
xnor U14191 (N_14191,N_13232,N_13344);
xor U14192 (N_14192,N_12202,N_12670);
nor U14193 (N_14193,N_12800,N_13205);
or U14194 (N_14194,N_12455,N_13342);
or U14195 (N_14195,N_12362,N_12954);
nand U14196 (N_14196,N_12315,N_13432);
nor U14197 (N_14197,N_12887,N_12544);
nand U14198 (N_14198,N_12641,N_13093);
nor U14199 (N_14199,N_12524,N_13006);
nand U14200 (N_14200,N_12470,N_13155);
nor U14201 (N_14201,N_13218,N_12077);
or U14202 (N_14202,N_12195,N_12414);
nand U14203 (N_14203,N_13427,N_12888);
and U14204 (N_14204,N_13322,N_12293);
xnor U14205 (N_14205,N_12409,N_13029);
xnor U14206 (N_14206,N_13114,N_13059);
nand U14207 (N_14207,N_12931,N_12711);
or U14208 (N_14208,N_12476,N_13496);
xnor U14209 (N_14209,N_12396,N_12322);
xor U14210 (N_14210,N_12875,N_12893);
and U14211 (N_14211,N_13466,N_12447);
nor U14212 (N_14212,N_13098,N_12801);
or U14213 (N_14213,N_12187,N_12070);
nor U14214 (N_14214,N_12716,N_12420);
or U14215 (N_14215,N_12730,N_13454);
nand U14216 (N_14216,N_12617,N_12111);
nand U14217 (N_14217,N_13144,N_12965);
nor U14218 (N_14218,N_12929,N_12303);
xnor U14219 (N_14219,N_13038,N_13253);
xnor U14220 (N_14220,N_12971,N_12210);
xor U14221 (N_14221,N_12593,N_12754);
or U14222 (N_14222,N_12039,N_13368);
or U14223 (N_14223,N_12867,N_12939);
or U14224 (N_14224,N_13325,N_12672);
nor U14225 (N_14225,N_13075,N_13056);
nand U14226 (N_14226,N_12190,N_12972);
nor U14227 (N_14227,N_13491,N_13396);
nand U14228 (N_14228,N_13199,N_12098);
and U14229 (N_14229,N_13492,N_13153);
nand U14230 (N_14230,N_12399,N_12242);
and U14231 (N_14231,N_13411,N_12675);
and U14232 (N_14232,N_12136,N_13134);
nor U14233 (N_14233,N_12984,N_12601);
and U14234 (N_14234,N_13211,N_12007);
and U14235 (N_14235,N_12808,N_12484);
nor U14236 (N_14236,N_12745,N_12876);
nor U14237 (N_14237,N_12545,N_13179);
nor U14238 (N_14238,N_12703,N_12127);
xor U14239 (N_14239,N_12517,N_13301);
and U14240 (N_14240,N_13298,N_13010);
nor U14241 (N_14241,N_13248,N_13405);
xor U14242 (N_14242,N_12890,N_13105);
and U14243 (N_14243,N_12728,N_12083);
nor U14244 (N_14244,N_12248,N_12105);
nor U14245 (N_14245,N_12766,N_13446);
and U14246 (N_14246,N_12634,N_12701);
or U14247 (N_14247,N_12050,N_12836);
or U14248 (N_14248,N_12499,N_13210);
or U14249 (N_14249,N_12117,N_12993);
or U14250 (N_14250,N_12583,N_13498);
xor U14251 (N_14251,N_12333,N_12727);
or U14252 (N_14252,N_13346,N_12840);
xnor U14253 (N_14253,N_12047,N_12531);
nor U14254 (N_14254,N_13325,N_12631);
xnor U14255 (N_14255,N_12943,N_13148);
nor U14256 (N_14256,N_12125,N_12336);
or U14257 (N_14257,N_12623,N_12082);
nor U14258 (N_14258,N_13019,N_12115);
or U14259 (N_14259,N_12230,N_12982);
and U14260 (N_14260,N_13399,N_12919);
nand U14261 (N_14261,N_13210,N_12578);
or U14262 (N_14262,N_12862,N_12411);
nor U14263 (N_14263,N_13428,N_12065);
nor U14264 (N_14264,N_13246,N_13423);
nor U14265 (N_14265,N_12877,N_12323);
nor U14266 (N_14266,N_13333,N_13169);
and U14267 (N_14267,N_12296,N_13190);
and U14268 (N_14268,N_13291,N_12045);
nor U14269 (N_14269,N_12126,N_12251);
xor U14270 (N_14270,N_12506,N_13086);
nor U14271 (N_14271,N_12640,N_12414);
nor U14272 (N_14272,N_13438,N_12066);
nor U14273 (N_14273,N_12520,N_12576);
xnor U14274 (N_14274,N_12374,N_13109);
nor U14275 (N_14275,N_12448,N_12494);
xnor U14276 (N_14276,N_13424,N_12673);
nor U14277 (N_14277,N_12744,N_12778);
or U14278 (N_14278,N_12527,N_12275);
and U14279 (N_14279,N_12709,N_13365);
nor U14280 (N_14280,N_12464,N_12575);
nor U14281 (N_14281,N_12092,N_13325);
nand U14282 (N_14282,N_13442,N_12802);
xor U14283 (N_14283,N_12641,N_12146);
or U14284 (N_14284,N_12064,N_13121);
nand U14285 (N_14285,N_12172,N_12202);
and U14286 (N_14286,N_12790,N_13432);
nor U14287 (N_14287,N_12735,N_13050);
and U14288 (N_14288,N_12788,N_13447);
and U14289 (N_14289,N_12108,N_12455);
and U14290 (N_14290,N_13429,N_12786);
nor U14291 (N_14291,N_12177,N_12027);
and U14292 (N_14292,N_13422,N_12780);
and U14293 (N_14293,N_12319,N_12975);
nand U14294 (N_14294,N_12997,N_13458);
and U14295 (N_14295,N_12442,N_13365);
or U14296 (N_14296,N_12901,N_12259);
or U14297 (N_14297,N_12310,N_13265);
and U14298 (N_14298,N_13120,N_13330);
and U14299 (N_14299,N_12637,N_12927);
xnor U14300 (N_14300,N_12850,N_12933);
nor U14301 (N_14301,N_12626,N_13430);
xor U14302 (N_14302,N_12148,N_12326);
xnor U14303 (N_14303,N_12425,N_12907);
nor U14304 (N_14304,N_12116,N_13465);
or U14305 (N_14305,N_12572,N_12897);
or U14306 (N_14306,N_12250,N_13196);
nand U14307 (N_14307,N_12858,N_12223);
xor U14308 (N_14308,N_13088,N_12211);
or U14309 (N_14309,N_12166,N_12190);
and U14310 (N_14310,N_12394,N_12374);
xor U14311 (N_14311,N_13217,N_13078);
and U14312 (N_14312,N_12464,N_12416);
nand U14313 (N_14313,N_12485,N_12775);
or U14314 (N_14314,N_12316,N_13310);
nor U14315 (N_14315,N_13238,N_12791);
and U14316 (N_14316,N_12058,N_12694);
or U14317 (N_14317,N_12477,N_12276);
xor U14318 (N_14318,N_13067,N_12065);
nand U14319 (N_14319,N_13462,N_12977);
or U14320 (N_14320,N_12039,N_12965);
nor U14321 (N_14321,N_13024,N_12021);
xor U14322 (N_14322,N_12119,N_12586);
nand U14323 (N_14323,N_12525,N_13404);
nand U14324 (N_14324,N_12906,N_13072);
and U14325 (N_14325,N_12851,N_12052);
nor U14326 (N_14326,N_12325,N_13295);
or U14327 (N_14327,N_13390,N_12500);
nor U14328 (N_14328,N_12591,N_12197);
nand U14329 (N_14329,N_12529,N_12866);
nor U14330 (N_14330,N_12884,N_12409);
or U14331 (N_14331,N_13221,N_12834);
nor U14332 (N_14332,N_12342,N_13101);
xor U14333 (N_14333,N_12857,N_12515);
nor U14334 (N_14334,N_12487,N_12947);
nor U14335 (N_14335,N_12161,N_12984);
nand U14336 (N_14336,N_13235,N_13246);
and U14337 (N_14337,N_12867,N_13072);
xor U14338 (N_14338,N_13008,N_12598);
nand U14339 (N_14339,N_13485,N_12886);
nand U14340 (N_14340,N_12737,N_12741);
xnor U14341 (N_14341,N_13181,N_12840);
xor U14342 (N_14342,N_12047,N_12096);
nand U14343 (N_14343,N_13409,N_12188);
or U14344 (N_14344,N_12873,N_13357);
nand U14345 (N_14345,N_12109,N_12504);
and U14346 (N_14346,N_13079,N_12782);
xnor U14347 (N_14347,N_13331,N_13410);
xor U14348 (N_14348,N_13168,N_12421);
xor U14349 (N_14349,N_12762,N_12319);
nand U14350 (N_14350,N_13109,N_12331);
and U14351 (N_14351,N_12891,N_12906);
and U14352 (N_14352,N_12780,N_13192);
or U14353 (N_14353,N_13417,N_12890);
and U14354 (N_14354,N_13221,N_12971);
nor U14355 (N_14355,N_12542,N_13462);
xor U14356 (N_14356,N_13274,N_12369);
or U14357 (N_14357,N_12795,N_12826);
nand U14358 (N_14358,N_12301,N_12174);
xnor U14359 (N_14359,N_12150,N_13205);
or U14360 (N_14360,N_12702,N_12819);
or U14361 (N_14361,N_12948,N_12327);
or U14362 (N_14362,N_13152,N_13139);
xnor U14363 (N_14363,N_13415,N_12563);
or U14364 (N_14364,N_12584,N_12929);
nand U14365 (N_14365,N_12956,N_12440);
and U14366 (N_14366,N_13492,N_12666);
nor U14367 (N_14367,N_12795,N_12841);
and U14368 (N_14368,N_12987,N_12433);
xor U14369 (N_14369,N_13257,N_12808);
xor U14370 (N_14370,N_12588,N_12417);
or U14371 (N_14371,N_13376,N_12582);
nand U14372 (N_14372,N_12937,N_12861);
xnor U14373 (N_14373,N_12834,N_12648);
xnor U14374 (N_14374,N_13389,N_12109);
or U14375 (N_14375,N_12226,N_13170);
or U14376 (N_14376,N_12546,N_12704);
and U14377 (N_14377,N_12771,N_12673);
nand U14378 (N_14378,N_12720,N_13095);
or U14379 (N_14379,N_13007,N_13167);
nor U14380 (N_14380,N_13198,N_12352);
nand U14381 (N_14381,N_13001,N_12161);
nor U14382 (N_14382,N_12370,N_12393);
or U14383 (N_14383,N_12643,N_12620);
nor U14384 (N_14384,N_12425,N_13311);
or U14385 (N_14385,N_12126,N_12372);
and U14386 (N_14386,N_12007,N_12694);
nor U14387 (N_14387,N_12529,N_12563);
nor U14388 (N_14388,N_13368,N_13191);
xor U14389 (N_14389,N_13329,N_13010);
xnor U14390 (N_14390,N_12809,N_12985);
and U14391 (N_14391,N_12837,N_13498);
and U14392 (N_14392,N_12210,N_12446);
nand U14393 (N_14393,N_12775,N_12968);
xor U14394 (N_14394,N_12477,N_13103);
and U14395 (N_14395,N_12997,N_13457);
or U14396 (N_14396,N_12609,N_12143);
nand U14397 (N_14397,N_12128,N_12216);
nor U14398 (N_14398,N_13296,N_13202);
or U14399 (N_14399,N_12156,N_12894);
and U14400 (N_14400,N_12282,N_12767);
nand U14401 (N_14401,N_12464,N_12972);
xor U14402 (N_14402,N_12471,N_12902);
nor U14403 (N_14403,N_12507,N_13367);
nor U14404 (N_14404,N_12585,N_12555);
and U14405 (N_14405,N_12497,N_12666);
xnor U14406 (N_14406,N_12970,N_12265);
or U14407 (N_14407,N_12617,N_12496);
nand U14408 (N_14408,N_12418,N_12072);
and U14409 (N_14409,N_13440,N_12662);
nand U14410 (N_14410,N_13182,N_13151);
nand U14411 (N_14411,N_13013,N_13166);
and U14412 (N_14412,N_12533,N_12365);
or U14413 (N_14413,N_12103,N_13309);
or U14414 (N_14414,N_13472,N_12045);
nand U14415 (N_14415,N_13213,N_12168);
nand U14416 (N_14416,N_12601,N_13285);
and U14417 (N_14417,N_12224,N_13323);
nor U14418 (N_14418,N_12545,N_13256);
or U14419 (N_14419,N_12057,N_13156);
and U14420 (N_14420,N_12914,N_13189);
nand U14421 (N_14421,N_13013,N_12480);
nor U14422 (N_14422,N_12204,N_13032);
or U14423 (N_14423,N_12224,N_13340);
nand U14424 (N_14424,N_12847,N_12017);
xor U14425 (N_14425,N_12660,N_12381);
nand U14426 (N_14426,N_12839,N_12931);
xor U14427 (N_14427,N_12444,N_13466);
xnor U14428 (N_14428,N_12151,N_12617);
or U14429 (N_14429,N_12851,N_12372);
nand U14430 (N_14430,N_12043,N_12762);
nand U14431 (N_14431,N_13479,N_13420);
or U14432 (N_14432,N_13328,N_12732);
nor U14433 (N_14433,N_12713,N_13405);
and U14434 (N_14434,N_13322,N_13292);
nand U14435 (N_14435,N_12505,N_12892);
or U14436 (N_14436,N_12713,N_12699);
nor U14437 (N_14437,N_12418,N_12011);
nor U14438 (N_14438,N_12722,N_12458);
or U14439 (N_14439,N_12229,N_12625);
or U14440 (N_14440,N_12733,N_12764);
and U14441 (N_14441,N_13050,N_12781);
xnor U14442 (N_14442,N_12819,N_12976);
nor U14443 (N_14443,N_13396,N_13114);
xor U14444 (N_14444,N_13295,N_13050);
nand U14445 (N_14445,N_12501,N_12451);
and U14446 (N_14446,N_12558,N_12753);
nand U14447 (N_14447,N_12275,N_13428);
and U14448 (N_14448,N_12144,N_12521);
nor U14449 (N_14449,N_12403,N_12200);
or U14450 (N_14450,N_12917,N_12809);
or U14451 (N_14451,N_12464,N_12832);
and U14452 (N_14452,N_13009,N_13364);
nor U14453 (N_14453,N_12066,N_12291);
nor U14454 (N_14454,N_13318,N_13048);
nor U14455 (N_14455,N_13411,N_13374);
or U14456 (N_14456,N_13118,N_12704);
or U14457 (N_14457,N_12630,N_12165);
or U14458 (N_14458,N_12491,N_12565);
xnor U14459 (N_14459,N_13188,N_12523);
and U14460 (N_14460,N_13144,N_13252);
xnor U14461 (N_14461,N_13337,N_13029);
xnor U14462 (N_14462,N_12414,N_12968);
xor U14463 (N_14463,N_12463,N_12524);
and U14464 (N_14464,N_12286,N_13494);
nor U14465 (N_14465,N_12858,N_12221);
xor U14466 (N_14466,N_12135,N_12942);
or U14467 (N_14467,N_13112,N_12208);
nand U14468 (N_14468,N_13219,N_13201);
and U14469 (N_14469,N_13488,N_12083);
or U14470 (N_14470,N_13467,N_13230);
or U14471 (N_14471,N_13498,N_12386);
and U14472 (N_14472,N_12655,N_12449);
xnor U14473 (N_14473,N_12623,N_13354);
nand U14474 (N_14474,N_12036,N_12493);
or U14475 (N_14475,N_12724,N_13043);
xnor U14476 (N_14476,N_12991,N_12507);
nor U14477 (N_14477,N_12442,N_12873);
nand U14478 (N_14478,N_12644,N_12884);
xor U14479 (N_14479,N_12213,N_13039);
nor U14480 (N_14480,N_12775,N_12572);
nand U14481 (N_14481,N_12161,N_13126);
xor U14482 (N_14482,N_12165,N_12810);
nor U14483 (N_14483,N_12586,N_12495);
or U14484 (N_14484,N_12447,N_12592);
or U14485 (N_14485,N_12066,N_12688);
nor U14486 (N_14486,N_12704,N_12592);
and U14487 (N_14487,N_12362,N_12191);
and U14488 (N_14488,N_12994,N_12936);
nand U14489 (N_14489,N_13382,N_12749);
nand U14490 (N_14490,N_13240,N_12080);
xor U14491 (N_14491,N_12343,N_12949);
nor U14492 (N_14492,N_13048,N_12279);
nor U14493 (N_14493,N_13275,N_13173);
nor U14494 (N_14494,N_13455,N_13350);
nand U14495 (N_14495,N_12600,N_12831);
or U14496 (N_14496,N_13490,N_12883);
or U14497 (N_14497,N_13228,N_13385);
or U14498 (N_14498,N_13057,N_13386);
nor U14499 (N_14499,N_12078,N_12476);
nor U14500 (N_14500,N_12664,N_12957);
nor U14501 (N_14501,N_12862,N_13438);
or U14502 (N_14502,N_12555,N_12982);
xor U14503 (N_14503,N_12927,N_12684);
xor U14504 (N_14504,N_13450,N_12920);
and U14505 (N_14505,N_12243,N_12132);
nand U14506 (N_14506,N_12923,N_12592);
nor U14507 (N_14507,N_12250,N_13423);
and U14508 (N_14508,N_12895,N_12532);
or U14509 (N_14509,N_12656,N_13067);
nand U14510 (N_14510,N_12243,N_12002);
nor U14511 (N_14511,N_12024,N_12468);
and U14512 (N_14512,N_13056,N_13447);
nand U14513 (N_14513,N_12140,N_12220);
nand U14514 (N_14514,N_12126,N_12322);
or U14515 (N_14515,N_12460,N_12398);
nor U14516 (N_14516,N_12819,N_12937);
and U14517 (N_14517,N_13407,N_12096);
nand U14518 (N_14518,N_12241,N_12202);
nor U14519 (N_14519,N_12336,N_12320);
nand U14520 (N_14520,N_13479,N_12985);
nand U14521 (N_14521,N_12738,N_12191);
or U14522 (N_14522,N_12031,N_13250);
and U14523 (N_14523,N_12229,N_12325);
nor U14524 (N_14524,N_12150,N_13126);
or U14525 (N_14525,N_12334,N_12309);
nand U14526 (N_14526,N_12113,N_12825);
xnor U14527 (N_14527,N_12725,N_12498);
nor U14528 (N_14528,N_12554,N_12756);
xnor U14529 (N_14529,N_13055,N_13438);
xor U14530 (N_14530,N_12142,N_12992);
and U14531 (N_14531,N_12845,N_12453);
or U14532 (N_14532,N_12765,N_13179);
nand U14533 (N_14533,N_13337,N_12120);
nand U14534 (N_14534,N_13130,N_13194);
xnor U14535 (N_14535,N_12315,N_12299);
nor U14536 (N_14536,N_12352,N_13333);
or U14537 (N_14537,N_12851,N_12261);
xor U14538 (N_14538,N_12683,N_13293);
nor U14539 (N_14539,N_12911,N_13477);
or U14540 (N_14540,N_12613,N_12553);
and U14541 (N_14541,N_13240,N_13301);
or U14542 (N_14542,N_12755,N_12560);
nor U14543 (N_14543,N_12181,N_13289);
and U14544 (N_14544,N_12713,N_12939);
and U14545 (N_14545,N_13418,N_13288);
xnor U14546 (N_14546,N_12496,N_13215);
xor U14547 (N_14547,N_12472,N_12060);
xor U14548 (N_14548,N_12286,N_12759);
xor U14549 (N_14549,N_13107,N_13118);
xnor U14550 (N_14550,N_13002,N_12949);
nor U14551 (N_14551,N_13418,N_12962);
nor U14552 (N_14552,N_12984,N_12330);
and U14553 (N_14553,N_13381,N_12125);
or U14554 (N_14554,N_13070,N_13476);
nand U14555 (N_14555,N_13335,N_12817);
nor U14556 (N_14556,N_12638,N_13363);
nand U14557 (N_14557,N_13048,N_12615);
nor U14558 (N_14558,N_13216,N_12666);
or U14559 (N_14559,N_13443,N_12021);
or U14560 (N_14560,N_13281,N_12406);
nand U14561 (N_14561,N_12982,N_12647);
nor U14562 (N_14562,N_12922,N_12879);
nor U14563 (N_14563,N_13016,N_12385);
nor U14564 (N_14564,N_12842,N_13477);
nor U14565 (N_14565,N_12322,N_12758);
xnor U14566 (N_14566,N_13259,N_13417);
and U14567 (N_14567,N_12716,N_12805);
nor U14568 (N_14568,N_12303,N_12791);
nand U14569 (N_14569,N_12199,N_12111);
nor U14570 (N_14570,N_12170,N_13007);
and U14571 (N_14571,N_12847,N_13056);
nand U14572 (N_14572,N_12753,N_13348);
nor U14573 (N_14573,N_12407,N_13445);
or U14574 (N_14574,N_12488,N_13094);
nor U14575 (N_14575,N_12862,N_12833);
xor U14576 (N_14576,N_12512,N_13241);
xnor U14577 (N_14577,N_12002,N_12142);
xor U14578 (N_14578,N_12323,N_13103);
nor U14579 (N_14579,N_12012,N_13222);
or U14580 (N_14580,N_13305,N_12506);
nand U14581 (N_14581,N_12740,N_12891);
or U14582 (N_14582,N_13348,N_13274);
xnor U14583 (N_14583,N_13037,N_12630);
and U14584 (N_14584,N_12807,N_12795);
nand U14585 (N_14585,N_13266,N_12005);
or U14586 (N_14586,N_12026,N_13095);
xnor U14587 (N_14587,N_12376,N_12594);
xnor U14588 (N_14588,N_12497,N_13181);
and U14589 (N_14589,N_12511,N_13114);
and U14590 (N_14590,N_12805,N_12115);
nor U14591 (N_14591,N_13418,N_13318);
nor U14592 (N_14592,N_12313,N_12130);
xnor U14593 (N_14593,N_12828,N_13453);
xnor U14594 (N_14594,N_12839,N_12115);
xnor U14595 (N_14595,N_12615,N_12448);
and U14596 (N_14596,N_12014,N_13438);
nand U14597 (N_14597,N_12113,N_13294);
nand U14598 (N_14598,N_12139,N_12069);
nor U14599 (N_14599,N_13313,N_13437);
or U14600 (N_14600,N_12301,N_12462);
xor U14601 (N_14601,N_12403,N_12409);
and U14602 (N_14602,N_13422,N_12615);
nor U14603 (N_14603,N_13408,N_12836);
xnor U14604 (N_14604,N_12693,N_12279);
nor U14605 (N_14605,N_12313,N_12012);
nor U14606 (N_14606,N_13471,N_13100);
and U14607 (N_14607,N_13056,N_13352);
and U14608 (N_14608,N_13274,N_12577);
nor U14609 (N_14609,N_13043,N_13223);
nor U14610 (N_14610,N_13011,N_13269);
and U14611 (N_14611,N_12848,N_12462);
xor U14612 (N_14612,N_13010,N_12975);
and U14613 (N_14613,N_12208,N_12241);
or U14614 (N_14614,N_12181,N_13276);
or U14615 (N_14615,N_13420,N_12207);
nor U14616 (N_14616,N_12790,N_12616);
or U14617 (N_14617,N_12607,N_12009);
and U14618 (N_14618,N_12836,N_12577);
xnor U14619 (N_14619,N_13453,N_12509);
and U14620 (N_14620,N_12445,N_12748);
or U14621 (N_14621,N_12409,N_13120);
nor U14622 (N_14622,N_12244,N_12583);
nor U14623 (N_14623,N_13441,N_13235);
xnor U14624 (N_14624,N_12985,N_12459);
nand U14625 (N_14625,N_12001,N_12313);
and U14626 (N_14626,N_12048,N_12338);
nor U14627 (N_14627,N_12243,N_12507);
or U14628 (N_14628,N_12761,N_12937);
and U14629 (N_14629,N_13079,N_12904);
and U14630 (N_14630,N_12128,N_12136);
nand U14631 (N_14631,N_12027,N_12403);
nor U14632 (N_14632,N_12187,N_12557);
xor U14633 (N_14633,N_12771,N_12328);
nand U14634 (N_14634,N_12650,N_12025);
nand U14635 (N_14635,N_13063,N_13478);
and U14636 (N_14636,N_12894,N_13154);
nand U14637 (N_14637,N_13280,N_12434);
or U14638 (N_14638,N_13468,N_12983);
and U14639 (N_14639,N_13248,N_13318);
or U14640 (N_14640,N_13064,N_12648);
xnor U14641 (N_14641,N_12905,N_12884);
and U14642 (N_14642,N_13097,N_13133);
xor U14643 (N_14643,N_12403,N_12657);
and U14644 (N_14644,N_12969,N_12215);
nand U14645 (N_14645,N_12775,N_12044);
nand U14646 (N_14646,N_12543,N_12941);
or U14647 (N_14647,N_12533,N_12339);
nor U14648 (N_14648,N_12529,N_12232);
and U14649 (N_14649,N_13478,N_13076);
or U14650 (N_14650,N_12882,N_12348);
nand U14651 (N_14651,N_12093,N_12666);
nor U14652 (N_14652,N_12664,N_12101);
and U14653 (N_14653,N_12972,N_12819);
nor U14654 (N_14654,N_13023,N_12673);
xor U14655 (N_14655,N_13233,N_12398);
nor U14656 (N_14656,N_12925,N_12496);
and U14657 (N_14657,N_13090,N_12386);
and U14658 (N_14658,N_13402,N_12885);
or U14659 (N_14659,N_12565,N_12479);
and U14660 (N_14660,N_13185,N_12482);
nand U14661 (N_14661,N_12861,N_13300);
nor U14662 (N_14662,N_12362,N_13400);
nor U14663 (N_14663,N_12882,N_12871);
xor U14664 (N_14664,N_12037,N_12992);
nand U14665 (N_14665,N_13297,N_13250);
xor U14666 (N_14666,N_13435,N_12807);
or U14667 (N_14667,N_13410,N_12937);
xor U14668 (N_14668,N_12069,N_12576);
nor U14669 (N_14669,N_12571,N_13321);
or U14670 (N_14670,N_13201,N_12867);
nor U14671 (N_14671,N_12312,N_13198);
nand U14672 (N_14672,N_13197,N_12615);
or U14673 (N_14673,N_12237,N_12191);
or U14674 (N_14674,N_13336,N_12028);
nor U14675 (N_14675,N_12319,N_13335);
and U14676 (N_14676,N_12514,N_12815);
and U14677 (N_14677,N_12498,N_12536);
or U14678 (N_14678,N_12921,N_12860);
and U14679 (N_14679,N_13460,N_12791);
nor U14680 (N_14680,N_13472,N_12336);
nor U14681 (N_14681,N_12118,N_12404);
or U14682 (N_14682,N_12044,N_13150);
or U14683 (N_14683,N_12504,N_12062);
nand U14684 (N_14684,N_12942,N_12206);
and U14685 (N_14685,N_12087,N_13414);
xor U14686 (N_14686,N_12371,N_13021);
xor U14687 (N_14687,N_12063,N_13386);
nand U14688 (N_14688,N_12150,N_13306);
xor U14689 (N_14689,N_12084,N_13047);
or U14690 (N_14690,N_12862,N_12106);
nor U14691 (N_14691,N_12477,N_12619);
and U14692 (N_14692,N_12718,N_12428);
nor U14693 (N_14693,N_13438,N_13159);
xor U14694 (N_14694,N_12651,N_12136);
nor U14695 (N_14695,N_12706,N_12985);
nand U14696 (N_14696,N_12103,N_13073);
xnor U14697 (N_14697,N_12073,N_13107);
nor U14698 (N_14698,N_12705,N_12935);
xor U14699 (N_14699,N_13368,N_12534);
nand U14700 (N_14700,N_12024,N_12987);
nor U14701 (N_14701,N_12913,N_12251);
or U14702 (N_14702,N_12427,N_13023);
nand U14703 (N_14703,N_12610,N_13260);
and U14704 (N_14704,N_13064,N_12453);
nand U14705 (N_14705,N_13292,N_12616);
and U14706 (N_14706,N_13472,N_12216);
nor U14707 (N_14707,N_12902,N_12579);
nand U14708 (N_14708,N_13481,N_12126);
nor U14709 (N_14709,N_12662,N_13340);
and U14710 (N_14710,N_13338,N_12617);
or U14711 (N_14711,N_13251,N_13355);
and U14712 (N_14712,N_12892,N_12357);
and U14713 (N_14713,N_12714,N_12438);
and U14714 (N_14714,N_12177,N_13181);
nor U14715 (N_14715,N_12465,N_12942);
or U14716 (N_14716,N_13016,N_13480);
nand U14717 (N_14717,N_12548,N_12155);
and U14718 (N_14718,N_12830,N_12549);
and U14719 (N_14719,N_12360,N_13114);
and U14720 (N_14720,N_12648,N_12624);
nand U14721 (N_14721,N_12022,N_12451);
nand U14722 (N_14722,N_12438,N_12380);
nand U14723 (N_14723,N_12071,N_12859);
and U14724 (N_14724,N_12612,N_13255);
and U14725 (N_14725,N_12471,N_12589);
nand U14726 (N_14726,N_12175,N_13054);
nand U14727 (N_14727,N_13232,N_12145);
or U14728 (N_14728,N_12329,N_13292);
and U14729 (N_14729,N_13382,N_13130);
and U14730 (N_14730,N_12318,N_12415);
xor U14731 (N_14731,N_12699,N_12790);
nor U14732 (N_14732,N_13444,N_12036);
nand U14733 (N_14733,N_13330,N_12228);
or U14734 (N_14734,N_12756,N_12743);
nor U14735 (N_14735,N_12983,N_13329);
or U14736 (N_14736,N_12315,N_12435);
nand U14737 (N_14737,N_12352,N_12271);
xnor U14738 (N_14738,N_12483,N_13201);
nand U14739 (N_14739,N_12210,N_12398);
xor U14740 (N_14740,N_13085,N_12616);
nor U14741 (N_14741,N_12803,N_12272);
and U14742 (N_14742,N_13250,N_12345);
nand U14743 (N_14743,N_13119,N_12239);
xnor U14744 (N_14744,N_12288,N_13330);
nand U14745 (N_14745,N_12257,N_13344);
nand U14746 (N_14746,N_12534,N_13082);
and U14747 (N_14747,N_13325,N_12097);
nand U14748 (N_14748,N_13480,N_13179);
nand U14749 (N_14749,N_12360,N_12938);
or U14750 (N_14750,N_12683,N_12205);
and U14751 (N_14751,N_12632,N_12922);
or U14752 (N_14752,N_13014,N_12468);
or U14753 (N_14753,N_12152,N_12407);
xor U14754 (N_14754,N_12526,N_13135);
and U14755 (N_14755,N_12122,N_13247);
or U14756 (N_14756,N_12122,N_12635);
xnor U14757 (N_14757,N_12487,N_13498);
and U14758 (N_14758,N_12514,N_13000);
nand U14759 (N_14759,N_13326,N_12416);
and U14760 (N_14760,N_13140,N_13180);
nand U14761 (N_14761,N_12495,N_12144);
or U14762 (N_14762,N_12351,N_13393);
nand U14763 (N_14763,N_12764,N_13174);
xnor U14764 (N_14764,N_13111,N_12150);
or U14765 (N_14765,N_12702,N_13318);
xor U14766 (N_14766,N_13329,N_12796);
xor U14767 (N_14767,N_12299,N_13495);
nand U14768 (N_14768,N_12565,N_12514);
nand U14769 (N_14769,N_12387,N_12750);
or U14770 (N_14770,N_12778,N_12801);
or U14771 (N_14771,N_12179,N_12079);
nand U14772 (N_14772,N_12079,N_12744);
nor U14773 (N_14773,N_12971,N_13056);
or U14774 (N_14774,N_12099,N_12221);
nand U14775 (N_14775,N_12551,N_12830);
nand U14776 (N_14776,N_13343,N_12471);
or U14777 (N_14777,N_13284,N_12535);
xnor U14778 (N_14778,N_12166,N_12574);
xnor U14779 (N_14779,N_12708,N_12736);
xnor U14780 (N_14780,N_12567,N_13383);
xnor U14781 (N_14781,N_12339,N_12216);
xnor U14782 (N_14782,N_12410,N_12203);
xnor U14783 (N_14783,N_13464,N_12817);
nand U14784 (N_14784,N_12918,N_12245);
or U14785 (N_14785,N_12287,N_12883);
and U14786 (N_14786,N_12222,N_12246);
nor U14787 (N_14787,N_13087,N_12413);
or U14788 (N_14788,N_12079,N_13190);
nor U14789 (N_14789,N_12594,N_12240);
nand U14790 (N_14790,N_12540,N_12386);
xnor U14791 (N_14791,N_13362,N_13038);
xnor U14792 (N_14792,N_13412,N_12068);
xor U14793 (N_14793,N_13487,N_12258);
and U14794 (N_14794,N_12604,N_13361);
and U14795 (N_14795,N_12804,N_12234);
or U14796 (N_14796,N_12436,N_12772);
and U14797 (N_14797,N_13006,N_13122);
nor U14798 (N_14798,N_13401,N_12487);
or U14799 (N_14799,N_13309,N_12487);
and U14800 (N_14800,N_12238,N_12533);
nand U14801 (N_14801,N_12760,N_12051);
or U14802 (N_14802,N_13251,N_12324);
nand U14803 (N_14803,N_13384,N_12193);
and U14804 (N_14804,N_12715,N_12622);
or U14805 (N_14805,N_12465,N_12047);
or U14806 (N_14806,N_12353,N_12332);
and U14807 (N_14807,N_12302,N_13072);
and U14808 (N_14808,N_12971,N_13349);
or U14809 (N_14809,N_12534,N_12114);
or U14810 (N_14810,N_13085,N_12700);
xnor U14811 (N_14811,N_13041,N_12542);
or U14812 (N_14812,N_12275,N_13172);
nand U14813 (N_14813,N_13446,N_13218);
nor U14814 (N_14814,N_12415,N_12549);
or U14815 (N_14815,N_12366,N_12242);
and U14816 (N_14816,N_13308,N_12547);
nor U14817 (N_14817,N_13192,N_12546);
nand U14818 (N_14818,N_12973,N_12883);
nor U14819 (N_14819,N_12072,N_12029);
and U14820 (N_14820,N_12468,N_12998);
xor U14821 (N_14821,N_13053,N_13456);
and U14822 (N_14822,N_13493,N_12923);
xnor U14823 (N_14823,N_13468,N_13397);
nor U14824 (N_14824,N_12128,N_12399);
and U14825 (N_14825,N_12649,N_12885);
nand U14826 (N_14826,N_13192,N_13467);
xor U14827 (N_14827,N_12976,N_13422);
xor U14828 (N_14828,N_12300,N_12041);
and U14829 (N_14829,N_12798,N_12901);
and U14830 (N_14830,N_13438,N_12914);
nor U14831 (N_14831,N_13112,N_12367);
nand U14832 (N_14832,N_12581,N_12411);
xnor U14833 (N_14833,N_12752,N_13038);
and U14834 (N_14834,N_12430,N_12523);
and U14835 (N_14835,N_13018,N_12838);
nand U14836 (N_14836,N_13223,N_12958);
or U14837 (N_14837,N_12341,N_12371);
nor U14838 (N_14838,N_13002,N_12479);
nor U14839 (N_14839,N_12000,N_12486);
nor U14840 (N_14840,N_12699,N_12042);
and U14841 (N_14841,N_12668,N_13044);
and U14842 (N_14842,N_13080,N_13419);
nor U14843 (N_14843,N_12714,N_13095);
nor U14844 (N_14844,N_12731,N_12098);
or U14845 (N_14845,N_13454,N_13342);
xnor U14846 (N_14846,N_12199,N_12012);
and U14847 (N_14847,N_13335,N_13079);
or U14848 (N_14848,N_13229,N_12933);
xnor U14849 (N_14849,N_12644,N_12466);
nor U14850 (N_14850,N_12531,N_12981);
xor U14851 (N_14851,N_12208,N_13353);
xnor U14852 (N_14852,N_12065,N_12380);
and U14853 (N_14853,N_13180,N_12805);
nand U14854 (N_14854,N_12098,N_13399);
nor U14855 (N_14855,N_12536,N_12261);
or U14856 (N_14856,N_12747,N_12935);
or U14857 (N_14857,N_13097,N_13438);
xor U14858 (N_14858,N_12198,N_13360);
xor U14859 (N_14859,N_13157,N_13333);
nand U14860 (N_14860,N_13218,N_12740);
nand U14861 (N_14861,N_12465,N_12149);
nor U14862 (N_14862,N_12847,N_13251);
xor U14863 (N_14863,N_12070,N_13350);
nor U14864 (N_14864,N_12380,N_12078);
xnor U14865 (N_14865,N_12457,N_12589);
nor U14866 (N_14866,N_12290,N_12138);
or U14867 (N_14867,N_13221,N_12649);
or U14868 (N_14868,N_13479,N_12502);
nor U14869 (N_14869,N_12365,N_12358);
and U14870 (N_14870,N_13066,N_13458);
xnor U14871 (N_14871,N_12608,N_12530);
nand U14872 (N_14872,N_12723,N_12045);
nand U14873 (N_14873,N_13401,N_12156);
or U14874 (N_14874,N_12314,N_12133);
nand U14875 (N_14875,N_13303,N_12870);
nand U14876 (N_14876,N_13090,N_12832);
xnor U14877 (N_14877,N_12904,N_12807);
or U14878 (N_14878,N_13220,N_13153);
xnor U14879 (N_14879,N_12556,N_12684);
nor U14880 (N_14880,N_12271,N_13068);
nand U14881 (N_14881,N_13262,N_12037);
nand U14882 (N_14882,N_12748,N_12280);
nor U14883 (N_14883,N_12680,N_13018);
nand U14884 (N_14884,N_12848,N_12104);
nand U14885 (N_14885,N_12368,N_12308);
nor U14886 (N_14886,N_12165,N_13482);
xnor U14887 (N_14887,N_12036,N_13236);
xnor U14888 (N_14888,N_12873,N_12248);
or U14889 (N_14889,N_12577,N_12746);
nand U14890 (N_14890,N_12653,N_12014);
nand U14891 (N_14891,N_12569,N_12621);
nor U14892 (N_14892,N_13329,N_13267);
and U14893 (N_14893,N_13208,N_12593);
xor U14894 (N_14894,N_13224,N_12946);
or U14895 (N_14895,N_12469,N_13388);
xor U14896 (N_14896,N_12054,N_12995);
and U14897 (N_14897,N_12008,N_13286);
and U14898 (N_14898,N_13060,N_13070);
and U14899 (N_14899,N_12267,N_13116);
or U14900 (N_14900,N_12162,N_12298);
nand U14901 (N_14901,N_12648,N_13458);
nor U14902 (N_14902,N_12343,N_12786);
and U14903 (N_14903,N_12165,N_12665);
nand U14904 (N_14904,N_12896,N_12785);
and U14905 (N_14905,N_12570,N_12816);
xnor U14906 (N_14906,N_13374,N_13348);
and U14907 (N_14907,N_13167,N_12370);
nor U14908 (N_14908,N_13084,N_12501);
nand U14909 (N_14909,N_12137,N_12551);
or U14910 (N_14910,N_12272,N_12670);
and U14911 (N_14911,N_12621,N_12299);
or U14912 (N_14912,N_13331,N_12403);
nand U14913 (N_14913,N_12130,N_12903);
or U14914 (N_14914,N_13230,N_12149);
nor U14915 (N_14915,N_12674,N_12782);
or U14916 (N_14916,N_13165,N_12741);
xnor U14917 (N_14917,N_12979,N_12082);
or U14918 (N_14918,N_12684,N_13174);
or U14919 (N_14919,N_12852,N_13346);
nor U14920 (N_14920,N_12986,N_12943);
and U14921 (N_14921,N_12823,N_12747);
or U14922 (N_14922,N_12947,N_12568);
nand U14923 (N_14923,N_13046,N_12517);
nor U14924 (N_14924,N_13195,N_12013);
and U14925 (N_14925,N_12917,N_12901);
or U14926 (N_14926,N_12294,N_12500);
nor U14927 (N_14927,N_12602,N_13289);
nor U14928 (N_14928,N_12599,N_12553);
xor U14929 (N_14929,N_13403,N_12056);
and U14930 (N_14930,N_12064,N_12185);
and U14931 (N_14931,N_13325,N_12613);
xnor U14932 (N_14932,N_13449,N_13100);
or U14933 (N_14933,N_13202,N_12062);
nor U14934 (N_14934,N_12858,N_12046);
nor U14935 (N_14935,N_12605,N_13102);
nand U14936 (N_14936,N_13392,N_12254);
nand U14937 (N_14937,N_13052,N_12055);
nand U14938 (N_14938,N_13163,N_12033);
nand U14939 (N_14939,N_12586,N_12377);
nor U14940 (N_14940,N_12510,N_12756);
xnor U14941 (N_14941,N_12075,N_13311);
xor U14942 (N_14942,N_12857,N_13029);
or U14943 (N_14943,N_13024,N_13102);
nor U14944 (N_14944,N_12416,N_12289);
nor U14945 (N_14945,N_12651,N_12156);
xnor U14946 (N_14946,N_12192,N_12844);
nor U14947 (N_14947,N_12247,N_12883);
or U14948 (N_14948,N_12436,N_12646);
or U14949 (N_14949,N_12161,N_12751);
nand U14950 (N_14950,N_12728,N_13074);
and U14951 (N_14951,N_12645,N_13154);
xnor U14952 (N_14952,N_12969,N_12329);
nor U14953 (N_14953,N_12717,N_12671);
or U14954 (N_14954,N_12002,N_12050);
nand U14955 (N_14955,N_13071,N_12116);
nand U14956 (N_14956,N_12064,N_12240);
and U14957 (N_14957,N_12553,N_12336);
nand U14958 (N_14958,N_13199,N_12575);
nand U14959 (N_14959,N_12918,N_13320);
xor U14960 (N_14960,N_12970,N_13064);
or U14961 (N_14961,N_12641,N_13010);
nand U14962 (N_14962,N_13412,N_12898);
xnor U14963 (N_14963,N_13167,N_13054);
or U14964 (N_14964,N_13410,N_12228);
or U14965 (N_14965,N_13418,N_13498);
nor U14966 (N_14966,N_13398,N_12919);
or U14967 (N_14967,N_12827,N_12145);
nor U14968 (N_14968,N_13175,N_12250);
or U14969 (N_14969,N_12680,N_13073);
xor U14970 (N_14970,N_12252,N_13186);
nor U14971 (N_14971,N_12008,N_13140);
or U14972 (N_14972,N_12566,N_13175);
xnor U14973 (N_14973,N_13373,N_12378);
or U14974 (N_14974,N_13149,N_13490);
nor U14975 (N_14975,N_13074,N_12511);
and U14976 (N_14976,N_13326,N_13484);
and U14977 (N_14977,N_13009,N_13076);
or U14978 (N_14978,N_12214,N_12595);
and U14979 (N_14979,N_13328,N_12715);
nand U14980 (N_14980,N_12929,N_13079);
or U14981 (N_14981,N_12523,N_12957);
nand U14982 (N_14982,N_12713,N_12149);
nor U14983 (N_14983,N_12138,N_13382);
nor U14984 (N_14984,N_12202,N_13048);
xnor U14985 (N_14985,N_13339,N_13387);
nor U14986 (N_14986,N_12999,N_12292);
or U14987 (N_14987,N_13397,N_13495);
and U14988 (N_14988,N_12561,N_12996);
nor U14989 (N_14989,N_13038,N_12136);
or U14990 (N_14990,N_12121,N_12887);
or U14991 (N_14991,N_12789,N_12823);
xor U14992 (N_14992,N_13081,N_13080);
or U14993 (N_14993,N_12842,N_12442);
nor U14994 (N_14994,N_12635,N_12940);
or U14995 (N_14995,N_13079,N_12504);
or U14996 (N_14996,N_12450,N_13126);
nor U14997 (N_14997,N_13016,N_12786);
nor U14998 (N_14998,N_13432,N_13451);
or U14999 (N_14999,N_12265,N_12956);
or U15000 (N_15000,N_14386,N_14896);
xnor U15001 (N_15001,N_14757,N_13539);
nand U15002 (N_15002,N_14216,N_13690);
xor U15003 (N_15003,N_14658,N_14233);
xor U15004 (N_15004,N_14945,N_13932);
or U15005 (N_15005,N_14287,N_14929);
nor U15006 (N_15006,N_14560,N_14306);
or U15007 (N_15007,N_14220,N_14048);
and U15008 (N_15008,N_13514,N_13988);
nor U15009 (N_15009,N_14650,N_14343);
or U15010 (N_15010,N_14175,N_14406);
xor U15011 (N_15011,N_14036,N_13583);
or U15012 (N_15012,N_14813,N_13635);
nand U15013 (N_15013,N_14814,N_13885);
nor U15014 (N_15014,N_13937,N_13557);
and U15015 (N_15015,N_13941,N_14689);
and U15016 (N_15016,N_14897,N_14071);
or U15017 (N_15017,N_13553,N_14482);
and U15018 (N_15018,N_13567,N_13964);
nand U15019 (N_15019,N_14179,N_14640);
or U15020 (N_15020,N_13748,N_13864);
and U15021 (N_15021,N_14189,N_14960);
nand U15022 (N_15022,N_14285,N_14350);
nor U15023 (N_15023,N_14054,N_14344);
or U15024 (N_15024,N_14114,N_14671);
or U15025 (N_15025,N_14496,N_14020);
nand U15026 (N_15026,N_14201,N_14436);
and U15027 (N_15027,N_14367,N_14052);
or U15028 (N_15028,N_13700,N_13596);
or U15029 (N_15029,N_14852,N_13966);
and U15030 (N_15030,N_14511,N_13836);
nor U15031 (N_15031,N_13907,N_14889);
xnor U15032 (N_15032,N_14510,N_14737);
xnor U15033 (N_15033,N_14474,N_13906);
xnor U15034 (N_15034,N_13779,N_14764);
nor U15035 (N_15035,N_14796,N_13564);
and U15036 (N_15036,N_13617,N_14383);
xor U15037 (N_15037,N_14711,N_14027);
nand U15038 (N_15038,N_13793,N_14248);
xor U15039 (N_15039,N_14636,N_14774);
nor U15040 (N_15040,N_13780,N_13684);
nand U15041 (N_15041,N_14789,N_13840);
nor U15042 (N_15042,N_14720,N_13512);
nand U15043 (N_15043,N_14151,N_14275);
or U15044 (N_15044,N_14728,N_14610);
nand U15045 (N_15045,N_14604,N_13650);
xnor U15046 (N_15046,N_14058,N_14932);
and U15047 (N_15047,N_13537,N_14663);
xor U15048 (N_15048,N_14319,N_14881);
nand U15049 (N_15049,N_13696,N_14119);
nand U15050 (N_15050,N_14688,N_14615);
xnor U15051 (N_15051,N_14296,N_13558);
and U15052 (N_15052,N_13532,N_14212);
or U15053 (N_15053,N_14846,N_13633);
xnor U15054 (N_15054,N_14930,N_14417);
or U15055 (N_15055,N_14270,N_14762);
or U15056 (N_15056,N_13587,N_14241);
or U15057 (N_15057,N_14810,N_13620);
nor U15058 (N_15058,N_13657,N_13502);
nor U15059 (N_15059,N_13627,N_14756);
xor U15060 (N_15060,N_14817,N_14237);
xnor U15061 (N_15061,N_14418,N_13586);
or U15062 (N_15062,N_13654,N_14706);
or U15063 (N_15063,N_14811,N_14642);
xor U15064 (N_15064,N_14007,N_14371);
or U15065 (N_15065,N_13738,N_14668);
nor U15066 (N_15066,N_13822,N_14978);
or U15067 (N_15067,N_14594,N_14529);
xnor U15068 (N_15068,N_14264,N_14825);
nor U15069 (N_15069,N_13718,N_14521);
xor U15070 (N_15070,N_14578,N_14065);
xnor U15071 (N_15071,N_14907,N_14605);
xnor U15072 (N_15072,N_13943,N_14533);
and U15073 (N_15073,N_13601,N_14039);
nand U15074 (N_15074,N_14991,N_13781);
nor U15075 (N_15075,N_14623,N_14758);
nor U15076 (N_15076,N_13820,N_14106);
or U15077 (N_15077,N_14419,N_14550);
nor U15078 (N_15078,N_13523,N_13649);
xor U15079 (N_15079,N_14281,N_14587);
xor U15080 (N_15080,N_14161,N_13956);
nand U15081 (N_15081,N_14193,N_14795);
xnor U15082 (N_15082,N_14935,N_14675);
nor U15083 (N_15083,N_14183,N_13554);
and U15084 (N_15084,N_13838,N_14635);
and U15085 (N_15085,N_14019,N_13984);
nor U15086 (N_15086,N_14704,N_13823);
xnor U15087 (N_15087,N_13761,N_13918);
and U15088 (N_15088,N_14246,N_14501);
xnor U15089 (N_15089,N_14738,N_14683);
xnor U15090 (N_15090,N_14583,N_14854);
and U15091 (N_15091,N_14911,N_13784);
or U15092 (N_15092,N_14776,N_14553);
or U15093 (N_15093,N_14745,N_13995);
xor U15094 (N_15094,N_14893,N_13971);
and U15095 (N_15095,N_14600,N_14385);
or U15096 (N_15096,N_13630,N_14310);
or U15097 (N_15097,N_14396,N_14855);
and U15098 (N_15098,N_14956,N_14621);
and U15099 (N_15099,N_14990,N_14392);
xnor U15100 (N_15100,N_14867,N_13763);
nor U15101 (N_15101,N_14925,N_13691);
nand U15102 (N_15102,N_14458,N_13876);
or U15103 (N_15103,N_14539,N_14850);
nor U15104 (N_15104,N_14934,N_13922);
nand U15105 (N_15105,N_13658,N_14444);
nand U15106 (N_15106,N_13874,N_14375);
xor U15107 (N_15107,N_14590,N_13800);
nand U15108 (N_15108,N_14651,N_14099);
xor U15109 (N_15109,N_14628,N_14185);
and U15110 (N_15110,N_14626,N_14705);
nand U15111 (N_15111,N_14992,N_14714);
or U15112 (N_15112,N_14870,N_14516);
nor U15113 (N_15113,N_13860,N_14221);
nand U15114 (N_15114,N_14423,N_14974);
and U15115 (N_15115,N_13768,N_13522);
nor U15116 (N_15116,N_14722,N_14359);
xor U15117 (N_15117,N_14749,N_14364);
and U15118 (N_15118,N_14228,N_13787);
and U15119 (N_15119,N_14674,N_13723);
or U15120 (N_15120,N_13737,N_14112);
nand U15121 (N_15121,N_14649,N_14519);
and U15122 (N_15122,N_13678,N_14414);
nand U15123 (N_15123,N_13694,N_14574);
nor U15124 (N_15124,N_13680,N_14888);
or U15125 (N_15125,N_13571,N_14291);
nand U15126 (N_15126,N_13529,N_14210);
or U15127 (N_15127,N_14912,N_14295);
and U15128 (N_15128,N_13968,N_14792);
nand U15129 (N_15129,N_14240,N_14089);
nor U15130 (N_15130,N_14110,N_13796);
and U15131 (N_15131,N_14128,N_13740);
or U15132 (N_15132,N_13607,N_14038);
xnor U15133 (N_15133,N_13891,N_14284);
and U15134 (N_15134,N_14329,N_14950);
nor U15135 (N_15135,N_14973,N_13766);
or U15136 (N_15136,N_14581,N_14834);
nand U15137 (N_15137,N_14464,N_14133);
xnor U15138 (N_15138,N_13750,N_13717);
or U15139 (N_15139,N_14126,N_14480);
nor U15140 (N_15140,N_14499,N_14890);
and U15141 (N_15141,N_13702,N_13786);
nand U15142 (N_15142,N_14546,N_13616);
and U15143 (N_15143,N_14802,N_14011);
xor U15144 (N_15144,N_13904,N_14339);
nor U15145 (N_15145,N_14779,N_14866);
nand U15146 (N_15146,N_14184,N_14765);
and U15147 (N_15147,N_14589,N_14378);
or U15148 (N_15148,N_13615,N_14862);
and U15149 (N_15149,N_13701,N_13520);
nor U15150 (N_15150,N_13928,N_14446);
or U15151 (N_15151,N_14715,N_14087);
and U15152 (N_15152,N_14354,N_13855);
or U15153 (N_15153,N_14025,N_13790);
nor U15154 (N_15154,N_14517,N_14009);
or U15155 (N_15155,N_14500,N_13703);
xnor U15156 (N_15156,N_14859,N_14819);
xnor U15157 (N_15157,N_14274,N_13955);
nand U15158 (N_15158,N_13612,N_14079);
nor U15159 (N_15159,N_14545,N_14638);
nor U15160 (N_15160,N_14209,N_13677);
xor U15161 (N_15161,N_13825,N_14777);
xnor U15162 (N_15162,N_14479,N_14767);
xor U15163 (N_15163,N_14556,N_13505);
or U15164 (N_15164,N_14968,N_14648);
xnor U15165 (N_15165,N_14491,N_14068);
nand U15166 (N_15166,N_14617,N_13921);
nand U15167 (N_15167,N_14980,N_13591);
nor U15168 (N_15168,N_14135,N_14681);
nor U15169 (N_15169,N_14677,N_14664);
nor U15170 (N_15170,N_14984,N_13683);
or U15171 (N_15171,N_13829,N_13791);
nor U15172 (N_15172,N_14450,N_14262);
xnor U15173 (N_15173,N_13705,N_14603);
or U15174 (N_15174,N_13912,N_14592);
xnor U15175 (N_15175,N_13555,N_14124);
and U15176 (N_15176,N_14914,N_14994);
or U15177 (N_15177,N_14780,N_14260);
and U15178 (N_15178,N_14254,N_13515);
or U15179 (N_15179,N_13863,N_14361);
nor U15180 (N_15180,N_14490,N_14559);
and U15181 (N_15181,N_13821,N_14709);
nor U15182 (N_15182,N_14131,N_13899);
xnor U15183 (N_15183,N_13714,N_14597);
nand U15184 (N_15184,N_14986,N_13903);
or U15185 (N_15185,N_14456,N_13660);
or U15186 (N_15186,N_13873,N_14407);
nand U15187 (N_15187,N_14646,N_13721);
nand U15188 (N_15188,N_14049,N_14257);
xnor U15189 (N_15189,N_13978,N_14477);
and U15190 (N_15190,N_13648,N_14729);
nor U15191 (N_15191,N_13983,N_14670);
and U15192 (N_15192,N_14614,N_14040);
and U15193 (N_15193,N_14271,N_14368);
or U15194 (N_15194,N_13746,N_14085);
xor U15195 (N_15195,N_14927,N_13656);
nand U15196 (N_15196,N_13655,N_13756);
xor U15197 (N_15197,N_13577,N_13887);
xnor U15198 (N_15198,N_13681,N_13896);
nand U15199 (N_15199,N_14759,N_13931);
and U15200 (N_15200,N_14886,N_14154);
xnor U15201 (N_15201,N_13826,N_13642);
or U15202 (N_15202,N_14379,N_13608);
nor U15203 (N_15203,N_14537,N_13913);
nand U15204 (N_15204,N_14008,N_14439);
and U15205 (N_15205,N_14384,N_14856);
xnor U15206 (N_15206,N_14946,N_13902);
or U15207 (N_15207,N_13996,N_14061);
and U15208 (N_15208,N_14461,N_14527);
xnor U15209 (N_15209,N_14043,N_13527);
nor U15210 (N_15210,N_13609,N_13933);
xnor U15211 (N_15211,N_14643,N_14791);
nand U15212 (N_15212,N_14506,N_13788);
and U15213 (N_15213,N_14966,N_14352);
xnor U15214 (N_15214,N_14066,N_14125);
or U15215 (N_15215,N_14272,N_14502);
nand U15216 (N_15216,N_14595,N_13862);
xnor U15217 (N_15217,N_13976,N_14957);
xnor U15218 (N_15218,N_14426,N_14719);
and U15219 (N_15219,N_14460,N_14144);
and U15220 (N_15220,N_13503,N_13831);
and U15221 (N_15221,N_14398,N_13946);
or U15222 (N_15222,N_14849,N_13954);
nand U15223 (N_15223,N_14931,N_13942);
nand U15224 (N_15224,N_14782,N_13603);
xor U15225 (N_15225,N_14687,N_14006);
xnor U15226 (N_15226,N_14826,N_14993);
xnor U15227 (N_15227,N_14402,N_14969);
or U15228 (N_15228,N_14425,N_13602);
nand U15229 (N_15229,N_14101,N_14665);
or U15230 (N_15230,N_13736,N_14568);
nand U15231 (N_15231,N_13715,N_14340);
nor U15232 (N_15232,N_13859,N_14454);
and U15233 (N_15233,N_14224,N_14732);
nor U15234 (N_15234,N_13731,N_13626);
xnor U15235 (N_15235,N_13911,N_14358);
xnor U15236 (N_15236,N_14013,N_14971);
nor U15237 (N_15237,N_14667,N_14998);
nand U15238 (N_15238,N_14744,N_13952);
xor U15239 (N_15239,N_14806,N_14843);
xnor U15240 (N_15240,N_14585,N_13592);
and U15241 (N_15241,N_13975,N_14899);
or U15242 (N_15242,N_13578,N_13854);
nor U15243 (N_15243,N_14050,N_14926);
or U15244 (N_15244,N_13651,N_13613);
and U15245 (N_15245,N_14678,N_13551);
or U15246 (N_15246,N_13751,N_13979);
or U15247 (N_15247,N_13594,N_14922);
nor U15248 (N_15248,N_14682,N_14466);
nor U15249 (N_15249,N_14472,N_14060);
xor U15250 (N_15250,N_14309,N_13687);
xnor U15251 (N_15251,N_14234,N_14147);
nor U15252 (N_15252,N_13764,N_13871);
xnor U15253 (N_15253,N_14959,N_14141);
or U15254 (N_15254,N_13560,N_13589);
xor U15255 (N_15255,N_13531,N_13919);
nor U15256 (N_15256,N_14955,N_14961);
nand U15257 (N_15257,N_14684,N_13518);
and U15258 (N_15258,N_13692,N_14443);
xor U15259 (N_15259,N_13628,N_13735);
nor U15260 (N_15260,N_14387,N_14057);
and U15261 (N_15261,N_14727,N_14067);
nand U15262 (N_15262,N_14647,N_14747);
xnor U15263 (N_15263,N_14740,N_13845);
or U15264 (N_15264,N_14278,N_14486);
nor U15265 (N_15265,N_14916,N_14077);
or U15266 (N_15266,N_13810,N_14967);
xor U15267 (N_15267,N_14140,N_14898);
xor U15268 (N_15268,N_13624,N_13980);
xor U15269 (N_15269,N_14962,N_14348);
and U15270 (N_15270,N_14430,N_14783);
nor U15271 (N_15271,N_14909,N_14253);
xnor U15272 (N_15272,N_14158,N_14988);
xor U15273 (N_15273,N_14523,N_14440);
nand U15274 (N_15274,N_14498,N_14534);
and U15275 (N_15275,N_13685,N_14794);
nand U15276 (N_15276,N_14422,N_14772);
or U15277 (N_15277,N_14321,N_13850);
xor U15278 (N_15278,N_14428,N_13501);
or U15279 (N_15279,N_13986,N_13948);
xor U15280 (N_15280,N_14939,N_13632);
or U15281 (N_15281,N_14541,N_13806);
nor U15282 (N_15282,N_14475,N_14768);
xor U15283 (N_15283,N_14434,N_14979);
nor U15284 (N_15284,N_13938,N_14718);
nand U15285 (N_15285,N_13789,N_14393);
nor U15286 (N_15286,N_14447,N_13546);
or U15287 (N_15287,N_14606,N_14573);
nor U15288 (N_15288,N_13879,N_14096);
nor U15289 (N_15289,N_14891,N_14508);
or U15290 (N_15290,N_13510,N_14676);
nor U15291 (N_15291,N_14997,N_14915);
and U15292 (N_15292,N_14238,N_14255);
xnor U15293 (N_15293,N_14908,N_14902);
nand U15294 (N_15294,N_14017,N_14380);
xnor U15295 (N_15295,N_13525,N_14847);
nand U15296 (N_15296,N_13797,N_13830);
or U15297 (N_15297,N_14503,N_13600);
xor U15298 (N_15298,N_13598,N_13550);
and U15299 (N_15299,N_14222,N_14163);
or U15300 (N_15300,N_13759,N_13727);
nand U15301 (N_15301,N_13851,N_14808);
or U15302 (N_15302,N_13910,N_14920);
and U15303 (N_15303,N_13623,N_14887);
nor U15304 (N_15304,N_13663,N_14044);
nand U15305 (N_15305,N_13892,N_14601);
or U15306 (N_15306,N_13524,N_13990);
or U15307 (N_15307,N_14411,N_13720);
nor U15308 (N_15308,N_13847,N_14235);
or U15309 (N_15309,N_14032,N_13569);
or U15310 (N_15310,N_13767,N_14416);
or U15311 (N_15311,N_14569,N_14232);
xnor U15312 (N_15312,N_14326,N_14552);
and U15313 (N_15313,N_14679,N_14243);
or U15314 (N_15314,N_14219,N_14473);
nor U15315 (N_15315,N_14356,N_13675);
nand U15316 (N_15316,N_14345,N_13724);
nand U15317 (N_15317,N_14165,N_14455);
or U15318 (N_15318,N_13568,N_14631);
and U15319 (N_15319,N_14069,N_14160);
or U15320 (N_15320,N_13534,N_14136);
nor U15321 (N_15321,N_13803,N_14882);
xnor U15322 (N_15322,N_14857,N_14696);
xor U15323 (N_15323,N_14283,N_13959);
or U15324 (N_15324,N_14338,N_14572);
xor U15325 (N_15325,N_13580,N_14880);
nor U15326 (N_15326,N_13940,N_13827);
xnor U15327 (N_15327,N_14204,N_14951);
xnor U15328 (N_15328,N_14410,N_13890);
xnor U15329 (N_15329,N_14304,N_14736);
and U15330 (N_15330,N_14143,N_13961);
nor U15331 (N_15331,N_13636,N_14972);
or U15332 (N_15332,N_14030,N_13745);
and U15333 (N_15333,N_14924,N_14536);
or U15334 (N_15334,N_13936,N_14525);
nor U15335 (N_15335,N_13590,N_14748);
and U15336 (N_15336,N_14730,N_14731);
or U15337 (N_15337,N_13993,N_13804);
and U15338 (N_15338,N_14644,N_14639);
nor U15339 (N_15339,N_13698,N_14839);
or U15340 (N_15340,N_14512,N_13950);
and U15341 (N_15341,N_14970,N_14487);
and U15342 (N_15342,N_14816,N_14325);
or U15343 (N_15343,N_14377,N_14835);
nor U15344 (N_15344,N_14016,N_14793);
nor U15345 (N_15345,N_13813,N_14943);
nor U15346 (N_15346,N_13856,N_14804);
xnor U15347 (N_15347,N_13849,N_14923);
and U15348 (N_15348,N_13639,N_14190);
and U15349 (N_15349,N_14493,N_14330);
xnor U15350 (N_15350,N_14632,N_14507);
or U15351 (N_15351,N_14755,N_14122);
nand U15352 (N_15352,N_14528,N_14494);
and U15353 (N_15353,N_14515,N_14865);
or U15354 (N_15354,N_14900,N_14137);
xnor U15355 (N_15355,N_13542,N_14435);
nor U15356 (N_15356,N_14168,N_14192);
nor U15357 (N_15357,N_14369,N_14815);
and U15358 (N_15358,N_14599,N_14029);
nor U15359 (N_15359,N_14024,N_14211);
nand U15360 (N_15360,N_14611,N_14342);
and U15361 (N_15361,N_13729,N_13593);
or U15362 (N_15362,N_14115,N_14483);
nand U15363 (N_15363,N_14797,N_14952);
nand U15364 (N_15364,N_13815,N_14072);
xnor U15365 (N_15365,N_13762,N_14273);
and U15366 (N_15366,N_14152,N_14659);
nor U15367 (N_15367,N_14906,N_13741);
nor U15368 (N_15368,N_14995,N_14015);
and U15369 (N_15369,N_14836,N_14596);
xnor U15370 (N_15370,N_14012,N_14186);
and U15371 (N_15371,N_13728,N_13917);
and U15372 (N_15372,N_13634,N_13670);
nand U15373 (N_15373,N_14509,N_14562);
nand U15374 (N_15374,N_13770,N_13604);
and U15375 (N_15375,N_14784,N_14723);
and U15376 (N_15376,N_13772,N_14874);
or U15377 (N_15377,N_14075,N_14018);
nor U15378 (N_15378,N_14231,N_14088);
xor U15379 (N_15379,N_14524,N_13570);
and U15380 (N_15380,N_14653,N_14641);
or U15381 (N_15381,N_14701,N_14177);
nand U15382 (N_15382,N_14975,N_14555);
xor U15383 (N_15383,N_14478,N_13595);
and U15384 (N_15384,N_13513,N_14206);
or U15385 (N_15385,N_14877,N_14520);
or U15386 (N_15386,N_14051,N_13758);
and U15387 (N_15387,N_14337,N_14708);
or U15388 (N_15388,N_14372,N_14002);
nor U15389 (N_15389,N_13844,N_14944);
or U15390 (N_15390,N_14362,N_14405);
and U15391 (N_15391,N_13755,N_14217);
or U15392 (N_15392,N_14551,N_14055);
or U15393 (N_15393,N_13629,N_13610);
xor U15394 (N_15394,N_14871,N_14307);
or U15395 (N_15395,N_14790,N_13884);
nand U15396 (N_15396,N_13834,N_14202);
or U15397 (N_15397,N_14063,N_14457);
or U15398 (N_15398,N_14563,N_13898);
nand U15399 (N_15399,N_13646,N_13519);
and U15400 (N_15400,N_13875,N_14420);
or U15401 (N_15401,N_14666,N_14170);
nor U15402 (N_15402,N_14250,N_14561);
or U15403 (N_15403,N_13953,N_14300);
and U15404 (N_15404,N_13753,N_14166);
nor U15405 (N_15405,N_13566,N_13915);
xnor U15406 (N_15406,N_14919,N_14251);
and U15407 (N_15407,N_14197,N_13504);
nand U15408 (N_15408,N_14225,N_14376);
and U15409 (N_15409,N_14070,N_13533);
and U15410 (N_15410,N_14513,N_14580);
and U15411 (N_15411,N_13599,N_13939);
xnor U15412 (N_15412,N_14937,N_13865);
xnor U15413 (N_15413,N_14276,N_14538);
and U15414 (N_15414,N_13857,N_14566);
xnor U15415 (N_15415,N_14108,N_14629);
xnor U15416 (N_15416,N_14860,N_13509);
nand U15417 (N_15417,N_13837,N_14150);
nand U15418 (N_15418,N_14540,N_13742);
nand U15419 (N_15419,N_14619,N_13638);
xor U15420 (N_15420,N_14894,N_14645);
or U15421 (N_15421,N_14695,N_14895);
nand U15422 (N_15422,N_14196,N_14633);
and U15423 (N_15423,N_13575,N_14288);
or U15424 (N_15424,N_13631,N_14181);
and U15425 (N_15425,N_14033,N_14770);
nand U15426 (N_15426,N_14109,N_14547);
nand U15427 (N_15427,N_13872,N_14370);
or U15428 (N_15428,N_13997,N_13671);
or U15429 (N_15429,N_14608,N_13977);
and U15430 (N_15430,N_13643,N_14786);
nor U15431 (N_15431,N_13511,N_14134);
or U15432 (N_15432,N_14987,N_14239);
or U15433 (N_15433,N_13726,N_13665);
nor U15434 (N_15434,N_14982,N_13982);
and U15435 (N_15435,N_13754,N_14468);
nor U15436 (N_15436,N_14242,N_14685);
nor U15437 (N_15437,N_13526,N_14218);
or U15438 (N_15438,N_14095,N_14699);
nor U15439 (N_15439,N_14864,N_14335);
nor U15440 (N_15440,N_13841,N_13916);
xnor U15441 (N_15441,N_14399,N_14053);
nor U15442 (N_15442,N_14167,N_13706);
or U15443 (N_15443,N_13926,N_14121);
nand U15444 (N_15444,N_14470,N_14227);
or U15445 (N_15445,N_14081,N_14169);
or U15446 (N_15446,N_13944,N_13565);
nor U15447 (N_15447,N_13878,N_13507);
or U15448 (N_15448,N_13969,N_13962);
nand U15449 (N_15449,N_14293,N_14964);
nor U15450 (N_15450,N_13693,N_14940);
or U15451 (N_15451,N_13802,N_14831);
xnor U15452 (N_15452,N_13500,N_14389);
or U15453 (N_15453,N_14693,N_14031);
nand U15454 (N_15454,N_14215,N_14236);
nand U15455 (N_15455,N_13757,N_14123);
xnor U15456 (N_15456,N_13819,N_14751);
or U15457 (N_15457,N_13981,N_14173);
nor U15458 (N_15458,N_14637,N_14948);
and U15459 (N_15459,N_13994,N_14820);
nand U15460 (N_15460,N_14421,N_14492);
xor U15461 (N_15461,N_13882,N_14901);
and U15462 (N_15462,N_13794,N_13773);
nor U15463 (N_15463,N_14876,N_14117);
or U15464 (N_15464,N_14145,N_14752);
nor U15465 (N_15465,N_13561,N_14721);
nand U15466 (N_15466,N_14766,N_13695);
nor U15467 (N_15467,N_13853,N_14413);
nand U15468 (N_15468,N_13645,N_14258);
and U15469 (N_15469,N_14602,N_14936);
and U15470 (N_15470,N_14607,N_13606);
or U15471 (N_15471,N_14333,N_13730);
xnor U15472 (N_15472,N_13579,N_13858);
nand U15473 (N_15473,N_14172,N_14153);
nand U15474 (N_15474,N_14958,N_14716);
and U15475 (N_15475,N_14408,N_14785);
nor U15476 (N_15476,N_14208,N_13782);
xnor U15477 (N_15477,N_14662,N_14471);
xor U15478 (N_15478,N_14037,N_13679);
and U15479 (N_15479,N_14848,N_13621);
nand U15480 (N_15480,N_14432,N_14741);
nor U15481 (N_15481,N_14195,N_13974);
nor U15482 (N_15482,N_14845,N_14981);
and U15483 (N_15483,N_13536,N_14954);
nor U15484 (N_15484,N_14199,N_13792);
and U15485 (N_15485,N_14686,N_13530);
or U15486 (N_15486,N_14698,N_13909);
or U15487 (N_15487,N_14489,N_14803);
nor U15488 (N_15488,N_14996,N_14700);
xnor U15489 (N_15489,N_13661,N_14022);
and U15490 (N_15490,N_14103,N_14388);
nor U15491 (N_15491,N_13894,N_14351);
nand U15492 (N_15492,N_14107,N_14842);
and U15493 (N_15493,N_14395,N_14827);
or U15494 (N_15494,N_14495,N_13676);
nor U15495 (N_15495,N_13664,N_13987);
nand U15496 (N_15496,N_14692,N_13704);
xor U15497 (N_15497,N_13930,N_14485);
xor U15498 (N_15498,N_13914,N_13833);
or U15499 (N_15499,N_14773,N_13732);
and U15500 (N_15500,N_14394,N_14484);
xor U15501 (N_15501,N_13895,N_14286);
nor U15502 (N_15502,N_14120,N_13541);
nand U15503 (N_15503,N_14775,N_14324);
or U15504 (N_15504,N_13795,N_14858);
xor U15505 (N_15505,N_13588,N_14365);
nand U15506 (N_15506,N_14837,N_14381);
nor U15507 (N_15507,N_14280,N_14263);
and U15508 (N_15508,N_14076,N_14869);
nor U15509 (N_15509,N_14656,N_14613);
nand U15510 (N_15510,N_14203,N_13548);
or U15511 (N_15511,N_13585,N_13809);
nor U15512 (N_15512,N_14965,N_14505);
and U15513 (N_15513,N_13958,N_14593);
and U15514 (N_15514,N_14347,N_14091);
or U15515 (N_15515,N_14207,N_14156);
or U15516 (N_15516,N_14609,N_14298);
or U15517 (N_15517,N_14294,N_13668);
or U15518 (N_15518,N_13998,N_14200);
or U15519 (N_15519,N_14431,N_13743);
or U15520 (N_15520,N_14297,N_14514);
nor U15521 (N_15521,N_14554,N_13799);
nor U15522 (N_15522,N_14266,N_13584);
and U15523 (N_15523,N_14360,N_13870);
xnor U15524 (N_15524,N_14724,N_13744);
nand U15525 (N_15525,N_14316,N_14373);
nand U15526 (N_15526,N_13707,N_14176);
nor U15527 (N_15527,N_14734,N_13970);
or U15528 (N_15528,N_13749,N_13777);
nand U15529 (N_15529,N_14873,N_14279);
or U15530 (N_15530,N_14247,N_14833);
or U15531 (N_15531,N_14575,N_13843);
and U15532 (N_15532,N_14320,N_13713);
or U15533 (N_15533,N_13963,N_13818);
and U15534 (N_15534,N_14760,N_13653);
nor U15535 (N_15535,N_13929,N_14059);
or U15536 (N_15536,N_13556,N_13672);
xnor U15537 (N_15537,N_14884,N_13625);
and U15538 (N_15538,N_14921,N_14159);
and U15539 (N_15539,N_13880,N_14442);
nand U15540 (N_15540,N_13562,N_14311);
xor U15541 (N_15541,N_14312,N_14750);
and U15542 (N_15542,N_14976,N_13908);
nor U15543 (N_15543,N_14074,N_14229);
and U15544 (N_15544,N_14463,N_14182);
and U15545 (N_15545,N_14710,N_13965);
and U15546 (N_15546,N_14164,N_14102);
or U15547 (N_15547,N_13733,N_14567);
nand U15548 (N_15548,N_14812,N_13771);
xnor U15549 (N_15549,N_14746,N_13785);
nor U15550 (N_15550,N_13920,N_14707);
nand U15551 (N_15551,N_14459,N_14357);
and U15552 (N_15552,N_14840,N_13798);
xor U15553 (N_15553,N_14001,N_14374);
nand U15554 (N_15554,N_14598,N_13549);
and U15555 (N_15555,N_14963,N_13618);
nand U15556 (N_15556,N_14548,N_13709);
xnor U15557 (N_15557,N_13506,N_14634);
nand U15558 (N_15558,N_14056,N_13640);
and U15559 (N_15559,N_13597,N_14577);
or U15560 (N_15560,N_14390,N_13852);
nor U15561 (N_15561,N_14449,N_14244);
nor U15562 (N_15562,N_13508,N_14346);
or U15563 (N_15563,N_13927,N_13538);
nor U15564 (N_15564,N_13712,N_13985);
nor U15565 (N_15565,N_14753,N_13828);
nor U15566 (N_15566,N_14669,N_14194);
and U15567 (N_15567,N_13708,N_13960);
and U15568 (N_15568,N_14078,N_13868);
and U15569 (N_15569,N_14532,N_14327);
or U15570 (N_15570,N_13543,N_14809);
and U15571 (N_15571,N_14712,N_14821);
nor U15572 (N_15572,N_14094,N_13725);
nand U15573 (N_15573,N_14113,N_14942);
nor U15574 (N_15574,N_14178,N_14267);
nor U15575 (N_15575,N_14875,N_14162);
xnor U15576 (N_15576,N_13807,N_14838);
or U15577 (N_15577,N_14130,N_14064);
nor U15578 (N_15578,N_14149,N_14465);
nand U15579 (N_15579,N_13774,N_14851);
and U15580 (N_15580,N_14082,N_14841);
xor U15581 (N_15581,N_13832,N_13805);
xnor U15582 (N_15582,N_13893,N_14132);
nor U15583 (N_15583,N_13776,N_14726);
or U15584 (N_15584,N_14832,N_14268);
and U15585 (N_15585,N_14542,N_13669);
and U15586 (N_15586,N_14148,N_14518);
and U15587 (N_15587,N_14249,N_13697);
and U15588 (N_15588,N_14269,N_14822);
xnor U15589 (N_15589,N_14497,N_14879);
or U15590 (N_15590,N_13667,N_13516);
xnor U15591 (N_15591,N_14171,N_14445);
and U15592 (N_15592,N_14933,N_14620);
xor U15593 (N_15593,N_14844,N_13824);
or U15594 (N_15594,N_14618,N_14308);
nor U15595 (N_15595,N_13752,N_14086);
or U15596 (N_15596,N_13719,N_14080);
xor U15597 (N_15597,N_14302,N_14366);
and U15598 (N_15598,N_14142,N_14315);
nand U15599 (N_15599,N_14448,N_13817);
and U15600 (N_15600,N_13582,N_14438);
nand U15601 (N_15601,N_14127,N_13528);
nor U15602 (N_15602,N_14823,N_13989);
xor U15603 (N_15603,N_13710,N_14469);
or U15604 (N_15604,N_13674,N_14047);
or U15605 (N_15605,N_14021,N_13637);
nand U15606 (N_15606,N_14046,N_13662);
nand U15607 (N_15607,N_14332,N_14863);
nand U15608 (N_15608,N_13897,N_14591);
nand U15609 (N_15609,N_14035,N_14624);
or U15610 (N_15610,N_13711,N_14928);
nor U15611 (N_15611,N_13686,N_14282);
nor U15612 (N_15612,N_14735,N_14522);
xor U15613 (N_15613,N_13957,N_14872);
nand U15614 (N_15614,N_13812,N_13547);
nor U15615 (N_15615,N_14116,N_13659);
nand U15616 (N_15616,N_13905,N_14256);
and U15617 (N_15617,N_13576,N_13747);
nand U15618 (N_15618,N_13605,N_13992);
nand U15619 (N_15619,N_13559,N_13716);
xnor U15620 (N_15620,N_14349,N_14026);
nand U15621 (N_15621,N_14277,N_14654);
xnor U15622 (N_15622,N_14083,N_14129);
nor U15623 (N_15623,N_14437,N_14328);
or U15624 (N_15624,N_14612,N_14363);
nand U15625 (N_15625,N_14073,N_14400);
and U15626 (N_15626,N_13947,N_13867);
and U15627 (N_15627,N_13783,N_14205);
or U15628 (N_15628,N_14885,N_13552);
xor U15629 (N_15629,N_14467,N_14391);
or U15630 (N_15630,N_14093,N_14322);
and U15631 (N_15631,N_14452,N_14042);
xnor U15632 (N_15632,N_13814,N_14763);
and U15633 (N_15633,N_14694,N_14424);
xnor U15634 (N_15634,N_14787,N_13999);
nand U15635 (N_15635,N_14985,N_14000);
nand U15636 (N_15636,N_14441,N_13574);
and U15637 (N_15637,N_14828,N_14010);
nor U15638 (N_15638,N_14868,N_13563);
nand U15639 (N_15639,N_14918,N_14622);
or U15640 (N_15640,N_13619,N_14703);
nand U15641 (N_15641,N_13808,N_14549);
or U15642 (N_15642,N_14481,N_14138);
and U15643 (N_15643,N_13682,N_13545);
nand U15644 (N_15644,N_13861,N_14230);
xnor U15645 (N_15645,N_14531,N_13699);
or U15646 (N_15646,N_13535,N_14265);
xnor U15647 (N_15647,N_13816,N_14586);
nor U15648 (N_15648,N_14259,N_13846);
nand U15649 (N_15649,N_13734,N_13967);
or U15650 (N_15650,N_14739,N_13622);
and U15651 (N_15651,N_14334,N_14652);
and U15652 (N_15652,N_13924,N_13835);
and U15653 (N_15653,N_13611,N_14830);
nor U15654 (N_15654,N_13934,N_14301);
or U15655 (N_15655,N_13973,N_13778);
nor U15656 (N_15656,N_14003,N_14801);
nor U15657 (N_15657,N_14245,N_13581);
or U15658 (N_15658,N_14355,N_13951);
nand U15659 (N_15659,N_14155,N_14409);
or U15660 (N_15660,N_14829,N_14453);
and U15661 (N_15661,N_14781,N_14799);
or U15662 (N_15662,N_14800,N_14903);
nand U15663 (N_15663,N_14382,N_14223);
nand U15664 (N_15664,N_14807,N_14878);
nor U15665 (N_15665,N_14824,N_14576);
or U15666 (N_15666,N_13760,N_14299);
xor U15667 (N_15667,N_14579,N_13688);
nor U15668 (N_15668,N_14625,N_14661);
xor U15669 (N_15669,N_14412,N_14028);
nand U15670 (N_15670,N_14104,N_14989);
nor U15671 (N_15671,N_14174,N_14097);
nor U15672 (N_15672,N_14761,N_14558);
and U15673 (N_15673,N_14892,N_14977);
nand U15674 (N_15674,N_14680,N_14725);
or U15675 (N_15675,N_14004,N_14754);
or U15676 (N_15676,N_14743,N_14616);
nand U15677 (N_15677,N_14292,N_14226);
and U15678 (N_15678,N_13811,N_13540);
or U15679 (N_15679,N_14353,N_14041);
nor U15680 (N_15680,N_13901,N_14341);
nor U15681 (N_15681,N_14630,N_13877);
or U15682 (N_15682,N_13848,N_14883);
nor U15683 (N_15683,N_13722,N_14100);
xnor U15684 (N_15684,N_13900,N_14717);
or U15685 (N_15685,N_14910,N_13881);
nand U15686 (N_15686,N_13666,N_14582);
xnor U15687 (N_15687,N_14290,N_14023);
nor U15688 (N_15688,N_14314,N_14938);
nor U15689 (N_15689,N_14157,N_13883);
nor U15690 (N_15690,N_14564,N_14289);
or U15691 (N_15691,N_14090,N_14588);
nor U15692 (N_15692,N_14672,N_14571);
nor U15693 (N_15693,N_14034,N_14526);
or U15694 (N_15694,N_14742,N_13614);
and U15695 (N_15695,N_14429,N_14146);
xor U15696 (N_15696,N_14118,N_14323);
xor U15697 (N_15697,N_13689,N_14660);
nor U15698 (N_15698,N_14702,N_14584);
xnor U15699 (N_15699,N_14401,N_14313);
or U15700 (N_15700,N_14476,N_13647);
nand U15701 (N_15701,N_14433,N_13889);
nand U15702 (N_15702,N_14697,N_14336);
and U15703 (N_15703,N_14657,N_14913);
and U15704 (N_15704,N_14673,N_14535);
xnor U15705 (N_15705,N_14999,N_14062);
xnor U15706 (N_15706,N_14557,N_14788);
and U15707 (N_15707,N_13769,N_14252);
or U15708 (N_15708,N_13544,N_13801);
xnor U15709 (N_15709,N_14180,N_14917);
xnor U15710 (N_15710,N_14462,N_13652);
nand U15711 (N_15711,N_14949,N_14983);
nor U15712 (N_15712,N_14397,N_14045);
and U15713 (N_15713,N_14331,N_13641);
nor U15714 (N_15714,N_14403,N_14098);
xor U15715 (N_15715,N_13923,N_14733);
nor U15716 (N_15716,N_14198,N_13869);
nand U15717 (N_15717,N_14861,N_14947);
or U15718 (N_15718,N_14778,N_13573);
nand U15719 (N_15719,N_14544,N_14139);
nand U15720 (N_15720,N_13673,N_14905);
and U15721 (N_15721,N_14941,N_14769);
or U15722 (N_15722,N_14305,N_14105);
and U15723 (N_15723,N_14427,N_13935);
or U15724 (N_15724,N_13839,N_13945);
and U15725 (N_15725,N_14504,N_14798);
nor U15726 (N_15726,N_14805,N_14690);
or U15727 (N_15727,N_14188,N_13517);
and U15728 (N_15728,N_14214,N_14451);
or U15729 (N_15729,N_13739,N_14318);
nor U15730 (N_15730,N_14691,N_14191);
xor U15731 (N_15731,N_14655,N_14530);
nor U15732 (N_15732,N_14570,N_13888);
and U15733 (N_15733,N_14213,N_13949);
xor U15734 (N_15734,N_13572,N_14853);
or U15735 (N_15735,N_14713,N_14953);
nand U15736 (N_15736,N_14084,N_14092);
nand U15737 (N_15737,N_13842,N_14303);
nand U15738 (N_15738,N_14771,N_14111);
or U15739 (N_15739,N_14543,N_14904);
nor U15740 (N_15740,N_13775,N_14488);
xnor U15741 (N_15741,N_14565,N_14404);
nor U15742 (N_15742,N_14415,N_13866);
and U15743 (N_15743,N_14261,N_13521);
and U15744 (N_15744,N_14187,N_13765);
nand U15745 (N_15745,N_14317,N_14005);
xor U15746 (N_15746,N_13644,N_14014);
and U15747 (N_15747,N_13886,N_13925);
nand U15748 (N_15748,N_14818,N_13972);
nor U15749 (N_15749,N_13991,N_14627);
nor U15750 (N_15750,N_14957,N_14517);
xnor U15751 (N_15751,N_13903,N_13922);
xnor U15752 (N_15752,N_14170,N_14626);
nand U15753 (N_15753,N_14244,N_13869);
nand U15754 (N_15754,N_14610,N_14352);
nand U15755 (N_15755,N_14807,N_14682);
nand U15756 (N_15756,N_14725,N_14062);
nand U15757 (N_15757,N_13530,N_13622);
nand U15758 (N_15758,N_14880,N_14246);
nand U15759 (N_15759,N_14809,N_13678);
or U15760 (N_15760,N_13612,N_14544);
and U15761 (N_15761,N_14998,N_14108);
and U15762 (N_15762,N_14369,N_14058);
and U15763 (N_15763,N_13926,N_14315);
and U15764 (N_15764,N_13521,N_14087);
nor U15765 (N_15765,N_14111,N_13972);
and U15766 (N_15766,N_13901,N_14451);
nor U15767 (N_15767,N_13806,N_14046);
nand U15768 (N_15768,N_13866,N_13892);
xnor U15769 (N_15769,N_13589,N_14740);
nand U15770 (N_15770,N_13929,N_13768);
or U15771 (N_15771,N_14165,N_14605);
nor U15772 (N_15772,N_14203,N_14639);
xor U15773 (N_15773,N_13749,N_14323);
or U15774 (N_15774,N_14700,N_13980);
nor U15775 (N_15775,N_14433,N_14904);
nor U15776 (N_15776,N_14109,N_13867);
xnor U15777 (N_15777,N_13581,N_14146);
or U15778 (N_15778,N_14027,N_13570);
nand U15779 (N_15779,N_14135,N_13640);
xor U15780 (N_15780,N_14184,N_14790);
nand U15781 (N_15781,N_14496,N_14291);
or U15782 (N_15782,N_14534,N_14119);
nand U15783 (N_15783,N_14973,N_13538);
and U15784 (N_15784,N_13558,N_14939);
and U15785 (N_15785,N_14896,N_14651);
and U15786 (N_15786,N_14922,N_13645);
xor U15787 (N_15787,N_14387,N_14710);
nor U15788 (N_15788,N_13624,N_13706);
nand U15789 (N_15789,N_14005,N_14679);
xnor U15790 (N_15790,N_14017,N_13821);
nand U15791 (N_15791,N_14012,N_14031);
xnor U15792 (N_15792,N_14923,N_13698);
xor U15793 (N_15793,N_14754,N_14426);
nand U15794 (N_15794,N_13981,N_14288);
xor U15795 (N_15795,N_14760,N_14770);
nor U15796 (N_15796,N_14667,N_14958);
xnor U15797 (N_15797,N_14302,N_14161);
and U15798 (N_15798,N_14708,N_14799);
nand U15799 (N_15799,N_13936,N_14330);
nand U15800 (N_15800,N_14215,N_13582);
or U15801 (N_15801,N_14699,N_13833);
nor U15802 (N_15802,N_13712,N_14615);
nand U15803 (N_15803,N_14846,N_13634);
nand U15804 (N_15804,N_14788,N_13984);
xor U15805 (N_15805,N_13778,N_14076);
xnor U15806 (N_15806,N_13580,N_14151);
and U15807 (N_15807,N_14424,N_14980);
nor U15808 (N_15808,N_13681,N_14959);
nand U15809 (N_15809,N_14018,N_14061);
xnor U15810 (N_15810,N_13730,N_14135);
nor U15811 (N_15811,N_14355,N_13644);
or U15812 (N_15812,N_14481,N_13917);
or U15813 (N_15813,N_14436,N_14163);
or U15814 (N_15814,N_13977,N_14631);
nand U15815 (N_15815,N_14622,N_14625);
nand U15816 (N_15816,N_14992,N_14989);
nor U15817 (N_15817,N_14595,N_13826);
or U15818 (N_15818,N_14588,N_14713);
xnor U15819 (N_15819,N_14678,N_13693);
and U15820 (N_15820,N_14181,N_14344);
nand U15821 (N_15821,N_13681,N_14306);
nand U15822 (N_15822,N_13721,N_14453);
or U15823 (N_15823,N_14298,N_14930);
nand U15824 (N_15824,N_14348,N_14874);
xor U15825 (N_15825,N_14765,N_14012);
nand U15826 (N_15826,N_14360,N_14993);
nand U15827 (N_15827,N_14717,N_14638);
and U15828 (N_15828,N_14679,N_14923);
xnor U15829 (N_15829,N_14677,N_13957);
nor U15830 (N_15830,N_14687,N_14299);
xor U15831 (N_15831,N_14343,N_14293);
and U15832 (N_15832,N_13661,N_14506);
xor U15833 (N_15833,N_13623,N_14400);
nand U15834 (N_15834,N_14361,N_14065);
nand U15835 (N_15835,N_14197,N_13541);
nand U15836 (N_15836,N_13991,N_14299);
nand U15837 (N_15837,N_14563,N_14069);
nor U15838 (N_15838,N_14635,N_13566);
and U15839 (N_15839,N_13519,N_14375);
xor U15840 (N_15840,N_13956,N_14150);
and U15841 (N_15841,N_13549,N_14460);
xnor U15842 (N_15842,N_14981,N_14178);
nor U15843 (N_15843,N_14950,N_14341);
or U15844 (N_15844,N_13905,N_13866);
nand U15845 (N_15845,N_14085,N_14633);
and U15846 (N_15846,N_13513,N_14337);
xnor U15847 (N_15847,N_14838,N_14359);
and U15848 (N_15848,N_14272,N_14755);
nor U15849 (N_15849,N_14332,N_14249);
and U15850 (N_15850,N_14126,N_13843);
and U15851 (N_15851,N_14507,N_14601);
nor U15852 (N_15852,N_14007,N_14204);
and U15853 (N_15853,N_13570,N_14510);
xor U15854 (N_15854,N_14725,N_14822);
and U15855 (N_15855,N_14685,N_14540);
xnor U15856 (N_15856,N_13969,N_14501);
nor U15857 (N_15857,N_14574,N_14344);
nor U15858 (N_15858,N_14394,N_14023);
nor U15859 (N_15859,N_14593,N_14654);
nor U15860 (N_15860,N_14432,N_13927);
nor U15861 (N_15861,N_13941,N_14473);
xnor U15862 (N_15862,N_13903,N_14583);
nor U15863 (N_15863,N_13686,N_14141);
xnor U15864 (N_15864,N_14755,N_14526);
nand U15865 (N_15865,N_14544,N_14938);
and U15866 (N_15866,N_14674,N_13526);
or U15867 (N_15867,N_14320,N_14840);
and U15868 (N_15868,N_13643,N_14409);
nand U15869 (N_15869,N_13883,N_14154);
xnor U15870 (N_15870,N_13938,N_14199);
or U15871 (N_15871,N_14413,N_13650);
or U15872 (N_15872,N_13777,N_14124);
nand U15873 (N_15873,N_14530,N_13983);
xnor U15874 (N_15874,N_13805,N_13795);
nor U15875 (N_15875,N_13564,N_13740);
and U15876 (N_15876,N_13802,N_14465);
nand U15877 (N_15877,N_14825,N_14242);
and U15878 (N_15878,N_14861,N_14500);
and U15879 (N_15879,N_14603,N_13824);
or U15880 (N_15880,N_14833,N_14311);
nand U15881 (N_15881,N_14904,N_13661);
nand U15882 (N_15882,N_14803,N_13687);
nor U15883 (N_15883,N_14562,N_13575);
nor U15884 (N_15884,N_14851,N_14816);
nand U15885 (N_15885,N_13965,N_13866);
or U15886 (N_15886,N_13979,N_14616);
or U15887 (N_15887,N_14901,N_14994);
xor U15888 (N_15888,N_14943,N_14392);
or U15889 (N_15889,N_14632,N_14533);
and U15890 (N_15890,N_14699,N_14251);
nand U15891 (N_15891,N_14459,N_14114);
or U15892 (N_15892,N_14947,N_14552);
and U15893 (N_15893,N_13876,N_14623);
or U15894 (N_15894,N_14575,N_14351);
nor U15895 (N_15895,N_14200,N_14650);
xnor U15896 (N_15896,N_14640,N_14506);
or U15897 (N_15897,N_14419,N_14842);
nand U15898 (N_15898,N_14484,N_14871);
xor U15899 (N_15899,N_14702,N_14921);
or U15900 (N_15900,N_13891,N_13627);
nor U15901 (N_15901,N_13560,N_13986);
nand U15902 (N_15902,N_14840,N_14895);
xor U15903 (N_15903,N_13888,N_14909);
or U15904 (N_15904,N_14758,N_14549);
xnor U15905 (N_15905,N_14394,N_14071);
xnor U15906 (N_15906,N_14822,N_14169);
nand U15907 (N_15907,N_14982,N_14256);
and U15908 (N_15908,N_14274,N_14466);
nand U15909 (N_15909,N_14470,N_14785);
and U15910 (N_15910,N_14484,N_14365);
xor U15911 (N_15911,N_13873,N_14925);
nand U15912 (N_15912,N_14524,N_13546);
xor U15913 (N_15913,N_13521,N_14680);
and U15914 (N_15914,N_14243,N_14981);
nand U15915 (N_15915,N_13942,N_14809);
xor U15916 (N_15916,N_14048,N_14834);
or U15917 (N_15917,N_14366,N_14694);
xor U15918 (N_15918,N_14559,N_14992);
xnor U15919 (N_15919,N_14804,N_13591);
or U15920 (N_15920,N_14666,N_14826);
nand U15921 (N_15921,N_13506,N_13855);
nand U15922 (N_15922,N_14550,N_14786);
nor U15923 (N_15923,N_14080,N_14320);
and U15924 (N_15924,N_13941,N_13736);
xnor U15925 (N_15925,N_13671,N_13851);
nor U15926 (N_15926,N_14365,N_13500);
or U15927 (N_15927,N_13931,N_13814);
xnor U15928 (N_15928,N_14949,N_13571);
xor U15929 (N_15929,N_13951,N_13811);
xor U15930 (N_15930,N_13547,N_13608);
or U15931 (N_15931,N_14928,N_14740);
or U15932 (N_15932,N_14723,N_14771);
and U15933 (N_15933,N_14017,N_13577);
xor U15934 (N_15934,N_14440,N_14800);
or U15935 (N_15935,N_14606,N_13502);
or U15936 (N_15936,N_13975,N_14406);
and U15937 (N_15937,N_13858,N_13652);
xnor U15938 (N_15938,N_14601,N_13878);
nor U15939 (N_15939,N_14184,N_13523);
or U15940 (N_15940,N_14798,N_14983);
nand U15941 (N_15941,N_13516,N_14701);
nand U15942 (N_15942,N_14098,N_14229);
and U15943 (N_15943,N_14053,N_14863);
and U15944 (N_15944,N_14731,N_14618);
and U15945 (N_15945,N_13661,N_14248);
or U15946 (N_15946,N_14449,N_14564);
nand U15947 (N_15947,N_14016,N_14658);
or U15948 (N_15948,N_13623,N_14427);
xor U15949 (N_15949,N_14786,N_13738);
nand U15950 (N_15950,N_14606,N_14347);
nand U15951 (N_15951,N_14854,N_13860);
xor U15952 (N_15952,N_13711,N_14703);
nor U15953 (N_15953,N_14248,N_14330);
and U15954 (N_15954,N_14541,N_14045);
or U15955 (N_15955,N_14273,N_14344);
and U15956 (N_15956,N_13607,N_14242);
or U15957 (N_15957,N_13710,N_14673);
nand U15958 (N_15958,N_14391,N_14454);
and U15959 (N_15959,N_14000,N_14123);
or U15960 (N_15960,N_14390,N_14419);
nand U15961 (N_15961,N_14308,N_14855);
xnor U15962 (N_15962,N_14206,N_14127);
nand U15963 (N_15963,N_13721,N_14377);
or U15964 (N_15964,N_14944,N_14312);
xnor U15965 (N_15965,N_13911,N_14128);
xnor U15966 (N_15966,N_13672,N_13669);
nor U15967 (N_15967,N_14549,N_14544);
or U15968 (N_15968,N_14891,N_14692);
xnor U15969 (N_15969,N_13739,N_14796);
nor U15970 (N_15970,N_14137,N_14983);
nor U15971 (N_15971,N_14244,N_14672);
or U15972 (N_15972,N_14641,N_13806);
nor U15973 (N_15973,N_14178,N_13593);
nand U15974 (N_15974,N_14194,N_13829);
xnor U15975 (N_15975,N_13955,N_14693);
xnor U15976 (N_15976,N_13905,N_14241);
or U15977 (N_15977,N_14361,N_14334);
nand U15978 (N_15978,N_14186,N_14082);
nor U15979 (N_15979,N_14256,N_14123);
xnor U15980 (N_15980,N_14118,N_13822);
and U15981 (N_15981,N_14900,N_13687);
nor U15982 (N_15982,N_14402,N_14513);
or U15983 (N_15983,N_13533,N_14481);
xor U15984 (N_15984,N_14872,N_13627);
or U15985 (N_15985,N_14856,N_14878);
nand U15986 (N_15986,N_14064,N_14841);
or U15987 (N_15987,N_14880,N_13542);
nor U15988 (N_15988,N_14068,N_14044);
nor U15989 (N_15989,N_14824,N_14170);
xnor U15990 (N_15990,N_14805,N_14354);
or U15991 (N_15991,N_14930,N_14861);
nor U15992 (N_15992,N_13683,N_13846);
nor U15993 (N_15993,N_13621,N_14371);
nor U15994 (N_15994,N_14076,N_14772);
nand U15995 (N_15995,N_14870,N_14855);
and U15996 (N_15996,N_14082,N_13999);
or U15997 (N_15997,N_14114,N_14235);
xnor U15998 (N_15998,N_13999,N_13736);
nand U15999 (N_15999,N_13846,N_14251);
nor U16000 (N_16000,N_13612,N_14694);
or U16001 (N_16001,N_13632,N_14781);
and U16002 (N_16002,N_14992,N_13695);
nor U16003 (N_16003,N_13618,N_13661);
or U16004 (N_16004,N_14430,N_14280);
xor U16005 (N_16005,N_14714,N_13939);
nor U16006 (N_16006,N_14160,N_14199);
nor U16007 (N_16007,N_14177,N_14045);
and U16008 (N_16008,N_14545,N_14873);
xnor U16009 (N_16009,N_14895,N_13918);
nor U16010 (N_16010,N_13760,N_13957);
nand U16011 (N_16011,N_14485,N_13569);
or U16012 (N_16012,N_13604,N_14584);
and U16013 (N_16013,N_13846,N_14451);
and U16014 (N_16014,N_14469,N_14353);
and U16015 (N_16015,N_13812,N_14665);
nor U16016 (N_16016,N_13924,N_13917);
and U16017 (N_16017,N_14236,N_14372);
xor U16018 (N_16018,N_13748,N_14648);
or U16019 (N_16019,N_14483,N_14204);
and U16020 (N_16020,N_14162,N_13758);
and U16021 (N_16021,N_14015,N_14063);
xor U16022 (N_16022,N_14533,N_14082);
or U16023 (N_16023,N_14128,N_13507);
nand U16024 (N_16024,N_13799,N_13715);
nand U16025 (N_16025,N_14878,N_14765);
nand U16026 (N_16026,N_14286,N_13725);
and U16027 (N_16027,N_13517,N_14574);
xor U16028 (N_16028,N_14520,N_14730);
nand U16029 (N_16029,N_14934,N_13651);
and U16030 (N_16030,N_14557,N_14113);
nand U16031 (N_16031,N_13511,N_14363);
or U16032 (N_16032,N_14075,N_13947);
nor U16033 (N_16033,N_14331,N_14660);
nor U16034 (N_16034,N_14054,N_14722);
nand U16035 (N_16035,N_13968,N_13777);
or U16036 (N_16036,N_13889,N_14582);
and U16037 (N_16037,N_14275,N_14036);
xor U16038 (N_16038,N_13672,N_14575);
nand U16039 (N_16039,N_14126,N_14588);
nand U16040 (N_16040,N_14169,N_14662);
nor U16041 (N_16041,N_14869,N_14543);
nor U16042 (N_16042,N_14087,N_14772);
nand U16043 (N_16043,N_14519,N_14564);
or U16044 (N_16044,N_14320,N_13911);
and U16045 (N_16045,N_14881,N_13765);
xnor U16046 (N_16046,N_13560,N_14851);
nor U16047 (N_16047,N_14736,N_14815);
and U16048 (N_16048,N_14869,N_13555);
nand U16049 (N_16049,N_14163,N_14040);
nor U16050 (N_16050,N_14536,N_14693);
and U16051 (N_16051,N_13741,N_14993);
nand U16052 (N_16052,N_14711,N_14835);
or U16053 (N_16053,N_14489,N_14420);
and U16054 (N_16054,N_13941,N_13640);
and U16055 (N_16055,N_13674,N_14450);
and U16056 (N_16056,N_14885,N_14319);
xnor U16057 (N_16057,N_13812,N_14168);
and U16058 (N_16058,N_13653,N_14769);
and U16059 (N_16059,N_13977,N_13756);
and U16060 (N_16060,N_14725,N_13546);
xnor U16061 (N_16061,N_13851,N_14653);
nor U16062 (N_16062,N_14055,N_13504);
and U16063 (N_16063,N_14675,N_14007);
or U16064 (N_16064,N_14681,N_14412);
xnor U16065 (N_16065,N_14127,N_13944);
nor U16066 (N_16066,N_13940,N_14938);
nor U16067 (N_16067,N_14933,N_14556);
nor U16068 (N_16068,N_14358,N_14972);
or U16069 (N_16069,N_13995,N_14467);
and U16070 (N_16070,N_13690,N_14575);
xnor U16071 (N_16071,N_14641,N_13957);
or U16072 (N_16072,N_13976,N_14160);
nand U16073 (N_16073,N_14526,N_14521);
xor U16074 (N_16074,N_14194,N_13791);
and U16075 (N_16075,N_13537,N_13630);
xnor U16076 (N_16076,N_14115,N_14060);
and U16077 (N_16077,N_13773,N_13531);
or U16078 (N_16078,N_13984,N_14671);
nor U16079 (N_16079,N_14617,N_13874);
or U16080 (N_16080,N_14157,N_14158);
or U16081 (N_16081,N_14691,N_13808);
nand U16082 (N_16082,N_13682,N_14120);
or U16083 (N_16083,N_14152,N_14678);
nor U16084 (N_16084,N_14999,N_13622);
nor U16085 (N_16085,N_14944,N_14986);
nand U16086 (N_16086,N_14466,N_14628);
and U16087 (N_16087,N_14411,N_14939);
or U16088 (N_16088,N_14836,N_14648);
xnor U16089 (N_16089,N_14303,N_13512);
xnor U16090 (N_16090,N_13628,N_14541);
xnor U16091 (N_16091,N_13961,N_14819);
or U16092 (N_16092,N_14933,N_14715);
or U16093 (N_16093,N_13979,N_14535);
nor U16094 (N_16094,N_14273,N_14575);
nor U16095 (N_16095,N_13512,N_14449);
xnor U16096 (N_16096,N_13873,N_14136);
xnor U16097 (N_16097,N_14992,N_13843);
and U16098 (N_16098,N_14347,N_14602);
or U16099 (N_16099,N_14337,N_13762);
nand U16100 (N_16100,N_14581,N_14965);
nand U16101 (N_16101,N_14848,N_14540);
or U16102 (N_16102,N_13593,N_14754);
nor U16103 (N_16103,N_13687,N_14312);
nand U16104 (N_16104,N_14107,N_13737);
nor U16105 (N_16105,N_14478,N_14995);
and U16106 (N_16106,N_14587,N_13713);
and U16107 (N_16107,N_14291,N_14337);
nand U16108 (N_16108,N_13882,N_14598);
nand U16109 (N_16109,N_14567,N_13929);
nor U16110 (N_16110,N_14543,N_14284);
or U16111 (N_16111,N_14002,N_14216);
or U16112 (N_16112,N_14396,N_14470);
or U16113 (N_16113,N_14298,N_14892);
xnor U16114 (N_16114,N_13500,N_14495);
nand U16115 (N_16115,N_13846,N_14385);
nor U16116 (N_16116,N_14591,N_14398);
xnor U16117 (N_16117,N_13866,N_14661);
nor U16118 (N_16118,N_14823,N_14900);
or U16119 (N_16119,N_13676,N_14894);
nand U16120 (N_16120,N_14392,N_13688);
nor U16121 (N_16121,N_14357,N_14431);
nor U16122 (N_16122,N_13994,N_14104);
nand U16123 (N_16123,N_14977,N_13868);
and U16124 (N_16124,N_14872,N_14515);
xnor U16125 (N_16125,N_14988,N_14520);
and U16126 (N_16126,N_14701,N_13836);
or U16127 (N_16127,N_13756,N_14092);
or U16128 (N_16128,N_14297,N_14733);
nand U16129 (N_16129,N_14105,N_14633);
and U16130 (N_16130,N_14370,N_14075);
xnor U16131 (N_16131,N_14162,N_14663);
and U16132 (N_16132,N_14053,N_14420);
and U16133 (N_16133,N_14726,N_14959);
and U16134 (N_16134,N_13739,N_14937);
nand U16135 (N_16135,N_14925,N_13683);
nand U16136 (N_16136,N_14708,N_14472);
or U16137 (N_16137,N_13770,N_14547);
xor U16138 (N_16138,N_14931,N_14348);
xnor U16139 (N_16139,N_14459,N_13562);
and U16140 (N_16140,N_14699,N_14716);
and U16141 (N_16141,N_14116,N_14358);
xnor U16142 (N_16142,N_13516,N_13512);
xor U16143 (N_16143,N_13591,N_13655);
nand U16144 (N_16144,N_13749,N_14051);
nand U16145 (N_16145,N_14486,N_13546);
nand U16146 (N_16146,N_14083,N_13585);
and U16147 (N_16147,N_13808,N_14193);
nor U16148 (N_16148,N_13837,N_14163);
nor U16149 (N_16149,N_13986,N_13536);
and U16150 (N_16150,N_13614,N_14212);
and U16151 (N_16151,N_14015,N_13552);
and U16152 (N_16152,N_13773,N_14702);
nand U16153 (N_16153,N_13730,N_14618);
nand U16154 (N_16154,N_13836,N_14321);
or U16155 (N_16155,N_13975,N_14461);
xor U16156 (N_16156,N_14632,N_14274);
and U16157 (N_16157,N_14074,N_14795);
nor U16158 (N_16158,N_14594,N_14890);
xnor U16159 (N_16159,N_13580,N_14232);
nand U16160 (N_16160,N_13854,N_14672);
and U16161 (N_16161,N_14300,N_14468);
xnor U16162 (N_16162,N_14668,N_14990);
or U16163 (N_16163,N_14558,N_14870);
xnor U16164 (N_16164,N_14857,N_14443);
nor U16165 (N_16165,N_14645,N_14631);
nor U16166 (N_16166,N_13837,N_14943);
and U16167 (N_16167,N_14060,N_14593);
nand U16168 (N_16168,N_14793,N_13800);
and U16169 (N_16169,N_13923,N_14818);
xnor U16170 (N_16170,N_13656,N_14537);
nor U16171 (N_16171,N_14361,N_14525);
or U16172 (N_16172,N_14808,N_14786);
and U16173 (N_16173,N_13770,N_14177);
or U16174 (N_16174,N_14228,N_14100);
and U16175 (N_16175,N_13900,N_14564);
and U16176 (N_16176,N_14808,N_13733);
nor U16177 (N_16177,N_13883,N_14991);
and U16178 (N_16178,N_13587,N_14937);
or U16179 (N_16179,N_14325,N_14168);
nor U16180 (N_16180,N_14487,N_14785);
nand U16181 (N_16181,N_14571,N_14356);
xnor U16182 (N_16182,N_13536,N_13522);
or U16183 (N_16183,N_13686,N_14109);
nand U16184 (N_16184,N_14641,N_14029);
or U16185 (N_16185,N_14502,N_14862);
xor U16186 (N_16186,N_14107,N_14426);
nand U16187 (N_16187,N_14647,N_13585);
nand U16188 (N_16188,N_14064,N_14718);
nand U16189 (N_16189,N_13948,N_14412);
or U16190 (N_16190,N_14803,N_13617);
nor U16191 (N_16191,N_14074,N_13903);
nand U16192 (N_16192,N_14689,N_14127);
nand U16193 (N_16193,N_13943,N_14007);
xnor U16194 (N_16194,N_14100,N_13974);
xnor U16195 (N_16195,N_14460,N_14602);
nor U16196 (N_16196,N_14939,N_13725);
nor U16197 (N_16197,N_13681,N_14622);
nand U16198 (N_16198,N_14570,N_14991);
and U16199 (N_16199,N_13864,N_14648);
nand U16200 (N_16200,N_14324,N_14604);
or U16201 (N_16201,N_13964,N_14827);
nand U16202 (N_16202,N_14363,N_14265);
nand U16203 (N_16203,N_14712,N_14870);
nor U16204 (N_16204,N_14350,N_13720);
xor U16205 (N_16205,N_13895,N_13590);
xnor U16206 (N_16206,N_13535,N_13794);
or U16207 (N_16207,N_13696,N_13792);
and U16208 (N_16208,N_14324,N_14968);
nand U16209 (N_16209,N_14194,N_14520);
xnor U16210 (N_16210,N_13925,N_14894);
and U16211 (N_16211,N_14192,N_14376);
or U16212 (N_16212,N_13998,N_13987);
nor U16213 (N_16213,N_14630,N_13795);
nand U16214 (N_16214,N_14542,N_14179);
nor U16215 (N_16215,N_13961,N_14445);
nand U16216 (N_16216,N_13524,N_14422);
xnor U16217 (N_16217,N_13748,N_14992);
xor U16218 (N_16218,N_14462,N_13743);
nor U16219 (N_16219,N_14181,N_14594);
xor U16220 (N_16220,N_13575,N_14962);
xor U16221 (N_16221,N_14334,N_14208);
and U16222 (N_16222,N_14700,N_13976);
and U16223 (N_16223,N_14353,N_13836);
nor U16224 (N_16224,N_14126,N_14628);
nand U16225 (N_16225,N_14085,N_13915);
or U16226 (N_16226,N_14416,N_14800);
and U16227 (N_16227,N_14490,N_14587);
and U16228 (N_16228,N_14401,N_13961);
and U16229 (N_16229,N_14473,N_13950);
nor U16230 (N_16230,N_14737,N_14829);
or U16231 (N_16231,N_14082,N_13809);
and U16232 (N_16232,N_14985,N_13616);
nand U16233 (N_16233,N_14316,N_14968);
nor U16234 (N_16234,N_14794,N_14484);
nor U16235 (N_16235,N_14683,N_14533);
nand U16236 (N_16236,N_14761,N_13639);
or U16237 (N_16237,N_13676,N_14581);
nor U16238 (N_16238,N_13933,N_14608);
or U16239 (N_16239,N_13588,N_14779);
xnor U16240 (N_16240,N_14792,N_14712);
xnor U16241 (N_16241,N_13840,N_14357);
or U16242 (N_16242,N_14233,N_14666);
nand U16243 (N_16243,N_14019,N_14378);
and U16244 (N_16244,N_14337,N_14808);
nor U16245 (N_16245,N_13929,N_14136);
nor U16246 (N_16246,N_14186,N_14325);
xor U16247 (N_16247,N_13607,N_14689);
xnor U16248 (N_16248,N_14006,N_13851);
nand U16249 (N_16249,N_14780,N_14222);
xor U16250 (N_16250,N_14356,N_13825);
nor U16251 (N_16251,N_14108,N_14485);
nand U16252 (N_16252,N_13608,N_14327);
xor U16253 (N_16253,N_14921,N_13704);
xnor U16254 (N_16254,N_14880,N_14864);
nand U16255 (N_16255,N_14297,N_13885);
xnor U16256 (N_16256,N_14647,N_14510);
or U16257 (N_16257,N_14614,N_14276);
and U16258 (N_16258,N_13663,N_14070);
nor U16259 (N_16259,N_14584,N_14158);
or U16260 (N_16260,N_14260,N_14621);
nor U16261 (N_16261,N_14290,N_14341);
and U16262 (N_16262,N_13591,N_14062);
xor U16263 (N_16263,N_14195,N_14819);
or U16264 (N_16264,N_13573,N_13729);
nor U16265 (N_16265,N_14405,N_14763);
xor U16266 (N_16266,N_14887,N_14125);
xnor U16267 (N_16267,N_14367,N_13980);
nor U16268 (N_16268,N_13784,N_13582);
and U16269 (N_16269,N_14650,N_14460);
nand U16270 (N_16270,N_14002,N_13814);
xor U16271 (N_16271,N_13860,N_14525);
or U16272 (N_16272,N_13656,N_13504);
nor U16273 (N_16273,N_14313,N_13736);
xor U16274 (N_16274,N_14095,N_13630);
and U16275 (N_16275,N_13640,N_14111);
and U16276 (N_16276,N_13660,N_14667);
nand U16277 (N_16277,N_13959,N_14204);
and U16278 (N_16278,N_14094,N_14447);
xor U16279 (N_16279,N_13910,N_13977);
or U16280 (N_16280,N_14139,N_13990);
nor U16281 (N_16281,N_13517,N_14646);
xor U16282 (N_16282,N_14991,N_14752);
nand U16283 (N_16283,N_14076,N_14657);
nor U16284 (N_16284,N_14763,N_14881);
nand U16285 (N_16285,N_14921,N_14877);
or U16286 (N_16286,N_13553,N_14076);
nor U16287 (N_16287,N_14841,N_13516);
xor U16288 (N_16288,N_14239,N_14954);
or U16289 (N_16289,N_13589,N_14496);
xnor U16290 (N_16290,N_13852,N_13620);
xnor U16291 (N_16291,N_13738,N_14383);
nand U16292 (N_16292,N_14947,N_14966);
and U16293 (N_16293,N_13712,N_13770);
and U16294 (N_16294,N_13504,N_13589);
nand U16295 (N_16295,N_14572,N_14047);
nor U16296 (N_16296,N_14296,N_14971);
nand U16297 (N_16297,N_14380,N_13659);
nand U16298 (N_16298,N_13925,N_14167);
and U16299 (N_16299,N_13647,N_13818);
nor U16300 (N_16300,N_14977,N_13676);
nand U16301 (N_16301,N_14846,N_13529);
nor U16302 (N_16302,N_13673,N_13912);
and U16303 (N_16303,N_14183,N_14185);
nor U16304 (N_16304,N_13758,N_14446);
or U16305 (N_16305,N_14559,N_14583);
xnor U16306 (N_16306,N_13501,N_14429);
nor U16307 (N_16307,N_13532,N_14090);
nand U16308 (N_16308,N_13534,N_14624);
or U16309 (N_16309,N_14366,N_13635);
and U16310 (N_16310,N_14419,N_14203);
or U16311 (N_16311,N_14732,N_14069);
nor U16312 (N_16312,N_13984,N_14908);
or U16313 (N_16313,N_13514,N_13513);
or U16314 (N_16314,N_14062,N_14754);
nand U16315 (N_16315,N_13697,N_14239);
or U16316 (N_16316,N_14154,N_14927);
or U16317 (N_16317,N_14147,N_14968);
nand U16318 (N_16318,N_13607,N_14149);
and U16319 (N_16319,N_14943,N_13719);
nand U16320 (N_16320,N_14980,N_14715);
or U16321 (N_16321,N_13630,N_13670);
nand U16322 (N_16322,N_13598,N_13644);
nor U16323 (N_16323,N_13902,N_13747);
xnor U16324 (N_16324,N_13986,N_14071);
and U16325 (N_16325,N_13644,N_14503);
and U16326 (N_16326,N_14049,N_13753);
or U16327 (N_16327,N_14157,N_13578);
xnor U16328 (N_16328,N_14824,N_14486);
nor U16329 (N_16329,N_14838,N_14377);
nand U16330 (N_16330,N_13600,N_14200);
nand U16331 (N_16331,N_13614,N_14283);
xor U16332 (N_16332,N_14833,N_14682);
or U16333 (N_16333,N_14828,N_14157);
or U16334 (N_16334,N_13507,N_14411);
nand U16335 (N_16335,N_13644,N_14025);
nor U16336 (N_16336,N_14506,N_13524);
nor U16337 (N_16337,N_14034,N_13933);
and U16338 (N_16338,N_13974,N_14054);
xor U16339 (N_16339,N_14934,N_14925);
xnor U16340 (N_16340,N_13626,N_13910);
nand U16341 (N_16341,N_14880,N_14798);
or U16342 (N_16342,N_14011,N_14440);
nor U16343 (N_16343,N_13519,N_14438);
nor U16344 (N_16344,N_13538,N_14073);
nand U16345 (N_16345,N_14067,N_13922);
and U16346 (N_16346,N_14772,N_14419);
nand U16347 (N_16347,N_14172,N_14377);
and U16348 (N_16348,N_13803,N_13975);
and U16349 (N_16349,N_14896,N_14445);
and U16350 (N_16350,N_14413,N_14516);
and U16351 (N_16351,N_14719,N_14758);
xnor U16352 (N_16352,N_13636,N_14216);
nor U16353 (N_16353,N_13869,N_14066);
nor U16354 (N_16354,N_13934,N_14906);
nand U16355 (N_16355,N_13558,N_13897);
and U16356 (N_16356,N_14193,N_13812);
and U16357 (N_16357,N_14260,N_13794);
xor U16358 (N_16358,N_14844,N_14529);
and U16359 (N_16359,N_14569,N_14493);
nor U16360 (N_16360,N_14730,N_14399);
xor U16361 (N_16361,N_14838,N_14572);
xor U16362 (N_16362,N_14439,N_13799);
and U16363 (N_16363,N_14101,N_14067);
or U16364 (N_16364,N_14569,N_14725);
xor U16365 (N_16365,N_14770,N_14708);
and U16366 (N_16366,N_14303,N_13727);
and U16367 (N_16367,N_13999,N_14063);
xor U16368 (N_16368,N_14775,N_14286);
nor U16369 (N_16369,N_14721,N_14149);
xor U16370 (N_16370,N_14331,N_14536);
xor U16371 (N_16371,N_13651,N_14772);
xor U16372 (N_16372,N_13735,N_14897);
and U16373 (N_16373,N_13562,N_13823);
xor U16374 (N_16374,N_14278,N_14745);
nor U16375 (N_16375,N_14527,N_14618);
xnor U16376 (N_16376,N_14456,N_14540);
nor U16377 (N_16377,N_13691,N_13849);
nand U16378 (N_16378,N_13504,N_14130);
and U16379 (N_16379,N_14915,N_13907);
or U16380 (N_16380,N_13718,N_14372);
nand U16381 (N_16381,N_13691,N_14230);
nand U16382 (N_16382,N_14913,N_13537);
and U16383 (N_16383,N_13901,N_14493);
nor U16384 (N_16384,N_13686,N_13567);
xor U16385 (N_16385,N_14340,N_14199);
nand U16386 (N_16386,N_14262,N_14309);
and U16387 (N_16387,N_14254,N_13865);
nand U16388 (N_16388,N_14742,N_13851);
nand U16389 (N_16389,N_14625,N_14973);
xnor U16390 (N_16390,N_13888,N_13995);
xnor U16391 (N_16391,N_14773,N_14041);
xor U16392 (N_16392,N_14505,N_14341);
or U16393 (N_16393,N_14057,N_14455);
or U16394 (N_16394,N_14582,N_14523);
nand U16395 (N_16395,N_14486,N_14722);
xor U16396 (N_16396,N_14886,N_14573);
nor U16397 (N_16397,N_13974,N_14511);
xnor U16398 (N_16398,N_13652,N_14908);
nor U16399 (N_16399,N_13661,N_14387);
or U16400 (N_16400,N_13853,N_14969);
nor U16401 (N_16401,N_13951,N_13964);
xnor U16402 (N_16402,N_13956,N_14564);
nand U16403 (N_16403,N_13761,N_14963);
nand U16404 (N_16404,N_13624,N_13843);
or U16405 (N_16405,N_13715,N_14366);
xor U16406 (N_16406,N_14809,N_14745);
nor U16407 (N_16407,N_13904,N_13796);
nor U16408 (N_16408,N_14783,N_14360);
nand U16409 (N_16409,N_13969,N_14508);
xnor U16410 (N_16410,N_14426,N_14994);
and U16411 (N_16411,N_14063,N_14123);
and U16412 (N_16412,N_14171,N_14189);
nor U16413 (N_16413,N_14322,N_14529);
and U16414 (N_16414,N_13982,N_13861);
nor U16415 (N_16415,N_14714,N_14005);
nand U16416 (N_16416,N_14616,N_14622);
nor U16417 (N_16417,N_14145,N_14931);
nand U16418 (N_16418,N_14315,N_14740);
nand U16419 (N_16419,N_14652,N_14630);
or U16420 (N_16420,N_13809,N_13690);
nand U16421 (N_16421,N_14220,N_13830);
xnor U16422 (N_16422,N_13566,N_14683);
or U16423 (N_16423,N_14576,N_14160);
and U16424 (N_16424,N_13892,N_13962);
nand U16425 (N_16425,N_14158,N_14446);
nand U16426 (N_16426,N_13663,N_13979);
and U16427 (N_16427,N_13776,N_14328);
nand U16428 (N_16428,N_13976,N_13543);
or U16429 (N_16429,N_14446,N_13621);
or U16430 (N_16430,N_13606,N_13755);
nand U16431 (N_16431,N_14292,N_14983);
or U16432 (N_16432,N_13649,N_13716);
or U16433 (N_16433,N_14442,N_14319);
or U16434 (N_16434,N_13567,N_14480);
nand U16435 (N_16435,N_14946,N_14405);
and U16436 (N_16436,N_14772,N_13940);
nor U16437 (N_16437,N_13748,N_14944);
xnor U16438 (N_16438,N_13801,N_14272);
and U16439 (N_16439,N_14976,N_13544);
nor U16440 (N_16440,N_14660,N_13871);
and U16441 (N_16441,N_14449,N_14885);
nor U16442 (N_16442,N_14071,N_14977);
or U16443 (N_16443,N_14642,N_14425);
and U16444 (N_16444,N_13623,N_14825);
xnor U16445 (N_16445,N_14446,N_14761);
or U16446 (N_16446,N_13664,N_14958);
xnor U16447 (N_16447,N_14607,N_14134);
nor U16448 (N_16448,N_13619,N_14136);
xor U16449 (N_16449,N_13888,N_14478);
and U16450 (N_16450,N_13764,N_14452);
and U16451 (N_16451,N_14279,N_13950);
nand U16452 (N_16452,N_13878,N_13811);
xnor U16453 (N_16453,N_13802,N_14102);
nor U16454 (N_16454,N_14659,N_14833);
or U16455 (N_16455,N_13514,N_14216);
nand U16456 (N_16456,N_13562,N_14692);
xor U16457 (N_16457,N_13645,N_14680);
xor U16458 (N_16458,N_13935,N_14422);
nand U16459 (N_16459,N_13926,N_14383);
and U16460 (N_16460,N_14897,N_14301);
nand U16461 (N_16461,N_13782,N_13722);
nand U16462 (N_16462,N_14767,N_14061);
xor U16463 (N_16463,N_13827,N_14800);
or U16464 (N_16464,N_14916,N_14779);
and U16465 (N_16465,N_14723,N_14704);
nand U16466 (N_16466,N_13934,N_13966);
nor U16467 (N_16467,N_14178,N_13827);
nand U16468 (N_16468,N_14194,N_14567);
and U16469 (N_16469,N_13909,N_14452);
nor U16470 (N_16470,N_13606,N_13677);
xnor U16471 (N_16471,N_14345,N_14599);
nand U16472 (N_16472,N_13832,N_14471);
xnor U16473 (N_16473,N_13893,N_13862);
or U16474 (N_16474,N_14028,N_13534);
and U16475 (N_16475,N_14012,N_13751);
nand U16476 (N_16476,N_13645,N_14943);
nor U16477 (N_16477,N_14517,N_14232);
and U16478 (N_16478,N_14727,N_13610);
nand U16479 (N_16479,N_14069,N_14116);
and U16480 (N_16480,N_13650,N_13958);
and U16481 (N_16481,N_13665,N_14886);
and U16482 (N_16482,N_13566,N_13902);
or U16483 (N_16483,N_14065,N_14296);
nor U16484 (N_16484,N_13748,N_13663);
nand U16485 (N_16485,N_13713,N_14427);
nand U16486 (N_16486,N_13658,N_14768);
or U16487 (N_16487,N_14035,N_13980);
nand U16488 (N_16488,N_13996,N_14176);
nor U16489 (N_16489,N_14756,N_13719);
nand U16490 (N_16490,N_14337,N_14373);
nor U16491 (N_16491,N_13915,N_13919);
nor U16492 (N_16492,N_13615,N_14755);
and U16493 (N_16493,N_14182,N_14559);
xor U16494 (N_16494,N_14944,N_14317);
nor U16495 (N_16495,N_13570,N_14532);
nor U16496 (N_16496,N_14280,N_14243);
nor U16497 (N_16497,N_14759,N_14235);
nor U16498 (N_16498,N_14407,N_14204);
nor U16499 (N_16499,N_14228,N_14639);
nor U16500 (N_16500,N_16132,N_16232);
nand U16501 (N_16501,N_15230,N_15849);
or U16502 (N_16502,N_15876,N_16116);
or U16503 (N_16503,N_15620,N_15551);
or U16504 (N_16504,N_16380,N_16356);
nor U16505 (N_16505,N_15441,N_15522);
and U16506 (N_16506,N_16076,N_16145);
nand U16507 (N_16507,N_15310,N_15650);
or U16508 (N_16508,N_15611,N_16150);
nor U16509 (N_16509,N_16174,N_16233);
and U16510 (N_16510,N_16276,N_15332);
nand U16511 (N_16511,N_15245,N_16321);
nor U16512 (N_16512,N_15878,N_15300);
xnor U16513 (N_16513,N_15739,N_15419);
or U16514 (N_16514,N_15277,N_15690);
or U16515 (N_16515,N_15965,N_15284);
nand U16516 (N_16516,N_16400,N_16399);
nand U16517 (N_16517,N_15854,N_16240);
nor U16518 (N_16518,N_15773,N_16197);
nand U16519 (N_16519,N_15409,N_16191);
nand U16520 (N_16520,N_16318,N_15774);
nand U16521 (N_16521,N_16015,N_16242);
nand U16522 (N_16522,N_15320,N_15346);
and U16523 (N_16523,N_16139,N_16391);
and U16524 (N_16524,N_16311,N_15660);
xor U16525 (N_16525,N_16325,N_15406);
nand U16526 (N_16526,N_15543,N_15555);
nor U16527 (N_16527,N_15973,N_15116);
xnor U16528 (N_16528,N_16433,N_15343);
or U16529 (N_16529,N_15323,N_16342);
xor U16530 (N_16530,N_15192,N_15266);
or U16531 (N_16531,N_16291,N_15338);
nor U16532 (N_16532,N_16450,N_15091);
or U16533 (N_16533,N_15162,N_15279);
nand U16534 (N_16534,N_15259,N_16292);
nand U16535 (N_16535,N_15122,N_16498);
or U16536 (N_16536,N_15499,N_15726);
and U16537 (N_16537,N_16331,N_15354);
and U16538 (N_16538,N_16141,N_15313);
nor U16539 (N_16539,N_16268,N_15483);
and U16540 (N_16540,N_16146,N_15949);
and U16541 (N_16541,N_15516,N_15582);
or U16542 (N_16542,N_15943,N_15901);
xnor U16543 (N_16543,N_15378,N_15534);
xor U16544 (N_16544,N_15857,N_15956);
nand U16545 (N_16545,N_16248,N_16102);
xnor U16546 (N_16546,N_16396,N_16065);
and U16547 (N_16547,N_15256,N_15570);
xor U16548 (N_16548,N_15134,N_15634);
and U16549 (N_16549,N_15141,N_15584);
xnor U16550 (N_16550,N_15655,N_16209);
nor U16551 (N_16551,N_15271,N_16219);
nand U16552 (N_16552,N_16206,N_16029);
nand U16553 (N_16553,N_15238,N_16130);
nor U16554 (N_16554,N_15561,N_15251);
and U16555 (N_16555,N_15647,N_15940);
nand U16556 (N_16556,N_15178,N_15540);
xor U16557 (N_16557,N_16301,N_16364);
nand U16558 (N_16558,N_15765,N_15776);
and U16559 (N_16559,N_15485,N_15128);
or U16560 (N_16560,N_15491,N_16290);
nor U16561 (N_16561,N_15045,N_15903);
or U16562 (N_16562,N_16459,N_15113);
xnor U16563 (N_16563,N_15403,N_16460);
xor U16564 (N_16564,N_16271,N_15630);
nor U16565 (N_16565,N_16363,N_15865);
or U16566 (N_16566,N_15598,N_16479);
nand U16567 (N_16567,N_15775,N_16448);
nand U16568 (N_16568,N_15923,N_15741);
xnor U16569 (N_16569,N_15109,N_16135);
nor U16570 (N_16570,N_15674,N_15010);
and U16571 (N_16571,N_15467,N_15411);
nor U16572 (N_16572,N_15732,N_15131);
nor U16573 (N_16573,N_15846,N_15575);
nor U16574 (N_16574,N_15676,N_16062);
nor U16575 (N_16575,N_15100,N_15526);
nand U16576 (N_16576,N_15695,N_16298);
or U16577 (N_16577,N_15054,N_15662);
or U16578 (N_16578,N_15760,N_16078);
and U16579 (N_16579,N_15050,N_16402);
nand U16580 (N_16580,N_15175,N_15214);
xnor U16581 (N_16581,N_15980,N_15104);
and U16582 (N_16582,N_15476,N_15188);
nand U16583 (N_16583,N_16277,N_16004);
nor U16584 (N_16584,N_15914,N_15318);
and U16585 (N_16585,N_15426,N_15077);
nor U16586 (N_16586,N_15324,N_15458);
nor U16587 (N_16587,N_16368,N_15623);
nor U16588 (N_16588,N_16072,N_15282);
nand U16589 (N_16589,N_16208,N_16243);
and U16590 (N_16590,N_16317,N_15288);
xor U16591 (N_16591,N_15585,N_16278);
nand U16592 (N_16592,N_16495,N_15811);
xor U16593 (N_16593,N_15112,N_15766);
nor U16594 (N_16594,N_15734,N_15761);
and U16595 (N_16595,N_15533,N_16079);
nand U16596 (N_16596,N_15462,N_15799);
nand U16597 (N_16597,N_16234,N_15843);
nand U16598 (N_16598,N_15578,N_15442);
nand U16599 (N_16599,N_15405,N_15964);
or U16600 (N_16600,N_16121,N_15912);
xor U16601 (N_16601,N_16251,N_16198);
nor U16602 (N_16602,N_15201,N_15853);
and U16603 (N_16603,N_16172,N_15357);
nor U16604 (N_16604,N_16069,N_15363);
and U16605 (N_16605,N_15446,N_15482);
xor U16606 (N_16606,N_15142,N_16404);
and U16607 (N_16607,N_15506,N_16073);
nor U16608 (N_16608,N_15029,N_15339);
nor U16609 (N_16609,N_15212,N_16403);
nor U16610 (N_16610,N_15168,N_16094);
xnor U16611 (N_16611,N_15422,N_15280);
nor U16612 (N_16612,N_16068,N_16293);
nand U16613 (N_16613,N_16047,N_15750);
xnor U16614 (N_16614,N_15012,N_15831);
xnor U16615 (N_16615,N_15334,N_15631);
and U16616 (N_16616,N_15132,N_15538);
nand U16617 (N_16617,N_15547,N_15869);
nand U16618 (N_16618,N_15353,N_15167);
or U16619 (N_16619,N_15082,N_16468);
nand U16620 (N_16620,N_15769,N_15718);
and U16621 (N_16621,N_15033,N_15093);
nand U16622 (N_16622,N_16222,N_15215);
or U16623 (N_16623,N_16417,N_16114);
or U16624 (N_16624,N_15840,N_15920);
xnor U16625 (N_16625,N_15566,N_15730);
and U16626 (N_16626,N_15402,N_15152);
and U16627 (N_16627,N_15759,N_16013);
and U16628 (N_16628,N_15355,N_15145);
xnor U16629 (N_16629,N_15392,N_15687);
and U16630 (N_16630,N_16085,N_15124);
and U16631 (N_16631,N_15548,N_15723);
or U16632 (N_16632,N_15706,N_15821);
xor U16633 (N_16633,N_16118,N_15616);
nand U16634 (N_16634,N_15729,N_15042);
and U16635 (N_16635,N_16453,N_15580);
or U16636 (N_16636,N_15743,N_16335);
nand U16637 (N_16637,N_15569,N_16482);
nor U16638 (N_16638,N_15546,N_15997);
xor U16639 (N_16639,N_15470,N_15244);
xor U16640 (N_16640,N_15413,N_16412);
nor U16641 (N_16641,N_16049,N_16185);
xor U16642 (N_16642,N_15816,N_15902);
and U16643 (N_16643,N_15782,N_15797);
or U16644 (N_16644,N_15269,N_15000);
nand U16645 (N_16645,N_16186,N_16159);
nand U16646 (N_16646,N_15897,N_15531);
xor U16647 (N_16647,N_15407,N_15672);
nand U16648 (N_16648,N_16218,N_16398);
nor U16649 (N_16649,N_15438,N_15423);
nor U16650 (N_16650,N_16048,N_15473);
nand U16651 (N_16651,N_15263,N_16456);
nor U16652 (N_16652,N_15233,N_16432);
nor U16653 (N_16653,N_15250,N_15958);
xor U16654 (N_16654,N_16452,N_15115);
nor U16655 (N_16655,N_15254,N_15733);
xor U16656 (N_16656,N_15607,N_15500);
nand U16657 (N_16657,N_15767,N_15264);
nor U16658 (N_16658,N_15437,N_15589);
xnor U16659 (N_16659,N_15118,N_16389);
xnor U16660 (N_16660,N_16143,N_15989);
or U16661 (N_16661,N_16044,N_15048);
xnor U16662 (N_16662,N_15410,N_15779);
nor U16663 (N_16663,N_15833,N_16093);
or U16664 (N_16664,N_15475,N_15839);
xor U16665 (N_16665,N_16095,N_16151);
nand U16666 (N_16666,N_16499,N_15879);
nor U16667 (N_16667,N_16435,N_16211);
or U16668 (N_16668,N_15632,N_16046);
and U16669 (N_16669,N_15868,N_15636);
and U16670 (N_16670,N_15993,N_16273);
and U16671 (N_16671,N_15751,N_15460);
or U16672 (N_16672,N_16312,N_15837);
xor U16673 (N_16673,N_16051,N_15796);
and U16674 (N_16674,N_16324,N_15536);
nand U16675 (N_16675,N_15348,N_15183);
nor U16676 (N_16676,N_15702,N_15891);
xor U16677 (N_16677,N_15040,N_16147);
and U16678 (N_16678,N_16226,N_15758);
nand U16679 (N_16679,N_15260,N_15870);
or U16680 (N_16680,N_16279,N_15521);
xor U16681 (N_16681,N_16465,N_16036);
or U16682 (N_16682,N_15638,N_16425);
xnor U16683 (N_16683,N_15179,N_15014);
nand U16684 (N_16684,N_15713,N_16107);
and U16685 (N_16685,N_16012,N_15977);
xor U16686 (N_16686,N_15968,N_15641);
or U16687 (N_16687,N_15421,N_16264);
nor U16688 (N_16688,N_15311,N_16039);
xor U16689 (N_16689,N_15568,N_15424);
or U16690 (N_16690,N_15369,N_16199);
and U16691 (N_16691,N_16351,N_15668);
and U16692 (N_16692,N_15382,N_15390);
xnor U16693 (N_16693,N_15295,N_15185);
or U16694 (N_16694,N_15812,N_15916);
and U16695 (N_16695,N_16481,N_16131);
nand U16696 (N_16696,N_15592,N_16379);
and U16697 (N_16697,N_16451,N_16006);
nand U16698 (N_16698,N_15314,N_15972);
or U16699 (N_16699,N_15858,N_16386);
nand U16700 (N_16700,N_16097,N_16122);
or U16701 (N_16701,N_15756,N_16269);
nand U16702 (N_16702,N_15350,N_15140);
and U16703 (N_16703,N_15125,N_15560);
nor U16704 (N_16704,N_16415,N_15747);
or U16705 (N_16705,N_15149,N_16144);
nand U16706 (N_16706,N_15608,N_16314);
nor U16707 (N_16707,N_15213,N_16326);
and U16708 (N_16708,N_16419,N_16464);
or U16709 (N_16709,N_15567,N_15810);
or U16710 (N_16710,N_15319,N_15825);
nand U16711 (N_16711,N_16098,N_16252);
or U16712 (N_16712,N_16173,N_16244);
xnor U16713 (N_16713,N_16024,N_15487);
or U16714 (N_16714,N_15067,N_15105);
nor U16715 (N_16715,N_15925,N_16421);
nand U16716 (N_16716,N_15177,N_15190);
and U16717 (N_16717,N_16125,N_15015);
and U16718 (N_16718,N_15737,N_15193);
nand U16719 (N_16719,N_15326,N_16050);
or U16720 (N_16720,N_16469,N_15913);
nand U16721 (N_16721,N_15789,N_16087);
nor U16722 (N_16722,N_15978,N_15746);
and U16723 (N_16723,N_16408,N_15283);
or U16724 (N_16724,N_15685,N_15621);
and U16725 (N_16725,N_16103,N_15996);
nor U16726 (N_16726,N_16307,N_15671);
nand U16727 (N_16727,N_15241,N_15712);
or U16728 (N_16728,N_16349,N_15614);
or U16729 (N_16729,N_16040,N_15772);
or U16730 (N_16730,N_15023,N_15497);
or U16731 (N_16731,N_15204,N_16213);
nand U16732 (N_16732,N_15165,N_16395);
nor U16733 (N_16733,N_15838,N_15880);
and U16734 (N_16734,N_16165,N_15006);
xor U16735 (N_16735,N_16203,N_16035);
or U16736 (N_16736,N_15449,N_15160);
and U16737 (N_16737,N_15342,N_15762);
and U16738 (N_16738,N_16330,N_15684);
nor U16739 (N_16739,N_16045,N_16060);
xnor U16740 (N_16740,N_15911,N_16055);
xnor U16741 (N_16741,N_16176,N_16353);
xnor U16742 (N_16742,N_15716,N_16362);
nor U16743 (N_16743,N_15217,N_15080);
nand U16744 (N_16744,N_15594,N_16295);
and U16745 (N_16745,N_16148,N_15290);
xnor U16746 (N_16746,N_15558,N_15975);
or U16747 (N_16747,N_15976,N_16101);
xor U16748 (N_16748,N_16322,N_15076);
nand U16749 (N_16749,N_16250,N_15520);
nand U16750 (N_16750,N_16205,N_15133);
nand U16751 (N_16751,N_15863,N_16091);
nand U16752 (N_16752,N_16470,N_16265);
nor U16753 (N_16753,N_16308,N_15929);
xnor U16754 (N_16754,N_15532,N_16200);
nand U16755 (N_16755,N_16007,N_16296);
and U16756 (N_16756,N_15866,N_15087);
or U16757 (N_16757,N_15699,N_15347);
nand U16758 (N_16758,N_15220,N_15439);
xnor U16759 (N_16759,N_15431,N_15110);
nand U16760 (N_16760,N_16299,N_15794);
nor U16761 (N_16761,N_15399,N_15917);
nor U16762 (N_16762,N_16297,N_15709);
and U16763 (N_16763,N_15302,N_15447);
xor U16764 (N_16764,N_16134,N_15844);
or U16765 (N_16765,N_16410,N_15479);
nor U16766 (N_16766,N_15951,N_15457);
xor U16767 (N_16767,N_16361,N_16347);
and U16768 (N_16768,N_15325,N_16074);
nand U16769 (N_16769,N_16009,N_15053);
nor U16770 (N_16770,N_15824,N_15386);
or U16771 (N_16771,N_16155,N_15604);
xnor U16772 (N_16772,N_15221,N_16057);
nor U16773 (N_16773,N_16056,N_15166);
nand U16774 (N_16774,N_15025,N_16424);
or U16775 (N_16775,N_15539,N_15564);
or U16776 (N_16776,N_16043,N_15315);
or U16777 (N_16777,N_16328,N_15478);
xor U16778 (N_16778,N_15804,N_15096);
nor U16779 (N_16779,N_15574,N_15512);
nand U16780 (N_16780,N_15807,N_15187);
xnor U16781 (N_16781,N_15159,N_15389);
and U16782 (N_16782,N_15545,N_15523);
or U16783 (N_16783,N_15253,N_16315);
or U16784 (N_16784,N_15967,N_15947);
xor U16785 (N_16785,N_15686,N_15344);
or U16786 (N_16786,N_16111,N_15137);
nand U16787 (N_16787,N_15802,N_15306);
nor U16788 (N_16788,N_15101,N_15586);
xnor U16789 (N_16789,N_15654,N_16027);
or U16790 (N_16790,N_16332,N_15404);
nor U16791 (N_16791,N_15908,N_15186);
xnor U16792 (N_16792,N_15194,N_16287);
nand U16793 (N_16793,N_15525,N_15021);
xor U16794 (N_16794,N_15652,N_16017);
xnor U16795 (N_16795,N_15845,N_16346);
xor U16796 (N_16796,N_15366,N_15697);
xor U16797 (N_16797,N_15541,N_16323);
xor U16798 (N_16798,N_15609,N_15107);
nand U16799 (N_16799,N_16231,N_15725);
nor U16800 (N_16800,N_16449,N_15896);
or U16801 (N_16801,N_16397,N_16104);
xnor U16802 (N_16802,N_15031,N_15368);
nand U16803 (N_16803,N_15888,N_16042);
nor U16804 (N_16804,N_15835,N_16071);
and U16805 (N_16805,N_15717,N_15679);
or U16806 (N_16806,N_16423,N_15017);
and U16807 (N_16807,N_15139,N_15498);
nor U16808 (N_16808,N_15795,N_16373);
nor U16809 (N_16809,N_15991,N_16457);
xor U16810 (N_16810,N_15784,N_16466);
nor U16811 (N_16811,N_15603,N_15657);
nor U16812 (N_16812,N_15164,N_15452);
or U16813 (N_16813,N_15983,N_15384);
nand U16814 (N_16814,N_15433,N_15090);
and U16815 (N_16815,N_15553,N_16088);
or U16816 (N_16816,N_16003,N_15905);
xor U16817 (N_16817,N_15352,N_16136);
xor U16818 (N_16818,N_16154,N_15819);
xor U16819 (N_16819,N_16261,N_16434);
nand U16820 (N_16820,N_15704,N_16305);
nor U16821 (N_16821,N_15815,N_15581);
xnor U16822 (N_16822,N_16089,N_16306);
nor U16823 (N_16823,N_15335,N_15544);
and U16824 (N_16824,N_15084,N_15692);
xor U16825 (N_16825,N_15788,N_16262);
nand U16826 (N_16826,N_15918,N_15727);
or U16827 (N_16827,N_15554,N_16018);
nand U16828 (N_16828,N_15872,N_16021);
or U16829 (N_16829,N_16140,N_15337);
or U16830 (N_16830,N_16249,N_16184);
nand U16831 (N_16831,N_15875,N_16192);
nand U16832 (N_16832,N_16375,N_15443);
xnor U16833 (N_16833,N_15229,N_15207);
xor U16834 (N_16834,N_15184,N_16216);
and U16835 (N_16835,N_16281,N_15262);
nand U16836 (N_16836,N_16259,N_15393);
nand U16837 (N_16837,N_16224,N_16473);
and U16838 (N_16838,N_15210,N_15293);
xnor U16839 (N_16839,N_15150,N_15651);
nor U16840 (N_16840,N_15020,N_16339);
or U16841 (N_16841,N_15327,N_16038);
nand U16842 (N_16842,N_16493,N_15330);
and U16843 (N_16843,N_16436,N_15856);
xnor U16844 (N_16844,N_15635,N_15365);
and U16845 (N_16845,N_15994,N_15493);
and U16846 (N_16846,N_15236,N_16336);
nor U16847 (N_16847,N_15571,N_16034);
or U16848 (N_16848,N_15345,N_15793);
nand U16849 (N_16849,N_16019,N_16392);
xor U16850 (N_16850,N_15735,N_15754);
nor U16851 (N_16851,N_16310,N_15341);
nor U16852 (N_16852,N_16066,N_15008);
nand U16853 (N_16853,N_15617,N_15272);
nor U16854 (N_16854,N_15719,N_16282);
and U16855 (N_16855,N_15990,N_15764);
or U16856 (N_16856,N_15001,N_15009);
nor U16857 (N_16857,N_15061,N_15011);
xnor U16858 (N_16858,N_15089,N_16082);
nor U16859 (N_16859,N_16246,N_15196);
xnor U16860 (N_16860,N_15664,N_16355);
or U16861 (N_16861,N_15226,N_15962);
xor U16862 (N_16862,N_15075,N_16357);
or U16863 (N_16863,N_16407,N_16284);
nor U16864 (N_16864,N_15890,N_15926);
nor U16865 (N_16865,N_15261,N_15783);
nand U16866 (N_16866,N_16426,N_15044);
nand U16867 (N_16867,N_15514,N_15862);
nand U16868 (N_16868,N_15157,N_15711);
and U16869 (N_16869,N_15851,N_16316);
or U16870 (N_16870,N_15590,N_15024);
nor U16871 (N_16871,N_15883,N_15069);
and U16872 (N_16872,N_15291,N_15097);
or U16873 (N_16873,N_16420,N_15477);
nand U16874 (N_16874,N_16334,N_15155);
or U16875 (N_16875,N_16230,N_16254);
xor U16876 (N_16876,N_15791,N_15693);
or U16877 (N_16877,N_16294,N_15199);
or U16878 (N_16878,N_15073,N_15731);
and U16879 (N_16879,N_15301,N_16359);
and U16880 (N_16880,N_15316,N_15591);
or U16881 (N_16881,N_15273,N_15834);
nor U16882 (N_16882,N_15955,N_16105);
nor U16883 (N_16883,N_15753,N_16360);
nor U16884 (N_16884,N_15928,N_15995);
nand U16885 (N_16885,N_16204,N_16390);
and U16886 (N_16886,N_15919,N_16106);
nand U16887 (N_16887,N_15689,N_15563);
xor U16888 (N_16888,N_15736,N_15117);
nor U16889 (N_16889,N_15593,N_15946);
and U16890 (N_16890,N_15710,N_15867);
xnor U16891 (N_16891,N_16090,N_16474);
nand U16892 (N_16892,N_16394,N_15884);
xor U16893 (N_16893,N_15328,N_15036);
xor U16894 (N_16894,N_15740,N_15046);
nor U16895 (N_16895,N_15708,N_15127);
nor U16896 (N_16896,N_15808,N_15228);
and U16897 (N_16897,N_16366,N_16388);
xnor U16898 (N_16898,N_16053,N_16327);
and U16899 (N_16899,N_15786,N_15135);
xor U16900 (N_16900,N_15742,N_16446);
and U16901 (N_16901,N_15900,N_15683);
or U16902 (N_16902,N_15573,N_16194);
nor U16903 (N_16903,N_16329,N_15942);
nor U16904 (N_16904,N_15049,N_15806);
xnor U16905 (N_16905,N_15126,N_15496);
or U16906 (N_16906,N_15969,N_15847);
and U16907 (N_16907,N_16228,N_16171);
and U16908 (N_16908,N_16166,N_16486);
or U16909 (N_16909,N_15071,N_16160);
xor U16910 (N_16910,N_15827,N_16274);
or U16911 (N_16911,N_15971,N_15813);
and U16912 (N_16912,N_15007,N_15618);
nand U16913 (N_16913,N_15270,N_15234);
nand U16914 (N_16914,N_15530,N_15208);
nand U16915 (N_16915,N_15257,N_15985);
nor U16916 (N_16916,N_15275,N_16117);
nand U16917 (N_16917,N_15083,N_15388);
xor U16918 (N_16918,N_16350,N_16164);
xnor U16919 (N_16919,N_15777,N_16472);
and U16920 (N_16920,N_15243,N_15944);
or U16921 (N_16921,N_15286,N_15231);
or U16922 (N_16922,N_15351,N_15982);
nand U16923 (N_16923,N_15448,N_15216);
and U16924 (N_16924,N_16494,N_15871);
nand U16925 (N_16925,N_15146,N_15941);
and U16926 (N_16926,N_15715,N_15542);
nor U16927 (N_16927,N_16214,N_15787);
nand U16928 (N_16928,N_16447,N_16406);
xnor U16929 (N_16929,N_16223,N_15887);
or U16930 (N_16930,N_15503,N_16341);
xnor U16931 (N_16931,N_15209,N_15752);
or U16932 (N_16932,N_16454,N_15030);
and U16933 (N_16933,N_15667,N_16485);
nand U16934 (N_16934,N_15239,N_15158);
xor U16935 (N_16935,N_16092,N_15016);
xor U16936 (N_16936,N_15309,N_15180);
xor U16937 (N_16937,N_15848,N_15202);
nor U16938 (N_16938,N_15970,N_16257);
xnor U16939 (N_16939,N_16058,N_16431);
nand U16940 (N_16940,N_15106,N_16245);
nand U16941 (N_16941,N_15056,N_15535);
and U16942 (N_16942,N_15507,N_15757);
nor U16943 (N_16943,N_15170,N_15622);
or U16944 (N_16944,N_15665,N_15287);
or U16945 (N_16945,N_16212,N_15026);
xnor U16946 (N_16946,N_15892,N_16063);
and U16947 (N_16947,N_15454,N_15161);
xor U16948 (N_16948,N_15877,N_16187);
nor U16949 (N_16949,N_16227,N_15924);
or U16950 (N_16950,N_16471,N_16175);
or U16951 (N_16951,N_15189,N_15416);
or U16952 (N_16952,N_16476,N_15034);
nor U16953 (N_16953,N_15637,N_15893);
or U16954 (N_16954,N_16032,N_16384);
and U16955 (N_16955,N_16225,N_15596);
xnor U16956 (N_16956,N_16458,N_15842);
nand U16957 (N_16957,N_16113,N_16487);
nand U16958 (N_16958,N_16011,N_15304);
and U16959 (N_16959,N_15200,N_15331);
and U16960 (N_16960,N_15550,N_15803);
nor U16961 (N_16961,N_15889,N_15829);
nand U16962 (N_16962,N_15663,N_16455);
or U16963 (N_16963,N_16195,N_15785);
and U16964 (N_16964,N_15798,N_16026);
or U16965 (N_16965,N_15108,N_15644);
nor U16966 (N_16966,N_15169,N_15666);
xor U16967 (N_16967,N_16483,N_16124);
and U16968 (N_16968,N_15267,N_16272);
nand U16969 (N_16969,N_16182,N_16477);
xnor U16970 (N_16970,N_15882,N_15988);
nand U16971 (N_16971,N_15237,N_16115);
nand U16972 (N_16972,N_15361,N_15123);
nor U16973 (N_16973,N_15894,N_16100);
or U16974 (N_16974,N_15153,N_15249);
or U16975 (N_16975,N_16289,N_15383);
or U16976 (N_16976,N_15999,N_16112);
and U16977 (N_16977,N_15412,N_15370);
or U16978 (N_16978,N_15721,N_16333);
nor U16979 (N_16979,N_15182,N_15062);
and U16980 (N_16980,N_15154,N_15203);
nand U16981 (N_16981,N_15602,N_15680);
xor U16982 (N_16982,N_16490,N_16215);
xor U16983 (N_16983,N_15572,N_16304);
nand U16984 (N_16984,N_16157,N_15445);
xnor U16985 (N_16985,N_15143,N_15677);
xnor U16986 (N_16986,N_15434,N_15092);
nand U16987 (N_16987,N_16023,N_16030);
or U16988 (N_16988,N_15780,N_16158);
nand U16989 (N_16989,N_15886,N_15296);
and U16990 (N_16990,N_15455,N_16418);
nor U16991 (N_16991,N_15562,N_15932);
nand U16992 (N_16992,N_16382,N_16033);
and U16993 (N_16993,N_15379,N_15397);
xor U16994 (N_16994,N_16267,N_16285);
nand U16995 (N_16995,N_16084,N_16239);
nor U16996 (N_16996,N_16478,N_16137);
xnor U16997 (N_16997,N_16387,N_15395);
and U16998 (N_16998,N_15755,N_16280);
and U16999 (N_16999,N_16283,N_16345);
xnor U17000 (N_17000,N_16381,N_16300);
and U17001 (N_17001,N_16480,N_15349);
or U17002 (N_17002,N_15595,N_16126);
nand U17003 (N_17003,N_15163,N_15376);
xnor U17004 (N_17004,N_16221,N_15218);
xnor U17005 (N_17005,N_15966,N_15633);
and U17006 (N_17006,N_15909,N_15285);
or U17007 (N_17007,N_16429,N_16376);
nand U17008 (N_17008,N_15933,N_15874);
nand U17009 (N_17009,N_15624,N_15950);
nand U17010 (N_17010,N_15444,N_16496);
or U17011 (N_17011,N_15222,N_15147);
or U17012 (N_17012,N_15492,N_15329);
nor U17013 (N_17013,N_15037,N_15678);
and U17014 (N_17014,N_15700,N_15148);
or U17015 (N_17015,N_15289,N_15432);
nor U17016 (N_17016,N_16302,N_15640);
and U17017 (N_17017,N_16247,N_15645);
and U17018 (N_17018,N_16337,N_15022);
and U17019 (N_17019,N_15694,N_16401);
and U17020 (N_17020,N_15052,N_15066);
and U17021 (N_17021,N_15696,N_15173);
xnor U17022 (N_17022,N_15722,N_16275);
nor U17023 (N_17023,N_15364,N_16041);
nand U17024 (N_17024,N_15002,N_16442);
xor U17025 (N_17025,N_15181,N_15504);
xnor U17026 (N_17026,N_15307,N_16054);
and U17027 (N_17027,N_15265,N_15385);
xor U17028 (N_17028,N_16491,N_15881);
nand U17029 (N_17029,N_16343,N_15469);
or U17030 (N_17030,N_16083,N_15770);
xor U17031 (N_17031,N_15579,N_16266);
nor U17032 (N_17032,N_16253,N_16077);
or U17033 (N_17033,N_15745,N_16260);
nand U17034 (N_17034,N_16263,N_15549);
nand U17035 (N_17035,N_16064,N_15832);
xnor U17036 (N_17036,N_15099,N_15673);
and U17037 (N_17037,N_15490,N_15653);
nor U17038 (N_17038,N_16461,N_15247);
or U17039 (N_17039,N_15018,N_15576);
or U17040 (N_17040,N_15986,N_15144);
xnor U17041 (N_17041,N_15321,N_16441);
nand U17042 (N_17042,N_15610,N_15992);
nor U17043 (N_17043,N_15800,N_15906);
nor U17044 (N_17044,N_15197,N_15508);
nand U17045 (N_17045,N_16133,N_16467);
or U17046 (N_17046,N_15373,N_16180);
or U17047 (N_17047,N_16405,N_16149);
nor U17048 (N_17048,N_15427,N_15081);
nor U17049 (N_17049,N_15111,N_15248);
and U17050 (N_17050,N_16489,N_15281);
xnor U17051 (N_17051,N_15714,N_15927);
nand U17052 (N_17052,N_16378,N_16344);
or U17053 (N_17053,N_15600,N_15060);
nand U17054 (N_17054,N_15915,N_16220);
xor U17055 (N_17055,N_15171,N_16168);
xor U17056 (N_17056,N_15515,N_15820);
xor U17057 (N_17057,N_16475,N_16169);
and U17058 (N_17058,N_15428,N_15688);
xnor U17059 (N_17059,N_15648,N_15957);
and U17060 (N_17060,N_15489,N_15377);
nor U17061 (N_17061,N_16178,N_15391);
xor U17062 (N_17062,N_15059,N_15484);
nand U17063 (N_17063,N_16463,N_16086);
nand U17064 (N_17064,N_15415,N_16438);
xor U17065 (N_17065,N_15763,N_16161);
xor U17066 (N_17066,N_15121,N_15809);
xor U17067 (N_17067,N_15450,N_15292);
or U17068 (N_17068,N_16025,N_15453);
nand U17069 (N_17069,N_15055,N_16201);
xor U17070 (N_17070,N_15322,N_15979);
nor U17071 (N_17071,N_15805,N_15235);
xor U17072 (N_17072,N_15274,N_15625);
xor U17073 (N_17073,N_16002,N_15705);
nand U17074 (N_17074,N_16016,N_15138);
xor U17075 (N_17075,N_16156,N_16422);
and U17076 (N_17076,N_15480,N_15861);
or U17077 (N_17077,N_15639,N_15003);
or U17078 (N_17078,N_15027,N_16070);
nand U17079 (N_17079,N_16190,N_15305);
nand U17080 (N_17080,N_16005,N_15120);
nor U17081 (N_17081,N_16256,N_15461);
and U17082 (N_17082,N_16416,N_16152);
nand U17083 (N_17083,N_16217,N_15088);
nor U17084 (N_17084,N_15509,N_15464);
nor U17085 (N_17085,N_16445,N_15079);
or U17086 (N_17086,N_15276,N_16348);
or U17087 (N_17087,N_15401,N_15629);
nor U17088 (N_17088,N_15904,N_16128);
and U17089 (N_17089,N_15661,N_15822);
nand U17090 (N_17090,N_15468,N_15771);
or U17091 (N_17091,N_15703,N_15268);
or U17092 (N_17092,N_15098,N_15242);
and U17093 (N_17093,N_16258,N_15519);
and U17094 (N_17094,N_16167,N_16270);
nor U17095 (N_17095,N_15252,N_15830);
and U17096 (N_17096,N_15963,N_15565);
and U17097 (N_17097,N_16080,N_16427);
nand U17098 (N_17098,N_15255,N_15481);
xor U17099 (N_17099,N_16439,N_15058);
nand U17100 (N_17100,N_15937,N_15948);
or U17101 (N_17101,N_15394,N_16207);
nor U17102 (N_17102,N_16255,N_15400);
nand U17103 (N_17103,N_16462,N_15094);
or U17104 (N_17104,N_15524,N_15720);
xnor U17105 (N_17105,N_16031,N_15981);
nor U17106 (N_17106,N_15206,N_15086);
or U17107 (N_17107,N_15907,N_15959);
and U17108 (N_17108,N_15068,N_16236);
and U17109 (N_17109,N_15070,N_15038);
nand U17110 (N_17110,N_16383,N_15649);
nor U17111 (N_17111,N_15556,N_15205);
and U17112 (N_17112,N_15615,N_15768);
nor U17113 (N_17113,N_16052,N_15367);
xnor U17114 (N_17114,N_15669,N_15312);
nand U17115 (N_17115,N_15518,N_16037);
xnor U17116 (N_17116,N_15103,N_15939);
nor U17117 (N_17117,N_15019,N_16371);
xor U17118 (N_17118,N_15557,N_15095);
or U17119 (N_17119,N_15032,N_16059);
nor U17120 (N_17120,N_15474,N_15828);
nand U17121 (N_17121,N_15380,N_16153);
or U17122 (N_17122,N_15472,N_15998);
or U17123 (N_17123,N_15074,N_15360);
and U17124 (N_17124,N_16008,N_15278);
nor U17125 (N_17125,N_15898,N_16369);
and U17126 (N_17126,N_15744,N_15195);
nor U17127 (N_17127,N_15790,N_16413);
and U17128 (N_17128,N_15961,N_15613);
xnor U17129 (N_17129,N_15801,N_15294);
and U17130 (N_17130,N_15529,N_16138);
nor U17131 (N_17131,N_15488,N_16229);
or U17132 (N_17132,N_16120,N_15072);
nand U17133 (N_17133,N_16162,N_15921);
or U17134 (N_17134,N_16288,N_15681);
nand U17135 (N_17135,N_15028,N_16020);
nand U17136 (N_17136,N_15945,N_16411);
or U17137 (N_17137,N_15748,N_15826);
and U17138 (N_17138,N_15859,N_15051);
nor U17139 (N_17139,N_15517,N_15606);
nor U17140 (N_17140,N_16183,N_15043);
nor U17141 (N_17141,N_15471,N_15701);
nand U17142 (N_17142,N_16443,N_16241);
or U17143 (N_17143,N_15129,N_16428);
nand U17144 (N_17144,N_15864,N_15938);
nand U17145 (N_17145,N_16022,N_16370);
xnor U17146 (N_17146,N_15387,N_15818);
nor U17147 (N_17147,N_16320,N_15505);
nand U17148 (N_17148,N_15792,N_15430);
xnor U17149 (N_17149,N_16075,N_16061);
nor U17150 (N_17150,N_16303,N_15174);
xor U17151 (N_17151,N_16374,N_15258);
xnor U17152 (N_17152,N_15513,N_16393);
and U17153 (N_17153,N_16189,N_15298);
or U17154 (N_17154,N_16129,N_15246);
xor U17155 (N_17155,N_15417,N_15974);
nand U17156 (N_17156,N_15065,N_15130);
nor U17157 (N_17157,N_15873,N_15910);
or U17158 (N_17158,N_15047,N_16385);
and U17159 (N_17159,N_15728,N_15960);
nor U17160 (N_17160,N_16181,N_16367);
or U17161 (N_17161,N_15643,N_15035);
xnor U17162 (N_17162,N_15749,N_15336);
nor U17163 (N_17163,N_15987,N_16096);
xnor U17164 (N_17164,N_15642,N_15781);
nand U17165 (N_17165,N_15724,N_15078);
xnor U17166 (N_17166,N_16177,N_15358);
xor U17167 (N_17167,N_15778,N_15004);
or U17168 (N_17168,N_16354,N_15852);
nand U17169 (N_17169,N_15501,N_15414);
and U17170 (N_17170,N_15340,N_16010);
xor U17171 (N_17171,N_15659,N_15308);
nor U17172 (N_17172,N_16110,N_15396);
nand U17173 (N_17173,N_15219,N_16488);
nor U17174 (N_17174,N_15953,N_15656);
xor U17175 (N_17175,N_15005,N_16309);
xnor U17176 (N_17176,N_15612,N_16484);
nand U17177 (N_17177,N_15013,N_16028);
and U17178 (N_17178,N_15420,N_15936);
and U17179 (N_17179,N_15418,N_15041);
xor U17180 (N_17180,N_16440,N_15191);
or U17181 (N_17181,N_16127,N_16414);
or U17182 (N_17182,N_15465,N_16319);
nand U17183 (N_17183,N_16179,N_16163);
nand U17184 (N_17184,N_15675,N_15738);
xor U17185 (N_17185,N_16119,N_15583);
nand U17186 (N_17186,N_15836,N_15682);
or U17187 (N_17187,N_15063,N_15176);
nand U17188 (N_17188,N_15670,N_15930);
and U17189 (N_17189,N_15172,N_15362);
xor U17190 (N_17190,N_15303,N_16099);
nor U17191 (N_17191,N_15954,N_16352);
and U17192 (N_17192,N_16000,N_15463);
nor U17193 (N_17193,N_15502,N_15359);
nand U17194 (N_17194,N_15601,N_15599);
or U17195 (N_17195,N_15211,N_15227);
nand U17196 (N_17196,N_15136,N_15646);
and U17197 (N_17197,N_15372,N_15619);
nand U17198 (N_17198,N_15587,N_15597);
and U17199 (N_17199,N_15375,N_15885);
xor U17200 (N_17200,N_16081,N_15559);
or U17201 (N_17201,N_15371,N_15299);
nand U17202 (N_17202,N_16014,N_15398);
xnor U17203 (N_17203,N_16444,N_15628);
nor U17204 (N_17204,N_15374,N_15588);
xor U17205 (N_17205,N_16235,N_15156);
or U17206 (N_17206,N_15931,N_16237);
and U17207 (N_17207,N_15232,N_15935);
xnor U17208 (N_17208,N_15456,N_15855);
or U17209 (N_17209,N_15552,N_15223);
or U17210 (N_17210,N_15356,N_16358);
xor U17211 (N_17211,N_16372,N_15899);
nor U17212 (N_17212,N_16196,N_15922);
nand U17213 (N_17213,N_16338,N_16109);
and U17214 (N_17214,N_15626,N_15119);
and U17215 (N_17215,N_15085,N_15317);
or U17216 (N_17216,N_15408,N_15495);
nor U17217 (N_17217,N_15823,N_15605);
or U17218 (N_17218,N_15486,N_15627);
and U17219 (N_17219,N_15333,N_15440);
and U17220 (N_17220,N_15814,N_15707);
and U17221 (N_17221,N_16238,N_15451);
nand U17222 (N_17222,N_16377,N_16001);
nand U17223 (N_17223,N_16188,N_16210);
nor U17224 (N_17224,N_15064,N_15895);
and U17225 (N_17225,N_16430,N_15297);
or U17226 (N_17226,N_15435,N_15698);
and U17227 (N_17227,N_16142,N_15425);
or U17228 (N_17228,N_15527,N_15511);
nor U17229 (N_17229,N_15224,N_15225);
or U17230 (N_17230,N_15952,N_16365);
nand U17231 (N_17231,N_16067,N_15510);
and U17232 (N_17232,N_15691,N_15528);
or U17233 (N_17233,N_15841,N_15198);
nand U17234 (N_17234,N_15057,N_16202);
xnor U17235 (N_17235,N_16313,N_15817);
xor U17236 (N_17236,N_15984,N_15381);
and U17237 (N_17237,N_15537,N_15466);
xnor U17238 (N_17238,N_15151,N_16193);
and U17239 (N_17239,N_15459,N_15850);
or U17240 (N_17240,N_15494,N_15039);
and U17241 (N_17241,N_15429,N_16340);
xor U17242 (N_17242,N_15102,N_16170);
and U17243 (N_17243,N_15436,N_16123);
nand U17244 (N_17244,N_15577,N_15658);
nand U17245 (N_17245,N_16409,N_15240);
xnor U17246 (N_17246,N_16437,N_16286);
nor U17247 (N_17247,N_16492,N_16108);
nand U17248 (N_17248,N_15934,N_15114);
and U17249 (N_17249,N_16497,N_15860);
and U17250 (N_17250,N_15260,N_16293);
or U17251 (N_17251,N_15864,N_15743);
nor U17252 (N_17252,N_15307,N_15944);
xnor U17253 (N_17253,N_16036,N_15837);
xor U17254 (N_17254,N_15293,N_16170);
xor U17255 (N_17255,N_15278,N_15017);
or U17256 (N_17256,N_15047,N_15374);
nand U17257 (N_17257,N_15949,N_16076);
nand U17258 (N_17258,N_16274,N_15667);
xnor U17259 (N_17259,N_15753,N_16496);
xnor U17260 (N_17260,N_16160,N_15626);
xor U17261 (N_17261,N_16118,N_15988);
and U17262 (N_17262,N_15278,N_15584);
or U17263 (N_17263,N_15039,N_15993);
xor U17264 (N_17264,N_16166,N_15010);
and U17265 (N_17265,N_15423,N_16400);
nor U17266 (N_17266,N_15768,N_15955);
nor U17267 (N_17267,N_15642,N_15446);
or U17268 (N_17268,N_15652,N_15626);
nand U17269 (N_17269,N_15987,N_15267);
nor U17270 (N_17270,N_15134,N_16137);
xor U17271 (N_17271,N_15978,N_16348);
nor U17272 (N_17272,N_16469,N_15734);
nor U17273 (N_17273,N_16087,N_15027);
nand U17274 (N_17274,N_16197,N_15248);
nor U17275 (N_17275,N_15060,N_15849);
xnor U17276 (N_17276,N_16348,N_15380);
xnor U17277 (N_17277,N_16479,N_15546);
nand U17278 (N_17278,N_16082,N_16255);
nand U17279 (N_17279,N_16119,N_16191);
xnor U17280 (N_17280,N_15255,N_15821);
and U17281 (N_17281,N_16312,N_15867);
xnor U17282 (N_17282,N_15517,N_15699);
and U17283 (N_17283,N_15956,N_15536);
nand U17284 (N_17284,N_15700,N_16232);
xnor U17285 (N_17285,N_15758,N_15845);
and U17286 (N_17286,N_16218,N_15819);
nand U17287 (N_17287,N_15077,N_15297);
nand U17288 (N_17288,N_15578,N_16345);
or U17289 (N_17289,N_15512,N_16467);
xor U17290 (N_17290,N_15198,N_15210);
nor U17291 (N_17291,N_15063,N_15392);
nand U17292 (N_17292,N_16135,N_16448);
nand U17293 (N_17293,N_15628,N_16211);
nor U17294 (N_17294,N_15265,N_16267);
and U17295 (N_17295,N_16098,N_15229);
nand U17296 (N_17296,N_16094,N_15198);
or U17297 (N_17297,N_16460,N_16040);
nand U17298 (N_17298,N_15075,N_15568);
or U17299 (N_17299,N_15846,N_15148);
or U17300 (N_17300,N_15230,N_15060);
and U17301 (N_17301,N_15525,N_15762);
xnor U17302 (N_17302,N_15543,N_15570);
xnor U17303 (N_17303,N_15243,N_15539);
nor U17304 (N_17304,N_15969,N_16346);
nor U17305 (N_17305,N_15291,N_15939);
and U17306 (N_17306,N_15205,N_15938);
or U17307 (N_17307,N_16222,N_15397);
and U17308 (N_17308,N_15171,N_16096);
xnor U17309 (N_17309,N_15064,N_16179);
xor U17310 (N_17310,N_15200,N_16306);
or U17311 (N_17311,N_16363,N_16050);
and U17312 (N_17312,N_15597,N_15256);
or U17313 (N_17313,N_16261,N_15802);
and U17314 (N_17314,N_16345,N_15282);
nand U17315 (N_17315,N_16464,N_15763);
or U17316 (N_17316,N_15934,N_15481);
xor U17317 (N_17317,N_15071,N_15987);
and U17318 (N_17318,N_16458,N_15206);
or U17319 (N_17319,N_15523,N_15856);
and U17320 (N_17320,N_16012,N_15617);
nor U17321 (N_17321,N_15678,N_15714);
nand U17322 (N_17322,N_16190,N_16272);
xor U17323 (N_17323,N_15939,N_15402);
or U17324 (N_17324,N_15863,N_15185);
or U17325 (N_17325,N_15458,N_15244);
or U17326 (N_17326,N_15795,N_15809);
and U17327 (N_17327,N_15780,N_15675);
xnor U17328 (N_17328,N_15037,N_15828);
nor U17329 (N_17329,N_15110,N_15208);
nor U17330 (N_17330,N_16267,N_15931);
nor U17331 (N_17331,N_15663,N_16437);
or U17332 (N_17332,N_15833,N_16032);
nor U17333 (N_17333,N_15420,N_16066);
nor U17334 (N_17334,N_15314,N_16285);
and U17335 (N_17335,N_15837,N_16315);
nor U17336 (N_17336,N_15492,N_15065);
and U17337 (N_17337,N_16119,N_15497);
nor U17338 (N_17338,N_16116,N_16184);
nand U17339 (N_17339,N_15012,N_16207);
xor U17340 (N_17340,N_16346,N_15690);
or U17341 (N_17341,N_15058,N_15497);
and U17342 (N_17342,N_16159,N_15747);
xor U17343 (N_17343,N_15050,N_15391);
nand U17344 (N_17344,N_16088,N_15350);
or U17345 (N_17345,N_16455,N_15855);
nand U17346 (N_17346,N_15763,N_15543);
or U17347 (N_17347,N_16417,N_15202);
nor U17348 (N_17348,N_16352,N_15288);
nand U17349 (N_17349,N_15280,N_15705);
or U17350 (N_17350,N_15908,N_16336);
nand U17351 (N_17351,N_16156,N_15858);
or U17352 (N_17352,N_15844,N_15677);
nor U17353 (N_17353,N_15124,N_15807);
nand U17354 (N_17354,N_15286,N_16473);
nand U17355 (N_17355,N_15390,N_15253);
and U17356 (N_17356,N_15181,N_15035);
or U17357 (N_17357,N_16205,N_15274);
or U17358 (N_17358,N_15222,N_16086);
nand U17359 (N_17359,N_15866,N_16241);
xnor U17360 (N_17360,N_16443,N_15509);
or U17361 (N_17361,N_15141,N_15956);
nor U17362 (N_17362,N_15760,N_15046);
nand U17363 (N_17363,N_16020,N_15159);
nor U17364 (N_17364,N_16049,N_16267);
nor U17365 (N_17365,N_15507,N_15433);
and U17366 (N_17366,N_15879,N_15912);
xor U17367 (N_17367,N_16206,N_15757);
or U17368 (N_17368,N_15030,N_15486);
and U17369 (N_17369,N_15209,N_15845);
xor U17370 (N_17370,N_15278,N_16077);
xor U17371 (N_17371,N_16407,N_16415);
or U17372 (N_17372,N_15102,N_16352);
nor U17373 (N_17373,N_16442,N_15006);
xor U17374 (N_17374,N_15498,N_15899);
or U17375 (N_17375,N_16037,N_15804);
and U17376 (N_17376,N_15553,N_15274);
xor U17377 (N_17377,N_15661,N_15858);
nand U17378 (N_17378,N_16113,N_16280);
or U17379 (N_17379,N_16302,N_15081);
nand U17380 (N_17380,N_16362,N_15646);
and U17381 (N_17381,N_15392,N_15417);
xnor U17382 (N_17382,N_15191,N_15185);
nand U17383 (N_17383,N_15177,N_15138);
and U17384 (N_17384,N_15491,N_16191);
xnor U17385 (N_17385,N_15077,N_16144);
and U17386 (N_17386,N_15342,N_15439);
and U17387 (N_17387,N_16194,N_16237);
nor U17388 (N_17388,N_16346,N_15874);
nor U17389 (N_17389,N_15679,N_16238);
xor U17390 (N_17390,N_15961,N_16120);
nor U17391 (N_17391,N_15461,N_16474);
xor U17392 (N_17392,N_16033,N_15096);
and U17393 (N_17393,N_16310,N_15343);
and U17394 (N_17394,N_16150,N_16194);
nor U17395 (N_17395,N_15507,N_16176);
nor U17396 (N_17396,N_15682,N_15548);
and U17397 (N_17397,N_15721,N_16088);
or U17398 (N_17398,N_15251,N_15159);
nor U17399 (N_17399,N_15722,N_15374);
xor U17400 (N_17400,N_15210,N_15318);
nor U17401 (N_17401,N_16107,N_15672);
and U17402 (N_17402,N_15569,N_15242);
or U17403 (N_17403,N_15609,N_15966);
nor U17404 (N_17404,N_16017,N_15661);
nor U17405 (N_17405,N_15365,N_15663);
and U17406 (N_17406,N_16398,N_15085);
or U17407 (N_17407,N_15611,N_16067);
and U17408 (N_17408,N_15664,N_15284);
xnor U17409 (N_17409,N_15635,N_15938);
nor U17410 (N_17410,N_15165,N_15375);
and U17411 (N_17411,N_15724,N_15002);
nor U17412 (N_17412,N_15087,N_16354);
xnor U17413 (N_17413,N_16029,N_15265);
xor U17414 (N_17414,N_15849,N_15585);
and U17415 (N_17415,N_16250,N_16165);
nand U17416 (N_17416,N_16161,N_15836);
nand U17417 (N_17417,N_15409,N_15628);
and U17418 (N_17418,N_16054,N_16447);
xnor U17419 (N_17419,N_16201,N_16040);
nor U17420 (N_17420,N_15115,N_15266);
nor U17421 (N_17421,N_16297,N_16193);
xor U17422 (N_17422,N_15619,N_16017);
nor U17423 (N_17423,N_16377,N_15015);
xnor U17424 (N_17424,N_16259,N_15376);
nand U17425 (N_17425,N_16139,N_15486);
nor U17426 (N_17426,N_15855,N_16309);
and U17427 (N_17427,N_15361,N_16133);
and U17428 (N_17428,N_16197,N_16267);
or U17429 (N_17429,N_16272,N_16321);
xnor U17430 (N_17430,N_16148,N_15542);
xor U17431 (N_17431,N_16114,N_15372);
nor U17432 (N_17432,N_16196,N_15933);
xor U17433 (N_17433,N_15601,N_15147);
or U17434 (N_17434,N_16363,N_15853);
and U17435 (N_17435,N_15993,N_16419);
nand U17436 (N_17436,N_15518,N_16163);
and U17437 (N_17437,N_16250,N_15592);
and U17438 (N_17438,N_16225,N_15148);
and U17439 (N_17439,N_15645,N_15845);
or U17440 (N_17440,N_15402,N_15424);
and U17441 (N_17441,N_16375,N_15811);
nand U17442 (N_17442,N_15180,N_15284);
nor U17443 (N_17443,N_15370,N_16145);
or U17444 (N_17444,N_15682,N_15123);
xnor U17445 (N_17445,N_15204,N_16057);
xnor U17446 (N_17446,N_16072,N_15735);
or U17447 (N_17447,N_16177,N_15672);
or U17448 (N_17448,N_16347,N_16175);
and U17449 (N_17449,N_15289,N_15578);
or U17450 (N_17450,N_16166,N_15243);
xnor U17451 (N_17451,N_15006,N_15821);
and U17452 (N_17452,N_15281,N_15049);
nor U17453 (N_17453,N_16377,N_15800);
nor U17454 (N_17454,N_16141,N_16120);
or U17455 (N_17455,N_15367,N_16114);
and U17456 (N_17456,N_15179,N_15284);
xnor U17457 (N_17457,N_16111,N_15186);
or U17458 (N_17458,N_16462,N_16180);
nor U17459 (N_17459,N_15150,N_16342);
xnor U17460 (N_17460,N_16497,N_15671);
nand U17461 (N_17461,N_15874,N_15141);
nor U17462 (N_17462,N_15231,N_15558);
or U17463 (N_17463,N_15602,N_15473);
or U17464 (N_17464,N_15918,N_16040);
and U17465 (N_17465,N_15081,N_15220);
or U17466 (N_17466,N_15195,N_15812);
xor U17467 (N_17467,N_16184,N_16084);
nand U17468 (N_17468,N_15366,N_15802);
or U17469 (N_17469,N_16385,N_15094);
nor U17470 (N_17470,N_15588,N_16448);
nor U17471 (N_17471,N_16244,N_15346);
xnor U17472 (N_17472,N_16078,N_16319);
and U17473 (N_17473,N_15755,N_15441);
xor U17474 (N_17474,N_15793,N_16483);
nand U17475 (N_17475,N_15708,N_15674);
xor U17476 (N_17476,N_15493,N_16429);
or U17477 (N_17477,N_16086,N_15563);
or U17478 (N_17478,N_16057,N_16376);
nand U17479 (N_17479,N_15560,N_15299);
nand U17480 (N_17480,N_15399,N_15648);
nor U17481 (N_17481,N_15142,N_16215);
nand U17482 (N_17482,N_15628,N_16145);
nand U17483 (N_17483,N_15901,N_15694);
nor U17484 (N_17484,N_16040,N_16402);
nor U17485 (N_17485,N_16137,N_15263);
nand U17486 (N_17486,N_15896,N_15759);
nand U17487 (N_17487,N_15057,N_16439);
or U17488 (N_17488,N_15835,N_15104);
nor U17489 (N_17489,N_16279,N_15075);
nor U17490 (N_17490,N_15502,N_15384);
nand U17491 (N_17491,N_16235,N_15509);
and U17492 (N_17492,N_15560,N_15984);
and U17493 (N_17493,N_16370,N_15182);
or U17494 (N_17494,N_15234,N_15592);
nor U17495 (N_17495,N_16171,N_16369);
and U17496 (N_17496,N_15063,N_15342);
nand U17497 (N_17497,N_16345,N_15556);
or U17498 (N_17498,N_16352,N_16319);
xor U17499 (N_17499,N_15508,N_16410);
xor U17500 (N_17500,N_16365,N_15235);
xnor U17501 (N_17501,N_16277,N_15379);
nor U17502 (N_17502,N_15433,N_15995);
and U17503 (N_17503,N_16206,N_16498);
xnor U17504 (N_17504,N_15879,N_15645);
nor U17505 (N_17505,N_15851,N_16394);
xor U17506 (N_17506,N_15452,N_15600);
nand U17507 (N_17507,N_15531,N_16494);
and U17508 (N_17508,N_15145,N_15554);
nand U17509 (N_17509,N_16081,N_15785);
nand U17510 (N_17510,N_15344,N_16263);
nand U17511 (N_17511,N_15489,N_16369);
nand U17512 (N_17512,N_16219,N_15880);
or U17513 (N_17513,N_15644,N_15225);
nor U17514 (N_17514,N_15703,N_15479);
or U17515 (N_17515,N_15084,N_15670);
and U17516 (N_17516,N_16084,N_16319);
and U17517 (N_17517,N_16463,N_15424);
nand U17518 (N_17518,N_15273,N_15904);
nand U17519 (N_17519,N_15540,N_15154);
xor U17520 (N_17520,N_15116,N_16359);
xor U17521 (N_17521,N_15323,N_15900);
and U17522 (N_17522,N_15149,N_15605);
and U17523 (N_17523,N_16103,N_15645);
nand U17524 (N_17524,N_15428,N_16069);
or U17525 (N_17525,N_15317,N_16277);
or U17526 (N_17526,N_15112,N_15338);
nor U17527 (N_17527,N_16378,N_16078);
xor U17528 (N_17528,N_16375,N_15624);
and U17529 (N_17529,N_15649,N_15699);
nor U17530 (N_17530,N_15711,N_15767);
or U17531 (N_17531,N_15630,N_15397);
nor U17532 (N_17532,N_16492,N_15861);
or U17533 (N_17533,N_15841,N_16130);
nor U17534 (N_17534,N_16346,N_16379);
xnor U17535 (N_17535,N_16154,N_15569);
nand U17536 (N_17536,N_15903,N_16296);
nor U17537 (N_17537,N_15261,N_16408);
xnor U17538 (N_17538,N_16180,N_15558);
and U17539 (N_17539,N_15801,N_15127);
or U17540 (N_17540,N_15707,N_15909);
nand U17541 (N_17541,N_16303,N_15696);
nor U17542 (N_17542,N_16293,N_15201);
nor U17543 (N_17543,N_15446,N_16329);
or U17544 (N_17544,N_15837,N_16482);
xnor U17545 (N_17545,N_15532,N_16383);
xor U17546 (N_17546,N_15604,N_15202);
and U17547 (N_17547,N_15948,N_16185);
nor U17548 (N_17548,N_15291,N_15802);
nand U17549 (N_17549,N_15433,N_15552);
or U17550 (N_17550,N_16358,N_15817);
or U17551 (N_17551,N_15640,N_15010);
or U17552 (N_17552,N_16056,N_16153);
nand U17553 (N_17553,N_16208,N_15118);
nor U17554 (N_17554,N_16246,N_15328);
and U17555 (N_17555,N_15217,N_15186);
or U17556 (N_17556,N_16459,N_15164);
and U17557 (N_17557,N_15928,N_16098);
and U17558 (N_17558,N_15530,N_16355);
nand U17559 (N_17559,N_15520,N_15521);
xor U17560 (N_17560,N_15395,N_15269);
nor U17561 (N_17561,N_15145,N_15742);
nand U17562 (N_17562,N_15359,N_16487);
nand U17563 (N_17563,N_15116,N_15345);
nand U17564 (N_17564,N_15947,N_16113);
nand U17565 (N_17565,N_15453,N_15219);
and U17566 (N_17566,N_15362,N_15991);
nand U17567 (N_17567,N_15139,N_15476);
nand U17568 (N_17568,N_15146,N_16008);
and U17569 (N_17569,N_15435,N_15594);
nor U17570 (N_17570,N_15616,N_16244);
xor U17571 (N_17571,N_15444,N_16328);
or U17572 (N_17572,N_15259,N_16168);
nor U17573 (N_17573,N_15337,N_16272);
xor U17574 (N_17574,N_15246,N_15677);
nand U17575 (N_17575,N_15264,N_15684);
nand U17576 (N_17576,N_15404,N_15148);
or U17577 (N_17577,N_15717,N_16224);
or U17578 (N_17578,N_15369,N_15946);
nor U17579 (N_17579,N_16361,N_15933);
or U17580 (N_17580,N_15395,N_16277);
or U17581 (N_17581,N_16242,N_15123);
xnor U17582 (N_17582,N_16432,N_15840);
and U17583 (N_17583,N_15436,N_15109);
xnor U17584 (N_17584,N_15045,N_15726);
nand U17585 (N_17585,N_16300,N_15826);
nor U17586 (N_17586,N_15796,N_16484);
nand U17587 (N_17587,N_16380,N_15857);
and U17588 (N_17588,N_16322,N_16281);
and U17589 (N_17589,N_15971,N_15576);
xnor U17590 (N_17590,N_15492,N_15071);
xor U17591 (N_17591,N_16127,N_15864);
and U17592 (N_17592,N_15940,N_15731);
and U17593 (N_17593,N_15423,N_16095);
nor U17594 (N_17594,N_16380,N_15110);
xnor U17595 (N_17595,N_15192,N_15101);
nand U17596 (N_17596,N_16058,N_16289);
nor U17597 (N_17597,N_16280,N_15340);
nand U17598 (N_17598,N_15729,N_15199);
and U17599 (N_17599,N_15671,N_16131);
nor U17600 (N_17600,N_15582,N_15036);
nor U17601 (N_17601,N_15304,N_16465);
nand U17602 (N_17602,N_16084,N_15751);
xnor U17603 (N_17603,N_15086,N_15358);
nor U17604 (N_17604,N_15200,N_15922);
nor U17605 (N_17605,N_16405,N_15897);
nor U17606 (N_17606,N_15288,N_16032);
nor U17607 (N_17607,N_15500,N_16091);
xnor U17608 (N_17608,N_15448,N_16178);
xnor U17609 (N_17609,N_15668,N_15086);
and U17610 (N_17610,N_15395,N_16419);
nor U17611 (N_17611,N_16171,N_16367);
or U17612 (N_17612,N_16353,N_16458);
nor U17613 (N_17613,N_16233,N_16100);
and U17614 (N_17614,N_15237,N_15784);
nand U17615 (N_17615,N_15341,N_16199);
nand U17616 (N_17616,N_16361,N_15857);
nor U17617 (N_17617,N_15724,N_15725);
or U17618 (N_17618,N_15911,N_15695);
xor U17619 (N_17619,N_15733,N_15200);
nand U17620 (N_17620,N_15636,N_15620);
xor U17621 (N_17621,N_16366,N_15933);
nand U17622 (N_17622,N_15105,N_16351);
or U17623 (N_17623,N_16357,N_15334);
nor U17624 (N_17624,N_15664,N_15107);
nor U17625 (N_17625,N_16324,N_16072);
nor U17626 (N_17626,N_15241,N_15771);
xnor U17627 (N_17627,N_16330,N_15177);
xor U17628 (N_17628,N_15296,N_15257);
nor U17629 (N_17629,N_15479,N_15297);
nand U17630 (N_17630,N_16066,N_15641);
or U17631 (N_17631,N_16189,N_15043);
nor U17632 (N_17632,N_15436,N_15956);
xnor U17633 (N_17633,N_16489,N_15064);
xor U17634 (N_17634,N_15368,N_15343);
or U17635 (N_17635,N_15806,N_15552);
and U17636 (N_17636,N_15505,N_15935);
or U17637 (N_17637,N_15580,N_15719);
or U17638 (N_17638,N_15997,N_15627);
nand U17639 (N_17639,N_16369,N_15227);
nand U17640 (N_17640,N_15539,N_15961);
or U17641 (N_17641,N_15868,N_15278);
nand U17642 (N_17642,N_15474,N_16008);
or U17643 (N_17643,N_15187,N_15449);
xnor U17644 (N_17644,N_16472,N_16085);
and U17645 (N_17645,N_16327,N_16281);
or U17646 (N_17646,N_15064,N_16138);
or U17647 (N_17647,N_16175,N_15715);
and U17648 (N_17648,N_15797,N_15921);
or U17649 (N_17649,N_15746,N_15851);
xor U17650 (N_17650,N_16359,N_16114);
nor U17651 (N_17651,N_16383,N_15002);
nand U17652 (N_17652,N_15264,N_15617);
xnor U17653 (N_17653,N_16372,N_15798);
and U17654 (N_17654,N_15653,N_15353);
nor U17655 (N_17655,N_15029,N_15937);
nand U17656 (N_17656,N_15665,N_16047);
nor U17657 (N_17657,N_16482,N_15839);
xor U17658 (N_17658,N_16138,N_15801);
nand U17659 (N_17659,N_15388,N_15557);
nor U17660 (N_17660,N_15340,N_15872);
xnor U17661 (N_17661,N_15630,N_16133);
or U17662 (N_17662,N_15379,N_16052);
xnor U17663 (N_17663,N_15876,N_16015);
nor U17664 (N_17664,N_15522,N_15115);
nor U17665 (N_17665,N_15613,N_15209);
xnor U17666 (N_17666,N_16354,N_15552);
nor U17667 (N_17667,N_15373,N_15686);
nor U17668 (N_17668,N_15775,N_16129);
nor U17669 (N_17669,N_15518,N_16242);
and U17670 (N_17670,N_15352,N_15412);
or U17671 (N_17671,N_15644,N_15149);
nand U17672 (N_17672,N_16254,N_15737);
nor U17673 (N_17673,N_15618,N_15692);
and U17674 (N_17674,N_15478,N_16163);
xnor U17675 (N_17675,N_15736,N_15462);
nor U17676 (N_17676,N_16191,N_15546);
and U17677 (N_17677,N_15974,N_15539);
xor U17678 (N_17678,N_15627,N_15681);
or U17679 (N_17679,N_15646,N_16427);
and U17680 (N_17680,N_15161,N_16213);
nand U17681 (N_17681,N_16444,N_16403);
or U17682 (N_17682,N_15730,N_15960);
nor U17683 (N_17683,N_15249,N_15564);
and U17684 (N_17684,N_16171,N_15167);
xor U17685 (N_17685,N_15471,N_15513);
nor U17686 (N_17686,N_15948,N_16198);
nor U17687 (N_17687,N_15787,N_15109);
or U17688 (N_17688,N_15287,N_15995);
and U17689 (N_17689,N_16221,N_15746);
or U17690 (N_17690,N_15634,N_15513);
nor U17691 (N_17691,N_16218,N_16046);
or U17692 (N_17692,N_15089,N_15432);
nor U17693 (N_17693,N_16047,N_15992);
nand U17694 (N_17694,N_16443,N_15990);
nor U17695 (N_17695,N_16242,N_15503);
or U17696 (N_17696,N_15085,N_15849);
nor U17697 (N_17697,N_16018,N_15579);
xnor U17698 (N_17698,N_16091,N_15786);
nor U17699 (N_17699,N_16499,N_16081);
and U17700 (N_17700,N_16088,N_15679);
and U17701 (N_17701,N_16266,N_16419);
and U17702 (N_17702,N_16033,N_15868);
nor U17703 (N_17703,N_15472,N_15340);
nor U17704 (N_17704,N_15641,N_16499);
or U17705 (N_17705,N_16312,N_16423);
nand U17706 (N_17706,N_15567,N_16022);
nand U17707 (N_17707,N_15655,N_15871);
nand U17708 (N_17708,N_15861,N_15746);
or U17709 (N_17709,N_15984,N_15458);
xor U17710 (N_17710,N_16031,N_15079);
and U17711 (N_17711,N_15793,N_15776);
and U17712 (N_17712,N_15136,N_16256);
nand U17713 (N_17713,N_15051,N_15164);
and U17714 (N_17714,N_16272,N_15796);
xnor U17715 (N_17715,N_16095,N_16116);
or U17716 (N_17716,N_15163,N_15382);
nand U17717 (N_17717,N_15199,N_16028);
nand U17718 (N_17718,N_16377,N_15667);
nand U17719 (N_17719,N_16301,N_15592);
or U17720 (N_17720,N_15720,N_16470);
xor U17721 (N_17721,N_15159,N_15989);
nand U17722 (N_17722,N_16451,N_15679);
or U17723 (N_17723,N_15683,N_15681);
and U17724 (N_17724,N_16301,N_16090);
xor U17725 (N_17725,N_15427,N_15234);
and U17726 (N_17726,N_16033,N_15657);
or U17727 (N_17727,N_16021,N_16218);
nand U17728 (N_17728,N_16139,N_16189);
nand U17729 (N_17729,N_15110,N_16148);
xor U17730 (N_17730,N_16495,N_15741);
nor U17731 (N_17731,N_15484,N_15990);
nand U17732 (N_17732,N_15839,N_15020);
and U17733 (N_17733,N_15655,N_16307);
nor U17734 (N_17734,N_15569,N_15352);
or U17735 (N_17735,N_16322,N_15688);
nand U17736 (N_17736,N_16075,N_15071);
or U17737 (N_17737,N_16052,N_16383);
nand U17738 (N_17738,N_16096,N_15784);
nor U17739 (N_17739,N_15329,N_16143);
xnor U17740 (N_17740,N_16381,N_15359);
nand U17741 (N_17741,N_15101,N_15079);
nor U17742 (N_17742,N_15256,N_15998);
and U17743 (N_17743,N_15011,N_16313);
or U17744 (N_17744,N_16019,N_16177);
and U17745 (N_17745,N_15826,N_15713);
nor U17746 (N_17746,N_15573,N_16265);
nor U17747 (N_17747,N_15221,N_15986);
xor U17748 (N_17748,N_15200,N_16257);
or U17749 (N_17749,N_16212,N_16268);
nor U17750 (N_17750,N_16053,N_16146);
or U17751 (N_17751,N_15171,N_15505);
xor U17752 (N_17752,N_16285,N_15475);
xor U17753 (N_17753,N_16130,N_15535);
nor U17754 (N_17754,N_16453,N_16340);
and U17755 (N_17755,N_15876,N_15918);
and U17756 (N_17756,N_15143,N_16484);
nand U17757 (N_17757,N_16009,N_15135);
nor U17758 (N_17758,N_15947,N_16129);
nor U17759 (N_17759,N_15154,N_15547);
and U17760 (N_17760,N_15728,N_15597);
nor U17761 (N_17761,N_15008,N_15083);
and U17762 (N_17762,N_15305,N_15903);
and U17763 (N_17763,N_15436,N_16371);
nor U17764 (N_17764,N_15887,N_15654);
and U17765 (N_17765,N_15341,N_15813);
nand U17766 (N_17766,N_16203,N_15219);
nand U17767 (N_17767,N_16314,N_15601);
xnor U17768 (N_17768,N_15333,N_15664);
or U17769 (N_17769,N_15035,N_16238);
and U17770 (N_17770,N_15735,N_16021);
nand U17771 (N_17771,N_15607,N_15663);
nor U17772 (N_17772,N_15555,N_16249);
or U17773 (N_17773,N_15374,N_15367);
nand U17774 (N_17774,N_15010,N_15195);
and U17775 (N_17775,N_15581,N_15239);
xor U17776 (N_17776,N_16476,N_16477);
xnor U17777 (N_17777,N_16321,N_16226);
or U17778 (N_17778,N_15442,N_16430);
xor U17779 (N_17779,N_16009,N_15956);
or U17780 (N_17780,N_15658,N_15744);
xor U17781 (N_17781,N_16307,N_15306);
and U17782 (N_17782,N_15672,N_15683);
nor U17783 (N_17783,N_15049,N_16302);
nor U17784 (N_17784,N_15480,N_15388);
nand U17785 (N_17785,N_15112,N_16427);
or U17786 (N_17786,N_15611,N_16162);
nand U17787 (N_17787,N_16397,N_16481);
and U17788 (N_17788,N_16124,N_15654);
xnor U17789 (N_17789,N_15417,N_16068);
and U17790 (N_17790,N_15635,N_15123);
nand U17791 (N_17791,N_15160,N_16310);
xor U17792 (N_17792,N_15566,N_15523);
or U17793 (N_17793,N_16481,N_15006);
or U17794 (N_17794,N_15191,N_15068);
nand U17795 (N_17795,N_16132,N_16104);
xnor U17796 (N_17796,N_15570,N_15330);
xor U17797 (N_17797,N_16340,N_16216);
nand U17798 (N_17798,N_16213,N_15519);
xnor U17799 (N_17799,N_16126,N_16132);
xor U17800 (N_17800,N_15156,N_15940);
and U17801 (N_17801,N_15381,N_15063);
and U17802 (N_17802,N_15771,N_16141);
and U17803 (N_17803,N_16479,N_16487);
nand U17804 (N_17804,N_15880,N_15584);
or U17805 (N_17805,N_15216,N_15921);
and U17806 (N_17806,N_15250,N_15880);
xnor U17807 (N_17807,N_15133,N_15890);
or U17808 (N_17808,N_15070,N_15253);
xnor U17809 (N_17809,N_15625,N_15519);
nand U17810 (N_17810,N_16158,N_16085);
and U17811 (N_17811,N_16382,N_16388);
or U17812 (N_17812,N_16154,N_16068);
nand U17813 (N_17813,N_15674,N_15062);
xnor U17814 (N_17814,N_16195,N_16217);
nand U17815 (N_17815,N_16156,N_15272);
or U17816 (N_17816,N_15231,N_16091);
or U17817 (N_17817,N_15404,N_16473);
nand U17818 (N_17818,N_15825,N_16145);
nor U17819 (N_17819,N_16337,N_15404);
xor U17820 (N_17820,N_15700,N_16371);
or U17821 (N_17821,N_16373,N_15855);
xnor U17822 (N_17822,N_15543,N_16125);
or U17823 (N_17823,N_16315,N_16455);
and U17824 (N_17824,N_15342,N_15214);
nor U17825 (N_17825,N_15951,N_15683);
and U17826 (N_17826,N_15157,N_15447);
or U17827 (N_17827,N_15343,N_15775);
nor U17828 (N_17828,N_15748,N_16232);
nor U17829 (N_17829,N_15545,N_15325);
nand U17830 (N_17830,N_15964,N_15054);
or U17831 (N_17831,N_16233,N_16449);
nor U17832 (N_17832,N_16261,N_16309);
or U17833 (N_17833,N_15959,N_15166);
nand U17834 (N_17834,N_15546,N_16297);
nor U17835 (N_17835,N_15955,N_15031);
nor U17836 (N_17836,N_15746,N_16282);
or U17837 (N_17837,N_15229,N_15029);
nor U17838 (N_17838,N_16019,N_15761);
and U17839 (N_17839,N_15676,N_15379);
nand U17840 (N_17840,N_16207,N_16357);
and U17841 (N_17841,N_16165,N_16483);
or U17842 (N_17842,N_16385,N_15457);
nand U17843 (N_17843,N_16058,N_15225);
and U17844 (N_17844,N_16034,N_16431);
nand U17845 (N_17845,N_16021,N_16460);
and U17846 (N_17846,N_15841,N_15470);
and U17847 (N_17847,N_16138,N_15284);
nor U17848 (N_17848,N_15860,N_15577);
or U17849 (N_17849,N_16318,N_15886);
or U17850 (N_17850,N_15383,N_15573);
xnor U17851 (N_17851,N_15769,N_15231);
nor U17852 (N_17852,N_16195,N_15140);
nand U17853 (N_17853,N_16368,N_15947);
and U17854 (N_17854,N_16191,N_15077);
nor U17855 (N_17855,N_15577,N_15372);
nor U17856 (N_17856,N_16057,N_15390);
nand U17857 (N_17857,N_15968,N_15405);
xnor U17858 (N_17858,N_15357,N_16181);
xnor U17859 (N_17859,N_15261,N_15317);
nor U17860 (N_17860,N_15723,N_15390);
xor U17861 (N_17861,N_16215,N_15210);
nor U17862 (N_17862,N_16390,N_16202);
or U17863 (N_17863,N_16129,N_15730);
nor U17864 (N_17864,N_15770,N_16225);
xor U17865 (N_17865,N_15382,N_16021);
nand U17866 (N_17866,N_15815,N_15217);
or U17867 (N_17867,N_15346,N_15241);
and U17868 (N_17868,N_15604,N_16497);
nand U17869 (N_17869,N_16019,N_16199);
xor U17870 (N_17870,N_16240,N_16246);
or U17871 (N_17871,N_15347,N_15458);
and U17872 (N_17872,N_15710,N_15654);
nand U17873 (N_17873,N_16288,N_16101);
or U17874 (N_17874,N_15009,N_15379);
nor U17875 (N_17875,N_15196,N_16267);
nor U17876 (N_17876,N_15172,N_15001);
nor U17877 (N_17877,N_15371,N_15379);
or U17878 (N_17878,N_15237,N_15592);
nor U17879 (N_17879,N_15889,N_15517);
or U17880 (N_17880,N_16032,N_15098);
nor U17881 (N_17881,N_15366,N_15359);
nor U17882 (N_17882,N_15750,N_15071);
and U17883 (N_17883,N_16002,N_15678);
nor U17884 (N_17884,N_15734,N_15307);
nor U17885 (N_17885,N_15357,N_15450);
or U17886 (N_17886,N_15309,N_15239);
nor U17887 (N_17887,N_16098,N_15517);
or U17888 (N_17888,N_15443,N_16386);
xnor U17889 (N_17889,N_16212,N_15909);
xnor U17890 (N_17890,N_16392,N_15912);
nor U17891 (N_17891,N_15951,N_15479);
and U17892 (N_17892,N_16302,N_16303);
and U17893 (N_17893,N_15172,N_16225);
nor U17894 (N_17894,N_15582,N_15687);
nor U17895 (N_17895,N_15895,N_16315);
nor U17896 (N_17896,N_15904,N_15811);
nand U17897 (N_17897,N_16012,N_16214);
and U17898 (N_17898,N_16262,N_15252);
or U17899 (N_17899,N_16301,N_15373);
or U17900 (N_17900,N_15833,N_16066);
nand U17901 (N_17901,N_16476,N_16311);
nor U17902 (N_17902,N_15894,N_15977);
and U17903 (N_17903,N_15689,N_15834);
nor U17904 (N_17904,N_16314,N_15158);
or U17905 (N_17905,N_15471,N_15015);
nand U17906 (N_17906,N_15369,N_15452);
nand U17907 (N_17907,N_15639,N_15179);
nand U17908 (N_17908,N_15601,N_15900);
nor U17909 (N_17909,N_16433,N_16165);
and U17910 (N_17910,N_15477,N_16275);
xor U17911 (N_17911,N_16206,N_16181);
xor U17912 (N_17912,N_16260,N_15692);
nand U17913 (N_17913,N_15041,N_15810);
and U17914 (N_17914,N_15217,N_15535);
or U17915 (N_17915,N_15117,N_15938);
nand U17916 (N_17916,N_15768,N_15155);
and U17917 (N_17917,N_15394,N_16198);
or U17918 (N_17918,N_16038,N_15552);
xnor U17919 (N_17919,N_15738,N_15701);
nor U17920 (N_17920,N_16197,N_16294);
xor U17921 (N_17921,N_16268,N_16276);
nand U17922 (N_17922,N_16154,N_16410);
nand U17923 (N_17923,N_15574,N_16108);
xnor U17924 (N_17924,N_16183,N_15703);
or U17925 (N_17925,N_15694,N_16357);
xor U17926 (N_17926,N_15426,N_15969);
or U17927 (N_17927,N_15648,N_15144);
nor U17928 (N_17928,N_15148,N_15530);
nand U17929 (N_17929,N_15551,N_15739);
and U17930 (N_17930,N_16199,N_15865);
nor U17931 (N_17931,N_16088,N_15554);
and U17932 (N_17932,N_15594,N_16156);
and U17933 (N_17933,N_15551,N_15576);
nand U17934 (N_17934,N_16264,N_15890);
or U17935 (N_17935,N_15165,N_15449);
xnor U17936 (N_17936,N_16496,N_15385);
and U17937 (N_17937,N_15295,N_15576);
nor U17938 (N_17938,N_16049,N_16195);
nand U17939 (N_17939,N_15622,N_15470);
nor U17940 (N_17940,N_16057,N_16414);
xnor U17941 (N_17941,N_15912,N_16338);
and U17942 (N_17942,N_15884,N_15155);
or U17943 (N_17943,N_16075,N_16169);
xor U17944 (N_17944,N_15002,N_15723);
nand U17945 (N_17945,N_15689,N_16363);
and U17946 (N_17946,N_15321,N_16210);
and U17947 (N_17947,N_16456,N_16181);
xnor U17948 (N_17948,N_15157,N_15500);
or U17949 (N_17949,N_15830,N_15750);
or U17950 (N_17950,N_15146,N_16000);
xor U17951 (N_17951,N_16324,N_16196);
and U17952 (N_17952,N_15379,N_15288);
xnor U17953 (N_17953,N_16403,N_16263);
xnor U17954 (N_17954,N_15906,N_16129);
and U17955 (N_17955,N_15342,N_15637);
xnor U17956 (N_17956,N_16353,N_15141);
or U17957 (N_17957,N_15611,N_16387);
or U17958 (N_17958,N_15427,N_15846);
or U17959 (N_17959,N_16102,N_15067);
xor U17960 (N_17960,N_16279,N_16297);
and U17961 (N_17961,N_16280,N_16489);
xor U17962 (N_17962,N_16341,N_15365);
nor U17963 (N_17963,N_15241,N_15946);
and U17964 (N_17964,N_16491,N_16137);
xor U17965 (N_17965,N_16237,N_16494);
xor U17966 (N_17966,N_16498,N_16151);
or U17967 (N_17967,N_15348,N_15121);
nand U17968 (N_17968,N_15374,N_15392);
and U17969 (N_17969,N_15995,N_15661);
nand U17970 (N_17970,N_16462,N_15450);
nor U17971 (N_17971,N_15201,N_15239);
nand U17972 (N_17972,N_15821,N_16248);
nor U17973 (N_17973,N_16045,N_15816);
or U17974 (N_17974,N_16246,N_15261);
xor U17975 (N_17975,N_15134,N_15521);
nand U17976 (N_17976,N_16123,N_15961);
or U17977 (N_17977,N_15943,N_15180);
and U17978 (N_17978,N_15381,N_15845);
nor U17979 (N_17979,N_15612,N_15370);
and U17980 (N_17980,N_15181,N_15698);
nor U17981 (N_17981,N_15381,N_15058);
xnor U17982 (N_17982,N_15001,N_15813);
nand U17983 (N_17983,N_16082,N_16291);
xor U17984 (N_17984,N_15089,N_15436);
nor U17985 (N_17985,N_15982,N_15225);
nand U17986 (N_17986,N_16001,N_15090);
and U17987 (N_17987,N_16445,N_16106);
or U17988 (N_17988,N_15211,N_15877);
nand U17989 (N_17989,N_16290,N_15818);
xor U17990 (N_17990,N_15161,N_15578);
nor U17991 (N_17991,N_16033,N_15224);
nand U17992 (N_17992,N_15521,N_15377);
nor U17993 (N_17993,N_15266,N_16473);
or U17994 (N_17994,N_15947,N_15239);
or U17995 (N_17995,N_15804,N_15553);
nor U17996 (N_17996,N_16016,N_15050);
nand U17997 (N_17997,N_15957,N_15598);
and U17998 (N_17998,N_16050,N_15179);
and U17999 (N_17999,N_15170,N_15792);
xnor U18000 (N_18000,N_17751,N_17783);
nand U18001 (N_18001,N_17288,N_17667);
nand U18002 (N_18002,N_17886,N_17771);
xnor U18003 (N_18003,N_16983,N_17488);
or U18004 (N_18004,N_16921,N_17290);
or U18005 (N_18005,N_17407,N_17187);
xor U18006 (N_18006,N_16932,N_16667);
and U18007 (N_18007,N_16890,N_17547);
nand U18008 (N_18008,N_17732,N_17349);
xnor U18009 (N_18009,N_16939,N_16869);
nand U18010 (N_18010,N_17515,N_17276);
nor U18011 (N_18011,N_17611,N_17089);
or U18012 (N_18012,N_17400,N_17500);
nand U18013 (N_18013,N_16982,N_17970);
nor U18014 (N_18014,N_16878,N_17828);
and U18015 (N_18015,N_17758,N_17412);
nor U18016 (N_18016,N_16906,N_16828);
nand U18017 (N_18017,N_17922,N_17910);
xnor U18018 (N_18018,N_16537,N_17733);
nor U18019 (N_18019,N_16898,N_17190);
nor U18020 (N_18020,N_16839,N_17087);
xor U18021 (N_18021,N_16822,N_16716);
xor U18022 (N_18022,N_17084,N_16611);
nand U18023 (N_18023,N_16666,N_17120);
nor U18024 (N_18024,N_17062,N_16953);
and U18025 (N_18025,N_16527,N_17868);
nand U18026 (N_18026,N_16914,N_17191);
nand U18027 (N_18027,N_17449,N_17620);
nor U18028 (N_18028,N_16686,N_17638);
nor U18029 (N_18029,N_17273,N_17432);
nor U18030 (N_18030,N_17720,N_17919);
xnor U18031 (N_18031,N_17865,N_17260);
and U18032 (N_18032,N_17074,N_17607);
xnor U18033 (N_18033,N_16560,N_17477);
nand U18034 (N_18034,N_17418,N_17567);
nand U18035 (N_18035,N_17099,N_17197);
nand U18036 (N_18036,N_17364,N_17461);
nand U18037 (N_18037,N_17007,N_16947);
and U18038 (N_18038,N_16991,N_16619);
nor U18039 (N_18039,N_17148,N_17929);
or U18040 (N_18040,N_17544,N_17326);
or U18041 (N_18041,N_16661,N_17822);
xor U18042 (N_18042,N_16863,N_16808);
nor U18043 (N_18043,N_17646,N_16987);
xnor U18044 (N_18044,N_17269,N_16996);
nor U18045 (N_18045,N_17000,N_17870);
xnor U18046 (N_18046,N_17329,N_16521);
xnor U18047 (N_18047,N_17813,N_17243);
and U18048 (N_18048,N_17593,N_17641);
xnor U18049 (N_18049,N_17416,N_17127);
xor U18050 (N_18050,N_17721,N_17832);
nand U18051 (N_18051,N_16500,N_17305);
or U18052 (N_18052,N_16675,N_17272);
nor U18053 (N_18053,N_16931,N_16979);
xor U18054 (N_18054,N_16706,N_17592);
xor U18055 (N_18055,N_17845,N_17314);
and U18056 (N_18056,N_17092,N_17510);
or U18057 (N_18057,N_17268,N_17601);
nor U18058 (N_18058,N_17403,N_17614);
nor U18059 (N_18059,N_16951,N_17193);
nand U18060 (N_18060,N_16781,N_17212);
and U18061 (N_18061,N_17222,N_17093);
and U18062 (N_18062,N_17158,N_17053);
or U18063 (N_18063,N_17178,N_17583);
and U18064 (N_18064,N_17317,N_17621);
and U18065 (N_18065,N_17737,N_16606);
nor U18066 (N_18066,N_16962,N_17256);
nand U18067 (N_18067,N_17275,N_16782);
or U18068 (N_18068,N_17220,N_16620);
and U18069 (N_18069,N_17430,N_16720);
and U18070 (N_18070,N_17591,N_16817);
nand U18071 (N_18071,N_17226,N_16819);
or U18072 (N_18072,N_16602,N_17224);
xor U18073 (N_18073,N_17232,N_16566);
or U18074 (N_18074,N_17128,N_16525);
and U18075 (N_18075,N_17896,N_16629);
nor U18076 (N_18076,N_16825,N_17951);
nand U18077 (N_18077,N_17686,N_17787);
xnor U18078 (N_18078,N_17457,N_16758);
nand U18079 (N_18079,N_17453,N_17709);
or U18080 (N_18080,N_17112,N_17223);
and U18081 (N_18081,N_17928,N_16844);
or U18082 (N_18082,N_17790,N_16829);
or U18083 (N_18083,N_17930,N_17377);
nand U18084 (N_18084,N_17631,N_16649);
or U18085 (N_18085,N_17892,N_17316);
xor U18086 (N_18086,N_17576,N_17878);
xnor U18087 (N_18087,N_17693,N_16528);
nor U18088 (N_18088,N_16504,N_17078);
nand U18089 (N_18089,N_16816,N_16992);
and U18090 (N_18090,N_17997,N_17494);
nor U18091 (N_18091,N_17509,N_17956);
and U18092 (N_18092,N_17059,N_16514);
nand U18093 (N_18093,N_16793,N_16920);
and U18094 (N_18094,N_17531,N_17271);
or U18095 (N_18095,N_17634,N_17152);
nand U18096 (N_18096,N_17935,N_17069);
nor U18097 (N_18097,N_17528,N_16830);
xor U18098 (N_18098,N_16506,N_17300);
xnor U18099 (N_18099,N_17436,N_17283);
nor U18100 (N_18100,N_17451,N_16807);
or U18101 (N_18101,N_17789,N_17920);
nor U18102 (N_18102,N_17114,N_17372);
and U18103 (N_18103,N_17924,N_17331);
nand U18104 (N_18104,N_16981,N_17570);
xnor U18105 (N_18105,N_17590,N_17360);
nor U18106 (N_18106,N_17119,N_17802);
xor U18107 (N_18107,N_16750,N_17881);
nor U18108 (N_18108,N_16895,N_17140);
nand U18109 (N_18109,N_16590,N_17839);
nor U18110 (N_18110,N_17947,N_17218);
nor U18111 (N_18111,N_17976,N_17773);
nand U18112 (N_18112,N_16763,N_16545);
and U18113 (N_18113,N_17766,N_17991);
nor U18114 (N_18114,N_17060,N_16700);
or U18115 (N_18115,N_17526,N_17473);
nand U18116 (N_18116,N_17350,N_17653);
nor U18117 (N_18117,N_17309,N_17524);
nor U18118 (N_18118,N_17475,N_17808);
nand U18119 (N_18119,N_17353,N_17677);
xnor U18120 (N_18120,N_16569,N_16744);
xor U18121 (N_18121,N_17707,N_17033);
nand U18122 (N_18122,N_17998,N_16613);
and U18123 (N_18123,N_17036,N_16645);
and U18124 (N_18124,N_16964,N_17841);
nand U18125 (N_18125,N_16880,N_17810);
nor U18126 (N_18126,N_17303,N_17995);
nand U18127 (N_18127,N_16938,N_17957);
and U18128 (N_18128,N_16955,N_16591);
xor U18129 (N_18129,N_17444,N_16838);
nand U18130 (N_18130,N_17577,N_17723);
nor U18131 (N_18131,N_17645,N_17625);
xor U18132 (N_18132,N_17126,N_16974);
or U18133 (N_18133,N_16636,N_16553);
nor U18134 (N_18134,N_17393,N_17067);
or U18135 (N_18135,N_16954,N_16815);
or U18136 (N_18136,N_17167,N_17934);
nand U18137 (N_18137,N_17949,N_16865);
nand U18138 (N_18138,N_17312,N_16638);
nor U18139 (N_18139,N_16940,N_17748);
nand U18140 (N_18140,N_16663,N_17792);
and U18141 (N_18141,N_16845,N_16797);
xnor U18142 (N_18142,N_17107,N_17565);
nor U18143 (N_18143,N_16631,N_17972);
and U18144 (N_18144,N_16729,N_17031);
nor U18145 (N_18145,N_17992,N_17405);
nor U18146 (N_18146,N_17295,N_16725);
nor U18147 (N_18147,N_17354,N_16988);
and U18148 (N_18148,N_17159,N_17237);
or U18149 (N_18149,N_17980,N_17698);
nand U18150 (N_18150,N_16710,N_17936);
and U18151 (N_18151,N_17803,N_17595);
and U18152 (N_18152,N_16643,N_17826);
nand U18153 (N_18153,N_17780,N_17566);
xor U18154 (N_18154,N_16832,N_17108);
and U18155 (N_18155,N_17355,N_16544);
or U18156 (N_18156,N_16733,N_16640);
or U18157 (N_18157,N_17977,N_16579);
xnor U18158 (N_18158,N_17145,N_16775);
and U18159 (N_18159,N_17796,N_17013);
and U18160 (N_18160,N_17043,N_17993);
nor U18161 (N_18161,N_17888,N_16507);
nand U18162 (N_18162,N_17616,N_17650);
xor U18163 (N_18163,N_17753,N_16884);
or U18164 (N_18164,N_16668,N_17111);
nand U18165 (N_18165,N_17666,N_17613);
and U18166 (N_18166,N_17959,N_16572);
and U18167 (N_18167,N_16670,N_17437);
xor U18168 (N_18168,N_17076,N_17724);
xor U18169 (N_18169,N_16599,N_16760);
nor U18170 (N_18170,N_17287,N_17550);
nor U18171 (N_18171,N_17632,N_17670);
and U18172 (N_18172,N_17537,N_16912);
and U18173 (N_18173,N_17628,N_17551);
and U18174 (N_18174,N_17011,N_16823);
nand U18175 (N_18175,N_17596,N_17768);
and U18176 (N_18176,N_17603,N_17851);
xor U18177 (N_18177,N_17923,N_16766);
xnor U18178 (N_18178,N_17756,N_17793);
nand U18179 (N_18179,N_16646,N_16798);
and U18180 (N_18180,N_17296,N_17482);
and U18181 (N_18181,N_17597,N_17738);
and U18182 (N_18182,N_17688,N_17410);
and U18183 (N_18183,N_16524,N_17156);
nor U18184 (N_18184,N_17985,N_17598);
or U18185 (N_18185,N_17521,N_17209);
xor U18186 (N_18186,N_16586,N_16770);
nor U18187 (N_18187,N_17830,N_17659);
nand U18188 (N_18188,N_16723,N_17447);
xnor U18189 (N_18189,N_16576,N_17216);
and U18190 (N_18190,N_16834,N_16764);
xor U18191 (N_18191,N_17760,N_17857);
nand U18192 (N_18192,N_17887,N_17710);
nand U18193 (N_18193,N_17366,N_17090);
xor U18194 (N_18194,N_17495,N_16598);
and U18195 (N_18195,N_16887,N_16627);
or U18196 (N_18196,N_16737,N_17825);
and U18197 (N_18197,N_17138,N_17278);
and U18198 (N_18198,N_17974,N_17681);
xor U18199 (N_18199,N_17533,N_17622);
nand U18200 (N_18200,N_17683,N_16874);
xnor U18201 (N_18201,N_17065,N_17425);
xnor U18202 (N_18202,N_17781,N_17859);
nand U18203 (N_18203,N_17012,N_17088);
nor U18204 (N_18204,N_17195,N_16847);
nor U18205 (N_18205,N_16900,N_17261);
and U18206 (N_18206,N_17882,N_17945);
nor U18207 (N_18207,N_17522,N_16600);
or U18208 (N_18208,N_16945,N_17361);
and U18209 (N_18209,N_16818,N_17807);
and U18210 (N_18210,N_17440,N_16742);
or U18211 (N_18211,N_16583,N_16897);
or U18212 (N_18212,N_16970,N_16989);
and U18213 (N_18213,N_16980,N_17340);
xnor U18214 (N_18214,N_17809,N_16969);
xnor U18215 (N_18215,N_17151,N_17179);
nand U18216 (N_18216,N_17755,N_16730);
and U18217 (N_18217,N_17101,N_17814);
nand U18218 (N_18218,N_17198,N_16849);
nor U18219 (N_18219,N_17042,N_17313);
xnor U18220 (N_18220,N_17502,N_17767);
nor U18221 (N_18221,N_17530,N_16871);
and U18222 (N_18222,N_16573,N_16685);
xnor U18223 (N_18223,N_17694,N_17030);
xnor U18224 (N_18224,N_16997,N_16549);
xor U18225 (N_18225,N_17328,N_17774);
nor U18226 (N_18226,N_17679,N_17692);
nand U18227 (N_18227,N_17820,N_16893);
nor U18228 (N_18228,N_16536,N_17912);
and U18229 (N_18229,N_16555,N_17335);
or U18230 (N_18230,N_17701,N_17916);
nand U18231 (N_18231,N_17045,N_16628);
or U18232 (N_18232,N_17499,N_17827);
nor U18233 (N_18233,N_16949,N_16713);
xor U18234 (N_18234,N_17409,N_17286);
nor U18235 (N_18235,N_17978,N_17337);
xor U18236 (N_18236,N_17989,N_17587);
nor U18237 (N_18237,N_16673,N_17899);
and U18238 (N_18238,N_17394,N_17635);
nor U18239 (N_18239,N_17389,N_17086);
nand U18240 (N_18240,N_17657,N_16747);
xnor U18241 (N_18241,N_17474,N_17162);
or U18242 (N_18242,N_16707,N_16575);
nor U18243 (N_18243,N_17381,N_17610);
xnor U18244 (N_18244,N_16718,N_16704);
and U18245 (N_18245,N_16965,N_16811);
nor U18246 (N_18246,N_16609,N_17308);
or U18247 (N_18247,N_16977,N_17623);
nand U18248 (N_18248,N_17015,N_17734);
nand U18249 (N_18249,N_17619,N_17175);
nand U18250 (N_18250,N_17096,N_16915);
and U18251 (N_18251,N_16772,N_16712);
and U18252 (N_18252,N_17382,N_17266);
nor U18253 (N_18253,N_17588,N_16681);
and U18254 (N_18254,N_17471,N_17948);
nand U18255 (N_18255,N_17208,N_17081);
and U18256 (N_18256,N_16625,N_17519);
or U18257 (N_18257,N_16754,N_17426);
nand U18258 (N_18258,N_16547,N_17306);
xor U18259 (N_18259,N_16872,N_16526);
or U18260 (N_18260,N_17456,N_17343);
and U18261 (N_18261,N_16593,N_17523);
xor U18262 (N_18262,N_16642,N_17624);
nand U18263 (N_18263,N_17068,N_17445);
xor U18264 (N_18264,N_17648,N_17571);
nand U18265 (N_18265,N_16836,N_17245);
xor U18266 (N_18266,N_17911,N_17246);
and U18267 (N_18267,N_17134,N_17630);
xor U18268 (N_18268,N_17754,N_17640);
nand U18269 (N_18269,N_17302,N_17493);
xnor U18270 (N_18270,N_17016,N_17580);
xnor U18271 (N_18271,N_17219,N_17722);
and U18272 (N_18272,N_17772,N_17642);
nand U18273 (N_18273,N_17250,N_17898);
or U18274 (N_18274,N_17417,N_16570);
nand U18275 (N_18275,N_16655,N_17582);
or U18276 (N_18276,N_17536,N_17066);
xnor U18277 (N_18277,N_17357,N_16867);
and U18278 (N_18278,N_16594,N_17029);
and U18279 (N_18279,N_17113,N_17649);
or U18280 (N_18280,N_17231,N_16891);
nand U18281 (N_18281,N_17885,N_16904);
nand U18282 (N_18282,N_16944,N_17804);
and U18283 (N_18283,N_17821,N_17540);
nand U18284 (N_18284,N_16892,N_16703);
nor U18285 (N_18285,N_17265,N_17740);
and U18286 (N_18286,N_16903,N_17687);
xnor U18287 (N_18287,N_17166,N_17284);
and U18288 (N_18288,N_16896,N_17952);
or U18289 (N_18289,N_17664,N_17719);
and U18290 (N_18290,N_17183,N_17546);
nor U18291 (N_18291,N_16952,N_17848);
nor U18292 (N_18292,N_16910,N_16672);
nand U18293 (N_18293,N_17873,N_17342);
and U18294 (N_18294,N_17652,N_17946);
and U18295 (N_18295,N_17291,N_17319);
xor U18296 (N_18296,N_17044,N_16581);
nand U18297 (N_18297,N_16790,N_17600);
and U18298 (N_18298,N_16632,N_17429);
nor U18299 (N_18299,N_17806,N_17396);
nand U18300 (N_18300,N_17019,N_17174);
xnor U18301 (N_18301,N_17020,N_17795);
and U18302 (N_18302,N_16842,N_17564);
and U18303 (N_18303,N_17717,N_17380);
xnor U18304 (N_18304,N_16559,N_17371);
and U18305 (N_18305,N_17230,N_17647);
or U18306 (N_18306,N_17501,N_17629);
nor U18307 (N_18307,N_17121,N_17491);
xor U18308 (N_18308,N_17263,N_17633);
nor U18309 (N_18309,N_17759,N_17146);
or U18310 (N_18310,N_17039,N_17214);
xor U18311 (N_18311,N_16926,N_16533);
or U18312 (N_18312,N_17866,N_17233);
nand U18313 (N_18313,N_17324,N_17026);
xnor U18314 (N_18314,N_17712,N_17289);
or U18315 (N_18315,N_17439,N_16935);
or U18316 (N_18316,N_16922,N_17966);
or U18317 (N_18317,N_17805,N_17292);
xnor U18318 (N_18318,N_17858,N_17154);
or U18319 (N_18319,N_17915,N_16616);
nand U18320 (N_18320,N_17040,N_17661);
nand U18321 (N_18321,N_17904,N_17215);
or U18322 (N_18322,N_17070,N_16595);
nor U18323 (N_18323,N_17763,N_17006);
nor U18324 (N_18324,N_16868,N_17572);
nor U18325 (N_18325,N_17708,N_17125);
xnor U18326 (N_18326,N_17902,N_17569);
nor U18327 (N_18327,N_16956,N_17498);
or U18328 (N_18328,N_17367,N_17579);
nand U18329 (N_18329,N_17847,N_16662);
and U18330 (N_18330,N_17744,N_16837);
xor U18331 (N_18331,N_16588,N_16928);
nor U18332 (N_18332,N_17351,N_17508);
or U18333 (N_18333,N_17055,N_16833);
or U18334 (N_18334,N_16959,N_17248);
nand U18335 (N_18335,N_16578,N_17749);
or U18336 (N_18336,N_17718,N_16788);
or U18337 (N_18337,N_17189,N_16711);
and U18338 (N_18338,N_16810,N_17446);
and U18339 (N_18339,N_17942,N_17987);
or U18340 (N_18340,N_17251,N_17983);
xor U18341 (N_18341,N_17889,N_17129);
nor U18342 (N_18342,N_16881,N_16902);
nand U18343 (N_18343,N_17815,N_16736);
xor U18344 (N_18344,N_16794,N_16624);
nor U18345 (N_18345,N_17842,N_17095);
nand U18346 (N_18346,N_17714,N_17347);
nor U18347 (N_18347,N_16683,N_16513);
and U18348 (N_18348,N_16592,N_17257);
nor U18349 (N_18349,N_16787,N_17050);
xnor U18350 (N_18350,N_17901,N_17585);
nor U18351 (N_18351,N_17404,N_17010);
xnor U18352 (N_18352,N_17655,N_17321);
and U18353 (N_18353,N_17383,N_16659);
xor U18354 (N_18354,N_17241,N_16757);
or U18355 (N_18355,N_16994,N_16759);
nand U18356 (N_18356,N_17205,N_17696);
or U18357 (N_18357,N_17702,N_16615);
or U18358 (N_18358,N_16950,N_16674);
nand U18359 (N_18359,N_17589,N_17665);
nor U18360 (N_18360,N_17575,N_17034);
nand U18361 (N_18361,N_16966,N_17227);
nand U18362 (N_18362,N_17812,N_16857);
xnor U18363 (N_18363,N_16905,N_17336);
and U18364 (N_18364,N_17764,N_17411);
or U18365 (N_18365,N_16948,N_17188);
and U18366 (N_18366,N_16773,N_17875);
and U18367 (N_18367,N_17906,N_16585);
nand U18368 (N_18368,N_17549,N_17235);
and U18369 (N_18369,N_17448,N_17713);
nand U18370 (N_18370,N_16690,N_17786);
and U18371 (N_18371,N_17164,N_17489);
and U18372 (N_18372,N_17395,N_16864);
xor U18373 (N_18373,N_17855,N_17176);
nand U18374 (N_18374,N_17467,N_16925);
nand U18375 (N_18375,N_17891,N_17204);
xor U18376 (N_18376,N_17542,N_17385);
xor U18377 (N_18377,N_17890,N_17797);
nor U18378 (N_18378,N_17003,N_17727);
or U18379 (N_18379,N_17264,N_17990);
nand U18380 (N_18380,N_17478,N_17561);
xor U18381 (N_18381,N_16806,N_17373);
nand U18382 (N_18382,N_17777,N_16508);
and U18383 (N_18383,N_17386,N_17856);
xnor U18384 (N_18384,N_17527,N_17085);
or U18385 (N_18385,N_17153,N_16777);
and U18386 (N_18386,N_17715,N_16501);
or U18387 (N_18387,N_17578,N_17413);
nor U18388 (N_18388,N_17075,N_16567);
and U18389 (N_18389,N_17487,N_17184);
nand U18390 (N_18390,N_17017,N_16622);
nand U18391 (N_18391,N_17455,N_17917);
nand U18392 (N_18392,N_17518,N_16677);
nand U18393 (N_18393,N_17211,N_17027);
xor U18394 (N_18394,N_16603,N_17525);
xnor U18395 (N_18395,N_16582,N_17926);
xnor U18396 (N_18396,N_17757,N_16692);
nand U18397 (N_18397,N_16705,N_16739);
nand U18398 (N_18398,N_16973,N_17048);
xor U18399 (N_18399,N_17047,N_17770);
nand U18400 (N_18400,N_17716,N_17548);
nand U18401 (N_18401,N_17669,N_17893);
and U18402 (N_18402,N_17676,N_17318);
xnor U18403 (N_18403,N_16557,N_17529);
nor U18404 (N_18404,N_17492,N_17105);
nor U18405 (N_18405,N_17249,N_17077);
nand U18406 (N_18406,N_16552,N_17333);
nor U18407 (N_18407,N_16639,N_16676);
or U18408 (N_18408,N_16605,N_17950);
xor U18409 (N_18409,N_17872,N_16937);
and U18410 (N_18410,N_17674,N_17969);
xor U18411 (N_18411,N_16924,N_17562);
and U18412 (N_18412,N_16743,N_16546);
nor U18413 (N_18413,N_17867,N_17532);
nor U18414 (N_18414,N_16913,N_16765);
nor U18415 (N_18415,N_17979,N_17109);
nand U18416 (N_18416,N_17267,N_17160);
or U18417 (N_18417,N_17330,N_17869);
nand U18418 (N_18418,N_17785,N_16853);
and U18419 (N_18419,N_16843,N_17862);
nor U18420 (N_18420,N_17021,N_17791);
xnor U18421 (N_18421,N_17481,N_17379);
nor U18422 (N_18422,N_16774,N_17880);
and U18423 (N_18423,N_16534,N_17141);
or U18424 (N_18424,N_17051,N_17463);
nand U18425 (N_18425,N_17293,N_16732);
nor U18426 (N_18426,N_17434,N_17046);
or U18427 (N_18427,N_17513,N_17541);
nand U18428 (N_18428,N_17836,N_17871);
and U18429 (N_18429,N_17079,N_16540);
xor U18430 (N_18430,N_16637,N_17057);
nand U18431 (N_18431,N_16799,N_17225);
nand U18432 (N_18432,N_17699,N_17169);
and U18433 (N_18433,N_17484,N_16584);
or U18434 (N_18434,N_17943,N_16708);
nand U18435 (N_18435,N_16587,N_17091);
nor U18436 (N_18436,N_16614,N_17940);
xor U18437 (N_18437,N_16516,N_16522);
xnor U18438 (N_18438,N_16800,N_17639);
and U18439 (N_18439,N_17742,N_16976);
and U18440 (N_18440,N_17516,N_16551);
and U18441 (N_18441,N_17480,N_16610);
xor U18442 (N_18442,N_17961,N_17363);
and U18443 (N_18443,N_17672,N_17255);
or U18444 (N_18444,N_16715,N_17462);
nand U18445 (N_18445,N_16985,N_17356);
or U18446 (N_18446,N_17874,N_17776);
nor U18447 (N_18447,N_16679,N_17282);
and U18448 (N_18448,N_17654,N_17964);
nor U18449 (N_18449,N_16568,N_16907);
or U18450 (N_18450,N_17894,N_17769);
xnor U18451 (N_18451,N_17765,N_16734);
or U18452 (N_18452,N_17304,N_17643);
nor U18453 (N_18453,N_17252,N_17194);
or U18454 (N_18454,N_17837,N_17483);
nand U18455 (N_18455,N_17103,N_17925);
nand U18456 (N_18456,N_16535,N_17636);
or U18457 (N_18457,N_17311,N_16728);
or U18458 (N_18458,N_16888,N_16856);
nor U18459 (N_18459,N_17270,N_17281);
and U18460 (N_18460,N_17939,N_17903);
xnor U18461 (N_18461,N_17280,N_17504);
nand U18462 (N_18462,N_17254,N_17374);
nand U18463 (N_18463,N_16776,N_17999);
and U18464 (N_18464,N_16580,N_17102);
and U18465 (N_18465,N_17346,N_17782);
xnor U18466 (N_18466,N_17035,N_16740);
nor U18467 (N_18467,N_16917,N_17323);
and U18468 (N_18468,N_17644,N_16517);
or U18469 (N_18469,N_17049,N_17967);
and U18470 (N_18470,N_16556,N_16756);
and U18471 (N_18471,N_17008,N_17853);
nor U18472 (N_18472,N_17517,N_16682);
or U18473 (N_18473,N_17391,N_16824);
or U18474 (N_18474,N_16565,N_16644);
nand U18475 (N_18475,N_17401,N_17149);
nand U18476 (N_18476,N_16696,N_16827);
and U18477 (N_18477,N_17507,N_16660);
and U18478 (N_18478,N_16509,N_16751);
xor U18479 (N_18479,N_17838,N_16768);
or U18480 (N_18480,N_17420,N_17799);
nor U18481 (N_18481,N_17794,N_16698);
nor U18482 (N_18482,N_17442,N_17450);
xnor U18483 (N_18483,N_16911,N_17490);
nand U18484 (N_18484,N_17143,N_17443);
xor U18485 (N_18485,N_17852,N_16873);
nand U18486 (N_18486,N_17711,N_16647);
and U18487 (N_18487,N_17207,N_17421);
and U18488 (N_18488,N_16943,N_16652);
or U18489 (N_18489,N_17344,N_17656);
nand U18490 (N_18490,N_17554,N_17009);
xnor U18491 (N_18491,N_16597,N_17390);
nor U18492 (N_18492,N_17466,N_16748);
nand U18493 (N_18493,N_17900,N_16654);
nand U18494 (N_18494,N_16826,N_16876);
or U18495 (N_18495,N_17063,N_17277);
nor U18496 (N_18496,N_17663,N_17937);
and U18497 (N_18497,N_16804,N_17298);
xnor U18498 (N_18498,N_17726,N_17496);
nand U18499 (N_18499,N_17135,N_16780);
and U18500 (N_18500,N_16618,N_17725);
nor U18501 (N_18501,N_17229,N_16762);
nor U18502 (N_18502,N_17163,N_17840);
xnor U18503 (N_18503,N_16866,N_16721);
xnor U18504 (N_18504,N_17118,N_17365);
xnor U18505 (N_18505,N_16852,N_17459);
xnor U18506 (N_18506,N_17362,N_16995);
nor U18507 (N_18507,N_17428,N_17514);
and U18508 (N_18508,N_17690,N_17944);
nand U18509 (N_18509,N_17685,N_16571);
nor U18510 (N_18510,N_17778,N_16812);
xnor U18511 (N_18511,N_17028,N_17376);
nand U18512 (N_18512,N_17730,N_17877);
nor U18513 (N_18513,N_17824,N_17743);
nand U18514 (N_18514,N_17876,N_16651);
nand U18515 (N_18515,N_17637,N_17370);
or U18516 (N_18516,N_17419,N_17700);
or U18517 (N_18517,N_17503,N_17986);
nor U18518 (N_18518,N_16848,N_16741);
nand U18519 (N_18519,N_17627,N_16820);
xor U18520 (N_18520,N_16862,N_17083);
or U18521 (N_18521,N_17139,N_17762);
or U18522 (N_18522,N_17788,N_17973);
nor U18523 (N_18523,N_17913,N_17071);
and U18524 (N_18524,N_17602,N_17180);
nand U18525 (N_18525,N_16870,N_16785);
nand U18526 (N_18526,N_17752,N_17801);
and U18527 (N_18527,N_16731,N_17157);
and U18528 (N_18528,N_17918,N_17941);
or U18529 (N_18529,N_17673,N_17253);
nor U18530 (N_18530,N_16529,N_16719);
xnor U18531 (N_18531,N_17130,N_17996);
and U18532 (N_18532,N_17122,N_17558);
and U18533 (N_18533,N_16745,N_17779);
nand U18534 (N_18534,N_17662,N_17322);
or U18535 (N_18535,N_17199,N_16564);
nand U18536 (N_18536,N_17294,N_17117);
nand U18537 (N_18537,N_16877,N_17604);
or U18538 (N_18538,N_17884,N_17962);
nand U18539 (N_18539,N_17921,N_17606);
or U18540 (N_18540,N_17556,N_17080);
or U18541 (N_18541,N_17106,N_17750);
nand U18542 (N_18542,N_16783,N_17142);
nand U18543 (N_18543,N_17240,N_17001);
nand U18544 (N_18544,N_17505,N_16635);
xnor U18545 (N_18545,N_17689,N_17131);
xnor U18546 (N_18546,N_16669,N_17775);
or U18547 (N_18547,N_16523,N_16680);
xor U18548 (N_18548,N_16805,N_16548);
nand U18549 (N_18549,N_16554,N_17955);
and U18550 (N_18550,N_16753,N_17186);
and U18551 (N_18551,N_17818,N_17338);
nand U18552 (N_18552,N_16854,N_17684);
nand U18553 (N_18553,N_17835,N_16778);
and U18554 (N_18554,N_17058,N_17668);
nor U18555 (N_18555,N_16971,N_16650);
and U18556 (N_18556,N_17965,N_16879);
or U18557 (N_18557,N_17147,N_16531);
nand U18558 (N_18558,N_17022,N_17861);
nor U18559 (N_18559,N_17054,N_17052);
or U18560 (N_18560,N_16755,N_17746);
and U18561 (N_18561,N_16998,N_17441);
xnor U18562 (N_18562,N_17651,N_16695);
and U18563 (N_18563,N_17399,N_17234);
nand U18564 (N_18564,N_17850,N_16861);
nor U18565 (N_18565,N_17975,N_16786);
nand U18566 (N_18566,N_17392,N_17626);
or U18567 (N_18567,N_16701,N_16779);
or U18568 (N_18568,N_17538,N_17297);
nand U18569 (N_18569,N_17422,N_17301);
xor U18570 (N_18570,N_17170,N_17931);
or U18571 (N_18571,N_16738,N_16761);
nand U18572 (N_18572,N_16941,N_17883);
nor U18573 (N_18573,N_16539,N_17747);
nand U18574 (N_18574,N_17658,N_17932);
xor U18575 (N_18575,N_17217,N_16821);
xor U18576 (N_18576,N_17981,N_16678);
xor U18577 (N_18577,N_16831,N_17560);
nand U18578 (N_18578,N_16769,N_17543);
nand U18579 (N_18579,N_16543,N_17221);
nand U18580 (N_18580,N_17691,N_17553);
nor U18581 (N_18581,N_16801,N_17454);
or U18582 (N_18582,N_16607,N_17279);
and U18583 (N_18583,N_17994,N_16978);
and U18584 (N_18584,N_17479,N_17433);
nor U18585 (N_18585,N_16752,N_16883);
xnor U18586 (N_18586,N_17023,N_17675);
nor U18587 (N_18587,N_17458,N_16860);
xnor U18588 (N_18588,N_16601,N_17056);
xor U18589 (N_18589,N_17615,N_17415);
nand U18590 (N_18590,N_16671,N_16960);
and U18591 (N_18591,N_17552,N_17061);
nor U18592 (N_18592,N_16512,N_17327);
xnor U18593 (N_18593,N_17609,N_17506);
and U18594 (N_18594,N_16889,N_17435);
nand U18595 (N_18595,N_17954,N_17299);
nor U18596 (N_18596,N_17739,N_16727);
xnor U18597 (N_18597,N_16664,N_16617);
nor U18598 (N_18598,N_17823,N_17005);
xor U18599 (N_18599,N_17860,N_16658);
nand U18600 (N_18600,N_17368,N_17247);
xor U18601 (N_18601,N_17414,N_16814);
or U18602 (N_18602,N_16919,N_16722);
xor U18603 (N_18603,N_16608,N_17239);
xnor U18604 (N_18604,N_17206,N_16558);
or U18605 (N_18605,N_17242,N_17895);
and U18606 (N_18606,N_17817,N_16702);
and U18607 (N_18607,N_16541,N_17469);
nor U18608 (N_18608,N_16851,N_17854);
or U18609 (N_18609,N_17037,N_17397);
xor U18610 (N_18610,N_17695,N_17369);
nand U18611 (N_18611,N_17398,N_17038);
nor U18612 (N_18612,N_17563,N_16621);
nor U18613 (N_18613,N_17172,N_17897);
nor U18614 (N_18614,N_17472,N_17660);
xnor U18615 (N_18615,N_16724,N_17465);
and U18616 (N_18616,N_16909,N_16641);
or U18617 (N_18617,N_17497,N_17960);
xor U18618 (N_18618,N_17310,N_17002);
or U18619 (N_18619,N_17704,N_17617);
or U18620 (N_18620,N_17082,N_16532);
xnor U18621 (N_18621,N_17697,N_16596);
or U18622 (N_18622,N_16767,N_17375);
xor U18623 (N_18623,N_16936,N_17608);
and U18624 (N_18624,N_17200,N_17161);
nand U18625 (N_18625,N_16795,N_16930);
or U18626 (N_18626,N_17819,N_16612);
and U18627 (N_18627,N_16519,N_16946);
xor U18628 (N_18628,N_17334,N_16665);
and U18629 (N_18629,N_17816,N_17171);
nand U18630 (N_18630,N_16693,N_17203);
and U18631 (N_18631,N_17238,N_16542);
xor U18632 (N_18632,N_17144,N_17905);
nor U18633 (N_18633,N_17307,N_16850);
and U18634 (N_18634,N_16993,N_16840);
nand U18635 (N_18635,N_17798,N_17339);
nand U18636 (N_18636,N_16923,N_16520);
xor U18637 (N_18637,N_17460,N_17844);
xor U18638 (N_18638,N_16746,N_17424);
nor U18639 (N_18639,N_16975,N_17618);
xor U18640 (N_18640,N_16934,N_17938);
nor U18641 (N_18641,N_17511,N_16589);
nand U18642 (N_18642,N_17953,N_16894);
and U18643 (N_18643,N_17914,N_17784);
xor U18644 (N_18644,N_16859,N_17133);
or U18645 (N_18645,N_17682,N_17064);
nor U18646 (N_18646,N_17341,N_17387);
xor U18647 (N_18647,N_17116,N_17406);
nand U18648 (N_18648,N_17388,N_17735);
nand U18649 (N_18649,N_16577,N_17464);
or U18650 (N_18650,N_16648,N_17182);
or U18651 (N_18651,N_17210,N_16518);
xor U18652 (N_18652,N_16942,N_17032);
and U18653 (N_18653,N_17402,N_16561);
nor U18654 (N_18654,N_17971,N_17908);
xnor U18655 (N_18655,N_17468,N_16999);
nor U18656 (N_18656,N_17833,N_17438);
xnor U18657 (N_18657,N_17123,N_17846);
or U18658 (N_18658,N_17320,N_17285);
nor U18659 (N_18659,N_16510,N_16901);
or U18660 (N_18660,N_16630,N_16687);
nand U18661 (N_18661,N_17907,N_17678);
nand U18662 (N_18662,N_17731,N_17427);
nor U18663 (N_18663,N_16908,N_16657);
nor U18664 (N_18664,N_16858,N_17196);
or U18665 (N_18665,N_16697,N_17181);
xnor U18666 (N_18666,N_17165,N_16963);
or U18667 (N_18667,N_16653,N_16709);
and U18668 (N_18668,N_17559,N_17982);
and U18669 (N_18669,N_16791,N_17100);
nand U18670 (N_18670,N_16574,N_17831);
nor U18671 (N_18671,N_17485,N_17018);
nor U18672 (N_18672,N_17927,N_16846);
nand U18673 (N_18673,N_17834,N_17843);
nand U18674 (N_18674,N_16633,N_17094);
and U18675 (N_18675,N_17431,N_17829);
xnor U18676 (N_18676,N_17168,N_17104);
nor U18677 (N_18677,N_16714,N_16933);
nand U18678 (N_18678,N_17680,N_16505);
nor U18679 (N_18679,N_16984,N_17706);
nor U18680 (N_18680,N_17705,N_16511);
xnor U18681 (N_18681,N_16813,N_17097);
or U18682 (N_18682,N_17024,N_17452);
nor U18683 (N_18683,N_17545,N_17863);
or U18684 (N_18684,N_17584,N_16990);
nand U18685 (N_18685,N_17259,N_17849);
nor U18686 (N_18686,N_16885,N_16841);
nand U18687 (N_18687,N_17345,N_17535);
nor U18688 (N_18688,N_16550,N_17745);
nor U18689 (N_18689,N_16562,N_17741);
nor U18690 (N_18690,N_16502,N_17408);
xor U18691 (N_18691,N_16986,N_16530);
nor U18692 (N_18692,N_17555,N_16784);
nand U18693 (N_18693,N_17202,N_17137);
nor U18694 (N_18694,N_17185,N_17599);
or U18695 (N_18695,N_16796,N_17073);
nor U18696 (N_18696,N_17072,N_17384);
nand U18697 (N_18697,N_17262,N_17568);
and U18698 (N_18698,N_17358,N_16882);
xnor U18699 (N_18699,N_17228,N_17879);
or U18700 (N_18700,N_17136,N_17811);
nand U18701 (N_18701,N_17581,N_17761);
or U18702 (N_18702,N_17728,N_17378);
xor U18703 (N_18703,N_17574,N_16875);
and U18704 (N_18704,N_16929,N_17703);
nand U18705 (N_18705,N_16855,N_16691);
and U18706 (N_18706,N_16749,N_17115);
xor U18707 (N_18707,N_17155,N_17963);
and U18708 (N_18708,N_16563,N_16958);
nand U18709 (N_18709,N_16538,N_16735);
nor U18710 (N_18710,N_17958,N_17150);
and U18711 (N_18711,N_17332,N_16916);
nand U18712 (N_18712,N_17520,N_17258);
nand U18713 (N_18713,N_17124,N_17352);
and U18714 (N_18714,N_16809,N_17864);
and U18715 (N_18715,N_16886,N_16899);
or U18716 (N_18716,N_17988,N_17132);
nor U18717 (N_18717,N_17573,N_17512);
nand U18718 (N_18718,N_16957,N_17213);
nor U18719 (N_18719,N_17984,N_16771);
nand U18720 (N_18720,N_16503,N_17177);
xnor U18721 (N_18721,N_17423,N_16694);
xnor U18722 (N_18722,N_17539,N_17014);
xnor U18723 (N_18723,N_16688,N_17325);
or U18724 (N_18724,N_17098,N_17025);
xor U18725 (N_18725,N_17110,N_16918);
nor U18726 (N_18726,N_17909,N_17470);
nor U18727 (N_18727,N_16789,N_17557);
nand U18728 (N_18728,N_16515,N_17348);
xor U18729 (N_18729,N_17476,N_17671);
nor U18730 (N_18730,N_17359,N_16689);
nand U18731 (N_18731,N_17486,N_17315);
xnor U18732 (N_18732,N_17192,N_16803);
and U18733 (N_18733,N_16792,N_16972);
nor U18734 (N_18734,N_17274,N_17800);
or U18735 (N_18735,N_17244,N_16717);
nand U18736 (N_18736,N_17729,N_17594);
nand U18737 (N_18737,N_16604,N_16656);
nand U18738 (N_18738,N_16967,N_17933);
or U18739 (N_18739,N_17041,N_17605);
nor U18740 (N_18740,N_17201,N_17968);
or U18741 (N_18741,N_17236,N_17004);
nand U18742 (N_18742,N_16968,N_16726);
nor U18743 (N_18743,N_17612,N_16634);
nand U18744 (N_18744,N_16623,N_16699);
or U18745 (N_18745,N_16835,N_17736);
and U18746 (N_18746,N_17173,N_16684);
xor U18747 (N_18747,N_17586,N_16927);
nand U18748 (N_18748,N_16626,N_16802);
or U18749 (N_18749,N_17534,N_16961);
nor U18750 (N_18750,N_17693,N_16675);
nand U18751 (N_18751,N_16670,N_17404);
or U18752 (N_18752,N_16683,N_16756);
or U18753 (N_18753,N_17087,N_17953);
nor U18754 (N_18754,N_17906,N_17360);
and U18755 (N_18755,N_17457,N_17206);
nand U18756 (N_18756,N_16658,N_17434);
nand U18757 (N_18757,N_17701,N_16891);
nor U18758 (N_18758,N_17503,N_16688);
or U18759 (N_18759,N_17040,N_16579);
nor U18760 (N_18760,N_17784,N_17285);
nand U18761 (N_18761,N_16901,N_16740);
nand U18762 (N_18762,N_16901,N_17624);
or U18763 (N_18763,N_17265,N_17827);
nand U18764 (N_18764,N_16533,N_17391);
nor U18765 (N_18765,N_17636,N_17690);
or U18766 (N_18766,N_17090,N_17936);
xor U18767 (N_18767,N_17410,N_17644);
xnor U18768 (N_18768,N_17846,N_17514);
or U18769 (N_18769,N_16577,N_16810);
xnor U18770 (N_18770,N_17076,N_17150);
nor U18771 (N_18771,N_16553,N_17220);
xor U18772 (N_18772,N_17437,N_17877);
and U18773 (N_18773,N_16826,N_16904);
and U18774 (N_18774,N_17837,N_17587);
nand U18775 (N_18775,N_17826,N_17457);
nand U18776 (N_18776,N_16676,N_17932);
nor U18777 (N_18777,N_16541,N_17414);
and U18778 (N_18778,N_17736,N_17055);
nor U18779 (N_18779,N_17886,N_16553);
xor U18780 (N_18780,N_17129,N_17344);
and U18781 (N_18781,N_17502,N_17373);
nand U18782 (N_18782,N_17333,N_17399);
xor U18783 (N_18783,N_17018,N_16765);
xnor U18784 (N_18784,N_16576,N_16902);
and U18785 (N_18785,N_17527,N_16745);
xnor U18786 (N_18786,N_17687,N_17039);
or U18787 (N_18787,N_16764,N_16570);
or U18788 (N_18788,N_17946,N_16715);
or U18789 (N_18789,N_17058,N_17536);
nand U18790 (N_18790,N_16508,N_16777);
and U18791 (N_18791,N_16799,N_17454);
or U18792 (N_18792,N_17140,N_16846);
or U18793 (N_18793,N_16727,N_17474);
nand U18794 (N_18794,N_16762,N_16829);
and U18795 (N_18795,N_17996,N_17663);
and U18796 (N_18796,N_17859,N_17810);
nor U18797 (N_18797,N_16718,N_16822);
nand U18798 (N_18798,N_17753,N_17467);
xor U18799 (N_18799,N_17600,N_17559);
xnor U18800 (N_18800,N_17718,N_17159);
or U18801 (N_18801,N_16696,N_17912);
nor U18802 (N_18802,N_16590,N_17691);
nand U18803 (N_18803,N_17056,N_17484);
and U18804 (N_18804,N_16889,N_16655);
and U18805 (N_18805,N_16829,N_16823);
nor U18806 (N_18806,N_17646,N_17494);
and U18807 (N_18807,N_17770,N_16966);
and U18808 (N_18808,N_17498,N_17710);
xor U18809 (N_18809,N_17273,N_17649);
and U18810 (N_18810,N_16771,N_17115);
nand U18811 (N_18811,N_17013,N_17051);
xor U18812 (N_18812,N_17558,N_16674);
nor U18813 (N_18813,N_17303,N_17549);
xor U18814 (N_18814,N_16619,N_16840);
xnor U18815 (N_18815,N_17005,N_16638);
nor U18816 (N_18816,N_17642,N_16954);
xor U18817 (N_18817,N_17116,N_17449);
nand U18818 (N_18818,N_16957,N_17478);
or U18819 (N_18819,N_17473,N_17206);
and U18820 (N_18820,N_17740,N_16866);
and U18821 (N_18821,N_17156,N_16820);
or U18822 (N_18822,N_17715,N_16683);
xnor U18823 (N_18823,N_17251,N_17431);
or U18824 (N_18824,N_16557,N_17619);
nor U18825 (N_18825,N_17660,N_17666);
or U18826 (N_18826,N_16997,N_17884);
nand U18827 (N_18827,N_17179,N_17020);
nand U18828 (N_18828,N_16617,N_17918);
or U18829 (N_18829,N_16745,N_17335);
or U18830 (N_18830,N_17029,N_16844);
nand U18831 (N_18831,N_17451,N_17537);
nor U18832 (N_18832,N_16930,N_16553);
xor U18833 (N_18833,N_16995,N_17566);
nor U18834 (N_18834,N_17153,N_17027);
nand U18835 (N_18835,N_17929,N_17580);
nand U18836 (N_18836,N_17322,N_16969);
or U18837 (N_18837,N_17869,N_17986);
or U18838 (N_18838,N_16885,N_17581);
or U18839 (N_18839,N_16955,N_17999);
nor U18840 (N_18840,N_17858,N_16708);
nand U18841 (N_18841,N_17258,N_17017);
and U18842 (N_18842,N_17902,N_16969);
xor U18843 (N_18843,N_17072,N_17215);
or U18844 (N_18844,N_17597,N_17515);
and U18845 (N_18845,N_17117,N_17537);
and U18846 (N_18846,N_17717,N_17682);
and U18847 (N_18847,N_17150,N_16556);
or U18848 (N_18848,N_17733,N_17524);
or U18849 (N_18849,N_17042,N_16634);
nor U18850 (N_18850,N_17840,N_16771);
nand U18851 (N_18851,N_16577,N_17500);
and U18852 (N_18852,N_16862,N_16961);
xor U18853 (N_18853,N_17784,N_17156);
or U18854 (N_18854,N_16851,N_17054);
and U18855 (N_18855,N_17925,N_17942);
and U18856 (N_18856,N_16946,N_17370);
nor U18857 (N_18857,N_17386,N_17125);
and U18858 (N_18858,N_17199,N_17404);
nor U18859 (N_18859,N_16950,N_16804);
nand U18860 (N_18860,N_17950,N_16948);
nor U18861 (N_18861,N_17539,N_17863);
xnor U18862 (N_18862,N_16742,N_17967);
and U18863 (N_18863,N_16752,N_17465);
nand U18864 (N_18864,N_16701,N_16677);
and U18865 (N_18865,N_16577,N_17928);
or U18866 (N_18866,N_17466,N_16607);
or U18867 (N_18867,N_17345,N_16761);
xnor U18868 (N_18868,N_16932,N_17198);
or U18869 (N_18869,N_17976,N_17104);
or U18870 (N_18870,N_17968,N_17473);
or U18871 (N_18871,N_16503,N_17984);
xor U18872 (N_18872,N_17431,N_17305);
and U18873 (N_18873,N_16658,N_16763);
xor U18874 (N_18874,N_16978,N_17639);
nand U18875 (N_18875,N_16586,N_17737);
or U18876 (N_18876,N_17168,N_17130);
nand U18877 (N_18877,N_17437,N_17659);
nor U18878 (N_18878,N_17478,N_16748);
or U18879 (N_18879,N_16812,N_16614);
xnor U18880 (N_18880,N_17181,N_16911);
xnor U18881 (N_18881,N_17099,N_16529);
xnor U18882 (N_18882,N_17426,N_16848);
or U18883 (N_18883,N_16906,N_16633);
xnor U18884 (N_18884,N_17764,N_17097);
or U18885 (N_18885,N_17087,N_17522);
and U18886 (N_18886,N_17310,N_16868);
nand U18887 (N_18887,N_16625,N_17927);
and U18888 (N_18888,N_17478,N_16665);
nor U18889 (N_18889,N_17672,N_16955);
or U18890 (N_18890,N_17288,N_17190);
nand U18891 (N_18891,N_17863,N_17117);
xor U18892 (N_18892,N_17854,N_16905);
or U18893 (N_18893,N_17150,N_17983);
and U18894 (N_18894,N_17506,N_17816);
xor U18895 (N_18895,N_17824,N_17656);
nor U18896 (N_18896,N_17006,N_17400);
nand U18897 (N_18897,N_17134,N_17848);
or U18898 (N_18898,N_16528,N_17085);
nor U18899 (N_18899,N_17443,N_17424);
nand U18900 (N_18900,N_17671,N_17625);
xnor U18901 (N_18901,N_17079,N_16569);
nand U18902 (N_18902,N_17155,N_17766);
nand U18903 (N_18903,N_17357,N_17398);
and U18904 (N_18904,N_17746,N_16652);
and U18905 (N_18905,N_17336,N_17127);
nor U18906 (N_18906,N_17276,N_16941);
nand U18907 (N_18907,N_17064,N_17729);
nor U18908 (N_18908,N_17473,N_17368);
nand U18909 (N_18909,N_17536,N_16697);
nand U18910 (N_18910,N_17002,N_17695);
nand U18911 (N_18911,N_17784,N_16626);
xnor U18912 (N_18912,N_17726,N_17925);
or U18913 (N_18913,N_16857,N_17668);
nand U18914 (N_18914,N_17586,N_17409);
and U18915 (N_18915,N_17624,N_17066);
and U18916 (N_18916,N_17585,N_16579);
and U18917 (N_18917,N_16963,N_16809);
nor U18918 (N_18918,N_16518,N_17194);
nand U18919 (N_18919,N_16920,N_17877);
nor U18920 (N_18920,N_17297,N_17174);
or U18921 (N_18921,N_17410,N_16739);
or U18922 (N_18922,N_17275,N_17550);
nand U18923 (N_18923,N_17454,N_17914);
nand U18924 (N_18924,N_17969,N_17679);
or U18925 (N_18925,N_17404,N_17121);
and U18926 (N_18926,N_17441,N_16730);
nand U18927 (N_18927,N_17856,N_17267);
or U18928 (N_18928,N_16861,N_17445);
xor U18929 (N_18929,N_16531,N_17890);
and U18930 (N_18930,N_16765,N_17310);
nor U18931 (N_18931,N_16584,N_16626);
xnor U18932 (N_18932,N_17550,N_17508);
and U18933 (N_18933,N_16873,N_17949);
and U18934 (N_18934,N_17625,N_17155);
and U18935 (N_18935,N_17407,N_17520);
nor U18936 (N_18936,N_17811,N_17292);
xor U18937 (N_18937,N_17648,N_16569);
nand U18938 (N_18938,N_17232,N_17929);
nor U18939 (N_18939,N_16691,N_16788);
xnor U18940 (N_18940,N_16927,N_17983);
and U18941 (N_18941,N_17365,N_16519);
and U18942 (N_18942,N_16781,N_17824);
nor U18943 (N_18943,N_17733,N_17205);
xor U18944 (N_18944,N_16596,N_17163);
or U18945 (N_18945,N_17537,N_17839);
nor U18946 (N_18946,N_17759,N_17433);
nand U18947 (N_18947,N_16985,N_16634);
nand U18948 (N_18948,N_17751,N_17175);
and U18949 (N_18949,N_17474,N_17294);
nand U18950 (N_18950,N_17063,N_16785);
or U18951 (N_18951,N_16842,N_17183);
nor U18952 (N_18952,N_17566,N_16854);
xor U18953 (N_18953,N_17070,N_17820);
xnor U18954 (N_18954,N_17007,N_17535);
nand U18955 (N_18955,N_17832,N_17897);
xor U18956 (N_18956,N_17376,N_17450);
and U18957 (N_18957,N_16599,N_17596);
and U18958 (N_18958,N_17177,N_17332);
and U18959 (N_18959,N_17346,N_16938);
and U18960 (N_18960,N_16522,N_16558);
or U18961 (N_18961,N_17390,N_17574);
xnor U18962 (N_18962,N_16979,N_17357);
or U18963 (N_18963,N_16668,N_17489);
nor U18964 (N_18964,N_16868,N_16580);
or U18965 (N_18965,N_17617,N_16784);
and U18966 (N_18966,N_16959,N_16530);
or U18967 (N_18967,N_16615,N_16740);
nand U18968 (N_18968,N_16944,N_17276);
and U18969 (N_18969,N_17010,N_17990);
xor U18970 (N_18970,N_17478,N_17948);
and U18971 (N_18971,N_17328,N_17957);
or U18972 (N_18972,N_17849,N_17118);
and U18973 (N_18973,N_17129,N_17160);
or U18974 (N_18974,N_17464,N_17785);
and U18975 (N_18975,N_16526,N_17559);
and U18976 (N_18976,N_16546,N_16607);
xnor U18977 (N_18977,N_16975,N_16536);
nand U18978 (N_18978,N_17322,N_17643);
nand U18979 (N_18979,N_17977,N_17687);
nor U18980 (N_18980,N_17935,N_16579);
or U18981 (N_18981,N_16657,N_16744);
nand U18982 (N_18982,N_17844,N_17850);
nand U18983 (N_18983,N_17022,N_17092);
nand U18984 (N_18984,N_17311,N_17987);
and U18985 (N_18985,N_17809,N_17566);
nor U18986 (N_18986,N_17946,N_17128);
nand U18987 (N_18987,N_17139,N_17454);
or U18988 (N_18988,N_17638,N_16699);
nand U18989 (N_18989,N_16792,N_17364);
or U18990 (N_18990,N_17929,N_17119);
or U18991 (N_18991,N_16848,N_17523);
xor U18992 (N_18992,N_16607,N_17768);
xor U18993 (N_18993,N_17403,N_17562);
xnor U18994 (N_18994,N_16705,N_17312);
or U18995 (N_18995,N_17373,N_17434);
nor U18996 (N_18996,N_17268,N_16580);
nor U18997 (N_18997,N_17387,N_17191);
nand U18998 (N_18998,N_17396,N_17631);
nor U18999 (N_18999,N_17349,N_16536);
xor U19000 (N_19000,N_16868,N_17147);
and U19001 (N_19001,N_17643,N_17778);
nand U19002 (N_19002,N_17462,N_17818);
nand U19003 (N_19003,N_16946,N_17407);
or U19004 (N_19004,N_17659,N_16740);
nand U19005 (N_19005,N_16730,N_16554);
xor U19006 (N_19006,N_16677,N_17081);
nand U19007 (N_19007,N_17906,N_17923);
nand U19008 (N_19008,N_16873,N_17093);
and U19009 (N_19009,N_17133,N_17893);
nand U19010 (N_19010,N_17859,N_17768);
nand U19011 (N_19011,N_17392,N_16752);
nor U19012 (N_19012,N_17685,N_16955);
nand U19013 (N_19013,N_17466,N_17241);
or U19014 (N_19014,N_16759,N_17253);
nand U19015 (N_19015,N_16985,N_17894);
nor U19016 (N_19016,N_17158,N_16986);
and U19017 (N_19017,N_16672,N_16663);
nand U19018 (N_19018,N_17554,N_17685);
nand U19019 (N_19019,N_17269,N_17626);
nor U19020 (N_19020,N_17909,N_17586);
nor U19021 (N_19021,N_17712,N_17614);
and U19022 (N_19022,N_16918,N_17084);
and U19023 (N_19023,N_16520,N_16674);
nand U19024 (N_19024,N_17421,N_16833);
and U19025 (N_19025,N_17106,N_17343);
xnor U19026 (N_19026,N_16747,N_17467);
or U19027 (N_19027,N_17837,N_17828);
nand U19028 (N_19028,N_16830,N_17770);
and U19029 (N_19029,N_17755,N_16514);
or U19030 (N_19030,N_16817,N_17322);
nand U19031 (N_19031,N_17246,N_17021);
nor U19032 (N_19032,N_17993,N_16681);
nor U19033 (N_19033,N_16837,N_17297);
nor U19034 (N_19034,N_17849,N_17422);
nand U19035 (N_19035,N_17253,N_17884);
and U19036 (N_19036,N_17986,N_17286);
and U19037 (N_19037,N_17381,N_17867);
nand U19038 (N_19038,N_17195,N_17854);
or U19039 (N_19039,N_16531,N_17154);
and U19040 (N_19040,N_16857,N_17949);
nand U19041 (N_19041,N_17577,N_16514);
xor U19042 (N_19042,N_16827,N_16654);
nor U19043 (N_19043,N_16546,N_17574);
nor U19044 (N_19044,N_16799,N_17540);
nand U19045 (N_19045,N_17583,N_17569);
nor U19046 (N_19046,N_17212,N_17415);
or U19047 (N_19047,N_16527,N_16763);
nand U19048 (N_19048,N_16766,N_17812);
or U19049 (N_19049,N_16946,N_17519);
or U19050 (N_19050,N_17437,N_16876);
or U19051 (N_19051,N_17338,N_17795);
and U19052 (N_19052,N_17939,N_17422);
or U19053 (N_19053,N_17546,N_17273);
and U19054 (N_19054,N_17013,N_17312);
and U19055 (N_19055,N_16646,N_16531);
xnor U19056 (N_19056,N_16527,N_16721);
or U19057 (N_19057,N_16622,N_16530);
nor U19058 (N_19058,N_17762,N_17973);
and U19059 (N_19059,N_17873,N_17796);
and U19060 (N_19060,N_16931,N_17978);
nand U19061 (N_19061,N_17897,N_17240);
xnor U19062 (N_19062,N_17099,N_17194);
or U19063 (N_19063,N_17779,N_17647);
or U19064 (N_19064,N_17009,N_17403);
or U19065 (N_19065,N_17773,N_16964);
nor U19066 (N_19066,N_17237,N_17323);
or U19067 (N_19067,N_17064,N_17626);
and U19068 (N_19068,N_17447,N_17875);
and U19069 (N_19069,N_17869,N_17956);
nand U19070 (N_19070,N_17176,N_17876);
nand U19071 (N_19071,N_16747,N_17582);
nor U19072 (N_19072,N_16663,N_17810);
nor U19073 (N_19073,N_16501,N_16962);
nand U19074 (N_19074,N_17802,N_17640);
nor U19075 (N_19075,N_16765,N_17304);
nor U19076 (N_19076,N_17913,N_16769);
nor U19077 (N_19077,N_17094,N_17519);
nor U19078 (N_19078,N_16736,N_16542);
nor U19079 (N_19079,N_17464,N_16778);
nand U19080 (N_19080,N_17216,N_16704);
nand U19081 (N_19081,N_17732,N_17033);
nor U19082 (N_19082,N_16741,N_16718);
nor U19083 (N_19083,N_17738,N_17405);
or U19084 (N_19084,N_17559,N_16980);
and U19085 (N_19085,N_17417,N_17967);
and U19086 (N_19086,N_16577,N_17905);
and U19087 (N_19087,N_17843,N_17635);
nor U19088 (N_19088,N_17047,N_17242);
nor U19089 (N_19089,N_17825,N_16596);
nor U19090 (N_19090,N_16773,N_17676);
xor U19091 (N_19091,N_16627,N_17878);
or U19092 (N_19092,N_17579,N_17405);
or U19093 (N_19093,N_17878,N_17847);
nand U19094 (N_19094,N_16574,N_16513);
nor U19095 (N_19095,N_17409,N_17238);
nand U19096 (N_19096,N_17936,N_17868);
or U19097 (N_19097,N_17148,N_17203);
nand U19098 (N_19098,N_17438,N_17199);
nand U19099 (N_19099,N_17955,N_17942);
xnor U19100 (N_19100,N_17111,N_17594);
and U19101 (N_19101,N_17596,N_17436);
nand U19102 (N_19102,N_16513,N_17980);
nor U19103 (N_19103,N_17144,N_17438);
nand U19104 (N_19104,N_17710,N_16688);
and U19105 (N_19105,N_17805,N_17831);
or U19106 (N_19106,N_17274,N_17039);
nor U19107 (N_19107,N_17720,N_17883);
and U19108 (N_19108,N_17618,N_16637);
and U19109 (N_19109,N_17442,N_16956);
or U19110 (N_19110,N_16611,N_17086);
nor U19111 (N_19111,N_17059,N_17281);
nand U19112 (N_19112,N_17659,N_17194);
and U19113 (N_19113,N_17498,N_17588);
nand U19114 (N_19114,N_17502,N_17577);
xnor U19115 (N_19115,N_16690,N_16678);
nor U19116 (N_19116,N_17164,N_17565);
nor U19117 (N_19117,N_17957,N_16646);
or U19118 (N_19118,N_16722,N_17756);
xnor U19119 (N_19119,N_17996,N_17260);
nand U19120 (N_19120,N_17533,N_17073);
nor U19121 (N_19121,N_17457,N_17302);
and U19122 (N_19122,N_16719,N_17516);
or U19123 (N_19123,N_17299,N_16563);
or U19124 (N_19124,N_16596,N_17094);
xor U19125 (N_19125,N_17929,N_16771);
nand U19126 (N_19126,N_17980,N_17065);
nor U19127 (N_19127,N_17839,N_17847);
xor U19128 (N_19128,N_16965,N_17456);
xnor U19129 (N_19129,N_16805,N_17369);
nand U19130 (N_19130,N_17200,N_17007);
and U19131 (N_19131,N_16661,N_17727);
or U19132 (N_19132,N_17329,N_17514);
nand U19133 (N_19133,N_17504,N_16824);
or U19134 (N_19134,N_17973,N_17971);
and U19135 (N_19135,N_16559,N_17340);
or U19136 (N_19136,N_17897,N_17507);
nor U19137 (N_19137,N_17769,N_17166);
and U19138 (N_19138,N_16738,N_17054);
nand U19139 (N_19139,N_17203,N_16895);
nand U19140 (N_19140,N_17811,N_16878);
or U19141 (N_19141,N_16840,N_17515);
nand U19142 (N_19142,N_17752,N_17588);
nand U19143 (N_19143,N_17384,N_16843);
nor U19144 (N_19144,N_17479,N_16500);
nor U19145 (N_19145,N_16519,N_16978);
xnor U19146 (N_19146,N_17492,N_17193);
and U19147 (N_19147,N_17483,N_17554);
or U19148 (N_19148,N_17437,N_16594);
and U19149 (N_19149,N_17301,N_17664);
and U19150 (N_19150,N_17039,N_16971);
nor U19151 (N_19151,N_17239,N_17029);
and U19152 (N_19152,N_17850,N_17562);
xor U19153 (N_19153,N_16587,N_16915);
and U19154 (N_19154,N_17740,N_17260);
nor U19155 (N_19155,N_17349,N_17501);
and U19156 (N_19156,N_17987,N_17095);
and U19157 (N_19157,N_17697,N_16505);
nor U19158 (N_19158,N_16593,N_17815);
or U19159 (N_19159,N_16645,N_16860);
nor U19160 (N_19160,N_17822,N_17496);
xnor U19161 (N_19161,N_17610,N_16860);
and U19162 (N_19162,N_17264,N_17647);
nor U19163 (N_19163,N_17399,N_16918);
and U19164 (N_19164,N_17918,N_17979);
and U19165 (N_19165,N_17879,N_17556);
xnor U19166 (N_19166,N_17868,N_17778);
xnor U19167 (N_19167,N_17454,N_17418);
or U19168 (N_19168,N_17462,N_17838);
nor U19169 (N_19169,N_17597,N_17866);
or U19170 (N_19170,N_17768,N_17056);
or U19171 (N_19171,N_17228,N_16658);
and U19172 (N_19172,N_17309,N_17449);
or U19173 (N_19173,N_16871,N_16901);
nor U19174 (N_19174,N_16948,N_17524);
nor U19175 (N_19175,N_16821,N_17431);
and U19176 (N_19176,N_16920,N_16689);
and U19177 (N_19177,N_17246,N_17302);
and U19178 (N_19178,N_17248,N_16526);
nand U19179 (N_19179,N_17226,N_16873);
nand U19180 (N_19180,N_16541,N_17196);
nor U19181 (N_19181,N_17896,N_17657);
and U19182 (N_19182,N_17557,N_16661);
xnor U19183 (N_19183,N_16923,N_17844);
nor U19184 (N_19184,N_16940,N_17053);
or U19185 (N_19185,N_17458,N_17050);
nand U19186 (N_19186,N_16927,N_17976);
or U19187 (N_19187,N_17662,N_16708);
nor U19188 (N_19188,N_17219,N_17147);
nand U19189 (N_19189,N_17451,N_17810);
and U19190 (N_19190,N_17077,N_16982);
nor U19191 (N_19191,N_17046,N_16670);
or U19192 (N_19192,N_17760,N_16819);
or U19193 (N_19193,N_17670,N_16609);
nand U19194 (N_19194,N_17567,N_17497);
or U19195 (N_19195,N_16581,N_16965);
and U19196 (N_19196,N_17550,N_17645);
nand U19197 (N_19197,N_17905,N_16596);
xnor U19198 (N_19198,N_17447,N_17050);
or U19199 (N_19199,N_17479,N_17439);
or U19200 (N_19200,N_16922,N_17822);
nor U19201 (N_19201,N_17831,N_17546);
nor U19202 (N_19202,N_17602,N_17951);
nor U19203 (N_19203,N_16806,N_17470);
nand U19204 (N_19204,N_16769,N_17359);
and U19205 (N_19205,N_16704,N_17280);
or U19206 (N_19206,N_17274,N_17919);
xor U19207 (N_19207,N_16931,N_16591);
nand U19208 (N_19208,N_16978,N_16959);
xnor U19209 (N_19209,N_17420,N_16943);
and U19210 (N_19210,N_17717,N_16777);
nor U19211 (N_19211,N_16682,N_17099);
nor U19212 (N_19212,N_17204,N_17802);
xor U19213 (N_19213,N_17800,N_16698);
xor U19214 (N_19214,N_17070,N_17799);
nand U19215 (N_19215,N_17966,N_17909);
nor U19216 (N_19216,N_16862,N_17099);
and U19217 (N_19217,N_17811,N_17171);
nor U19218 (N_19218,N_16723,N_17288);
and U19219 (N_19219,N_16598,N_16632);
xnor U19220 (N_19220,N_17189,N_16712);
xor U19221 (N_19221,N_17612,N_17604);
or U19222 (N_19222,N_16847,N_17198);
and U19223 (N_19223,N_16686,N_17829);
xnor U19224 (N_19224,N_16623,N_16553);
nor U19225 (N_19225,N_16776,N_17859);
and U19226 (N_19226,N_17492,N_16800);
and U19227 (N_19227,N_17225,N_16924);
nand U19228 (N_19228,N_17446,N_17359);
and U19229 (N_19229,N_16553,N_17665);
nand U19230 (N_19230,N_16932,N_17422);
nor U19231 (N_19231,N_17781,N_16756);
nand U19232 (N_19232,N_17226,N_16821);
or U19233 (N_19233,N_17402,N_16970);
xor U19234 (N_19234,N_16654,N_17194);
nand U19235 (N_19235,N_17596,N_17220);
xnor U19236 (N_19236,N_17671,N_17282);
or U19237 (N_19237,N_16811,N_17363);
xnor U19238 (N_19238,N_17142,N_17986);
or U19239 (N_19239,N_16614,N_17968);
or U19240 (N_19240,N_16818,N_17093);
nand U19241 (N_19241,N_16610,N_17653);
nand U19242 (N_19242,N_17794,N_17443);
and U19243 (N_19243,N_17363,N_16870);
nor U19244 (N_19244,N_16777,N_16547);
xor U19245 (N_19245,N_17723,N_17423);
nor U19246 (N_19246,N_16745,N_16856);
nand U19247 (N_19247,N_16778,N_17771);
xnor U19248 (N_19248,N_17467,N_16981);
and U19249 (N_19249,N_17411,N_16888);
nand U19250 (N_19250,N_17022,N_17199);
xnor U19251 (N_19251,N_17554,N_16896);
nor U19252 (N_19252,N_16582,N_16962);
xor U19253 (N_19253,N_17918,N_17255);
nand U19254 (N_19254,N_17256,N_17516);
nand U19255 (N_19255,N_17250,N_16749);
and U19256 (N_19256,N_17653,N_17824);
nor U19257 (N_19257,N_17727,N_16786);
nand U19258 (N_19258,N_17287,N_17974);
xor U19259 (N_19259,N_17783,N_17465);
or U19260 (N_19260,N_17655,N_16762);
nand U19261 (N_19261,N_17638,N_17057);
and U19262 (N_19262,N_17593,N_17492);
nand U19263 (N_19263,N_17916,N_16986);
and U19264 (N_19264,N_17701,N_16710);
nor U19265 (N_19265,N_16684,N_17603);
nor U19266 (N_19266,N_16839,N_16592);
nand U19267 (N_19267,N_16721,N_17802);
and U19268 (N_19268,N_17952,N_17880);
and U19269 (N_19269,N_16757,N_17660);
nand U19270 (N_19270,N_17639,N_17068);
or U19271 (N_19271,N_17439,N_17550);
xor U19272 (N_19272,N_16737,N_16873);
xnor U19273 (N_19273,N_17670,N_17281);
xnor U19274 (N_19274,N_16858,N_17452);
or U19275 (N_19275,N_17411,N_16588);
or U19276 (N_19276,N_16591,N_17537);
and U19277 (N_19277,N_17692,N_17902);
nand U19278 (N_19278,N_17443,N_17267);
or U19279 (N_19279,N_17032,N_16856);
and U19280 (N_19280,N_17098,N_17552);
nor U19281 (N_19281,N_17619,N_17916);
and U19282 (N_19282,N_17064,N_17293);
nor U19283 (N_19283,N_16734,N_17290);
nor U19284 (N_19284,N_16825,N_17082);
or U19285 (N_19285,N_17477,N_16804);
nand U19286 (N_19286,N_17335,N_17363);
xnor U19287 (N_19287,N_17733,N_17223);
xor U19288 (N_19288,N_16882,N_16533);
and U19289 (N_19289,N_16541,N_16509);
and U19290 (N_19290,N_17633,N_16504);
nor U19291 (N_19291,N_17693,N_17645);
nor U19292 (N_19292,N_16683,N_17718);
or U19293 (N_19293,N_16871,N_17593);
nand U19294 (N_19294,N_17195,N_17371);
nor U19295 (N_19295,N_17144,N_17948);
and U19296 (N_19296,N_16804,N_17685);
and U19297 (N_19297,N_17163,N_16523);
and U19298 (N_19298,N_17926,N_17106);
or U19299 (N_19299,N_17382,N_17133);
or U19300 (N_19300,N_17474,N_17644);
or U19301 (N_19301,N_16695,N_16739);
nor U19302 (N_19302,N_17107,N_17072);
nor U19303 (N_19303,N_17388,N_17904);
nand U19304 (N_19304,N_17761,N_16963);
or U19305 (N_19305,N_17655,N_17394);
or U19306 (N_19306,N_17231,N_17060);
nand U19307 (N_19307,N_16573,N_17510);
xor U19308 (N_19308,N_17326,N_16634);
xnor U19309 (N_19309,N_16737,N_16756);
xnor U19310 (N_19310,N_16663,N_16824);
or U19311 (N_19311,N_17124,N_17869);
and U19312 (N_19312,N_17963,N_16739);
and U19313 (N_19313,N_17862,N_17277);
xor U19314 (N_19314,N_17334,N_17603);
nand U19315 (N_19315,N_17620,N_17204);
xor U19316 (N_19316,N_16893,N_17664);
nor U19317 (N_19317,N_16823,N_17117);
and U19318 (N_19318,N_16507,N_16915);
or U19319 (N_19319,N_17426,N_17389);
xor U19320 (N_19320,N_17411,N_17147);
nor U19321 (N_19321,N_16984,N_17095);
and U19322 (N_19322,N_16803,N_17283);
xnor U19323 (N_19323,N_16739,N_17368);
nor U19324 (N_19324,N_17826,N_17342);
or U19325 (N_19325,N_16889,N_16980);
and U19326 (N_19326,N_17615,N_17102);
nand U19327 (N_19327,N_17194,N_17945);
or U19328 (N_19328,N_17299,N_17915);
nor U19329 (N_19329,N_17582,N_17258);
nand U19330 (N_19330,N_17649,N_17512);
nand U19331 (N_19331,N_16822,N_16570);
nand U19332 (N_19332,N_16529,N_17909);
or U19333 (N_19333,N_16738,N_17531);
nand U19334 (N_19334,N_17394,N_16884);
and U19335 (N_19335,N_16738,N_16892);
nor U19336 (N_19336,N_16743,N_16756);
nor U19337 (N_19337,N_16914,N_17216);
and U19338 (N_19338,N_16734,N_16719);
and U19339 (N_19339,N_17551,N_17241);
nor U19340 (N_19340,N_17855,N_17205);
xnor U19341 (N_19341,N_17769,N_17329);
nand U19342 (N_19342,N_17396,N_17303);
and U19343 (N_19343,N_16749,N_17953);
nor U19344 (N_19344,N_17378,N_16756);
xor U19345 (N_19345,N_16906,N_17322);
nand U19346 (N_19346,N_17611,N_17029);
nor U19347 (N_19347,N_16881,N_17868);
nand U19348 (N_19348,N_17451,N_16858);
xnor U19349 (N_19349,N_17448,N_17210);
nand U19350 (N_19350,N_17322,N_17169);
or U19351 (N_19351,N_16507,N_17264);
and U19352 (N_19352,N_16751,N_17318);
xnor U19353 (N_19353,N_17969,N_17959);
nand U19354 (N_19354,N_17639,N_17954);
nor U19355 (N_19355,N_16924,N_16710);
or U19356 (N_19356,N_17390,N_16770);
and U19357 (N_19357,N_17191,N_16621);
nor U19358 (N_19358,N_17054,N_16979);
xor U19359 (N_19359,N_17829,N_16645);
and U19360 (N_19360,N_17569,N_17565);
nand U19361 (N_19361,N_16881,N_17009);
nand U19362 (N_19362,N_17597,N_17509);
xor U19363 (N_19363,N_17699,N_17886);
nand U19364 (N_19364,N_16585,N_17574);
or U19365 (N_19365,N_16618,N_17034);
nand U19366 (N_19366,N_17312,N_17904);
or U19367 (N_19367,N_16816,N_17459);
xor U19368 (N_19368,N_17915,N_17160);
or U19369 (N_19369,N_17696,N_17031);
xnor U19370 (N_19370,N_17991,N_16972);
xor U19371 (N_19371,N_17559,N_16993);
and U19372 (N_19372,N_16749,N_17672);
nand U19373 (N_19373,N_17731,N_17609);
or U19374 (N_19374,N_16598,N_17371);
nand U19375 (N_19375,N_17494,N_17253);
or U19376 (N_19376,N_17623,N_17212);
or U19377 (N_19377,N_16945,N_17234);
nor U19378 (N_19378,N_16903,N_17218);
nand U19379 (N_19379,N_17957,N_17426);
nand U19380 (N_19380,N_16742,N_17747);
and U19381 (N_19381,N_16639,N_17365);
nand U19382 (N_19382,N_16554,N_16649);
or U19383 (N_19383,N_16901,N_17464);
or U19384 (N_19384,N_17527,N_17553);
nand U19385 (N_19385,N_17856,N_17034);
or U19386 (N_19386,N_17872,N_16705);
or U19387 (N_19387,N_17670,N_16584);
nor U19388 (N_19388,N_16590,N_17845);
nand U19389 (N_19389,N_16859,N_16930);
and U19390 (N_19390,N_16917,N_17867);
nor U19391 (N_19391,N_16658,N_17522);
nand U19392 (N_19392,N_17292,N_16754);
or U19393 (N_19393,N_17097,N_16807);
nand U19394 (N_19394,N_16645,N_17087);
xnor U19395 (N_19395,N_16579,N_16717);
and U19396 (N_19396,N_17954,N_17078);
nand U19397 (N_19397,N_16799,N_16820);
nor U19398 (N_19398,N_16541,N_16876);
nand U19399 (N_19399,N_17104,N_16972);
and U19400 (N_19400,N_16819,N_16522);
xor U19401 (N_19401,N_17880,N_17679);
nand U19402 (N_19402,N_17179,N_16523);
and U19403 (N_19403,N_17669,N_17155);
nor U19404 (N_19404,N_17745,N_17657);
or U19405 (N_19405,N_16785,N_16548);
nor U19406 (N_19406,N_17569,N_17689);
nor U19407 (N_19407,N_17542,N_16714);
nor U19408 (N_19408,N_16817,N_17426);
and U19409 (N_19409,N_17808,N_17231);
xnor U19410 (N_19410,N_17349,N_16921);
and U19411 (N_19411,N_16883,N_16636);
xor U19412 (N_19412,N_17336,N_16543);
and U19413 (N_19413,N_17617,N_17212);
xor U19414 (N_19414,N_17328,N_16889);
xor U19415 (N_19415,N_17549,N_17477);
nor U19416 (N_19416,N_17124,N_16702);
nor U19417 (N_19417,N_17334,N_17796);
nor U19418 (N_19418,N_17963,N_17906);
nor U19419 (N_19419,N_17293,N_16675);
xnor U19420 (N_19420,N_17953,N_17135);
nand U19421 (N_19421,N_16579,N_17831);
nor U19422 (N_19422,N_17738,N_17126);
and U19423 (N_19423,N_17837,N_17619);
or U19424 (N_19424,N_17437,N_17149);
or U19425 (N_19425,N_17664,N_17090);
or U19426 (N_19426,N_16867,N_16985);
nor U19427 (N_19427,N_16789,N_17195);
nor U19428 (N_19428,N_17754,N_17675);
xor U19429 (N_19429,N_17458,N_17492);
and U19430 (N_19430,N_17724,N_17122);
or U19431 (N_19431,N_16524,N_16696);
nand U19432 (N_19432,N_17846,N_16867);
nand U19433 (N_19433,N_17569,N_16677);
nand U19434 (N_19434,N_17202,N_17705);
nand U19435 (N_19435,N_17685,N_16673);
or U19436 (N_19436,N_17745,N_17452);
or U19437 (N_19437,N_17341,N_16865);
nand U19438 (N_19438,N_17501,N_16893);
and U19439 (N_19439,N_16687,N_17033);
xor U19440 (N_19440,N_17845,N_17492);
nor U19441 (N_19441,N_17242,N_17401);
xnor U19442 (N_19442,N_16877,N_16724);
xnor U19443 (N_19443,N_17999,N_17712);
nor U19444 (N_19444,N_17299,N_17429);
nand U19445 (N_19445,N_16824,N_16819);
and U19446 (N_19446,N_17050,N_17585);
or U19447 (N_19447,N_17267,N_17311);
nand U19448 (N_19448,N_17619,N_16579);
or U19449 (N_19449,N_16656,N_17753);
nand U19450 (N_19450,N_17142,N_17433);
nand U19451 (N_19451,N_17300,N_16532);
xnor U19452 (N_19452,N_16932,N_17419);
xor U19453 (N_19453,N_17982,N_17927);
xnor U19454 (N_19454,N_17366,N_17871);
nand U19455 (N_19455,N_17490,N_17956);
nor U19456 (N_19456,N_17556,N_16884);
or U19457 (N_19457,N_17731,N_16589);
and U19458 (N_19458,N_17986,N_17163);
nand U19459 (N_19459,N_16660,N_17572);
nand U19460 (N_19460,N_16694,N_17383);
and U19461 (N_19461,N_16966,N_17979);
or U19462 (N_19462,N_17123,N_17032);
xnor U19463 (N_19463,N_16702,N_17902);
or U19464 (N_19464,N_16507,N_16953);
xor U19465 (N_19465,N_16958,N_17208);
and U19466 (N_19466,N_16736,N_17902);
nand U19467 (N_19467,N_17250,N_16922);
nand U19468 (N_19468,N_16814,N_17590);
and U19469 (N_19469,N_16999,N_17243);
xor U19470 (N_19470,N_16899,N_17793);
xnor U19471 (N_19471,N_17261,N_17814);
nand U19472 (N_19472,N_17833,N_17395);
or U19473 (N_19473,N_17609,N_17161);
xnor U19474 (N_19474,N_17250,N_17080);
or U19475 (N_19475,N_17520,N_17532);
and U19476 (N_19476,N_17707,N_17853);
nand U19477 (N_19477,N_16588,N_17976);
or U19478 (N_19478,N_17590,N_17930);
or U19479 (N_19479,N_17054,N_17921);
nand U19480 (N_19480,N_17073,N_17580);
nand U19481 (N_19481,N_16986,N_16853);
and U19482 (N_19482,N_16909,N_17882);
xnor U19483 (N_19483,N_16619,N_17151);
nand U19484 (N_19484,N_17115,N_17427);
nand U19485 (N_19485,N_17410,N_17723);
nand U19486 (N_19486,N_16952,N_17294);
nor U19487 (N_19487,N_16535,N_16829);
xor U19488 (N_19488,N_16925,N_16622);
nor U19489 (N_19489,N_17361,N_17184);
or U19490 (N_19490,N_16800,N_17140);
nand U19491 (N_19491,N_17251,N_17864);
xor U19492 (N_19492,N_16972,N_16878);
xor U19493 (N_19493,N_16928,N_17098);
or U19494 (N_19494,N_17217,N_16774);
nor U19495 (N_19495,N_16679,N_17918);
nand U19496 (N_19496,N_17867,N_17677);
xnor U19497 (N_19497,N_17786,N_17013);
nand U19498 (N_19498,N_17706,N_17423);
nand U19499 (N_19499,N_16724,N_16676);
and U19500 (N_19500,N_19484,N_18033);
and U19501 (N_19501,N_18329,N_18762);
xnor U19502 (N_19502,N_18618,N_18357);
nor U19503 (N_19503,N_18967,N_18547);
or U19504 (N_19504,N_18541,N_18933);
nor U19505 (N_19505,N_18778,N_18442);
and U19506 (N_19506,N_18632,N_18270);
or U19507 (N_19507,N_18435,N_19055);
nor U19508 (N_19508,N_18663,N_18101);
xnor U19509 (N_19509,N_19033,N_18828);
xnor U19510 (N_19510,N_19043,N_18091);
and U19511 (N_19511,N_18893,N_18903);
nor U19512 (N_19512,N_18815,N_18816);
xnor U19513 (N_19513,N_18793,N_18196);
or U19514 (N_19514,N_19105,N_18365);
nor U19515 (N_19515,N_18086,N_18892);
or U19516 (N_19516,N_18684,N_19236);
xnor U19517 (N_19517,N_19145,N_18532);
nor U19518 (N_19518,N_18886,N_18368);
and U19519 (N_19519,N_19310,N_18773);
nor U19520 (N_19520,N_18508,N_18078);
nor U19521 (N_19521,N_18163,N_19030);
or U19522 (N_19522,N_18154,N_19262);
nand U19523 (N_19523,N_18550,N_18012);
and U19524 (N_19524,N_19406,N_18022);
nor U19525 (N_19525,N_18428,N_19231);
nor U19526 (N_19526,N_18512,N_19106);
xnor U19527 (N_19527,N_18617,N_18981);
and U19528 (N_19528,N_19127,N_19048);
or U19529 (N_19529,N_18352,N_18305);
and U19530 (N_19530,N_18569,N_19166);
xnor U19531 (N_19531,N_19379,N_18956);
nand U19532 (N_19532,N_19342,N_18349);
or U19533 (N_19533,N_19355,N_18955);
nor U19534 (N_19534,N_19478,N_18462);
nor U19535 (N_19535,N_18283,N_19025);
nand U19536 (N_19536,N_18314,N_19137);
nor U19537 (N_19537,N_18176,N_19164);
and U19538 (N_19538,N_18958,N_18876);
nor U19539 (N_19539,N_19135,N_18579);
nand U19540 (N_19540,N_18273,N_19283);
xnor U19541 (N_19541,N_19375,N_19093);
nand U19542 (N_19542,N_18069,N_18571);
xnor U19543 (N_19543,N_19394,N_18709);
nor U19544 (N_19544,N_18346,N_19068);
and U19545 (N_19545,N_19157,N_18714);
nand U19546 (N_19546,N_19083,N_18953);
xnor U19547 (N_19547,N_18850,N_18043);
nand U19548 (N_19548,N_19273,N_18340);
xor U19549 (N_19549,N_19405,N_18947);
nor U19550 (N_19550,N_19334,N_18244);
or U19551 (N_19551,N_19423,N_19208);
or U19552 (N_19552,N_18467,N_18590);
nor U19553 (N_19553,N_18831,N_18100);
or U19554 (N_19554,N_19018,N_19466);
or U19555 (N_19555,N_18738,N_19100);
and U19556 (N_19556,N_18463,N_19403);
and U19557 (N_19557,N_18434,N_18611);
nand U19558 (N_19558,N_19380,N_18990);
xnor U19559 (N_19559,N_18194,N_18080);
and U19560 (N_19560,N_18320,N_18070);
and U19561 (N_19561,N_19343,N_18897);
and U19562 (N_19562,N_18806,N_18603);
and U19563 (N_19563,N_18654,N_18792);
nand U19564 (N_19564,N_18392,N_18090);
nand U19565 (N_19565,N_18197,N_19427);
and U19566 (N_19566,N_18874,N_19097);
xnor U19567 (N_19567,N_18891,N_18476);
xnor U19568 (N_19568,N_18740,N_19229);
or U19569 (N_19569,N_18339,N_19170);
and U19570 (N_19570,N_18545,N_18992);
xnor U19571 (N_19571,N_19404,N_18253);
and U19572 (N_19572,N_18810,N_18011);
nor U19573 (N_19573,N_19429,N_19425);
and U19574 (N_19574,N_18307,N_18420);
nand U19575 (N_19575,N_18358,N_19369);
or U19576 (N_19576,N_18516,N_18864);
nand U19577 (N_19577,N_19315,N_18664);
or U19578 (N_19578,N_19333,N_18628);
or U19579 (N_19579,N_18289,N_18426);
or U19580 (N_19580,N_18267,N_19435);
xor U19581 (N_19581,N_18539,N_18821);
or U19582 (N_19582,N_19089,N_18345);
nand U19583 (N_19583,N_19250,N_18199);
or U19584 (N_19584,N_18556,N_18524);
xnor U19585 (N_19585,N_19475,N_18797);
or U19586 (N_19586,N_19426,N_18491);
and U19587 (N_19587,N_19268,N_18877);
or U19588 (N_19588,N_18366,N_18728);
nand U19589 (N_19589,N_19209,N_18148);
or U19590 (N_19590,N_19196,N_19226);
and U19591 (N_19591,N_18093,N_19330);
and U19592 (N_19592,N_18631,N_18483);
xor U19593 (N_19593,N_18334,N_19362);
and U19594 (N_19594,N_18814,N_19143);
nor U19595 (N_19595,N_19275,N_19265);
xnor U19596 (N_19596,N_18919,N_18837);
xnor U19597 (N_19597,N_18888,N_18730);
nand U19598 (N_19598,N_18984,N_18771);
xor U19599 (N_19599,N_18700,N_19180);
or U19600 (N_19600,N_18985,N_19282);
nor U19601 (N_19601,N_18901,N_19156);
nor U19602 (N_19602,N_18690,N_19059);
nor U19603 (N_19603,N_18131,N_18688);
nand U19604 (N_19604,N_18326,N_18776);
and U19605 (N_19605,N_18162,N_19297);
nor U19606 (N_19606,N_18455,N_18324);
and U19607 (N_19607,N_18068,N_19247);
nand U19608 (N_19608,N_19324,N_18586);
xor U19609 (N_19609,N_18694,N_18546);
nor U19610 (N_19610,N_18059,N_18920);
and U19611 (N_19611,N_19378,N_18923);
xnor U19612 (N_19612,N_19173,N_18446);
xor U19613 (N_19613,N_18717,N_18959);
and U19614 (N_19614,N_18585,N_19306);
or U19615 (N_19615,N_18486,N_19281);
and U19616 (N_19616,N_18904,N_19351);
nor U19617 (N_19617,N_18336,N_18280);
nand U19618 (N_19618,N_19266,N_19431);
xnor U19619 (N_19619,N_19468,N_18139);
nand U19620 (N_19620,N_19108,N_19128);
xnor U19621 (N_19621,N_18045,N_19136);
nor U19622 (N_19622,N_18950,N_18029);
nor U19623 (N_19623,N_19348,N_18480);
xor U19624 (N_19624,N_18034,N_19201);
or U19625 (N_19625,N_18800,N_18871);
nor U19626 (N_19626,N_18582,N_19304);
xor U19627 (N_19627,N_19194,N_18922);
nand U19628 (N_19628,N_18023,N_18658);
and U19629 (N_19629,N_18386,N_18974);
xnor U19630 (N_19630,N_18272,N_18848);
xnor U19631 (N_19631,N_19412,N_18859);
xnor U19632 (N_19632,N_19473,N_18318);
xor U19633 (N_19633,N_18393,N_18453);
xor U19634 (N_19634,N_18062,N_18666);
nor U19635 (N_19635,N_18794,N_18211);
and U19636 (N_19636,N_18936,N_18121);
nand U19637 (N_19637,N_18064,N_18879);
or U19638 (N_19638,N_18406,N_18661);
nor U19639 (N_19639,N_18998,N_19460);
and U19640 (N_19640,N_18543,N_19174);
nand U19641 (N_19641,N_18482,N_19420);
xor U19642 (N_19642,N_18777,N_18041);
nand U19643 (N_19643,N_18566,N_19121);
and U19644 (N_19644,N_18402,N_19045);
nor U19645 (N_19645,N_19418,N_18494);
nor U19646 (N_19646,N_19274,N_18911);
and U19647 (N_19647,N_18843,N_19260);
xnor U19648 (N_19648,N_18264,N_18248);
xor U19649 (N_19649,N_19177,N_18328);
and U19650 (N_19650,N_19487,N_18535);
nand U19651 (N_19651,N_19467,N_19214);
nand U19652 (N_19652,N_18790,N_18077);
xnor U19653 (N_19653,N_18916,N_18284);
xnor U19654 (N_19654,N_18994,N_19248);
xnor U19655 (N_19655,N_19091,N_18622);
and U19656 (N_19656,N_18454,N_18503);
nor U19657 (N_19657,N_19027,N_18942);
or U19658 (N_19658,N_18220,N_18655);
xnor U19659 (N_19659,N_18088,N_18887);
nand U19660 (N_19660,N_18819,N_18997);
nand U19661 (N_19661,N_18878,N_19211);
or U19662 (N_19662,N_18063,N_18254);
nor U19663 (N_19663,N_19354,N_18867);
nand U19664 (N_19664,N_18593,N_18475);
xor U19665 (N_19665,N_18000,N_18360);
and U19666 (N_19666,N_18051,N_18559);
xnor U19667 (N_19667,N_18962,N_19175);
or U19668 (N_19668,N_19116,N_18146);
or U19669 (N_19669,N_18609,N_18301);
nand U19670 (N_19670,N_18114,N_18854);
and U19671 (N_19671,N_18321,N_18239);
or U19672 (N_19672,N_18975,N_19325);
and U19673 (N_19673,N_18676,N_19279);
or U19674 (N_19674,N_18281,N_18941);
xor U19675 (N_19675,N_18432,N_18497);
nand U19676 (N_19676,N_18753,N_18509);
nor U19677 (N_19677,N_19452,N_19336);
nor U19678 (N_19678,N_18662,N_19181);
and U19679 (N_19679,N_18247,N_18869);
xor U19680 (N_19680,N_18583,N_18926);
and U19681 (N_19681,N_18642,N_18506);
and U19682 (N_19682,N_19125,N_19437);
nand U19683 (N_19683,N_18161,N_19316);
nor U19684 (N_19684,N_18774,N_18637);
or U19685 (N_19685,N_19090,N_18173);
or U19686 (N_19686,N_19439,N_18372);
xor U19687 (N_19687,N_19399,N_18474);
xor U19688 (N_19688,N_18287,N_18822);
nor U19689 (N_19689,N_18423,N_19360);
nand U19690 (N_19690,N_19232,N_18180);
or U19691 (N_19691,N_18110,N_18748);
xor U19692 (N_19692,N_18803,N_19398);
xnor U19693 (N_19693,N_19036,N_18779);
nor U19694 (N_19694,N_18531,N_18987);
nand U19695 (N_19695,N_18518,N_18747);
nor U19696 (N_19696,N_18206,N_18589);
and U19697 (N_19697,N_18844,N_19227);
nand U19698 (N_19698,N_18501,N_18931);
nand U19699 (N_19699,N_18652,N_18175);
xor U19700 (N_19700,N_18373,N_18081);
nor U19701 (N_19701,N_18572,N_18650);
and U19702 (N_19702,N_18374,N_19142);
nand U19703 (N_19703,N_19115,N_19332);
and U19704 (N_19704,N_18613,N_18028);
nor U19705 (N_19705,N_18145,N_19359);
nand U19706 (N_19706,N_19044,N_18278);
nand U19707 (N_19707,N_19086,N_19396);
or U19708 (N_19708,N_18095,N_18102);
or U19709 (N_19709,N_18332,N_18404);
xor U19710 (N_19710,N_18370,N_18945);
xnor U19711 (N_19711,N_19470,N_19414);
and U19712 (N_19712,N_18979,N_19041);
nor U19713 (N_19713,N_18355,N_18193);
or U19714 (N_19714,N_18898,N_18251);
nor U19715 (N_19715,N_18493,N_19222);
nand U19716 (N_19716,N_18460,N_18066);
nand U19717 (N_19717,N_19184,N_18087);
nand U19718 (N_19718,N_18948,N_18939);
nand U19719 (N_19719,N_18192,N_18761);
xnor U19720 (N_19720,N_18016,N_18515);
and U19721 (N_19721,N_18563,N_18565);
nand U19722 (N_19722,N_18678,N_19293);
nor U19723 (N_19723,N_19016,N_18217);
nor U19724 (N_19724,N_19462,N_18243);
nor U19725 (N_19725,N_18096,N_18050);
nor U19726 (N_19726,N_18699,N_18723);
xnor U19727 (N_19727,N_18380,N_19186);
nor U19728 (N_19728,N_19472,N_18834);
nand U19729 (N_19729,N_18001,N_18057);
nand U19730 (N_19730,N_19482,N_19474);
xor U19731 (N_19731,N_19497,N_18513);
or U19732 (N_19732,N_19493,N_18549);
and U19733 (N_19733,N_19317,N_18147);
xnor U19734 (N_19734,N_18238,N_19070);
xor U19735 (N_19735,N_18913,N_19308);
nor U19736 (N_19736,N_19329,N_19067);
nor U19737 (N_19737,N_18444,N_18484);
nand U19738 (N_19738,N_18781,N_18303);
or U19739 (N_19739,N_19147,N_18179);
nand U19740 (N_19740,N_18689,N_19081);
and U19741 (N_19741,N_19216,N_18884);
xnor U19742 (N_19742,N_19331,N_19239);
xor U19743 (N_19743,N_18245,N_18604);
nor U19744 (N_19744,N_18969,N_19276);
and U19745 (N_19745,N_19202,N_19010);
xor U19746 (N_19746,N_19243,N_18588);
nand U19747 (N_19747,N_18805,N_18205);
and U19748 (N_19748,N_18561,N_19490);
nor U19749 (N_19749,N_18846,N_18259);
or U19750 (N_19750,N_18276,N_19213);
nand U19751 (N_19751,N_18500,N_18744);
or U19752 (N_19752,N_18249,N_19047);
nand U19753 (N_19753,N_19134,N_18938);
xnor U19754 (N_19754,N_19159,N_18852);
xnor U19755 (N_19755,N_18924,N_18782);
or U19756 (N_19756,N_18692,N_18711);
xor U19757 (N_19757,N_18918,N_19032);
and U19758 (N_19758,N_19168,N_19294);
and U19759 (N_19759,N_18930,N_18377);
xor U19760 (N_19760,N_18416,N_19154);
xor U19761 (N_19761,N_19060,N_19352);
nand U19762 (N_19762,N_18350,N_18388);
nand U19763 (N_19763,N_19272,N_18004);
or U19764 (N_19764,N_18808,N_18167);
nand U19765 (N_19765,N_19075,N_18469);
or U19766 (N_19766,N_19280,N_18129);
xor U19767 (N_19767,N_19225,N_19193);
nor U19768 (N_19768,N_18542,N_18659);
xor U19769 (N_19769,N_18555,N_18651);
and U19770 (N_19770,N_18448,N_18046);
or U19771 (N_19771,N_19483,N_19249);
or U19772 (N_19772,N_18452,N_19320);
or U19773 (N_19773,N_19263,N_18682);
nor U19774 (N_19774,N_18492,N_19046);
nor U19775 (N_19775,N_19099,N_18246);
nor U19776 (N_19776,N_19062,N_18390);
and U19777 (N_19777,N_18451,N_19498);
and U19778 (N_19778,N_18643,N_19295);
xor U19779 (N_19779,N_18725,N_19189);
nor U19780 (N_19780,N_19411,N_19071);
nor U19781 (N_19781,N_18823,N_18519);
nand U19782 (N_19782,N_18534,N_19117);
nor U19783 (N_19783,N_18255,N_18413);
and U19784 (N_19784,N_18319,N_18219);
nand U19785 (N_19785,N_19087,N_18645);
nor U19786 (N_19786,N_18602,N_18548);
and U19787 (N_19787,N_19450,N_18980);
or U19788 (N_19788,N_18520,N_18098);
xnor U19789 (N_19789,N_19040,N_18302);
and U19790 (N_19790,N_18032,N_19428);
or U19791 (N_19791,N_18252,N_18209);
xor U19792 (N_19792,N_19064,N_18616);
or U19793 (N_19793,N_18839,N_19284);
and U19794 (N_19794,N_18256,N_18149);
or U19795 (N_19795,N_18499,N_18921);
and U19796 (N_19796,N_19422,N_18218);
xnor U19797 (N_19797,N_18424,N_18934);
nand U19798 (N_19798,N_18530,N_18067);
nor U19799 (N_19799,N_18596,N_18989);
xor U19800 (N_19800,N_18890,N_18450);
xor U19801 (N_19801,N_18932,N_18759);
or U19802 (N_19802,N_19499,N_18758);
xnor U19803 (N_19803,N_18809,N_19095);
or U19804 (N_19804,N_19447,N_18140);
nand U19805 (N_19805,N_18840,N_18168);
xor U19806 (N_19806,N_18250,N_19442);
nor U19807 (N_19807,N_18234,N_19084);
and U19808 (N_19808,N_19053,N_19436);
nor U19809 (N_19809,N_18159,N_18660);
nand U19810 (N_19810,N_19148,N_18310);
nand U19811 (N_19811,N_19311,N_18872);
or U19812 (N_19812,N_19357,N_18418);
xor U19813 (N_19813,N_19344,N_18943);
nand U19814 (N_19814,N_19102,N_19008);
and U19815 (N_19815,N_18718,N_18181);
nor U19816 (N_19816,N_18038,N_18915);
nor U19817 (N_19817,N_18798,N_18174);
xor U19818 (N_19818,N_18914,N_19123);
and U19819 (N_19819,N_18082,N_18210);
or U19820 (N_19820,N_18802,N_18860);
nand U19821 (N_19821,N_19491,N_18641);
xnor U19822 (N_19822,N_19037,N_18060);
xor U19823 (N_19823,N_19277,N_18010);
nor U19824 (N_19824,N_19119,N_18459);
nor U19825 (N_19825,N_18624,N_18019);
and U19826 (N_19826,N_18780,N_18130);
and U19827 (N_19827,N_18061,N_18395);
xor U19828 (N_19828,N_18657,N_18269);
and U19829 (N_19829,N_19035,N_19014);
nor U19830 (N_19830,N_19223,N_19113);
or U19831 (N_19831,N_19171,N_18623);
xnor U19832 (N_19832,N_18615,N_19353);
nand U19833 (N_19833,N_18411,N_19361);
nand U19834 (N_19834,N_18853,N_18526);
nand U19835 (N_19835,N_18675,N_19217);
nor U19836 (N_19836,N_18737,N_19419);
nor U19837 (N_19837,N_19221,N_19421);
or U19838 (N_19838,N_19078,N_18732);
or U19839 (N_19839,N_19079,N_18529);
nand U19840 (N_19840,N_18036,N_19118);
nor U19841 (N_19841,N_19395,N_19058);
nor U19842 (N_19842,N_19479,N_18083);
nor U19843 (N_19843,N_18568,N_18905);
and U19844 (N_19844,N_19219,N_18387);
xor U19845 (N_19845,N_18580,N_18035);
nand U19846 (N_19846,N_18191,N_18736);
nand U19847 (N_19847,N_19074,N_18594);
or U19848 (N_19848,N_18075,N_19096);
nand U19849 (N_19849,N_18713,N_19402);
and U19850 (N_19850,N_19288,N_18620);
and U19851 (N_19851,N_18553,N_18047);
nor U19852 (N_19852,N_19237,N_19434);
and U19853 (N_19853,N_18973,N_18382);
nand U19854 (N_19854,N_18300,N_18863);
nand U19855 (N_19855,N_18907,N_19131);
or U19856 (N_19856,N_18039,N_18788);
or U19857 (N_19857,N_18412,N_18785);
nor U19858 (N_19858,N_19443,N_18207);
nor U19859 (N_19859,N_18222,N_18313);
xnor U19860 (N_19860,N_18695,N_18026);
nor U19861 (N_19861,N_18295,N_18221);
nor U19862 (N_19862,N_18674,N_19269);
xor U19863 (N_19863,N_18203,N_18008);
nand U19864 (N_19864,N_18710,N_19372);
nand U19865 (N_19865,N_18361,N_19261);
or U19866 (N_19866,N_18749,N_19176);
nor U19867 (N_19867,N_19165,N_19347);
nor U19868 (N_19868,N_18719,N_18708);
xnor U19869 (N_19869,N_18362,N_18304);
and U19870 (N_19870,N_19069,N_18707);
nor U19871 (N_19871,N_18824,N_18436);
and U19872 (N_19872,N_18697,N_18232);
and U19873 (N_19873,N_19291,N_18461);
nor U19874 (N_19874,N_19230,N_18917);
nand U19875 (N_19875,N_18044,N_18605);
or U19876 (N_19876,N_18621,N_18136);
nand U19877 (N_19877,N_18909,N_18118);
or U19878 (N_19878,N_18775,N_18649);
nor U19879 (N_19879,N_18286,N_18669);
nand U19880 (N_19880,N_19377,N_19464);
and U19881 (N_19881,N_18410,N_18795);
or U19882 (N_19882,N_18341,N_19101);
and U19883 (N_19883,N_18257,N_19477);
nand U19884 (N_19884,N_18160,N_18094);
nand U19885 (N_19885,N_18384,N_19407);
and U19886 (N_19886,N_18165,N_18517);
and U19887 (N_19887,N_19271,N_18972);
xor U19888 (N_19888,N_18408,N_18433);
nor U19889 (N_19889,N_19022,N_19188);
xor U19890 (N_19890,N_19433,N_19386);
and U19891 (N_19891,N_18299,N_18223);
and U19892 (N_19892,N_18477,N_18940);
nor U19893 (N_19893,N_18521,N_18268);
nand U19894 (N_19894,N_18472,N_18048);
nand U19895 (N_19895,N_18971,N_18626);
or U19896 (N_19896,N_19387,N_18963);
xor U19897 (N_19897,N_19393,N_18108);
nor U19898 (N_19898,N_19356,N_18085);
nand U19899 (N_19899,N_18449,N_19312);
and U19900 (N_19900,N_18567,N_18498);
or U19901 (N_19901,N_18113,N_19107);
or U19902 (N_19902,N_18369,N_19251);
and U19903 (N_19903,N_18703,N_18007);
xor U19904 (N_19904,N_18441,N_18236);
xor U19905 (N_19905,N_19061,N_18644);
nor U19906 (N_19906,N_18241,N_19258);
or U19907 (N_19907,N_18097,N_18906);
or U19908 (N_19908,N_18421,N_18755);
and U19909 (N_19909,N_18478,N_19339);
nand U19910 (N_19910,N_18528,N_19178);
nor U19911 (N_19911,N_18342,N_19314);
or U19912 (N_19912,N_18564,N_19163);
nor U19913 (N_19913,N_18949,N_19072);
nor U19914 (N_19914,N_18182,N_19082);
xnor U19915 (N_19915,N_18151,N_18638);
xnor U19916 (N_19916,N_18055,N_18152);
nand U19917 (N_19917,N_19388,N_18505);
nor U19918 (N_19918,N_18306,N_19124);
xnor U19919 (N_19919,N_19459,N_19409);
nand U19920 (N_19920,N_18665,N_18999);
xor U19921 (N_19921,N_19120,N_19203);
nand U19922 (N_19922,N_19323,N_18419);
and U19923 (N_19923,N_18851,N_19368);
xnor U19924 (N_19924,N_18458,N_19210);
or U19925 (N_19925,N_18673,N_19007);
and U19926 (N_19926,N_18685,N_18470);
nand U19927 (N_19927,N_18827,N_19256);
and U19928 (N_19928,N_19149,N_19088);
nand U19929 (N_19929,N_19384,N_18002);
nand U19930 (N_19930,N_19065,N_19289);
nor U19931 (N_19931,N_19192,N_18347);
nand U19932 (N_19932,N_18807,N_18544);
and U19933 (N_19933,N_18186,N_18504);
nand U19934 (N_19934,N_18190,N_19004);
xor U19935 (N_19935,N_19257,N_18353);
xnor U19936 (N_19936,N_18954,N_18899);
xnor U19937 (N_19937,N_19471,N_18635);
or U19938 (N_19938,N_19092,N_19307);
nand U19939 (N_19939,N_18811,N_18201);
xor U19940 (N_19940,N_18224,N_19441);
nand U19941 (N_19941,N_18601,N_19296);
and U19942 (N_19942,N_18274,N_18275);
nand U19943 (N_19943,N_18414,N_19410);
or U19944 (N_19944,N_18634,N_19207);
or U19945 (N_19945,N_18204,N_19397);
or U19946 (N_19946,N_18171,N_18523);
nand U19947 (N_19947,N_19321,N_18229);
nor U19948 (N_19948,N_19322,N_19050);
nand U19949 (N_19949,N_18178,N_18003);
nand U19950 (N_19950,N_18693,N_19455);
or U19951 (N_19951,N_18522,N_18716);
nand U19952 (N_19952,N_19114,N_18263);
or U19953 (N_19953,N_18351,N_18595);
nor U19954 (N_19954,N_18715,N_18344);
nand U19955 (N_19955,N_18683,N_18630);
or U19956 (N_19956,N_18213,N_18801);
or U19957 (N_19957,N_19158,N_18466);
nor U19958 (N_19958,N_18396,N_18399);
nor U19959 (N_19959,N_18538,N_18479);
and U19960 (N_19960,N_18786,N_18142);
nand U19961 (N_19961,N_18376,N_18488);
or U19962 (N_19962,N_18597,N_19302);
or U19963 (N_19963,N_19300,N_18896);
xor U19964 (N_19964,N_18970,N_18183);
or U19965 (N_19965,N_18902,N_19346);
nor U19966 (N_19966,N_19140,N_18883);
nor U19967 (N_19967,N_18293,N_18966);
xnor U19968 (N_19968,N_18875,N_19246);
or U19969 (N_19969,N_19029,N_18185);
and U19970 (N_19970,N_19382,N_18394);
or U19971 (N_19971,N_18951,N_19005);
nor U19972 (N_19972,N_18783,N_18670);
and U19973 (N_19973,N_18712,N_18187);
xnor U19974 (N_19974,N_18405,N_18079);
and U19975 (N_19975,N_19039,N_18726);
nand U19976 (N_19976,N_18215,N_18681);
nor U19977 (N_19977,N_18415,N_18667);
and U19978 (N_19978,N_19021,N_18849);
nor U19979 (N_19979,N_19456,N_18364);
xor U19980 (N_19980,N_18978,N_18440);
nand U19981 (N_19981,N_18671,N_18889);
xor U19982 (N_19982,N_19287,N_18056);
or U19983 (N_19983,N_18608,N_19153);
or U19984 (N_19984,N_19011,N_18053);
nor U19985 (N_19985,N_18610,N_19486);
and U19986 (N_19986,N_18125,N_19109);
xor U19987 (N_19987,N_19430,N_18552);
nand U19988 (N_19988,N_18495,N_18993);
nand U19989 (N_19989,N_18338,N_18705);
xor U19990 (N_19990,N_19345,N_18836);
and U19991 (N_19991,N_18071,N_19370);
nor U19992 (N_19992,N_18076,N_19390);
or U19993 (N_19993,N_18262,N_18578);
and U19994 (N_19994,N_18024,N_18829);
nand U19995 (N_19995,N_19286,N_19367);
or U19996 (N_19996,N_18225,N_18865);
or U19997 (N_19997,N_18741,N_18323);
nor U19998 (N_19998,N_18111,N_18636);
or U19999 (N_19999,N_18367,N_18633);
xor U20000 (N_20000,N_18763,N_18908);
xnor U20001 (N_20001,N_18170,N_19408);
or U20002 (N_20002,N_18156,N_19066);
xor U20003 (N_20003,N_18957,N_18983);
nor U20004 (N_20004,N_18018,N_19241);
or U20005 (N_20005,N_18430,N_18084);
nor U20006 (N_20006,N_19416,N_18912);
nand U20007 (N_20007,N_18237,N_18507);
nand U20008 (N_20008,N_18866,N_18261);
or U20009 (N_20009,N_19042,N_19438);
xnor U20010 (N_20010,N_18481,N_18540);
nor U20011 (N_20011,N_18724,N_18935);
nand U20012 (N_20012,N_19152,N_19358);
nand U20013 (N_20013,N_19126,N_18857);
xnor U20014 (N_20014,N_19328,N_19376);
and U20015 (N_20015,N_19495,N_19112);
nand U20016 (N_20016,N_19244,N_19389);
and U20017 (N_20017,N_18398,N_19363);
or U20018 (N_20018,N_18233,N_18260);
or U20019 (N_20019,N_18733,N_18348);
nand U20020 (N_20020,N_19417,N_18104);
or U20021 (N_20021,N_18818,N_18389);
and U20022 (N_20022,N_18760,N_19098);
or U20023 (N_20023,N_19489,N_18214);
nor U20024 (N_20024,N_19488,N_18784);
and U20025 (N_20025,N_19335,N_18285);
xnor U20026 (N_20026,N_18443,N_18115);
xnor U20027 (N_20027,N_19160,N_18052);
nor U20028 (N_20028,N_18577,N_19206);
nand U20029 (N_20029,N_19401,N_18629);
xnor U20030 (N_20030,N_18769,N_18438);
or U20031 (N_20031,N_18054,N_19038);
or U20032 (N_20032,N_19138,N_18031);
xor U20033 (N_20033,N_19267,N_18537);
nor U20034 (N_20034,N_18294,N_18751);
nor U20035 (N_20035,N_18292,N_18073);
nand U20036 (N_20036,N_19150,N_18005);
nor U20037 (N_20037,N_19197,N_18812);
xor U20038 (N_20038,N_19234,N_19264);
nor U20039 (N_20039,N_18381,N_18074);
nand U20040 (N_20040,N_19292,N_18437);
nor U20041 (N_20041,N_19270,N_19017);
and U20042 (N_20042,N_18465,N_19000);
and U20043 (N_20043,N_18439,N_18177);
nor U20044 (N_20044,N_18551,N_18401);
xnor U20045 (N_20045,N_19111,N_19233);
nand U20046 (N_20046,N_19028,N_18135);
or U20047 (N_20047,N_18212,N_19235);
and U20048 (N_20048,N_19204,N_18485);
xnor U20049 (N_20049,N_18489,N_19187);
nand U20050 (N_20050,N_18166,N_19104);
xor U20051 (N_20051,N_19319,N_18471);
and U20052 (N_20052,N_18457,N_19212);
nor U20053 (N_20053,N_18040,N_18487);
xor U20054 (N_20054,N_19015,N_18473);
nor U20055 (N_20055,N_18648,N_18581);
nand U20056 (N_20056,N_19278,N_19446);
and U20057 (N_20057,N_19063,N_19132);
nor U20058 (N_20058,N_19026,N_18072);
and U20059 (N_20059,N_19020,N_18216);
or U20060 (N_20060,N_18625,N_18144);
nand U20061 (N_20061,N_18189,N_19023);
and U20062 (N_20062,N_18562,N_19337);
or U20063 (N_20063,N_19019,N_18025);
nand U20064 (N_20064,N_19327,N_19094);
xor U20065 (N_20065,N_18153,N_18290);
and U20066 (N_20066,N_18756,N_18188);
nor U20067 (N_20067,N_19200,N_18928);
nor U20068 (N_20068,N_18720,N_18359);
or U20069 (N_20069,N_18639,N_18570);
xor U20070 (N_20070,N_18258,N_18606);
nand U20071 (N_20071,N_18787,N_18862);
nor U20072 (N_20072,N_18870,N_19162);
nand U20073 (N_20073,N_18838,N_18881);
nand U20074 (N_20074,N_18965,N_19054);
and U20075 (N_20075,N_18614,N_18640);
nor U20076 (N_20076,N_19013,N_18742);
nor U20077 (N_20077,N_18735,N_18230);
nand U20078 (N_20078,N_18308,N_18680);
nand U20079 (N_20079,N_18722,N_18169);
nand U20080 (N_20080,N_19253,N_19444);
nand U20081 (N_20081,N_19364,N_18977);
or U20082 (N_20082,N_19303,N_18927);
nand U20083 (N_20083,N_18982,N_18172);
nor U20084 (N_20084,N_19298,N_18006);
nand U20085 (N_20085,N_18195,N_19391);
xor U20086 (N_20086,N_18375,N_18991);
xnor U20087 (N_20087,N_18727,N_18653);
and U20088 (N_20088,N_18058,N_18696);
nand U20089 (N_20089,N_19338,N_18835);
xor U20090 (N_20090,N_19413,N_18894);
nor U20091 (N_20091,N_18986,N_19305);
and U20092 (N_20092,N_19012,N_18845);
xnor U20093 (N_20093,N_18138,N_18330);
xor U20094 (N_20094,N_18929,N_19299);
xnor U20095 (N_20095,N_18335,N_18830);
nand U20096 (N_20096,N_18825,N_18317);
and U20097 (N_20097,N_19242,N_19290);
nand U20098 (N_20098,N_18356,N_19009);
nand U20099 (N_20099,N_19205,N_19366);
nor U20100 (N_20100,N_19496,N_18995);
nor U20101 (N_20101,N_19463,N_18873);
xnor U20102 (N_20102,N_19340,N_18745);
or U20103 (N_20103,N_18202,N_18855);
xnor U20104 (N_20104,N_18799,N_18228);
nor U20105 (N_20105,N_18820,N_18030);
xor U20106 (N_20106,N_18333,N_18968);
nand U20107 (N_20107,N_18961,N_19432);
or U20108 (N_20108,N_19003,N_18976);
nor U20109 (N_20109,N_19469,N_18015);
nand U20110 (N_20110,N_18952,N_18841);
or U20111 (N_20111,N_18668,N_19220);
xnor U20112 (N_20112,N_18910,N_18882);
nor U20113 (N_20113,N_18227,N_18164);
nand U20114 (N_20114,N_18691,N_19400);
xnor U20115 (N_20115,N_19285,N_18445);
or U20116 (N_20116,N_18558,N_18288);
xnor U20117 (N_20117,N_18960,N_18946);
nand U20118 (N_20118,N_18157,N_18198);
and U20119 (N_20119,N_19190,N_18385);
xor U20120 (N_20120,N_19129,N_19476);
nor U20121 (N_20121,N_18431,N_19034);
or U20122 (N_20122,N_18842,N_18309);
or U20123 (N_20123,N_18847,N_18880);
xor U20124 (N_20124,N_18813,N_18143);
xnor U20125 (N_20125,N_18772,N_18576);
nand U20126 (N_20126,N_19218,N_19198);
or U20127 (N_20127,N_18944,N_18009);
nor U20128 (N_20128,N_18117,N_18619);
and U20129 (N_20129,N_18679,N_19195);
nor U20130 (N_20130,N_19494,N_19341);
nand U20131 (N_20131,N_18427,N_19024);
nor U20132 (N_20132,N_19146,N_18584);
nand U20133 (N_20133,N_18765,N_18832);
nand U20134 (N_20134,N_19049,N_19458);
or U20135 (N_20135,N_18686,N_19169);
xor U20136 (N_20136,N_18021,N_18311);
or U20137 (N_20137,N_18764,N_18729);
or U20138 (N_20138,N_19385,N_18297);
nand U20139 (N_20139,N_18124,N_18591);
nor U20140 (N_20140,N_18937,N_18120);
or U20141 (N_20141,N_19080,N_18925);
nor U20142 (N_20142,N_18277,N_19238);
xor U20143 (N_20143,N_18354,N_18510);
xnor U20144 (N_20144,N_19057,N_18383);
nand U20145 (N_20145,N_18242,N_18575);
nand U20146 (N_20146,N_18804,N_18833);
xnor U20147 (N_20147,N_18721,N_18282);
or U20148 (N_20148,N_18134,N_18525);
nor U20149 (N_20149,N_18698,N_18900);
xor U20150 (N_20150,N_19448,N_18468);
xor U20151 (N_20151,N_18327,N_19415);
nor U20152 (N_20152,N_18706,N_19001);
and U20153 (N_20153,N_18533,N_18647);
nand U20154 (N_20154,N_18514,N_18791);
or U20155 (N_20155,N_19313,N_18119);
nand U20156 (N_20156,N_18379,N_18013);
nor U20157 (N_20157,N_18996,N_18378);
nand U20158 (N_20158,N_18343,N_18291);
and U20159 (N_20159,N_18155,N_19185);
nand U20160 (N_20160,N_18133,N_18766);
nor U20161 (N_20161,N_19144,N_18646);
and U20162 (N_20162,N_19240,N_18109);
nor U20163 (N_20163,N_18116,N_18743);
xnor U20164 (N_20164,N_18123,N_19392);
nand U20165 (N_20165,N_18316,N_19301);
and U20166 (N_20166,N_18964,N_18754);
or U20167 (N_20167,N_18049,N_19374);
xor U20168 (N_20168,N_19051,N_18296);
nand U20169 (N_20169,N_18325,N_19373);
or U20170 (N_20170,N_18536,N_18122);
xnor U20171 (N_20171,N_19454,N_19224);
xnor U20172 (N_20172,N_19461,N_18105);
nor U20173 (N_20173,N_19085,N_18014);
and U20174 (N_20174,N_19424,N_19139);
nand U20175 (N_20175,N_18128,N_18511);
or U20176 (N_20176,N_18092,N_18701);
or U20177 (N_20177,N_18363,N_18112);
nand U20178 (N_20178,N_18099,N_18496);
nand U20179 (N_20179,N_18861,N_18599);
or U20180 (N_20180,N_19191,N_18767);
and U20181 (N_20181,N_18627,N_19451);
and U20182 (N_20182,N_19453,N_19199);
nor U20183 (N_20183,N_18208,N_18331);
xor U20184 (N_20184,N_19133,N_19110);
and U20185 (N_20185,N_18266,N_19076);
or U20186 (N_20186,N_18150,N_18600);
nor U20187 (N_20187,N_18020,N_18240);
nand U20188 (N_20188,N_19349,N_19309);
xor U20189 (N_20189,N_19457,N_19383);
or U20190 (N_20190,N_18065,N_18397);
and U20191 (N_20191,N_18315,N_18235);
and U20192 (N_20192,N_18502,N_18103);
and U20193 (N_20193,N_18560,N_18885);
or U20194 (N_20194,N_18527,N_19056);
xnor U20195 (N_20195,N_18768,N_18858);
nand U20196 (N_20196,N_18573,N_18126);
or U20197 (N_20197,N_19151,N_19052);
xor U20198 (N_20198,N_19318,N_18574);
or U20199 (N_20199,N_18557,N_19141);
and U20200 (N_20200,N_18417,N_19122);
nand U20201 (N_20201,N_18127,N_18037);
and U20202 (N_20202,N_18422,N_19254);
nor U20203 (N_20203,N_18312,N_18429);
nand U20204 (N_20204,N_18587,N_18988);
and U20205 (N_20205,N_19167,N_18107);
and U20206 (N_20206,N_18447,N_18042);
nand U20207 (N_20207,N_18456,N_19179);
nor U20208 (N_20208,N_19371,N_18796);
or U20209 (N_20209,N_18089,N_19103);
xnor U20210 (N_20210,N_19252,N_18826);
xnor U20211 (N_20211,N_19255,N_18757);
nor U20212 (N_20212,N_18731,N_18425);
xnor U20213 (N_20213,N_18704,N_18739);
nand U20214 (N_20214,N_18017,N_19002);
and U20215 (N_20215,N_18687,N_19326);
or U20216 (N_20216,N_18598,N_19245);
nand U20217 (N_20217,N_18490,N_18132);
nor U20218 (N_20218,N_18407,N_19445);
xor U20219 (N_20219,N_19259,N_18677);
nor U20220 (N_20220,N_18371,N_18298);
xnor U20221 (N_20221,N_19492,N_19365);
xnor U20222 (N_20222,N_19130,N_18226);
nand U20223 (N_20223,N_19155,N_19077);
and U20224 (N_20224,N_19183,N_18672);
and U20225 (N_20225,N_18554,N_19215);
and U20226 (N_20226,N_19465,N_19449);
xor U20227 (N_20227,N_18158,N_18656);
or U20228 (N_20228,N_18746,N_18607);
nor U20229 (N_20229,N_19485,N_18403);
and U20230 (N_20230,N_18265,N_19228);
nand U20231 (N_20231,N_18789,N_18464);
nor U20232 (N_20232,N_18734,N_18141);
xnor U20233 (N_20233,N_18391,N_18752);
xnor U20234 (N_20234,N_19440,N_19480);
nand U20235 (N_20235,N_18322,N_18200);
and U20236 (N_20236,N_19031,N_18750);
xor U20237 (N_20237,N_18400,N_18184);
and U20238 (N_20238,N_18612,N_19161);
xnor U20239 (N_20239,N_19006,N_18592);
xnor U20240 (N_20240,N_18770,N_18027);
or U20241 (N_20241,N_19182,N_19073);
xor U20242 (N_20242,N_18231,N_18137);
and U20243 (N_20243,N_19172,N_18409);
xor U20244 (N_20244,N_18271,N_18106);
and U20245 (N_20245,N_19381,N_19481);
xor U20246 (N_20246,N_18856,N_18337);
nor U20247 (N_20247,N_18702,N_19350);
nand U20248 (N_20248,N_18868,N_18817);
nand U20249 (N_20249,N_18279,N_18895);
xor U20250 (N_20250,N_19350,N_18006);
xor U20251 (N_20251,N_19019,N_18162);
xor U20252 (N_20252,N_18984,N_19341);
xnor U20253 (N_20253,N_19158,N_18015);
and U20254 (N_20254,N_19411,N_19338);
nor U20255 (N_20255,N_18169,N_19149);
and U20256 (N_20256,N_18888,N_18015);
nor U20257 (N_20257,N_19279,N_18689);
or U20258 (N_20258,N_18671,N_18103);
xnor U20259 (N_20259,N_18333,N_19045);
nor U20260 (N_20260,N_19240,N_18551);
nand U20261 (N_20261,N_18757,N_18675);
nor U20262 (N_20262,N_18878,N_18993);
nand U20263 (N_20263,N_18797,N_19336);
and U20264 (N_20264,N_18862,N_18084);
nand U20265 (N_20265,N_19136,N_19369);
nor U20266 (N_20266,N_19267,N_18575);
xor U20267 (N_20267,N_19027,N_18913);
and U20268 (N_20268,N_19261,N_18105);
or U20269 (N_20269,N_18442,N_18109);
nor U20270 (N_20270,N_18926,N_18668);
and U20271 (N_20271,N_18182,N_18434);
xor U20272 (N_20272,N_18783,N_19371);
and U20273 (N_20273,N_18848,N_19001);
xor U20274 (N_20274,N_19214,N_19344);
nand U20275 (N_20275,N_18909,N_18503);
or U20276 (N_20276,N_19281,N_18588);
or U20277 (N_20277,N_18931,N_18560);
or U20278 (N_20278,N_18642,N_18847);
and U20279 (N_20279,N_18638,N_18265);
nand U20280 (N_20280,N_18251,N_18109);
nand U20281 (N_20281,N_18526,N_18427);
nand U20282 (N_20282,N_19050,N_18234);
nor U20283 (N_20283,N_18466,N_18346);
nor U20284 (N_20284,N_19237,N_19192);
and U20285 (N_20285,N_18311,N_19188);
or U20286 (N_20286,N_18840,N_18069);
or U20287 (N_20287,N_18617,N_18921);
nor U20288 (N_20288,N_19467,N_19380);
xnor U20289 (N_20289,N_19488,N_18698);
xor U20290 (N_20290,N_18621,N_18246);
or U20291 (N_20291,N_18619,N_18876);
nor U20292 (N_20292,N_19415,N_18938);
or U20293 (N_20293,N_19307,N_19462);
xnor U20294 (N_20294,N_18904,N_19136);
and U20295 (N_20295,N_18268,N_18664);
nand U20296 (N_20296,N_18071,N_18870);
nor U20297 (N_20297,N_18443,N_19075);
nor U20298 (N_20298,N_18919,N_19324);
or U20299 (N_20299,N_19088,N_19377);
xor U20300 (N_20300,N_19480,N_19419);
or U20301 (N_20301,N_18949,N_18684);
nand U20302 (N_20302,N_19194,N_18029);
xor U20303 (N_20303,N_18974,N_18968);
or U20304 (N_20304,N_18141,N_18649);
and U20305 (N_20305,N_19204,N_19100);
xor U20306 (N_20306,N_19206,N_18195);
nor U20307 (N_20307,N_18089,N_18751);
nor U20308 (N_20308,N_18231,N_19287);
xnor U20309 (N_20309,N_18617,N_18664);
nor U20310 (N_20310,N_18441,N_18535);
or U20311 (N_20311,N_18597,N_18106);
nand U20312 (N_20312,N_18999,N_18971);
xnor U20313 (N_20313,N_18525,N_18168);
nor U20314 (N_20314,N_18804,N_18741);
nor U20315 (N_20315,N_19406,N_19023);
xor U20316 (N_20316,N_18803,N_19066);
nor U20317 (N_20317,N_18399,N_19085);
and U20318 (N_20318,N_19350,N_18537);
or U20319 (N_20319,N_18547,N_19151);
nand U20320 (N_20320,N_18980,N_19211);
and U20321 (N_20321,N_18820,N_18699);
or U20322 (N_20322,N_19473,N_18230);
xor U20323 (N_20323,N_18091,N_19188);
nand U20324 (N_20324,N_18992,N_18986);
nand U20325 (N_20325,N_19163,N_18215);
or U20326 (N_20326,N_19154,N_18848);
xnor U20327 (N_20327,N_18725,N_18216);
and U20328 (N_20328,N_18135,N_18974);
nand U20329 (N_20329,N_19078,N_18634);
xor U20330 (N_20330,N_18016,N_18318);
or U20331 (N_20331,N_19052,N_19195);
nor U20332 (N_20332,N_19451,N_18332);
nor U20333 (N_20333,N_18448,N_18099);
or U20334 (N_20334,N_18391,N_18018);
or U20335 (N_20335,N_19035,N_18664);
or U20336 (N_20336,N_18497,N_19363);
or U20337 (N_20337,N_18376,N_18293);
or U20338 (N_20338,N_18817,N_18899);
nor U20339 (N_20339,N_19009,N_18435);
and U20340 (N_20340,N_19272,N_18258);
nor U20341 (N_20341,N_18618,N_19253);
nor U20342 (N_20342,N_18423,N_18363);
xnor U20343 (N_20343,N_18698,N_18036);
nand U20344 (N_20344,N_18398,N_19391);
xnor U20345 (N_20345,N_18194,N_18850);
or U20346 (N_20346,N_18682,N_19389);
nor U20347 (N_20347,N_18608,N_18654);
nor U20348 (N_20348,N_18719,N_18178);
nand U20349 (N_20349,N_18170,N_18607);
and U20350 (N_20350,N_18657,N_19010);
xnor U20351 (N_20351,N_18702,N_18740);
nor U20352 (N_20352,N_18552,N_18752);
nor U20353 (N_20353,N_18595,N_19142);
and U20354 (N_20354,N_18921,N_18608);
and U20355 (N_20355,N_18303,N_19284);
xnor U20356 (N_20356,N_19123,N_18776);
nand U20357 (N_20357,N_18083,N_18004);
nor U20358 (N_20358,N_18641,N_19207);
and U20359 (N_20359,N_18450,N_19446);
nor U20360 (N_20360,N_19244,N_18484);
nor U20361 (N_20361,N_19307,N_18235);
xor U20362 (N_20362,N_19271,N_18783);
xnor U20363 (N_20363,N_19427,N_18640);
or U20364 (N_20364,N_18980,N_18111);
or U20365 (N_20365,N_18649,N_19068);
and U20366 (N_20366,N_18983,N_18176);
xnor U20367 (N_20367,N_19212,N_18686);
nand U20368 (N_20368,N_19425,N_18256);
nor U20369 (N_20369,N_18816,N_19248);
xnor U20370 (N_20370,N_18906,N_18193);
nand U20371 (N_20371,N_18114,N_19280);
nor U20372 (N_20372,N_18264,N_18329);
nor U20373 (N_20373,N_19435,N_18102);
nand U20374 (N_20374,N_18871,N_18327);
nor U20375 (N_20375,N_18169,N_18051);
and U20376 (N_20376,N_18567,N_19130);
xnor U20377 (N_20377,N_18298,N_19290);
xor U20378 (N_20378,N_18019,N_18385);
or U20379 (N_20379,N_18024,N_18306);
and U20380 (N_20380,N_19183,N_18314);
xnor U20381 (N_20381,N_18373,N_18297);
xor U20382 (N_20382,N_19106,N_19091);
or U20383 (N_20383,N_19401,N_18743);
xor U20384 (N_20384,N_18271,N_19305);
nand U20385 (N_20385,N_19372,N_18040);
and U20386 (N_20386,N_18676,N_18130);
nand U20387 (N_20387,N_18874,N_18011);
nand U20388 (N_20388,N_18806,N_19360);
or U20389 (N_20389,N_18377,N_18301);
and U20390 (N_20390,N_18888,N_18814);
or U20391 (N_20391,N_18053,N_18439);
xnor U20392 (N_20392,N_18132,N_19308);
xnor U20393 (N_20393,N_18513,N_18446);
and U20394 (N_20394,N_18887,N_19064);
and U20395 (N_20395,N_18765,N_19064);
xnor U20396 (N_20396,N_18091,N_19192);
and U20397 (N_20397,N_19332,N_18803);
nand U20398 (N_20398,N_18763,N_18379);
and U20399 (N_20399,N_18636,N_18570);
or U20400 (N_20400,N_19444,N_18776);
nand U20401 (N_20401,N_18856,N_19070);
nor U20402 (N_20402,N_19320,N_18515);
or U20403 (N_20403,N_18142,N_18977);
nor U20404 (N_20404,N_18171,N_19104);
and U20405 (N_20405,N_19025,N_18314);
nor U20406 (N_20406,N_18185,N_18420);
nand U20407 (N_20407,N_18183,N_18140);
nand U20408 (N_20408,N_18601,N_19213);
xnor U20409 (N_20409,N_18662,N_18440);
nor U20410 (N_20410,N_18873,N_18384);
nand U20411 (N_20411,N_19126,N_18436);
xnor U20412 (N_20412,N_19097,N_18383);
nor U20413 (N_20413,N_19016,N_18477);
or U20414 (N_20414,N_19195,N_18629);
and U20415 (N_20415,N_19388,N_18910);
nand U20416 (N_20416,N_19319,N_18984);
or U20417 (N_20417,N_18348,N_18863);
nand U20418 (N_20418,N_19290,N_19024);
nand U20419 (N_20419,N_19188,N_18746);
nor U20420 (N_20420,N_18922,N_19109);
nor U20421 (N_20421,N_18542,N_18000);
and U20422 (N_20422,N_18617,N_18171);
and U20423 (N_20423,N_19130,N_18737);
nor U20424 (N_20424,N_18960,N_18335);
xnor U20425 (N_20425,N_18245,N_18777);
or U20426 (N_20426,N_18463,N_18095);
or U20427 (N_20427,N_19137,N_19422);
nor U20428 (N_20428,N_18273,N_18011);
nand U20429 (N_20429,N_18563,N_19279);
xnor U20430 (N_20430,N_19454,N_19313);
xor U20431 (N_20431,N_18201,N_18479);
nand U20432 (N_20432,N_18722,N_18599);
or U20433 (N_20433,N_18299,N_18694);
or U20434 (N_20434,N_18399,N_19224);
nor U20435 (N_20435,N_18600,N_18838);
and U20436 (N_20436,N_18656,N_18868);
or U20437 (N_20437,N_18464,N_19127);
xnor U20438 (N_20438,N_19350,N_19323);
xnor U20439 (N_20439,N_18277,N_18577);
and U20440 (N_20440,N_18419,N_18281);
nand U20441 (N_20441,N_18450,N_18113);
nand U20442 (N_20442,N_19346,N_18806);
nand U20443 (N_20443,N_18143,N_18072);
xnor U20444 (N_20444,N_19215,N_19255);
or U20445 (N_20445,N_18543,N_19463);
or U20446 (N_20446,N_19229,N_19038);
xor U20447 (N_20447,N_18122,N_18978);
and U20448 (N_20448,N_18849,N_18994);
nand U20449 (N_20449,N_18410,N_19325);
nor U20450 (N_20450,N_19340,N_18412);
nand U20451 (N_20451,N_19187,N_18598);
and U20452 (N_20452,N_18116,N_19260);
nor U20453 (N_20453,N_19253,N_19161);
or U20454 (N_20454,N_18701,N_18204);
xor U20455 (N_20455,N_19102,N_19105);
nand U20456 (N_20456,N_18016,N_18201);
and U20457 (N_20457,N_18967,N_18074);
nor U20458 (N_20458,N_18128,N_19101);
nor U20459 (N_20459,N_18749,N_18279);
nand U20460 (N_20460,N_18570,N_19469);
nand U20461 (N_20461,N_18988,N_18899);
nor U20462 (N_20462,N_18994,N_19474);
nor U20463 (N_20463,N_18653,N_19139);
and U20464 (N_20464,N_18607,N_18446);
or U20465 (N_20465,N_18529,N_19114);
nor U20466 (N_20466,N_18954,N_19431);
nand U20467 (N_20467,N_18842,N_19090);
nor U20468 (N_20468,N_18329,N_18697);
or U20469 (N_20469,N_18704,N_18995);
and U20470 (N_20470,N_18891,N_18367);
and U20471 (N_20471,N_18129,N_19102);
nand U20472 (N_20472,N_19481,N_19059);
xnor U20473 (N_20473,N_18684,N_18796);
nor U20474 (N_20474,N_18067,N_18296);
xnor U20475 (N_20475,N_19383,N_18303);
and U20476 (N_20476,N_18283,N_18848);
nand U20477 (N_20477,N_18916,N_19066);
or U20478 (N_20478,N_19407,N_18645);
and U20479 (N_20479,N_19166,N_19245);
and U20480 (N_20480,N_18278,N_18152);
and U20481 (N_20481,N_18630,N_18873);
nor U20482 (N_20482,N_18280,N_18711);
nor U20483 (N_20483,N_18363,N_18540);
xor U20484 (N_20484,N_19451,N_18018);
nor U20485 (N_20485,N_18557,N_19261);
nand U20486 (N_20486,N_18774,N_19126);
and U20487 (N_20487,N_18030,N_18195);
nand U20488 (N_20488,N_18296,N_19022);
or U20489 (N_20489,N_18655,N_18443);
nor U20490 (N_20490,N_19450,N_18421);
and U20491 (N_20491,N_19450,N_18944);
and U20492 (N_20492,N_19347,N_18071);
nand U20493 (N_20493,N_19011,N_18243);
nor U20494 (N_20494,N_19140,N_19424);
nand U20495 (N_20495,N_19339,N_18651);
nor U20496 (N_20496,N_18777,N_18917);
nand U20497 (N_20497,N_18968,N_18223);
nor U20498 (N_20498,N_18984,N_18195);
or U20499 (N_20499,N_18682,N_19292);
or U20500 (N_20500,N_18692,N_18823);
nand U20501 (N_20501,N_19397,N_18444);
and U20502 (N_20502,N_19302,N_18233);
and U20503 (N_20503,N_19372,N_19319);
and U20504 (N_20504,N_19305,N_18237);
xor U20505 (N_20505,N_18640,N_18394);
nand U20506 (N_20506,N_19420,N_19377);
nor U20507 (N_20507,N_18650,N_18482);
xnor U20508 (N_20508,N_19469,N_18667);
and U20509 (N_20509,N_18136,N_18184);
nor U20510 (N_20510,N_19131,N_18118);
xor U20511 (N_20511,N_18987,N_18918);
and U20512 (N_20512,N_18485,N_19488);
nor U20513 (N_20513,N_18320,N_18885);
nand U20514 (N_20514,N_18875,N_18997);
nor U20515 (N_20515,N_18476,N_18187);
xor U20516 (N_20516,N_19431,N_18370);
xnor U20517 (N_20517,N_18894,N_19486);
nand U20518 (N_20518,N_19286,N_18426);
or U20519 (N_20519,N_18088,N_18616);
or U20520 (N_20520,N_19236,N_18803);
or U20521 (N_20521,N_19173,N_19184);
xor U20522 (N_20522,N_18006,N_18754);
and U20523 (N_20523,N_18746,N_18787);
or U20524 (N_20524,N_18977,N_18747);
nor U20525 (N_20525,N_18123,N_19422);
or U20526 (N_20526,N_18473,N_18938);
or U20527 (N_20527,N_19435,N_18758);
xnor U20528 (N_20528,N_18262,N_19220);
nand U20529 (N_20529,N_19449,N_18291);
or U20530 (N_20530,N_19398,N_18740);
or U20531 (N_20531,N_18472,N_18250);
and U20532 (N_20532,N_19391,N_18357);
or U20533 (N_20533,N_19145,N_19192);
xnor U20534 (N_20534,N_18352,N_18751);
or U20535 (N_20535,N_18023,N_18647);
or U20536 (N_20536,N_19107,N_18535);
and U20537 (N_20537,N_18972,N_19386);
and U20538 (N_20538,N_18235,N_18343);
and U20539 (N_20539,N_18017,N_18085);
nand U20540 (N_20540,N_19097,N_18048);
or U20541 (N_20541,N_18603,N_18650);
nand U20542 (N_20542,N_18269,N_18588);
nor U20543 (N_20543,N_19124,N_18987);
xnor U20544 (N_20544,N_18971,N_18008);
nand U20545 (N_20545,N_18663,N_18837);
nand U20546 (N_20546,N_18161,N_19308);
xor U20547 (N_20547,N_18869,N_18030);
nand U20548 (N_20548,N_18553,N_19044);
nor U20549 (N_20549,N_18614,N_18558);
xor U20550 (N_20550,N_18414,N_19182);
or U20551 (N_20551,N_18546,N_18471);
nand U20552 (N_20552,N_18475,N_18939);
nor U20553 (N_20553,N_18403,N_18825);
nor U20554 (N_20554,N_18226,N_18776);
and U20555 (N_20555,N_18179,N_19126);
or U20556 (N_20556,N_18466,N_18140);
nor U20557 (N_20557,N_18569,N_19434);
xor U20558 (N_20558,N_18340,N_18310);
nand U20559 (N_20559,N_19475,N_18986);
nand U20560 (N_20560,N_18068,N_19153);
xnor U20561 (N_20561,N_18303,N_18141);
nand U20562 (N_20562,N_18147,N_18669);
nor U20563 (N_20563,N_19119,N_18141);
nand U20564 (N_20564,N_18855,N_18352);
xnor U20565 (N_20565,N_19188,N_19113);
or U20566 (N_20566,N_18918,N_18158);
nand U20567 (N_20567,N_18305,N_18809);
nor U20568 (N_20568,N_19408,N_18443);
nor U20569 (N_20569,N_18287,N_18078);
and U20570 (N_20570,N_19179,N_18017);
or U20571 (N_20571,N_19007,N_19493);
and U20572 (N_20572,N_18719,N_18224);
or U20573 (N_20573,N_18655,N_18047);
nor U20574 (N_20574,N_18862,N_18378);
nand U20575 (N_20575,N_19399,N_19015);
nand U20576 (N_20576,N_18847,N_18721);
and U20577 (N_20577,N_18905,N_19072);
xnor U20578 (N_20578,N_18834,N_19452);
or U20579 (N_20579,N_18198,N_19425);
nor U20580 (N_20580,N_18813,N_18594);
nor U20581 (N_20581,N_19362,N_18277);
nand U20582 (N_20582,N_19409,N_18563);
nor U20583 (N_20583,N_19458,N_18374);
xor U20584 (N_20584,N_18969,N_18362);
and U20585 (N_20585,N_18572,N_19431);
nand U20586 (N_20586,N_19461,N_18214);
nor U20587 (N_20587,N_18613,N_18189);
nand U20588 (N_20588,N_18422,N_18606);
xor U20589 (N_20589,N_18890,N_18899);
nor U20590 (N_20590,N_18772,N_18147);
nand U20591 (N_20591,N_19434,N_19176);
and U20592 (N_20592,N_19278,N_18380);
nor U20593 (N_20593,N_18733,N_18448);
nor U20594 (N_20594,N_18622,N_18547);
nand U20595 (N_20595,N_18086,N_19272);
nor U20596 (N_20596,N_18489,N_18178);
and U20597 (N_20597,N_18308,N_18431);
nor U20598 (N_20598,N_18719,N_18511);
nor U20599 (N_20599,N_18337,N_19295);
and U20600 (N_20600,N_19254,N_18663);
nor U20601 (N_20601,N_18763,N_18236);
and U20602 (N_20602,N_18847,N_18212);
and U20603 (N_20603,N_18572,N_19399);
or U20604 (N_20604,N_19464,N_19154);
and U20605 (N_20605,N_18478,N_18372);
xnor U20606 (N_20606,N_18113,N_18851);
nand U20607 (N_20607,N_18029,N_18180);
nand U20608 (N_20608,N_18576,N_18783);
or U20609 (N_20609,N_18601,N_18366);
nor U20610 (N_20610,N_19492,N_18414);
and U20611 (N_20611,N_19251,N_18875);
nand U20612 (N_20612,N_18206,N_18526);
xor U20613 (N_20613,N_18356,N_18010);
or U20614 (N_20614,N_19394,N_19104);
xnor U20615 (N_20615,N_19408,N_18978);
xnor U20616 (N_20616,N_18127,N_18272);
and U20617 (N_20617,N_18149,N_19185);
nand U20618 (N_20618,N_18153,N_19046);
or U20619 (N_20619,N_19067,N_18843);
nor U20620 (N_20620,N_19163,N_18143);
or U20621 (N_20621,N_18838,N_18247);
or U20622 (N_20622,N_19206,N_18472);
nand U20623 (N_20623,N_19283,N_18809);
nand U20624 (N_20624,N_18124,N_18463);
or U20625 (N_20625,N_18635,N_19325);
xor U20626 (N_20626,N_18272,N_19209);
nor U20627 (N_20627,N_18594,N_19294);
and U20628 (N_20628,N_18577,N_18767);
nand U20629 (N_20629,N_18352,N_18083);
nor U20630 (N_20630,N_18223,N_18604);
and U20631 (N_20631,N_18438,N_18956);
and U20632 (N_20632,N_19167,N_18457);
nor U20633 (N_20633,N_18247,N_18849);
or U20634 (N_20634,N_19151,N_18791);
xnor U20635 (N_20635,N_18529,N_18900);
xor U20636 (N_20636,N_19366,N_18827);
and U20637 (N_20637,N_18312,N_18938);
xnor U20638 (N_20638,N_19122,N_19317);
and U20639 (N_20639,N_18881,N_18633);
or U20640 (N_20640,N_18793,N_18481);
nand U20641 (N_20641,N_19052,N_18567);
xor U20642 (N_20642,N_18299,N_18763);
or U20643 (N_20643,N_18976,N_18651);
and U20644 (N_20644,N_18691,N_18857);
nor U20645 (N_20645,N_18804,N_18532);
or U20646 (N_20646,N_18831,N_18010);
or U20647 (N_20647,N_19204,N_18207);
nor U20648 (N_20648,N_19046,N_19464);
nor U20649 (N_20649,N_18045,N_18505);
or U20650 (N_20650,N_18393,N_18993);
nor U20651 (N_20651,N_18561,N_18467);
nand U20652 (N_20652,N_18213,N_19418);
and U20653 (N_20653,N_18499,N_19356);
or U20654 (N_20654,N_19370,N_18479);
nor U20655 (N_20655,N_19205,N_18551);
and U20656 (N_20656,N_18791,N_19252);
nand U20657 (N_20657,N_19298,N_19028);
or U20658 (N_20658,N_19342,N_18272);
xnor U20659 (N_20659,N_18085,N_19223);
nand U20660 (N_20660,N_18493,N_18750);
or U20661 (N_20661,N_19227,N_19214);
xor U20662 (N_20662,N_18406,N_18223);
or U20663 (N_20663,N_19396,N_19198);
nor U20664 (N_20664,N_19310,N_18115);
or U20665 (N_20665,N_19125,N_18809);
nand U20666 (N_20666,N_18358,N_18347);
nand U20667 (N_20667,N_18950,N_18010);
and U20668 (N_20668,N_19338,N_18324);
or U20669 (N_20669,N_18325,N_18432);
nand U20670 (N_20670,N_18300,N_18094);
xnor U20671 (N_20671,N_19273,N_18931);
or U20672 (N_20672,N_18566,N_18623);
and U20673 (N_20673,N_18047,N_18551);
nand U20674 (N_20674,N_18716,N_18086);
and U20675 (N_20675,N_19243,N_19025);
nor U20676 (N_20676,N_18080,N_18444);
and U20677 (N_20677,N_18820,N_18871);
nand U20678 (N_20678,N_18993,N_18961);
xnor U20679 (N_20679,N_18950,N_19319);
nor U20680 (N_20680,N_19478,N_18999);
and U20681 (N_20681,N_19095,N_18302);
nor U20682 (N_20682,N_18760,N_19396);
xnor U20683 (N_20683,N_19150,N_19283);
and U20684 (N_20684,N_19213,N_18483);
nor U20685 (N_20685,N_19230,N_18090);
nand U20686 (N_20686,N_18646,N_19392);
xor U20687 (N_20687,N_19307,N_18302);
nor U20688 (N_20688,N_18345,N_18069);
or U20689 (N_20689,N_18976,N_18436);
xnor U20690 (N_20690,N_18631,N_18035);
nor U20691 (N_20691,N_18047,N_19469);
xor U20692 (N_20692,N_19167,N_18309);
and U20693 (N_20693,N_19487,N_18153);
nor U20694 (N_20694,N_18638,N_18833);
and U20695 (N_20695,N_18105,N_18346);
and U20696 (N_20696,N_18535,N_18486);
or U20697 (N_20697,N_18149,N_18167);
and U20698 (N_20698,N_19252,N_19281);
xnor U20699 (N_20699,N_18317,N_19435);
and U20700 (N_20700,N_19181,N_18574);
nand U20701 (N_20701,N_18789,N_18877);
xor U20702 (N_20702,N_18611,N_18243);
xnor U20703 (N_20703,N_18452,N_19305);
or U20704 (N_20704,N_19153,N_18863);
nand U20705 (N_20705,N_19050,N_18943);
nor U20706 (N_20706,N_18159,N_18685);
and U20707 (N_20707,N_18663,N_18375);
xor U20708 (N_20708,N_18095,N_18928);
and U20709 (N_20709,N_18808,N_19267);
nor U20710 (N_20710,N_18775,N_18235);
and U20711 (N_20711,N_18668,N_19335);
xor U20712 (N_20712,N_18778,N_18024);
and U20713 (N_20713,N_19010,N_19191);
xnor U20714 (N_20714,N_18538,N_18723);
and U20715 (N_20715,N_18381,N_18307);
and U20716 (N_20716,N_19100,N_18717);
or U20717 (N_20717,N_18101,N_19227);
xor U20718 (N_20718,N_19415,N_19455);
nand U20719 (N_20719,N_18620,N_18264);
nor U20720 (N_20720,N_18217,N_18021);
nand U20721 (N_20721,N_18365,N_19399);
nand U20722 (N_20722,N_18918,N_19062);
nand U20723 (N_20723,N_19469,N_18542);
and U20724 (N_20724,N_19078,N_19113);
xnor U20725 (N_20725,N_19109,N_19354);
nor U20726 (N_20726,N_19328,N_18796);
nand U20727 (N_20727,N_18097,N_19126);
or U20728 (N_20728,N_19256,N_18494);
nor U20729 (N_20729,N_19257,N_18768);
nor U20730 (N_20730,N_18190,N_18831);
xor U20731 (N_20731,N_19375,N_18931);
nand U20732 (N_20732,N_18229,N_19051);
nand U20733 (N_20733,N_18134,N_19285);
or U20734 (N_20734,N_18944,N_19313);
nand U20735 (N_20735,N_18166,N_18140);
xor U20736 (N_20736,N_18723,N_18940);
and U20737 (N_20737,N_18673,N_18710);
xor U20738 (N_20738,N_18695,N_18728);
xor U20739 (N_20739,N_18602,N_18192);
nor U20740 (N_20740,N_19404,N_19024);
or U20741 (N_20741,N_18139,N_18936);
and U20742 (N_20742,N_18452,N_18697);
xor U20743 (N_20743,N_18747,N_19320);
and U20744 (N_20744,N_19430,N_18639);
and U20745 (N_20745,N_19122,N_18011);
nor U20746 (N_20746,N_18429,N_19285);
nor U20747 (N_20747,N_19071,N_18491);
nand U20748 (N_20748,N_19083,N_18209);
xnor U20749 (N_20749,N_18165,N_18251);
nor U20750 (N_20750,N_18983,N_19365);
or U20751 (N_20751,N_18283,N_18734);
and U20752 (N_20752,N_18647,N_19304);
xor U20753 (N_20753,N_18833,N_18313);
nand U20754 (N_20754,N_18419,N_18843);
and U20755 (N_20755,N_18281,N_18545);
or U20756 (N_20756,N_18549,N_18565);
nor U20757 (N_20757,N_18119,N_18887);
or U20758 (N_20758,N_19333,N_18918);
nand U20759 (N_20759,N_18536,N_18443);
xor U20760 (N_20760,N_19072,N_18130);
and U20761 (N_20761,N_18018,N_18175);
nor U20762 (N_20762,N_19164,N_19356);
xnor U20763 (N_20763,N_18314,N_19168);
xnor U20764 (N_20764,N_18639,N_18017);
nor U20765 (N_20765,N_18698,N_18045);
nand U20766 (N_20766,N_18618,N_19276);
or U20767 (N_20767,N_18138,N_18458);
and U20768 (N_20768,N_19129,N_18946);
nand U20769 (N_20769,N_18420,N_19363);
or U20770 (N_20770,N_18943,N_19143);
xnor U20771 (N_20771,N_19364,N_18784);
nor U20772 (N_20772,N_19429,N_19441);
nand U20773 (N_20773,N_19084,N_18131);
nor U20774 (N_20774,N_18355,N_18670);
nand U20775 (N_20775,N_19109,N_18793);
or U20776 (N_20776,N_18182,N_18515);
xor U20777 (N_20777,N_18731,N_19018);
nor U20778 (N_20778,N_19494,N_18725);
nor U20779 (N_20779,N_18973,N_18646);
xnor U20780 (N_20780,N_18938,N_19175);
xor U20781 (N_20781,N_19327,N_18925);
xnor U20782 (N_20782,N_18422,N_18759);
nand U20783 (N_20783,N_18626,N_18716);
or U20784 (N_20784,N_19156,N_18336);
nand U20785 (N_20785,N_19305,N_19060);
or U20786 (N_20786,N_18560,N_19237);
and U20787 (N_20787,N_18976,N_19485);
nand U20788 (N_20788,N_18125,N_19413);
xor U20789 (N_20789,N_18240,N_18503);
or U20790 (N_20790,N_18265,N_18398);
xor U20791 (N_20791,N_18937,N_18639);
nor U20792 (N_20792,N_18436,N_18079);
nand U20793 (N_20793,N_18230,N_18237);
and U20794 (N_20794,N_18319,N_18055);
nor U20795 (N_20795,N_18923,N_18637);
or U20796 (N_20796,N_19258,N_18082);
nor U20797 (N_20797,N_19345,N_18703);
nor U20798 (N_20798,N_19232,N_18636);
xnor U20799 (N_20799,N_18145,N_18190);
and U20800 (N_20800,N_19240,N_18317);
nand U20801 (N_20801,N_18921,N_18839);
or U20802 (N_20802,N_18230,N_19403);
or U20803 (N_20803,N_19148,N_19039);
nor U20804 (N_20804,N_19187,N_19047);
and U20805 (N_20805,N_18980,N_18193);
nor U20806 (N_20806,N_18888,N_18984);
nand U20807 (N_20807,N_18273,N_19097);
or U20808 (N_20808,N_18906,N_18044);
or U20809 (N_20809,N_18705,N_18165);
or U20810 (N_20810,N_19076,N_19292);
and U20811 (N_20811,N_18859,N_18040);
and U20812 (N_20812,N_18809,N_18732);
and U20813 (N_20813,N_19488,N_18802);
and U20814 (N_20814,N_19096,N_19231);
or U20815 (N_20815,N_18185,N_18902);
nand U20816 (N_20816,N_18633,N_19464);
nor U20817 (N_20817,N_18540,N_19436);
nand U20818 (N_20818,N_18379,N_18990);
nor U20819 (N_20819,N_18176,N_18044);
nor U20820 (N_20820,N_18717,N_19175);
and U20821 (N_20821,N_18618,N_18135);
and U20822 (N_20822,N_19496,N_19052);
and U20823 (N_20823,N_18896,N_18253);
and U20824 (N_20824,N_18851,N_18229);
and U20825 (N_20825,N_18467,N_19321);
xnor U20826 (N_20826,N_18441,N_18822);
and U20827 (N_20827,N_19384,N_18906);
nor U20828 (N_20828,N_18145,N_19179);
and U20829 (N_20829,N_18433,N_18923);
nor U20830 (N_20830,N_18461,N_18093);
xnor U20831 (N_20831,N_19323,N_18928);
and U20832 (N_20832,N_18637,N_18607);
nor U20833 (N_20833,N_18319,N_18557);
and U20834 (N_20834,N_18424,N_19433);
nand U20835 (N_20835,N_19282,N_19001);
nor U20836 (N_20836,N_19292,N_18838);
nand U20837 (N_20837,N_18871,N_18762);
and U20838 (N_20838,N_18850,N_19012);
and U20839 (N_20839,N_18211,N_18295);
xnor U20840 (N_20840,N_18615,N_18425);
nand U20841 (N_20841,N_19182,N_18366);
and U20842 (N_20842,N_18396,N_18593);
or U20843 (N_20843,N_18595,N_18863);
or U20844 (N_20844,N_18875,N_19213);
nand U20845 (N_20845,N_18161,N_19379);
xor U20846 (N_20846,N_18564,N_19243);
nand U20847 (N_20847,N_18504,N_18061);
and U20848 (N_20848,N_19270,N_18175);
and U20849 (N_20849,N_19395,N_19393);
xnor U20850 (N_20850,N_19032,N_18430);
nand U20851 (N_20851,N_19006,N_18331);
xor U20852 (N_20852,N_19328,N_19395);
xor U20853 (N_20853,N_18284,N_18400);
and U20854 (N_20854,N_18434,N_18479);
nor U20855 (N_20855,N_19354,N_18296);
or U20856 (N_20856,N_18920,N_19179);
or U20857 (N_20857,N_18109,N_18837);
or U20858 (N_20858,N_19044,N_18292);
nor U20859 (N_20859,N_18110,N_18822);
nor U20860 (N_20860,N_19117,N_19308);
nand U20861 (N_20861,N_18016,N_18443);
nand U20862 (N_20862,N_18751,N_19353);
and U20863 (N_20863,N_18946,N_18028);
xor U20864 (N_20864,N_18523,N_18424);
or U20865 (N_20865,N_18185,N_19061);
nand U20866 (N_20866,N_19225,N_19154);
or U20867 (N_20867,N_18049,N_18824);
and U20868 (N_20868,N_18373,N_18969);
nor U20869 (N_20869,N_18281,N_18089);
or U20870 (N_20870,N_18485,N_19455);
nand U20871 (N_20871,N_18449,N_19170);
xor U20872 (N_20872,N_18832,N_18995);
or U20873 (N_20873,N_18805,N_19274);
or U20874 (N_20874,N_18386,N_18957);
nor U20875 (N_20875,N_18387,N_18702);
and U20876 (N_20876,N_19274,N_18678);
nor U20877 (N_20877,N_18714,N_18678);
nand U20878 (N_20878,N_19101,N_18204);
and U20879 (N_20879,N_19069,N_18432);
nand U20880 (N_20880,N_18401,N_18680);
and U20881 (N_20881,N_18881,N_18426);
nor U20882 (N_20882,N_19143,N_18784);
or U20883 (N_20883,N_19248,N_18813);
or U20884 (N_20884,N_18159,N_18055);
and U20885 (N_20885,N_18975,N_19420);
nand U20886 (N_20886,N_19243,N_18230);
or U20887 (N_20887,N_18892,N_19050);
nor U20888 (N_20888,N_18136,N_19145);
nand U20889 (N_20889,N_19414,N_19001);
nand U20890 (N_20890,N_18690,N_18043);
xnor U20891 (N_20891,N_18730,N_18328);
xnor U20892 (N_20892,N_18530,N_18785);
nand U20893 (N_20893,N_18704,N_18776);
and U20894 (N_20894,N_18458,N_19366);
or U20895 (N_20895,N_19404,N_19207);
xor U20896 (N_20896,N_19338,N_18769);
and U20897 (N_20897,N_18780,N_18140);
xnor U20898 (N_20898,N_19197,N_18115);
or U20899 (N_20899,N_18053,N_18327);
xnor U20900 (N_20900,N_18101,N_18246);
and U20901 (N_20901,N_18158,N_18228);
and U20902 (N_20902,N_18187,N_19348);
or U20903 (N_20903,N_19123,N_18649);
and U20904 (N_20904,N_19184,N_19491);
xnor U20905 (N_20905,N_19048,N_18884);
and U20906 (N_20906,N_18285,N_18458);
nand U20907 (N_20907,N_18842,N_18326);
and U20908 (N_20908,N_19192,N_19367);
xor U20909 (N_20909,N_18966,N_18918);
nor U20910 (N_20910,N_18929,N_19122);
and U20911 (N_20911,N_19318,N_18193);
nand U20912 (N_20912,N_18591,N_18318);
nor U20913 (N_20913,N_19391,N_18032);
nand U20914 (N_20914,N_19151,N_18801);
xnor U20915 (N_20915,N_18741,N_18528);
nor U20916 (N_20916,N_18505,N_18321);
and U20917 (N_20917,N_18894,N_19113);
and U20918 (N_20918,N_19386,N_19225);
and U20919 (N_20919,N_19313,N_18544);
or U20920 (N_20920,N_18409,N_18913);
and U20921 (N_20921,N_19202,N_19404);
or U20922 (N_20922,N_18500,N_19039);
nor U20923 (N_20923,N_18116,N_19322);
xor U20924 (N_20924,N_19038,N_18817);
nand U20925 (N_20925,N_18991,N_18466);
nand U20926 (N_20926,N_18399,N_18659);
and U20927 (N_20927,N_18145,N_18640);
and U20928 (N_20928,N_18652,N_19070);
xor U20929 (N_20929,N_18424,N_18962);
and U20930 (N_20930,N_18753,N_19359);
and U20931 (N_20931,N_18016,N_18189);
nor U20932 (N_20932,N_19210,N_18061);
or U20933 (N_20933,N_19169,N_18992);
nand U20934 (N_20934,N_18935,N_18763);
nor U20935 (N_20935,N_18763,N_19235);
or U20936 (N_20936,N_19209,N_18602);
nor U20937 (N_20937,N_18287,N_18037);
nor U20938 (N_20938,N_18806,N_18892);
nand U20939 (N_20939,N_18038,N_19329);
nand U20940 (N_20940,N_18982,N_18509);
nand U20941 (N_20941,N_19086,N_18407);
and U20942 (N_20942,N_18453,N_19116);
nand U20943 (N_20943,N_19260,N_19175);
nor U20944 (N_20944,N_19427,N_18310);
and U20945 (N_20945,N_18038,N_18572);
and U20946 (N_20946,N_18147,N_18612);
or U20947 (N_20947,N_18726,N_18807);
xnor U20948 (N_20948,N_18827,N_18775);
xnor U20949 (N_20949,N_18089,N_18861);
and U20950 (N_20950,N_18543,N_18096);
or U20951 (N_20951,N_18943,N_19476);
xnor U20952 (N_20952,N_18575,N_19307);
or U20953 (N_20953,N_18743,N_18834);
xnor U20954 (N_20954,N_19282,N_18721);
nor U20955 (N_20955,N_18846,N_19298);
nor U20956 (N_20956,N_18994,N_19272);
nand U20957 (N_20957,N_19305,N_18623);
nand U20958 (N_20958,N_18187,N_18594);
xnor U20959 (N_20959,N_19145,N_18806);
nor U20960 (N_20960,N_18859,N_18085);
nor U20961 (N_20961,N_18415,N_18085);
nand U20962 (N_20962,N_18930,N_19009);
and U20963 (N_20963,N_18782,N_19056);
nor U20964 (N_20964,N_19342,N_19353);
nand U20965 (N_20965,N_18612,N_18540);
and U20966 (N_20966,N_18189,N_18983);
and U20967 (N_20967,N_18833,N_18881);
or U20968 (N_20968,N_18596,N_19019);
nor U20969 (N_20969,N_19286,N_18323);
nor U20970 (N_20970,N_18643,N_18023);
and U20971 (N_20971,N_18922,N_19390);
and U20972 (N_20972,N_18890,N_19478);
and U20973 (N_20973,N_18587,N_18131);
xnor U20974 (N_20974,N_18326,N_18756);
xnor U20975 (N_20975,N_19173,N_19460);
nand U20976 (N_20976,N_18941,N_19482);
nor U20977 (N_20977,N_18368,N_18607);
or U20978 (N_20978,N_18920,N_19135);
nor U20979 (N_20979,N_19239,N_18825);
nor U20980 (N_20980,N_19135,N_18672);
and U20981 (N_20981,N_18939,N_18545);
and U20982 (N_20982,N_19272,N_19130);
nand U20983 (N_20983,N_19098,N_18611);
nand U20984 (N_20984,N_18382,N_18242);
xor U20985 (N_20985,N_19331,N_18354);
and U20986 (N_20986,N_18288,N_18875);
nor U20987 (N_20987,N_18992,N_19481);
or U20988 (N_20988,N_19098,N_18672);
nand U20989 (N_20989,N_19472,N_18218);
and U20990 (N_20990,N_19405,N_18637);
nand U20991 (N_20991,N_19156,N_18904);
or U20992 (N_20992,N_18397,N_18752);
or U20993 (N_20993,N_18529,N_19243);
xor U20994 (N_20994,N_18022,N_19077);
or U20995 (N_20995,N_18242,N_18935);
or U20996 (N_20996,N_18647,N_18529);
xor U20997 (N_20997,N_18985,N_19127);
xnor U20998 (N_20998,N_18499,N_19495);
or U20999 (N_20999,N_18183,N_18627);
or U21000 (N_21000,N_19994,N_19504);
nand U21001 (N_21001,N_20048,N_20450);
and U21002 (N_21002,N_20725,N_19765);
and U21003 (N_21003,N_20094,N_19606);
and U21004 (N_21004,N_20702,N_20408);
and U21005 (N_21005,N_20994,N_20834);
or U21006 (N_21006,N_20555,N_19851);
and U21007 (N_21007,N_19691,N_20789);
and U21008 (N_21008,N_20115,N_19710);
xnor U21009 (N_21009,N_20985,N_20025);
and U21010 (N_21010,N_20545,N_19758);
xnor U21011 (N_21011,N_20047,N_19783);
and U21012 (N_21012,N_20589,N_20677);
and U21013 (N_21013,N_20977,N_20631);
xnor U21014 (N_21014,N_20179,N_20422);
or U21015 (N_21015,N_19701,N_19870);
and U21016 (N_21016,N_19595,N_20301);
or U21017 (N_21017,N_20437,N_20142);
nand U21018 (N_21018,N_20594,N_20817);
or U21019 (N_21019,N_20137,N_20608);
and U21020 (N_21020,N_19978,N_19873);
and U21021 (N_21021,N_20713,N_20127);
or U21022 (N_21022,N_20723,N_20694);
nand U21023 (N_21023,N_19850,N_20225);
or U21024 (N_21024,N_20216,N_19591);
xor U21025 (N_21025,N_20377,N_20925);
nand U21026 (N_21026,N_20520,N_20051);
nand U21027 (N_21027,N_19807,N_20507);
nor U21028 (N_21028,N_20685,N_19541);
xor U21029 (N_21029,N_20361,N_20891);
or U21030 (N_21030,N_20903,N_20476);
xor U21031 (N_21031,N_20441,N_20270);
xnor U21032 (N_21032,N_19611,N_20168);
xnor U21033 (N_21033,N_20544,N_20705);
nand U21034 (N_21034,N_20516,N_20350);
nor U21035 (N_21035,N_19587,N_20799);
nand U21036 (N_21036,N_20831,N_20488);
nor U21037 (N_21037,N_20633,N_19969);
nand U21038 (N_21038,N_20921,N_20731);
or U21039 (N_21039,N_19584,N_19776);
xor U21040 (N_21040,N_19906,N_20104);
nor U21041 (N_21041,N_20357,N_20315);
or U21042 (N_21042,N_20280,N_20808);
or U21043 (N_21043,N_19703,N_20021);
or U21044 (N_21044,N_20722,N_20889);
nand U21045 (N_21045,N_20401,N_20188);
xor U21046 (N_21046,N_19940,N_20390);
xnor U21047 (N_21047,N_20071,N_19980);
nor U21048 (N_21048,N_20346,N_20648);
xor U21049 (N_21049,N_19853,N_20468);
or U21050 (N_21050,N_19864,N_19986);
nor U21051 (N_21051,N_20028,N_20046);
nor U21052 (N_21052,N_19533,N_20656);
and U21053 (N_21053,N_20867,N_20974);
xnor U21054 (N_21054,N_20861,N_20165);
or U21055 (N_21055,N_20029,N_20269);
xnor U21056 (N_21056,N_20092,N_20768);
and U21057 (N_21057,N_20879,N_20514);
nand U21058 (N_21058,N_19550,N_20440);
xnor U21059 (N_21059,N_20014,N_20411);
nor U21060 (N_21060,N_20463,N_19734);
nand U21061 (N_21061,N_20486,N_20090);
or U21062 (N_21062,N_20982,N_20676);
nand U21063 (N_21063,N_20809,N_20709);
and U21064 (N_21064,N_19952,N_20885);
and U21065 (N_21065,N_20583,N_20192);
and U21066 (N_21066,N_20948,N_19542);
or U21067 (N_21067,N_19847,N_20448);
xnor U21068 (N_21068,N_20250,N_19804);
and U21069 (N_21069,N_19823,N_20968);
xor U21070 (N_21070,N_19537,N_20642);
xor U21071 (N_21071,N_19732,N_20240);
xnor U21072 (N_21072,N_20329,N_20851);
or U21073 (N_21073,N_20364,N_20863);
and U21074 (N_21074,N_19770,N_20752);
or U21075 (N_21075,N_20331,N_20060);
nor U21076 (N_21076,N_20193,N_20595);
nand U21077 (N_21077,N_20576,N_19661);
or U21078 (N_21078,N_20271,N_20763);
nor U21079 (N_21079,N_20119,N_20133);
nand U21080 (N_21080,N_19996,N_20996);
and U21081 (N_21081,N_19902,N_19859);
nor U21082 (N_21082,N_20610,N_20614);
nand U21083 (N_21083,N_19630,N_20868);
xnor U21084 (N_21084,N_20366,N_19957);
nor U21085 (N_21085,N_19757,N_20762);
xor U21086 (N_21086,N_20181,N_20754);
nand U21087 (N_21087,N_19811,N_20393);
nor U21088 (N_21088,N_20522,N_20016);
and U21089 (N_21089,N_20637,N_20742);
xnor U21090 (N_21090,N_20805,N_19547);
xnor U21091 (N_21091,N_19916,N_19764);
xor U21092 (N_21092,N_20811,N_20733);
nor U21093 (N_21093,N_20321,N_20382);
nor U21094 (N_21094,N_19545,N_20551);
xor U21095 (N_21095,N_19627,N_20552);
and U21096 (N_21096,N_19629,N_20509);
nand U21097 (N_21097,N_20939,N_19888);
nand U21098 (N_21098,N_20954,N_20823);
and U21099 (N_21099,N_20207,N_19683);
and U21100 (N_21100,N_20340,N_20553);
or U21101 (N_21101,N_20532,N_20945);
and U21102 (N_21102,N_20353,N_20936);
or U21103 (N_21103,N_19785,N_20172);
or U21104 (N_21104,N_19670,N_20730);
xor U21105 (N_21105,N_20955,N_20472);
xnor U21106 (N_21106,N_20881,N_20727);
or U21107 (N_21107,N_19941,N_20276);
and U21108 (N_21108,N_20618,N_20537);
and U21109 (N_21109,N_20989,N_20031);
and U21110 (N_21110,N_19604,N_19919);
nor U21111 (N_21111,N_19860,N_20132);
nand U21112 (N_21112,N_19731,N_19886);
nand U21113 (N_21113,N_20083,N_19557);
xor U21114 (N_21114,N_19838,N_20547);
nor U21115 (N_21115,N_19963,N_20420);
nand U21116 (N_21116,N_20439,N_20452);
and U21117 (N_21117,N_19951,N_19964);
nand U21118 (N_21118,N_20004,N_20086);
xor U21119 (N_21119,N_20371,N_20026);
and U21120 (N_21120,N_20978,N_19645);
xnor U21121 (N_21121,N_19740,N_19707);
xnor U21122 (N_21122,N_20146,N_20466);
nand U21123 (N_21123,N_20233,N_19700);
nand U21124 (N_21124,N_20624,N_20895);
nand U21125 (N_21125,N_19928,N_19739);
nor U21126 (N_21126,N_19997,N_19880);
or U21127 (N_21127,N_19631,N_20039);
or U21128 (N_21128,N_20123,N_19531);
and U21129 (N_21129,N_19846,N_20342);
and U21130 (N_21130,N_20375,N_20517);
and U21131 (N_21131,N_20980,N_20592);
nor U21132 (N_21132,N_20061,N_20419);
or U21133 (N_21133,N_20432,N_20647);
and U21134 (N_21134,N_19681,N_19946);
nand U21135 (N_21135,N_20837,N_20523);
xnor U21136 (N_21136,N_20822,N_20926);
xor U21137 (N_21137,N_20332,N_19589);
nor U21138 (N_21138,N_20510,N_20367);
xnor U21139 (N_21139,N_20392,N_20971);
xnor U21140 (N_21140,N_20764,N_19500);
nor U21141 (N_21141,N_20872,N_20780);
nor U21142 (N_21142,N_20154,N_19634);
and U21143 (N_21143,N_20745,N_19717);
nand U21144 (N_21144,N_19521,N_19721);
nand U21145 (N_21145,N_20447,N_20562);
or U21146 (N_21146,N_20120,N_19948);
or U21147 (N_21147,N_19979,N_20044);
nor U21148 (N_21148,N_19876,N_19834);
xnor U21149 (N_21149,N_20384,N_20087);
and U21150 (N_21150,N_19745,N_19741);
xor U21151 (N_21151,N_20534,N_20473);
or U21152 (N_21152,N_19861,N_20904);
or U21153 (N_21153,N_19865,N_20073);
nand U21154 (N_21154,N_19883,N_19802);
nand U21155 (N_21155,N_20591,N_19977);
nor U21156 (N_21156,N_20857,N_19844);
and U21157 (N_21157,N_19815,N_19863);
nor U21158 (N_21158,N_20289,N_20222);
xnor U21159 (N_21159,N_20006,N_19644);
and U21160 (N_21160,N_20674,N_19839);
xnor U21161 (N_21161,N_19666,N_19549);
or U21162 (N_21162,N_19506,N_20063);
or U21163 (N_21163,N_20178,N_19563);
nor U21164 (N_21164,N_19704,N_20295);
xnor U21165 (N_21165,N_20262,N_20721);
nor U21166 (N_21166,N_19773,N_20199);
xnor U21167 (N_21167,N_19760,N_19821);
nor U21168 (N_21168,N_19950,N_20264);
and U21169 (N_21169,N_19553,N_20910);
nand U21170 (N_21170,N_20296,N_20404);
or U21171 (N_21171,N_20502,N_19752);
or U21172 (N_21172,N_20882,N_20573);
or U21173 (N_21173,N_20140,N_19778);
nor U21174 (N_21174,N_20932,N_20457);
nor U21175 (N_21175,N_20878,N_20117);
or U21176 (N_21176,N_19830,N_20659);
nand U21177 (N_21177,N_19782,N_20958);
nand U21178 (N_21178,N_20256,N_20690);
nand U21179 (N_21179,N_20229,N_20859);
and U21180 (N_21180,N_20265,N_19827);
or U21181 (N_21181,N_20002,N_20600);
nor U21182 (N_21182,N_20456,N_20728);
or U21183 (N_21183,N_19726,N_20325);
xnor U21184 (N_21184,N_20266,N_20771);
or U21185 (N_21185,N_19967,N_19738);
or U21186 (N_21186,N_19788,N_20009);
and U21187 (N_21187,N_20409,N_20241);
xor U21188 (N_21188,N_20348,N_19640);
nor U21189 (N_21189,N_19771,N_20913);
nor U21190 (N_21190,N_20309,N_19842);
nand U21191 (N_21191,N_19914,N_20224);
or U21192 (N_21192,N_20308,N_19926);
xnor U21193 (N_21193,N_20686,N_19620);
xnor U21194 (N_21194,N_20635,N_20159);
and U21195 (N_21195,N_20578,N_20144);
xnor U21196 (N_21196,N_20906,N_19889);
and U21197 (N_21197,N_19548,N_20673);
nand U21198 (N_21198,N_20483,N_19737);
or U21199 (N_21199,N_20679,N_19517);
nand U21200 (N_21200,N_19988,N_20849);
or U21201 (N_21201,N_20698,N_20407);
nand U21202 (N_21202,N_20281,N_19992);
xnor U21203 (N_21203,N_20305,N_19971);
or U21204 (N_21204,N_20124,N_20615);
and U21205 (N_21205,N_20223,N_20482);
and U21206 (N_21206,N_20118,N_20757);
nor U21207 (N_21207,N_19891,N_20535);
or U21208 (N_21208,N_19956,N_20991);
nand U21209 (N_21209,N_20424,N_19649);
and U21210 (N_21210,N_20726,N_20036);
and U21211 (N_21211,N_19754,N_20755);
nand U21212 (N_21212,N_19826,N_20511);
xnor U21213 (N_21213,N_19949,N_20391);
and U21214 (N_21214,N_20961,N_19590);
xor U21215 (N_21215,N_20639,N_20912);
xor U21216 (N_21216,N_20970,N_19791);
xor U21217 (N_21217,N_20915,N_20521);
xor U21218 (N_21218,N_20983,N_20838);
and U21219 (N_21219,N_20819,N_20164);
nand U21220 (N_21220,N_20102,N_19655);
xor U21221 (N_21221,N_20972,N_20328);
nand U21222 (N_21222,N_20274,N_20998);
nor U21223 (N_21223,N_19808,N_19862);
xnor U21224 (N_21224,N_20792,N_20290);
nand U21225 (N_21225,N_19689,N_20103);
xnor U21226 (N_21226,N_20155,N_19762);
and U21227 (N_21227,N_20692,N_20494);
nor U21228 (N_21228,N_20737,N_19510);
nand U21229 (N_21229,N_20560,N_20369);
nand U21230 (N_21230,N_20273,N_20152);
nor U21231 (N_21231,N_19903,N_19796);
nor U21232 (N_21232,N_20662,N_20148);
or U21233 (N_21233,N_19943,N_20888);
nand U21234 (N_21234,N_19509,N_19831);
xnor U21235 (N_21235,N_19768,N_20130);
or U21236 (N_21236,N_19803,N_20979);
or U21237 (N_21237,N_20937,N_19800);
nor U21238 (N_21238,N_20848,N_19718);
xor U21239 (N_21239,N_20492,N_20701);
or U21240 (N_21240,N_20641,N_20605);
nor U21241 (N_21241,N_20952,N_20446);
xor U21242 (N_21242,N_19512,N_20593);
nor U21243 (N_21243,N_20068,N_20963);
or U21244 (N_21244,N_20194,N_20777);
nand U21245 (N_21245,N_19608,N_19678);
and U21246 (N_21246,N_20368,N_20640);
nor U21247 (N_21247,N_20924,N_19935);
and U21248 (N_21248,N_20294,N_20478);
xor U21249 (N_21249,N_19518,N_19784);
and U21250 (N_21250,N_19805,N_19650);
xor U21251 (N_21251,N_19639,N_20170);
nor U21252 (N_21252,N_19698,N_19597);
and U21253 (N_21253,N_20966,N_19702);
xnor U21254 (N_21254,N_20897,N_20345);
nand U21255 (N_21255,N_20835,N_20729);
and U21256 (N_21256,N_20333,N_20042);
nand U21257 (N_21257,N_19641,N_20606);
or U21258 (N_21258,N_20195,N_19897);
nor U21259 (N_21259,N_20682,N_20530);
or U21260 (N_21260,N_20097,N_20652);
xor U21261 (N_21261,N_19665,N_19600);
and U21262 (N_21262,N_19723,N_19662);
and U21263 (N_21263,N_19982,N_20110);
xor U21264 (N_21264,N_19915,N_20012);
nor U21265 (N_21265,N_20079,N_19633);
xnor U21266 (N_21266,N_20693,N_19930);
xor U21267 (N_21267,N_20257,N_19570);
and U21268 (N_21268,N_20810,N_20571);
or U21269 (N_21269,N_20358,N_19984);
nand U21270 (N_21270,N_20561,N_20750);
nand U21271 (N_21271,N_20900,N_20284);
or U21272 (N_21272,N_20663,N_19931);
xnor U21273 (N_21273,N_20548,N_20556);
xor U21274 (N_21274,N_20748,N_20344);
nand U21275 (N_21275,N_20540,N_19564);
nor U21276 (N_21276,N_20088,N_20942);
nor U21277 (N_21277,N_20854,N_19699);
or U21278 (N_21278,N_20666,N_20360);
xnor U21279 (N_21279,N_19923,N_19544);
or U21280 (N_21280,N_19554,N_19676);
nor U21281 (N_21281,N_20204,N_19965);
and U21282 (N_21282,N_19687,N_20609);
nand U21283 (N_21283,N_19656,N_19841);
and U21284 (N_21284,N_20202,N_20052);
nor U21285 (N_21285,N_20054,N_19622);
or U21286 (N_21286,N_20795,N_20251);
nand U21287 (N_21287,N_19905,N_20526);
nand U21288 (N_21288,N_19652,N_20376);
and U21289 (N_21289,N_20860,N_20828);
and U21290 (N_21290,N_19538,N_19884);
and U21291 (N_21291,N_20883,N_19857);
xnor U21292 (N_21292,N_20049,N_19513);
xnor U21293 (N_21293,N_19818,N_19532);
xnor U21294 (N_21294,N_20965,N_20969);
nor U21295 (N_21295,N_19955,N_20538);
nor U21296 (N_21296,N_19552,N_20570);
xor U21297 (N_21297,N_20268,N_20203);
or U21298 (N_21298,N_19638,N_20964);
nand U21299 (N_21299,N_20394,N_20248);
xor U21300 (N_21300,N_20992,N_20261);
or U21301 (N_21301,N_19562,N_20043);
or U21302 (N_21302,N_20313,N_20493);
or U21303 (N_21303,N_20425,N_20161);
or U21304 (N_21304,N_19934,N_20770);
nor U21305 (N_21305,N_20173,N_20818);
and U21306 (N_21306,N_20703,N_20769);
nand U21307 (N_21307,N_20585,N_20464);
or U21308 (N_21308,N_20234,N_20612);
or U21309 (N_21309,N_20417,N_20776);
and U21310 (N_21310,N_20291,N_20773);
xor U21311 (N_21311,N_19626,N_20542);
xnor U21312 (N_21312,N_19871,N_20629);
nor U21313 (N_21313,N_20349,N_20967);
xor U21314 (N_21314,N_19690,N_19602);
xor U21315 (N_21315,N_20681,N_20832);
xor U21316 (N_21316,N_20059,N_19609);
nand U21317 (N_21317,N_20714,N_20877);
xnor U21318 (N_21318,N_20765,N_19706);
nand U21319 (N_21319,N_20827,N_19536);
xor U21320 (N_21320,N_20699,N_20070);
and U21321 (N_21321,N_20338,N_20318);
xor U21322 (N_21322,N_19716,N_19806);
or U21323 (N_21323,N_20718,N_20797);
or U21324 (N_21324,N_20374,N_20053);
nor U21325 (N_21325,N_20667,N_19920);
and U21326 (N_21326,N_19836,N_20947);
nor U21327 (N_21327,N_20064,N_20235);
xor U21328 (N_21328,N_20536,N_20398);
or U21329 (N_21329,N_19991,N_20470);
nor U21330 (N_21330,N_20105,N_20311);
nand U21331 (N_21331,N_19987,N_20406);
xor U21332 (N_21332,N_19664,N_19983);
and U21333 (N_21333,N_20938,N_20581);
and U21334 (N_21334,N_20469,N_20423);
nand U21335 (N_21335,N_20803,N_20584);
nand U21336 (N_21336,N_20628,N_20020);
and U21337 (N_21337,N_20712,N_20244);
or U21338 (N_21338,N_19932,N_20249);
or U21339 (N_21339,N_19947,N_20798);
nand U21340 (N_21340,N_19603,N_20267);
xnor U21341 (N_21341,N_20672,N_20449);
and U21342 (N_21342,N_20356,N_20580);
or U21343 (N_21343,N_19907,N_20490);
nand U21344 (N_21344,N_19790,N_20370);
and U21345 (N_21345,N_19972,N_20237);
nor U21346 (N_21346,N_20246,N_20632);
xor U21347 (N_21347,N_20150,N_19917);
nand U21348 (N_21348,N_20793,N_19714);
nor U21349 (N_21349,N_19912,N_20232);
and U21350 (N_21350,N_20003,N_19660);
and U21351 (N_21351,N_19684,N_19894);
or U21352 (N_21352,N_20804,N_19503);
and U21353 (N_21353,N_19960,N_20747);
or U21354 (N_21354,N_20539,N_19730);
or U21355 (N_21355,N_20217,N_19774);
nand U21356 (N_21356,N_20820,N_19763);
and U21357 (N_21357,N_20310,N_19581);
or U21358 (N_21358,N_19601,N_19797);
xor U21359 (N_21359,N_20153,N_20697);
nor U21360 (N_21360,N_20214,N_20351);
xor U21361 (N_21361,N_19502,N_19646);
or U21362 (N_21362,N_20871,N_20352);
and U21363 (N_21363,N_19571,N_20474);
or U21364 (N_21364,N_19733,N_20880);
xnor U21365 (N_21365,N_19612,N_19578);
nand U21366 (N_21366,N_20226,N_20101);
or U21367 (N_21367,N_20190,N_19753);
or U21368 (N_21368,N_20221,N_20128);
nand U21369 (N_21369,N_20987,N_20515);
nor U21370 (N_21370,N_19682,N_19648);
and U21371 (N_21371,N_20744,N_19896);
xnor U21372 (N_21372,N_20191,N_20435);
or U21373 (N_21373,N_20100,N_20024);
nor U21374 (N_21374,N_19720,N_19793);
nand U21375 (N_21375,N_19913,N_20533);
and U21376 (N_21376,N_20920,N_19874);
xnor U21377 (N_21377,N_20324,N_19848);
and U21378 (N_21378,N_20129,N_20431);
or U21379 (N_21379,N_20541,N_19922);
nor U21380 (N_21380,N_20706,N_20711);
nor U21381 (N_21381,N_20846,N_20767);
or U21382 (N_21382,N_20602,N_20171);
or U21383 (N_21383,N_20825,N_20787);
nor U21384 (N_21384,N_19772,N_20413);
or U21385 (N_21385,N_19614,N_19879);
xor U21386 (N_21386,N_19748,N_20162);
and U21387 (N_21387,N_19743,N_19540);
and U21388 (N_21388,N_20160,N_20461);
and U21389 (N_21389,N_20689,N_20389);
nor U21390 (N_21390,N_20000,N_20506);
xor U21391 (N_21391,N_20343,N_20017);
nand U21392 (N_21392,N_19523,N_19901);
nor U21393 (N_21393,N_20876,N_20180);
xor U21394 (N_21394,N_20844,N_19744);
nand U21395 (N_21395,N_20208,N_20231);
and U21396 (N_21396,N_20887,N_20922);
or U21397 (N_21397,N_20157,N_19696);
and U21398 (N_21398,N_19671,N_19514);
or U21399 (N_21399,N_20136,N_20444);
nand U21400 (N_21400,N_19792,N_20372);
nand U21401 (N_21401,N_20396,N_20916);
and U21402 (N_21402,N_20907,N_19594);
xnor U21403 (N_21403,N_20106,N_19520);
nand U21404 (N_21404,N_20497,N_20184);
nor U21405 (N_21405,N_19973,N_19843);
xnor U21406 (N_21406,N_20563,N_20316);
or U21407 (N_21407,N_20625,N_20458);
nand U21408 (N_21408,N_20323,N_20081);
and U21409 (N_21409,N_19724,N_20962);
nand U21410 (N_21410,N_19933,N_20738);
nand U21411 (N_21411,N_20527,N_19995);
nor U21412 (N_21412,N_20277,N_20076);
and U21413 (N_21413,N_19534,N_20732);
xnor U21414 (N_21414,N_19705,N_20275);
and U21415 (N_21415,N_19695,N_20695);
xor U21416 (N_21416,N_19749,N_20442);
or U21417 (N_21417,N_19728,N_20056);
nor U21418 (N_21418,N_19647,N_19756);
or U21419 (N_21419,N_20107,N_19735);
xor U21420 (N_21420,N_20976,N_20986);
xnor U21421 (N_21421,N_20499,N_20761);
nor U21422 (N_21422,N_19643,N_20829);
nand U21423 (N_21423,N_20287,N_19574);
nor U21424 (N_21424,N_20588,N_20143);
nor U21425 (N_21425,N_20720,N_20599);
nand U21426 (N_21426,N_20781,N_20559);
nand U21427 (N_21427,N_19736,N_20505);
xor U21428 (N_21428,N_20412,N_20312);
or U21429 (N_21429,N_20210,N_20095);
or U21430 (N_21430,N_19507,N_20981);
nor U21431 (N_21431,N_20950,N_20138);
nor U21432 (N_21432,N_20428,N_19990);
xnor U21433 (N_21433,N_20688,N_19801);
and U21434 (N_21434,N_19677,N_20577);
nor U21435 (N_21435,N_20365,N_20018);
nor U21436 (N_21436,N_19529,N_20495);
nor U21437 (N_21437,N_20869,N_20219);
and U21438 (N_21438,N_20041,N_19767);
nand U21439 (N_21439,N_20794,N_20397);
nor U21440 (N_21440,N_19668,N_20596);
and U21441 (N_21441,N_20038,N_20512);
and U21442 (N_21442,N_20959,N_20491);
or U21443 (N_21443,N_20035,N_20660);
nor U21444 (N_21444,N_19593,N_20116);
or U21445 (N_21445,N_19918,N_20700);
or U21446 (N_21446,N_20568,N_19908);
and U21447 (N_21447,N_20678,N_20518);
and U21448 (N_21448,N_20260,N_20513);
nand U21449 (N_21449,N_20373,N_19795);
xnor U21450 (N_21450,N_20759,N_20953);
and U21451 (N_21451,N_20200,N_20091);
nor U21452 (N_21452,N_19794,N_20902);
nand U21453 (N_21453,N_20929,N_20022);
xnor U21454 (N_21454,N_20388,N_19875);
or U21455 (N_21455,N_19976,N_20856);
and U21456 (N_21456,N_19712,N_20306);
nand U21457 (N_21457,N_20255,N_20015);
or U21458 (N_21458,N_20341,N_20665);
nor U21459 (N_21459,N_19787,N_20201);
xor U21460 (N_21460,N_19944,N_20176);
or U21461 (N_21461,N_20905,N_20023);
nand U21462 (N_21462,N_20812,N_19527);
or U21463 (N_21463,N_20653,N_20740);
nor U21464 (N_21464,N_19692,N_20598);
and U21465 (N_21465,N_20756,N_20783);
or U21466 (N_21466,N_20252,N_20862);
nand U21467 (N_21467,N_19722,N_20993);
xnor U21468 (N_21468,N_19777,N_19572);
or U21469 (N_21469,N_20243,N_19837);
xnor U21470 (N_21470,N_19599,N_19673);
or U21471 (N_21471,N_20399,N_19809);
nand U21472 (N_21472,N_20259,N_20749);
xnor U21473 (N_21473,N_19598,N_20574);
and U21474 (N_21474,N_20113,N_20034);
nand U21475 (N_21475,N_20304,N_20928);
xnor U21476 (N_21476,N_19927,N_20855);
or U21477 (N_21477,N_19866,N_19898);
xor U21478 (N_21478,N_20498,N_20427);
nor U21479 (N_21479,N_19766,N_20320);
and U21480 (N_21480,N_20451,N_20841);
and U21481 (N_21481,N_20183,N_19881);
nand U21482 (N_21482,N_19567,N_20379);
nand U21483 (N_21483,N_20504,N_20645);
or U21484 (N_21484,N_20286,N_20297);
nor U21485 (N_21485,N_19868,N_20644);
xor U21486 (N_21486,N_20032,N_19755);
nand U21487 (N_21487,N_19653,N_20843);
xnor U21488 (N_21488,N_20946,N_19887);
nand U21489 (N_21489,N_20824,N_19680);
or U21490 (N_21490,N_20746,N_19628);
nor U21491 (N_21491,N_20131,N_19872);
and U21492 (N_21492,N_20802,N_20030);
nor U21493 (N_21493,N_20317,N_20227);
nand U21494 (N_21494,N_20156,N_20347);
or U21495 (N_21495,N_20800,N_19501);
or U21496 (N_21496,N_20719,N_20099);
nand U21497 (N_21497,N_20279,N_19747);
nand U21498 (N_21498,N_20901,N_20613);
or U21499 (N_21499,N_20433,N_20847);
nand U21500 (N_21500,N_19679,N_19751);
nor U21501 (N_21501,N_20973,N_20187);
or U21502 (N_21502,N_19852,N_19623);
and U21503 (N_21503,N_20421,N_20634);
nand U21504 (N_21504,N_20247,N_20687);
nand U21505 (N_21505,N_20484,N_20013);
or U21506 (N_21506,N_19663,N_20151);
or U21507 (N_21507,N_20182,N_20326);
nand U21508 (N_21508,N_19816,N_19686);
xor U21509 (N_21509,N_20935,N_20141);
xnor U21510 (N_21510,N_20760,N_20033);
or U21511 (N_21511,N_20826,N_19892);
xor U21512 (N_21512,N_20707,N_19719);
nand U21513 (N_21513,N_19925,N_20114);
nor U21514 (N_21514,N_19899,N_20957);
xnor U21515 (N_21515,N_20302,N_20557);
nand U21516 (N_21516,N_20299,N_19508);
nand U21517 (N_21517,N_19693,N_20716);
xor U21518 (N_21518,N_20941,N_19966);
xnor U21519 (N_21519,N_19832,N_19835);
xnor U21520 (N_21520,N_19558,N_19729);
nand U21521 (N_21521,N_20475,N_19900);
nor U21522 (N_21522,N_20158,N_20416);
and U21523 (N_21523,N_19632,N_19709);
nand U21524 (N_21524,N_20930,N_19968);
and U21525 (N_21525,N_20185,N_20567);
nand U21526 (N_21526,N_20405,N_20300);
xor U21527 (N_21527,N_19577,N_20566);
and U21528 (N_21528,N_20664,N_20334);
or U21529 (N_21529,N_20438,N_20460);
xor U21530 (N_21530,N_19658,N_20951);
and U21531 (N_21531,N_20496,N_20112);
nor U21532 (N_21532,N_19539,N_20292);
and U21533 (N_21533,N_20418,N_20385);
xnor U21534 (N_21534,N_19659,N_20646);
nor U21535 (N_21535,N_20298,N_20430);
and U21536 (N_21536,N_20807,N_19621);
nor U21537 (N_21537,N_19878,N_19576);
nand U21538 (N_21538,N_19654,N_20093);
nor U21539 (N_21539,N_19817,N_19959);
or U21540 (N_21540,N_20355,N_20480);
nor U21541 (N_21541,N_20471,N_19575);
nand U21542 (N_21542,N_19781,N_20359);
xor U21543 (N_21543,N_20383,N_20842);
nand U21544 (N_21544,N_19708,N_19511);
xnor U21545 (N_21545,N_20845,N_19561);
or U21546 (N_21546,N_19877,N_19535);
and U21547 (N_21547,N_20943,N_20622);
and U21548 (N_21548,N_20546,N_20908);
nand U21549 (N_21549,N_19845,N_20481);
nor U21550 (N_21550,N_20649,N_20791);
xnor U21551 (N_21551,N_20873,N_20501);
xor U21552 (N_21552,N_20211,N_20263);
nor U21553 (N_21553,N_20096,N_19582);
nand U21554 (N_21554,N_20670,N_19592);
and U21555 (N_21555,N_20931,N_20293);
nand U21556 (N_21556,N_20134,N_20683);
nand U21557 (N_21557,N_19828,N_20062);
xor U21558 (N_21558,N_20303,N_19619);
nor U21559 (N_21559,N_20378,N_20801);
xnor U21560 (N_21560,N_19607,N_20875);
xor U21561 (N_21561,N_19780,N_20668);
nand U21562 (N_21562,N_19715,N_20636);
and U21563 (N_21563,N_20569,N_20661);
nor U21564 (N_21564,N_20899,N_19938);
or U21565 (N_21565,N_20285,N_20549);
nor U21566 (N_21566,N_20055,N_20960);
nor U21567 (N_21567,N_20206,N_20840);
nand U21568 (N_21568,N_19560,N_19909);
nand U21569 (N_21569,N_20467,N_20796);
nand U21570 (N_21570,N_19775,N_20813);
and U21571 (N_21571,N_20554,N_20314);
nand U21572 (N_21572,N_20582,N_20228);
nand U21573 (N_21573,N_20893,N_20339);
and U21574 (N_21574,N_20080,N_20597);
or U21575 (N_21575,N_20058,N_19929);
or U21576 (N_21576,N_20619,N_20078);
and U21577 (N_21577,N_20166,N_20209);
or U21578 (N_21578,N_20858,N_20785);
xnor U21579 (N_21579,N_19858,N_19840);
xnor U21580 (N_21580,N_19910,N_20784);
nand U21581 (N_21581,N_20975,N_20657);
and U21582 (N_21582,N_20019,N_20434);
xor U21583 (N_21583,N_20999,N_20330);
nand U21584 (N_21584,N_20717,N_20620);
and U21585 (N_21585,N_20734,N_20704);
and U21586 (N_21586,N_20236,N_20196);
xor U21587 (N_21587,N_20626,N_19882);
and U21588 (N_21588,N_20575,N_20715);
nand U21589 (N_21589,N_20779,N_19516);
nor U21590 (N_21590,N_20739,N_20621);
nor U21591 (N_21591,N_19985,N_20917);
xnor U21592 (N_21592,N_19789,N_20774);
or U21593 (N_21593,N_19522,N_20319);
and U21594 (N_21594,N_20218,N_20524);
and U21595 (N_21595,N_20696,N_20508);
nor U21596 (N_21596,N_19746,N_20215);
xor U21597 (N_21597,N_20821,N_20485);
nand U21598 (N_21598,N_20586,N_20616);
nand U21599 (N_21599,N_20327,N_20402);
and U21600 (N_21600,N_20282,N_19636);
and U21601 (N_21601,N_20395,N_20617);
or U21602 (N_21602,N_20919,N_19822);
nor U21603 (N_21603,N_19727,N_20050);
xnor U21604 (N_21604,N_20381,N_20623);
and U21605 (N_21605,N_20866,N_19530);
and U21606 (N_21606,N_20654,N_20543);
nand U21607 (N_21607,N_19667,N_20077);
nand U21608 (N_21608,N_20918,N_20230);
xnor U21609 (N_21609,N_20239,N_20531);
nand U21610 (N_21610,N_19635,N_19742);
xnor U21611 (N_21611,N_20008,N_20169);
or U21612 (N_21612,N_20098,N_19769);
and U21613 (N_21613,N_20045,N_20065);
nand U21614 (N_21614,N_19596,N_19613);
xnor U21615 (N_21615,N_19855,N_19580);
nor U21616 (N_21616,N_20175,N_20830);
or U21617 (N_21617,N_20564,N_20944);
nand U21618 (N_21618,N_19833,N_20850);
nor U21619 (N_21619,N_19849,N_20066);
or U21620 (N_21620,N_20529,N_20806);
nand U21621 (N_21621,N_20684,N_19911);
nor U21622 (N_21622,N_19970,N_19954);
nor U21623 (N_21623,N_20010,N_19583);
or U21624 (N_21624,N_20519,N_19694);
xor U21625 (N_21625,N_20139,N_19579);
nand U21626 (N_21626,N_19624,N_20894);
nand U21627 (N_21627,N_19993,N_20477);
or U21628 (N_21628,N_19605,N_19974);
nand U21629 (N_21629,N_19981,N_19936);
xor U21630 (N_21630,N_19505,N_19642);
nand U21631 (N_21631,N_19515,N_20708);
xor U21632 (N_21632,N_19566,N_19559);
or U21633 (N_21633,N_20337,N_19779);
or U21634 (N_21634,N_19856,N_20753);
xnor U21635 (N_21635,N_20927,N_20604);
xor U21636 (N_21636,N_20786,N_19921);
nor U21637 (N_21637,N_19810,N_20459);
or U21638 (N_21638,N_20565,N_19961);
and U21639 (N_21639,N_19945,N_19625);
or U21640 (N_21640,N_19989,N_20380);
nand U21641 (N_21641,N_19975,N_20775);
and U21642 (N_21642,N_20735,N_19829);
nand U21643 (N_21643,N_19524,N_19812);
and U21644 (N_21644,N_20089,N_20126);
nand U21645 (N_21645,N_20220,N_20815);
nand U21646 (N_21646,N_20782,N_19820);
or U21647 (N_21647,N_20288,N_20892);
nand U21648 (N_21648,N_19750,N_20415);
and U21649 (N_21649,N_20057,N_19586);
or U21650 (N_21650,N_20736,N_20410);
and U21651 (N_21651,N_20611,N_20550);
nand U21652 (N_21652,N_20177,N_20122);
xnor U21653 (N_21653,N_19869,N_20627);
xnor U21654 (N_21654,N_20558,N_19813);
xnor U21655 (N_21655,N_19761,N_20426);
or U21656 (N_21656,N_19568,N_19867);
and U21657 (N_21657,N_19685,N_19697);
or U21658 (N_21658,N_20198,N_19519);
or U21659 (N_21659,N_20865,N_19674);
nor U21660 (N_21660,N_19711,N_20001);
or U21661 (N_21661,N_20572,N_20934);
nand U21662 (N_21662,N_20839,N_20479);
nand U21663 (N_21663,N_20362,N_20743);
nand U21664 (N_21664,N_20007,N_20741);
nand U21665 (N_21665,N_20691,N_20272);
nor U21666 (N_21666,N_19825,N_20205);
and U21667 (N_21667,N_20238,N_20528);
nor U21668 (N_21668,N_19617,N_20307);
and U21669 (N_21669,N_19939,N_20669);
nand U21670 (N_21670,N_20084,N_20601);
and U21671 (N_21671,N_20650,N_19937);
nor U21672 (N_21672,N_20245,N_19525);
and U21673 (N_21673,N_20724,N_20607);
or U21674 (N_21674,N_19556,N_20011);
or U21675 (N_21675,N_20603,N_19998);
xor U21676 (N_21676,N_20075,N_19526);
xnor U21677 (N_21677,N_20655,N_20658);
and U21678 (N_21678,N_20167,N_20363);
and U21679 (N_21679,N_20336,N_19585);
xor U21680 (N_21680,N_19798,N_20109);
xor U21681 (N_21681,N_20121,N_19713);
and U21682 (N_21682,N_19573,N_20354);
nor U21683 (N_21683,N_19657,N_20069);
and U21684 (N_21684,N_20197,N_20213);
nor U21685 (N_21685,N_20886,N_20147);
nand U21686 (N_21686,N_19675,N_19953);
and U21687 (N_21687,N_20772,N_20940);
or U21688 (N_21688,N_20643,N_20852);
nor U21689 (N_21689,N_20455,N_20462);
or U21690 (N_21690,N_20283,N_20671);
nor U21691 (N_21691,N_20864,N_20933);
or U21692 (N_21692,N_20988,N_19824);
xnor U21693 (N_21693,N_20414,N_20870);
xnor U21694 (N_21694,N_20125,N_20135);
or U21695 (N_21695,N_20500,N_20680);
or U21696 (N_21696,N_20949,N_20778);
nand U21697 (N_21697,N_19569,N_19819);
xnor U21698 (N_21698,N_20111,N_20212);
and U21699 (N_21699,N_19551,N_20956);
nand U21700 (N_21700,N_20253,N_20027);
nor U21701 (N_21701,N_19616,N_19543);
xnor U21702 (N_21702,N_20751,N_20836);
xor U21703 (N_21703,N_20242,N_20710);
xnor U21704 (N_21704,N_20630,N_20816);
or U21705 (N_21705,N_20590,N_20453);
nand U21706 (N_21706,N_20525,N_20898);
nor U21707 (N_21707,N_20387,N_19637);
or U21708 (N_21708,N_20072,N_19854);
or U21709 (N_21709,N_20445,N_20108);
or U21710 (N_21710,N_20911,N_20465);
nor U21711 (N_21711,N_19999,N_19885);
nor U21712 (N_21712,N_20909,N_19890);
or U21713 (N_21713,N_19610,N_20487);
xor U21714 (N_21714,N_20429,N_19942);
xnor U21715 (N_21715,N_20788,N_20436);
xor U21716 (N_21716,N_19618,N_19814);
and U21717 (N_21717,N_19799,N_20040);
or U21718 (N_21718,N_19725,N_19669);
and U21719 (N_21719,N_20258,N_20074);
nand U21720 (N_21720,N_20874,N_19904);
or U21721 (N_21721,N_19651,N_20189);
nand U21722 (N_21722,N_20067,N_19528);
or U21723 (N_21723,N_20890,N_19546);
xnor U21724 (N_21724,N_20085,N_20587);
xnor U21725 (N_21725,N_20914,N_19588);
or U21726 (N_21726,N_20833,N_20454);
nor U21727 (N_21727,N_20335,N_20400);
nor U21728 (N_21728,N_19759,N_20923);
nor U21729 (N_21729,N_20082,N_20186);
xor U21730 (N_21730,N_20163,N_20579);
nor U21731 (N_21731,N_20638,N_20675);
nor U21732 (N_21732,N_19688,N_20814);
nor U21733 (N_21733,N_20853,N_20884);
nand U21734 (N_21734,N_20403,N_20997);
nor U21735 (N_21735,N_20790,N_20278);
or U21736 (N_21736,N_20037,N_19962);
nand U21737 (N_21737,N_20651,N_19924);
xor U21738 (N_21738,N_20149,N_20984);
xnor U21739 (N_21739,N_20990,N_20145);
nor U21740 (N_21740,N_19895,N_20174);
or U21741 (N_21741,N_20766,N_20443);
nand U21742 (N_21742,N_19958,N_20254);
nor U21743 (N_21743,N_19615,N_20386);
and U21744 (N_21744,N_20005,N_20503);
or U21745 (N_21745,N_20322,N_19893);
xor U21746 (N_21746,N_19555,N_20995);
nor U21747 (N_21747,N_20758,N_19565);
and U21748 (N_21748,N_19672,N_20489);
or U21749 (N_21749,N_20896,N_19786);
nor U21750 (N_21750,N_19880,N_20300);
nor U21751 (N_21751,N_20924,N_19654);
nand U21752 (N_21752,N_20112,N_20600);
or U21753 (N_21753,N_20928,N_20349);
or U21754 (N_21754,N_20728,N_19695);
nor U21755 (N_21755,N_19881,N_20879);
nand U21756 (N_21756,N_20654,N_20567);
or U21757 (N_21757,N_20540,N_20377);
xor U21758 (N_21758,N_19857,N_19711);
xor U21759 (N_21759,N_19879,N_20858);
nand U21760 (N_21760,N_20760,N_20620);
xor U21761 (N_21761,N_20198,N_19914);
nand U21762 (N_21762,N_19714,N_19535);
and U21763 (N_21763,N_20343,N_20236);
or U21764 (N_21764,N_20995,N_19963);
and U21765 (N_21765,N_20118,N_20311);
nand U21766 (N_21766,N_20891,N_19773);
and U21767 (N_21767,N_19969,N_20028);
xor U21768 (N_21768,N_20961,N_20627);
nand U21769 (N_21769,N_20271,N_19931);
xnor U21770 (N_21770,N_20043,N_19948);
nand U21771 (N_21771,N_20937,N_20507);
nor U21772 (N_21772,N_20860,N_19873);
or U21773 (N_21773,N_20596,N_20912);
xnor U21774 (N_21774,N_20432,N_20079);
or U21775 (N_21775,N_20779,N_19827);
nand U21776 (N_21776,N_20231,N_20369);
nor U21777 (N_21777,N_20855,N_20329);
nor U21778 (N_21778,N_20207,N_19917);
xor U21779 (N_21779,N_19908,N_20979);
and U21780 (N_21780,N_20103,N_19805);
xnor U21781 (N_21781,N_20901,N_20786);
xor U21782 (N_21782,N_20441,N_20512);
xnor U21783 (N_21783,N_19879,N_20330);
nand U21784 (N_21784,N_19727,N_19675);
or U21785 (N_21785,N_19834,N_20681);
and U21786 (N_21786,N_20439,N_20429);
nand U21787 (N_21787,N_19861,N_20594);
nand U21788 (N_21788,N_19568,N_20891);
nor U21789 (N_21789,N_20519,N_20199);
or U21790 (N_21790,N_20028,N_20819);
xor U21791 (N_21791,N_20643,N_20921);
or U21792 (N_21792,N_19895,N_20148);
nand U21793 (N_21793,N_19781,N_19752);
and U21794 (N_21794,N_20372,N_20934);
and U21795 (N_21795,N_19740,N_19933);
nand U21796 (N_21796,N_20279,N_20640);
xnor U21797 (N_21797,N_20574,N_20817);
or U21798 (N_21798,N_20402,N_19878);
nand U21799 (N_21799,N_19925,N_20345);
nand U21800 (N_21800,N_20879,N_20121);
and U21801 (N_21801,N_20594,N_20575);
or U21802 (N_21802,N_20261,N_20043);
nand U21803 (N_21803,N_20197,N_20462);
nor U21804 (N_21804,N_20661,N_20431);
and U21805 (N_21805,N_19584,N_20056);
xor U21806 (N_21806,N_19939,N_20619);
or U21807 (N_21807,N_20615,N_20149);
or U21808 (N_21808,N_20025,N_20051);
xnor U21809 (N_21809,N_19682,N_19533);
or U21810 (N_21810,N_20542,N_19900);
nand U21811 (N_21811,N_19948,N_19558);
nor U21812 (N_21812,N_20819,N_20444);
or U21813 (N_21813,N_20928,N_19788);
nor U21814 (N_21814,N_20837,N_20759);
xor U21815 (N_21815,N_20487,N_20581);
xor U21816 (N_21816,N_20083,N_19929);
nand U21817 (N_21817,N_20622,N_19544);
nand U21818 (N_21818,N_20969,N_20020);
xor U21819 (N_21819,N_19766,N_20398);
nor U21820 (N_21820,N_20537,N_20825);
or U21821 (N_21821,N_19787,N_20047);
xor U21822 (N_21822,N_20522,N_20785);
or U21823 (N_21823,N_20103,N_20951);
and U21824 (N_21824,N_20663,N_19750);
and U21825 (N_21825,N_19622,N_20519);
xnor U21826 (N_21826,N_20288,N_19668);
nand U21827 (N_21827,N_19864,N_20167);
and U21828 (N_21828,N_19596,N_20978);
or U21829 (N_21829,N_19829,N_20448);
or U21830 (N_21830,N_20160,N_19556);
xor U21831 (N_21831,N_20218,N_20917);
and U21832 (N_21832,N_20480,N_19533);
or U21833 (N_21833,N_19559,N_19815);
or U21834 (N_21834,N_20453,N_19858);
nor U21835 (N_21835,N_20869,N_19882);
and U21836 (N_21836,N_19672,N_20008);
nand U21837 (N_21837,N_19812,N_20725);
xnor U21838 (N_21838,N_19574,N_19535);
or U21839 (N_21839,N_20487,N_19703);
or U21840 (N_21840,N_20665,N_19865);
xor U21841 (N_21841,N_19872,N_19530);
and U21842 (N_21842,N_20834,N_20765);
and U21843 (N_21843,N_20759,N_19959);
nor U21844 (N_21844,N_20493,N_20511);
xor U21845 (N_21845,N_19751,N_19726);
and U21846 (N_21846,N_19833,N_19828);
nand U21847 (N_21847,N_19851,N_20047);
xor U21848 (N_21848,N_20581,N_20630);
nand U21849 (N_21849,N_19703,N_19959);
nor U21850 (N_21850,N_20928,N_20321);
xor U21851 (N_21851,N_20340,N_20031);
nor U21852 (N_21852,N_20994,N_20497);
xor U21853 (N_21853,N_20624,N_20819);
nand U21854 (N_21854,N_20914,N_20648);
nand U21855 (N_21855,N_20967,N_20440);
and U21856 (N_21856,N_20149,N_19590);
nor U21857 (N_21857,N_19935,N_20396);
nand U21858 (N_21858,N_20494,N_19578);
and U21859 (N_21859,N_20848,N_19933);
and U21860 (N_21860,N_19569,N_20980);
nand U21861 (N_21861,N_19633,N_20240);
nor U21862 (N_21862,N_20536,N_19775);
or U21863 (N_21863,N_20923,N_20807);
nor U21864 (N_21864,N_20373,N_20863);
xor U21865 (N_21865,N_20546,N_19527);
xnor U21866 (N_21866,N_19891,N_20592);
nor U21867 (N_21867,N_20935,N_19742);
and U21868 (N_21868,N_20228,N_19971);
xor U21869 (N_21869,N_20076,N_19518);
nand U21870 (N_21870,N_19583,N_20711);
or U21871 (N_21871,N_20858,N_20543);
and U21872 (N_21872,N_19706,N_19655);
or U21873 (N_21873,N_19586,N_20558);
xor U21874 (N_21874,N_20488,N_20174);
xnor U21875 (N_21875,N_20937,N_20659);
and U21876 (N_21876,N_20608,N_19870);
nand U21877 (N_21877,N_20204,N_20685);
xor U21878 (N_21878,N_19935,N_20516);
nor U21879 (N_21879,N_20447,N_20079);
and U21880 (N_21880,N_19520,N_20977);
or U21881 (N_21881,N_19591,N_19788);
or U21882 (N_21882,N_20863,N_20626);
nand U21883 (N_21883,N_20160,N_20513);
nor U21884 (N_21884,N_19789,N_19577);
nand U21885 (N_21885,N_20087,N_19815);
and U21886 (N_21886,N_19700,N_19659);
nor U21887 (N_21887,N_20507,N_19956);
xor U21888 (N_21888,N_19916,N_20021);
nand U21889 (N_21889,N_19532,N_20834);
nor U21890 (N_21890,N_19636,N_19644);
nor U21891 (N_21891,N_20490,N_20209);
or U21892 (N_21892,N_20239,N_20548);
or U21893 (N_21893,N_20571,N_20242);
xnor U21894 (N_21894,N_20110,N_19570);
and U21895 (N_21895,N_20116,N_19778);
xor U21896 (N_21896,N_20896,N_20061);
nor U21897 (N_21897,N_19804,N_20715);
xor U21898 (N_21898,N_20720,N_19709);
nor U21899 (N_21899,N_20179,N_19830);
nand U21900 (N_21900,N_20811,N_19713);
and U21901 (N_21901,N_19936,N_20360);
or U21902 (N_21902,N_20534,N_20280);
or U21903 (N_21903,N_20829,N_19564);
and U21904 (N_21904,N_20200,N_20310);
or U21905 (N_21905,N_20659,N_19529);
or U21906 (N_21906,N_20140,N_19513);
nor U21907 (N_21907,N_20426,N_19565);
or U21908 (N_21908,N_20519,N_20546);
and U21909 (N_21909,N_19556,N_20130);
nor U21910 (N_21910,N_20390,N_20196);
nor U21911 (N_21911,N_19618,N_20205);
xnor U21912 (N_21912,N_20167,N_20676);
xor U21913 (N_21913,N_19665,N_20255);
nand U21914 (N_21914,N_20175,N_20338);
or U21915 (N_21915,N_20183,N_20137);
xor U21916 (N_21916,N_20080,N_19814);
nor U21917 (N_21917,N_19916,N_20647);
nor U21918 (N_21918,N_20481,N_20366);
nor U21919 (N_21919,N_19751,N_20204);
and U21920 (N_21920,N_20448,N_20687);
or U21921 (N_21921,N_19867,N_20655);
and U21922 (N_21922,N_20424,N_20984);
or U21923 (N_21923,N_19545,N_20404);
xnor U21924 (N_21924,N_20516,N_20923);
nand U21925 (N_21925,N_19509,N_20266);
nor U21926 (N_21926,N_19888,N_20012);
or U21927 (N_21927,N_20496,N_19967);
and U21928 (N_21928,N_20167,N_20646);
or U21929 (N_21929,N_20792,N_20278);
nor U21930 (N_21930,N_20636,N_20346);
nor U21931 (N_21931,N_19743,N_20086);
xor U21932 (N_21932,N_20083,N_19945);
nand U21933 (N_21933,N_19762,N_20186);
or U21934 (N_21934,N_20188,N_19609);
xnor U21935 (N_21935,N_20428,N_19705);
or U21936 (N_21936,N_20499,N_20220);
nor U21937 (N_21937,N_20005,N_19849);
and U21938 (N_21938,N_20662,N_19990);
and U21939 (N_21939,N_20572,N_19995);
nand U21940 (N_21940,N_19580,N_20030);
nor U21941 (N_21941,N_20349,N_20180);
xnor U21942 (N_21942,N_20901,N_19658);
nand U21943 (N_21943,N_20312,N_19928);
or U21944 (N_21944,N_20074,N_19622);
nor U21945 (N_21945,N_19992,N_20667);
xor U21946 (N_21946,N_20694,N_19933);
and U21947 (N_21947,N_20768,N_19822);
xnor U21948 (N_21948,N_20245,N_19848);
xor U21949 (N_21949,N_20942,N_20565);
or U21950 (N_21950,N_20461,N_19884);
nand U21951 (N_21951,N_20277,N_20931);
or U21952 (N_21952,N_19874,N_19833);
xnor U21953 (N_21953,N_19623,N_19813);
nor U21954 (N_21954,N_20181,N_19733);
nor U21955 (N_21955,N_19581,N_20789);
or U21956 (N_21956,N_20984,N_19868);
xor U21957 (N_21957,N_19871,N_19600);
nand U21958 (N_21958,N_20767,N_20581);
and U21959 (N_21959,N_19575,N_20078);
or U21960 (N_21960,N_19630,N_20245);
xor U21961 (N_21961,N_20340,N_20819);
nand U21962 (N_21962,N_19976,N_20056);
and U21963 (N_21963,N_20976,N_20330);
and U21964 (N_21964,N_19580,N_19517);
or U21965 (N_21965,N_19816,N_20296);
or U21966 (N_21966,N_20558,N_20427);
and U21967 (N_21967,N_20257,N_19709);
nor U21968 (N_21968,N_20701,N_20217);
and U21969 (N_21969,N_20247,N_20136);
or U21970 (N_21970,N_20297,N_20178);
nor U21971 (N_21971,N_19508,N_20975);
or U21972 (N_21972,N_20782,N_19633);
nor U21973 (N_21973,N_20651,N_19650);
xor U21974 (N_21974,N_20331,N_19597);
nand U21975 (N_21975,N_20743,N_20675);
or U21976 (N_21976,N_20254,N_20438);
nor U21977 (N_21977,N_20505,N_20611);
xnor U21978 (N_21978,N_20078,N_19849);
nor U21979 (N_21979,N_20286,N_20247);
and U21980 (N_21980,N_20155,N_19505);
xor U21981 (N_21981,N_19677,N_19826);
nor U21982 (N_21982,N_19873,N_19699);
or U21983 (N_21983,N_20052,N_19596);
or U21984 (N_21984,N_20443,N_19549);
nand U21985 (N_21985,N_20509,N_20966);
xor U21986 (N_21986,N_20220,N_19830);
xnor U21987 (N_21987,N_20395,N_20443);
and U21988 (N_21988,N_20951,N_19925);
xor U21989 (N_21989,N_20525,N_20682);
xnor U21990 (N_21990,N_20247,N_20540);
nand U21991 (N_21991,N_20402,N_20877);
or U21992 (N_21992,N_20296,N_19998);
and U21993 (N_21993,N_20270,N_20009);
nor U21994 (N_21994,N_19747,N_20822);
nor U21995 (N_21995,N_20608,N_19578);
nand U21996 (N_21996,N_20497,N_19646);
xor U21997 (N_21997,N_20056,N_19527);
nor U21998 (N_21998,N_19755,N_19712);
nor U21999 (N_21999,N_19638,N_19868);
or U22000 (N_22000,N_19650,N_19671);
and U22001 (N_22001,N_19966,N_20806);
or U22002 (N_22002,N_20745,N_19840);
nand U22003 (N_22003,N_20956,N_20833);
and U22004 (N_22004,N_20566,N_20256);
xnor U22005 (N_22005,N_20164,N_20680);
nand U22006 (N_22006,N_20971,N_19690);
or U22007 (N_22007,N_19598,N_20024);
or U22008 (N_22008,N_20420,N_20072);
nor U22009 (N_22009,N_19868,N_19771);
xor U22010 (N_22010,N_20681,N_19685);
or U22011 (N_22011,N_20863,N_20455);
or U22012 (N_22012,N_19724,N_20361);
or U22013 (N_22013,N_19990,N_20912);
xor U22014 (N_22014,N_19935,N_19962);
xnor U22015 (N_22015,N_19969,N_20182);
xnor U22016 (N_22016,N_19709,N_20988);
xor U22017 (N_22017,N_19624,N_19509);
nand U22018 (N_22018,N_20444,N_20555);
nand U22019 (N_22019,N_20626,N_19907);
and U22020 (N_22020,N_20459,N_19627);
or U22021 (N_22021,N_19683,N_19617);
or U22022 (N_22022,N_19621,N_20814);
xor U22023 (N_22023,N_19758,N_19693);
nor U22024 (N_22024,N_20964,N_20019);
or U22025 (N_22025,N_20608,N_20452);
nand U22026 (N_22026,N_20859,N_20005);
nand U22027 (N_22027,N_20507,N_20975);
nand U22028 (N_22028,N_20814,N_20889);
or U22029 (N_22029,N_20392,N_19525);
nand U22030 (N_22030,N_20180,N_19993);
nand U22031 (N_22031,N_19742,N_20442);
xnor U22032 (N_22032,N_20268,N_20365);
and U22033 (N_22033,N_20753,N_19784);
xnor U22034 (N_22034,N_20100,N_20026);
nand U22035 (N_22035,N_19509,N_20078);
and U22036 (N_22036,N_19514,N_20704);
nand U22037 (N_22037,N_20044,N_20211);
nor U22038 (N_22038,N_20381,N_20966);
nand U22039 (N_22039,N_20860,N_19572);
and U22040 (N_22040,N_20058,N_20175);
nor U22041 (N_22041,N_19712,N_20209);
and U22042 (N_22042,N_20556,N_20824);
and U22043 (N_22043,N_20010,N_20830);
or U22044 (N_22044,N_20000,N_19883);
nand U22045 (N_22045,N_19824,N_20706);
nor U22046 (N_22046,N_20905,N_20923);
nand U22047 (N_22047,N_20316,N_19946);
nand U22048 (N_22048,N_19531,N_19564);
nor U22049 (N_22049,N_20621,N_19585);
or U22050 (N_22050,N_20718,N_19712);
nor U22051 (N_22051,N_20700,N_20573);
or U22052 (N_22052,N_20603,N_20407);
and U22053 (N_22053,N_20361,N_20510);
xor U22054 (N_22054,N_20567,N_20424);
and U22055 (N_22055,N_19933,N_20349);
xnor U22056 (N_22056,N_20467,N_19579);
nor U22057 (N_22057,N_19902,N_20601);
xnor U22058 (N_22058,N_20722,N_19832);
and U22059 (N_22059,N_20273,N_20485);
nand U22060 (N_22060,N_20962,N_19503);
nor U22061 (N_22061,N_20373,N_19740);
nor U22062 (N_22062,N_19634,N_20309);
xor U22063 (N_22063,N_19868,N_20544);
nand U22064 (N_22064,N_19589,N_20792);
nand U22065 (N_22065,N_20722,N_20894);
xnor U22066 (N_22066,N_20796,N_19661);
xor U22067 (N_22067,N_20279,N_20878);
xnor U22068 (N_22068,N_20064,N_20363);
xor U22069 (N_22069,N_20700,N_20805);
and U22070 (N_22070,N_20826,N_20267);
nand U22071 (N_22071,N_20430,N_20442);
and U22072 (N_22072,N_20264,N_20297);
nor U22073 (N_22073,N_20458,N_19597);
xor U22074 (N_22074,N_19785,N_20252);
and U22075 (N_22075,N_19903,N_19709);
nand U22076 (N_22076,N_20034,N_20205);
xor U22077 (N_22077,N_19932,N_20914);
nand U22078 (N_22078,N_20861,N_20983);
nand U22079 (N_22079,N_19722,N_20208);
nor U22080 (N_22080,N_20928,N_19805);
and U22081 (N_22081,N_20247,N_20783);
nand U22082 (N_22082,N_20422,N_20693);
nand U22083 (N_22083,N_19613,N_19761);
or U22084 (N_22084,N_19553,N_19614);
nor U22085 (N_22085,N_20820,N_20780);
nor U22086 (N_22086,N_20260,N_20616);
and U22087 (N_22087,N_20976,N_20933);
nand U22088 (N_22088,N_20728,N_20899);
and U22089 (N_22089,N_20532,N_20736);
nand U22090 (N_22090,N_20959,N_20267);
nor U22091 (N_22091,N_20991,N_20264);
and U22092 (N_22092,N_19657,N_20022);
or U22093 (N_22093,N_19674,N_20923);
nand U22094 (N_22094,N_19800,N_20622);
nor U22095 (N_22095,N_20476,N_20787);
xnor U22096 (N_22096,N_20654,N_20618);
xor U22097 (N_22097,N_20796,N_20567);
and U22098 (N_22098,N_20382,N_20007);
or U22099 (N_22099,N_20755,N_19646);
or U22100 (N_22100,N_20529,N_20789);
or U22101 (N_22101,N_20077,N_20003);
or U22102 (N_22102,N_20822,N_20394);
or U22103 (N_22103,N_20604,N_19588);
xnor U22104 (N_22104,N_20970,N_20632);
xnor U22105 (N_22105,N_19656,N_20108);
xnor U22106 (N_22106,N_19637,N_19743);
or U22107 (N_22107,N_19818,N_20886);
nand U22108 (N_22108,N_20385,N_20912);
nand U22109 (N_22109,N_20882,N_20232);
nor U22110 (N_22110,N_19825,N_20396);
nor U22111 (N_22111,N_20334,N_20728);
nor U22112 (N_22112,N_20704,N_20333);
or U22113 (N_22113,N_19656,N_19504);
or U22114 (N_22114,N_20280,N_19788);
nor U22115 (N_22115,N_19866,N_20640);
xor U22116 (N_22116,N_19703,N_20045);
xnor U22117 (N_22117,N_20303,N_20823);
xor U22118 (N_22118,N_20716,N_19774);
or U22119 (N_22119,N_20186,N_19602);
xnor U22120 (N_22120,N_19709,N_19889);
and U22121 (N_22121,N_19902,N_20339);
or U22122 (N_22122,N_20106,N_19866);
or U22123 (N_22123,N_20313,N_20316);
or U22124 (N_22124,N_20316,N_20859);
or U22125 (N_22125,N_20687,N_20427);
nand U22126 (N_22126,N_19808,N_20529);
nor U22127 (N_22127,N_20860,N_20300);
or U22128 (N_22128,N_20569,N_19697);
xnor U22129 (N_22129,N_20493,N_20018);
nand U22130 (N_22130,N_19836,N_20995);
nand U22131 (N_22131,N_20519,N_20909);
xnor U22132 (N_22132,N_20028,N_20658);
nor U22133 (N_22133,N_20041,N_20829);
or U22134 (N_22134,N_19580,N_19920);
xor U22135 (N_22135,N_20246,N_20640);
nand U22136 (N_22136,N_20179,N_19671);
nor U22137 (N_22137,N_19932,N_19733);
nand U22138 (N_22138,N_19562,N_19611);
and U22139 (N_22139,N_20420,N_19842);
and U22140 (N_22140,N_20262,N_20654);
nand U22141 (N_22141,N_20168,N_20263);
or U22142 (N_22142,N_20897,N_19890);
and U22143 (N_22143,N_19907,N_20270);
and U22144 (N_22144,N_20213,N_20720);
xnor U22145 (N_22145,N_20962,N_19840);
xor U22146 (N_22146,N_20175,N_19956);
or U22147 (N_22147,N_20904,N_19666);
nand U22148 (N_22148,N_20894,N_20058);
or U22149 (N_22149,N_19746,N_20064);
and U22150 (N_22150,N_20012,N_20252);
or U22151 (N_22151,N_20517,N_20981);
xor U22152 (N_22152,N_20402,N_20207);
xnor U22153 (N_22153,N_19986,N_20035);
nor U22154 (N_22154,N_20100,N_20190);
and U22155 (N_22155,N_20819,N_19890);
xor U22156 (N_22156,N_20889,N_19646);
nor U22157 (N_22157,N_20229,N_19704);
xnor U22158 (N_22158,N_20284,N_20849);
and U22159 (N_22159,N_20873,N_19519);
xor U22160 (N_22160,N_20637,N_20243);
xor U22161 (N_22161,N_20218,N_19713);
xnor U22162 (N_22162,N_20899,N_20990);
and U22163 (N_22163,N_20400,N_20240);
or U22164 (N_22164,N_20273,N_20303);
nand U22165 (N_22165,N_20274,N_20351);
xnor U22166 (N_22166,N_19964,N_19599);
nand U22167 (N_22167,N_20910,N_20891);
and U22168 (N_22168,N_19562,N_20039);
nand U22169 (N_22169,N_19663,N_20621);
and U22170 (N_22170,N_20356,N_20014);
xnor U22171 (N_22171,N_20718,N_20673);
or U22172 (N_22172,N_20270,N_19632);
xnor U22173 (N_22173,N_20155,N_20643);
and U22174 (N_22174,N_20995,N_20217);
xor U22175 (N_22175,N_20985,N_20602);
nand U22176 (N_22176,N_20440,N_20414);
xor U22177 (N_22177,N_19729,N_19526);
and U22178 (N_22178,N_20904,N_20731);
or U22179 (N_22179,N_20448,N_20298);
nor U22180 (N_22180,N_20060,N_20543);
or U22181 (N_22181,N_20052,N_20205);
nor U22182 (N_22182,N_20760,N_19768);
nor U22183 (N_22183,N_20876,N_19730);
nor U22184 (N_22184,N_19759,N_20030);
xor U22185 (N_22185,N_19869,N_19820);
or U22186 (N_22186,N_19783,N_19843);
and U22187 (N_22187,N_20036,N_19837);
and U22188 (N_22188,N_19664,N_20763);
or U22189 (N_22189,N_19565,N_19745);
and U22190 (N_22190,N_20877,N_20724);
nand U22191 (N_22191,N_20579,N_19944);
nand U22192 (N_22192,N_19666,N_20644);
nor U22193 (N_22193,N_19838,N_20672);
nor U22194 (N_22194,N_20432,N_20405);
nand U22195 (N_22195,N_20986,N_19635);
nor U22196 (N_22196,N_20474,N_20505);
or U22197 (N_22197,N_20074,N_20879);
xnor U22198 (N_22198,N_20283,N_20385);
xnor U22199 (N_22199,N_20440,N_20674);
nor U22200 (N_22200,N_19591,N_20951);
nor U22201 (N_22201,N_20556,N_20942);
or U22202 (N_22202,N_19783,N_19589);
and U22203 (N_22203,N_19576,N_20586);
xor U22204 (N_22204,N_19866,N_20799);
and U22205 (N_22205,N_20903,N_20729);
nor U22206 (N_22206,N_20494,N_19917);
or U22207 (N_22207,N_20898,N_20943);
or U22208 (N_22208,N_19766,N_20602);
nor U22209 (N_22209,N_19981,N_20253);
xor U22210 (N_22210,N_20773,N_20535);
nor U22211 (N_22211,N_20845,N_20349);
or U22212 (N_22212,N_19787,N_20185);
nor U22213 (N_22213,N_20096,N_20408);
xnor U22214 (N_22214,N_20363,N_20746);
nor U22215 (N_22215,N_20892,N_19966);
nand U22216 (N_22216,N_19656,N_19528);
xnor U22217 (N_22217,N_20373,N_19914);
xnor U22218 (N_22218,N_20181,N_19505);
xnor U22219 (N_22219,N_20458,N_20951);
or U22220 (N_22220,N_20986,N_20399);
nand U22221 (N_22221,N_20435,N_20808);
and U22222 (N_22222,N_20484,N_20143);
xor U22223 (N_22223,N_20734,N_20190);
or U22224 (N_22224,N_20837,N_20096);
or U22225 (N_22225,N_20576,N_20772);
nor U22226 (N_22226,N_19620,N_19935);
nand U22227 (N_22227,N_20762,N_19793);
or U22228 (N_22228,N_20459,N_20641);
nand U22229 (N_22229,N_20452,N_19597);
nand U22230 (N_22230,N_19691,N_19560);
nand U22231 (N_22231,N_20774,N_20297);
and U22232 (N_22232,N_20019,N_20643);
nand U22233 (N_22233,N_20195,N_19991);
nand U22234 (N_22234,N_20718,N_20193);
nor U22235 (N_22235,N_19789,N_20861);
nand U22236 (N_22236,N_20605,N_20272);
nor U22237 (N_22237,N_20564,N_20800);
and U22238 (N_22238,N_19791,N_20342);
and U22239 (N_22239,N_20395,N_20709);
or U22240 (N_22240,N_19507,N_19706);
or U22241 (N_22241,N_20466,N_20024);
or U22242 (N_22242,N_19782,N_20551);
nor U22243 (N_22243,N_19633,N_19856);
and U22244 (N_22244,N_20053,N_20360);
nor U22245 (N_22245,N_19821,N_19676);
or U22246 (N_22246,N_20138,N_20683);
nand U22247 (N_22247,N_20465,N_20744);
or U22248 (N_22248,N_20866,N_20643);
nor U22249 (N_22249,N_20745,N_20550);
and U22250 (N_22250,N_20333,N_20881);
nor U22251 (N_22251,N_20996,N_19922);
and U22252 (N_22252,N_20754,N_19636);
nor U22253 (N_22253,N_19772,N_20814);
and U22254 (N_22254,N_19799,N_20996);
nand U22255 (N_22255,N_19589,N_20343);
or U22256 (N_22256,N_20055,N_19699);
and U22257 (N_22257,N_20527,N_20797);
or U22258 (N_22258,N_19760,N_20526);
and U22259 (N_22259,N_20693,N_20908);
nor U22260 (N_22260,N_20642,N_19787);
nor U22261 (N_22261,N_19705,N_20977);
or U22262 (N_22262,N_20577,N_19710);
nand U22263 (N_22263,N_19897,N_20956);
nand U22264 (N_22264,N_19700,N_20350);
xor U22265 (N_22265,N_20959,N_20189);
nor U22266 (N_22266,N_20834,N_20016);
or U22267 (N_22267,N_20327,N_20255);
and U22268 (N_22268,N_20222,N_19563);
and U22269 (N_22269,N_20300,N_19588);
nor U22270 (N_22270,N_20010,N_20396);
nand U22271 (N_22271,N_19710,N_20804);
or U22272 (N_22272,N_19798,N_20056);
and U22273 (N_22273,N_19761,N_19775);
nor U22274 (N_22274,N_20564,N_19904);
or U22275 (N_22275,N_19861,N_20576);
and U22276 (N_22276,N_19940,N_20064);
and U22277 (N_22277,N_20730,N_19979);
nor U22278 (N_22278,N_20126,N_20326);
nor U22279 (N_22279,N_19892,N_19660);
nand U22280 (N_22280,N_20845,N_19563);
xor U22281 (N_22281,N_20153,N_19729);
and U22282 (N_22282,N_20210,N_20931);
nand U22283 (N_22283,N_19936,N_20729);
xnor U22284 (N_22284,N_19695,N_19674);
nand U22285 (N_22285,N_20614,N_20222);
xor U22286 (N_22286,N_20421,N_20727);
or U22287 (N_22287,N_20930,N_20203);
or U22288 (N_22288,N_20201,N_20655);
or U22289 (N_22289,N_19808,N_19561);
xnor U22290 (N_22290,N_20947,N_20738);
nand U22291 (N_22291,N_20929,N_20817);
or U22292 (N_22292,N_19778,N_20807);
nor U22293 (N_22293,N_20888,N_19989);
nand U22294 (N_22294,N_20909,N_20391);
nor U22295 (N_22295,N_20753,N_20976);
nor U22296 (N_22296,N_20705,N_20497);
nand U22297 (N_22297,N_20446,N_19508);
or U22298 (N_22298,N_19792,N_20623);
nor U22299 (N_22299,N_19671,N_20224);
or U22300 (N_22300,N_19575,N_20296);
nand U22301 (N_22301,N_19650,N_20113);
and U22302 (N_22302,N_19732,N_20035);
and U22303 (N_22303,N_20891,N_20453);
nand U22304 (N_22304,N_20591,N_20104);
nand U22305 (N_22305,N_20800,N_20452);
xor U22306 (N_22306,N_20082,N_19925);
and U22307 (N_22307,N_19920,N_20318);
xor U22308 (N_22308,N_20448,N_20835);
or U22309 (N_22309,N_19710,N_20359);
and U22310 (N_22310,N_19638,N_20375);
xnor U22311 (N_22311,N_19931,N_20191);
or U22312 (N_22312,N_20076,N_20932);
nand U22313 (N_22313,N_19963,N_19669);
xnor U22314 (N_22314,N_20200,N_20725);
or U22315 (N_22315,N_20527,N_20400);
xor U22316 (N_22316,N_19762,N_20810);
nor U22317 (N_22317,N_19707,N_20959);
and U22318 (N_22318,N_19795,N_19782);
nand U22319 (N_22319,N_20846,N_19955);
nor U22320 (N_22320,N_20080,N_20946);
and U22321 (N_22321,N_20169,N_20475);
or U22322 (N_22322,N_20437,N_20823);
and U22323 (N_22323,N_19551,N_20939);
or U22324 (N_22324,N_20122,N_19653);
xor U22325 (N_22325,N_20202,N_20486);
and U22326 (N_22326,N_20577,N_20288);
or U22327 (N_22327,N_20546,N_20979);
nand U22328 (N_22328,N_19734,N_19889);
xnor U22329 (N_22329,N_20364,N_20598);
or U22330 (N_22330,N_19702,N_20776);
nand U22331 (N_22331,N_20781,N_20289);
and U22332 (N_22332,N_19894,N_20964);
nor U22333 (N_22333,N_20545,N_20027);
xnor U22334 (N_22334,N_20867,N_20144);
and U22335 (N_22335,N_20186,N_20683);
nor U22336 (N_22336,N_20114,N_20300);
nand U22337 (N_22337,N_19667,N_19917);
xor U22338 (N_22338,N_20245,N_20058);
nand U22339 (N_22339,N_19936,N_20806);
or U22340 (N_22340,N_20713,N_20711);
and U22341 (N_22341,N_20600,N_20987);
nand U22342 (N_22342,N_20917,N_20179);
and U22343 (N_22343,N_20064,N_20430);
or U22344 (N_22344,N_20455,N_20745);
nand U22345 (N_22345,N_20347,N_20901);
or U22346 (N_22346,N_19907,N_19505);
xnor U22347 (N_22347,N_19622,N_19818);
and U22348 (N_22348,N_20945,N_19963);
nor U22349 (N_22349,N_20809,N_20917);
nand U22350 (N_22350,N_20426,N_20688);
xor U22351 (N_22351,N_19879,N_19809);
nand U22352 (N_22352,N_19988,N_19810);
or U22353 (N_22353,N_20991,N_20408);
or U22354 (N_22354,N_20649,N_19634);
or U22355 (N_22355,N_19621,N_20802);
and U22356 (N_22356,N_19550,N_20096);
nor U22357 (N_22357,N_19697,N_20919);
nor U22358 (N_22358,N_19702,N_20294);
nor U22359 (N_22359,N_20666,N_19759);
or U22360 (N_22360,N_20024,N_20052);
nand U22361 (N_22361,N_20658,N_20821);
nand U22362 (N_22362,N_20276,N_20267);
nor U22363 (N_22363,N_19811,N_20692);
and U22364 (N_22364,N_20127,N_19794);
and U22365 (N_22365,N_20192,N_20791);
xor U22366 (N_22366,N_20571,N_19994);
nor U22367 (N_22367,N_20434,N_20352);
nor U22368 (N_22368,N_19863,N_20888);
nand U22369 (N_22369,N_20415,N_20708);
or U22370 (N_22370,N_20061,N_19896);
or U22371 (N_22371,N_20506,N_20740);
nor U22372 (N_22372,N_20270,N_19543);
nor U22373 (N_22373,N_19731,N_20664);
or U22374 (N_22374,N_20485,N_19911);
nor U22375 (N_22375,N_19517,N_20208);
xor U22376 (N_22376,N_20907,N_20626);
xnor U22377 (N_22377,N_19798,N_19650);
xor U22378 (N_22378,N_20175,N_19740);
or U22379 (N_22379,N_20117,N_20900);
and U22380 (N_22380,N_20651,N_20004);
nor U22381 (N_22381,N_20692,N_20708);
and U22382 (N_22382,N_20836,N_20243);
nand U22383 (N_22383,N_20592,N_19666);
nor U22384 (N_22384,N_19868,N_20481);
or U22385 (N_22385,N_20334,N_20583);
and U22386 (N_22386,N_19978,N_20425);
and U22387 (N_22387,N_19729,N_20810);
or U22388 (N_22388,N_19730,N_20683);
xnor U22389 (N_22389,N_20292,N_19664);
nand U22390 (N_22390,N_20079,N_20396);
xor U22391 (N_22391,N_20648,N_19811);
nand U22392 (N_22392,N_20401,N_20534);
nor U22393 (N_22393,N_20263,N_19688);
nand U22394 (N_22394,N_20345,N_20365);
or U22395 (N_22395,N_20396,N_19782);
nor U22396 (N_22396,N_20511,N_20731);
and U22397 (N_22397,N_20982,N_20650);
and U22398 (N_22398,N_20803,N_20683);
xnor U22399 (N_22399,N_20243,N_20944);
and U22400 (N_22400,N_19578,N_20642);
or U22401 (N_22401,N_19670,N_19806);
nand U22402 (N_22402,N_19606,N_20932);
nor U22403 (N_22403,N_20609,N_20213);
xnor U22404 (N_22404,N_19676,N_19801);
xnor U22405 (N_22405,N_20470,N_19700);
and U22406 (N_22406,N_20771,N_20874);
nor U22407 (N_22407,N_19853,N_20302);
and U22408 (N_22408,N_20238,N_20451);
nor U22409 (N_22409,N_20949,N_20867);
or U22410 (N_22410,N_20572,N_20097);
xnor U22411 (N_22411,N_19892,N_19541);
or U22412 (N_22412,N_20918,N_20588);
nor U22413 (N_22413,N_20496,N_20519);
xnor U22414 (N_22414,N_19787,N_19669);
xor U22415 (N_22415,N_20580,N_19616);
xnor U22416 (N_22416,N_20713,N_19657);
nor U22417 (N_22417,N_19742,N_20242);
xor U22418 (N_22418,N_20464,N_20143);
and U22419 (N_22419,N_20044,N_19829);
and U22420 (N_22420,N_20997,N_20994);
nor U22421 (N_22421,N_20539,N_20421);
and U22422 (N_22422,N_20996,N_19975);
xor U22423 (N_22423,N_20599,N_19592);
or U22424 (N_22424,N_19650,N_20461);
xnor U22425 (N_22425,N_19829,N_20549);
nor U22426 (N_22426,N_20653,N_20332);
xor U22427 (N_22427,N_19795,N_19508);
and U22428 (N_22428,N_20949,N_19998);
or U22429 (N_22429,N_20095,N_19857);
or U22430 (N_22430,N_20798,N_20155);
or U22431 (N_22431,N_20729,N_19823);
and U22432 (N_22432,N_20452,N_20338);
or U22433 (N_22433,N_19745,N_20745);
or U22434 (N_22434,N_20186,N_20794);
xor U22435 (N_22435,N_20670,N_20253);
or U22436 (N_22436,N_19620,N_19706);
xor U22437 (N_22437,N_20075,N_20959);
or U22438 (N_22438,N_20100,N_19776);
xnor U22439 (N_22439,N_20421,N_20201);
xor U22440 (N_22440,N_19514,N_20931);
xnor U22441 (N_22441,N_20410,N_20210);
xnor U22442 (N_22442,N_19987,N_20548);
and U22443 (N_22443,N_20661,N_19990);
xor U22444 (N_22444,N_20890,N_19874);
xnor U22445 (N_22445,N_20820,N_20639);
nand U22446 (N_22446,N_20766,N_20977);
or U22447 (N_22447,N_20426,N_20763);
or U22448 (N_22448,N_20737,N_20462);
xnor U22449 (N_22449,N_20035,N_20364);
or U22450 (N_22450,N_20583,N_20396);
or U22451 (N_22451,N_19843,N_20525);
and U22452 (N_22452,N_20532,N_20849);
and U22453 (N_22453,N_20746,N_20520);
xnor U22454 (N_22454,N_20278,N_20428);
and U22455 (N_22455,N_20424,N_19702);
and U22456 (N_22456,N_20168,N_20490);
nand U22457 (N_22457,N_19517,N_19796);
nand U22458 (N_22458,N_20266,N_19774);
xnor U22459 (N_22459,N_20898,N_20460);
xor U22460 (N_22460,N_20416,N_19688);
nor U22461 (N_22461,N_19743,N_19615);
or U22462 (N_22462,N_20293,N_19642);
nor U22463 (N_22463,N_19698,N_19566);
and U22464 (N_22464,N_20177,N_20856);
xor U22465 (N_22465,N_19857,N_20988);
and U22466 (N_22466,N_20620,N_19755);
xnor U22467 (N_22467,N_19586,N_20294);
xnor U22468 (N_22468,N_20906,N_19640);
and U22469 (N_22469,N_19987,N_19618);
xnor U22470 (N_22470,N_19768,N_20790);
xor U22471 (N_22471,N_19982,N_20285);
and U22472 (N_22472,N_19579,N_19576);
nand U22473 (N_22473,N_20466,N_19606);
xor U22474 (N_22474,N_20799,N_20703);
nor U22475 (N_22475,N_20076,N_19947);
xnor U22476 (N_22476,N_20158,N_19858);
or U22477 (N_22477,N_19715,N_20376);
nand U22478 (N_22478,N_20180,N_19875);
nor U22479 (N_22479,N_19559,N_19712);
nand U22480 (N_22480,N_19504,N_19630);
or U22481 (N_22481,N_20156,N_20494);
or U22482 (N_22482,N_20045,N_20819);
and U22483 (N_22483,N_19687,N_19927);
xnor U22484 (N_22484,N_20301,N_19722);
and U22485 (N_22485,N_20775,N_20904);
or U22486 (N_22486,N_20929,N_19518);
and U22487 (N_22487,N_20426,N_20406);
nor U22488 (N_22488,N_19825,N_20616);
and U22489 (N_22489,N_19689,N_20257);
or U22490 (N_22490,N_19838,N_19718);
nand U22491 (N_22491,N_20457,N_19835);
nand U22492 (N_22492,N_19937,N_20120);
nand U22493 (N_22493,N_20021,N_19689);
or U22494 (N_22494,N_20911,N_20153);
xor U22495 (N_22495,N_19981,N_20234);
nand U22496 (N_22496,N_19816,N_19661);
nand U22497 (N_22497,N_20604,N_19739);
and U22498 (N_22498,N_20516,N_19800);
xnor U22499 (N_22499,N_20345,N_20053);
xnor U22500 (N_22500,N_21015,N_21654);
nand U22501 (N_22501,N_22213,N_22227);
and U22502 (N_22502,N_22115,N_21609);
nor U22503 (N_22503,N_21788,N_22149);
or U22504 (N_22504,N_22049,N_21324);
nor U22505 (N_22505,N_22377,N_22247);
nor U22506 (N_22506,N_22085,N_21519);
xnor U22507 (N_22507,N_22343,N_21247);
xnor U22508 (N_22508,N_21532,N_21351);
or U22509 (N_22509,N_21093,N_21781);
or U22510 (N_22510,N_22361,N_21742);
nor U22511 (N_22511,N_21523,N_21619);
and U22512 (N_22512,N_21293,N_21566);
nor U22513 (N_22513,N_21848,N_21049);
or U22514 (N_22514,N_21269,N_21320);
and U22515 (N_22515,N_21404,N_21747);
nand U22516 (N_22516,N_21348,N_21760);
xnor U22517 (N_22517,N_22367,N_22057);
nor U22518 (N_22518,N_22028,N_22417);
nor U22519 (N_22519,N_21514,N_21004);
or U22520 (N_22520,N_21708,N_22069);
xnor U22521 (N_22521,N_21211,N_21309);
and U22522 (N_22522,N_21575,N_22114);
or U22523 (N_22523,N_21552,N_21969);
nor U22524 (N_22524,N_22026,N_21393);
and U22525 (N_22525,N_22186,N_21664);
or U22526 (N_22526,N_21653,N_21376);
nor U22527 (N_22527,N_21895,N_22283);
nor U22528 (N_22528,N_21524,N_21463);
or U22529 (N_22529,N_21974,N_21581);
xor U22530 (N_22530,N_21028,N_21938);
xor U22531 (N_22531,N_21842,N_21407);
nor U22532 (N_22532,N_21190,N_22230);
nand U22533 (N_22533,N_21952,N_21037);
and U22534 (N_22534,N_21979,N_21606);
or U22535 (N_22535,N_22233,N_21198);
nand U22536 (N_22536,N_21806,N_21216);
nor U22537 (N_22537,N_21985,N_22051);
and U22538 (N_22538,N_22327,N_21713);
or U22539 (N_22539,N_21888,N_22487);
nand U22540 (N_22540,N_21811,N_22393);
or U22541 (N_22541,N_21295,N_22324);
and U22542 (N_22542,N_22300,N_21438);
or U22543 (N_22543,N_21744,N_21548);
and U22544 (N_22544,N_21573,N_22212);
nand U22545 (N_22545,N_21262,N_22007);
or U22546 (N_22546,N_21599,N_21264);
xor U22547 (N_22547,N_21927,N_21214);
nor U22548 (N_22548,N_21425,N_22036);
and U22549 (N_22549,N_21650,N_21821);
or U22550 (N_22550,N_22365,N_21881);
nor U22551 (N_22551,N_21586,N_22265);
xor U22552 (N_22552,N_22132,N_21521);
and U22553 (N_22553,N_21738,N_21671);
nand U22554 (N_22554,N_21851,N_21899);
nor U22555 (N_22555,N_21535,N_21601);
nand U22556 (N_22556,N_22122,N_22474);
or U22557 (N_22557,N_21017,N_21836);
and U22558 (N_22558,N_22158,N_21429);
or U22559 (N_22559,N_22496,N_21593);
xnor U22560 (N_22560,N_21477,N_21000);
nor U22561 (N_22561,N_21580,N_21166);
nand U22562 (N_22562,N_21560,N_22145);
and U22563 (N_22563,N_21289,N_22330);
nand U22564 (N_22564,N_22329,N_22005);
and U22565 (N_22565,N_21648,N_21319);
nor U22566 (N_22566,N_21427,N_21499);
nand U22567 (N_22567,N_22254,N_21106);
nor U22568 (N_22568,N_21456,N_21423);
xnor U22569 (N_22569,N_21692,N_21257);
nand U22570 (N_22570,N_21200,N_21873);
and U22571 (N_22571,N_22066,N_22205);
or U22572 (N_22572,N_22086,N_22054);
nor U22573 (N_22573,N_21870,N_21451);
and U22574 (N_22574,N_21646,N_22434);
and U22575 (N_22575,N_21364,N_21547);
and U22576 (N_22576,N_22243,N_22075);
nand U22577 (N_22577,N_21164,N_21074);
nor U22578 (N_22578,N_21911,N_22134);
nand U22579 (N_22579,N_22137,N_22295);
nand U22580 (N_22580,N_21255,N_22299);
or U22581 (N_22581,N_21623,N_21071);
and U22582 (N_22582,N_21468,N_22089);
and U22583 (N_22583,N_21131,N_21626);
nand U22584 (N_22584,N_21943,N_22201);
nand U22585 (N_22585,N_22091,N_21909);
nor U22586 (N_22586,N_22311,N_22237);
nand U22587 (N_22587,N_21600,N_21119);
nand U22588 (N_22588,N_21445,N_21908);
and U22589 (N_22589,N_21898,N_21259);
and U22590 (N_22590,N_21687,N_22152);
xor U22591 (N_22591,N_21805,N_21418);
and U22592 (N_22592,N_21414,N_21210);
nor U22593 (N_22593,N_21267,N_21602);
nand U22594 (N_22594,N_21256,N_21750);
and U22595 (N_22595,N_21780,N_21428);
xnor U22596 (N_22596,N_21276,N_22498);
xor U22597 (N_22597,N_22409,N_21820);
nor U22598 (N_22598,N_21622,N_22470);
and U22599 (N_22599,N_21846,N_21349);
nor U22600 (N_22600,N_21857,N_22154);
or U22601 (N_22601,N_21534,N_22253);
or U22602 (N_22602,N_21620,N_21834);
nor U22603 (N_22603,N_22079,N_21167);
and U22604 (N_22604,N_21745,N_21641);
xor U22605 (N_22605,N_21125,N_22339);
nor U22606 (N_22606,N_21040,N_21545);
nor U22607 (N_22607,N_21287,N_21826);
nand U22608 (N_22608,N_21946,N_21053);
or U22609 (N_22609,N_22484,N_21526);
nor U22610 (N_22610,N_22156,N_22387);
and U22611 (N_22611,N_22379,N_22298);
nor U22612 (N_22612,N_21582,N_22171);
nand U22613 (N_22613,N_22297,N_21371);
nand U22614 (N_22614,N_21486,N_21512);
and U22615 (N_22615,N_21789,N_21239);
xnor U22616 (N_22616,N_21224,N_21151);
nand U22617 (N_22617,N_22406,N_22431);
xor U22618 (N_22618,N_22194,N_21841);
xnor U22619 (N_22619,N_21629,N_21241);
or U22620 (N_22620,N_22155,N_21921);
nor U22621 (N_22621,N_22053,N_22002);
or U22622 (N_22622,N_21882,N_21819);
or U22623 (N_22623,N_21672,N_21301);
or U22624 (N_22624,N_22466,N_21492);
xnor U22625 (N_22625,N_21448,N_21591);
and U22626 (N_22626,N_22318,N_21651);
nand U22627 (N_22627,N_22123,N_21299);
or U22628 (N_22628,N_21402,N_22317);
or U22629 (N_22629,N_21929,N_21060);
nand U22630 (N_22630,N_22314,N_22306);
xnor U22631 (N_22631,N_21459,N_21977);
nand U22632 (N_22632,N_21139,N_22142);
and U22633 (N_22633,N_22093,N_21073);
nand U22634 (N_22634,N_21827,N_22218);
or U22635 (N_22635,N_21755,N_21122);
or U22636 (N_22636,N_21507,N_22364);
nand U22637 (N_22637,N_22291,N_21416);
nand U22638 (N_22638,N_21022,N_21754);
and U22639 (N_22639,N_21003,N_22178);
xnor U22640 (N_22640,N_21987,N_21808);
nand U22641 (N_22641,N_21598,N_22337);
nand U22642 (N_22642,N_22479,N_21809);
nand U22643 (N_22643,N_21767,N_21434);
nor U22644 (N_22644,N_21610,N_22362);
and U22645 (N_22645,N_21368,N_22183);
nand U22646 (N_22646,N_21978,N_22457);
nor U22647 (N_22647,N_22344,N_21705);
nand U22648 (N_22648,N_21104,N_21226);
or U22649 (N_22649,N_22226,N_21678);
xnor U22650 (N_22650,N_21695,N_22217);
xor U22651 (N_22651,N_21587,N_21147);
xnor U22652 (N_22652,N_21994,N_22032);
and U22653 (N_22653,N_21859,N_22220);
or U22654 (N_22654,N_22181,N_22354);
or U22655 (N_22655,N_22133,N_21197);
nor U22656 (N_22656,N_21454,N_22004);
nand U22657 (N_22657,N_21718,N_21730);
nor U22658 (N_22658,N_21904,N_21172);
or U22659 (N_22659,N_21228,N_22196);
nor U22660 (N_22660,N_21694,N_21174);
nand U22661 (N_22661,N_21719,N_22430);
nor U22662 (N_22662,N_21607,N_21018);
nor U22663 (N_22663,N_21356,N_21288);
nor U22664 (N_22664,N_22222,N_21035);
xor U22665 (N_22665,N_22296,N_21799);
nor U22666 (N_22666,N_22141,N_21594);
and U22667 (N_22667,N_22232,N_21530);
xor U22668 (N_22668,N_21373,N_21308);
nand U22669 (N_22669,N_21564,N_21922);
and U22670 (N_22670,N_21081,N_21885);
nand U22671 (N_22671,N_22353,N_22103);
xnor U22672 (N_22672,N_22345,N_21871);
and U22673 (N_22673,N_22485,N_21618);
and U22674 (N_22674,N_22424,N_21804);
nand U22675 (N_22675,N_21701,N_22419);
xnor U22676 (N_22676,N_22094,N_21362);
nand U22677 (N_22677,N_21070,N_21441);
nor U22678 (N_22678,N_21382,N_22476);
xnor U22679 (N_22679,N_22077,N_22308);
xnor U22680 (N_22680,N_21406,N_21966);
nor U22681 (N_22681,N_21115,N_21274);
xnor U22682 (N_22682,N_21249,N_21891);
or U22683 (N_22683,N_22463,N_21931);
nor U22684 (N_22684,N_21263,N_21075);
or U22685 (N_22685,N_21498,N_21945);
xnor U22686 (N_22686,N_21509,N_22246);
or U22687 (N_22687,N_21177,N_21778);
nand U22688 (N_22688,N_21518,N_21111);
or U22689 (N_22689,N_22319,N_21457);
and U22690 (N_22690,N_21220,N_21996);
nor U22691 (N_22691,N_22411,N_21307);
nand U22692 (N_22692,N_22348,N_21019);
and U22693 (N_22693,N_21900,N_21417);
nand U22694 (N_22694,N_21689,N_22277);
nor U22695 (N_22695,N_21387,N_21967);
nand U22696 (N_22696,N_22003,N_21411);
and U22697 (N_22697,N_21655,N_21658);
nor U22698 (N_22698,N_21303,N_21992);
and U22699 (N_22699,N_21148,N_22366);
nor U22700 (N_22700,N_21331,N_21500);
nand U22701 (N_22701,N_21325,N_21849);
nand U22702 (N_22702,N_21143,N_22428);
nand U22703 (N_22703,N_21699,N_21209);
or U22704 (N_22704,N_21076,N_21732);
nand U22705 (N_22705,N_22398,N_21603);
nor U22706 (N_22706,N_22280,N_22396);
xor U22707 (N_22707,N_22322,N_21686);
and U22708 (N_22708,N_22199,N_21085);
nor U22709 (N_22709,N_22117,N_21196);
nand U22710 (N_22710,N_21972,N_22017);
or U22711 (N_22711,N_22260,N_21893);
nand U22712 (N_22712,N_21522,N_21207);
or U22713 (N_22713,N_22432,N_21752);
nor U22714 (N_22714,N_22338,N_22235);
xor U22715 (N_22715,N_22302,N_21481);
and U22716 (N_22716,N_21777,N_22106);
or U22717 (N_22717,N_22349,N_21999);
xnor U22718 (N_22718,N_22290,N_21424);
xor U22719 (N_22719,N_22058,N_22207);
or U22720 (N_22720,N_22165,N_22175);
and U22721 (N_22721,N_21916,N_21579);
or U22722 (N_22722,N_21092,N_21171);
xnor U22723 (N_22723,N_22381,N_21627);
nand U22724 (N_22724,N_22261,N_22346);
nand U22725 (N_22725,N_21940,N_22064);
nor U22726 (N_22726,N_21828,N_21543);
and U22727 (N_22727,N_21229,N_21991);
xnor U22728 (N_22728,N_21219,N_21011);
or U22729 (N_22729,N_21935,N_21300);
nor U22730 (N_22730,N_21791,N_22000);
or U22731 (N_22731,N_21185,N_21955);
xnor U22732 (N_22732,N_22489,N_21989);
nor U22733 (N_22733,N_22334,N_21926);
and U22734 (N_22734,N_21915,N_21595);
xnor U22735 (N_22735,N_22259,N_21298);
or U22736 (N_22736,N_22042,N_21258);
xnor U22737 (N_22737,N_21964,N_22011);
nor U22738 (N_22738,N_21659,N_21772);
nand U22739 (N_22739,N_21690,N_21234);
or U22740 (N_22740,N_22073,N_22124);
and U22741 (N_22741,N_21390,N_22138);
nand U22742 (N_22742,N_21735,N_22391);
and U22743 (N_22743,N_22458,N_22490);
nand U22744 (N_22744,N_22161,N_21831);
nor U22745 (N_22745,N_22090,N_22030);
nor U22746 (N_22746,N_22150,N_21867);
and U22747 (N_22747,N_21576,N_21050);
nand U22748 (N_22748,N_21759,N_22013);
nand U22749 (N_22749,N_21322,N_21124);
or U22750 (N_22750,N_21715,N_22310);
xnor U22751 (N_22751,N_21910,N_21795);
xor U22752 (N_22752,N_21557,N_22410);
and U22753 (N_22753,N_21590,N_21561);
nand U22754 (N_22754,N_22376,N_21936);
and U22755 (N_22755,N_21728,N_21956);
and U22756 (N_22756,N_21639,N_22080);
nor U22757 (N_22757,N_21923,N_21397);
nand U22758 (N_22758,N_21511,N_21473);
nand U22759 (N_22759,N_21129,N_21311);
xor U22760 (N_22760,N_21764,N_21377);
xor U22761 (N_22761,N_22021,N_22435);
and U22762 (N_22762,N_22200,N_21367);
and U22763 (N_22763,N_21178,N_22350);
nor U22764 (N_22764,N_21769,N_21027);
xor U22765 (N_22765,N_21890,N_21845);
xnor U22766 (N_22766,N_21903,N_21280);
xor U22767 (N_22767,N_22284,N_22305);
nand U22768 (N_22768,N_22228,N_22481);
xnor U22769 (N_22769,N_21879,N_21152);
nor U22770 (N_22770,N_22016,N_21674);
nand U22771 (N_22771,N_21538,N_22340);
nand U22772 (N_22772,N_22312,N_22245);
xor U22773 (N_22773,N_21757,N_21458);
or U22774 (N_22774,N_22369,N_22068);
or U22775 (N_22775,N_21937,N_22275);
nand U22776 (N_22776,N_21297,N_22048);
or U22777 (N_22777,N_21822,N_21201);
or U22778 (N_22778,N_21496,N_21688);
nand U22779 (N_22779,N_21057,N_21948);
and U22780 (N_22780,N_21268,N_21230);
and U22781 (N_22781,N_21608,N_21774);
nor U22782 (N_22782,N_21472,N_21170);
xnor U22783 (N_22783,N_21012,N_21634);
xnor U22784 (N_22784,N_22143,N_21874);
nor U22785 (N_22785,N_21612,N_22110);
xor U22786 (N_22786,N_22486,N_22234);
and U22787 (N_22787,N_22248,N_21667);
nor U22788 (N_22788,N_21635,N_21140);
or U22789 (N_22789,N_22015,N_21829);
and U22790 (N_22790,N_21852,N_21316);
nor U22791 (N_22791,N_21668,N_21630);
xor U22792 (N_22792,N_22440,N_21254);
or U22793 (N_22793,N_21624,N_21340);
or U22794 (N_22794,N_21783,N_21768);
xnor U22795 (N_22795,N_22482,N_21717);
and U22796 (N_22796,N_21984,N_22425);
and U22797 (N_22797,N_21408,N_21782);
and U22798 (N_22798,N_21370,N_21285);
and U22799 (N_22799,N_21026,N_21702);
and U22800 (N_22800,N_22444,N_22426);
xnor U22801 (N_22801,N_22266,N_21327);
or U22802 (N_22802,N_21378,N_22179);
or U22803 (N_22803,N_21313,N_21491);
nor U22804 (N_22804,N_22169,N_21628);
xor U22805 (N_22805,N_21998,N_22342);
nor U22806 (N_22806,N_21227,N_22413);
or U22807 (N_22807,N_21321,N_21054);
and U22808 (N_22808,N_22109,N_22383);
nand U22809 (N_22809,N_22006,N_21246);
xnor U22810 (N_22810,N_21539,N_21217);
and U22811 (N_22811,N_21918,N_21968);
nand U22812 (N_22812,N_21310,N_21508);
nor U22813 (N_22813,N_21711,N_21913);
nand U22814 (N_22814,N_21181,N_22164);
xor U22815 (N_22815,N_21030,N_21120);
nand U22816 (N_22816,N_22400,N_22035);
and U22817 (N_22817,N_21160,N_22041);
nand U22818 (N_22818,N_21363,N_22174);
nor U22819 (N_22819,N_22416,N_21208);
and U22820 (N_22820,N_21105,N_21133);
xor U22821 (N_22821,N_22162,N_22148);
or U22822 (N_22822,N_22371,N_21475);
or U22823 (N_22823,N_21957,N_21381);
nor U22824 (N_22824,N_21415,N_22412);
and U22825 (N_22825,N_21064,N_22188);
nand U22826 (N_22826,N_21965,N_21544);
and U22827 (N_22827,N_21880,N_21676);
xor U22828 (N_22828,N_21329,N_21856);
or U22829 (N_22829,N_21215,N_21592);
nor U22830 (N_22830,N_22325,N_22304);
xnor U22831 (N_22831,N_21596,N_22039);
or U22832 (N_22832,N_21084,N_21047);
or U22833 (N_22833,N_21981,N_21951);
or U22834 (N_22834,N_21565,N_21335);
or U22835 (N_22835,N_21077,N_22257);
or U22836 (N_22836,N_22214,N_21248);
or U22837 (N_22837,N_21144,N_21088);
nor U22838 (N_22838,N_21420,N_22076);
nor U22839 (N_22839,N_21005,N_21354);
nand U22840 (N_22840,N_22018,N_21396);
or U22841 (N_22841,N_21095,N_21398);
and U22842 (N_22842,N_21155,N_22052);
and U22843 (N_22843,N_21275,N_22352);
nand U22844 (N_22844,N_22001,N_21912);
xor U22845 (N_22845,N_22014,N_21533);
nor U22846 (N_22846,N_21680,N_21621);
xnor U22847 (N_22847,N_22384,N_21282);
xnor U22848 (N_22848,N_21542,N_21344);
nand U22849 (N_22849,N_22388,N_22336);
nor U22850 (N_22850,N_21357,N_22170);
nand U22851 (N_22851,N_22236,N_21379);
or U22852 (N_22852,N_21640,N_21684);
nor U22853 (N_22853,N_21839,N_22159);
xnor U22854 (N_22854,N_21787,N_22357);
or U22855 (N_22855,N_21366,N_22370);
nand U22856 (N_22856,N_21691,N_21986);
or U22857 (N_22857,N_22099,N_21555);
nor U22858 (N_22858,N_21665,N_21644);
xor U22859 (N_22859,N_21273,N_21189);
or U22860 (N_22860,N_22456,N_21703);
nor U22861 (N_22861,N_21146,N_21698);
nor U22862 (N_22862,N_22439,N_22111);
and U22863 (N_22863,N_21484,N_21920);
or U22864 (N_22864,N_22081,N_22211);
and U22865 (N_22865,N_21260,N_21212);
xor U22866 (N_22866,N_21505,N_21221);
and U22867 (N_22867,N_22125,N_22373);
nand U22868 (N_22868,N_22009,N_22022);
nor U22869 (N_22869,N_21961,N_21014);
and U22870 (N_22870,N_21504,N_21435);
nor U22871 (N_22871,N_21816,N_22475);
and U22872 (N_22872,N_22287,N_22210);
nor U22873 (N_22873,N_21034,N_21007);
xor U22874 (N_22874,N_22151,N_22157);
xnor U22875 (N_22875,N_21461,N_21862);
nand U22876 (N_22876,N_21589,N_22182);
nor U22877 (N_22877,N_21110,N_21163);
nor U22878 (N_22878,N_21860,N_22029);
nor U22879 (N_22879,N_21008,N_21103);
xnor U22880 (N_22880,N_21467,N_21765);
nor U22881 (N_22881,N_21825,N_22092);
nand U22882 (N_22882,N_22119,N_21339);
nand U22883 (N_22883,N_22395,N_21696);
nand U22884 (N_22884,N_22040,N_21089);
and U22885 (N_22885,N_22067,N_21520);
nor U22886 (N_22886,N_21240,N_22140);
or U22887 (N_22887,N_22131,N_21395);
nor U22888 (N_22888,N_21854,N_21059);
xnor U22889 (N_22889,N_21213,N_21182);
nand U22890 (N_22890,N_21355,N_21063);
nand U22891 (N_22891,N_22368,N_21305);
and U22892 (N_22892,N_21066,N_22043);
and U22893 (N_22893,N_21290,N_21959);
or U22894 (N_22894,N_22065,N_22045);
xnor U22895 (N_22895,N_21261,N_22445);
xnor U22896 (N_22896,N_22269,N_21332);
nor U22897 (N_22897,N_21861,N_21494);
and U22898 (N_22898,N_21412,N_21479);
nor U22899 (N_22899,N_21315,N_22191);
and U22900 (N_22900,N_22087,N_21132);
nor U22901 (N_22901,N_21531,N_21675);
and U22902 (N_22902,N_21374,N_21361);
and U22903 (N_22903,N_22146,N_21540);
or U22904 (N_22904,N_21762,N_21384);
xor U22905 (N_22905,N_21932,N_21126);
nand U22906 (N_22906,N_21934,N_22168);
xnor U22907 (N_22907,N_21562,N_22184);
or U22908 (N_22908,N_21453,N_22378);
nor U22909 (N_22909,N_21942,N_22027);
and U22910 (N_22910,N_21058,N_21121);
or U22911 (N_22911,N_21569,N_22126);
or U22912 (N_22912,N_22448,N_22315);
and U22913 (N_22913,N_21469,N_21286);
xor U22914 (N_22914,N_22112,N_21941);
nor U22915 (N_22915,N_21123,N_21734);
nand U22916 (N_22916,N_22460,N_21117);
nor U22917 (N_22917,N_21740,N_21889);
or U22918 (N_22918,N_22452,N_21794);
xnor U22919 (N_22919,N_22034,N_22250);
and U22920 (N_22920,N_21096,N_21223);
xnor U22921 (N_22921,N_21847,N_21790);
nand U22922 (N_22922,N_21585,N_22229);
or U22923 (N_22923,N_22494,N_22447);
nor U22924 (N_22924,N_21232,N_21277);
and U22925 (N_22925,N_21460,N_21697);
nor U22926 (N_22926,N_21086,N_21488);
and U22927 (N_22927,N_22038,N_21950);
and U22928 (N_22928,N_22478,N_21036);
and U22929 (N_22929,N_22403,N_21489);
and U22930 (N_22930,N_21449,N_21328);
and U22931 (N_22931,N_22118,N_22242);
xor U22932 (N_22932,N_21497,N_21010);
nor U22933 (N_22933,N_21098,N_21038);
nor U22934 (N_22934,N_21495,N_22240);
nor U22935 (N_22935,N_21243,N_22392);
nand U22936 (N_22936,N_22449,N_21817);
and U22937 (N_22937,N_21250,N_21976);
or U22938 (N_22938,N_22394,N_22104);
xor U22939 (N_22939,N_22056,N_22055);
nor U22940 (N_22940,N_21638,N_21118);
nor U22941 (N_22941,N_22189,N_21238);
nand U22942 (N_22942,N_21430,N_21693);
xnor U22943 (N_22943,N_22173,N_21225);
or U22944 (N_22944,N_22267,N_21737);
nand U22945 (N_22945,N_21180,N_21662);
or U22946 (N_22946,N_21436,N_21113);
or U22947 (N_22947,N_22282,N_21850);
xor U22948 (N_22948,N_21471,N_21578);
or U22949 (N_22949,N_22355,N_21766);
or U22950 (N_22950,N_22390,N_22136);
or U22951 (N_22951,N_21517,N_21761);
nand U22952 (N_22952,N_22167,N_21168);
and U22953 (N_22953,N_22144,N_21797);
or U22954 (N_22954,N_22221,N_22397);
xor U22955 (N_22955,N_21145,N_22386);
xor U22956 (N_22956,N_21611,N_21753);
xnor U22957 (N_22957,N_21202,N_21279);
nand U22958 (N_22958,N_22187,N_22465);
and U22959 (N_22959,N_21067,N_21814);
nor U22960 (N_22960,N_21270,N_21266);
nand U22961 (N_22961,N_21983,N_22095);
or U22962 (N_22962,N_21995,N_21815);
nand U22963 (N_22963,N_21506,N_21326);
nor U22964 (N_22964,N_22382,N_22215);
or U22965 (N_22965,N_21389,N_21043);
nor U22966 (N_22966,N_21771,N_21206);
and U22967 (N_22967,N_21149,N_22096);
or U22968 (N_22968,N_21588,N_21529);
or U22969 (N_22969,N_22071,N_21549);
nand U22970 (N_22970,N_21872,N_21157);
nand U22971 (N_22971,N_22468,N_22461);
and U22972 (N_22972,N_22402,N_21350);
and U22973 (N_22973,N_21020,N_21385);
nor U22974 (N_22974,N_21731,N_21099);
nand U22975 (N_22975,N_21452,N_21878);
or U22976 (N_22976,N_22084,N_21527);
nand U22977 (N_22977,N_22438,N_21410);
and U22978 (N_22978,N_21818,N_22307);
nor U22979 (N_22979,N_22333,N_21501);
nor U22980 (N_22980,N_21341,N_21204);
or U22981 (N_22981,N_21917,N_21291);
and U22982 (N_22982,N_21554,N_22271);
nor U22983 (N_22983,N_21864,N_22241);
and U22984 (N_22984,N_22127,N_21837);
xnor U22985 (N_22985,N_21055,N_22060);
nand U22986 (N_22986,N_21082,N_22270);
and U22987 (N_22987,N_21858,N_22480);
xor U22988 (N_22988,N_21709,N_21466);
xor U22989 (N_22989,N_21312,N_22256);
and U22990 (N_22990,N_22285,N_21072);
nor U22991 (N_22991,N_21843,N_21342);
xor U22992 (N_22992,N_21485,N_22421);
and U22993 (N_22993,N_21925,N_21330);
xor U22994 (N_22994,N_22491,N_22062);
or U22995 (N_22995,N_22294,N_21162);
or U22996 (N_22996,N_21724,N_21470);
and U22997 (N_22997,N_22272,N_21186);
nand U22998 (N_22998,N_21502,N_22020);
or U22999 (N_22999,N_22313,N_21156);
xnor U23000 (N_23000,N_22225,N_21079);
and U23001 (N_23001,N_21068,N_22202);
xor U23002 (N_23002,N_21334,N_21748);
xnor U23003 (N_23003,N_21437,N_21838);
nor U23004 (N_23004,N_21800,N_21714);
and U23005 (N_23005,N_21218,N_21556);
or U23006 (N_23006,N_21306,N_22172);
nand U23007 (N_23007,N_21683,N_21480);
and U23008 (N_23008,N_21632,N_21877);
nand U23009 (N_23009,N_22128,N_22008);
xor U23010 (N_23010,N_21625,N_21563);
or U23011 (N_23011,N_21392,N_21685);
or U23012 (N_23012,N_21700,N_22375);
and U23013 (N_23013,N_21061,N_21725);
or U23014 (N_23014,N_22046,N_21546);
and U23015 (N_23015,N_21175,N_22433);
and U23016 (N_23016,N_21763,N_21136);
nor U23017 (N_23017,N_22303,N_21107);
or U23018 (N_23018,N_22446,N_22262);
nand U23019 (N_23019,N_22195,N_22139);
and U23020 (N_23020,N_22405,N_21191);
or U23021 (N_23021,N_21736,N_22209);
nand U23022 (N_23022,N_22328,N_21323);
xnor U23023 (N_23023,N_21770,N_21252);
or U23024 (N_23024,N_21975,N_22429);
or U23025 (N_23025,N_22208,N_21572);
nand U23026 (N_23026,N_21930,N_21652);
or U23027 (N_23027,N_21169,N_22332);
nor U23028 (N_23028,N_21345,N_21577);
or U23029 (N_23029,N_21963,N_22427);
nor U23030 (N_23030,N_21786,N_22160);
nor U23031 (N_23031,N_21906,N_21803);
and U23032 (N_23032,N_21812,N_21729);
xor U23033 (N_23033,N_21231,N_21751);
nand U23034 (N_23034,N_21150,N_21840);
nor U23035 (N_23035,N_21663,N_21021);
nand U23036 (N_23036,N_21884,N_21944);
xor U23037 (N_23037,N_22477,N_21080);
or U23038 (N_23038,N_22273,N_21962);
xnor U23039 (N_23039,N_21346,N_21464);
and U23040 (N_23040,N_21296,N_21159);
and U23041 (N_23041,N_21097,N_21432);
nand U23042 (N_23042,N_21394,N_22483);
nor U23043 (N_23043,N_22203,N_22418);
nand U23044 (N_23044,N_21281,N_21785);
or U23045 (N_23045,N_21679,N_22356);
xor U23046 (N_23046,N_21465,N_21013);
and U23047 (N_23047,N_21571,N_21493);
or U23048 (N_23048,N_22414,N_21673);
xnor U23049 (N_23049,N_22288,N_21029);
nand U23050 (N_23050,N_21090,N_22063);
and U23051 (N_23051,N_21914,N_21048);
and U23052 (N_23052,N_21982,N_21525);
and U23053 (N_23053,N_22252,N_22190);
and U23054 (N_23054,N_22258,N_22059);
nor U23055 (N_23055,N_22044,N_21314);
and U23056 (N_23056,N_21681,N_21866);
nand U23057 (N_23057,N_21284,N_22374);
nand U23058 (N_23058,N_22031,N_21433);
and U23059 (N_23059,N_22453,N_21939);
nor U23060 (N_23060,N_21830,N_22107);
xnor U23061 (N_23061,N_21101,N_22488);
xor U23062 (N_23062,N_21633,N_21741);
or U23063 (N_23063,N_21758,N_21973);
or U23064 (N_23064,N_22471,N_21283);
xor U23065 (N_23065,N_22441,N_21360);
nor U23066 (N_23066,N_21947,N_22078);
or U23067 (N_23067,N_21863,N_22360);
and U23068 (N_23068,N_21649,N_21720);
nand U23069 (N_23069,N_22098,N_22495);
nand U23070 (N_23070,N_21960,N_22105);
and U23071 (N_23071,N_21835,N_22363);
xnor U23072 (N_23072,N_22197,N_21924);
nor U23073 (N_23073,N_21025,N_21743);
and U23074 (N_23074,N_21704,N_22097);
xor U23075 (N_23075,N_22347,N_21677);
xor U23076 (N_23076,N_21798,N_21102);
nor U23077 (N_23077,N_22047,N_21135);
and U23078 (N_23078,N_21265,N_22286);
and U23079 (N_23079,N_22289,N_22401);
nand U23080 (N_23080,N_22192,N_21443);
or U23081 (N_23081,N_22292,N_21887);
nor U23082 (N_23082,N_21388,N_21242);
or U23083 (N_23083,N_21399,N_21510);
or U23084 (N_23084,N_21318,N_22010);
nor U23085 (N_23085,N_22108,N_21033);
and U23086 (N_23086,N_21617,N_21183);
nand U23087 (N_23087,N_22423,N_22193);
and U23088 (N_23088,N_21865,N_21894);
nor U23089 (N_23089,N_22380,N_22012);
xnor U23090 (N_23090,N_22415,N_21116);
nand U23091 (N_23091,N_21237,N_21490);
and U23092 (N_23092,N_21426,N_21775);
or U23093 (N_23093,N_21756,N_21338);
nor U23094 (N_23094,N_22204,N_21905);
or U23095 (N_23095,N_22372,N_22101);
and U23096 (N_23096,N_21195,N_22467);
nand U23097 (N_23097,N_22231,N_21065);
xnor U23098 (N_23098,N_21980,N_22050);
and U23099 (N_23099,N_21023,N_22177);
nor U23100 (N_23100,N_21721,N_22493);
nor U23101 (N_23101,N_22472,N_21087);
or U23102 (N_23102,N_21933,N_22454);
xor U23103 (N_23103,N_22462,N_21137);
nand U23104 (N_23104,N_21666,N_22335);
nand U23105 (N_23105,N_21041,N_21707);
or U23106 (N_23106,N_22264,N_21272);
and U23107 (N_23107,N_21188,N_22351);
xor U23108 (N_23108,N_21161,N_22130);
and U23109 (N_23109,N_21359,N_21727);
or U23110 (N_23110,N_22072,N_21541);
and U23111 (N_23111,N_22216,N_21352);
xnor U23112 (N_23112,N_22455,N_21516);
nand U23113 (N_23113,N_22301,N_21176);
xor U23114 (N_23114,N_21833,N_21251);
or U23115 (N_23115,N_21896,N_21187);
or U23116 (N_23116,N_21141,N_21776);
and U23117 (N_23117,N_22279,N_21813);
nand U23118 (N_23118,N_21205,N_21478);
xor U23119 (N_23119,N_21997,N_21138);
or U23120 (N_23120,N_22185,N_21405);
nor U23121 (N_23121,N_22163,N_21876);
nand U23122 (N_23122,N_21193,N_21645);
or U23123 (N_23123,N_22385,N_21710);
or U23124 (N_23124,N_22251,N_21184);
nor U23125 (N_23125,N_21446,N_21400);
and U23126 (N_23126,N_22100,N_21439);
or U23127 (N_23127,N_22037,N_21515);
xnor U23128 (N_23128,N_21807,N_21083);
nand U23129 (N_23129,N_21333,N_22025);
nor U23130 (N_23130,N_21375,N_21109);
xor U23131 (N_23131,N_22293,N_22244);
nor U23132 (N_23132,N_22153,N_21570);
nor U23133 (N_23133,N_21199,N_21801);
nor U23134 (N_23134,N_21537,N_21051);
xnor U23135 (N_23135,N_21844,N_21604);
nand U23136 (N_23136,N_22399,N_22082);
nand U23137 (N_23137,N_22083,N_21442);
xnor U23138 (N_23138,N_21482,N_22321);
and U23139 (N_23139,N_21158,N_21024);
nand U23140 (N_23140,N_22389,N_21723);
xnor U23141 (N_23141,N_21749,N_21583);
nand U23142 (N_23142,N_21503,N_22274);
or U23143 (N_23143,N_22166,N_21567);
and U23144 (N_23144,N_21892,N_22088);
xnor U23145 (N_23145,N_22263,N_21365);
nor U23146 (N_23146,N_21528,N_21990);
or U23147 (N_23147,N_22473,N_22436);
xor U23148 (N_23148,N_21637,N_22102);
or U23149 (N_23149,N_21222,N_21802);
nor U23150 (N_23150,N_21928,N_21712);
nand U23151 (N_23151,N_22281,N_21643);
xnor U23152 (N_23152,N_22359,N_22113);
xor U23153 (N_23153,N_21883,N_21294);
nand U23154 (N_23154,N_21153,N_21716);
and U23155 (N_23155,N_21855,N_21773);
or U23156 (N_23156,N_22420,N_22497);
xor U23157 (N_23157,N_21902,N_22135);
and U23158 (N_23158,N_21233,N_21401);
or U23159 (N_23159,N_21347,N_21154);
or U23160 (N_23160,N_21660,N_21958);
nand U23161 (N_23161,N_21391,N_21369);
xor U23162 (N_23162,N_21419,N_21726);
nand U23163 (N_23163,N_21203,N_22278);
nand U23164 (N_23164,N_21128,N_21134);
nor U23165 (N_23165,N_21304,N_22408);
or U23166 (N_23166,N_21631,N_21616);
xnor U23167 (N_23167,N_21421,N_22074);
or U23168 (N_23168,N_22443,N_21253);
nand U23169 (N_23169,N_21824,N_21657);
or U23170 (N_23170,N_21413,N_22469);
nor U23171 (N_23171,N_22404,N_21235);
xor U23172 (N_23172,N_21032,N_21094);
nor U23173 (N_23173,N_22316,N_21009);
or U23174 (N_23174,N_21045,N_22206);
nand U23175 (N_23175,N_21558,N_21422);
nand U23176 (N_23176,N_21383,N_21919);
xnor U23177 (N_23177,N_22023,N_21069);
nand U23178 (N_23178,N_21832,N_21006);
nand U23179 (N_23179,N_21142,N_21614);
xor U23180 (N_23180,N_21553,N_21386);
nand U23181 (N_23181,N_21302,N_21031);
nor U23182 (N_23182,N_21192,N_21271);
xor U23183 (N_23183,N_21245,N_22276);
or U23184 (N_23184,N_21444,N_21907);
nor U23185 (N_23185,N_22492,N_21868);
nand U23186 (N_23186,N_21584,N_22176);
xor U23187 (N_23187,N_21046,N_21642);
nand U23188 (N_23188,N_21091,N_21661);
xor U23189 (N_23189,N_21056,N_21574);
nor U23190 (N_23190,N_22223,N_21615);
xnor U23191 (N_23191,N_21739,N_21597);
and U23192 (N_23192,N_22180,N_21853);
nor U23193 (N_23193,N_21173,N_21078);
nand U23194 (N_23194,N_21559,N_21656);
xor U23195 (N_23195,N_21447,N_21988);
nor U23196 (N_23196,N_21886,N_22459);
and U23197 (N_23197,N_22219,N_21970);
and U23198 (N_23198,N_22019,N_22116);
xnor U23199 (N_23199,N_21568,N_21042);
nand U23200 (N_23200,N_21901,N_21810);
nor U23201 (N_23201,N_21779,N_21409);
and U23202 (N_23202,N_22326,N_22249);
xor U23203 (N_23203,N_22309,N_21130);
or U23204 (N_23204,N_21993,N_21044);
nor U23205 (N_23205,N_21403,N_22033);
and U23206 (N_23206,N_22238,N_22341);
xnor U23207 (N_23207,N_22121,N_22061);
nand U23208 (N_23208,N_22070,N_21244);
or U23209 (N_23209,N_21450,N_21462);
or U23210 (N_23210,N_21179,N_22331);
xor U23211 (N_23211,N_21317,N_22198);
or U23212 (N_23212,N_22442,N_21358);
nand U23213 (N_23213,N_22407,N_21016);
xor U23214 (N_23214,N_21100,N_22120);
or U23215 (N_23215,N_22464,N_21605);
or U23216 (N_23216,N_21875,N_21476);
xor U23217 (N_23217,N_21869,N_21792);
xor U23218 (N_23218,N_22422,N_21062);
nor U23219 (N_23219,N_22255,N_21002);
or U23220 (N_23220,N_21669,N_21746);
xor U23221 (N_23221,N_21647,N_21551);
nor U23222 (N_23222,N_21784,N_21052);
or U23223 (N_23223,N_21513,N_21953);
nand U23224 (N_23224,N_21440,N_21108);
or U23225 (N_23225,N_22147,N_21483);
and U23226 (N_23226,N_22268,N_21353);
nand U23227 (N_23227,N_21706,N_21278);
xor U23228 (N_23228,N_21474,N_21954);
nand U23229 (N_23229,N_21670,N_21536);
xor U23230 (N_23230,N_22320,N_21550);
and U23231 (N_23231,N_21336,N_21897);
or U23232 (N_23232,N_21431,N_21039);
nand U23233 (N_23233,N_21613,N_21682);
nor U23234 (N_23234,N_21114,N_21636);
xnor U23235 (N_23235,N_21949,N_22499);
nor U23236 (N_23236,N_22450,N_22437);
or U23237 (N_23237,N_22224,N_21455);
or U23238 (N_23238,N_21165,N_21380);
nor U23239 (N_23239,N_21343,N_22358);
nor U23240 (N_23240,N_22129,N_21001);
nor U23241 (N_23241,N_21127,N_22323);
and U23242 (N_23242,N_21194,N_21793);
and U23243 (N_23243,N_21372,N_21722);
and U23244 (N_23244,N_21971,N_21292);
or U23245 (N_23245,N_21487,N_21823);
nor U23246 (N_23246,N_22451,N_21112);
nor U23247 (N_23247,N_21337,N_21733);
nand U23248 (N_23248,N_22024,N_21796);
and U23249 (N_23249,N_22239,N_21236);
nor U23250 (N_23250,N_21318,N_21140);
xor U23251 (N_23251,N_22431,N_21723);
nand U23252 (N_23252,N_21056,N_21194);
nand U23253 (N_23253,N_21768,N_21188);
nor U23254 (N_23254,N_21906,N_21920);
xor U23255 (N_23255,N_21930,N_21226);
nor U23256 (N_23256,N_21113,N_21205);
nor U23257 (N_23257,N_22236,N_22159);
or U23258 (N_23258,N_21231,N_22080);
and U23259 (N_23259,N_21961,N_22464);
xnor U23260 (N_23260,N_21751,N_22115);
nor U23261 (N_23261,N_21649,N_21686);
xnor U23262 (N_23262,N_22207,N_21637);
nor U23263 (N_23263,N_22445,N_21897);
nand U23264 (N_23264,N_21637,N_21493);
nand U23265 (N_23265,N_21966,N_21222);
nand U23266 (N_23266,N_21899,N_21929);
nor U23267 (N_23267,N_22279,N_22156);
or U23268 (N_23268,N_21897,N_21380);
nor U23269 (N_23269,N_21446,N_21815);
xnor U23270 (N_23270,N_21923,N_22348);
or U23271 (N_23271,N_21661,N_21663);
or U23272 (N_23272,N_22338,N_22416);
nand U23273 (N_23273,N_21871,N_21106);
and U23274 (N_23274,N_21268,N_21350);
or U23275 (N_23275,N_21258,N_21132);
or U23276 (N_23276,N_21388,N_22457);
nor U23277 (N_23277,N_22313,N_21097);
nand U23278 (N_23278,N_21109,N_21330);
nor U23279 (N_23279,N_21953,N_21702);
nand U23280 (N_23280,N_21938,N_21462);
and U23281 (N_23281,N_22098,N_21337);
nand U23282 (N_23282,N_21567,N_21781);
xor U23283 (N_23283,N_21213,N_22147);
xor U23284 (N_23284,N_21236,N_21228);
nand U23285 (N_23285,N_21448,N_21561);
nand U23286 (N_23286,N_21170,N_21386);
nor U23287 (N_23287,N_21742,N_21499);
or U23288 (N_23288,N_22341,N_22170);
and U23289 (N_23289,N_21139,N_22149);
and U23290 (N_23290,N_21707,N_21042);
or U23291 (N_23291,N_21094,N_21914);
and U23292 (N_23292,N_21774,N_21630);
nor U23293 (N_23293,N_21414,N_21624);
nand U23294 (N_23294,N_21204,N_22209);
nand U23295 (N_23295,N_22160,N_22198);
and U23296 (N_23296,N_21641,N_21909);
nand U23297 (N_23297,N_21309,N_22408);
xnor U23298 (N_23298,N_22067,N_22248);
nand U23299 (N_23299,N_21771,N_22406);
and U23300 (N_23300,N_21181,N_21299);
or U23301 (N_23301,N_22087,N_22431);
or U23302 (N_23302,N_22361,N_21696);
and U23303 (N_23303,N_22091,N_21458);
xor U23304 (N_23304,N_22222,N_21605);
nand U23305 (N_23305,N_21107,N_21352);
and U23306 (N_23306,N_22494,N_22139);
or U23307 (N_23307,N_22480,N_21457);
nand U23308 (N_23308,N_21878,N_22415);
and U23309 (N_23309,N_22029,N_21423);
nand U23310 (N_23310,N_22144,N_21429);
nor U23311 (N_23311,N_22082,N_21326);
nand U23312 (N_23312,N_21281,N_21719);
nand U23313 (N_23313,N_22029,N_21361);
or U23314 (N_23314,N_21182,N_22058);
xnor U23315 (N_23315,N_21824,N_21666);
or U23316 (N_23316,N_21890,N_22303);
nor U23317 (N_23317,N_21859,N_22299);
xor U23318 (N_23318,N_21044,N_21255);
or U23319 (N_23319,N_22174,N_21423);
and U23320 (N_23320,N_21653,N_21996);
or U23321 (N_23321,N_22280,N_21257);
or U23322 (N_23322,N_21822,N_22360);
or U23323 (N_23323,N_22315,N_21364);
or U23324 (N_23324,N_21505,N_21873);
or U23325 (N_23325,N_22338,N_22350);
and U23326 (N_23326,N_21457,N_21009);
nor U23327 (N_23327,N_21085,N_21887);
or U23328 (N_23328,N_21798,N_22244);
xnor U23329 (N_23329,N_21193,N_21538);
nor U23330 (N_23330,N_21312,N_21260);
and U23331 (N_23331,N_21762,N_21653);
xor U23332 (N_23332,N_21158,N_21336);
nor U23333 (N_23333,N_21678,N_21978);
nor U23334 (N_23334,N_22243,N_22233);
nand U23335 (N_23335,N_22103,N_21673);
xor U23336 (N_23336,N_21060,N_22241);
nor U23337 (N_23337,N_22071,N_21749);
nor U23338 (N_23338,N_21644,N_22201);
nand U23339 (N_23339,N_21622,N_21663);
and U23340 (N_23340,N_22336,N_21882);
xnor U23341 (N_23341,N_22050,N_22027);
nand U23342 (N_23342,N_22065,N_21177);
and U23343 (N_23343,N_22100,N_21635);
or U23344 (N_23344,N_21715,N_21877);
nor U23345 (N_23345,N_21132,N_22053);
nand U23346 (N_23346,N_22450,N_22250);
xor U23347 (N_23347,N_22108,N_21772);
nor U23348 (N_23348,N_21865,N_22027);
nor U23349 (N_23349,N_21621,N_21017);
nor U23350 (N_23350,N_21022,N_21051);
and U23351 (N_23351,N_21782,N_21200);
nand U23352 (N_23352,N_21563,N_21440);
and U23353 (N_23353,N_21981,N_21127);
or U23354 (N_23354,N_22413,N_22058);
nand U23355 (N_23355,N_22301,N_21953);
or U23356 (N_23356,N_21115,N_22477);
xor U23357 (N_23357,N_21185,N_21686);
or U23358 (N_23358,N_22341,N_21703);
or U23359 (N_23359,N_22043,N_22319);
nand U23360 (N_23360,N_21640,N_21100);
and U23361 (N_23361,N_22001,N_21123);
xnor U23362 (N_23362,N_21688,N_22269);
and U23363 (N_23363,N_21231,N_21408);
xnor U23364 (N_23364,N_21994,N_22257);
nor U23365 (N_23365,N_21370,N_21266);
or U23366 (N_23366,N_21485,N_21393);
or U23367 (N_23367,N_21405,N_22474);
xor U23368 (N_23368,N_21315,N_21985);
nand U23369 (N_23369,N_22269,N_22384);
xnor U23370 (N_23370,N_21555,N_21233);
xor U23371 (N_23371,N_21274,N_21009);
nand U23372 (N_23372,N_22301,N_21781);
or U23373 (N_23373,N_22409,N_21774);
nand U23374 (N_23374,N_22265,N_21291);
and U23375 (N_23375,N_21542,N_22156);
or U23376 (N_23376,N_22493,N_21630);
and U23377 (N_23377,N_21338,N_21519);
and U23378 (N_23378,N_21530,N_22358);
nand U23379 (N_23379,N_22021,N_21265);
xnor U23380 (N_23380,N_22421,N_21797);
xor U23381 (N_23381,N_21509,N_21214);
nand U23382 (N_23382,N_22032,N_21040);
nor U23383 (N_23383,N_21520,N_21327);
nand U23384 (N_23384,N_22043,N_21333);
nand U23385 (N_23385,N_22454,N_22073);
and U23386 (N_23386,N_21257,N_21715);
nand U23387 (N_23387,N_21222,N_22089);
nor U23388 (N_23388,N_21147,N_21583);
xnor U23389 (N_23389,N_21094,N_21831);
nand U23390 (N_23390,N_21442,N_21473);
nand U23391 (N_23391,N_21657,N_21720);
xor U23392 (N_23392,N_21677,N_22099);
nor U23393 (N_23393,N_22072,N_21079);
xor U23394 (N_23394,N_21729,N_21833);
nor U23395 (N_23395,N_21180,N_22244);
or U23396 (N_23396,N_22065,N_21694);
xnor U23397 (N_23397,N_21882,N_21651);
and U23398 (N_23398,N_21501,N_21825);
and U23399 (N_23399,N_22407,N_21983);
or U23400 (N_23400,N_21866,N_22462);
xor U23401 (N_23401,N_21691,N_22350);
nand U23402 (N_23402,N_21832,N_21866);
xnor U23403 (N_23403,N_22126,N_22434);
and U23404 (N_23404,N_21935,N_21957);
nor U23405 (N_23405,N_21457,N_21335);
and U23406 (N_23406,N_21378,N_21863);
nor U23407 (N_23407,N_22021,N_21446);
xor U23408 (N_23408,N_22210,N_21479);
nand U23409 (N_23409,N_21777,N_22173);
nand U23410 (N_23410,N_21072,N_21219);
nand U23411 (N_23411,N_21072,N_21504);
or U23412 (N_23412,N_22351,N_21721);
nor U23413 (N_23413,N_21543,N_21117);
nor U23414 (N_23414,N_21530,N_21513);
or U23415 (N_23415,N_22489,N_21811);
nand U23416 (N_23416,N_21423,N_21345);
or U23417 (N_23417,N_22266,N_21941);
xor U23418 (N_23418,N_22337,N_21727);
and U23419 (N_23419,N_21079,N_21239);
or U23420 (N_23420,N_21012,N_21137);
nor U23421 (N_23421,N_21110,N_22214);
or U23422 (N_23422,N_21293,N_21213);
nor U23423 (N_23423,N_22040,N_21466);
and U23424 (N_23424,N_22047,N_21574);
xnor U23425 (N_23425,N_22263,N_21097);
and U23426 (N_23426,N_21674,N_21276);
nor U23427 (N_23427,N_21352,N_21231);
xnor U23428 (N_23428,N_21658,N_22318);
nand U23429 (N_23429,N_21969,N_22390);
nand U23430 (N_23430,N_21666,N_22195);
nor U23431 (N_23431,N_21838,N_21642);
nor U23432 (N_23432,N_21847,N_21932);
xor U23433 (N_23433,N_22164,N_21394);
or U23434 (N_23434,N_22010,N_21043);
and U23435 (N_23435,N_21711,N_21855);
or U23436 (N_23436,N_21189,N_21845);
nand U23437 (N_23437,N_21317,N_21829);
and U23438 (N_23438,N_21672,N_21230);
xnor U23439 (N_23439,N_22412,N_21633);
nand U23440 (N_23440,N_21975,N_21084);
xor U23441 (N_23441,N_21852,N_22194);
nand U23442 (N_23442,N_22468,N_22474);
or U23443 (N_23443,N_22365,N_21721);
xnor U23444 (N_23444,N_21185,N_21550);
nand U23445 (N_23445,N_21191,N_21041);
or U23446 (N_23446,N_21312,N_21226);
and U23447 (N_23447,N_22395,N_22264);
or U23448 (N_23448,N_21735,N_21340);
and U23449 (N_23449,N_22302,N_21760);
nor U23450 (N_23450,N_21851,N_22355);
or U23451 (N_23451,N_22428,N_21086);
or U23452 (N_23452,N_21682,N_21217);
and U23453 (N_23453,N_21723,N_21528);
xnor U23454 (N_23454,N_21021,N_21508);
nor U23455 (N_23455,N_21423,N_22048);
or U23456 (N_23456,N_21274,N_21364);
or U23457 (N_23457,N_22454,N_21392);
xnor U23458 (N_23458,N_21085,N_22156);
or U23459 (N_23459,N_21930,N_22483);
xnor U23460 (N_23460,N_22461,N_21737);
or U23461 (N_23461,N_21937,N_22042);
xnor U23462 (N_23462,N_21548,N_21494);
or U23463 (N_23463,N_22088,N_21952);
xor U23464 (N_23464,N_22057,N_22408);
nor U23465 (N_23465,N_21685,N_21036);
and U23466 (N_23466,N_21313,N_21591);
xnor U23467 (N_23467,N_21316,N_21584);
and U23468 (N_23468,N_21314,N_21005);
or U23469 (N_23469,N_21088,N_22191);
xor U23470 (N_23470,N_21296,N_21140);
xnor U23471 (N_23471,N_21512,N_21614);
xnor U23472 (N_23472,N_22222,N_21598);
or U23473 (N_23473,N_21431,N_21706);
and U23474 (N_23474,N_21939,N_21429);
nand U23475 (N_23475,N_22311,N_21405);
nand U23476 (N_23476,N_21811,N_21879);
nor U23477 (N_23477,N_21825,N_21784);
nand U23478 (N_23478,N_21825,N_21752);
nand U23479 (N_23479,N_21320,N_21365);
nor U23480 (N_23480,N_22236,N_21145);
nand U23481 (N_23481,N_22079,N_21113);
nand U23482 (N_23482,N_21447,N_22437);
nor U23483 (N_23483,N_22134,N_22128);
xnor U23484 (N_23484,N_21541,N_22486);
xor U23485 (N_23485,N_21316,N_21939);
nand U23486 (N_23486,N_21534,N_22349);
xor U23487 (N_23487,N_22134,N_21757);
xnor U23488 (N_23488,N_21765,N_21853);
nand U23489 (N_23489,N_21684,N_21194);
nor U23490 (N_23490,N_21405,N_22462);
and U23491 (N_23491,N_22234,N_21627);
xor U23492 (N_23492,N_21253,N_22071);
nand U23493 (N_23493,N_22470,N_21434);
nand U23494 (N_23494,N_21801,N_21566);
xnor U23495 (N_23495,N_22329,N_21494);
or U23496 (N_23496,N_22416,N_21437);
nor U23497 (N_23497,N_22187,N_21242);
xnor U23498 (N_23498,N_21652,N_22087);
nor U23499 (N_23499,N_21392,N_21877);
nand U23500 (N_23500,N_21126,N_21836);
nand U23501 (N_23501,N_21627,N_22022);
nor U23502 (N_23502,N_21455,N_21436);
or U23503 (N_23503,N_21685,N_21558);
nand U23504 (N_23504,N_22313,N_22144);
nand U23505 (N_23505,N_22144,N_22080);
nor U23506 (N_23506,N_21008,N_21546);
or U23507 (N_23507,N_21483,N_22277);
and U23508 (N_23508,N_22059,N_21130);
or U23509 (N_23509,N_21137,N_21992);
nand U23510 (N_23510,N_22314,N_22102);
nand U23511 (N_23511,N_22327,N_22128);
xor U23512 (N_23512,N_21145,N_21182);
nand U23513 (N_23513,N_21646,N_21704);
and U23514 (N_23514,N_22336,N_21474);
and U23515 (N_23515,N_21118,N_21799);
or U23516 (N_23516,N_21809,N_22444);
nor U23517 (N_23517,N_21475,N_21864);
xor U23518 (N_23518,N_21681,N_21971);
nor U23519 (N_23519,N_21391,N_21447);
or U23520 (N_23520,N_21486,N_21294);
and U23521 (N_23521,N_21005,N_21070);
nand U23522 (N_23522,N_22477,N_22322);
and U23523 (N_23523,N_21115,N_21756);
nor U23524 (N_23524,N_21634,N_22292);
nor U23525 (N_23525,N_22036,N_21947);
xnor U23526 (N_23526,N_22134,N_21916);
nor U23527 (N_23527,N_22365,N_22063);
xor U23528 (N_23528,N_22043,N_21437);
nand U23529 (N_23529,N_22322,N_22402);
and U23530 (N_23530,N_21133,N_22058);
nand U23531 (N_23531,N_21300,N_21477);
nand U23532 (N_23532,N_21534,N_21706);
or U23533 (N_23533,N_22202,N_21790);
or U23534 (N_23534,N_21068,N_22003);
or U23535 (N_23535,N_21973,N_22184);
nand U23536 (N_23536,N_22429,N_21620);
nand U23537 (N_23537,N_22398,N_21192);
or U23538 (N_23538,N_21986,N_21027);
nand U23539 (N_23539,N_21330,N_21470);
nor U23540 (N_23540,N_21181,N_21706);
xor U23541 (N_23541,N_21842,N_21830);
or U23542 (N_23542,N_21549,N_21706);
xnor U23543 (N_23543,N_22433,N_21753);
xnor U23544 (N_23544,N_21084,N_21173);
or U23545 (N_23545,N_22258,N_21142);
nor U23546 (N_23546,N_22246,N_21423);
xnor U23547 (N_23547,N_21053,N_21024);
xor U23548 (N_23548,N_21297,N_22426);
nand U23549 (N_23549,N_21536,N_21274);
xnor U23550 (N_23550,N_21783,N_22372);
and U23551 (N_23551,N_22033,N_22412);
or U23552 (N_23552,N_22172,N_21444);
and U23553 (N_23553,N_22003,N_21180);
xor U23554 (N_23554,N_21860,N_21935);
or U23555 (N_23555,N_21025,N_22093);
nand U23556 (N_23556,N_22005,N_21707);
and U23557 (N_23557,N_22448,N_21488);
nor U23558 (N_23558,N_21837,N_21525);
xor U23559 (N_23559,N_22245,N_21206);
xor U23560 (N_23560,N_22295,N_21117);
nor U23561 (N_23561,N_22388,N_22448);
nand U23562 (N_23562,N_22499,N_21785);
or U23563 (N_23563,N_21493,N_22466);
nor U23564 (N_23564,N_21072,N_22315);
nand U23565 (N_23565,N_21179,N_21338);
and U23566 (N_23566,N_21610,N_21640);
and U23567 (N_23567,N_21658,N_21408);
and U23568 (N_23568,N_21813,N_21313);
xnor U23569 (N_23569,N_21909,N_22073);
and U23570 (N_23570,N_21835,N_21074);
and U23571 (N_23571,N_21863,N_22480);
xor U23572 (N_23572,N_21086,N_21628);
and U23573 (N_23573,N_21078,N_22356);
or U23574 (N_23574,N_22487,N_21711);
nand U23575 (N_23575,N_21464,N_21066);
or U23576 (N_23576,N_21016,N_21219);
or U23577 (N_23577,N_21831,N_21412);
and U23578 (N_23578,N_22184,N_21871);
or U23579 (N_23579,N_22180,N_21225);
xor U23580 (N_23580,N_22346,N_22001);
nor U23581 (N_23581,N_21612,N_21061);
nand U23582 (N_23582,N_21892,N_21960);
or U23583 (N_23583,N_21699,N_21342);
or U23584 (N_23584,N_21328,N_21078);
xor U23585 (N_23585,N_22358,N_21408);
nor U23586 (N_23586,N_21060,N_22380);
nand U23587 (N_23587,N_22386,N_21027);
xor U23588 (N_23588,N_22223,N_21197);
and U23589 (N_23589,N_21428,N_21341);
xor U23590 (N_23590,N_22232,N_21814);
xnor U23591 (N_23591,N_21566,N_21446);
nor U23592 (N_23592,N_22324,N_21764);
nand U23593 (N_23593,N_21927,N_22330);
nand U23594 (N_23594,N_22069,N_21461);
nand U23595 (N_23595,N_21059,N_21543);
xnor U23596 (N_23596,N_22495,N_21663);
nand U23597 (N_23597,N_22017,N_22090);
and U23598 (N_23598,N_22205,N_21432);
nor U23599 (N_23599,N_21501,N_21759);
nand U23600 (N_23600,N_21959,N_22177);
xnor U23601 (N_23601,N_22290,N_21715);
nand U23602 (N_23602,N_22448,N_22105);
xor U23603 (N_23603,N_21957,N_21305);
nand U23604 (N_23604,N_22426,N_21689);
nand U23605 (N_23605,N_21291,N_22206);
nand U23606 (N_23606,N_21224,N_21843);
or U23607 (N_23607,N_22181,N_21511);
xnor U23608 (N_23608,N_21144,N_21891);
and U23609 (N_23609,N_21540,N_21242);
and U23610 (N_23610,N_21202,N_21929);
xor U23611 (N_23611,N_21052,N_21098);
nand U23612 (N_23612,N_22201,N_21783);
nand U23613 (N_23613,N_22474,N_22247);
xnor U23614 (N_23614,N_21282,N_21040);
or U23615 (N_23615,N_21665,N_22206);
nor U23616 (N_23616,N_21017,N_21147);
or U23617 (N_23617,N_21043,N_21170);
nand U23618 (N_23618,N_21615,N_21080);
nor U23619 (N_23619,N_21558,N_22497);
or U23620 (N_23620,N_21209,N_21082);
nor U23621 (N_23621,N_21743,N_22393);
xnor U23622 (N_23622,N_21225,N_21298);
or U23623 (N_23623,N_21266,N_22027);
and U23624 (N_23624,N_21752,N_21808);
or U23625 (N_23625,N_21513,N_21771);
and U23626 (N_23626,N_21582,N_21816);
or U23627 (N_23627,N_22310,N_21249);
and U23628 (N_23628,N_21570,N_21827);
nor U23629 (N_23629,N_21377,N_21223);
xor U23630 (N_23630,N_21139,N_21143);
nand U23631 (N_23631,N_21859,N_22398);
xnor U23632 (N_23632,N_21750,N_21199);
or U23633 (N_23633,N_22272,N_22142);
nor U23634 (N_23634,N_21285,N_21711);
nor U23635 (N_23635,N_22488,N_21558);
or U23636 (N_23636,N_21676,N_21981);
nor U23637 (N_23637,N_21316,N_21946);
xor U23638 (N_23638,N_21201,N_21369);
nor U23639 (N_23639,N_21632,N_21068);
nand U23640 (N_23640,N_21405,N_21044);
nand U23641 (N_23641,N_22162,N_21942);
or U23642 (N_23642,N_21038,N_21881);
and U23643 (N_23643,N_22470,N_21528);
xor U23644 (N_23644,N_21537,N_21667);
and U23645 (N_23645,N_21552,N_22394);
xnor U23646 (N_23646,N_21501,N_21916);
or U23647 (N_23647,N_21546,N_21730);
nor U23648 (N_23648,N_22158,N_21064);
xor U23649 (N_23649,N_22152,N_21492);
and U23650 (N_23650,N_22496,N_22015);
xor U23651 (N_23651,N_21210,N_22288);
nor U23652 (N_23652,N_21092,N_21139);
and U23653 (N_23653,N_21042,N_21457);
nor U23654 (N_23654,N_21491,N_22205);
or U23655 (N_23655,N_21926,N_21661);
and U23656 (N_23656,N_21867,N_21136);
xnor U23657 (N_23657,N_21184,N_21959);
xor U23658 (N_23658,N_22122,N_22351);
nor U23659 (N_23659,N_21357,N_21792);
nor U23660 (N_23660,N_21073,N_22463);
xnor U23661 (N_23661,N_21293,N_22062);
and U23662 (N_23662,N_21265,N_21129);
or U23663 (N_23663,N_21522,N_21523);
xor U23664 (N_23664,N_21242,N_21346);
and U23665 (N_23665,N_21736,N_22161);
or U23666 (N_23666,N_22296,N_22415);
and U23667 (N_23667,N_21183,N_21256);
and U23668 (N_23668,N_22348,N_21536);
nand U23669 (N_23669,N_21565,N_21681);
or U23670 (N_23670,N_22407,N_22366);
and U23671 (N_23671,N_21252,N_21777);
nand U23672 (N_23672,N_22445,N_22408);
and U23673 (N_23673,N_21772,N_22398);
xor U23674 (N_23674,N_21866,N_21121);
xnor U23675 (N_23675,N_21897,N_22057);
nand U23676 (N_23676,N_21918,N_21570);
or U23677 (N_23677,N_22390,N_22056);
xor U23678 (N_23678,N_21214,N_21464);
or U23679 (N_23679,N_21493,N_21369);
xnor U23680 (N_23680,N_21413,N_21356);
nor U23681 (N_23681,N_21624,N_22283);
and U23682 (N_23682,N_21788,N_21158);
nor U23683 (N_23683,N_22169,N_22357);
nand U23684 (N_23684,N_21841,N_21295);
and U23685 (N_23685,N_21942,N_22323);
and U23686 (N_23686,N_22020,N_21569);
nand U23687 (N_23687,N_21493,N_22493);
xnor U23688 (N_23688,N_21932,N_21317);
and U23689 (N_23689,N_22171,N_21403);
and U23690 (N_23690,N_22264,N_21299);
and U23691 (N_23691,N_21924,N_22115);
nand U23692 (N_23692,N_21929,N_21463);
nor U23693 (N_23693,N_21003,N_21815);
nand U23694 (N_23694,N_22159,N_22140);
nand U23695 (N_23695,N_22443,N_21787);
and U23696 (N_23696,N_22332,N_21465);
nand U23697 (N_23697,N_21731,N_21790);
and U23698 (N_23698,N_21388,N_21279);
or U23699 (N_23699,N_21816,N_22212);
xnor U23700 (N_23700,N_22055,N_22369);
xor U23701 (N_23701,N_22449,N_22203);
xor U23702 (N_23702,N_22284,N_22159);
nor U23703 (N_23703,N_21521,N_21349);
or U23704 (N_23704,N_21884,N_21710);
nor U23705 (N_23705,N_21030,N_21905);
nor U23706 (N_23706,N_21968,N_21782);
nand U23707 (N_23707,N_22238,N_22076);
nand U23708 (N_23708,N_21930,N_21221);
and U23709 (N_23709,N_21943,N_22177);
or U23710 (N_23710,N_21047,N_22186);
xnor U23711 (N_23711,N_21763,N_21142);
or U23712 (N_23712,N_21129,N_21238);
nand U23713 (N_23713,N_22214,N_22315);
and U23714 (N_23714,N_21621,N_22264);
or U23715 (N_23715,N_21637,N_21670);
or U23716 (N_23716,N_22299,N_21325);
or U23717 (N_23717,N_22129,N_21796);
xnor U23718 (N_23718,N_21494,N_21710);
or U23719 (N_23719,N_22373,N_22303);
xor U23720 (N_23720,N_21461,N_21902);
xnor U23721 (N_23721,N_21351,N_21139);
nor U23722 (N_23722,N_21110,N_22324);
xor U23723 (N_23723,N_21938,N_21186);
or U23724 (N_23724,N_21736,N_21360);
xor U23725 (N_23725,N_21262,N_22206);
or U23726 (N_23726,N_21211,N_21269);
nor U23727 (N_23727,N_21567,N_21391);
or U23728 (N_23728,N_21494,N_21603);
xnor U23729 (N_23729,N_21619,N_22473);
nor U23730 (N_23730,N_21311,N_21508);
xnor U23731 (N_23731,N_21541,N_21133);
and U23732 (N_23732,N_21531,N_22094);
or U23733 (N_23733,N_21091,N_21573);
nand U23734 (N_23734,N_22081,N_22394);
and U23735 (N_23735,N_22455,N_21154);
nand U23736 (N_23736,N_21504,N_21495);
or U23737 (N_23737,N_22295,N_22176);
nand U23738 (N_23738,N_21191,N_22049);
nand U23739 (N_23739,N_21727,N_22052);
or U23740 (N_23740,N_21599,N_21501);
and U23741 (N_23741,N_22341,N_22475);
nand U23742 (N_23742,N_21506,N_22450);
and U23743 (N_23743,N_21770,N_21138);
xor U23744 (N_23744,N_21289,N_21245);
nand U23745 (N_23745,N_21442,N_21208);
nor U23746 (N_23746,N_21305,N_21186);
nor U23747 (N_23747,N_21494,N_21168);
or U23748 (N_23748,N_22005,N_22211);
xor U23749 (N_23749,N_21555,N_21628);
and U23750 (N_23750,N_21709,N_21791);
nor U23751 (N_23751,N_21295,N_21953);
and U23752 (N_23752,N_22019,N_21351);
nor U23753 (N_23753,N_21391,N_21241);
nand U23754 (N_23754,N_21358,N_21341);
or U23755 (N_23755,N_22331,N_21005);
nor U23756 (N_23756,N_22052,N_22415);
nor U23757 (N_23757,N_22182,N_21058);
xnor U23758 (N_23758,N_22291,N_21357);
nor U23759 (N_23759,N_22057,N_21330);
or U23760 (N_23760,N_21281,N_21716);
nand U23761 (N_23761,N_21609,N_21396);
and U23762 (N_23762,N_21440,N_21179);
nor U23763 (N_23763,N_21070,N_21159);
or U23764 (N_23764,N_21292,N_21437);
nor U23765 (N_23765,N_21317,N_22395);
xor U23766 (N_23766,N_21411,N_22171);
or U23767 (N_23767,N_22223,N_21374);
or U23768 (N_23768,N_21610,N_22096);
or U23769 (N_23769,N_21535,N_21992);
nand U23770 (N_23770,N_21173,N_21182);
nor U23771 (N_23771,N_21049,N_21895);
xnor U23772 (N_23772,N_21809,N_22462);
and U23773 (N_23773,N_21272,N_22388);
nand U23774 (N_23774,N_21024,N_22105);
and U23775 (N_23775,N_22199,N_22347);
nor U23776 (N_23776,N_21982,N_22175);
nand U23777 (N_23777,N_22190,N_21034);
and U23778 (N_23778,N_21220,N_21916);
and U23779 (N_23779,N_22115,N_21060);
or U23780 (N_23780,N_22361,N_21204);
and U23781 (N_23781,N_21858,N_22048);
nand U23782 (N_23782,N_21181,N_21764);
xnor U23783 (N_23783,N_21165,N_22243);
nor U23784 (N_23784,N_22358,N_22050);
or U23785 (N_23785,N_21567,N_21706);
xnor U23786 (N_23786,N_21685,N_21511);
xor U23787 (N_23787,N_21827,N_22403);
nand U23788 (N_23788,N_21684,N_22358);
nand U23789 (N_23789,N_21570,N_21145);
and U23790 (N_23790,N_22085,N_22228);
and U23791 (N_23791,N_21301,N_21219);
xor U23792 (N_23792,N_21803,N_21707);
nand U23793 (N_23793,N_22363,N_21945);
and U23794 (N_23794,N_21252,N_21507);
nor U23795 (N_23795,N_21204,N_22488);
and U23796 (N_23796,N_21027,N_22442);
or U23797 (N_23797,N_21244,N_21299);
or U23798 (N_23798,N_22499,N_22038);
xor U23799 (N_23799,N_21750,N_21230);
xor U23800 (N_23800,N_21218,N_22454);
and U23801 (N_23801,N_22343,N_22165);
or U23802 (N_23802,N_21407,N_21019);
or U23803 (N_23803,N_21561,N_21602);
xor U23804 (N_23804,N_21085,N_21922);
xnor U23805 (N_23805,N_21383,N_21089);
and U23806 (N_23806,N_21502,N_21927);
nand U23807 (N_23807,N_21139,N_21787);
nor U23808 (N_23808,N_21601,N_22335);
nor U23809 (N_23809,N_21032,N_22036);
or U23810 (N_23810,N_21898,N_21965);
and U23811 (N_23811,N_21571,N_21710);
nand U23812 (N_23812,N_21375,N_21111);
xor U23813 (N_23813,N_21769,N_21140);
nand U23814 (N_23814,N_22415,N_22241);
xnor U23815 (N_23815,N_21027,N_22464);
nor U23816 (N_23816,N_21000,N_21338);
and U23817 (N_23817,N_21972,N_21246);
and U23818 (N_23818,N_22170,N_22498);
or U23819 (N_23819,N_21671,N_21058);
or U23820 (N_23820,N_21438,N_21397);
xnor U23821 (N_23821,N_22499,N_21082);
xnor U23822 (N_23822,N_22169,N_22157);
xnor U23823 (N_23823,N_21543,N_22210);
and U23824 (N_23824,N_22138,N_21636);
nand U23825 (N_23825,N_21121,N_21756);
nand U23826 (N_23826,N_22450,N_21527);
nor U23827 (N_23827,N_21952,N_22034);
and U23828 (N_23828,N_21623,N_22373);
and U23829 (N_23829,N_21698,N_21525);
xor U23830 (N_23830,N_22066,N_21149);
nor U23831 (N_23831,N_22303,N_22032);
nand U23832 (N_23832,N_21706,N_21210);
xor U23833 (N_23833,N_21108,N_22442);
nor U23834 (N_23834,N_21025,N_21437);
and U23835 (N_23835,N_21897,N_21886);
nor U23836 (N_23836,N_21383,N_21916);
nand U23837 (N_23837,N_22405,N_22146);
nor U23838 (N_23838,N_21674,N_21236);
and U23839 (N_23839,N_22155,N_22427);
and U23840 (N_23840,N_21980,N_22009);
nand U23841 (N_23841,N_21100,N_21283);
or U23842 (N_23842,N_21865,N_21361);
and U23843 (N_23843,N_22085,N_21474);
nor U23844 (N_23844,N_21837,N_21445);
nand U23845 (N_23845,N_21501,N_21888);
nand U23846 (N_23846,N_22079,N_22085);
and U23847 (N_23847,N_21175,N_22109);
and U23848 (N_23848,N_22162,N_22326);
and U23849 (N_23849,N_22230,N_22392);
and U23850 (N_23850,N_21509,N_22243);
or U23851 (N_23851,N_21413,N_21575);
nor U23852 (N_23852,N_22165,N_22154);
nand U23853 (N_23853,N_22309,N_22038);
nand U23854 (N_23854,N_21154,N_21036);
xor U23855 (N_23855,N_21413,N_21747);
and U23856 (N_23856,N_22148,N_22383);
xnor U23857 (N_23857,N_22011,N_21277);
nand U23858 (N_23858,N_21227,N_21202);
nor U23859 (N_23859,N_22277,N_21525);
xor U23860 (N_23860,N_22326,N_21969);
nor U23861 (N_23861,N_21322,N_22156);
and U23862 (N_23862,N_22019,N_21571);
xnor U23863 (N_23863,N_21965,N_21045);
nor U23864 (N_23864,N_21461,N_21170);
and U23865 (N_23865,N_21982,N_21929);
nor U23866 (N_23866,N_22404,N_21398);
and U23867 (N_23867,N_22317,N_21418);
nand U23868 (N_23868,N_22012,N_22350);
xnor U23869 (N_23869,N_21272,N_22398);
or U23870 (N_23870,N_21935,N_21220);
nand U23871 (N_23871,N_21441,N_21176);
or U23872 (N_23872,N_22480,N_21273);
nand U23873 (N_23873,N_22072,N_21840);
or U23874 (N_23874,N_22253,N_21544);
nand U23875 (N_23875,N_21838,N_21471);
nand U23876 (N_23876,N_22398,N_22392);
or U23877 (N_23877,N_21881,N_21187);
nand U23878 (N_23878,N_21448,N_22346);
nor U23879 (N_23879,N_21714,N_21258);
xnor U23880 (N_23880,N_21579,N_22116);
xnor U23881 (N_23881,N_21759,N_21215);
xor U23882 (N_23882,N_21533,N_21570);
or U23883 (N_23883,N_21876,N_22357);
nor U23884 (N_23884,N_22197,N_21884);
xor U23885 (N_23885,N_21805,N_21531);
xor U23886 (N_23886,N_21736,N_21431);
xnor U23887 (N_23887,N_21453,N_22054);
xor U23888 (N_23888,N_21125,N_22192);
nand U23889 (N_23889,N_22426,N_21959);
xnor U23890 (N_23890,N_22487,N_21511);
and U23891 (N_23891,N_21915,N_22427);
nor U23892 (N_23892,N_21200,N_22173);
and U23893 (N_23893,N_22484,N_22110);
nor U23894 (N_23894,N_22141,N_21963);
nor U23895 (N_23895,N_21899,N_21973);
xnor U23896 (N_23896,N_21271,N_21414);
nor U23897 (N_23897,N_21865,N_21397);
nand U23898 (N_23898,N_22104,N_22033);
nand U23899 (N_23899,N_21209,N_22031);
nand U23900 (N_23900,N_22136,N_21036);
xnor U23901 (N_23901,N_21538,N_21548);
xor U23902 (N_23902,N_22338,N_22257);
nor U23903 (N_23903,N_22264,N_22055);
nor U23904 (N_23904,N_21746,N_22013);
or U23905 (N_23905,N_21592,N_22200);
or U23906 (N_23906,N_22007,N_21332);
nand U23907 (N_23907,N_21559,N_22339);
nor U23908 (N_23908,N_21021,N_22338);
nand U23909 (N_23909,N_21107,N_22074);
xnor U23910 (N_23910,N_21048,N_21168);
nor U23911 (N_23911,N_21018,N_21084);
nand U23912 (N_23912,N_22090,N_21127);
or U23913 (N_23913,N_22423,N_22311);
or U23914 (N_23914,N_22327,N_22236);
nor U23915 (N_23915,N_22010,N_22168);
nor U23916 (N_23916,N_21167,N_21890);
or U23917 (N_23917,N_21733,N_22389);
nor U23918 (N_23918,N_21092,N_22005);
and U23919 (N_23919,N_22116,N_21038);
nor U23920 (N_23920,N_21013,N_21846);
and U23921 (N_23921,N_21492,N_22151);
nand U23922 (N_23922,N_22407,N_22185);
nand U23923 (N_23923,N_21319,N_21896);
xnor U23924 (N_23924,N_21607,N_22135);
or U23925 (N_23925,N_22499,N_21148);
or U23926 (N_23926,N_21357,N_21824);
and U23927 (N_23927,N_21505,N_22028);
xor U23928 (N_23928,N_21147,N_21526);
and U23929 (N_23929,N_22419,N_22382);
nand U23930 (N_23930,N_21426,N_22124);
nand U23931 (N_23931,N_22389,N_21206);
nor U23932 (N_23932,N_21976,N_21135);
nor U23933 (N_23933,N_22289,N_22147);
nand U23934 (N_23934,N_22472,N_22031);
nand U23935 (N_23935,N_22465,N_21975);
xor U23936 (N_23936,N_21248,N_22015);
xor U23937 (N_23937,N_21922,N_21546);
xnor U23938 (N_23938,N_22389,N_22238);
and U23939 (N_23939,N_21028,N_22291);
or U23940 (N_23940,N_21755,N_22030);
nand U23941 (N_23941,N_21884,N_21432);
or U23942 (N_23942,N_21100,N_21988);
nand U23943 (N_23943,N_21269,N_22103);
xnor U23944 (N_23944,N_22385,N_22293);
or U23945 (N_23945,N_21113,N_22408);
nor U23946 (N_23946,N_22366,N_22241);
or U23947 (N_23947,N_21626,N_22445);
and U23948 (N_23948,N_22221,N_21888);
nand U23949 (N_23949,N_21346,N_21421);
xor U23950 (N_23950,N_21377,N_22204);
or U23951 (N_23951,N_21835,N_22066);
or U23952 (N_23952,N_21243,N_21317);
and U23953 (N_23953,N_21043,N_22252);
or U23954 (N_23954,N_21614,N_21434);
and U23955 (N_23955,N_21112,N_21538);
xnor U23956 (N_23956,N_21734,N_21466);
and U23957 (N_23957,N_22052,N_21858);
nand U23958 (N_23958,N_22050,N_21583);
xnor U23959 (N_23959,N_22490,N_22123);
xor U23960 (N_23960,N_22151,N_21107);
and U23961 (N_23961,N_21011,N_21646);
xor U23962 (N_23962,N_21804,N_22479);
nor U23963 (N_23963,N_21256,N_21965);
nand U23964 (N_23964,N_22046,N_21931);
nor U23965 (N_23965,N_21680,N_21393);
and U23966 (N_23966,N_21003,N_22477);
nor U23967 (N_23967,N_21871,N_22283);
nand U23968 (N_23968,N_22059,N_21870);
xor U23969 (N_23969,N_21886,N_21020);
nor U23970 (N_23970,N_21083,N_21642);
xnor U23971 (N_23971,N_22256,N_21638);
xnor U23972 (N_23972,N_21985,N_21712);
or U23973 (N_23973,N_21317,N_21605);
xor U23974 (N_23974,N_21806,N_22149);
nor U23975 (N_23975,N_21248,N_22073);
nor U23976 (N_23976,N_21025,N_22457);
nand U23977 (N_23977,N_21411,N_21731);
and U23978 (N_23978,N_22061,N_22334);
nand U23979 (N_23979,N_21933,N_22430);
nor U23980 (N_23980,N_21887,N_22154);
and U23981 (N_23981,N_21538,N_22254);
nor U23982 (N_23982,N_22071,N_22293);
nor U23983 (N_23983,N_21801,N_21596);
nor U23984 (N_23984,N_22380,N_22331);
xnor U23985 (N_23985,N_21945,N_21354);
nor U23986 (N_23986,N_21972,N_21479);
nor U23987 (N_23987,N_22442,N_21944);
nand U23988 (N_23988,N_21380,N_21163);
nand U23989 (N_23989,N_21581,N_21686);
nand U23990 (N_23990,N_21507,N_21272);
or U23991 (N_23991,N_21393,N_22072);
xnor U23992 (N_23992,N_21004,N_21416);
nor U23993 (N_23993,N_21575,N_21018);
nor U23994 (N_23994,N_21362,N_22419);
or U23995 (N_23995,N_21801,N_21095);
and U23996 (N_23996,N_21540,N_21515);
and U23997 (N_23997,N_21704,N_22192);
and U23998 (N_23998,N_21188,N_21349);
and U23999 (N_23999,N_21759,N_21838);
xnor U24000 (N_24000,N_23029,N_23850);
xor U24001 (N_24001,N_23962,N_23133);
nand U24002 (N_24002,N_23307,N_22597);
and U24003 (N_24003,N_22984,N_23628);
or U24004 (N_24004,N_22588,N_23811);
nor U24005 (N_24005,N_22853,N_22961);
nand U24006 (N_24006,N_23641,N_22725);
and U24007 (N_24007,N_23639,N_23555);
and U24008 (N_24008,N_23214,N_23827);
or U24009 (N_24009,N_23763,N_23288);
and U24010 (N_24010,N_22920,N_22932);
and U24011 (N_24011,N_22598,N_23551);
and U24012 (N_24012,N_23670,N_22902);
nand U24013 (N_24013,N_23908,N_23479);
or U24014 (N_24014,N_22560,N_23729);
or U24015 (N_24015,N_22757,N_23887);
nand U24016 (N_24016,N_23566,N_22847);
nand U24017 (N_24017,N_23971,N_22618);
nand U24018 (N_24018,N_23302,N_22651);
or U24019 (N_24019,N_23078,N_23810);
and U24020 (N_24020,N_23535,N_22698);
or U24021 (N_24021,N_23591,N_23070);
and U24022 (N_24022,N_22604,N_23043);
nor U24023 (N_24023,N_23859,N_22953);
or U24024 (N_24024,N_23634,N_23703);
or U24025 (N_24025,N_23538,N_22811);
and U24026 (N_24026,N_23780,N_23685);
and U24027 (N_24027,N_23212,N_23734);
or U24028 (N_24028,N_23612,N_23171);
xnor U24029 (N_24029,N_22638,N_23032);
nor U24030 (N_24030,N_23438,N_23477);
or U24031 (N_24031,N_23838,N_23167);
or U24032 (N_24032,N_23650,N_23161);
nand U24033 (N_24033,N_23320,N_23107);
nand U24034 (N_24034,N_23226,N_22599);
xnor U24035 (N_24035,N_23541,N_23829);
nand U24036 (N_24036,N_23943,N_22855);
nor U24037 (N_24037,N_22892,N_23697);
and U24038 (N_24038,N_22985,N_23651);
xor U24039 (N_24039,N_23820,N_22515);
nand U24040 (N_24040,N_22539,N_22772);
nor U24041 (N_24041,N_23385,N_23751);
nor U24042 (N_24042,N_22843,N_22538);
or U24043 (N_24043,N_23286,N_22529);
and U24044 (N_24044,N_23548,N_23278);
xor U24045 (N_24045,N_22729,N_23809);
nor U24046 (N_24046,N_23244,N_23946);
nand U24047 (N_24047,N_22986,N_23969);
nand U24048 (N_24048,N_23353,N_23545);
nor U24049 (N_24049,N_23679,N_22681);
xnor U24050 (N_24050,N_22754,N_22937);
nor U24051 (N_24051,N_22643,N_23778);
xor U24052 (N_24052,N_23276,N_23457);
or U24053 (N_24053,N_23413,N_23414);
or U24054 (N_24054,N_22886,N_23588);
or U24055 (N_24055,N_23877,N_23916);
and U24056 (N_24056,N_23681,N_23671);
nand U24057 (N_24057,N_23382,N_22722);
and U24058 (N_24058,N_23439,N_23303);
or U24059 (N_24059,N_22590,N_22734);
nor U24060 (N_24060,N_23726,N_22871);
and U24061 (N_24061,N_23243,N_23649);
and U24062 (N_24062,N_23567,N_23259);
nand U24063 (N_24063,N_23949,N_23915);
and U24064 (N_24064,N_22827,N_22600);
and U24065 (N_24065,N_23404,N_22688);
nor U24066 (N_24066,N_23098,N_22756);
nor U24067 (N_24067,N_23415,N_23062);
and U24068 (N_24068,N_23507,N_22851);
nand U24069 (N_24069,N_22607,N_23396);
and U24070 (N_24070,N_22662,N_23981);
or U24071 (N_24071,N_22728,N_22894);
xor U24072 (N_24072,N_22965,N_22803);
nor U24073 (N_24073,N_23722,N_23909);
and U24074 (N_24074,N_23818,N_23669);
or U24075 (N_24075,N_23749,N_23356);
nand U24076 (N_24076,N_23633,N_23805);
nor U24077 (N_24077,N_23732,N_22969);
and U24078 (N_24078,N_23448,N_22667);
nor U24079 (N_24079,N_23550,N_23026);
or U24080 (N_24080,N_22699,N_23883);
nand U24081 (N_24081,N_22925,N_22812);
nor U24082 (N_24082,N_23018,N_23322);
nand U24083 (N_24083,N_23424,N_23505);
xnor U24084 (N_24084,N_22720,N_23088);
nand U24085 (N_24085,N_23642,N_23592);
xor U24086 (N_24086,N_22747,N_23035);
nand U24087 (N_24087,N_23761,N_23084);
nand U24088 (N_24088,N_23125,N_22613);
xor U24089 (N_24089,N_23123,N_23512);
and U24090 (N_24090,N_23436,N_23624);
or U24091 (N_24091,N_22779,N_23037);
and U24092 (N_24092,N_23155,N_23766);
nor U24093 (N_24093,N_23991,N_23914);
nor U24094 (N_24094,N_22594,N_22608);
or U24095 (N_24095,N_23713,N_23750);
xor U24096 (N_24096,N_23179,N_23926);
nand U24097 (N_24097,N_22556,N_23400);
and U24098 (N_24098,N_23597,N_23611);
and U24099 (N_24099,N_23274,N_22610);
nand U24100 (N_24100,N_23998,N_23019);
or U24101 (N_24101,N_22629,N_23851);
nand U24102 (N_24102,N_23701,N_22842);
and U24103 (N_24103,N_22702,N_23562);
and U24104 (N_24104,N_22921,N_23573);
and U24105 (N_24105,N_23565,N_23475);
nand U24106 (N_24106,N_23618,N_22806);
and U24107 (N_24107,N_22758,N_23326);
nand U24108 (N_24108,N_23379,N_23518);
or U24109 (N_24109,N_23373,N_22506);
and U24110 (N_24110,N_23406,N_23557);
nand U24111 (N_24111,N_22861,N_23483);
or U24112 (N_24112,N_23896,N_23452);
and U24113 (N_24113,N_22958,N_22791);
nand U24114 (N_24114,N_23394,N_23901);
xor U24115 (N_24115,N_23773,N_23849);
xnor U24116 (N_24116,N_22577,N_22711);
nand U24117 (N_24117,N_23783,N_23100);
xnor U24118 (N_24118,N_23159,N_23271);
xnor U24119 (N_24119,N_23246,N_22879);
or U24120 (N_24120,N_23927,N_22971);
or U24121 (N_24121,N_22573,N_22690);
and U24122 (N_24122,N_23339,N_23637);
xor U24123 (N_24123,N_22963,N_23707);
nor U24124 (N_24124,N_22752,N_23038);
and U24125 (N_24125,N_23273,N_22907);
nand U24126 (N_24126,N_22676,N_22586);
and U24127 (N_24127,N_22605,N_23407);
xor U24128 (N_24128,N_23210,N_22959);
and U24129 (N_24129,N_22947,N_23539);
nand U24130 (N_24130,N_23529,N_23644);
nor U24131 (N_24131,N_23886,N_23963);
xor U24132 (N_24132,N_23925,N_23229);
or U24133 (N_24133,N_23769,N_23245);
or U24134 (N_24134,N_23675,N_23635);
nor U24135 (N_24135,N_22825,N_23081);
or U24136 (N_24136,N_22622,N_23022);
xor U24137 (N_24137,N_23762,N_22889);
xor U24138 (N_24138,N_23678,N_23305);
xor U24139 (N_24139,N_23623,N_23420);
and U24140 (N_24140,N_23145,N_23281);
nand U24141 (N_24141,N_23711,N_23103);
or U24142 (N_24142,N_22555,N_23940);
or U24143 (N_24143,N_22708,N_23499);
nor U24144 (N_24144,N_22991,N_22578);
or U24145 (N_24145,N_23702,N_23387);
or U24146 (N_24146,N_23324,N_23252);
nand U24147 (N_24147,N_23461,N_23730);
and U24148 (N_24148,N_22931,N_23298);
nand U24149 (N_24149,N_23710,N_22521);
xor U24150 (N_24150,N_23426,N_22735);
xnor U24151 (N_24151,N_22761,N_23254);
or U24152 (N_24152,N_23073,N_23453);
or U24153 (N_24153,N_23357,N_22888);
nor U24154 (N_24154,N_23826,N_23282);
and U24155 (N_24155,N_23606,N_23141);
xnor U24156 (N_24156,N_23277,N_23012);
nor U24157 (N_24157,N_23848,N_22798);
and U24158 (N_24158,N_22505,N_22763);
nand U24159 (N_24159,N_23176,N_23525);
or U24160 (N_24160,N_23837,N_22621);
xnor U24161 (N_24161,N_23640,N_23304);
and U24162 (N_24162,N_22983,N_23542);
nor U24163 (N_24163,N_23131,N_23777);
xor U24164 (N_24164,N_23972,N_23311);
or U24165 (N_24165,N_22684,N_22721);
nor U24166 (N_24166,N_23690,N_23348);
and U24167 (N_24167,N_23884,N_22956);
nor U24168 (N_24168,N_22541,N_22949);
xnor U24169 (N_24169,N_22609,N_23262);
nand U24170 (N_24170,N_22778,N_23636);
nand U24171 (N_24171,N_23048,N_22633);
nor U24172 (N_24172,N_23683,N_22703);
xor U24173 (N_24173,N_23359,N_23920);
nor U24174 (N_24174,N_23197,N_23417);
xor U24175 (N_24175,N_23794,N_23832);
and U24176 (N_24176,N_22693,N_23815);
xor U24177 (N_24177,N_23275,N_23008);
nand U24178 (N_24178,N_22796,N_22775);
and U24179 (N_24179,N_23381,N_23742);
nor U24180 (N_24180,N_22966,N_23934);
nand U24181 (N_24181,N_23121,N_23570);
nor U24182 (N_24182,N_23705,N_23792);
xnor U24183 (N_24183,N_22628,N_23405);
nand U24184 (N_24184,N_22845,N_23568);
and U24185 (N_24185,N_22639,N_23030);
nor U24186 (N_24186,N_22615,N_23075);
xor U24187 (N_24187,N_23833,N_22786);
nor U24188 (N_24188,N_23027,N_22550);
nor U24189 (N_24189,N_22687,N_22789);
nor U24190 (N_24190,N_23362,N_23494);
nand U24191 (N_24191,N_23596,N_23992);
and U24192 (N_24192,N_23437,N_23817);
nand U24193 (N_24193,N_22664,N_22527);
and U24194 (N_24194,N_23497,N_23552);
nand U24195 (N_24195,N_22741,N_23208);
nor U24196 (N_24196,N_22792,N_23203);
or U24197 (N_24197,N_23115,N_23409);
or U24198 (N_24198,N_23631,N_23323);
nand U24199 (N_24199,N_23435,N_23451);
or U24200 (N_24200,N_23042,N_22895);
nor U24201 (N_24201,N_23266,N_23543);
nand U24202 (N_24202,N_23031,N_22942);
or U24203 (N_24203,N_23137,N_22546);
nor U24204 (N_24204,N_22522,N_22862);
nand U24205 (N_24205,N_23964,N_22948);
xor U24206 (N_24206,N_22558,N_22706);
or U24207 (N_24207,N_22717,N_23124);
xor U24208 (N_24208,N_23186,N_23626);
nor U24209 (N_24209,N_22813,N_23071);
nand U24210 (N_24210,N_22869,N_22714);
nand U24211 (N_24211,N_22704,N_23411);
and U24212 (N_24212,N_23268,N_23661);
nor U24213 (N_24213,N_23938,N_23412);
nor U24214 (N_24214,N_22850,N_23139);
and U24215 (N_24215,N_23283,N_23600);
nor U24216 (N_24216,N_23263,N_23113);
or U24217 (N_24217,N_23188,N_23738);
and U24218 (N_24218,N_23955,N_22910);
or U24219 (N_24219,N_23057,N_23072);
and U24220 (N_24220,N_22509,N_22526);
nor U24221 (N_24221,N_23608,N_23109);
or U24222 (N_24222,N_23754,N_23063);
xnor U24223 (N_24223,N_22832,N_23853);
or U24224 (N_24224,N_22970,N_23478);
xnor U24225 (N_24225,N_23051,N_22611);
nor U24226 (N_24226,N_22957,N_22890);
xnor U24227 (N_24227,N_22569,N_22982);
nor U24228 (N_24228,N_23345,N_23201);
nand U24229 (N_24229,N_23911,N_23735);
nand U24230 (N_24230,N_22887,N_23892);
nand U24231 (N_24231,N_23882,N_23044);
and U24232 (N_24232,N_23249,N_22885);
nand U24233 (N_24233,N_22893,N_22570);
nor U24234 (N_24234,N_22990,N_22807);
xor U24235 (N_24235,N_22954,N_22666);
nor U24236 (N_24236,N_22659,N_23010);
or U24237 (N_24237,N_22863,N_22750);
nor U24238 (N_24238,N_23610,N_22809);
xor U24239 (N_24239,N_23054,N_22719);
and U24240 (N_24240,N_23194,N_23490);
nand U24241 (N_24241,N_23772,N_23001);
xnor U24242 (N_24242,N_23480,N_23745);
nand U24243 (N_24243,N_23684,N_22999);
xnor U24244 (N_24244,N_23090,N_23270);
nor U24245 (N_24245,N_23594,N_23489);
and U24246 (N_24246,N_22748,N_23787);
and U24247 (N_24247,N_23758,N_23069);
xor U24248 (N_24248,N_22656,N_22952);
and U24249 (N_24249,N_22564,N_23845);
or U24250 (N_24250,N_23560,N_23673);
nand U24251 (N_24251,N_23554,N_23575);
nor U24252 (N_24252,N_23096,N_23973);
or U24253 (N_24253,N_23248,N_23349);
or U24254 (N_24254,N_23388,N_23039);
nor U24255 (N_24255,N_23721,N_22762);
nand U24256 (N_24256,N_23727,N_22649);
nand U24257 (N_24257,N_22767,N_23747);
and U24258 (N_24258,N_23045,N_23146);
or U24259 (N_24259,N_22883,N_22926);
nor U24260 (N_24260,N_23770,N_22661);
or U24261 (N_24261,N_23272,N_23930);
or U24262 (N_24262,N_22545,N_23168);
and U24263 (N_24263,N_22930,N_23143);
or U24264 (N_24264,N_22914,N_23374);
nand U24265 (N_24265,N_23013,N_23583);
nand U24266 (N_24266,N_22631,N_23421);
xnor U24267 (N_24267,N_22502,N_22595);
and U24268 (N_24268,N_22612,N_23046);
xnor U24269 (N_24269,N_22822,N_22606);
or U24270 (N_24270,N_23524,N_22870);
or U24271 (N_24271,N_23185,N_23351);
xnor U24272 (N_24272,N_22975,N_23813);
xor U24273 (N_24273,N_22940,N_22776);
nor U24274 (N_24274,N_23983,N_23174);
nand U24275 (N_24275,N_22857,N_23935);
and U24276 (N_24276,N_23432,N_22830);
xnor U24277 (N_24277,N_23757,N_22933);
or U24278 (N_24278,N_23774,N_22927);
xnor U24279 (N_24279,N_23513,N_23578);
or U24280 (N_24280,N_23875,N_22510);
nor U24281 (N_24281,N_22995,N_23907);
and U24282 (N_24282,N_23257,N_22524);
and U24283 (N_24283,N_22616,N_23181);
nor U24284 (N_24284,N_23067,N_23719);
or U24285 (N_24285,N_23872,N_23528);
and U24286 (N_24286,N_23343,N_22749);
and U24287 (N_24287,N_23547,N_23686);
xor U24288 (N_24288,N_23433,N_23170);
nand U24289 (N_24289,N_23091,N_23785);
or U24290 (N_24290,N_22686,N_23236);
xor U24291 (N_24291,N_23215,N_23843);
and U24292 (N_24292,N_23790,N_22903);
xor U24293 (N_24293,N_22977,N_23736);
nor U24294 (N_24294,N_22774,N_22777);
and U24295 (N_24295,N_23632,N_23468);
xnor U24296 (N_24296,N_22634,N_22877);
xnor U24297 (N_24297,N_23050,N_23680);
or U24298 (N_24298,N_22673,N_22897);
nand U24299 (N_24299,N_23017,N_23918);
nand U24300 (N_24300,N_23308,N_23863);
nor U24301 (N_24301,N_23163,N_23173);
nand U24302 (N_24302,N_23313,N_22800);
nand U24303 (N_24303,N_23590,N_23280);
xor U24304 (N_24304,N_22922,N_22553);
nand U24305 (N_24305,N_22860,N_23445);
nand U24306 (N_24306,N_23693,N_22519);
xnor U24307 (N_24307,N_23332,N_22632);
and U24308 (N_24308,N_23237,N_22795);
xnor U24309 (N_24309,N_23645,N_23999);
xnor U24310 (N_24310,N_23799,N_23423);
or U24311 (N_24311,N_23162,N_22962);
and U24312 (N_24312,N_23984,N_23672);
or U24313 (N_24313,N_22884,N_22784);
nand U24314 (N_24314,N_23134,N_23341);
nand U24315 (N_24315,N_23430,N_22918);
xor U24316 (N_24316,N_23654,N_22878);
nor U24317 (N_24317,N_23878,N_22973);
or U24318 (N_24318,N_23699,N_23950);
and U24319 (N_24319,N_22572,N_23440);
and U24320 (N_24320,N_23114,N_23897);
or U24321 (N_24321,N_22880,N_22978);
or U24322 (N_24322,N_23363,N_23040);
nor U24323 (N_24323,N_22710,N_22773);
xnor U24324 (N_24324,N_23912,N_23354);
nor U24325 (N_24325,N_22517,N_23970);
or U24326 (N_24326,N_23676,N_22769);
nand U24327 (N_24327,N_22650,N_23571);
xor U24328 (N_24328,N_23260,N_23997);
nand U24329 (N_24329,N_23982,N_22520);
xor U24330 (N_24330,N_23517,N_22653);
or U24331 (N_24331,N_23668,N_23398);
or U24332 (N_24332,N_23888,N_23002);
nand U24333 (N_24333,N_23136,N_23976);
or U24334 (N_24334,N_23009,N_23016);
or U24335 (N_24335,N_22713,N_23368);
or U24336 (N_24336,N_23160,N_22797);
nand U24337 (N_24337,N_23344,N_23102);
xor U24338 (N_24338,N_23255,N_23965);
or U24339 (N_24339,N_23924,N_23961);
xor U24340 (N_24340,N_23933,N_22938);
nand U24341 (N_24341,N_23110,N_23410);
or U24342 (N_24342,N_23979,N_22866);
or U24343 (N_24343,N_22856,N_22818);
xnor U24344 (N_24344,N_22707,N_23293);
or U24345 (N_24345,N_22705,N_23759);
or U24346 (N_24346,N_23023,N_23889);
and U24347 (N_24347,N_22837,N_22655);
nand U24348 (N_24348,N_23211,N_23442);
or U24349 (N_24349,N_23097,N_23151);
and U24350 (N_24350,N_22768,N_22709);
and U24351 (N_24351,N_22617,N_23240);
xnor U24352 (N_24352,N_22911,N_23496);
nand U24353 (N_24353,N_23372,N_22872);
nor U24354 (N_24354,N_23666,N_23191);
nand U24355 (N_24355,N_23416,N_23369);
nand U24356 (N_24356,N_23314,N_22696);
nand U24357 (N_24357,N_23172,N_23222);
nand U24358 (N_24358,N_23804,N_22782);
nand U24359 (N_24359,N_23688,N_23881);
xnor U24360 (N_24360,N_23643,N_23111);
nor U24361 (N_24361,N_22587,N_23085);
xor U24362 (N_24362,N_23775,N_23166);
or U24363 (N_24363,N_23036,N_23209);
xnor U24364 (N_24364,N_22746,N_22876);
xnor U24365 (N_24365,N_23198,N_22602);
xor U24366 (N_24366,N_23947,N_23331);
nor U24367 (N_24367,N_23144,N_23418);
xnor U24368 (N_24368,N_23885,N_22858);
or U24369 (N_24369,N_22759,N_22674);
or U24370 (N_24370,N_23764,N_22751);
xnor U24371 (N_24371,N_23523,N_22591);
nand U24372 (N_24372,N_23056,N_22682);
nor U24373 (N_24373,N_22589,N_22581);
or U24374 (N_24374,N_22891,N_22755);
nand U24375 (N_24375,N_23515,N_23797);
xnor U24376 (N_24376,N_22514,N_22540);
and U24377 (N_24377,N_22808,N_22997);
xnor U24378 (N_24378,N_23183,N_23251);
nand U24379 (N_24379,N_23708,N_22625);
nor U24380 (N_24380,N_23455,N_22815);
xor U24381 (N_24381,N_23020,N_23053);
xor U24382 (N_24382,N_23492,N_23617);
nand U24383 (N_24383,N_22793,N_22697);
xnor U24384 (N_24384,N_23462,N_23549);
nand U24385 (N_24385,N_23715,N_23358);
nand U24386 (N_24386,N_22919,N_23465);
or U24387 (N_24387,N_23692,N_22584);
or U24388 (N_24388,N_23190,N_23205);
nand U24389 (N_24389,N_23028,N_23390);
or U24390 (N_24390,N_23621,N_23932);
xor U24391 (N_24391,N_23361,N_23698);
xnor U24392 (N_24392,N_22685,N_23220);
and U24393 (N_24393,N_22998,N_23342);
or U24394 (N_24394,N_23501,N_23367);
nand U24395 (N_24395,N_23104,N_23138);
nor U24396 (N_24396,N_23422,N_23917);
or U24397 (N_24397,N_23953,N_22771);
xor U24398 (N_24398,N_22934,N_23204);
and U24399 (N_24399,N_23428,N_23855);
and U24400 (N_24400,N_22571,N_22993);
nor U24401 (N_24401,N_23402,N_22660);
nand U24402 (N_24402,N_23857,N_23835);
and U24403 (N_24403,N_22531,N_23488);
and U24404 (N_24404,N_23140,N_23511);
nor U24405 (N_24405,N_23861,N_22996);
and U24406 (N_24406,N_23223,N_22523);
and U24407 (N_24407,N_23870,N_22908);
and U24408 (N_24408,N_22652,N_22554);
and U24409 (N_24409,N_22726,N_23954);
nand U24410 (N_24410,N_22551,N_23537);
and U24411 (N_24411,N_22972,N_23401);
nor U24412 (N_24412,N_23238,N_23177);
xnor U24413 (N_24413,N_23980,N_23740);
nor U24414 (N_24414,N_22575,N_22941);
xnor U24415 (N_24415,N_23383,N_22831);
and U24416 (N_24416,N_23265,N_23502);
or U24417 (N_24417,N_23629,N_22603);
and U24418 (N_24418,N_23371,N_23250);
or U24419 (N_24419,N_22753,N_22592);
nand U24420 (N_24420,N_23466,N_23842);
or U24421 (N_24421,N_22936,N_22692);
xnor U24422 (N_24422,N_23328,N_22740);
and U24423 (N_24423,N_23395,N_23744);
nor U24424 (N_24424,N_23099,N_23674);
or U24425 (N_24425,N_23819,N_23024);
xor U24426 (N_24426,N_22727,N_22989);
or U24427 (N_24427,N_23450,N_23586);
nand U24428 (N_24428,N_23200,N_22533);
nand U24429 (N_24429,N_23856,N_23656);
or U24430 (N_24430,N_22542,N_22787);
or U24431 (N_24431,N_23728,N_23365);
xnor U24432 (N_24432,N_23309,N_23495);
nand U24433 (N_24433,N_22641,N_23902);
or U24434 (N_24434,N_23956,N_23391);
xnor U24435 (N_24435,N_23891,N_23622);
and U24436 (N_24436,N_23052,N_23660);
and U24437 (N_24437,N_22901,N_23653);
nand U24438 (N_24438,N_23472,N_22881);
or U24439 (N_24439,N_23092,N_22736);
xor U24440 (N_24440,N_22783,N_23380);
or U24441 (N_24441,N_23184,N_23169);
xnor U24442 (N_24442,N_23798,N_23831);
and U24443 (N_24443,N_22950,N_22864);
nor U24444 (N_24444,N_23559,N_23944);
nor U24445 (N_24445,N_23064,N_23325);
xnor U24446 (N_24446,N_22583,N_23444);
or U24447 (N_24447,N_23795,N_23714);
and U24448 (N_24448,N_23034,N_23994);
and U24449 (N_24449,N_23858,N_23087);
nand U24450 (N_24450,N_23193,N_23269);
nand U24451 (N_24451,N_23256,N_23360);
nor U24452 (N_24452,N_22516,N_22645);
xnor U24453 (N_24453,N_23105,N_23604);
or U24454 (N_24454,N_22689,N_23526);
nand U24455 (N_24455,N_23948,N_23021);
or U24456 (N_24456,N_23366,N_23598);
nand U24457 (N_24457,N_23334,N_22548);
xor U24458 (N_24458,N_23306,N_22582);
nand U24459 (N_24459,N_22764,N_23895);
nand U24460 (N_24460,N_23975,N_23589);
and U24461 (N_24461,N_23284,N_22742);
nor U24462 (N_24462,N_23840,N_23093);
or U24463 (N_24463,N_23846,N_22623);
nand U24464 (N_24464,N_22501,N_22816);
nand U24465 (N_24465,N_23952,N_23393);
nor U24466 (N_24466,N_23335,N_23945);
nor U24467 (N_24467,N_22557,N_23487);
xnor U24468 (N_24468,N_23287,N_22723);
or U24469 (N_24469,N_22928,N_22504);
or U24470 (N_24470,N_22943,N_23553);
nor U24471 (N_24471,N_22658,N_23126);
or U24472 (N_24472,N_23004,N_23990);
xnor U24473 (N_24473,N_22974,N_23292);
or U24474 (N_24474,N_23869,N_23871);
nand U24475 (N_24475,N_23630,N_23602);
and U24476 (N_24476,N_23521,N_22547);
and U24477 (N_24477,N_23261,N_23665);
or U24478 (N_24478,N_22534,N_23725);
or U24479 (N_24479,N_23285,N_23913);
or U24480 (N_24480,N_23147,N_23330);
nor U24481 (N_24481,N_23338,N_23294);
and U24482 (N_24482,N_23978,N_22946);
or U24483 (N_24483,N_23207,N_23929);
or U24484 (N_24484,N_23469,N_22859);
or U24485 (N_24485,N_23425,N_22619);
xnor U24486 (N_24486,N_22835,N_23609);
and U24487 (N_24487,N_23049,N_22819);
and U24488 (N_24488,N_23300,N_23060);
xnor U24489 (N_24489,N_23704,N_23786);
or U24490 (N_24490,N_23217,N_23206);
and U24491 (N_24491,N_23867,N_23296);
nand U24492 (N_24492,N_23716,N_23985);
or U24493 (N_24493,N_22899,N_23158);
and U24494 (N_24494,N_22817,N_23847);
nand U24495 (N_24495,N_22820,N_22620);
nor U24496 (N_24496,N_23149,N_23419);
xor U24497 (N_24497,N_22677,N_23695);
and U24498 (N_24498,N_23801,N_23564);
nor U24499 (N_24499,N_22657,N_23153);
nand U24500 (N_24500,N_23221,N_23905);
nor U24501 (N_24501,N_23556,N_22955);
and U24502 (N_24502,N_23977,N_23746);
nand U24503 (N_24503,N_22525,N_23936);
xor U24504 (N_24504,N_23491,N_22810);
nand U24505 (N_24505,N_23723,N_23830);
nor U24506 (N_24506,N_23696,N_23350);
xor U24507 (N_24507,N_23864,N_23482);
xor U24508 (N_24508,N_23706,N_22601);
nand U24509 (N_24509,N_23951,N_23967);
and U24510 (N_24510,N_23011,N_23005);
nor U24511 (N_24511,N_22566,N_23906);
and U24512 (N_24512,N_22916,N_23677);
xor U24513 (N_24513,N_23312,N_23403);
and U24514 (N_24514,N_23329,N_23803);
xnor U24515 (N_24515,N_22642,N_22596);
and U24516 (N_24516,N_23120,N_23601);
and U24517 (N_24517,N_23605,N_23664);
and U24518 (N_24518,N_23572,N_22680);
xor U24519 (N_24519,N_23291,N_22732);
or U24520 (N_24520,N_23068,N_23106);
or U24521 (N_24521,N_23454,N_23816);
nor U24522 (N_24522,N_23224,N_22637);
nor U24523 (N_24523,N_22544,N_23587);
and U24524 (N_24524,N_23493,N_22665);
or U24525 (N_24525,N_23192,N_23836);
xor U24526 (N_24526,N_22737,N_22760);
xor U24527 (N_24527,N_22896,N_23033);
xor U24528 (N_24528,N_23336,N_23752);
nand U24529 (N_24529,N_22839,N_23239);
xnor U24530 (N_24530,N_23658,N_22865);
xor U24531 (N_24531,N_23232,N_22691);
and U24532 (N_24532,N_22960,N_22563);
nor U24533 (N_24533,N_22900,N_23247);
or U24534 (N_24534,N_23429,N_23456);
nor U24535 (N_24535,N_23655,N_23127);
nor U24536 (N_24536,N_23995,N_23822);
nor U24537 (N_24537,N_23315,N_23007);
nor U24538 (N_24538,N_23333,N_23218);
nor U24539 (N_24539,N_22718,N_23868);
and U24540 (N_24540,N_23130,N_23408);
or U24541 (N_24541,N_22781,N_22824);
or U24542 (N_24542,N_22552,N_23989);
nor U24543 (N_24543,N_22805,N_23648);
nand U24544 (N_24544,N_22846,N_23784);
nor U24545 (N_24545,N_23866,N_23900);
or U24546 (N_24546,N_23061,N_22695);
or U24547 (N_24547,N_23536,N_23473);
and U24548 (N_24548,N_23446,N_23663);
nand U24549 (N_24549,N_23231,N_23463);
xnor U24550 (N_24550,N_23731,N_23377);
xnor U24551 (N_24551,N_23316,N_22935);
xor U24552 (N_24552,N_23370,N_23593);
nor U24553 (N_24553,N_23389,N_23733);
or U24554 (N_24554,N_23899,N_23854);
nand U24555 (N_24555,N_23299,N_23993);
nor U24556 (N_24556,N_23712,N_23095);
and U24557 (N_24557,N_23922,N_23180);
nor U24558 (N_24558,N_22814,N_22849);
and U24559 (N_24559,N_23647,N_23152);
and U24560 (N_24560,N_23957,N_23129);
or U24561 (N_24561,N_22874,N_22882);
or U24562 (N_24562,N_23834,N_23006);
xnor U24563 (N_24563,N_22574,N_22647);
or U24564 (N_24564,N_23996,N_22875);
and U24565 (N_24565,N_23903,N_23397);
and U24566 (N_24566,N_23148,N_23150);
nand U24567 (N_24567,N_23142,N_23667);
nand U24568 (N_24568,N_23756,N_22967);
xor U24569 (N_24569,N_23844,N_22904);
nor U24570 (N_24570,N_22712,N_23470);
and U24571 (N_24571,N_23364,N_23059);
nand U24572 (N_24572,N_23625,N_23310);
nand U24573 (N_24573,N_22568,N_22909);
or U24574 (N_24574,N_23584,N_22559);
or U24575 (N_24575,N_23852,N_22905);
or U24576 (N_24576,N_23295,N_23821);
nor U24577 (N_24577,N_23481,N_23937);
and U24578 (N_24578,N_23616,N_23116);
nor U24579 (N_24579,N_23657,N_23014);
nand U24580 (N_24580,N_23958,N_22679);
or U24581 (N_24581,N_22648,N_23646);
nand U24582 (N_24582,N_23375,N_22829);
nand U24583 (N_24583,N_23928,N_22976);
or U24584 (N_24584,N_22979,N_23219);
nand U24585 (N_24585,N_23119,N_23510);
xnor U24586 (N_24586,N_23862,N_23808);
nor U24587 (N_24587,N_22549,N_23319);
nand U24588 (N_24588,N_22821,N_23720);
xnor U24589 (N_24589,N_23279,N_22694);
and U24590 (N_24590,N_22701,N_22898);
nor U24591 (N_24591,N_23199,N_23768);
xor U24592 (N_24592,N_22654,N_22987);
and U24593 (N_24593,N_23460,N_23659);
or U24594 (N_24594,N_22530,N_22964);
nand U24595 (N_24595,N_23814,N_22670);
nand U24596 (N_24596,N_22511,N_23189);
and U24597 (N_24597,N_23789,N_23579);
nand U24598 (N_24598,N_22672,N_23802);
or U24599 (N_24599,N_22579,N_23599);
nand U24600 (N_24600,N_22770,N_22794);
nand U24601 (N_24601,N_23522,N_23561);
nor U24602 (N_24602,N_23988,N_23615);
or U24603 (N_24603,N_22733,N_23519);
nor U24604 (N_24604,N_23117,N_22627);
and U24605 (N_24605,N_23431,N_22840);
nor U24606 (N_24606,N_23687,N_23476);
nor U24607 (N_24607,N_23202,N_23253);
xnor U24608 (N_24608,N_22500,N_22636);
or U24609 (N_24609,N_23443,N_23384);
nor U24610 (N_24610,N_22683,N_22640);
nand U24611 (N_24611,N_23165,N_23083);
or U24612 (N_24612,N_22834,N_23779);
nand U24613 (N_24613,N_23434,N_22867);
and U24614 (N_24614,N_23718,N_23919);
nand U24615 (N_24615,N_22537,N_23258);
nor U24616 (N_24616,N_23297,N_22968);
xnor U24617 (N_24617,N_22944,N_23378);
nand U24618 (N_24618,N_22913,N_22745);
or U24619 (N_24619,N_23748,N_23796);
and U24620 (N_24620,N_22799,N_23025);
and U24621 (N_24621,N_23485,N_23791);
or U24622 (N_24622,N_23484,N_23077);
xnor U24623 (N_24623,N_23662,N_22585);
nor U24624 (N_24624,N_22724,N_23241);
or U24625 (N_24625,N_23065,N_23755);
nor U24626 (N_24626,N_23318,N_23504);
nand U24627 (N_24627,N_23508,N_23074);
xnor U24628 (N_24628,N_23576,N_23399);
or U24629 (N_24629,N_23327,N_23873);
or U24630 (N_24630,N_23709,N_23347);
and U24631 (N_24631,N_23966,N_23865);
or U24632 (N_24632,N_23880,N_22565);
and U24633 (N_24633,N_22823,N_23569);
or U24634 (N_24634,N_22646,N_23337);
nor U24635 (N_24635,N_22804,N_23771);
and U24636 (N_24636,N_23321,N_23782);
or U24637 (N_24637,N_23156,N_22738);
nand U24638 (N_24638,N_23691,N_22739);
nand U24639 (N_24639,N_23753,N_23516);
and U24640 (N_24640,N_23824,N_22715);
nand U24641 (N_24641,N_23694,N_23923);
or U24642 (N_24642,N_23839,N_22671);
xor U24643 (N_24643,N_23267,N_23290);
or U24644 (N_24644,N_23893,N_23942);
or U24645 (N_24645,N_23066,N_23227);
nor U24646 (N_24646,N_22700,N_23289);
xor U24647 (N_24647,N_22543,N_22765);
and U24648 (N_24648,N_23986,N_22561);
or U24649 (N_24649,N_22833,N_23213);
nand U24650 (N_24650,N_23638,N_23582);
nand U24651 (N_24651,N_23486,N_23717);
and U24652 (N_24652,N_23135,N_22507);
nor U24653 (N_24653,N_23094,N_22593);
and U24654 (N_24654,N_22906,N_22873);
and U24655 (N_24655,N_22945,N_23242);
xor U24656 (N_24656,N_23041,N_23355);
xor U24657 (N_24657,N_22790,N_23828);
nand U24658 (N_24658,N_22630,N_23216);
xnor U24659 (N_24659,N_22678,N_23739);
xor U24660 (N_24660,N_23960,N_22923);
and U24661 (N_24661,N_23122,N_22518);
xor U24662 (N_24662,N_23503,N_23534);
xor U24663 (N_24663,N_23825,N_23807);
nor U24664 (N_24664,N_22730,N_23182);
nor U24665 (N_24665,N_22668,N_23921);
nand U24666 (N_24666,N_23540,N_22802);
or U24667 (N_24667,N_22785,N_22788);
nand U24668 (N_24668,N_23767,N_23910);
nor U24669 (N_24669,N_22854,N_22828);
or U24670 (N_24670,N_22576,N_23941);
and U24671 (N_24671,N_22981,N_23264);
or U24672 (N_24672,N_23894,N_23235);
xnor U24673 (N_24673,N_23580,N_22743);
nand U24674 (N_24674,N_22826,N_22915);
or U24675 (N_24675,N_22939,N_23225);
xnor U24676 (N_24676,N_23793,N_23471);
and U24677 (N_24677,N_23700,N_22980);
or U24678 (N_24678,N_22716,N_23781);
and U24679 (N_24679,N_23898,N_23800);
and U24680 (N_24680,N_23301,N_23959);
xor U24681 (N_24681,N_23558,N_23765);
nand U24682 (N_24682,N_22744,N_22614);
nor U24683 (N_24683,N_23233,N_23392);
nand U24684 (N_24684,N_23154,N_23464);
xnor U24685 (N_24685,N_23447,N_23585);
or U24686 (N_24686,N_23546,N_23082);
nand U24687 (N_24687,N_23076,N_23876);
nor U24688 (N_24688,N_23458,N_23080);
nor U24689 (N_24689,N_23128,N_23652);
or U24690 (N_24690,N_22663,N_22780);
nand U24691 (N_24691,N_23860,N_23544);
nor U24692 (N_24692,N_22503,N_22994);
xnor U24693 (N_24693,N_23931,N_23108);
nand U24694 (N_24694,N_22532,N_23879);
xor U24695 (N_24695,N_23386,N_22567);
or U24696 (N_24696,N_22841,N_23157);
nor U24697 (N_24697,N_23187,N_22868);
or U24698 (N_24698,N_23614,N_23603);
or U24699 (N_24699,N_23427,N_22852);
xor U24700 (N_24700,N_22513,N_22580);
nand U24701 (N_24701,N_23175,N_23939);
nand U24702 (N_24702,N_22528,N_23530);
nor U24703 (N_24703,N_23228,N_23234);
xnor U24704 (N_24704,N_23340,N_23118);
nand U24705 (N_24705,N_23619,N_23904);
xor U24706 (N_24706,N_23196,N_22836);
and U24707 (N_24707,N_23987,N_23079);
xor U24708 (N_24708,N_23532,N_23806);
and U24709 (N_24709,N_23531,N_23178);
or U24710 (N_24710,N_23015,N_22929);
or U24711 (N_24711,N_23689,N_23620);
nand U24712 (N_24712,N_23230,N_23974);
nor U24713 (N_24713,N_23577,N_23788);
and U24714 (N_24714,N_23164,N_22848);
nor U24715 (N_24715,N_22912,N_22535);
nand U24716 (N_24716,N_23352,N_23195);
or U24717 (N_24717,N_22988,N_23467);
nor U24718 (N_24718,N_23132,N_23890);
or U24719 (N_24719,N_22626,N_23509);
nor U24720 (N_24720,N_23741,N_23812);
nor U24721 (N_24721,N_23574,N_23743);
nand U24722 (N_24722,N_23058,N_22675);
and U24723 (N_24723,N_23627,N_23520);
nor U24724 (N_24724,N_23682,N_23441);
nor U24725 (N_24725,N_23874,N_23047);
and U24726 (N_24726,N_22508,N_22844);
xnor U24727 (N_24727,N_23112,N_22536);
and U24728 (N_24728,N_22924,N_22644);
and U24729 (N_24729,N_23563,N_23101);
and U24730 (N_24730,N_22801,N_22731);
xor U24731 (N_24731,N_22669,N_23607);
xor U24732 (N_24732,N_23000,N_23595);
or U24733 (N_24733,N_23581,N_23474);
or U24734 (N_24734,N_23449,N_22838);
or U24735 (N_24735,N_23737,N_23506);
nand U24736 (N_24736,N_22512,N_22766);
or U24737 (N_24737,N_23003,N_23613);
and U24738 (N_24738,N_23514,N_23055);
or U24739 (N_24739,N_22624,N_23089);
and U24740 (N_24740,N_23527,N_22951);
and U24741 (N_24741,N_23498,N_23968);
and U24742 (N_24742,N_23346,N_23724);
xnor U24743 (N_24743,N_22992,N_22562);
and U24744 (N_24744,N_22635,N_23376);
or U24745 (N_24745,N_23459,N_23533);
and U24746 (N_24746,N_23841,N_23823);
and U24747 (N_24747,N_23500,N_23760);
and U24748 (N_24748,N_23776,N_22917);
nand U24749 (N_24749,N_23317,N_23086);
and U24750 (N_24750,N_23607,N_22714);
xor U24751 (N_24751,N_23015,N_22559);
or U24752 (N_24752,N_23449,N_22570);
nand U24753 (N_24753,N_23207,N_22524);
xor U24754 (N_24754,N_23552,N_23869);
or U24755 (N_24755,N_23404,N_22681);
xor U24756 (N_24756,N_22919,N_23256);
or U24757 (N_24757,N_23909,N_22662);
nor U24758 (N_24758,N_23002,N_23254);
nand U24759 (N_24759,N_23894,N_22540);
and U24760 (N_24760,N_23282,N_23254);
xor U24761 (N_24761,N_22630,N_23073);
nand U24762 (N_24762,N_22749,N_22971);
or U24763 (N_24763,N_22871,N_23243);
nor U24764 (N_24764,N_23773,N_22598);
nor U24765 (N_24765,N_22971,N_23425);
or U24766 (N_24766,N_23261,N_23440);
and U24767 (N_24767,N_23404,N_23050);
nor U24768 (N_24768,N_23336,N_22633);
and U24769 (N_24769,N_23379,N_23686);
xor U24770 (N_24770,N_23027,N_23173);
and U24771 (N_24771,N_23000,N_23529);
xnor U24772 (N_24772,N_23526,N_23093);
or U24773 (N_24773,N_23494,N_23346);
or U24774 (N_24774,N_23430,N_22940);
nand U24775 (N_24775,N_22667,N_23170);
xor U24776 (N_24776,N_22598,N_23483);
or U24777 (N_24777,N_23102,N_23426);
or U24778 (N_24778,N_23342,N_22761);
xnor U24779 (N_24779,N_22951,N_23940);
nor U24780 (N_24780,N_23724,N_23813);
nor U24781 (N_24781,N_23944,N_23448);
xnor U24782 (N_24782,N_23486,N_23375);
or U24783 (N_24783,N_22583,N_23829);
and U24784 (N_24784,N_23899,N_23508);
and U24785 (N_24785,N_23976,N_23578);
and U24786 (N_24786,N_23876,N_23282);
nor U24787 (N_24787,N_23345,N_22698);
nor U24788 (N_24788,N_23338,N_23486);
or U24789 (N_24789,N_23554,N_22938);
nor U24790 (N_24790,N_23959,N_22949);
nor U24791 (N_24791,N_23606,N_22719);
and U24792 (N_24792,N_23843,N_23381);
nand U24793 (N_24793,N_23422,N_23846);
and U24794 (N_24794,N_23594,N_23272);
xnor U24795 (N_24795,N_22788,N_22933);
nand U24796 (N_24796,N_22839,N_22736);
nor U24797 (N_24797,N_22943,N_23170);
and U24798 (N_24798,N_23317,N_23379);
and U24799 (N_24799,N_23812,N_23452);
or U24800 (N_24800,N_22966,N_23849);
nor U24801 (N_24801,N_22889,N_23110);
and U24802 (N_24802,N_22583,N_22550);
and U24803 (N_24803,N_23316,N_23360);
or U24804 (N_24804,N_22590,N_22784);
nand U24805 (N_24805,N_22867,N_23162);
nand U24806 (N_24806,N_23547,N_22867);
and U24807 (N_24807,N_23891,N_23141);
or U24808 (N_24808,N_23204,N_23398);
or U24809 (N_24809,N_23050,N_23777);
and U24810 (N_24810,N_23079,N_22638);
nand U24811 (N_24811,N_23976,N_22752);
or U24812 (N_24812,N_23543,N_23313);
xor U24813 (N_24813,N_23361,N_22952);
nor U24814 (N_24814,N_23320,N_23777);
nand U24815 (N_24815,N_23925,N_22721);
nand U24816 (N_24816,N_23477,N_22678);
nand U24817 (N_24817,N_23973,N_23782);
or U24818 (N_24818,N_22662,N_22903);
and U24819 (N_24819,N_23229,N_23989);
and U24820 (N_24820,N_23660,N_22515);
nor U24821 (N_24821,N_23886,N_23900);
nor U24822 (N_24822,N_22825,N_23827);
xor U24823 (N_24823,N_23277,N_22750);
or U24824 (N_24824,N_22773,N_23920);
or U24825 (N_24825,N_23124,N_22533);
xor U24826 (N_24826,N_23109,N_22677);
xnor U24827 (N_24827,N_22578,N_23174);
xnor U24828 (N_24828,N_23333,N_23608);
nand U24829 (N_24829,N_23235,N_23314);
or U24830 (N_24830,N_23464,N_23407);
xnor U24831 (N_24831,N_23632,N_23617);
or U24832 (N_24832,N_23285,N_22971);
nand U24833 (N_24833,N_23880,N_22636);
nor U24834 (N_24834,N_23821,N_23328);
xnor U24835 (N_24835,N_22781,N_22991);
or U24836 (N_24836,N_22680,N_23822);
nand U24837 (N_24837,N_22541,N_22913);
nor U24838 (N_24838,N_22559,N_23715);
or U24839 (N_24839,N_22611,N_22630);
and U24840 (N_24840,N_23550,N_23044);
or U24841 (N_24841,N_22631,N_23539);
and U24842 (N_24842,N_22618,N_22633);
or U24843 (N_24843,N_22789,N_23567);
nand U24844 (N_24844,N_23846,N_22943);
nand U24845 (N_24845,N_23158,N_23100);
or U24846 (N_24846,N_22509,N_23621);
and U24847 (N_24847,N_22713,N_23674);
nand U24848 (N_24848,N_23162,N_23213);
and U24849 (N_24849,N_23727,N_23141);
nand U24850 (N_24850,N_22900,N_23046);
nor U24851 (N_24851,N_23868,N_23070);
nand U24852 (N_24852,N_23227,N_23398);
and U24853 (N_24853,N_22747,N_23667);
nand U24854 (N_24854,N_23509,N_23479);
nand U24855 (N_24855,N_23662,N_22746);
nand U24856 (N_24856,N_22925,N_22939);
nand U24857 (N_24857,N_22706,N_23544);
xor U24858 (N_24858,N_23592,N_22682);
and U24859 (N_24859,N_22846,N_22987);
nand U24860 (N_24860,N_23064,N_23792);
xnor U24861 (N_24861,N_23094,N_22865);
nand U24862 (N_24862,N_23279,N_23444);
xnor U24863 (N_24863,N_23153,N_23231);
and U24864 (N_24864,N_22810,N_23487);
nand U24865 (N_24865,N_23021,N_23081);
or U24866 (N_24866,N_22708,N_23050);
nand U24867 (N_24867,N_23659,N_23840);
or U24868 (N_24868,N_22892,N_23127);
xor U24869 (N_24869,N_23267,N_23252);
nor U24870 (N_24870,N_23728,N_23028);
or U24871 (N_24871,N_23254,N_23054);
or U24872 (N_24872,N_22768,N_22990);
nor U24873 (N_24873,N_23804,N_23970);
xor U24874 (N_24874,N_23558,N_23630);
xor U24875 (N_24875,N_22986,N_23071);
and U24876 (N_24876,N_22509,N_23880);
xor U24877 (N_24877,N_23853,N_23836);
and U24878 (N_24878,N_23294,N_22893);
nand U24879 (N_24879,N_23151,N_23138);
nor U24880 (N_24880,N_23062,N_23328);
xor U24881 (N_24881,N_22647,N_23481);
and U24882 (N_24882,N_22644,N_23304);
and U24883 (N_24883,N_23885,N_23556);
nand U24884 (N_24884,N_23583,N_23622);
nor U24885 (N_24885,N_22907,N_23894);
xor U24886 (N_24886,N_23667,N_22506);
or U24887 (N_24887,N_23168,N_23351);
nand U24888 (N_24888,N_23359,N_23721);
nor U24889 (N_24889,N_23803,N_23683);
nor U24890 (N_24890,N_23471,N_22628);
nand U24891 (N_24891,N_23518,N_22841);
xor U24892 (N_24892,N_22979,N_23994);
or U24893 (N_24893,N_23002,N_23721);
nand U24894 (N_24894,N_23275,N_22663);
xor U24895 (N_24895,N_22719,N_23632);
or U24896 (N_24896,N_23493,N_23363);
nand U24897 (N_24897,N_22671,N_23403);
or U24898 (N_24898,N_22885,N_23407);
nor U24899 (N_24899,N_23855,N_23176);
nor U24900 (N_24900,N_23168,N_23089);
or U24901 (N_24901,N_23412,N_23650);
or U24902 (N_24902,N_23048,N_23200);
xnor U24903 (N_24903,N_23238,N_22685);
nand U24904 (N_24904,N_23489,N_22630);
or U24905 (N_24905,N_22773,N_23890);
nand U24906 (N_24906,N_22955,N_22754);
xnor U24907 (N_24907,N_22822,N_22906);
xnor U24908 (N_24908,N_22693,N_23394);
xnor U24909 (N_24909,N_23155,N_22887);
nor U24910 (N_24910,N_23051,N_22875);
or U24911 (N_24911,N_22534,N_22689);
nor U24912 (N_24912,N_23100,N_23278);
and U24913 (N_24913,N_23826,N_22923);
and U24914 (N_24914,N_23135,N_23206);
and U24915 (N_24915,N_22634,N_23031);
xnor U24916 (N_24916,N_23947,N_23447);
nand U24917 (N_24917,N_22914,N_23338);
or U24918 (N_24918,N_23386,N_23797);
nor U24919 (N_24919,N_23500,N_23029);
xor U24920 (N_24920,N_22669,N_23671);
and U24921 (N_24921,N_23195,N_22845);
or U24922 (N_24922,N_22931,N_23247);
or U24923 (N_24923,N_23586,N_23889);
and U24924 (N_24924,N_23271,N_22637);
nor U24925 (N_24925,N_23253,N_23628);
and U24926 (N_24926,N_23784,N_22758);
nor U24927 (N_24927,N_22842,N_23006);
and U24928 (N_24928,N_23755,N_23672);
xor U24929 (N_24929,N_22862,N_23453);
and U24930 (N_24930,N_23006,N_22923);
and U24931 (N_24931,N_22741,N_23727);
or U24932 (N_24932,N_23117,N_23896);
nand U24933 (N_24933,N_23647,N_23163);
or U24934 (N_24934,N_22906,N_23351);
or U24935 (N_24935,N_22676,N_23958);
xnor U24936 (N_24936,N_23159,N_23463);
nand U24937 (N_24937,N_23545,N_23808);
or U24938 (N_24938,N_23054,N_23682);
and U24939 (N_24939,N_23069,N_23964);
nor U24940 (N_24940,N_23091,N_22632);
and U24941 (N_24941,N_22998,N_22736);
and U24942 (N_24942,N_23302,N_23384);
nor U24943 (N_24943,N_23729,N_22907);
nand U24944 (N_24944,N_22946,N_23784);
xor U24945 (N_24945,N_22680,N_23942);
or U24946 (N_24946,N_23503,N_22674);
nand U24947 (N_24947,N_22681,N_23276);
or U24948 (N_24948,N_23067,N_23328);
and U24949 (N_24949,N_23421,N_22917);
nor U24950 (N_24950,N_22646,N_23815);
or U24951 (N_24951,N_23175,N_23450);
nor U24952 (N_24952,N_23892,N_23686);
nor U24953 (N_24953,N_23901,N_22516);
and U24954 (N_24954,N_23528,N_23331);
xnor U24955 (N_24955,N_22647,N_22925);
or U24956 (N_24956,N_22856,N_22849);
and U24957 (N_24957,N_23599,N_23027);
or U24958 (N_24958,N_23117,N_23789);
or U24959 (N_24959,N_22595,N_22848);
nor U24960 (N_24960,N_23669,N_22578);
and U24961 (N_24961,N_23477,N_23880);
and U24962 (N_24962,N_22980,N_23537);
nor U24963 (N_24963,N_23851,N_22817);
and U24964 (N_24964,N_23878,N_22758);
xnor U24965 (N_24965,N_22590,N_22828);
nor U24966 (N_24966,N_23544,N_23285);
nand U24967 (N_24967,N_23704,N_23827);
nor U24968 (N_24968,N_22899,N_23322);
or U24969 (N_24969,N_23183,N_23749);
or U24970 (N_24970,N_23242,N_22694);
nor U24971 (N_24971,N_23260,N_22974);
nor U24972 (N_24972,N_23089,N_22866);
or U24973 (N_24973,N_23582,N_23067);
nor U24974 (N_24974,N_22674,N_23801);
and U24975 (N_24975,N_23530,N_23094);
and U24976 (N_24976,N_23561,N_23536);
nor U24977 (N_24977,N_23800,N_22570);
and U24978 (N_24978,N_23994,N_23691);
nor U24979 (N_24979,N_22636,N_23126);
nor U24980 (N_24980,N_23399,N_22943);
and U24981 (N_24981,N_23935,N_23426);
xor U24982 (N_24982,N_22771,N_23111);
or U24983 (N_24983,N_23780,N_22658);
nand U24984 (N_24984,N_23266,N_23097);
nor U24985 (N_24985,N_23914,N_23690);
and U24986 (N_24986,N_22949,N_23247);
xnor U24987 (N_24987,N_22855,N_22952);
xor U24988 (N_24988,N_23491,N_22615);
xnor U24989 (N_24989,N_23363,N_23187);
or U24990 (N_24990,N_23519,N_23486);
nor U24991 (N_24991,N_23490,N_23548);
xor U24992 (N_24992,N_22943,N_22647);
or U24993 (N_24993,N_23033,N_23749);
nand U24994 (N_24994,N_23032,N_23255);
xnor U24995 (N_24995,N_22900,N_23114);
and U24996 (N_24996,N_23735,N_23061);
nand U24997 (N_24997,N_22885,N_23776);
and U24998 (N_24998,N_22775,N_23913);
xnor U24999 (N_24999,N_22846,N_22959);
and U25000 (N_25000,N_23339,N_23078);
or U25001 (N_25001,N_23288,N_22694);
and U25002 (N_25002,N_23692,N_22976);
or U25003 (N_25003,N_22765,N_22681);
or U25004 (N_25004,N_22717,N_23519);
nand U25005 (N_25005,N_23052,N_23288);
nand U25006 (N_25006,N_23529,N_23361);
xor U25007 (N_25007,N_23620,N_23993);
xnor U25008 (N_25008,N_23079,N_23748);
nor U25009 (N_25009,N_22835,N_23193);
or U25010 (N_25010,N_23004,N_22590);
or U25011 (N_25011,N_22887,N_22574);
xnor U25012 (N_25012,N_23864,N_23439);
and U25013 (N_25013,N_23994,N_22907);
xor U25014 (N_25014,N_23104,N_22595);
xor U25015 (N_25015,N_23232,N_22940);
xnor U25016 (N_25016,N_22680,N_23795);
and U25017 (N_25017,N_23469,N_23161);
xor U25018 (N_25018,N_22646,N_23655);
nand U25019 (N_25019,N_23720,N_22789);
nand U25020 (N_25020,N_22542,N_23434);
xnor U25021 (N_25021,N_23229,N_23959);
xor U25022 (N_25022,N_23012,N_22779);
xor U25023 (N_25023,N_23169,N_23833);
nand U25024 (N_25024,N_23564,N_23490);
nor U25025 (N_25025,N_23691,N_23420);
nor U25026 (N_25026,N_22695,N_23633);
and U25027 (N_25027,N_22864,N_23480);
nand U25028 (N_25028,N_22970,N_22594);
xnor U25029 (N_25029,N_22585,N_22718);
or U25030 (N_25030,N_23023,N_23710);
nor U25031 (N_25031,N_23346,N_22955);
xor U25032 (N_25032,N_23942,N_23774);
or U25033 (N_25033,N_23841,N_22814);
nand U25034 (N_25034,N_23981,N_23760);
or U25035 (N_25035,N_23723,N_23443);
xor U25036 (N_25036,N_23620,N_23097);
and U25037 (N_25037,N_23385,N_23394);
or U25038 (N_25038,N_23813,N_22593);
nand U25039 (N_25039,N_23561,N_22831);
xnor U25040 (N_25040,N_23395,N_22587);
nand U25041 (N_25041,N_22983,N_23084);
xor U25042 (N_25042,N_23851,N_22862);
nand U25043 (N_25043,N_23185,N_23747);
xnor U25044 (N_25044,N_23077,N_22673);
nor U25045 (N_25045,N_22569,N_22853);
and U25046 (N_25046,N_23986,N_22989);
and U25047 (N_25047,N_22877,N_23219);
nor U25048 (N_25048,N_23957,N_23504);
and U25049 (N_25049,N_23882,N_22932);
or U25050 (N_25050,N_23129,N_23930);
or U25051 (N_25051,N_23234,N_23019);
nor U25052 (N_25052,N_23755,N_23796);
xor U25053 (N_25053,N_22863,N_23580);
and U25054 (N_25054,N_23483,N_23654);
xnor U25055 (N_25055,N_22804,N_22847);
and U25056 (N_25056,N_23445,N_23702);
nor U25057 (N_25057,N_23377,N_23923);
nor U25058 (N_25058,N_23213,N_23671);
or U25059 (N_25059,N_23923,N_23003);
and U25060 (N_25060,N_23645,N_23949);
xnor U25061 (N_25061,N_23475,N_22584);
and U25062 (N_25062,N_22581,N_23907);
and U25063 (N_25063,N_23219,N_22712);
nor U25064 (N_25064,N_23185,N_22933);
or U25065 (N_25065,N_23347,N_23844);
nand U25066 (N_25066,N_22915,N_22995);
xor U25067 (N_25067,N_22599,N_22956);
or U25068 (N_25068,N_23391,N_22915);
nor U25069 (N_25069,N_22851,N_23988);
nor U25070 (N_25070,N_22532,N_23564);
and U25071 (N_25071,N_22510,N_23775);
and U25072 (N_25072,N_23984,N_23719);
nor U25073 (N_25073,N_22591,N_23057);
and U25074 (N_25074,N_22687,N_22811);
nand U25075 (N_25075,N_22914,N_22589);
nand U25076 (N_25076,N_23648,N_22951);
xnor U25077 (N_25077,N_23554,N_23660);
or U25078 (N_25078,N_23067,N_22837);
or U25079 (N_25079,N_23547,N_22744);
xor U25080 (N_25080,N_23960,N_22746);
xnor U25081 (N_25081,N_22795,N_22790);
or U25082 (N_25082,N_23929,N_23142);
xnor U25083 (N_25083,N_23741,N_23405);
nand U25084 (N_25084,N_23918,N_23916);
nand U25085 (N_25085,N_23441,N_23246);
or U25086 (N_25086,N_23753,N_23471);
nor U25087 (N_25087,N_23111,N_22643);
and U25088 (N_25088,N_22531,N_23248);
nor U25089 (N_25089,N_23689,N_23186);
and U25090 (N_25090,N_22835,N_22540);
and U25091 (N_25091,N_22932,N_22904);
nand U25092 (N_25092,N_23713,N_23915);
nor U25093 (N_25093,N_23663,N_23007);
xor U25094 (N_25094,N_23009,N_23847);
nor U25095 (N_25095,N_23120,N_23180);
nor U25096 (N_25096,N_23657,N_23454);
xnor U25097 (N_25097,N_23613,N_22607);
xnor U25098 (N_25098,N_23503,N_23852);
and U25099 (N_25099,N_22826,N_23814);
or U25100 (N_25100,N_22862,N_23212);
and U25101 (N_25101,N_23036,N_23958);
xor U25102 (N_25102,N_23289,N_23967);
xnor U25103 (N_25103,N_23712,N_23793);
and U25104 (N_25104,N_23289,N_23797);
xor U25105 (N_25105,N_23044,N_22603);
and U25106 (N_25106,N_23427,N_23987);
or U25107 (N_25107,N_23207,N_23891);
nor U25108 (N_25108,N_23687,N_23506);
nand U25109 (N_25109,N_23989,N_22889);
xnor U25110 (N_25110,N_23066,N_23731);
nor U25111 (N_25111,N_23373,N_23853);
xnor U25112 (N_25112,N_22539,N_23558);
or U25113 (N_25113,N_22811,N_23016);
nand U25114 (N_25114,N_23047,N_23074);
nand U25115 (N_25115,N_23859,N_23652);
and U25116 (N_25116,N_23404,N_23338);
and U25117 (N_25117,N_23915,N_22837);
and U25118 (N_25118,N_23665,N_22906);
and U25119 (N_25119,N_23284,N_22830);
nand U25120 (N_25120,N_23297,N_22730);
nand U25121 (N_25121,N_23781,N_23249);
or U25122 (N_25122,N_22533,N_23021);
or U25123 (N_25123,N_22968,N_22907);
and U25124 (N_25124,N_23829,N_23352);
xnor U25125 (N_25125,N_22757,N_23094);
xnor U25126 (N_25126,N_23508,N_23542);
xor U25127 (N_25127,N_23488,N_23595);
and U25128 (N_25128,N_23742,N_22595);
or U25129 (N_25129,N_22907,N_23777);
or U25130 (N_25130,N_23279,N_23064);
nor U25131 (N_25131,N_23144,N_22533);
or U25132 (N_25132,N_23803,N_23244);
and U25133 (N_25133,N_23798,N_22892);
nand U25134 (N_25134,N_23381,N_23367);
or U25135 (N_25135,N_23298,N_23189);
nand U25136 (N_25136,N_23779,N_23604);
or U25137 (N_25137,N_23670,N_23173);
xor U25138 (N_25138,N_23634,N_23100);
xor U25139 (N_25139,N_23376,N_22830);
xnor U25140 (N_25140,N_22987,N_22662);
nor U25141 (N_25141,N_23920,N_23846);
or U25142 (N_25142,N_23009,N_22924);
nand U25143 (N_25143,N_22866,N_22643);
nand U25144 (N_25144,N_22919,N_23016);
or U25145 (N_25145,N_23194,N_23564);
or U25146 (N_25146,N_23330,N_22712);
or U25147 (N_25147,N_23970,N_23323);
xor U25148 (N_25148,N_22631,N_22875);
or U25149 (N_25149,N_23823,N_23363);
or U25150 (N_25150,N_22886,N_22926);
nor U25151 (N_25151,N_22646,N_23973);
or U25152 (N_25152,N_22844,N_23894);
nand U25153 (N_25153,N_23916,N_23056);
nor U25154 (N_25154,N_23437,N_22792);
xor U25155 (N_25155,N_23619,N_23469);
nand U25156 (N_25156,N_23131,N_22936);
nor U25157 (N_25157,N_23051,N_23616);
and U25158 (N_25158,N_22630,N_23313);
nor U25159 (N_25159,N_23505,N_23899);
and U25160 (N_25160,N_23349,N_22531);
nand U25161 (N_25161,N_23353,N_23879);
nor U25162 (N_25162,N_23931,N_22713);
xor U25163 (N_25163,N_22819,N_23863);
nor U25164 (N_25164,N_23563,N_23576);
or U25165 (N_25165,N_23254,N_23998);
xor U25166 (N_25166,N_23844,N_23527);
xnor U25167 (N_25167,N_22941,N_23552);
or U25168 (N_25168,N_22902,N_23215);
or U25169 (N_25169,N_23181,N_23273);
xnor U25170 (N_25170,N_22818,N_23842);
nor U25171 (N_25171,N_23458,N_23488);
nor U25172 (N_25172,N_23856,N_23780);
and U25173 (N_25173,N_22938,N_23207);
nand U25174 (N_25174,N_23061,N_22863);
or U25175 (N_25175,N_22967,N_23328);
nor U25176 (N_25176,N_23127,N_23141);
or U25177 (N_25177,N_22825,N_23333);
and U25178 (N_25178,N_23445,N_23081);
xor U25179 (N_25179,N_23871,N_22951);
or U25180 (N_25180,N_22542,N_23425);
nor U25181 (N_25181,N_23697,N_23756);
xor U25182 (N_25182,N_23119,N_23844);
and U25183 (N_25183,N_23839,N_22589);
or U25184 (N_25184,N_23260,N_23918);
and U25185 (N_25185,N_23964,N_22567);
nor U25186 (N_25186,N_23938,N_23200);
nor U25187 (N_25187,N_23231,N_22706);
xnor U25188 (N_25188,N_23460,N_22770);
and U25189 (N_25189,N_22828,N_23243);
xor U25190 (N_25190,N_23042,N_22772);
xnor U25191 (N_25191,N_22669,N_22808);
or U25192 (N_25192,N_23303,N_23625);
and U25193 (N_25193,N_23604,N_22909);
or U25194 (N_25194,N_22968,N_23346);
and U25195 (N_25195,N_23704,N_22705);
nand U25196 (N_25196,N_23291,N_23941);
or U25197 (N_25197,N_22674,N_23905);
xnor U25198 (N_25198,N_23574,N_23165);
nand U25199 (N_25199,N_23897,N_23117);
xnor U25200 (N_25200,N_23118,N_23820);
nor U25201 (N_25201,N_23102,N_22758);
and U25202 (N_25202,N_22855,N_22548);
or U25203 (N_25203,N_23952,N_23324);
nand U25204 (N_25204,N_22957,N_23273);
nand U25205 (N_25205,N_23762,N_23871);
xnor U25206 (N_25206,N_23916,N_22620);
nor U25207 (N_25207,N_23536,N_23276);
nand U25208 (N_25208,N_23684,N_22703);
nor U25209 (N_25209,N_22673,N_23962);
nand U25210 (N_25210,N_23613,N_23297);
or U25211 (N_25211,N_23695,N_23225);
nor U25212 (N_25212,N_22574,N_23958);
and U25213 (N_25213,N_22725,N_23127);
nand U25214 (N_25214,N_23834,N_22574);
nor U25215 (N_25215,N_23825,N_23832);
or U25216 (N_25216,N_23000,N_23965);
xor U25217 (N_25217,N_22597,N_23888);
nor U25218 (N_25218,N_23577,N_23556);
xor U25219 (N_25219,N_22708,N_23173);
xor U25220 (N_25220,N_23587,N_23638);
and U25221 (N_25221,N_22676,N_23023);
nand U25222 (N_25222,N_22904,N_23514);
and U25223 (N_25223,N_23179,N_22813);
and U25224 (N_25224,N_23194,N_22698);
nand U25225 (N_25225,N_23625,N_22643);
or U25226 (N_25226,N_23882,N_23726);
nand U25227 (N_25227,N_22959,N_23811);
and U25228 (N_25228,N_22854,N_22582);
and U25229 (N_25229,N_23631,N_22527);
and U25230 (N_25230,N_22768,N_23178);
or U25231 (N_25231,N_23413,N_22504);
nor U25232 (N_25232,N_23231,N_23064);
nand U25233 (N_25233,N_23134,N_22519);
nor U25234 (N_25234,N_23733,N_22783);
nand U25235 (N_25235,N_23368,N_23766);
or U25236 (N_25236,N_23714,N_23733);
and U25237 (N_25237,N_23111,N_23095);
and U25238 (N_25238,N_22797,N_23826);
nor U25239 (N_25239,N_23885,N_22784);
or U25240 (N_25240,N_23774,N_23641);
or U25241 (N_25241,N_22998,N_22625);
xor U25242 (N_25242,N_22757,N_23306);
or U25243 (N_25243,N_22997,N_23759);
nand U25244 (N_25244,N_23776,N_23417);
and U25245 (N_25245,N_22847,N_23058);
nor U25246 (N_25246,N_23811,N_23372);
and U25247 (N_25247,N_23060,N_22910);
or U25248 (N_25248,N_22683,N_23813);
nand U25249 (N_25249,N_23255,N_22836);
and U25250 (N_25250,N_23114,N_23265);
and U25251 (N_25251,N_22733,N_22923);
and U25252 (N_25252,N_22950,N_23616);
or U25253 (N_25253,N_23666,N_22602);
nand U25254 (N_25254,N_23874,N_23876);
and U25255 (N_25255,N_23915,N_22566);
nor U25256 (N_25256,N_22985,N_23889);
nor U25257 (N_25257,N_23730,N_22950);
and U25258 (N_25258,N_23505,N_22780);
and U25259 (N_25259,N_23699,N_23458);
or U25260 (N_25260,N_23956,N_23754);
nand U25261 (N_25261,N_23180,N_22830);
nand U25262 (N_25262,N_22952,N_23680);
nor U25263 (N_25263,N_22592,N_23083);
xnor U25264 (N_25264,N_22776,N_23620);
xnor U25265 (N_25265,N_23189,N_22531);
and U25266 (N_25266,N_23435,N_22603);
xor U25267 (N_25267,N_22697,N_23542);
xor U25268 (N_25268,N_23450,N_22824);
and U25269 (N_25269,N_22983,N_23699);
and U25270 (N_25270,N_22962,N_23130);
xor U25271 (N_25271,N_23395,N_23788);
nand U25272 (N_25272,N_23050,N_23801);
nor U25273 (N_25273,N_22528,N_22563);
xnor U25274 (N_25274,N_23208,N_23897);
xor U25275 (N_25275,N_23496,N_23149);
nand U25276 (N_25276,N_22565,N_23105);
nor U25277 (N_25277,N_23519,N_23650);
nand U25278 (N_25278,N_22984,N_23133);
xor U25279 (N_25279,N_22702,N_23017);
or U25280 (N_25280,N_22744,N_23487);
and U25281 (N_25281,N_22571,N_23867);
nor U25282 (N_25282,N_22822,N_22746);
and U25283 (N_25283,N_23364,N_22890);
nand U25284 (N_25284,N_23231,N_23220);
nand U25285 (N_25285,N_22681,N_23605);
xnor U25286 (N_25286,N_23238,N_23979);
or U25287 (N_25287,N_23559,N_23713);
or U25288 (N_25288,N_23118,N_23309);
xor U25289 (N_25289,N_23191,N_23416);
and U25290 (N_25290,N_23124,N_23120);
or U25291 (N_25291,N_23813,N_23417);
nor U25292 (N_25292,N_22900,N_22646);
xor U25293 (N_25293,N_22573,N_23919);
and U25294 (N_25294,N_23634,N_23807);
or U25295 (N_25295,N_22672,N_23816);
and U25296 (N_25296,N_22727,N_22917);
nor U25297 (N_25297,N_23265,N_23698);
and U25298 (N_25298,N_23919,N_22746);
xor U25299 (N_25299,N_23313,N_22502);
nor U25300 (N_25300,N_23734,N_23525);
nor U25301 (N_25301,N_23342,N_22633);
nor U25302 (N_25302,N_23980,N_23260);
nor U25303 (N_25303,N_23807,N_23165);
nor U25304 (N_25304,N_22660,N_23437);
nor U25305 (N_25305,N_23775,N_23165);
or U25306 (N_25306,N_22884,N_23146);
nor U25307 (N_25307,N_23776,N_23114);
xor U25308 (N_25308,N_23301,N_23857);
nor U25309 (N_25309,N_22663,N_22661);
nand U25310 (N_25310,N_22955,N_23702);
nor U25311 (N_25311,N_22748,N_23436);
and U25312 (N_25312,N_23691,N_23538);
and U25313 (N_25313,N_23466,N_23509);
and U25314 (N_25314,N_23879,N_23116);
and U25315 (N_25315,N_22681,N_23671);
and U25316 (N_25316,N_22693,N_23396);
xnor U25317 (N_25317,N_23685,N_23581);
nor U25318 (N_25318,N_23895,N_23178);
and U25319 (N_25319,N_23065,N_23604);
xnor U25320 (N_25320,N_22877,N_23445);
nand U25321 (N_25321,N_22924,N_23397);
and U25322 (N_25322,N_22700,N_23923);
nor U25323 (N_25323,N_23117,N_23839);
or U25324 (N_25324,N_23990,N_22804);
xnor U25325 (N_25325,N_23107,N_23451);
nor U25326 (N_25326,N_22886,N_23022);
nand U25327 (N_25327,N_23023,N_22860);
and U25328 (N_25328,N_23322,N_22888);
and U25329 (N_25329,N_23543,N_23940);
nand U25330 (N_25330,N_22725,N_23855);
or U25331 (N_25331,N_23078,N_22800);
and U25332 (N_25332,N_23047,N_23208);
and U25333 (N_25333,N_23304,N_23035);
nor U25334 (N_25334,N_23943,N_23753);
or U25335 (N_25335,N_22776,N_23929);
xor U25336 (N_25336,N_23632,N_23707);
and U25337 (N_25337,N_22712,N_22816);
and U25338 (N_25338,N_23393,N_22565);
and U25339 (N_25339,N_23379,N_23722);
nand U25340 (N_25340,N_23773,N_22968);
nor U25341 (N_25341,N_23087,N_22582);
and U25342 (N_25342,N_23905,N_23368);
nor U25343 (N_25343,N_23389,N_23294);
nand U25344 (N_25344,N_23213,N_23027);
or U25345 (N_25345,N_23549,N_22509);
xnor U25346 (N_25346,N_23864,N_23454);
nand U25347 (N_25347,N_22863,N_23241);
and U25348 (N_25348,N_23572,N_22961);
or U25349 (N_25349,N_23621,N_23905);
and U25350 (N_25350,N_22901,N_23615);
or U25351 (N_25351,N_23626,N_23734);
and U25352 (N_25352,N_23879,N_23279);
xnor U25353 (N_25353,N_22561,N_22801);
nor U25354 (N_25354,N_22809,N_22858);
nand U25355 (N_25355,N_22791,N_23389);
nor U25356 (N_25356,N_23322,N_23946);
and U25357 (N_25357,N_23096,N_22701);
xnor U25358 (N_25358,N_23470,N_23978);
or U25359 (N_25359,N_23604,N_22533);
xor U25360 (N_25360,N_22596,N_22877);
nor U25361 (N_25361,N_22539,N_22770);
xnor U25362 (N_25362,N_23541,N_23839);
or U25363 (N_25363,N_22573,N_22877);
xnor U25364 (N_25364,N_23687,N_23301);
nand U25365 (N_25365,N_23242,N_23215);
or U25366 (N_25366,N_23234,N_23844);
nor U25367 (N_25367,N_23367,N_23119);
xnor U25368 (N_25368,N_22752,N_23254);
nand U25369 (N_25369,N_22811,N_22876);
nand U25370 (N_25370,N_23213,N_23896);
nor U25371 (N_25371,N_23049,N_23513);
nand U25372 (N_25372,N_23228,N_23780);
or U25373 (N_25373,N_23771,N_23656);
nor U25374 (N_25374,N_23501,N_23066);
nor U25375 (N_25375,N_22705,N_22840);
or U25376 (N_25376,N_23744,N_23726);
and U25377 (N_25377,N_23282,N_22856);
nor U25378 (N_25378,N_23596,N_23410);
xnor U25379 (N_25379,N_23240,N_23772);
xnor U25380 (N_25380,N_23175,N_22513);
xor U25381 (N_25381,N_22986,N_22981);
and U25382 (N_25382,N_23394,N_23764);
nand U25383 (N_25383,N_22908,N_23555);
nor U25384 (N_25384,N_22794,N_23498);
or U25385 (N_25385,N_23868,N_23832);
or U25386 (N_25386,N_23128,N_23598);
nor U25387 (N_25387,N_23759,N_22691);
and U25388 (N_25388,N_23855,N_23275);
nand U25389 (N_25389,N_23900,N_22571);
and U25390 (N_25390,N_23555,N_22701);
nand U25391 (N_25391,N_23545,N_23104);
xor U25392 (N_25392,N_23399,N_22822);
nor U25393 (N_25393,N_23396,N_23743);
or U25394 (N_25394,N_22582,N_23285);
and U25395 (N_25395,N_22918,N_23096);
nand U25396 (N_25396,N_23532,N_23388);
nor U25397 (N_25397,N_23842,N_23373);
and U25398 (N_25398,N_23868,N_23043);
xor U25399 (N_25399,N_23780,N_22512);
nand U25400 (N_25400,N_22707,N_22816);
or U25401 (N_25401,N_23906,N_23026);
and U25402 (N_25402,N_23238,N_22932);
xnor U25403 (N_25403,N_23362,N_23367);
nand U25404 (N_25404,N_23283,N_23097);
or U25405 (N_25405,N_23721,N_23102);
or U25406 (N_25406,N_23144,N_22522);
xor U25407 (N_25407,N_22713,N_23358);
or U25408 (N_25408,N_23722,N_23077);
nand U25409 (N_25409,N_23705,N_22861);
nand U25410 (N_25410,N_22663,N_22584);
or U25411 (N_25411,N_23453,N_23366);
xnor U25412 (N_25412,N_22885,N_22611);
and U25413 (N_25413,N_23343,N_22845);
and U25414 (N_25414,N_23120,N_23484);
xnor U25415 (N_25415,N_22553,N_23920);
xnor U25416 (N_25416,N_23369,N_23868);
xnor U25417 (N_25417,N_22510,N_23338);
nor U25418 (N_25418,N_23691,N_23456);
nand U25419 (N_25419,N_23675,N_23331);
or U25420 (N_25420,N_23338,N_22592);
xnor U25421 (N_25421,N_22755,N_22838);
nand U25422 (N_25422,N_23816,N_23396);
and U25423 (N_25423,N_22793,N_23733);
nor U25424 (N_25424,N_23959,N_23736);
or U25425 (N_25425,N_22731,N_23862);
and U25426 (N_25426,N_23975,N_23305);
nand U25427 (N_25427,N_23221,N_23024);
nand U25428 (N_25428,N_22566,N_22654);
xor U25429 (N_25429,N_23355,N_23391);
nand U25430 (N_25430,N_23968,N_23679);
nand U25431 (N_25431,N_23258,N_23988);
or U25432 (N_25432,N_23306,N_23115);
and U25433 (N_25433,N_23605,N_23732);
nand U25434 (N_25434,N_23499,N_23967);
and U25435 (N_25435,N_23779,N_23707);
and U25436 (N_25436,N_23652,N_23034);
nand U25437 (N_25437,N_23996,N_23611);
or U25438 (N_25438,N_23685,N_22521);
and U25439 (N_25439,N_23115,N_22957);
nor U25440 (N_25440,N_22859,N_22976);
and U25441 (N_25441,N_23883,N_23787);
and U25442 (N_25442,N_22811,N_23984);
and U25443 (N_25443,N_22898,N_23737);
nor U25444 (N_25444,N_23690,N_23387);
and U25445 (N_25445,N_23399,N_23612);
or U25446 (N_25446,N_23321,N_23258);
or U25447 (N_25447,N_23019,N_22842);
nor U25448 (N_25448,N_23691,N_22551);
nand U25449 (N_25449,N_23978,N_22560);
or U25450 (N_25450,N_23018,N_23635);
or U25451 (N_25451,N_23765,N_22620);
nand U25452 (N_25452,N_22761,N_23180);
and U25453 (N_25453,N_23062,N_22987);
and U25454 (N_25454,N_23360,N_22970);
and U25455 (N_25455,N_23073,N_22663);
xor U25456 (N_25456,N_22706,N_23619);
nor U25457 (N_25457,N_23630,N_23871);
or U25458 (N_25458,N_23412,N_23253);
xor U25459 (N_25459,N_23969,N_22583);
or U25460 (N_25460,N_23338,N_22887);
xor U25461 (N_25461,N_22960,N_23308);
xor U25462 (N_25462,N_22566,N_22828);
and U25463 (N_25463,N_23855,N_23139);
and U25464 (N_25464,N_23457,N_23650);
nor U25465 (N_25465,N_23165,N_23253);
and U25466 (N_25466,N_23296,N_22867);
or U25467 (N_25467,N_23811,N_23953);
nor U25468 (N_25468,N_23470,N_22858);
nor U25469 (N_25469,N_22749,N_23356);
or U25470 (N_25470,N_23812,N_23044);
nand U25471 (N_25471,N_23629,N_23812);
xor U25472 (N_25472,N_22586,N_22759);
or U25473 (N_25473,N_22665,N_22841);
nand U25474 (N_25474,N_23717,N_23720);
and U25475 (N_25475,N_22688,N_22653);
nand U25476 (N_25476,N_22751,N_22641);
nand U25477 (N_25477,N_23417,N_23843);
nand U25478 (N_25478,N_23635,N_22825);
xnor U25479 (N_25479,N_22811,N_23460);
nand U25480 (N_25480,N_22557,N_22803);
nand U25481 (N_25481,N_23464,N_22515);
nand U25482 (N_25482,N_22862,N_22515);
or U25483 (N_25483,N_22896,N_23956);
nand U25484 (N_25484,N_22953,N_23557);
nand U25485 (N_25485,N_23449,N_23172);
or U25486 (N_25486,N_23119,N_22627);
nor U25487 (N_25487,N_22650,N_22888);
nand U25488 (N_25488,N_22504,N_22947);
nor U25489 (N_25489,N_23507,N_22512);
or U25490 (N_25490,N_23897,N_22748);
and U25491 (N_25491,N_23899,N_22604);
and U25492 (N_25492,N_22518,N_22582);
nand U25493 (N_25493,N_23222,N_23364);
nand U25494 (N_25494,N_23982,N_23796);
and U25495 (N_25495,N_23081,N_23501);
or U25496 (N_25496,N_23615,N_22525);
and U25497 (N_25497,N_23535,N_23534);
nor U25498 (N_25498,N_22556,N_23813);
or U25499 (N_25499,N_23995,N_22965);
nor U25500 (N_25500,N_25243,N_24360);
and U25501 (N_25501,N_24626,N_24432);
or U25502 (N_25502,N_24888,N_25020);
xnor U25503 (N_25503,N_24291,N_25039);
nand U25504 (N_25504,N_25366,N_24470);
nor U25505 (N_25505,N_24545,N_25419);
and U25506 (N_25506,N_24928,N_24905);
nand U25507 (N_25507,N_24944,N_24904);
and U25508 (N_25508,N_24224,N_24912);
nor U25509 (N_25509,N_24317,N_25403);
nor U25510 (N_25510,N_25188,N_25335);
xnor U25511 (N_25511,N_24733,N_24711);
nand U25512 (N_25512,N_25014,N_24040);
or U25513 (N_25513,N_24346,N_25393);
or U25514 (N_25514,N_24319,N_25061);
or U25515 (N_25515,N_24960,N_24191);
or U25516 (N_25516,N_24443,N_25030);
and U25517 (N_25517,N_25086,N_24018);
or U25518 (N_25518,N_24195,N_24741);
or U25519 (N_25519,N_24981,N_24431);
and U25520 (N_25520,N_24369,N_24838);
nor U25521 (N_25521,N_24720,N_24921);
xnor U25522 (N_25522,N_24868,N_24024);
xor U25523 (N_25523,N_24528,N_25161);
and U25524 (N_25524,N_25068,N_24990);
nand U25525 (N_25525,N_25043,N_25448);
nor U25526 (N_25526,N_25186,N_24232);
or U25527 (N_25527,N_24650,N_24541);
xor U25528 (N_25528,N_24568,N_24493);
nor U25529 (N_25529,N_24764,N_24697);
nor U25530 (N_25530,N_25128,N_24729);
nor U25531 (N_25531,N_24550,N_24236);
or U25532 (N_25532,N_24544,N_24211);
and U25533 (N_25533,N_25180,N_24495);
nand U25534 (N_25534,N_24925,N_24419);
or U25535 (N_25535,N_25492,N_24297);
or U25536 (N_25536,N_24758,N_24952);
xor U25537 (N_25537,N_24248,N_24060);
nor U25538 (N_25538,N_24813,N_24200);
xor U25539 (N_25539,N_24931,N_25425);
xor U25540 (N_25540,N_25050,N_24983);
nor U25541 (N_25541,N_24546,N_25034);
nand U25542 (N_25542,N_24889,N_24103);
nand U25543 (N_25543,N_24595,N_24911);
or U25544 (N_25544,N_24599,N_24272);
nor U25545 (N_25545,N_25088,N_25238);
nor U25546 (N_25546,N_24907,N_24365);
and U25547 (N_25547,N_25191,N_25071);
nor U25548 (N_25548,N_25377,N_25170);
nand U25549 (N_25549,N_25135,N_24779);
and U25550 (N_25550,N_25320,N_24352);
or U25551 (N_25551,N_24472,N_25137);
and U25552 (N_25552,N_24615,N_24149);
xnor U25553 (N_25553,N_24994,N_24454);
and U25554 (N_25554,N_24050,N_24334);
nor U25555 (N_25555,N_25465,N_24581);
nor U25556 (N_25556,N_25110,N_24806);
or U25557 (N_25557,N_24636,N_24832);
xnor U25558 (N_25558,N_24028,N_25368);
or U25559 (N_25559,N_24034,N_24869);
nand U25560 (N_25560,N_24481,N_24513);
xnor U25561 (N_25561,N_24266,N_25350);
nor U25562 (N_25562,N_24458,N_25459);
and U25563 (N_25563,N_24142,N_25358);
xor U25564 (N_25564,N_24135,N_25312);
or U25565 (N_25565,N_24392,N_25233);
and U25566 (N_25566,N_25227,N_24575);
or U25567 (N_25567,N_25055,N_25434);
and U25568 (N_25568,N_24939,N_24844);
or U25569 (N_25569,N_25232,N_24430);
nand U25570 (N_25570,N_24309,N_24000);
nand U25571 (N_25571,N_25131,N_24294);
and U25572 (N_25572,N_24478,N_24988);
and U25573 (N_25573,N_25431,N_24221);
nand U25574 (N_25574,N_24916,N_24755);
or U25575 (N_25575,N_24756,N_25417);
nand U25576 (N_25576,N_24652,N_25246);
xor U25577 (N_25577,N_25437,N_24721);
nand U25578 (N_25578,N_25079,N_25105);
and U25579 (N_25579,N_25252,N_25416);
and U25580 (N_25580,N_24753,N_24933);
or U25581 (N_25581,N_24605,N_24601);
nand U25582 (N_25582,N_24465,N_25331);
nand U25583 (N_25583,N_24304,N_25478);
nand U25584 (N_25584,N_25152,N_24915);
and U25585 (N_25585,N_25494,N_24836);
or U25586 (N_25586,N_24835,N_25495);
or U25587 (N_25587,N_24161,N_24416);
nor U25588 (N_25588,N_24453,N_25375);
nor U25589 (N_25589,N_24728,N_25329);
xnor U25590 (N_25590,N_24563,N_24260);
nor U25591 (N_25591,N_24680,N_25165);
xnor U25592 (N_25592,N_24945,N_25120);
and U25593 (N_25593,N_24937,N_24795);
and U25594 (N_25594,N_24651,N_24433);
nor U25595 (N_25595,N_24824,N_24850);
xnor U25596 (N_25596,N_25420,N_25209);
or U25597 (N_25597,N_25053,N_24586);
nor U25598 (N_25598,N_25452,N_24063);
or U25599 (N_25599,N_24131,N_25119);
and U25600 (N_25600,N_24705,N_24903);
nand U25601 (N_25601,N_25353,N_24881);
and U25602 (N_25602,N_24318,N_24398);
xnor U25603 (N_25603,N_24876,N_24415);
xnor U25604 (N_25604,N_24910,N_25107);
xnor U25605 (N_25605,N_24308,N_24709);
and U25606 (N_25606,N_24136,N_24509);
and U25607 (N_25607,N_24421,N_24716);
nor U25608 (N_25608,N_24106,N_24742);
or U25609 (N_25609,N_24022,N_24490);
nand U25610 (N_25610,N_24328,N_25025);
nand U25611 (N_25611,N_24710,N_25456);
nand U25612 (N_25612,N_24642,N_24547);
and U25613 (N_25613,N_24153,N_24234);
xnor U25614 (N_25614,N_24166,N_24088);
xor U25615 (N_25615,N_25241,N_24214);
or U25616 (N_25616,N_24897,N_24021);
or U25617 (N_25617,N_25266,N_24965);
nand U25618 (N_25618,N_24796,N_24781);
and U25619 (N_25619,N_25340,N_25258);
nand U25620 (N_25620,N_25482,N_24237);
and U25621 (N_25621,N_24357,N_24202);
nand U25622 (N_25622,N_24583,N_25468);
and U25623 (N_25623,N_24763,N_25112);
or U25624 (N_25624,N_24124,N_24985);
and U25625 (N_25625,N_25369,N_24084);
xor U25626 (N_25626,N_25432,N_25248);
xnor U25627 (N_25627,N_24657,N_24207);
or U25628 (N_25628,N_24263,N_24856);
xnor U25629 (N_25629,N_25346,N_25361);
nand U25630 (N_25630,N_25015,N_25294);
nand U25631 (N_25631,N_24048,N_24569);
nor U25632 (N_25632,N_24557,N_24479);
xnor U25633 (N_25633,N_24590,N_24695);
or U25634 (N_25634,N_24062,N_24058);
nand U25635 (N_25635,N_24957,N_24873);
nand U25636 (N_25636,N_25488,N_25210);
xnor U25637 (N_25637,N_24288,N_25096);
and U25638 (N_25638,N_24497,N_24420);
nor U25639 (N_25639,N_24193,N_25485);
nor U25640 (N_25640,N_24393,N_25264);
xnor U25641 (N_25641,N_24144,N_24205);
or U25642 (N_25642,N_24402,N_24025);
nand U25643 (N_25643,N_25024,N_24573);
and U25644 (N_25644,N_24165,N_25155);
and U25645 (N_25645,N_24871,N_25153);
xnor U25646 (N_25646,N_25136,N_24380);
or U25647 (N_25647,N_24370,N_25006);
nor U25648 (N_25648,N_24723,N_24313);
or U25649 (N_25649,N_24030,N_24774);
or U25650 (N_25650,N_25144,N_24958);
nor U25651 (N_25651,N_25216,N_25038);
xnor U25652 (N_25652,N_24858,N_24891);
nor U25653 (N_25653,N_24158,N_25115);
xor U25654 (N_25654,N_24638,N_25443);
nor U25655 (N_25655,N_24770,N_24475);
and U25656 (N_25656,N_24228,N_25262);
xnor U25657 (N_25657,N_25285,N_24932);
xnor U25658 (N_25658,N_24117,N_25111);
and U25659 (N_25659,N_24769,N_25421);
xnor U25660 (N_25660,N_25464,N_25057);
xnor U25661 (N_25661,N_25117,N_24137);
nor U25662 (N_25662,N_24198,N_24310);
or U25663 (N_25663,N_24512,N_24484);
nor U25664 (N_25664,N_24071,N_25220);
xnor U25665 (N_25665,N_24353,N_24209);
and U25666 (N_25666,N_24622,N_25173);
or U25667 (N_25667,N_24732,N_25479);
nor U25668 (N_25668,N_24655,N_25245);
nor U25669 (N_25669,N_25001,N_25439);
xor U25670 (N_25670,N_24505,N_25183);
or U25671 (N_25671,N_24726,N_24196);
xnor U25672 (N_25672,N_24056,N_24081);
xnor U25673 (N_25673,N_25208,N_24285);
nor U25674 (N_25674,N_25424,N_25225);
and U25675 (N_25675,N_24108,N_24148);
and U25676 (N_25676,N_25101,N_24610);
or U25677 (N_25677,N_24511,N_24621);
nor U25678 (N_25678,N_24345,N_24978);
or U25679 (N_25679,N_25298,N_24820);
and U25680 (N_25680,N_24768,N_25185);
xnor U25681 (N_25681,N_24699,N_25125);
nor U25682 (N_25682,N_25196,N_25189);
and U25683 (N_25683,N_24337,N_24080);
or U25684 (N_25684,N_25132,N_24589);
nor U25685 (N_25685,N_24325,N_24133);
nand U25686 (N_25686,N_24061,N_25436);
and U25687 (N_25687,N_24864,N_25476);
nor U25688 (N_25688,N_24016,N_24001);
or U25689 (N_25689,N_24999,N_24535);
nor U25690 (N_25690,N_25159,N_24611);
nor U25691 (N_25691,N_25442,N_24284);
nor U25692 (N_25692,N_24239,N_25281);
nand U25693 (N_25693,N_24576,N_24023);
xnor U25694 (N_25694,N_25092,N_24872);
or U25695 (N_25695,N_24130,N_24316);
nor U25696 (N_25696,N_25077,N_24390);
nand U25697 (N_25697,N_24703,N_25386);
and U25698 (N_25698,N_24155,N_25041);
nand U25699 (N_25699,N_25156,N_25106);
or U25700 (N_25700,N_25267,N_25451);
xor U25701 (N_25701,N_24087,N_24792);
nor U25702 (N_25702,N_24687,N_24953);
and U25703 (N_25703,N_24322,N_24057);
nand U25704 (N_25704,N_25414,N_24410);
or U25705 (N_25705,N_24855,N_24930);
and U25706 (N_25706,N_24292,N_25192);
and U25707 (N_25707,N_24669,N_25357);
and U25708 (N_25708,N_24900,N_25108);
nand U25709 (N_25709,N_25483,N_25205);
nor U25710 (N_25710,N_24307,N_24176);
or U25711 (N_25711,N_24554,N_24097);
or U25712 (N_25712,N_24217,N_25103);
nand U25713 (N_25713,N_24185,N_24388);
nor U25714 (N_25714,N_24139,N_24104);
nand U25715 (N_25715,N_25201,N_24457);
and U25716 (N_25716,N_25102,N_24029);
xnor U25717 (N_25717,N_25027,N_25422);
nand U25718 (N_25718,N_24092,N_24616);
and U25719 (N_25719,N_24004,N_24785);
nand U25720 (N_25720,N_25138,N_24434);
nor U25721 (N_25721,N_24629,N_24093);
xnor U25722 (N_25722,N_24109,N_24242);
nor U25723 (N_25723,N_25171,N_24761);
nand U25724 (N_25724,N_25322,N_24119);
and U25725 (N_25725,N_24805,N_24963);
nand U25726 (N_25726,N_24766,N_24719);
nand U25727 (N_25727,N_25054,N_24306);
nor U25728 (N_25728,N_24448,N_24730);
nor U25729 (N_25729,N_24438,N_24689);
or U25730 (N_25730,N_24518,N_24901);
nand U25731 (N_25731,N_25226,N_25090);
nor U25732 (N_25732,N_24287,N_25244);
nand U25733 (N_25733,N_24987,N_25166);
or U25734 (N_25734,N_24301,N_25072);
xor U25735 (N_25735,N_24258,N_24895);
xnor U25736 (N_25736,N_24678,N_25367);
or U25737 (N_25737,N_25401,N_25059);
and U25738 (N_25738,N_24336,N_25458);
and U25739 (N_25739,N_25430,N_25378);
or U25740 (N_25740,N_24885,N_24140);
nand U25741 (N_25741,N_24134,N_25497);
or U25742 (N_25742,N_24335,N_25113);
xor U25743 (N_25743,N_25299,N_24471);
nor U25744 (N_25744,N_24246,N_25147);
or U25745 (N_25745,N_24095,N_25154);
and U25746 (N_25746,N_24828,N_24101);
and U25747 (N_25747,N_25063,N_25118);
nand U25748 (N_25748,N_24673,N_24992);
and U25749 (N_25749,N_24100,N_24170);
or U25750 (N_25750,N_25036,N_25217);
xnor U25751 (N_25751,N_25418,N_24338);
nand U25752 (N_25752,N_24521,N_24647);
and U25753 (N_25753,N_24842,N_24789);
nor U25754 (N_25754,N_24967,N_25017);
nor U25755 (N_25755,N_24418,N_25130);
xor U25756 (N_25756,N_24231,N_24261);
nor U25757 (N_25757,N_24073,N_24537);
nor U25758 (N_25758,N_25388,N_25134);
xnor U25759 (N_25759,N_25409,N_25018);
and U25760 (N_25760,N_24808,N_24487);
nor U25761 (N_25761,N_25268,N_24278);
or U25762 (N_25762,N_25394,N_24997);
or U25763 (N_25763,N_24840,N_25163);
and U25764 (N_25764,N_24754,N_25237);
nor U25765 (N_25765,N_25215,N_24381);
and U25766 (N_25766,N_24233,N_25275);
or U25767 (N_25767,N_24055,N_24982);
or U25768 (N_25768,N_24520,N_25008);
xnor U25769 (N_25769,N_25087,N_24624);
or U25770 (N_25770,N_24943,N_24208);
or U25771 (N_25771,N_24035,N_24845);
or U25772 (N_25772,N_25257,N_24833);
or U25773 (N_25773,N_24603,N_24851);
or U25774 (N_25774,N_24302,N_24964);
nor U25775 (N_25775,N_24935,N_24694);
xnor U25776 (N_25776,N_24225,N_24817);
nand U25777 (N_25777,N_24474,N_24641);
nor U25778 (N_25778,N_24303,N_25129);
nor U25779 (N_25779,N_24251,N_24067);
nor U25780 (N_25780,N_24582,N_24556);
nor U25781 (N_25781,N_24950,N_24387);
nor U25782 (N_25782,N_24026,N_24909);
nand U25783 (N_25783,N_25391,N_24252);
xnor U25784 (N_25784,N_25318,N_24534);
nor U25785 (N_25785,N_24857,N_24070);
and U25786 (N_25786,N_25169,N_25460);
nor U25787 (N_25787,N_25028,N_25198);
nand U25788 (N_25788,N_24163,N_25250);
or U25789 (N_25789,N_24525,N_24600);
nor U25790 (N_25790,N_25289,N_24422);
nor U25791 (N_25791,N_24934,N_24218);
xor U25792 (N_25792,N_24374,N_24745);
and U25793 (N_25793,N_24017,N_25178);
xor U25794 (N_25794,N_24184,N_25440);
nand U25795 (N_25795,N_25195,N_24240);
nand U25796 (N_25796,N_24608,N_24244);
or U25797 (N_25797,N_24450,N_24899);
nand U25798 (N_25798,N_24739,N_25074);
nor U25799 (N_25799,N_24423,N_24107);
nor U25800 (N_25800,N_24002,N_24675);
xor U25801 (N_25801,N_24938,N_24323);
nand U25802 (N_25802,N_24507,N_24922);
nor U25803 (N_25803,N_24020,N_24271);
or U25804 (N_25804,N_24807,N_24046);
and U25805 (N_25805,N_25031,N_24386);
or U25806 (N_25806,N_24363,N_25313);
nor U25807 (N_25807,N_24923,N_25387);
nor U25808 (N_25808,N_25370,N_25235);
xor U25809 (N_25809,N_24286,N_25284);
nand U25810 (N_25810,N_24333,N_24414);
or U25811 (N_25811,N_24847,N_24690);
nand U25812 (N_25812,N_24849,N_24492);
or U25813 (N_25813,N_24666,N_24591);
and U25814 (N_25814,N_25175,N_24778);
nand U25815 (N_25815,N_24391,N_24371);
nand U25816 (N_25816,N_24010,N_24645);
and U25817 (N_25817,N_25247,N_24042);
nand U25818 (N_25818,N_24917,N_24255);
nor U25819 (N_25819,N_25221,N_24648);
and U25820 (N_25820,N_24801,N_24966);
xnor U25821 (N_25821,N_24700,N_25249);
or U25822 (N_25822,N_25306,N_25223);
or U25823 (N_25823,N_25081,N_24826);
or U25824 (N_25824,N_25265,N_24265);
and U25825 (N_25825,N_25260,N_24510);
xor U25826 (N_25826,N_24654,N_24052);
xor U25827 (N_25827,N_25080,N_24141);
xor U25828 (N_25828,N_25301,N_25012);
xnor U25829 (N_25829,N_24327,N_25202);
nor U25830 (N_25830,N_25213,N_24947);
or U25831 (N_25831,N_24853,N_24822);
or U25832 (N_25832,N_24339,N_24037);
or U25833 (N_25833,N_24105,N_25474);
and U25834 (N_25834,N_25314,N_25168);
nor U25835 (N_25835,N_24775,N_25098);
nand U25836 (N_25836,N_25450,N_25190);
and U25837 (N_25837,N_24969,N_24955);
xor U25838 (N_25838,N_25157,N_25083);
or U25839 (N_25839,N_24727,N_24598);
xor U25840 (N_25840,N_24749,N_24968);
and U25841 (N_25841,N_24574,N_25219);
nor U25842 (N_25842,N_25381,N_24126);
or U25843 (N_25843,N_25104,N_24526);
xnor U25844 (N_25844,N_25067,N_25073);
nor U25845 (N_25845,N_24083,N_24201);
xor U25846 (N_25846,N_25373,N_24315);
xnor U25847 (N_25847,N_24725,N_24777);
or U25848 (N_25848,N_24204,N_25032);
and U25849 (N_25849,N_24787,N_25415);
nand U25850 (N_25850,N_24441,N_24444);
nor U25851 (N_25851,N_24003,N_24708);
or U25852 (N_25852,N_24522,N_25214);
nor U25853 (N_25853,N_25179,N_24829);
nand U25854 (N_25854,N_24486,N_24340);
nand U25855 (N_25855,N_24321,N_25280);
xor U25856 (N_25856,N_25022,N_24115);
nor U25857 (N_25857,N_24283,N_25172);
nand U25858 (N_25858,N_24262,N_24098);
or U25859 (N_25859,N_24913,N_24919);
and U25860 (N_25860,N_24489,N_25286);
xnor U25861 (N_25861,N_24382,N_24397);
nor U25862 (N_25862,N_25097,N_24750);
or U25863 (N_25863,N_25349,N_25007);
nand U25864 (N_25864,N_24250,N_24800);
xor U25865 (N_25865,N_24394,N_24311);
nand U25866 (N_25866,N_24890,N_24408);
nor U25867 (N_25867,N_24906,N_24395);
and U25868 (N_25868,N_25288,N_24685);
nand U25869 (N_25869,N_25033,N_24435);
and U25870 (N_25870,N_25484,N_24956);
and U25871 (N_25871,N_24171,N_24693);
nor U25872 (N_25872,N_24918,N_24314);
nor U25873 (N_25873,N_24926,N_24082);
nor U25874 (N_25874,N_25141,N_24502);
nor U25875 (N_25875,N_25473,N_25078);
nand U25876 (N_25876,N_24661,N_24143);
and U25877 (N_25877,N_24878,N_25402);
xor U25878 (N_25878,N_24500,N_25251);
nand U25879 (N_25879,N_25274,N_25405);
nand U25880 (N_25880,N_24114,N_24993);
xnor U25881 (N_25881,N_24846,N_24235);
and U25882 (N_25882,N_24366,N_25095);
or U25883 (N_25883,N_24722,N_24210);
xnor U25884 (N_25884,N_24305,N_24530);
nor U25885 (N_25885,N_24663,N_25023);
nor U25886 (N_25886,N_24219,N_25142);
or U25887 (N_25887,N_25046,N_24632);
and U25888 (N_25888,N_24399,N_25290);
xnor U25889 (N_25889,N_24008,N_24861);
nand U25890 (N_25890,N_25158,N_24412);
xnor U25891 (N_25891,N_24914,N_24032);
nand U25892 (N_25892,N_24068,N_24536);
and U25893 (N_25893,N_25000,N_24480);
and U25894 (N_25894,N_24112,N_24998);
or U25895 (N_25895,N_25004,N_24403);
nor U25896 (N_25896,N_24679,N_24782);
nand U25897 (N_25897,N_25311,N_24194);
nand U25898 (N_25898,N_25362,N_24216);
xnor U25899 (N_25899,N_24122,N_25317);
xnor U25900 (N_25900,N_24767,N_25447);
nor U25901 (N_25901,N_24118,N_24962);
and U25902 (N_25902,N_25489,N_25376);
or U25903 (N_25903,N_24047,N_24893);
nand U25904 (N_25904,N_24883,N_24449);
or U25905 (N_25905,N_25399,N_25099);
nor U25906 (N_25906,N_24662,N_24186);
and U25907 (N_25907,N_24543,N_24190);
nand U25908 (N_25908,N_25021,N_24094);
nor U25909 (N_25909,N_25199,N_24355);
xor U25910 (N_25910,N_24946,N_25224);
nand U25911 (N_25911,N_25075,N_25374);
nand U25912 (N_25912,N_24159,N_25082);
and U25913 (N_25913,N_24637,N_24404);
and U25914 (N_25914,N_24954,N_24585);
and U25915 (N_25915,N_24887,N_24644);
and U25916 (N_25916,N_24524,N_24772);
nand U25917 (N_25917,N_24762,N_24238);
xnor U25918 (N_25918,N_24494,N_24451);
nand U25919 (N_25919,N_25297,N_24116);
nor U25920 (N_25920,N_24665,N_24974);
or U25921 (N_25921,N_24264,N_25167);
or U25922 (N_25922,N_24848,N_24941);
and U25923 (N_25923,N_25392,N_25446);
nor U25924 (N_25924,N_24863,N_24765);
nand U25925 (N_25925,N_24593,N_24776);
and U25926 (N_25926,N_25239,N_25383);
nand U25927 (N_25927,N_24455,N_25100);
and U25928 (N_25928,N_24596,N_24215);
xnor U25929 (N_25929,N_24014,N_24740);
and U25930 (N_25930,N_24396,N_24731);
nand U25931 (N_25931,N_24870,N_24971);
and U25932 (N_25932,N_24516,N_24614);
nor U25933 (N_25933,N_24332,N_24120);
nor U25934 (N_25934,N_25065,N_25240);
and U25935 (N_25935,N_24167,N_24377);
and U25936 (N_25936,N_24715,N_24169);
and U25937 (N_25937,N_25302,N_24091);
xnor U25938 (N_25938,N_24515,N_24157);
and U25939 (N_25939,N_24677,N_24877);
nand U25940 (N_25940,N_24588,N_24559);
or U25941 (N_25941,N_25457,N_25372);
nor U25942 (N_25942,N_25308,N_24179);
or U25943 (N_25943,N_24633,N_24676);
xor U25944 (N_25944,N_25413,N_24482);
nor U25945 (N_25945,N_24054,N_25019);
xnor U25946 (N_25946,N_24138,N_25332);
and U25947 (N_25947,N_24276,N_24558);
xnor U25948 (N_25948,N_24257,N_24797);
and U25949 (N_25949,N_25364,N_24199);
xnor U25950 (N_25950,N_24975,N_25321);
nor U25951 (N_25951,N_24940,N_25064);
nor U25952 (N_25952,N_25182,N_24439);
nor U25953 (N_25953,N_24446,N_24175);
nand U25954 (N_25954,N_24747,N_24951);
nand U25955 (N_25955,N_25058,N_24627);
xor U25956 (N_25956,N_24929,N_24426);
nand U25957 (N_25957,N_24213,N_25094);
and U25958 (N_25958,N_24223,N_24523);
xor U25959 (N_25959,N_24875,N_24780);
or U25960 (N_25960,N_25160,N_24013);
nor U25961 (N_25961,N_24075,N_25287);
nand U25962 (N_25962,N_24802,N_24936);
and U25963 (N_25963,N_25445,N_24049);
or U25964 (N_25964,N_24348,N_24174);
xnor U25965 (N_25965,N_24701,N_25200);
nand U25966 (N_25966,N_24734,N_24354);
nor U25967 (N_25967,N_24243,N_25319);
or U25968 (N_25968,N_24033,N_24274);
xnor U25969 (N_25969,N_25339,N_25062);
and U25970 (N_25970,N_25109,N_25016);
nand U25971 (N_25971,N_25122,N_24865);
nand U25972 (N_25972,N_24491,N_24656);
or U25973 (N_25973,N_24659,N_25255);
xor U25974 (N_25974,N_24125,N_24096);
and U25975 (N_25975,N_25400,N_24698);
nor U25976 (N_25976,N_25256,N_25408);
and U25977 (N_25977,N_24942,N_24587);
xor U25978 (N_25978,N_24692,N_24538);
xor U25979 (N_25979,N_24473,N_24841);
and U25980 (N_25980,N_25035,N_25231);
xnor U25981 (N_25981,N_25139,N_25384);
xnor U25982 (N_25982,N_24086,N_24065);
xor U25983 (N_25983,N_24406,N_24192);
nor U25984 (N_25984,N_24417,N_25176);
nor U25985 (N_25985,N_24821,N_25229);
nor U25986 (N_25986,N_24757,N_24226);
xor U25987 (N_25987,N_25276,N_24460);
xnor U25988 (N_25988,N_24059,N_24672);
and U25989 (N_25989,N_24247,N_25145);
xor U25990 (N_25990,N_25222,N_25469);
xnor U25991 (N_25991,N_24811,N_24639);
nor U25992 (N_25992,N_24533,N_25480);
or U25993 (N_25993,N_24241,N_25491);
xor U25994 (N_25994,N_25493,N_25441);
and U25995 (N_25995,N_24180,N_24702);
and U25996 (N_25996,N_25070,N_24799);
nand U25997 (N_25997,N_24362,N_24111);
or U25998 (N_25998,N_24977,N_24331);
xnor U25999 (N_25999,N_24445,N_25354);
nand U26000 (N_26000,N_24634,N_24385);
or U26001 (N_26001,N_24548,N_24290);
and U26002 (N_26002,N_24364,N_24784);
or U26003 (N_26003,N_24076,N_25228);
and U26004 (N_26004,N_24839,N_25151);
or U26005 (N_26005,N_25333,N_25150);
nor U26006 (N_26006,N_24074,N_24612);
nor U26007 (N_26007,N_24631,N_25300);
xnor U26008 (N_26008,N_24123,N_24467);
or U26009 (N_26009,N_25148,N_24625);
and U26010 (N_26010,N_25466,N_24688);
and U26011 (N_26011,N_24469,N_24718);
or U26012 (N_26012,N_25496,N_25093);
or U26013 (N_26013,N_24592,N_25292);
nand U26014 (N_26014,N_24009,N_25037);
and U26015 (N_26015,N_25123,N_24299);
nand U26016 (N_26016,N_25056,N_24580);
nor U26017 (N_26017,N_25143,N_24329);
nor U26018 (N_26018,N_24358,N_25271);
nor U26019 (N_26019,N_24866,N_24902);
nor U26020 (N_26020,N_24653,N_24831);
or U26021 (N_26021,N_25382,N_24649);
xor U26022 (N_26022,N_24532,N_25444);
xnor U26023 (N_26023,N_24830,N_25218);
xnor U26024 (N_26024,N_25325,N_24517);
nand U26025 (N_26025,N_25486,N_25426);
or U26026 (N_26026,N_24704,N_24724);
nand U26027 (N_26027,N_24085,N_25365);
nor U26028 (N_26028,N_24476,N_24594);
xor U26029 (N_26029,N_24862,N_24686);
or U26030 (N_26030,N_24597,N_24706);
nand U26031 (N_26031,N_24005,N_24976);
nor U26032 (N_26032,N_24671,N_24553);
nand U26033 (N_26033,N_24972,N_24442);
nor U26034 (N_26034,N_24043,N_24019);
xnor U26035 (N_26035,N_24463,N_24270);
nor U26036 (N_26036,N_25029,N_25498);
nor U26037 (N_26037,N_24168,N_25140);
nor U26038 (N_26038,N_24350,N_24300);
or U26039 (N_26039,N_24578,N_24810);
xnor U26040 (N_26040,N_25360,N_25323);
and U26041 (N_26041,N_24892,N_24011);
nor U26042 (N_26042,N_25475,N_24424);
xnor U26043 (N_26043,N_24401,N_24737);
nor U26044 (N_26044,N_24356,N_24584);
and U26045 (N_26045,N_24640,N_24496);
nand U26046 (N_26046,N_24110,N_25471);
or U26047 (N_26047,N_24039,N_24256);
xor U26048 (N_26048,N_25344,N_24786);
or U26049 (N_26049,N_24320,N_25277);
nor U26050 (N_26050,N_25005,N_24407);
and U26051 (N_26051,N_24425,N_24660);
and U26052 (N_26052,N_24613,N_24979);
or U26053 (N_26053,N_25091,N_25009);
or U26054 (N_26054,N_24189,N_24162);
nand U26055 (N_26055,N_25410,N_25211);
nand U26056 (N_26056,N_25395,N_24409);
or U26057 (N_26057,N_25042,N_25310);
or U26058 (N_26058,N_25455,N_24771);
nand U26059 (N_26059,N_25194,N_25291);
nand U26060 (N_26060,N_25114,N_25385);
nand U26061 (N_26061,N_24053,N_25380);
and U26062 (N_26062,N_25203,N_24289);
xor U26063 (N_26063,N_24735,N_24156);
nor U26064 (N_26064,N_25328,N_24330);
xnor U26065 (N_26065,N_24220,N_24326);
nand U26066 (N_26066,N_25272,N_24712);
nand U26067 (N_26067,N_24268,N_24324);
xor U26068 (N_26068,N_24312,N_24759);
xnor U26069 (N_26069,N_24531,N_24503);
nand U26070 (N_26070,N_24164,N_25206);
nor U26071 (N_26071,N_25487,N_25084);
or U26072 (N_26072,N_24884,N_24461);
nor U26073 (N_26073,N_24743,N_24436);
nand U26074 (N_26074,N_24411,N_24178);
nor U26075 (N_26075,N_25003,N_25398);
nor U26076 (N_26076,N_24882,N_24249);
nor U26077 (N_26077,N_24400,N_24012);
xnor U26078 (N_26078,N_25282,N_24986);
or U26079 (N_26079,N_24540,N_25047);
nor U26080 (N_26080,N_25293,N_24485);
and U26081 (N_26081,N_25359,N_25499);
nand U26082 (N_26082,N_25013,N_24160);
or U26083 (N_26083,N_24867,N_24379);
and U26084 (N_26084,N_24717,N_25406);
and U26085 (N_26085,N_25303,N_24670);
and U26086 (N_26086,N_25348,N_24619);
or U26087 (N_26087,N_24514,N_25454);
and U26088 (N_26088,N_24383,N_24646);
xnor U26089 (N_26089,N_25467,N_24466);
or U26090 (N_26090,N_25263,N_24519);
and U26091 (N_26091,N_25010,N_24714);
nand U26092 (N_26092,N_25040,N_24859);
and U26093 (N_26093,N_24007,N_25044);
and U26094 (N_26094,N_24015,N_24079);
nand U26095 (N_26095,N_25127,N_24121);
and U26096 (N_26096,N_25124,N_25428);
and U26097 (N_26097,N_24375,N_24529);
xor U26098 (N_26098,N_25026,N_24549);
nand U26099 (N_26099,N_24607,N_25146);
or U26100 (N_26100,N_25342,N_24874);
xor U26101 (N_26101,N_24267,N_25411);
nor U26102 (N_26102,N_24077,N_24683);
and U26103 (N_26103,N_24182,N_25253);
xor U26104 (N_26104,N_24681,N_25315);
nor U26105 (N_26105,N_25207,N_24468);
xnor U26106 (N_26106,N_24227,N_25181);
and U26107 (N_26107,N_24027,N_24696);
nand U26108 (N_26108,N_24295,N_25162);
and U26109 (N_26109,N_25347,N_24230);
and U26110 (N_26110,N_24823,N_25133);
or U26111 (N_26111,N_24794,N_24506);
nor U26112 (N_26112,N_24102,N_24560);
or U26113 (N_26113,N_24282,N_25316);
nand U26114 (N_26114,N_25345,N_25177);
or U26115 (N_26115,N_24552,N_24229);
nand U26116 (N_26116,N_24347,N_24539);
nand U26117 (N_26117,N_25296,N_25472);
or U26118 (N_26118,N_25069,N_24744);
nand U26119 (N_26119,N_24602,N_24961);
nor U26120 (N_26120,N_24854,N_25397);
and U26121 (N_26121,N_24041,N_24154);
or U26122 (N_26122,N_24405,N_25230);
nand U26123 (N_26123,N_24886,N_24793);
and U26124 (N_26124,N_25336,N_24452);
xnor U26125 (N_26125,N_24151,N_24825);
nand U26126 (N_26126,N_24989,N_25278);
nor U26127 (N_26127,N_25254,N_25462);
nand U26128 (N_26128,N_25273,N_25076);
nor U26129 (N_26129,N_25184,N_25334);
nor U26130 (N_26130,N_25121,N_24501);
or U26131 (N_26131,N_25356,N_24896);
or U26132 (N_26132,N_24389,N_24376);
and U26133 (N_26133,N_25438,N_24222);
and U26134 (N_26134,N_24372,N_24606);
nor U26135 (N_26135,N_24738,N_25389);
and U26136 (N_26136,N_24664,N_24948);
or U26137 (N_26137,N_25371,N_24038);
or U26138 (N_26138,N_24384,N_25174);
nand U26139 (N_26139,N_24150,N_25149);
xnor U26140 (N_26140,N_24643,N_24682);
or U26141 (N_26141,N_24736,N_25423);
nor U26142 (N_26142,N_24635,N_25407);
nand U26143 (N_26143,N_24924,N_24804);
and U26144 (N_26144,N_24275,N_24812);
or U26145 (N_26145,N_24751,N_24984);
nand U26146 (N_26146,N_24973,N_25066);
nor U26147 (N_26147,N_25261,N_24342);
and U26148 (N_26148,N_24064,N_24212);
nand U26149 (N_26149,N_25352,N_24341);
xnor U26150 (N_26150,N_24880,N_24031);
or U26151 (N_26151,N_24072,N_24277);
nor U26152 (N_26152,N_24609,N_24843);
nand U26153 (N_26153,N_25269,N_25490);
and U26154 (N_26154,N_24051,N_25412);
and U26155 (N_26155,N_24129,N_24783);
nand U26156 (N_26156,N_24127,N_24760);
nor U26157 (N_26157,N_24089,N_24748);
and U26158 (N_26158,N_24564,N_24970);
and U26159 (N_26159,N_25449,N_24296);
or U26160 (N_26160,N_25327,N_25351);
nand U26161 (N_26161,N_24628,N_24837);
nor U26162 (N_26162,N_25355,N_24620);
nor U26163 (N_26163,N_24344,N_24254);
xor U26164 (N_26164,N_25379,N_24790);
and U26165 (N_26165,N_25011,N_24281);
or U26166 (N_26166,N_25404,N_24440);
or U26167 (N_26167,N_24488,N_24368);
or U26168 (N_26168,N_24498,N_24099);
nor U26169 (N_26169,N_24188,N_25187);
xnor U26170 (N_26170,N_24788,N_25481);
nand U26171 (N_26171,N_25470,N_24044);
nor U26172 (N_26172,N_25197,N_25236);
and U26173 (N_26173,N_24570,N_24773);
and U26174 (N_26174,N_24181,N_24527);
nor U26175 (N_26175,N_25204,N_24667);
nor U26176 (N_26176,N_24707,N_24036);
xor U26177 (N_26177,N_24980,N_24090);
nand U26178 (N_26178,N_24604,N_24852);
and U26179 (N_26179,N_24464,N_25307);
nand U26180 (N_26180,N_24920,N_25089);
nand U26181 (N_26181,N_24145,N_24566);
nand U26182 (N_26182,N_25051,N_25433);
or U26183 (N_26183,N_24343,N_25295);
or U26184 (N_26184,N_24561,N_24551);
xor U26185 (N_26185,N_24819,N_24618);
and U26186 (N_26186,N_24197,N_24658);
nand U26187 (N_26187,N_24555,N_24152);
nand U26188 (N_26188,N_24577,N_24113);
xnor U26189 (N_26189,N_24045,N_25343);
or U26190 (N_26190,N_25283,N_24508);
xor U26191 (N_26191,N_24959,N_24879);
nand U26192 (N_26192,N_24827,N_25304);
nor U26193 (N_26193,N_24630,N_24860);
xnor U26194 (N_26194,N_25326,N_25341);
and U26195 (N_26195,N_25052,N_24269);
and U26196 (N_26196,N_24949,N_24579);
and U26197 (N_26197,N_24542,N_24206);
or U26198 (N_26198,N_24427,N_25048);
nand U26199 (N_26199,N_24146,N_24279);
and U26200 (N_26200,N_24809,N_24617);
or U26201 (N_26201,N_24894,N_25049);
nand U26202 (N_26202,N_24815,N_24177);
xnor U26203 (N_26203,N_24413,N_24429);
nor U26204 (N_26204,N_25427,N_25126);
nand U26205 (N_26205,N_25242,N_24814);
and U26206 (N_26206,N_25324,N_25477);
nor U26207 (N_26207,N_25164,N_24791);
xor U26208 (N_26208,N_25116,N_25193);
nor U26209 (N_26209,N_25337,N_24373);
xor U26210 (N_26210,N_24571,N_24746);
nand U26211 (N_26211,N_25259,N_24361);
xor U26212 (N_26212,N_24172,N_24273);
nand U26213 (N_26213,N_25330,N_25060);
xor U26214 (N_26214,N_24456,N_24996);
nor U26215 (N_26215,N_24991,N_24066);
nor U26216 (N_26216,N_24713,N_24818);
nor U26217 (N_26217,N_25429,N_24483);
and U26218 (N_26218,N_25309,N_24803);
nand U26219 (N_26219,N_25234,N_24691);
nor U26220 (N_26220,N_25085,N_24259);
and U26221 (N_26221,N_24203,N_24995);
nand U26222 (N_26222,N_24674,N_25396);
and U26223 (N_26223,N_25363,N_24816);
nor U26224 (N_26224,N_24447,N_24565);
or U26225 (N_26225,N_24187,N_24684);
and U26226 (N_26226,N_24359,N_25453);
and U26227 (N_26227,N_24351,N_24293);
nor U26228 (N_26228,N_24183,N_24477);
nand U26229 (N_26229,N_24437,N_24128);
xor U26230 (N_26230,N_24567,N_24459);
nand U26231 (N_26231,N_25435,N_24245);
xnor U26232 (N_26232,N_24572,N_24349);
xnor U26233 (N_26233,N_25270,N_24006);
nor U26234 (N_26234,N_24499,N_25390);
and U26235 (N_26235,N_24908,N_25045);
nand U26236 (N_26236,N_24078,N_24562);
nand U26237 (N_26237,N_25305,N_25002);
or U26238 (N_26238,N_24132,N_24834);
or U26239 (N_26239,N_24147,N_24798);
or U26240 (N_26240,N_24428,N_24173);
nor U26241 (N_26241,N_24298,N_24927);
nor U26242 (N_26242,N_24253,N_25461);
or U26243 (N_26243,N_24462,N_24623);
and U26244 (N_26244,N_24504,N_24668);
xnor U26245 (N_26245,N_24752,N_24367);
and U26246 (N_26246,N_24898,N_25212);
and U26247 (N_26247,N_24280,N_25463);
nor U26248 (N_26248,N_24378,N_25338);
and U26249 (N_26249,N_24069,N_25279);
xnor U26250 (N_26250,N_24300,N_24715);
nand U26251 (N_26251,N_24700,N_24174);
xnor U26252 (N_26252,N_24000,N_24140);
and U26253 (N_26253,N_24825,N_25085);
or U26254 (N_26254,N_24220,N_25336);
nand U26255 (N_26255,N_24476,N_24946);
and U26256 (N_26256,N_25082,N_24068);
nor U26257 (N_26257,N_24589,N_25104);
or U26258 (N_26258,N_25390,N_24881);
xor U26259 (N_26259,N_25414,N_25469);
or U26260 (N_26260,N_24298,N_25233);
nand U26261 (N_26261,N_24318,N_25325);
nand U26262 (N_26262,N_24606,N_25291);
nor U26263 (N_26263,N_24357,N_24893);
or U26264 (N_26264,N_24056,N_24881);
nor U26265 (N_26265,N_24271,N_24949);
nor U26266 (N_26266,N_24112,N_25246);
and U26267 (N_26267,N_25234,N_24114);
and U26268 (N_26268,N_25096,N_24816);
or U26269 (N_26269,N_25372,N_25384);
nand U26270 (N_26270,N_24506,N_24648);
nor U26271 (N_26271,N_25095,N_24647);
nor U26272 (N_26272,N_24159,N_24960);
nand U26273 (N_26273,N_25128,N_24324);
nor U26274 (N_26274,N_25453,N_25229);
nand U26275 (N_26275,N_25412,N_24254);
or U26276 (N_26276,N_24470,N_25185);
nor U26277 (N_26277,N_24050,N_24514);
and U26278 (N_26278,N_25171,N_24386);
xor U26279 (N_26279,N_25244,N_24356);
or U26280 (N_26280,N_25336,N_24829);
or U26281 (N_26281,N_25324,N_25191);
nor U26282 (N_26282,N_24532,N_24927);
or U26283 (N_26283,N_24975,N_25294);
and U26284 (N_26284,N_24950,N_24588);
nor U26285 (N_26285,N_24772,N_24266);
nor U26286 (N_26286,N_24980,N_24701);
xor U26287 (N_26287,N_24969,N_24373);
and U26288 (N_26288,N_24024,N_24249);
xnor U26289 (N_26289,N_24617,N_25481);
or U26290 (N_26290,N_24881,N_25019);
or U26291 (N_26291,N_24690,N_24203);
xor U26292 (N_26292,N_24553,N_24969);
xnor U26293 (N_26293,N_24228,N_25009);
xor U26294 (N_26294,N_24388,N_24093);
and U26295 (N_26295,N_24203,N_25347);
nand U26296 (N_26296,N_24365,N_24673);
and U26297 (N_26297,N_25248,N_24598);
nor U26298 (N_26298,N_24112,N_24968);
and U26299 (N_26299,N_24428,N_24743);
or U26300 (N_26300,N_24018,N_24468);
and U26301 (N_26301,N_24434,N_25295);
xnor U26302 (N_26302,N_24323,N_25362);
nand U26303 (N_26303,N_25401,N_24389);
nand U26304 (N_26304,N_24795,N_25018);
nor U26305 (N_26305,N_25216,N_24190);
nor U26306 (N_26306,N_25005,N_24030);
nor U26307 (N_26307,N_24663,N_25072);
and U26308 (N_26308,N_24297,N_24902);
nor U26309 (N_26309,N_25262,N_25289);
and U26310 (N_26310,N_25111,N_24581);
nand U26311 (N_26311,N_24258,N_25144);
nor U26312 (N_26312,N_25142,N_25478);
and U26313 (N_26313,N_25005,N_25258);
nand U26314 (N_26314,N_24404,N_24434);
or U26315 (N_26315,N_24076,N_24786);
or U26316 (N_26316,N_24358,N_24534);
nand U26317 (N_26317,N_25287,N_24859);
nor U26318 (N_26318,N_24009,N_24886);
and U26319 (N_26319,N_24589,N_24801);
and U26320 (N_26320,N_24253,N_24509);
or U26321 (N_26321,N_25075,N_24783);
xnor U26322 (N_26322,N_24222,N_24106);
or U26323 (N_26323,N_25392,N_25375);
xnor U26324 (N_26324,N_24344,N_25231);
or U26325 (N_26325,N_25323,N_24255);
nor U26326 (N_26326,N_24555,N_25126);
nand U26327 (N_26327,N_25121,N_24321);
and U26328 (N_26328,N_25261,N_25250);
xor U26329 (N_26329,N_25131,N_24222);
and U26330 (N_26330,N_25066,N_25457);
or U26331 (N_26331,N_24367,N_24545);
nor U26332 (N_26332,N_24928,N_24211);
or U26333 (N_26333,N_24504,N_24179);
and U26334 (N_26334,N_24832,N_24208);
xor U26335 (N_26335,N_24322,N_24925);
nor U26336 (N_26336,N_24769,N_24209);
and U26337 (N_26337,N_24390,N_25344);
and U26338 (N_26338,N_25160,N_24489);
or U26339 (N_26339,N_24994,N_24991);
or U26340 (N_26340,N_25492,N_25413);
nor U26341 (N_26341,N_25413,N_25419);
or U26342 (N_26342,N_25225,N_25140);
and U26343 (N_26343,N_25279,N_24229);
nand U26344 (N_26344,N_24292,N_24663);
nand U26345 (N_26345,N_25428,N_24389);
nand U26346 (N_26346,N_24493,N_24765);
or U26347 (N_26347,N_25346,N_24663);
nor U26348 (N_26348,N_24920,N_25392);
nor U26349 (N_26349,N_24415,N_24691);
nor U26350 (N_26350,N_25346,N_24288);
and U26351 (N_26351,N_25016,N_25012);
nand U26352 (N_26352,N_25057,N_24269);
and U26353 (N_26353,N_25456,N_25352);
and U26354 (N_26354,N_24531,N_24703);
nand U26355 (N_26355,N_24630,N_24701);
or U26356 (N_26356,N_25383,N_25407);
xnor U26357 (N_26357,N_24335,N_25043);
nand U26358 (N_26358,N_24168,N_25412);
and U26359 (N_26359,N_24711,N_24889);
or U26360 (N_26360,N_24455,N_25151);
or U26361 (N_26361,N_25173,N_25140);
xor U26362 (N_26362,N_25179,N_24140);
nor U26363 (N_26363,N_24056,N_24987);
nor U26364 (N_26364,N_24626,N_24741);
nand U26365 (N_26365,N_24982,N_25009);
xnor U26366 (N_26366,N_24089,N_24053);
nand U26367 (N_26367,N_25080,N_25167);
nand U26368 (N_26368,N_24702,N_24616);
and U26369 (N_26369,N_24158,N_24119);
xnor U26370 (N_26370,N_24620,N_25401);
and U26371 (N_26371,N_24674,N_25049);
nand U26372 (N_26372,N_24018,N_24833);
nand U26373 (N_26373,N_24680,N_24716);
nand U26374 (N_26374,N_25459,N_25286);
nand U26375 (N_26375,N_24720,N_24470);
or U26376 (N_26376,N_25078,N_24507);
nand U26377 (N_26377,N_24607,N_24376);
nor U26378 (N_26378,N_24792,N_24997);
nand U26379 (N_26379,N_24196,N_24752);
nor U26380 (N_26380,N_24072,N_25349);
or U26381 (N_26381,N_24433,N_24634);
xnor U26382 (N_26382,N_24254,N_25056);
and U26383 (N_26383,N_24663,N_25382);
and U26384 (N_26384,N_24329,N_24999);
and U26385 (N_26385,N_24413,N_24729);
and U26386 (N_26386,N_25099,N_25159);
and U26387 (N_26387,N_24400,N_25464);
xnor U26388 (N_26388,N_24272,N_25225);
nand U26389 (N_26389,N_24301,N_24322);
and U26390 (N_26390,N_24892,N_24516);
xor U26391 (N_26391,N_25497,N_25190);
nor U26392 (N_26392,N_24717,N_25352);
or U26393 (N_26393,N_24194,N_24747);
or U26394 (N_26394,N_24910,N_24825);
or U26395 (N_26395,N_24682,N_25264);
and U26396 (N_26396,N_24019,N_25168);
and U26397 (N_26397,N_24973,N_25053);
or U26398 (N_26398,N_24257,N_24085);
xnor U26399 (N_26399,N_24609,N_25494);
xor U26400 (N_26400,N_25064,N_24763);
nand U26401 (N_26401,N_24923,N_24812);
and U26402 (N_26402,N_25271,N_24729);
or U26403 (N_26403,N_24561,N_25217);
or U26404 (N_26404,N_24044,N_25328);
and U26405 (N_26405,N_25482,N_24182);
nor U26406 (N_26406,N_25025,N_24944);
xor U26407 (N_26407,N_24837,N_25473);
and U26408 (N_26408,N_25280,N_25046);
and U26409 (N_26409,N_24031,N_24074);
xor U26410 (N_26410,N_24465,N_24108);
and U26411 (N_26411,N_25240,N_24216);
nor U26412 (N_26412,N_24576,N_24710);
and U26413 (N_26413,N_24516,N_24469);
xor U26414 (N_26414,N_24953,N_25405);
or U26415 (N_26415,N_25100,N_24301);
xor U26416 (N_26416,N_25102,N_24605);
or U26417 (N_26417,N_24550,N_24563);
nor U26418 (N_26418,N_24751,N_25058);
or U26419 (N_26419,N_24408,N_24738);
nor U26420 (N_26420,N_24202,N_24850);
xnor U26421 (N_26421,N_25008,N_25202);
or U26422 (N_26422,N_24463,N_25255);
xnor U26423 (N_26423,N_24473,N_24529);
or U26424 (N_26424,N_24152,N_25473);
nand U26425 (N_26425,N_24902,N_24218);
nor U26426 (N_26426,N_24609,N_24256);
xnor U26427 (N_26427,N_24455,N_24057);
nor U26428 (N_26428,N_24278,N_25391);
nor U26429 (N_26429,N_24911,N_24176);
xor U26430 (N_26430,N_24352,N_25197);
or U26431 (N_26431,N_25185,N_25147);
xnor U26432 (N_26432,N_25065,N_24320);
nand U26433 (N_26433,N_24119,N_24810);
nand U26434 (N_26434,N_24020,N_25465);
nor U26435 (N_26435,N_24037,N_25153);
and U26436 (N_26436,N_24037,N_24214);
or U26437 (N_26437,N_25330,N_25335);
nand U26438 (N_26438,N_25497,N_24911);
nor U26439 (N_26439,N_24919,N_24859);
nand U26440 (N_26440,N_25162,N_25130);
or U26441 (N_26441,N_25131,N_24854);
nor U26442 (N_26442,N_25282,N_24837);
and U26443 (N_26443,N_25124,N_24432);
nor U26444 (N_26444,N_24546,N_24867);
or U26445 (N_26445,N_24555,N_24156);
xnor U26446 (N_26446,N_25405,N_25424);
nand U26447 (N_26447,N_24270,N_25338);
nor U26448 (N_26448,N_25434,N_24802);
nor U26449 (N_26449,N_24805,N_25445);
and U26450 (N_26450,N_24205,N_25491);
or U26451 (N_26451,N_25059,N_24176);
xnor U26452 (N_26452,N_24848,N_25477);
and U26453 (N_26453,N_24337,N_24129);
xnor U26454 (N_26454,N_24212,N_24196);
or U26455 (N_26455,N_24051,N_24673);
nand U26456 (N_26456,N_24873,N_24606);
or U26457 (N_26457,N_24899,N_24893);
xor U26458 (N_26458,N_24562,N_24605);
and U26459 (N_26459,N_24787,N_24064);
xor U26460 (N_26460,N_24105,N_25364);
nand U26461 (N_26461,N_24956,N_24581);
nand U26462 (N_26462,N_25228,N_24952);
xnor U26463 (N_26463,N_25254,N_24667);
nand U26464 (N_26464,N_25306,N_24012);
nor U26465 (N_26465,N_24798,N_24533);
nand U26466 (N_26466,N_24713,N_24863);
or U26467 (N_26467,N_24399,N_24943);
nand U26468 (N_26468,N_24533,N_24321);
and U26469 (N_26469,N_25385,N_25318);
and U26470 (N_26470,N_24917,N_24723);
and U26471 (N_26471,N_24430,N_25031);
and U26472 (N_26472,N_25483,N_24835);
nand U26473 (N_26473,N_24382,N_24998);
and U26474 (N_26474,N_25040,N_24694);
nor U26475 (N_26475,N_24315,N_25492);
and U26476 (N_26476,N_24933,N_25048);
nor U26477 (N_26477,N_25391,N_25290);
xor U26478 (N_26478,N_24939,N_24649);
nor U26479 (N_26479,N_25025,N_24422);
and U26480 (N_26480,N_25386,N_24292);
xnor U26481 (N_26481,N_24592,N_25263);
nand U26482 (N_26482,N_25303,N_24089);
or U26483 (N_26483,N_24319,N_24195);
nor U26484 (N_26484,N_24598,N_25214);
and U26485 (N_26485,N_25278,N_24067);
or U26486 (N_26486,N_24889,N_24791);
xnor U26487 (N_26487,N_24618,N_25285);
xor U26488 (N_26488,N_25077,N_25481);
nand U26489 (N_26489,N_25353,N_24078);
xnor U26490 (N_26490,N_24221,N_24414);
nor U26491 (N_26491,N_25164,N_25374);
xor U26492 (N_26492,N_25347,N_25088);
xnor U26493 (N_26493,N_24801,N_25181);
and U26494 (N_26494,N_24821,N_24881);
xnor U26495 (N_26495,N_24146,N_25036);
xor U26496 (N_26496,N_24846,N_24880);
nor U26497 (N_26497,N_25132,N_24629);
nand U26498 (N_26498,N_24073,N_25480);
nor U26499 (N_26499,N_24394,N_24161);
xnor U26500 (N_26500,N_25259,N_25410);
and U26501 (N_26501,N_24483,N_24017);
xor U26502 (N_26502,N_24617,N_24104);
xnor U26503 (N_26503,N_24102,N_25416);
xor U26504 (N_26504,N_24397,N_24016);
nor U26505 (N_26505,N_25162,N_24351);
or U26506 (N_26506,N_24861,N_24774);
xnor U26507 (N_26507,N_25022,N_25248);
nor U26508 (N_26508,N_25336,N_24677);
xnor U26509 (N_26509,N_24335,N_24714);
or U26510 (N_26510,N_24351,N_24751);
nand U26511 (N_26511,N_24797,N_24383);
and U26512 (N_26512,N_24074,N_24585);
or U26513 (N_26513,N_24021,N_24664);
and U26514 (N_26514,N_24684,N_24941);
or U26515 (N_26515,N_24949,N_24800);
nand U26516 (N_26516,N_24404,N_24730);
nor U26517 (N_26517,N_24677,N_24568);
or U26518 (N_26518,N_24909,N_25179);
nor U26519 (N_26519,N_24781,N_25284);
nand U26520 (N_26520,N_24517,N_24381);
nand U26521 (N_26521,N_25244,N_25200);
or U26522 (N_26522,N_24622,N_24039);
nand U26523 (N_26523,N_25117,N_24732);
or U26524 (N_26524,N_24118,N_24921);
or U26525 (N_26525,N_25268,N_25249);
nand U26526 (N_26526,N_24024,N_24749);
or U26527 (N_26527,N_25449,N_24268);
nand U26528 (N_26528,N_24572,N_24519);
nor U26529 (N_26529,N_24141,N_24219);
xnor U26530 (N_26530,N_24880,N_24668);
xor U26531 (N_26531,N_25469,N_25267);
or U26532 (N_26532,N_24618,N_24283);
nor U26533 (N_26533,N_24146,N_24297);
nor U26534 (N_26534,N_25212,N_24817);
xnor U26535 (N_26535,N_24038,N_25304);
xor U26536 (N_26536,N_24268,N_25102);
nand U26537 (N_26537,N_24696,N_24503);
nor U26538 (N_26538,N_25047,N_24063);
nand U26539 (N_26539,N_24014,N_24946);
nand U26540 (N_26540,N_24348,N_24256);
xor U26541 (N_26541,N_24888,N_24009);
and U26542 (N_26542,N_24266,N_25105);
and U26543 (N_26543,N_25494,N_24894);
or U26544 (N_26544,N_24404,N_24289);
and U26545 (N_26545,N_24456,N_25436);
xor U26546 (N_26546,N_24245,N_24788);
nand U26547 (N_26547,N_24055,N_24388);
xor U26548 (N_26548,N_24027,N_24426);
or U26549 (N_26549,N_25203,N_25263);
or U26550 (N_26550,N_24090,N_24595);
or U26551 (N_26551,N_25423,N_25453);
xor U26552 (N_26552,N_25028,N_24644);
or U26553 (N_26553,N_25072,N_24583);
xor U26554 (N_26554,N_24796,N_24348);
or U26555 (N_26555,N_24503,N_24516);
or U26556 (N_26556,N_24864,N_24628);
or U26557 (N_26557,N_24106,N_24240);
xor U26558 (N_26558,N_25271,N_24628);
and U26559 (N_26559,N_24431,N_24911);
nand U26560 (N_26560,N_24874,N_25362);
nor U26561 (N_26561,N_25302,N_25283);
xnor U26562 (N_26562,N_24713,N_24823);
nor U26563 (N_26563,N_25384,N_24041);
xnor U26564 (N_26564,N_24480,N_25065);
nand U26565 (N_26565,N_24584,N_24292);
nand U26566 (N_26566,N_25246,N_24503);
nand U26567 (N_26567,N_24268,N_24986);
nor U26568 (N_26568,N_24742,N_24900);
nor U26569 (N_26569,N_24991,N_25030);
and U26570 (N_26570,N_24444,N_24193);
and U26571 (N_26571,N_24901,N_24722);
and U26572 (N_26572,N_24574,N_25262);
xor U26573 (N_26573,N_24571,N_24902);
nand U26574 (N_26574,N_24944,N_24885);
xnor U26575 (N_26575,N_25064,N_24885);
xor U26576 (N_26576,N_25390,N_25171);
or U26577 (N_26577,N_24020,N_24959);
nand U26578 (N_26578,N_24011,N_24014);
and U26579 (N_26579,N_24325,N_24154);
and U26580 (N_26580,N_24270,N_24397);
nor U26581 (N_26581,N_24599,N_24106);
xnor U26582 (N_26582,N_25480,N_24597);
nand U26583 (N_26583,N_24045,N_24785);
nor U26584 (N_26584,N_24031,N_24300);
xnor U26585 (N_26585,N_25402,N_24400);
nand U26586 (N_26586,N_25363,N_24432);
and U26587 (N_26587,N_25205,N_24458);
xnor U26588 (N_26588,N_24061,N_24440);
xnor U26589 (N_26589,N_24541,N_25323);
nor U26590 (N_26590,N_24086,N_24815);
nand U26591 (N_26591,N_24980,N_24088);
or U26592 (N_26592,N_24021,N_24907);
nand U26593 (N_26593,N_24255,N_25492);
and U26594 (N_26594,N_24026,N_24712);
xor U26595 (N_26595,N_25392,N_25230);
nand U26596 (N_26596,N_25456,N_24587);
or U26597 (N_26597,N_25348,N_25340);
nor U26598 (N_26598,N_25078,N_24812);
xnor U26599 (N_26599,N_25065,N_24635);
nand U26600 (N_26600,N_24077,N_25215);
nor U26601 (N_26601,N_24870,N_25444);
or U26602 (N_26602,N_24691,N_24248);
xor U26603 (N_26603,N_25070,N_24837);
nor U26604 (N_26604,N_25461,N_24992);
nor U26605 (N_26605,N_24698,N_24267);
or U26606 (N_26606,N_24944,N_24356);
or U26607 (N_26607,N_24478,N_24684);
and U26608 (N_26608,N_24044,N_24721);
nor U26609 (N_26609,N_25422,N_25315);
and U26610 (N_26610,N_24230,N_24159);
xor U26611 (N_26611,N_24771,N_25381);
or U26612 (N_26612,N_24911,N_24469);
xor U26613 (N_26613,N_24182,N_25040);
xnor U26614 (N_26614,N_24118,N_24903);
and U26615 (N_26615,N_25376,N_24294);
xnor U26616 (N_26616,N_24249,N_24726);
nor U26617 (N_26617,N_25058,N_25048);
or U26618 (N_26618,N_24846,N_24760);
nor U26619 (N_26619,N_24546,N_24121);
or U26620 (N_26620,N_24618,N_25166);
nand U26621 (N_26621,N_24056,N_24334);
nor U26622 (N_26622,N_25158,N_25076);
xor U26623 (N_26623,N_24322,N_24639);
xnor U26624 (N_26624,N_25187,N_24947);
nand U26625 (N_26625,N_25423,N_25399);
and U26626 (N_26626,N_25231,N_24274);
xor U26627 (N_26627,N_24309,N_25428);
nor U26628 (N_26628,N_24458,N_25233);
nor U26629 (N_26629,N_25349,N_24594);
or U26630 (N_26630,N_25095,N_24811);
xor U26631 (N_26631,N_25247,N_24873);
nand U26632 (N_26632,N_24662,N_24441);
nor U26633 (N_26633,N_24988,N_24614);
and U26634 (N_26634,N_25056,N_25078);
xor U26635 (N_26635,N_25194,N_25319);
xor U26636 (N_26636,N_24278,N_24136);
nor U26637 (N_26637,N_25250,N_24936);
or U26638 (N_26638,N_24185,N_25314);
or U26639 (N_26639,N_24918,N_24619);
nand U26640 (N_26640,N_25474,N_24305);
nand U26641 (N_26641,N_24131,N_24752);
xnor U26642 (N_26642,N_25296,N_25080);
xor U26643 (N_26643,N_25040,N_25070);
or U26644 (N_26644,N_25438,N_24368);
nand U26645 (N_26645,N_24814,N_24464);
nand U26646 (N_26646,N_24180,N_24320);
nor U26647 (N_26647,N_24646,N_24361);
xnor U26648 (N_26648,N_25316,N_25128);
or U26649 (N_26649,N_24253,N_24575);
xor U26650 (N_26650,N_24411,N_24881);
xnor U26651 (N_26651,N_25492,N_25403);
nand U26652 (N_26652,N_24333,N_24045);
and U26653 (N_26653,N_25176,N_24208);
nor U26654 (N_26654,N_25266,N_25234);
nor U26655 (N_26655,N_24433,N_24700);
nor U26656 (N_26656,N_24690,N_25260);
nor U26657 (N_26657,N_25378,N_25114);
nor U26658 (N_26658,N_24425,N_24679);
nor U26659 (N_26659,N_25389,N_24897);
and U26660 (N_26660,N_25002,N_24605);
xor U26661 (N_26661,N_24332,N_24949);
or U26662 (N_26662,N_24920,N_25054);
and U26663 (N_26663,N_24407,N_24162);
or U26664 (N_26664,N_24518,N_25289);
or U26665 (N_26665,N_25495,N_25410);
and U26666 (N_26666,N_24819,N_24537);
and U26667 (N_26667,N_25189,N_24915);
nand U26668 (N_26668,N_24228,N_25393);
or U26669 (N_26669,N_24930,N_24163);
and U26670 (N_26670,N_25418,N_24983);
or U26671 (N_26671,N_24008,N_25137);
xnor U26672 (N_26672,N_24497,N_25145);
and U26673 (N_26673,N_24473,N_24303);
or U26674 (N_26674,N_25357,N_24264);
nor U26675 (N_26675,N_25424,N_24083);
nor U26676 (N_26676,N_25412,N_24284);
nor U26677 (N_26677,N_24822,N_24896);
xor U26678 (N_26678,N_24591,N_24844);
or U26679 (N_26679,N_24261,N_25421);
or U26680 (N_26680,N_24076,N_24101);
nand U26681 (N_26681,N_24885,N_25431);
xor U26682 (N_26682,N_24535,N_24593);
or U26683 (N_26683,N_25335,N_24998);
and U26684 (N_26684,N_24047,N_24820);
xor U26685 (N_26685,N_24794,N_24529);
or U26686 (N_26686,N_24200,N_24796);
xor U26687 (N_26687,N_25213,N_24618);
and U26688 (N_26688,N_24208,N_24028);
xnor U26689 (N_26689,N_25453,N_25118);
xor U26690 (N_26690,N_25251,N_24826);
nor U26691 (N_26691,N_24237,N_24490);
or U26692 (N_26692,N_24216,N_24292);
and U26693 (N_26693,N_24479,N_25138);
or U26694 (N_26694,N_24113,N_25235);
xnor U26695 (N_26695,N_24549,N_25346);
and U26696 (N_26696,N_24320,N_24025);
xor U26697 (N_26697,N_25185,N_24577);
or U26698 (N_26698,N_24826,N_25364);
nand U26699 (N_26699,N_24986,N_24664);
or U26700 (N_26700,N_24846,N_24767);
xor U26701 (N_26701,N_24319,N_24116);
and U26702 (N_26702,N_24144,N_24250);
nand U26703 (N_26703,N_24978,N_25130);
and U26704 (N_26704,N_25427,N_24562);
or U26705 (N_26705,N_24425,N_25409);
or U26706 (N_26706,N_24390,N_24773);
nand U26707 (N_26707,N_24032,N_25282);
nand U26708 (N_26708,N_24735,N_24337);
xnor U26709 (N_26709,N_25063,N_24641);
xor U26710 (N_26710,N_25282,N_24802);
and U26711 (N_26711,N_25242,N_24872);
nor U26712 (N_26712,N_24485,N_24738);
nand U26713 (N_26713,N_24355,N_24052);
nor U26714 (N_26714,N_24953,N_24775);
nand U26715 (N_26715,N_24306,N_24590);
xnor U26716 (N_26716,N_24024,N_24381);
and U26717 (N_26717,N_24835,N_24902);
nor U26718 (N_26718,N_25167,N_24318);
or U26719 (N_26719,N_24688,N_25227);
xor U26720 (N_26720,N_25289,N_24883);
and U26721 (N_26721,N_24020,N_24189);
or U26722 (N_26722,N_25280,N_25238);
nor U26723 (N_26723,N_25192,N_24078);
nor U26724 (N_26724,N_24453,N_25150);
and U26725 (N_26725,N_24641,N_24279);
nand U26726 (N_26726,N_24689,N_24009);
and U26727 (N_26727,N_24517,N_25248);
nand U26728 (N_26728,N_25035,N_24201);
or U26729 (N_26729,N_24782,N_25034);
and U26730 (N_26730,N_24504,N_25204);
nor U26731 (N_26731,N_24429,N_24338);
nand U26732 (N_26732,N_24774,N_24255);
nor U26733 (N_26733,N_24182,N_24901);
or U26734 (N_26734,N_25343,N_24509);
and U26735 (N_26735,N_24615,N_24516);
or U26736 (N_26736,N_24177,N_24754);
or U26737 (N_26737,N_24815,N_24746);
nor U26738 (N_26738,N_25299,N_24194);
or U26739 (N_26739,N_25347,N_25001);
nor U26740 (N_26740,N_24767,N_24327);
or U26741 (N_26741,N_24799,N_24362);
nand U26742 (N_26742,N_24807,N_24993);
nor U26743 (N_26743,N_25489,N_24281);
nor U26744 (N_26744,N_24182,N_24663);
xor U26745 (N_26745,N_24866,N_24508);
or U26746 (N_26746,N_24419,N_25471);
or U26747 (N_26747,N_24927,N_24644);
and U26748 (N_26748,N_24148,N_24963);
nor U26749 (N_26749,N_24655,N_24590);
nand U26750 (N_26750,N_24321,N_25449);
nand U26751 (N_26751,N_25224,N_25022);
xor U26752 (N_26752,N_25010,N_25293);
nor U26753 (N_26753,N_24688,N_24139);
nand U26754 (N_26754,N_25131,N_25291);
xor U26755 (N_26755,N_24457,N_24690);
xnor U26756 (N_26756,N_24048,N_24487);
or U26757 (N_26757,N_24178,N_24903);
and U26758 (N_26758,N_25328,N_25299);
nand U26759 (N_26759,N_25457,N_24100);
or U26760 (N_26760,N_24282,N_24102);
nor U26761 (N_26761,N_24828,N_25053);
and U26762 (N_26762,N_24255,N_24409);
xnor U26763 (N_26763,N_24458,N_24997);
xor U26764 (N_26764,N_24238,N_24833);
nand U26765 (N_26765,N_25093,N_24022);
nand U26766 (N_26766,N_24768,N_24398);
and U26767 (N_26767,N_24789,N_25316);
and U26768 (N_26768,N_24034,N_25202);
nor U26769 (N_26769,N_24376,N_24969);
nor U26770 (N_26770,N_24290,N_24985);
nand U26771 (N_26771,N_25257,N_24575);
nand U26772 (N_26772,N_25002,N_24039);
nor U26773 (N_26773,N_24238,N_24145);
or U26774 (N_26774,N_24289,N_24992);
xor U26775 (N_26775,N_25250,N_24439);
nand U26776 (N_26776,N_24090,N_25168);
nand U26777 (N_26777,N_25309,N_25191);
and U26778 (N_26778,N_24457,N_24052);
or U26779 (N_26779,N_24559,N_25441);
or U26780 (N_26780,N_24114,N_25083);
or U26781 (N_26781,N_24828,N_25076);
nand U26782 (N_26782,N_25191,N_25375);
nor U26783 (N_26783,N_24656,N_24698);
and U26784 (N_26784,N_24804,N_25298);
xor U26785 (N_26785,N_24618,N_25427);
xor U26786 (N_26786,N_25413,N_25355);
nand U26787 (N_26787,N_24249,N_24800);
nor U26788 (N_26788,N_25122,N_24220);
or U26789 (N_26789,N_24167,N_24258);
nor U26790 (N_26790,N_25335,N_24313);
xor U26791 (N_26791,N_24202,N_24606);
nor U26792 (N_26792,N_25037,N_24626);
nand U26793 (N_26793,N_25455,N_25422);
or U26794 (N_26794,N_24256,N_24349);
nor U26795 (N_26795,N_24877,N_24841);
nor U26796 (N_26796,N_24159,N_24448);
xor U26797 (N_26797,N_25365,N_24347);
xnor U26798 (N_26798,N_24591,N_25473);
or U26799 (N_26799,N_25398,N_25336);
nor U26800 (N_26800,N_24657,N_24294);
or U26801 (N_26801,N_25033,N_24599);
or U26802 (N_26802,N_24348,N_24782);
and U26803 (N_26803,N_24247,N_25188);
or U26804 (N_26804,N_25227,N_24954);
nor U26805 (N_26805,N_24554,N_24459);
or U26806 (N_26806,N_24565,N_24276);
nand U26807 (N_26807,N_25143,N_24550);
xnor U26808 (N_26808,N_25088,N_24812);
xnor U26809 (N_26809,N_25122,N_24690);
xnor U26810 (N_26810,N_25081,N_24753);
or U26811 (N_26811,N_24418,N_25464);
or U26812 (N_26812,N_24181,N_24272);
xnor U26813 (N_26813,N_24609,N_24280);
and U26814 (N_26814,N_24641,N_24125);
or U26815 (N_26815,N_24573,N_24743);
xor U26816 (N_26816,N_24311,N_24134);
nor U26817 (N_26817,N_25082,N_24866);
nand U26818 (N_26818,N_24620,N_24989);
xor U26819 (N_26819,N_24284,N_24075);
nand U26820 (N_26820,N_24513,N_25041);
xnor U26821 (N_26821,N_24598,N_24072);
nand U26822 (N_26822,N_24210,N_25191);
and U26823 (N_26823,N_24321,N_25235);
xor U26824 (N_26824,N_25172,N_25468);
nor U26825 (N_26825,N_25060,N_25328);
nand U26826 (N_26826,N_24208,N_24852);
nor U26827 (N_26827,N_24449,N_24442);
nand U26828 (N_26828,N_24101,N_25188);
and U26829 (N_26829,N_25394,N_24764);
nor U26830 (N_26830,N_25371,N_25434);
nand U26831 (N_26831,N_24706,N_24375);
xnor U26832 (N_26832,N_24974,N_24698);
nand U26833 (N_26833,N_24305,N_25284);
or U26834 (N_26834,N_24290,N_25159);
or U26835 (N_26835,N_24891,N_25077);
nand U26836 (N_26836,N_24921,N_25297);
nor U26837 (N_26837,N_24040,N_25028);
or U26838 (N_26838,N_25432,N_25218);
nor U26839 (N_26839,N_24205,N_24839);
xnor U26840 (N_26840,N_25418,N_25371);
nand U26841 (N_26841,N_25154,N_25394);
nand U26842 (N_26842,N_24277,N_25398);
and U26843 (N_26843,N_24992,N_24765);
xnor U26844 (N_26844,N_24610,N_24932);
nor U26845 (N_26845,N_24598,N_24742);
xor U26846 (N_26846,N_24078,N_25286);
or U26847 (N_26847,N_24531,N_24846);
nand U26848 (N_26848,N_24061,N_24643);
nor U26849 (N_26849,N_25498,N_24763);
or U26850 (N_26850,N_25148,N_25407);
or U26851 (N_26851,N_24702,N_24228);
and U26852 (N_26852,N_24420,N_24895);
and U26853 (N_26853,N_24776,N_24520);
and U26854 (N_26854,N_24061,N_24580);
or U26855 (N_26855,N_25196,N_25251);
or U26856 (N_26856,N_24025,N_25339);
and U26857 (N_26857,N_24002,N_25238);
and U26858 (N_26858,N_24670,N_24545);
or U26859 (N_26859,N_25027,N_24114);
nor U26860 (N_26860,N_25047,N_24504);
and U26861 (N_26861,N_24007,N_24738);
nor U26862 (N_26862,N_25099,N_24962);
or U26863 (N_26863,N_24209,N_24418);
xnor U26864 (N_26864,N_24751,N_25448);
and U26865 (N_26865,N_24730,N_25378);
or U26866 (N_26866,N_24313,N_25381);
and U26867 (N_26867,N_25346,N_24468);
nor U26868 (N_26868,N_25312,N_24906);
or U26869 (N_26869,N_24029,N_24347);
or U26870 (N_26870,N_24837,N_25260);
nand U26871 (N_26871,N_24083,N_24622);
nand U26872 (N_26872,N_25422,N_24888);
nand U26873 (N_26873,N_24615,N_24249);
nor U26874 (N_26874,N_24801,N_25288);
and U26875 (N_26875,N_24702,N_25383);
or U26876 (N_26876,N_24617,N_24289);
or U26877 (N_26877,N_25383,N_24248);
and U26878 (N_26878,N_25497,N_25341);
nor U26879 (N_26879,N_24918,N_24481);
xnor U26880 (N_26880,N_24037,N_24460);
nand U26881 (N_26881,N_25329,N_24082);
nor U26882 (N_26882,N_24762,N_24558);
xor U26883 (N_26883,N_24334,N_24504);
or U26884 (N_26884,N_24559,N_25219);
nor U26885 (N_26885,N_25417,N_25154);
or U26886 (N_26886,N_24749,N_25343);
nor U26887 (N_26887,N_24499,N_24057);
nor U26888 (N_26888,N_24217,N_24164);
or U26889 (N_26889,N_24392,N_24347);
or U26890 (N_26890,N_24941,N_25330);
or U26891 (N_26891,N_24506,N_24417);
nand U26892 (N_26892,N_24016,N_24863);
xor U26893 (N_26893,N_25220,N_25437);
nand U26894 (N_26894,N_24724,N_25142);
nand U26895 (N_26895,N_24889,N_24052);
nand U26896 (N_26896,N_24226,N_24348);
and U26897 (N_26897,N_25471,N_24998);
and U26898 (N_26898,N_24560,N_25386);
and U26899 (N_26899,N_24438,N_24569);
or U26900 (N_26900,N_24417,N_24228);
or U26901 (N_26901,N_25432,N_24749);
and U26902 (N_26902,N_24433,N_24967);
or U26903 (N_26903,N_24516,N_25159);
nand U26904 (N_26904,N_24042,N_24631);
nand U26905 (N_26905,N_24665,N_24998);
nor U26906 (N_26906,N_25084,N_24196);
nand U26907 (N_26907,N_24638,N_25183);
and U26908 (N_26908,N_25426,N_24799);
nand U26909 (N_26909,N_25227,N_24323);
and U26910 (N_26910,N_24967,N_24200);
and U26911 (N_26911,N_24230,N_24428);
xor U26912 (N_26912,N_24589,N_25272);
or U26913 (N_26913,N_24057,N_25187);
xnor U26914 (N_26914,N_24653,N_25084);
or U26915 (N_26915,N_25493,N_24841);
nand U26916 (N_26916,N_24464,N_24726);
or U26917 (N_26917,N_25009,N_24016);
nand U26918 (N_26918,N_24303,N_25205);
or U26919 (N_26919,N_24622,N_24533);
nor U26920 (N_26920,N_24388,N_24783);
xnor U26921 (N_26921,N_24873,N_24806);
nand U26922 (N_26922,N_25383,N_25145);
and U26923 (N_26923,N_25405,N_25385);
and U26924 (N_26924,N_24043,N_25236);
or U26925 (N_26925,N_24823,N_24339);
or U26926 (N_26926,N_24203,N_25148);
and U26927 (N_26927,N_24944,N_24360);
or U26928 (N_26928,N_24962,N_24022);
nand U26929 (N_26929,N_25083,N_24849);
nand U26930 (N_26930,N_24890,N_24524);
or U26931 (N_26931,N_25339,N_24924);
xor U26932 (N_26932,N_24395,N_25177);
or U26933 (N_26933,N_24989,N_25325);
or U26934 (N_26934,N_25045,N_24473);
nand U26935 (N_26935,N_24526,N_25457);
xnor U26936 (N_26936,N_24327,N_24491);
and U26937 (N_26937,N_25283,N_25076);
xor U26938 (N_26938,N_24890,N_24899);
and U26939 (N_26939,N_24061,N_24680);
xor U26940 (N_26940,N_24255,N_24363);
xnor U26941 (N_26941,N_24766,N_25120);
or U26942 (N_26942,N_24895,N_24631);
or U26943 (N_26943,N_24344,N_25061);
and U26944 (N_26944,N_24330,N_25356);
xor U26945 (N_26945,N_25387,N_25276);
and U26946 (N_26946,N_24479,N_25275);
nand U26947 (N_26947,N_24744,N_25424);
or U26948 (N_26948,N_25447,N_24092);
xnor U26949 (N_26949,N_24481,N_24375);
xor U26950 (N_26950,N_24043,N_24640);
or U26951 (N_26951,N_24127,N_24085);
xnor U26952 (N_26952,N_24232,N_25041);
and U26953 (N_26953,N_25286,N_24261);
xor U26954 (N_26954,N_25160,N_24233);
or U26955 (N_26955,N_24537,N_24836);
or U26956 (N_26956,N_24311,N_25169);
nand U26957 (N_26957,N_24456,N_24204);
and U26958 (N_26958,N_24459,N_24692);
nor U26959 (N_26959,N_25038,N_24294);
or U26960 (N_26960,N_24745,N_24798);
or U26961 (N_26961,N_25353,N_24850);
and U26962 (N_26962,N_24786,N_25402);
nand U26963 (N_26963,N_24718,N_25403);
nor U26964 (N_26964,N_24831,N_25343);
or U26965 (N_26965,N_24390,N_25495);
and U26966 (N_26966,N_24442,N_24478);
nand U26967 (N_26967,N_25204,N_25276);
xnor U26968 (N_26968,N_24747,N_25290);
xnor U26969 (N_26969,N_24394,N_24986);
nand U26970 (N_26970,N_24080,N_24857);
or U26971 (N_26971,N_24827,N_24460);
xor U26972 (N_26972,N_24076,N_25306);
and U26973 (N_26973,N_24852,N_24478);
and U26974 (N_26974,N_24054,N_25042);
nand U26975 (N_26975,N_25080,N_24365);
and U26976 (N_26976,N_24668,N_25481);
or U26977 (N_26977,N_24444,N_24751);
and U26978 (N_26978,N_24149,N_24527);
nor U26979 (N_26979,N_24306,N_24061);
xnor U26980 (N_26980,N_24194,N_24489);
or U26981 (N_26981,N_25060,N_25238);
nand U26982 (N_26982,N_24871,N_25341);
xnor U26983 (N_26983,N_25254,N_24945);
nor U26984 (N_26984,N_24066,N_24116);
nor U26985 (N_26985,N_24523,N_24592);
nand U26986 (N_26986,N_24483,N_24752);
or U26987 (N_26987,N_24998,N_24966);
nor U26988 (N_26988,N_24761,N_24052);
nand U26989 (N_26989,N_24161,N_25192);
xnor U26990 (N_26990,N_25393,N_24068);
xor U26991 (N_26991,N_24933,N_24328);
or U26992 (N_26992,N_24139,N_24880);
nor U26993 (N_26993,N_24681,N_24469);
xnor U26994 (N_26994,N_24247,N_25235);
and U26995 (N_26995,N_24441,N_24336);
xor U26996 (N_26996,N_24378,N_25009);
or U26997 (N_26997,N_24846,N_24643);
xnor U26998 (N_26998,N_24263,N_24244);
and U26999 (N_26999,N_24503,N_25278);
and U27000 (N_27000,N_26194,N_26448);
and U27001 (N_27001,N_26556,N_25531);
xor U27002 (N_27002,N_26784,N_25833);
and U27003 (N_27003,N_26352,N_26693);
and U27004 (N_27004,N_25637,N_26546);
nor U27005 (N_27005,N_26700,N_26409);
nand U27006 (N_27006,N_25764,N_26699);
nand U27007 (N_27007,N_25723,N_26379);
nand U27008 (N_27008,N_26196,N_25505);
xor U27009 (N_27009,N_25921,N_25856);
or U27010 (N_27010,N_26834,N_26513);
or U27011 (N_27011,N_25546,N_26113);
and U27012 (N_27012,N_26524,N_26628);
or U27013 (N_27013,N_26798,N_26708);
nor U27014 (N_27014,N_26161,N_25683);
or U27015 (N_27015,N_26520,N_25885);
nand U27016 (N_27016,N_26036,N_26721);
or U27017 (N_27017,N_25698,N_26820);
xnor U27018 (N_27018,N_25646,N_25613);
and U27019 (N_27019,N_26990,N_25570);
nand U27020 (N_27020,N_26559,N_25584);
or U27021 (N_27021,N_25781,N_26906);
nand U27022 (N_27022,N_25557,N_26537);
xor U27023 (N_27023,N_25862,N_25797);
or U27024 (N_27024,N_26970,N_25636);
nand U27025 (N_27025,N_26475,N_26376);
nor U27026 (N_27026,N_26143,N_26211);
and U27027 (N_27027,N_26770,N_26712);
nand U27028 (N_27028,N_26565,N_26627);
and U27029 (N_27029,N_25894,N_26213);
and U27030 (N_27030,N_25765,N_26681);
nor U27031 (N_27031,N_26014,N_25896);
nor U27032 (N_27032,N_25594,N_26724);
or U27033 (N_27033,N_26722,N_25848);
nand U27034 (N_27034,N_26315,N_26394);
and U27035 (N_27035,N_26363,N_26823);
and U27036 (N_27036,N_26868,N_26980);
nor U27037 (N_27037,N_26393,N_26821);
nor U27038 (N_27038,N_26054,N_25898);
xor U27039 (N_27039,N_26165,N_26610);
or U27040 (N_27040,N_25927,N_25759);
xor U27041 (N_27041,N_26479,N_26072);
nand U27042 (N_27042,N_26461,N_26971);
nand U27043 (N_27043,N_26824,N_26037);
xor U27044 (N_27044,N_26144,N_25631);
nand U27045 (N_27045,N_26274,N_26058);
nor U27046 (N_27046,N_26180,N_26382);
xnor U27047 (N_27047,N_26195,N_25974);
nand U27048 (N_27048,N_26728,N_26341);
or U27049 (N_27049,N_26273,N_26501);
nor U27050 (N_27050,N_26843,N_26313);
and U27051 (N_27051,N_25814,N_26988);
and U27052 (N_27052,N_26365,N_26127);
xor U27053 (N_27053,N_26793,N_26595);
nand U27054 (N_27054,N_26052,N_26119);
nor U27055 (N_27055,N_26239,N_26573);
or U27056 (N_27056,N_25605,N_26137);
and U27057 (N_27057,N_25753,N_25804);
or U27058 (N_27058,N_25558,N_26814);
or U27059 (N_27059,N_26328,N_26954);
or U27060 (N_27060,N_26308,N_26743);
xor U27061 (N_27061,N_26995,N_26011);
nor U27062 (N_27062,N_26283,N_25917);
nor U27063 (N_27063,N_26762,N_26282);
nor U27064 (N_27064,N_26992,N_26640);
or U27065 (N_27065,N_26083,N_26404);
or U27066 (N_27066,N_26355,N_25782);
xnor U27067 (N_27067,N_26185,N_25922);
or U27068 (N_27068,N_26764,N_25773);
nor U27069 (N_27069,N_25695,N_26181);
nor U27070 (N_27070,N_26476,N_25535);
nand U27071 (N_27071,N_26593,N_26487);
nand U27072 (N_27072,N_26269,N_25763);
and U27073 (N_27073,N_25831,N_26751);
nor U27074 (N_27074,N_25624,N_26013);
xnor U27075 (N_27075,N_26733,N_26601);
or U27076 (N_27076,N_26465,N_26342);
nor U27077 (N_27077,N_26103,N_26400);
or U27078 (N_27078,N_26430,N_26198);
or U27079 (N_27079,N_25714,N_26803);
xnor U27080 (N_27080,N_26596,N_26038);
nor U27081 (N_27081,N_25711,N_26248);
nor U27082 (N_27082,N_25815,N_25670);
nand U27083 (N_27083,N_26735,N_26934);
nand U27084 (N_27084,N_25778,N_26318);
nand U27085 (N_27085,N_26380,N_26809);
nand U27086 (N_27086,N_26490,N_26249);
and U27087 (N_27087,N_25902,N_26200);
xor U27088 (N_27088,N_26958,N_26081);
xnor U27089 (N_27089,N_26870,N_26648);
or U27090 (N_27090,N_26622,N_26949);
nor U27091 (N_27091,N_26514,N_26133);
nor U27092 (N_27092,N_25871,N_25843);
nand U27093 (N_27093,N_26689,N_26398);
xnor U27094 (N_27094,N_25543,N_26129);
xnor U27095 (N_27095,N_26043,N_25602);
nand U27096 (N_27096,N_25859,N_26940);
and U27097 (N_27097,N_26335,N_26157);
or U27098 (N_27098,N_26528,N_26948);
nor U27099 (N_27099,N_25530,N_26085);
xor U27100 (N_27100,N_25671,N_26900);
xnor U27101 (N_27101,N_25733,N_25527);
nor U27102 (N_27102,N_26962,N_26794);
and U27103 (N_27103,N_26406,N_25668);
nand U27104 (N_27104,N_25573,N_25736);
nand U27105 (N_27105,N_26719,N_25587);
and U27106 (N_27106,N_26874,N_25734);
nand U27107 (N_27107,N_25571,N_26332);
and U27108 (N_27108,N_26656,N_26295);
and U27109 (N_27109,N_25682,N_26401);
or U27110 (N_27110,N_25621,N_26303);
and U27111 (N_27111,N_25761,N_26366);
and U27112 (N_27112,N_25882,N_25891);
nand U27113 (N_27113,N_26463,N_26117);
and U27114 (N_27114,N_26496,N_26999);
nand U27115 (N_27115,N_26378,N_26894);
and U27116 (N_27116,N_26484,N_26760);
or U27117 (N_27117,N_26592,N_25887);
or U27118 (N_27118,N_26678,N_26732);
nand U27119 (N_27119,N_25817,N_25540);
and U27120 (N_27120,N_25715,N_26278);
nand U27121 (N_27121,N_26444,N_25672);
and U27122 (N_27122,N_26319,N_26073);
nor U27123 (N_27123,N_26292,N_26539);
and U27124 (N_27124,N_26612,N_26942);
or U27125 (N_27125,N_25823,N_26633);
nand U27126 (N_27126,N_25906,N_25800);
nor U27127 (N_27127,N_26788,N_25514);
nand U27128 (N_27128,N_26275,N_25533);
or U27129 (N_27129,N_26680,N_25549);
or U27130 (N_27130,N_25520,N_26474);
or U27131 (N_27131,N_26581,N_26545);
and U27132 (N_27132,N_26951,N_26397);
nand U27133 (N_27133,N_25526,N_26527);
and U27134 (N_27134,N_26854,N_25913);
and U27135 (N_27135,N_26092,N_26445);
nor U27136 (N_27136,N_26383,N_26881);
nand U27137 (N_27137,N_25623,N_25586);
or U27138 (N_27138,N_26647,N_26070);
nor U27139 (N_27139,N_25910,N_26405);
or U27140 (N_27140,N_26176,N_26774);
xnor U27141 (N_27141,N_26945,N_26585);
xnor U27142 (N_27142,N_26460,N_26550);
or U27143 (N_27143,N_25926,N_26336);
or U27144 (N_27144,N_26572,N_26158);
nand U27145 (N_27145,N_25740,N_25809);
nand U27146 (N_27146,N_26635,N_26146);
and U27147 (N_27147,N_26175,N_26168);
nor U27148 (N_27148,N_26234,N_26558);
nor U27149 (N_27149,N_25567,N_25725);
or U27150 (N_27150,N_26525,N_26367);
and U27151 (N_27151,N_26488,N_26502);
and U27152 (N_27152,N_26936,N_26755);
xor U27153 (N_27153,N_25941,N_26718);
xnor U27154 (N_27154,N_26626,N_26756);
nand U27155 (N_27155,N_26683,N_26028);
or U27156 (N_27156,N_26391,N_26048);
or U27157 (N_27157,N_26049,N_26167);
nor U27158 (N_27158,N_26829,N_26704);
or U27159 (N_27159,N_25643,N_26686);
or U27160 (N_27160,N_26260,N_26543);
or U27161 (N_27161,N_26782,N_26588);
nor U27162 (N_27162,N_26416,N_26511);
nor U27163 (N_27163,N_26613,N_26270);
nand U27164 (N_27164,N_26191,N_26608);
xnor U27165 (N_27165,N_26862,N_26122);
or U27166 (N_27166,N_26257,N_26657);
nand U27167 (N_27167,N_26171,N_26017);
and U27168 (N_27168,N_25966,N_26547);
nor U27169 (N_27169,N_26436,N_26553);
nand U27170 (N_27170,N_26884,N_26982);
xor U27171 (N_27171,N_26517,N_26716);
xor U27172 (N_27172,N_26026,N_26510);
and U27173 (N_27173,N_26482,N_25658);
nand U27174 (N_27174,N_26012,N_25789);
and U27175 (N_27175,N_26984,N_26882);
nor U27176 (N_27176,N_25529,N_26715);
or U27177 (N_27177,N_26675,N_25977);
and U27178 (N_27178,N_25750,N_26039);
and U27179 (N_27179,N_26023,N_25961);
nor U27180 (N_27180,N_26620,N_26123);
xnor U27181 (N_27181,N_26757,N_25840);
nor U27182 (N_27182,N_26768,N_26458);
and U27183 (N_27183,N_25730,N_26230);
nor U27184 (N_27184,N_25786,N_25615);
nand U27185 (N_27185,N_25609,N_25504);
or U27186 (N_27186,N_26529,N_25881);
xnor U27187 (N_27187,N_26251,N_26914);
xnor U27188 (N_27188,N_26826,N_26206);
xnor U27189 (N_27189,N_26896,N_26139);
nand U27190 (N_27190,N_26932,N_26493);
nand U27191 (N_27191,N_25721,N_25618);
xor U27192 (N_27192,N_26433,N_26202);
nor U27193 (N_27193,N_25738,N_26041);
nand U27194 (N_27194,N_26805,N_26521);
nand U27195 (N_27195,N_25627,N_25667);
xor U27196 (N_27196,N_26673,N_25818);
or U27197 (N_27197,N_26837,N_26228);
xor U27198 (N_27198,N_26399,N_25656);
nor U27199 (N_27199,N_25932,N_26421);
or U27200 (N_27200,N_26053,N_26464);
nor U27201 (N_27201,N_26388,N_26497);
or U27202 (N_27202,N_26816,N_26812);
nor U27203 (N_27203,N_26746,N_26979);
or U27204 (N_27204,N_26802,N_26918);
and U27205 (N_27205,N_26364,N_26549);
and U27206 (N_27206,N_26682,N_25691);
or U27207 (N_27207,N_26531,N_25710);
or U27208 (N_27208,N_26138,N_25564);
nor U27209 (N_27209,N_25767,N_26005);
and U27210 (N_27210,N_26575,N_26957);
and U27211 (N_27211,N_26907,N_26451);
xnor U27212 (N_27212,N_25747,N_26483);
and U27213 (N_27213,N_25869,N_25552);
xnor U27214 (N_27214,N_26076,N_26109);
and U27215 (N_27215,N_26231,N_25653);
nor U27216 (N_27216,N_26205,N_25641);
or U27217 (N_27217,N_26418,N_25807);
and U27218 (N_27218,N_26492,N_25728);
xnor U27219 (N_27219,N_26172,N_26062);
nor U27220 (N_27220,N_26885,N_25697);
nor U27221 (N_27221,N_26877,N_26773);
nand U27222 (N_27222,N_26557,N_26734);
nor U27223 (N_27223,N_25665,N_26845);
nor U27224 (N_27224,N_25518,N_25752);
xnor U27225 (N_27225,N_26093,N_25939);
nand U27226 (N_27226,N_26661,N_26199);
xnor U27227 (N_27227,N_25751,N_25745);
nor U27228 (N_27228,N_26901,N_26124);
and U27229 (N_27229,N_26969,N_26216);
or U27230 (N_27230,N_26035,N_25998);
or U27231 (N_27231,N_25940,N_26665);
or U27232 (N_27232,N_26259,N_26238);
nand U27233 (N_27233,N_26791,N_26761);
or U27234 (N_27234,N_25942,N_26783);
or U27235 (N_27235,N_26432,N_26452);
or U27236 (N_27236,N_26658,N_26311);
or U27237 (N_27237,N_26197,N_25937);
xnor U27238 (N_27238,N_25666,N_26915);
or U27239 (N_27239,N_26115,N_26615);
or U27240 (N_27240,N_25548,N_25598);
and U27241 (N_27241,N_26147,N_25978);
or U27242 (N_27242,N_25681,N_26417);
nor U27243 (N_27243,N_25562,N_26296);
nor U27244 (N_27244,N_25979,N_26107);
nor U27245 (N_27245,N_25991,N_26844);
and U27246 (N_27246,N_26747,N_25655);
xor U27247 (N_27247,N_26830,N_26214);
or U27248 (N_27248,N_26883,N_26852);
nand U27249 (N_27249,N_26672,N_25701);
or U27250 (N_27250,N_25805,N_26603);
nor U27251 (N_27251,N_25542,N_25669);
nand U27252 (N_27252,N_25886,N_26136);
xor U27253 (N_27253,N_25509,N_26201);
nand U27254 (N_27254,N_26368,N_26937);
xor U27255 (N_27255,N_26173,N_26560);
nor U27256 (N_27256,N_25645,N_26343);
nor U27257 (N_27257,N_25517,N_25685);
nor U27258 (N_27258,N_26655,N_26245);
nand U27259 (N_27259,N_26584,N_26390);
nor U27260 (N_27260,N_25957,N_26277);
nand U27261 (N_27261,N_25774,N_25739);
nand U27262 (N_27262,N_25617,N_25965);
and U27263 (N_27263,N_26972,N_26402);
nor U27264 (N_27264,N_26334,N_25718);
and U27265 (N_27265,N_26838,N_25565);
and U27266 (N_27266,N_26604,N_26486);
and U27267 (N_27267,N_26811,N_26674);
nand U27268 (N_27268,N_25729,N_26098);
xnor U27269 (N_27269,N_26912,N_25828);
nor U27270 (N_27270,N_26424,N_26462);
and U27271 (N_27271,N_26861,N_25703);
xor U27272 (N_27272,N_25716,N_26153);
xnor U27273 (N_27273,N_26684,N_26253);
nand U27274 (N_27274,N_25851,N_26044);
or U27275 (N_27275,N_25844,N_25888);
or U27276 (N_27276,N_26059,N_26410);
nor U27277 (N_27277,N_26019,N_26140);
nor U27278 (N_27278,N_26387,N_25625);
nand U27279 (N_27279,N_26569,N_26643);
and U27280 (N_27280,N_25560,N_26748);
nor U27281 (N_27281,N_26207,N_25528);
nor U27282 (N_27282,N_25663,N_26818);
xnor U27283 (N_27283,N_26159,N_25596);
nand U27284 (N_27284,N_25949,N_25630);
and U27285 (N_27285,N_25976,N_26047);
or U27286 (N_27286,N_25591,N_25892);
nor U27287 (N_27287,N_26375,N_26179);
nand U27288 (N_27288,N_26320,N_26022);
nand U27289 (N_27289,N_26340,N_26395);
and U27290 (N_27290,N_25792,N_25770);
nor U27291 (N_27291,N_26653,N_25821);
nor U27292 (N_27292,N_25628,N_25950);
xor U27293 (N_27293,N_25982,N_26056);
or U27294 (N_27294,N_25603,N_26169);
xor U27295 (N_27295,N_25948,N_26864);
or U27296 (N_27296,N_25633,N_26272);
or U27297 (N_27297,N_25787,N_26287);
and U27298 (N_27298,N_26926,N_26538);
nand U27299 (N_27299,N_26892,N_26920);
or U27300 (N_27300,N_26662,N_26533);
xor U27301 (N_27301,N_26536,N_26489);
nand U27302 (N_27302,N_26815,N_26166);
nand U27303 (N_27303,N_26899,N_26561);
nand U27304 (N_27304,N_26532,N_26714);
nor U27305 (N_27305,N_26978,N_25766);
or U27306 (N_27306,N_26411,N_26294);
nor U27307 (N_27307,N_26804,N_25769);
and U27308 (N_27308,N_25538,N_26254);
nand U27309 (N_27309,N_25574,N_26566);
or U27310 (N_27310,N_26099,N_26644);
nor U27311 (N_27311,N_25709,N_26905);
xor U27312 (N_27312,N_25554,N_26247);
and U27313 (N_27313,N_25849,N_26863);
or U27314 (N_27314,N_25513,N_26333);
nand U27315 (N_27315,N_25507,N_26706);
nor U27316 (N_27316,N_25614,N_25999);
nor U27317 (N_27317,N_26177,N_26141);
xnor U27318 (N_27318,N_26255,N_26021);
xnor U27319 (N_27319,N_26930,N_26720);
and U27320 (N_27320,N_25880,N_25600);
xnor U27321 (N_27321,N_25962,N_26504);
nor U27322 (N_27322,N_26232,N_25912);
nand U27323 (N_27323,N_26779,N_25577);
xnor U27324 (N_27324,N_25692,N_26729);
xor U27325 (N_27325,N_25502,N_26535);
nor U27326 (N_27326,N_26987,N_26841);
nor U27327 (N_27327,N_26944,N_26221);
nor U27328 (N_27328,N_26638,N_26745);
xnor U27329 (N_27329,N_25983,N_25972);
and U27330 (N_27330,N_25649,N_26636);
xnor U27331 (N_27331,N_25784,N_26346);
and U27332 (N_27332,N_25512,N_26797);
or U27333 (N_27333,N_26423,N_26965);
nand U27334 (N_27334,N_26562,N_26668);
or U27335 (N_27335,N_25951,N_25620);
nor U27336 (N_27336,N_26090,N_25662);
and U27337 (N_27337,N_26742,N_26664);
or U27338 (N_27338,N_26792,N_26835);
nand U27339 (N_27339,N_26850,N_25675);
or U27340 (N_27340,N_26289,N_25744);
nor U27341 (N_27341,N_25510,N_26904);
xnor U27342 (N_27342,N_25901,N_26454);
nor U27343 (N_27343,N_25973,N_25741);
xor U27344 (N_27344,N_26625,N_25676);
xnor U27345 (N_27345,N_26555,N_25595);
xor U27346 (N_27346,N_26121,N_26671);
and U27347 (N_27347,N_25634,N_25679);
xnor U27348 (N_27348,N_25712,N_26435);
and U27349 (N_27349,N_26084,N_26025);
nor U27350 (N_27350,N_25879,N_26749);
nor U27351 (N_27351,N_26220,N_26571);
nand U27352 (N_27352,N_25846,N_26691);
nand U27353 (N_27353,N_26500,N_26800);
nor U27354 (N_27354,N_26750,N_25678);
xor U27355 (N_27355,N_25827,N_26607);
and U27356 (N_27356,N_25619,N_25775);
nand U27357 (N_27357,N_26306,N_26941);
nor U27358 (N_27358,N_26246,N_26583);
and U27359 (N_27359,N_26078,N_26326);
nor U27360 (N_27360,N_26512,N_26590);
and U27361 (N_27361,N_25900,N_26676);
nor U27362 (N_27362,N_26789,N_25674);
xnor U27363 (N_27363,N_25858,N_26212);
xnor U27364 (N_27364,N_26917,N_26473);
nand U27365 (N_27365,N_26217,N_25987);
nand U27366 (N_27366,N_26096,N_26624);
nor U27367 (N_27367,N_25820,N_25593);
and U27368 (N_27368,N_26692,N_25608);
and U27369 (N_27369,N_26744,N_26976);
nor U27370 (N_27370,N_26086,N_26519);
nand U27371 (N_27371,N_26597,N_25632);
or U27372 (N_27372,N_26679,N_26996);
and U27373 (N_27373,N_26591,N_26243);
nor U27374 (N_27374,N_26040,N_25839);
or U27375 (N_27375,N_25606,N_26068);
or U27376 (N_27376,N_25661,N_26650);
and U27377 (N_27377,N_26856,N_26032);
or U27378 (N_27378,N_26867,N_26785);
or U27379 (N_27379,N_25995,N_25816);
and U27380 (N_27380,N_26840,N_26737);
or U27381 (N_27381,N_26865,N_26118);
and U27382 (N_27382,N_25933,N_26652);
and U27383 (N_27383,N_26235,N_25545);
nor U27384 (N_27384,N_26271,N_25929);
or U27385 (N_27385,N_25550,N_26414);
nor U27386 (N_27386,N_26403,N_26858);
nand U27387 (N_27387,N_26266,N_25523);
or U27388 (N_27388,N_26564,N_26778);
nor U27389 (N_27389,N_25762,N_25746);
and U27390 (N_27390,N_26786,N_25810);
nor U27391 (N_27391,N_26101,N_26097);
xnor U27392 (N_27392,N_26134,N_26832);
xnor U27393 (N_27393,N_26067,N_26468);
and U27394 (N_27394,N_26876,N_25980);
and U27395 (N_27395,N_25755,N_25657);
and U27396 (N_27396,N_26357,N_26002);
nor U27397 (N_27397,N_26589,N_25503);
nand U27398 (N_27398,N_25616,N_26983);
nand U27399 (N_27399,N_26425,N_26034);
nand U27400 (N_27400,N_26776,N_26050);
or U27401 (N_27401,N_25777,N_26188);
and U27402 (N_27402,N_26349,N_25639);
or U27403 (N_27403,N_26594,N_26371);
or U27404 (N_27404,N_25757,N_26413);
xor U27405 (N_27405,N_26522,N_26408);
or U27406 (N_27406,N_26518,N_26801);
and U27407 (N_27407,N_26509,N_25825);
nand U27408 (N_27408,N_25813,N_25754);
or U27409 (N_27409,N_26766,N_25583);
nand U27410 (N_27410,N_26089,N_25724);
and U27411 (N_27411,N_26112,N_25790);
and U27412 (N_27412,N_25988,N_25651);
xor U27413 (N_27413,N_26356,N_26300);
nor U27414 (N_27414,N_26694,N_25986);
and U27415 (N_27415,N_25705,N_25934);
xor U27416 (N_27416,N_25826,N_26007);
nand U27417 (N_27417,N_25629,N_25802);
xnor U27418 (N_27418,N_26066,N_26911);
and U27419 (N_27419,N_25946,N_26966);
and U27420 (N_27420,N_26579,N_26152);
or U27421 (N_27421,N_26069,N_26739);
xnor U27422 (N_27422,N_26888,N_25704);
xnor U27423 (N_27423,N_26329,N_25829);
and U27424 (N_27424,N_26859,N_26304);
nor U27425 (N_27425,N_26790,N_26775);
nand U27426 (N_27426,N_25909,N_25516);
nor U27427 (N_27427,N_26961,N_26100);
xor U27428 (N_27428,N_26377,N_26051);
nand U27429 (N_27429,N_26362,N_26227);
nand U27430 (N_27430,N_26384,N_25935);
or U27431 (N_27431,N_25954,N_26323);
or U27432 (N_27432,N_25911,N_26351);
and U27433 (N_27433,N_25664,N_26499);
xnor U27434 (N_27434,N_26752,N_26369);
nand U27435 (N_27435,N_25893,N_26781);
nand U27436 (N_27436,N_26860,N_25794);
and U27437 (N_27437,N_26046,N_26237);
nand U27438 (N_27438,N_26836,N_26736);
and U27439 (N_27439,N_26088,N_26286);
nand U27440 (N_27440,N_26981,N_25556);
nor U27441 (N_27441,N_26160,N_26309);
nand U27442 (N_27442,N_26889,N_25575);
or U27443 (N_27443,N_26710,N_26412);
nor U27444 (N_27444,N_26485,N_26225);
nor U27445 (N_27445,N_26471,N_26061);
xnor U27446 (N_27446,N_26419,N_25737);
and U27447 (N_27447,N_25680,N_25970);
nand U27448 (N_27448,N_26030,N_26869);
nand U27449 (N_27449,N_26960,N_26015);
or U27450 (N_27450,N_26910,N_25956);
nor U27451 (N_27451,N_25920,N_26447);
or U27452 (N_27452,N_25650,N_26909);
or U27453 (N_27453,N_25588,N_26924);
or U27454 (N_27454,N_26000,N_26261);
xor U27455 (N_27455,N_26064,N_26925);
and U27456 (N_27456,N_25511,N_25832);
xor U27457 (N_27457,N_26074,N_25532);
or U27458 (N_27458,N_26244,N_26219);
xnor U27459 (N_27459,N_25819,N_26297);
or U27460 (N_27460,N_25931,N_26893);
and U27461 (N_27461,N_26921,N_25553);
xnor U27462 (N_27462,N_26947,N_26939);
or U27463 (N_27463,N_26114,N_26938);
or U27464 (N_27464,N_26392,N_26163);
nand U27465 (N_27465,N_25963,N_26605);
nand U27466 (N_27466,N_26466,N_26902);
nand U27467 (N_27467,N_26717,N_26386);
and U27468 (N_27468,N_26370,N_26927);
or U27469 (N_27469,N_25611,N_26148);
nor U27470 (N_27470,N_25551,N_25857);
and U27471 (N_27471,N_25967,N_26293);
nor U27472 (N_27472,N_25559,N_26623);
nor U27473 (N_27473,N_26544,N_26631);
xnor U27474 (N_27474,N_25563,N_26279);
nand U27475 (N_27475,N_26629,N_26102);
and U27476 (N_27476,N_25544,N_26440);
nand U27477 (N_27477,N_26967,N_26077);
nor U27478 (N_27478,N_26372,N_25884);
nor U27479 (N_27479,N_26890,N_25521);
xnor U27480 (N_27480,N_25780,N_26407);
nand U27481 (N_27481,N_26457,N_25776);
nand U27482 (N_27482,N_25537,N_26851);
nor U27483 (N_27483,N_26991,N_26731);
nand U27484 (N_27484,N_26285,N_25694);
and U27485 (N_27485,N_26095,N_26866);
nor U27486 (N_27486,N_25944,N_26057);
or U27487 (N_27487,N_26651,N_26873);
nor U27488 (N_27488,N_25768,N_26331);
nor U27489 (N_27489,N_26598,N_26725);
and U27490 (N_27490,N_25785,N_26956);
and U27491 (N_27491,N_25735,N_26317);
nor U27492 (N_27492,N_26663,N_25799);
or U27493 (N_27493,N_26265,N_26848);
or U27494 (N_27494,N_26810,N_25506);
xor U27495 (N_27495,N_25500,N_26060);
nor U27496 (N_27496,N_25717,N_26325);
and U27497 (N_27497,N_25722,N_25660);
nand U27498 (N_27498,N_26688,N_26759);
or U27499 (N_27499,N_26645,N_26094);
nand U27500 (N_27500,N_26616,N_25938);
or U27501 (N_27501,N_26503,N_26577);
nand U27502 (N_27502,N_26570,N_26204);
or U27503 (N_27503,N_25748,N_26470);
and U27504 (N_27504,N_26817,N_26974);
xor U27505 (N_27505,N_25873,N_26027);
nor U27506 (N_27506,N_25865,N_26726);
nand U27507 (N_27507,N_26374,N_25989);
nand U27508 (N_27508,N_26441,N_25968);
xnor U27509 (N_27509,N_26156,N_25597);
nor U27510 (N_27510,N_25731,N_25836);
nand U27511 (N_27511,N_26576,N_25795);
or U27512 (N_27512,N_25803,N_25860);
nor U27513 (N_27513,N_26310,N_25515);
and U27514 (N_27514,N_26505,N_26469);
nor U27515 (N_27515,N_26437,N_26913);
nor U27516 (N_27516,N_26822,N_25578);
and U27517 (N_27517,N_26018,N_26373);
nand U27518 (N_27518,N_25953,N_26931);
nor U27519 (N_27519,N_25868,N_25812);
or U27520 (N_27520,N_26703,N_26337);
nand U27521 (N_27521,N_26130,N_25852);
or U27522 (N_27522,N_26164,N_25847);
xnor U27523 (N_27523,N_25654,N_25622);
and U27524 (N_27524,N_25904,N_26291);
and U27525 (N_27525,N_26641,N_26609);
and U27526 (N_27526,N_26080,N_25522);
and U27527 (N_27527,N_26314,N_26258);
xor U27528 (N_27528,N_26878,N_26606);
nand U27529 (N_27529,N_25756,N_26897);
or U27530 (N_27530,N_26660,N_25589);
nand U27531 (N_27531,N_26630,N_26828);
nor U27532 (N_27532,N_26857,N_26189);
and U27533 (N_27533,N_25635,N_25585);
xor U27534 (N_27534,N_25601,N_26250);
or U27535 (N_27535,N_25877,N_25796);
xnor U27536 (N_27536,N_26456,N_26438);
xnor U27537 (N_27537,N_26494,N_26186);
xor U27538 (N_27538,N_25878,N_26415);
and U27539 (N_27539,N_26455,N_25874);
xnor U27540 (N_27540,N_26919,N_26029);
or U27541 (N_27541,N_26955,N_25626);
or U27542 (N_27542,N_26707,N_26690);
nor U27543 (N_27543,N_26075,N_25875);
or U27544 (N_27544,N_26031,N_26498);
nor U27545 (N_27545,N_26055,N_26959);
xor U27546 (N_27546,N_25599,N_25534);
and U27547 (N_27547,N_26290,N_26687);
nor U27548 (N_27548,N_26478,N_26696);
xnor U27549 (N_27549,N_25719,N_25708);
nor U27550 (N_27550,N_26827,N_25647);
and U27551 (N_27551,N_26541,N_26145);
nand U27552 (N_27552,N_26358,N_25908);
nor U27553 (N_27553,N_25899,N_26359);
and U27554 (N_27554,N_26256,N_26701);
or U27555 (N_27555,N_26322,N_25822);
or U27556 (N_27556,N_26943,N_26554);
and U27557 (N_27557,N_26923,N_26670);
or U27558 (N_27558,N_26241,N_26666);
nand U27559 (N_27559,N_25808,N_25555);
and U27560 (N_27560,N_25811,N_26450);
and U27561 (N_27561,N_26299,N_26280);
or U27562 (N_27562,N_26895,N_25569);
nand U27563 (N_27563,N_26420,N_26695);
nand U27564 (N_27564,N_26229,N_26952);
nand U27565 (N_27565,N_25806,N_26713);
and U27566 (N_27566,N_26151,N_26087);
nand U27567 (N_27567,N_25975,N_25590);
nor U27568 (N_27568,N_26302,N_25801);
or U27569 (N_27569,N_25866,N_26020);
nand U27570 (N_27570,N_26042,N_25687);
or U27571 (N_27571,N_26993,N_26467);
and U27572 (N_27572,N_26621,N_26347);
xnor U27573 (N_27573,N_25861,N_25580);
and U27574 (N_27574,N_26209,N_26396);
nor U27575 (N_27575,N_26677,N_25889);
nor U27576 (N_27576,N_25783,N_25742);
and U27577 (N_27577,N_25581,N_26348);
or U27578 (N_27578,N_26552,N_26480);
and U27579 (N_27579,N_26758,N_26973);
and U27580 (N_27580,N_25855,N_26389);
xnor U27581 (N_27581,N_26116,N_26008);
nand U27582 (N_27582,N_26580,N_26298);
or U27583 (N_27583,N_26003,N_26472);
and U27584 (N_27584,N_26284,N_26875);
xor U27585 (N_27585,N_25981,N_26697);
nand U27586 (N_27586,N_25923,N_26618);
or U27587 (N_27587,N_26602,N_26542);
nand U27588 (N_27588,N_26642,N_25928);
nand U27589 (N_27589,N_26667,N_25890);
nor U27590 (N_27590,N_25732,N_26600);
nand U27591 (N_27591,N_26507,N_26033);
nand U27592 (N_27592,N_26659,N_25688);
xor U27593 (N_27593,N_26010,N_26654);
or U27594 (N_27594,N_26551,N_25876);
or U27595 (N_27595,N_26459,N_25870);
nor U27596 (N_27596,N_26842,N_26772);
nor U27597 (N_27597,N_26004,N_25568);
and U27598 (N_27598,N_26639,N_26428);
or U27599 (N_27599,N_26508,N_26024);
and U27600 (N_27600,N_25539,N_26685);
and U27601 (N_27601,N_26617,N_26174);
nor U27602 (N_27602,N_26730,N_26126);
and U27603 (N_27603,N_26345,N_26929);
nor U27604 (N_27604,N_25992,N_26252);
xnor U27605 (N_27605,N_26045,N_26833);
nor U27606 (N_27606,N_25536,N_26530);
nand U27607 (N_27607,N_25690,N_26305);
nand U27608 (N_27608,N_25713,N_25947);
nand U27609 (N_27609,N_26727,N_26193);
nor U27610 (N_27610,N_26891,N_26105);
nand U27611 (N_27611,N_26215,N_26307);
nand U27612 (N_27612,N_25955,N_26582);
xnor U27613 (N_27613,N_25758,N_26825);
xnor U27614 (N_27614,N_25945,N_26908);
or U27615 (N_27615,N_26698,N_25541);
or U27616 (N_27616,N_26935,N_25959);
and U27617 (N_27617,N_25689,N_25749);
nor U27618 (N_27618,N_26120,N_26953);
nor U27619 (N_27619,N_26106,N_26001);
xor U27620 (N_27620,N_25872,N_25915);
nor U27621 (N_27621,N_25592,N_26846);
or U27622 (N_27622,N_25960,N_26446);
nand U27623 (N_27623,N_26236,N_26267);
nand U27624 (N_27624,N_25642,N_26807);
and U27625 (N_27625,N_25579,N_26632);
nor U27626 (N_27626,N_26016,N_25699);
or U27627 (N_27627,N_25867,N_25519);
nand U27628 (N_27628,N_25925,N_26385);
nand U27629 (N_27629,N_25863,N_25996);
nand U27630 (N_27630,N_25952,N_26449);
and U27631 (N_27631,N_25693,N_26427);
nand U27632 (N_27632,N_26429,N_26540);
nor U27633 (N_27633,N_25525,N_26125);
nor U27634 (N_27634,N_26611,N_25798);
and U27635 (N_27635,N_26515,N_26771);
nor U27636 (N_27636,N_26330,N_26946);
nor U27637 (N_27637,N_26998,N_26637);
nor U27638 (N_27638,N_25684,N_26192);
and U27639 (N_27639,N_26208,N_26339);
xnor U27640 (N_27640,N_25743,N_25994);
xor U27641 (N_27641,N_25969,N_25924);
or U27642 (N_27642,N_26928,N_26361);
nor U27643 (N_27643,N_26276,N_26233);
nand U27644 (N_27644,N_26567,N_26183);
xnor U27645 (N_27645,N_26614,N_26149);
and U27646 (N_27646,N_25864,N_25726);
xnor U27647 (N_27647,N_26985,N_26963);
xnor U27648 (N_27648,N_26806,N_25850);
nor U27649 (N_27649,N_26506,N_26218);
nand U27650 (N_27650,N_26222,N_26702);
nor U27651 (N_27651,N_26646,N_26477);
nor U27652 (N_27652,N_26872,N_26344);
nand U27653 (N_27653,N_25958,N_25576);
nand U27654 (N_27654,N_26443,N_26104);
and U27655 (N_27655,N_25883,N_26381);
nand U27656 (N_27656,N_26767,N_25677);
nand U27657 (N_27657,N_26263,N_25791);
xnor U27658 (N_27658,N_26975,N_25582);
nand U27659 (N_27659,N_26634,N_26481);
or U27660 (N_27660,N_26796,N_26964);
nor U27661 (N_27661,N_25706,N_25919);
nor U27662 (N_27662,N_26350,N_26994);
xnor U27663 (N_27663,N_25985,N_25918);
nor U27664 (N_27664,N_26190,N_26354);
or U27665 (N_27665,N_26288,N_25779);
nor U27666 (N_27666,N_26787,N_25897);
nor U27667 (N_27667,N_26887,N_26649);
xnor U27668 (N_27668,N_25644,N_26777);
xor U27669 (N_27669,N_26977,N_26933);
or U27670 (N_27670,N_26568,N_26491);
nand U27671 (N_27671,N_26578,N_26009);
and U27672 (N_27672,N_25824,N_26006);
and U27673 (N_27673,N_26128,N_25659);
nor U27674 (N_27674,N_26203,N_25903);
xor U27675 (N_27675,N_26170,N_25990);
xor U27676 (N_27676,N_26808,N_25772);
nand U27677 (N_27677,N_26563,N_25696);
nand U27678 (N_27678,N_26178,N_26886);
or U27679 (N_27679,N_26226,N_26184);
or U27680 (N_27680,N_25845,N_25673);
and U27681 (N_27681,N_26795,N_26431);
or U27682 (N_27682,N_26240,N_25905);
or U27683 (N_27683,N_25936,N_25610);
and U27684 (N_27684,N_25547,N_25501);
nor U27685 (N_27685,N_26321,N_25835);
nor U27686 (N_27686,N_26989,N_25834);
and U27687 (N_27687,N_26439,N_26599);
or U27688 (N_27688,N_26301,N_26619);
nand U27689 (N_27689,N_26154,N_26922);
nand U27690 (N_27690,N_26753,N_26799);
or U27691 (N_27691,N_26898,N_26847);
or U27692 (N_27692,N_26110,N_26262);
xnor U27693 (N_27693,N_26324,N_25640);
xnor U27694 (N_27694,N_25727,N_25914);
and U27695 (N_27695,N_25793,N_26516);
nand U27696 (N_27696,N_26360,N_25971);
or U27697 (N_27697,N_26740,N_25607);
xor U27698 (N_27698,N_25702,N_26548);
or U27699 (N_27699,N_26434,N_26223);
nor U27700 (N_27700,N_25838,N_26849);
nand U27701 (N_27701,N_25648,N_26155);
xor U27702 (N_27702,N_26131,N_25524);
nand U27703 (N_27703,N_25907,N_26065);
nor U27704 (N_27704,N_26587,N_25566);
and U27705 (N_27705,N_26142,N_26738);
nor U27706 (N_27706,N_26997,N_25964);
and U27707 (N_27707,N_25895,N_25997);
nand U27708 (N_27708,N_26880,N_25854);
xnor U27709 (N_27709,N_26780,N_26741);
and U27710 (N_27710,N_26108,N_25760);
and U27711 (N_27711,N_26091,N_26495);
nor U27712 (N_27712,N_25720,N_26210);
nor U27713 (N_27713,N_26831,N_26082);
nand U27714 (N_27714,N_25842,N_25561);
and U27715 (N_27715,N_26709,N_26353);
nor U27716 (N_27716,N_26819,N_26264);
or U27717 (N_27717,N_26338,N_26813);
and U27718 (N_27718,N_26853,N_25837);
nor U27719 (N_27719,N_26669,N_26950);
nand U27720 (N_27720,N_26063,N_26968);
xnor U27721 (N_27721,N_25700,N_26162);
xnor U27722 (N_27722,N_26224,N_26242);
or U27723 (N_27723,N_26442,N_25771);
nand U27724 (N_27724,N_26327,N_26574);
and U27725 (N_27725,N_26268,N_26526);
or U27726 (N_27726,N_26187,N_25638);
or U27727 (N_27727,N_26855,N_26523);
nor U27728 (N_27728,N_26711,N_26839);
nand U27729 (N_27729,N_26132,N_25572);
or U27730 (N_27730,N_26903,N_26316);
nand U27731 (N_27731,N_25508,N_25652);
nor U27732 (N_27732,N_25984,N_26150);
or U27733 (N_27733,N_25830,N_25612);
nand U27734 (N_27734,N_26312,N_26135);
xor U27735 (N_27735,N_25943,N_25788);
or U27736 (N_27736,N_25686,N_26916);
xor U27737 (N_27737,N_26705,N_26182);
xor U27738 (N_27738,N_25604,N_26071);
or U27739 (N_27739,N_26586,N_26422);
nand U27740 (N_27740,N_26871,N_26986);
xor U27741 (N_27741,N_25841,N_26765);
xnor U27742 (N_27742,N_26079,N_26426);
nor U27743 (N_27743,N_26723,N_25707);
xor U27744 (N_27744,N_26534,N_25930);
nand U27745 (N_27745,N_26763,N_26281);
nand U27746 (N_27746,N_25916,N_25993);
nor U27747 (N_27747,N_26754,N_25853);
or U27748 (N_27748,N_26111,N_26769);
xor U27749 (N_27749,N_26879,N_26453);
nand U27750 (N_27750,N_26359,N_26539);
xor U27751 (N_27751,N_26619,N_26884);
or U27752 (N_27752,N_26193,N_26949);
nand U27753 (N_27753,N_25808,N_26241);
nor U27754 (N_27754,N_25716,N_25636);
nor U27755 (N_27755,N_25691,N_25559);
and U27756 (N_27756,N_26882,N_25877);
nand U27757 (N_27757,N_25997,N_25861);
and U27758 (N_27758,N_26098,N_25695);
or U27759 (N_27759,N_25832,N_25797);
nand U27760 (N_27760,N_25824,N_25743);
or U27761 (N_27761,N_25502,N_26976);
nand U27762 (N_27762,N_26929,N_26815);
nand U27763 (N_27763,N_26594,N_26897);
nand U27764 (N_27764,N_26111,N_25616);
nor U27765 (N_27765,N_26938,N_26724);
or U27766 (N_27766,N_26948,N_26842);
nor U27767 (N_27767,N_26519,N_26695);
or U27768 (N_27768,N_26996,N_26382);
nor U27769 (N_27769,N_26557,N_25793);
nor U27770 (N_27770,N_25931,N_26875);
xnor U27771 (N_27771,N_26713,N_26179);
xor U27772 (N_27772,N_26544,N_25965);
or U27773 (N_27773,N_26188,N_25570);
or U27774 (N_27774,N_26821,N_26034);
or U27775 (N_27775,N_25532,N_25983);
nand U27776 (N_27776,N_25639,N_26754);
or U27777 (N_27777,N_25713,N_25958);
nor U27778 (N_27778,N_26971,N_26037);
nand U27779 (N_27779,N_25892,N_25984);
xnor U27780 (N_27780,N_26802,N_26427);
and U27781 (N_27781,N_25856,N_25820);
nand U27782 (N_27782,N_26729,N_26623);
or U27783 (N_27783,N_25848,N_26691);
or U27784 (N_27784,N_26152,N_25904);
nand U27785 (N_27785,N_26082,N_26840);
or U27786 (N_27786,N_25643,N_25707);
nor U27787 (N_27787,N_26445,N_26846);
or U27788 (N_27788,N_26519,N_26952);
or U27789 (N_27789,N_26278,N_26938);
and U27790 (N_27790,N_26821,N_25942);
nand U27791 (N_27791,N_25539,N_26209);
nand U27792 (N_27792,N_25968,N_26521);
or U27793 (N_27793,N_26794,N_26441);
nor U27794 (N_27794,N_26812,N_25901);
nand U27795 (N_27795,N_25874,N_26777);
xor U27796 (N_27796,N_26385,N_26163);
xnor U27797 (N_27797,N_26862,N_25988);
nand U27798 (N_27798,N_26336,N_25565);
or U27799 (N_27799,N_26016,N_25513);
and U27800 (N_27800,N_26596,N_25818);
xnor U27801 (N_27801,N_25883,N_26658);
and U27802 (N_27802,N_26818,N_25909);
xnor U27803 (N_27803,N_25639,N_25699);
nand U27804 (N_27804,N_26779,N_26985);
or U27805 (N_27805,N_26394,N_26210);
nand U27806 (N_27806,N_26053,N_25848);
nand U27807 (N_27807,N_26719,N_26591);
xor U27808 (N_27808,N_26051,N_26118);
and U27809 (N_27809,N_26446,N_25682);
nand U27810 (N_27810,N_25680,N_26194);
xnor U27811 (N_27811,N_26970,N_26194);
xor U27812 (N_27812,N_25947,N_26608);
nor U27813 (N_27813,N_26834,N_25901);
nor U27814 (N_27814,N_26521,N_26369);
or U27815 (N_27815,N_26240,N_26188);
and U27816 (N_27816,N_26879,N_26530);
or U27817 (N_27817,N_26141,N_26532);
nor U27818 (N_27818,N_25573,N_26957);
xor U27819 (N_27819,N_26584,N_25841);
xor U27820 (N_27820,N_25503,N_26152);
or U27821 (N_27821,N_26336,N_25679);
nor U27822 (N_27822,N_26218,N_26661);
nor U27823 (N_27823,N_25835,N_26942);
or U27824 (N_27824,N_26775,N_25727);
or U27825 (N_27825,N_26667,N_26537);
xnor U27826 (N_27826,N_25876,N_26015);
or U27827 (N_27827,N_25521,N_25584);
and U27828 (N_27828,N_26554,N_26912);
or U27829 (N_27829,N_26587,N_26426);
and U27830 (N_27830,N_25960,N_26155);
and U27831 (N_27831,N_26985,N_25807);
and U27832 (N_27832,N_26291,N_25867);
or U27833 (N_27833,N_26663,N_25721);
nand U27834 (N_27834,N_26555,N_25954);
xor U27835 (N_27835,N_26019,N_26408);
nor U27836 (N_27836,N_25522,N_26051);
and U27837 (N_27837,N_26233,N_25993);
or U27838 (N_27838,N_26647,N_25717);
and U27839 (N_27839,N_26851,N_25901);
xor U27840 (N_27840,N_25905,N_26912);
nand U27841 (N_27841,N_26969,N_25969);
and U27842 (N_27842,N_26028,N_26911);
xor U27843 (N_27843,N_25948,N_26769);
or U27844 (N_27844,N_26514,N_26984);
nand U27845 (N_27845,N_26927,N_26373);
or U27846 (N_27846,N_25866,N_26995);
nor U27847 (N_27847,N_25971,N_26481);
or U27848 (N_27848,N_26154,N_26379);
xnor U27849 (N_27849,N_25871,N_26937);
nand U27850 (N_27850,N_25611,N_25561);
nor U27851 (N_27851,N_26468,N_25503);
or U27852 (N_27852,N_26948,N_25775);
xor U27853 (N_27853,N_25736,N_26457);
xor U27854 (N_27854,N_26090,N_25806);
and U27855 (N_27855,N_26441,N_26411);
or U27856 (N_27856,N_25561,N_26484);
xnor U27857 (N_27857,N_25617,N_26048);
and U27858 (N_27858,N_25810,N_25524);
xnor U27859 (N_27859,N_26005,N_26799);
nor U27860 (N_27860,N_26819,N_25874);
nor U27861 (N_27861,N_25594,N_25742);
or U27862 (N_27862,N_25823,N_26682);
xor U27863 (N_27863,N_26908,N_25985);
or U27864 (N_27864,N_26518,N_26410);
or U27865 (N_27865,N_26187,N_26664);
or U27866 (N_27866,N_25740,N_25566);
or U27867 (N_27867,N_26558,N_26285);
nor U27868 (N_27868,N_26416,N_25722);
and U27869 (N_27869,N_25862,N_26782);
nand U27870 (N_27870,N_25893,N_26327);
or U27871 (N_27871,N_25695,N_25939);
nand U27872 (N_27872,N_25985,N_26834);
nor U27873 (N_27873,N_25846,N_26060);
xnor U27874 (N_27874,N_26841,N_25569);
xnor U27875 (N_27875,N_25633,N_26586);
xor U27876 (N_27876,N_25837,N_26518);
or U27877 (N_27877,N_25576,N_26589);
or U27878 (N_27878,N_26576,N_26888);
and U27879 (N_27879,N_26956,N_25701);
or U27880 (N_27880,N_26260,N_25501);
or U27881 (N_27881,N_26003,N_26146);
or U27882 (N_27882,N_26313,N_26950);
nor U27883 (N_27883,N_25881,N_26381);
or U27884 (N_27884,N_26209,N_25684);
xnor U27885 (N_27885,N_26851,N_26914);
or U27886 (N_27886,N_25751,N_26630);
nor U27887 (N_27887,N_26619,N_25655);
xnor U27888 (N_27888,N_25981,N_25864);
xor U27889 (N_27889,N_26238,N_26699);
or U27890 (N_27890,N_25970,N_26143);
or U27891 (N_27891,N_26535,N_26030);
and U27892 (N_27892,N_25591,N_26102);
or U27893 (N_27893,N_26750,N_25934);
nor U27894 (N_27894,N_25652,N_26347);
xor U27895 (N_27895,N_26101,N_26466);
xor U27896 (N_27896,N_25729,N_25987);
xor U27897 (N_27897,N_26630,N_25527);
nand U27898 (N_27898,N_26376,N_26669);
or U27899 (N_27899,N_26849,N_25595);
nand U27900 (N_27900,N_26229,N_26689);
or U27901 (N_27901,N_26928,N_26853);
or U27902 (N_27902,N_26806,N_25883);
nand U27903 (N_27903,N_25885,N_26563);
nand U27904 (N_27904,N_26776,N_25594);
or U27905 (N_27905,N_25508,N_26672);
or U27906 (N_27906,N_26614,N_26259);
and U27907 (N_27907,N_26732,N_26560);
nand U27908 (N_27908,N_26696,N_25955);
or U27909 (N_27909,N_25790,N_26948);
or U27910 (N_27910,N_26181,N_26596);
nor U27911 (N_27911,N_26137,N_26726);
and U27912 (N_27912,N_25878,N_26416);
and U27913 (N_27913,N_26540,N_25615);
or U27914 (N_27914,N_26022,N_26090);
xor U27915 (N_27915,N_26789,N_25876);
and U27916 (N_27916,N_26851,N_26093);
nand U27917 (N_27917,N_26270,N_26403);
or U27918 (N_27918,N_26056,N_26593);
xnor U27919 (N_27919,N_25619,N_25869);
nand U27920 (N_27920,N_25567,N_26877);
and U27921 (N_27921,N_25510,N_26915);
xnor U27922 (N_27922,N_26466,N_26313);
nand U27923 (N_27923,N_26703,N_26971);
and U27924 (N_27924,N_25938,N_25971);
or U27925 (N_27925,N_25657,N_25949);
nor U27926 (N_27926,N_25801,N_26897);
xor U27927 (N_27927,N_26494,N_26646);
nor U27928 (N_27928,N_25773,N_26177);
xnor U27929 (N_27929,N_26307,N_26009);
xnor U27930 (N_27930,N_26678,N_26125);
nand U27931 (N_27931,N_26031,N_26096);
xor U27932 (N_27932,N_26105,N_26580);
nand U27933 (N_27933,N_25588,N_26190);
xnor U27934 (N_27934,N_26040,N_25939);
xnor U27935 (N_27935,N_25690,N_25934);
nor U27936 (N_27936,N_25524,N_26668);
or U27937 (N_27937,N_25519,N_26057);
nor U27938 (N_27938,N_25920,N_26071);
nand U27939 (N_27939,N_26790,N_26788);
and U27940 (N_27940,N_26962,N_26318);
and U27941 (N_27941,N_25921,N_25776);
or U27942 (N_27942,N_26881,N_26225);
and U27943 (N_27943,N_25804,N_26515);
and U27944 (N_27944,N_26788,N_26264);
nor U27945 (N_27945,N_25692,N_26706);
nand U27946 (N_27946,N_26443,N_26303);
or U27947 (N_27947,N_25549,N_26287);
or U27948 (N_27948,N_26559,N_26401);
or U27949 (N_27949,N_26734,N_26348);
or U27950 (N_27950,N_25690,N_26623);
xor U27951 (N_27951,N_26176,N_25657);
and U27952 (N_27952,N_25859,N_25745);
or U27953 (N_27953,N_26691,N_26963);
or U27954 (N_27954,N_25742,N_26210);
nor U27955 (N_27955,N_26855,N_26845);
nor U27956 (N_27956,N_25661,N_26181);
xor U27957 (N_27957,N_25685,N_26070);
nor U27958 (N_27958,N_26844,N_26443);
xor U27959 (N_27959,N_26442,N_26769);
and U27960 (N_27960,N_26321,N_26165);
and U27961 (N_27961,N_26294,N_26945);
or U27962 (N_27962,N_26839,N_26596);
nand U27963 (N_27963,N_26024,N_25544);
nor U27964 (N_27964,N_26321,N_25935);
or U27965 (N_27965,N_26105,N_26707);
and U27966 (N_27966,N_25665,N_26917);
nor U27967 (N_27967,N_25812,N_25863);
nand U27968 (N_27968,N_25953,N_26804);
or U27969 (N_27969,N_26619,N_26203);
and U27970 (N_27970,N_26147,N_26084);
xnor U27971 (N_27971,N_26749,N_26871);
nor U27972 (N_27972,N_25962,N_26601);
and U27973 (N_27973,N_26968,N_25971);
or U27974 (N_27974,N_25911,N_26657);
and U27975 (N_27975,N_25913,N_26461);
and U27976 (N_27976,N_26592,N_25583);
or U27977 (N_27977,N_26029,N_26653);
nand U27978 (N_27978,N_26869,N_25873);
or U27979 (N_27979,N_26190,N_26355);
nor U27980 (N_27980,N_25814,N_25891);
and U27981 (N_27981,N_25787,N_26794);
nor U27982 (N_27982,N_26363,N_25863);
or U27983 (N_27983,N_26130,N_25666);
nor U27984 (N_27984,N_25581,N_26171);
xor U27985 (N_27985,N_25907,N_26927);
xor U27986 (N_27986,N_25900,N_25938);
xnor U27987 (N_27987,N_26540,N_25659);
and U27988 (N_27988,N_26458,N_26838);
nand U27989 (N_27989,N_25829,N_25594);
nor U27990 (N_27990,N_25547,N_26058);
nand U27991 (N_27991,N_26527,N_26017);
nand U27992 (N_27992,N_26135,N_26025);
and U27993 (N_27993,N_25623,N_26279);
and U27994 (N_27994,N_26021,N_26930);
xnor U27995 (N_27995,N_26923,N_26533);
xnor U27996 (N_27996,N_25852,N_26361);
or U27997 (N_27997,N_25589,N_26314);
or U27998 (N_27998,N_25805,N_25886);
nor U27999 (N_27999,N_25616,N_26818);
and U28000 (N_28000,N_26658,N_25607);
xnor U28001 (N_28001,N_26328,N_26410);
or U28002 (N_28002,N_26592,N_25746);
xnor U28003 (N_28003,N_25821,N_26971);
and U28004 (N_28004,N_26005,N_26348);
nand U28005 (N_28005,N_26827,N_26824);
xnor U28006 (N_28006,N_26447,N_26822);
nand U28007 (N_28007,N_26138,N_25863);
and U28008 (N_28008,N_26752,N_25715);
xor U28009 (N_28009,N_26932,N_25958);
nor U28010 (N_28010,N_25511,N_26299);
or U28011 (N_28011,N_26539,N_26085);
and U28012 (N_28012,N_26625,N_25525);
nor U28013 (N_28013,N_26654,N_25992);
nor U28014 (N_28014,N_25606,N_26254);
and U28015 (N_28015,N_25971,N_26886);
nand U28016 (N_28016,N_26392,N_26458);
nand U28017 (N_28017,N_26109,N_26940);
or U28018 (N_28018,N_26328,N_26450);
and U28019 (N_28019,N_26541,N_26011);
xor U28020 (N_28020,N_25615,N_26596);
or U28021 (N_28021,N_26730,N_26559);
nor U28022 (N_28022,N_25516,N_26051);
and U28023 (N_28023,N_25632,N_25538);
nand U28024 (N_28024,N_26281,N_26886);
nor U28025 (N_28025,N_25608,N_26203);
or U28026 (N_28026,N_26431,N_25854);
xnor U28027 (N_28027,N_25555,N_26167);
nand U28028 (N_28028,N_25801,N_26682);
xnor U28029 (N_28029,N_26781,N_25790);
or U28030 (N_28030,N_26231,N_25657);
or U28031 (N_28031,N_26106,N_25813);
nor U28032 (N_28032,N_26980,N_25875);
and U28033 (N_28033,N_25827,N_26017);
xnor U28034 (N_28034,N_26532,N_26264);
and U28035 (N_28035,N_25790,N_26793);
nor U28036 (N_28036,N_26378,N_26882);
xnor U28037 (N_28037,N_26688,N_26246);
or U28038 (N_28038,N_25563,N_26769);
and U28039 (N_28039,N_25818,N_25606);
and U28040 (N_28040,N_25659,N_25948);
nand U28041 (N_28041,N_26261,N_25734);
xor U28042 (N_28042,N_26796,N_26828);
nor U28043 (N_28043,N_26392,N_26223);
nand U28044 (N_28044,N_25503,N_26597);
or U28045 (N_28045,N_26765,N_26149);
and U28046 (N_28046,N_26159,N_26023);
or U28047 (N_28047,N_25783,N_25781);
nand U28048 (N_28048,N_26877,N_25736);
and U28049 (N_28049,N_25731,N_26712);
xor U28050 (N_28050,N_26160,N_25933);
nand U28051 (N_28051,N_25651,N_26401);
nor U28052 (N_28052,N_26070,N_25556);
xor U28053 (N_28053,N_26333,N_26889);
nand U28054 (N_28054,N_26723,N_26638);
nor U28055 (N_28055,N_25838,N_26251);
nand U28056 (N_28056,N_26417,N_25712);
or U28057 (N_28057,N_26791,N_26107);
and U28058 (N_28058,N_26940,N_26159);
xor U28059 (N_28059,N_26902,N_25547);
nand U28060 (N_28060,N_26343,N_25521);
nor U28061 (N_28061,N_25817,N_26587);
nand U28062 (N_28062,N_26220,N_26918);
nand U28063 (N_28063,N_26089,N_26477);
nand U28064 (N_28064,N_25819,N_25975);
nor U28065 (N_28065,N_25692,N_26557);
and U28066 (N_28066,N_26130,N_26573);
xnor U28067 (N_28067,N_25759,N_26651);
xor U28068 (N_28068,N_26373,N_26928);
or U28069 (N_28069,N_26540,N_25524);
xor U28070 (N_28070,N_25696,N_25773);
nor U28071 (N_28071,N_25982,N_26256);
xnor U28072 (N_28072,N_26728,N_25925);
or U28073 (N_28073,N_26592,N_26787);
nor U28074 (N_28074,N_25590,N_25662);
nor U28075 (N_28075,N_26291,N_26546);
and U28076 (N_28076,N_26810,N_26137);
xor U28077 (N_28077,N_26205,N_26419);
or U28078 (N_28078,N_25689,N_26941);
nor U28079 (N_28079,N_26420,N_26774);
nor U28080 (N_28080,N_26272,N_26808);
or U28081 (N_28081,N_26576,N_26740);
or U28082 (N_28082,N_26445,N_26705);
and U28083 (N_28083,N_25742,N_25679);
and U28084 (N_28084,N_25952,N_26811);
or U28085 (N_28085,N_25887,N_25816);
and U28086 (N_28086,N_25999,N_25701);
and U28087 (N_28087,N_26251,N_26404);
nor U28088 (N_28088,N_26197,N_26106);
and U28089 (N_28089,N_26840,N_26750);
nand U28090 (N_28090,N_26295,N_26875);
nor U28091 (N_28091,N_26384,N_26381);
and U28092 (N_28092,N_26652,N_26084);
xnor U28093 (N_28093,N_25903,N_25611);
nand U28094 (N_28094,N_26653,N_26429);
nor U28095 (N_28095,N_26248,N_25690);
and U28096 (N_28096,N_25587,N_26445);
nand U28097 (N_28097,N_26510,N_25518);
nand U28098 (N_28098,N_26643,N_26640);
or U28099 (N_28099,N_26867,N_26511);
nand U28100 (N_28100,N_25969,N_25825);
or U28101 (N_28101,N_26091,N_26888);
nor U28102 (N_28102,N_25980,N_26575);
or U28103 (N_28103,N_25935,N_26290);
nor U28104 (N_28104,N_26853,N_26810);
xor U28105 (N_28105,N_25942,N_26859);
nor U28106 (N_28106,N_25883,N_26415);
xnor U28107 (N_28107,N_26473,N_26439);
nand U28108 (N_28108,N_25726,N_26626);
and U28109 (N_28109,N_26455,N_26440);
xor U28110 (N_28110,N_26924,N_26357);
nand U28111 (N_28111,N_26592,N_25615);
and U28112 (N_28112,N_26650,N_26287);
nor U28113 (N_28113,N_26560,N_25704);
nor U28114 (N_28114,N_26223,N_26985);
or U28115 (N_28115,N_26029,N_25817);
xor U28116 (N_28116,N_26554,N_26162);
nand U28117 (N_28117,N_26580,N_26228);
xnor U28118 (N_28118,N_26453,N_25530);
or U28119 (N_28119,N_25663,N_26947);
nand U28120 (N_28120,N_25850,N_26234);
and U28121 (N_28121,N_26809,N_26746);
nand U28122 (N_28122,N_26727,N_25969);
nand U28123 (N_28123,N_26679,N_25934);
or U28124 (N_28124,N_26522,N_25547);
or U28125 (N_28125,N_26092,N_25964);
nor U28126 (N_28126,N_25944,N_26635);
xor U28127 (N_28127,N_26997,N_26308);
or U28128 (N_28128,N_26054,N_26443);
or U28129 (N_28129,N_26197,N_26840);
or U28130 (N_28130,N_26051,N_26015);
or U28131 (N_28131,N_26825,N_26433);
and U28132 (N_28132,N_26284,N_25963);
xnor U28133 (N_28133,N_26884,N_25519);
nand U28134 (N_28134,N_25707,N_25646);
nor U28135 (N_28135,N_26627,N_25848);
or U28136 (N_28136,N_25610,N_26449);
and U28137 (N_28137,N_25791,N_25983);
xor U28138 (N_28138,N_25732,N_26261);
nand U28139 (N_28139,N_26608,N_25771);
nor U28140 (N_28140,N_26532,N_26176);
xor U28141 (N_28141,N_26180,N_26237);
xor U28142 (N_28142,N_26631,N_25816);
and U28143 (N_28143,N_25804,N_26616);
nor U28144 (N_28144,N_25884,N_25715);
nand U28145 (N_28145,N_26480,N_26978);
and U28146 (N_28146,N_25964,N_26977);
nor U28147 (N_28147,N_25820,N_25555);
nor U28148 (N_28148,N_25849,N_25710);
nand U28149 (N_28149,N_26159,N_26316);
or U28150 (N_28150,N_25625,N_26055);
and U28151 (N_28151,N_26739,N_26081);
nand U28152 (N_28152,N_26844,N_25551);
and U28153 (N_28153,N_26796,N_25701);
and U28154 (N_28154,N_26901,N_25867);
xor U28155 (N_28155,N_25672,N_25944);
xnor U28156 (N_28156,N_26769,N_25961);
and U28157 (N_28157,N_26499,N_26570);
nand U28158 (N_28158,N_26147,N_25865);
nor U28159 (N_28159,N_26238,N_25811);
or U28160 (N_28160,N_26482,N_26448);
or U28161 (N_28161,N_26981,N_26501);
or U28162 (N_28162,N_25794,N_26914);
nor U28163 (N_28163,N_25592,N_26752);
and U28164 (N_28164,N_26087,N_25986);
xor U28165 (N_28165,N_26673,N_25549);
nand U28166 (N_28166,N_26838,N_26639);
nand U28167 (N_28167,N_26683,N_25983);
or U28168 (N_28168,N_26620,N_26984);
and U28169 (N_28169,N_25610,N_25846);
nor U28170 (N_28170,N_26846,N_26860);
or U28171 (N_28171,N_26152,N_26449);
nor U28172 (N_28172,N_26823,N_26458);
xnor U28173 (N_28173,N_25836,N_26989);
and U28174 (N_28174,N_26925,N_25988);
and U28175 (N_28175,N_26473,N_26597);
nand U28176 (N_28176,N_26040,N_25729);
nor U28177 (N_28177,N_26497,N_26351);
nand U28178 (N_28178,N_25881,N_26273);
xnor U28179 (N_28179,N_26427,N_26208);
and U28180 (N_28180,N_25651,N_26118);
nand U28181 (N_28181,N_26806,N_25891);
xor U28182 (N_28182,N_26509,N_26493);
or U28183 (N_28183,N_26630,N_25563);
nor U28184 (N_28184,N_25833,N_26375);
nand U28185 (N_28185,N_26760,N_26478);
nand U28186 (N_28186,N_26796,N_26784);
nor U28187 (N_28187,N_25689,N_26267);
nor U28188 (N_28188,N_26275,N_26245);
and U28189 (N_28189,N_26973,N_25711);
nor U28190 (N_28190,N_25932,N_26434);
nor U28191 (N_28191,N_26670,N_25568);
nand U28192 (N_28192,N_26325,N_26629);
nor U28193 (N_28193,N_26596,N_26160);
nand U28194 (N_28194,N_26545,N_26585);
and U28195 (N_28195,N_26935,N_25728);
xnor U28196 (N_28196,N_25781,N_26515);
nand U28197 (N_28197,N_26728,N_26913);
and U28198 (N_28198,N_26292,N_26122);
nand U28199 (N_28199,N_26529,N_26445);
xor U28200 (N_28200,N_26604,N_25748);
xnor U28201 (N_28201,N_25502,N_26930);
nand U28202 (N_28202,N_26449,N_26430);
nand U28203 (N_28203,N_26088,N_26339);
xnor U28204 (N_28204,N_26455,N_25630);
xnor U28205 (N_28205,N_25815,N_26185);
and U28206 (N_28206,N_26614,N_26322);
xnor U28207 (N_28207,N_26401,N_25710);
and U28208 (N_28208,N_26792,N_25550);
nand U28209 (N_28209,N_26990,N_26536);
xnor U28210 (N_28210,N_25602,N_25556);
or U28211 (N_28211,N_26239,N_26567);
nand U28212 (N_28212,N_26012,N_26063);
and U28213 (N_28213,N_26499,N_26689);
nor U28214 (N_28214,N_25949,N_26566);
and U28215 (N_28215,N_26803,N_26688);
nand U28216 (N_28216,N_25974,N_25808);
or U28217 (N_28217,N_25610,N_26389);
or U28218 (N_28218,N_26433,N_26431);
xnor U28219 (N_28219,N_25809,N_26319);
and U28220 (N_28220,N_26211,N_26618);
and U28221 (N_28221,N_26314,N_26772);
and U28222 (N_28222,N_26006,N_26818);
nor U28223 (N_28223,N_25521,N_26051);
nand U28224 (N_28224,N_25799,N_26386);
or U28225 (N_28225,N_26447,N_26187);
and U28226 (N_28226,N_25852,N_26523);
xor U28227 (N_28227,N_25806,N_25673);
xor U28228 (N_28228,N_25905,N_26325);
nor U28229 (N_28229,N_26452,N_25884);
or U28230 (N_28230,N_25628,N_26194);
nor U28231 (N_28231,N_26229,N_26890);
or U28232 (N_28232,N_26322,N_25882);
nor U28233 (N_28233,N_26131,N_26000);
or U28234 (N_28234,N_25933,N_25972);
xnor U28235 (N_28235,N_26314,N_25970);
and U28236 (N_28236,N_26299,N_25640);
and U28237 (N_28237,N_26524,N_26075);
nor U28238 (N_28238,N_26423,N_26092);
and U28239 (N_28239,N_26167,N_26616);
xnor U28240 (N_28240,N_26596,N_26558);
and U28241 (N_28241,N_25520,N_25615);
nor U28242 (N_28242,N_26068,N_25969);
xnor U28243 (N_28243,N_26624,N_25687);
or U28244 (N_28244,N_25876,N_26159);
and U28245 (N_28245,N_26426,N_26784);
nand U28246 (N_28246,N_25983,N_25920);
and U28247 (N_28247,N_25894,N_25856);
nand U28248 (N_28248,N_26206,N_26616);
and U28249 (N_28249,N_26868,N_26175);
and U28250 (N_28250,N_26553,N_26355);
nor U28251 (N_28251,N_25504,N_26093);
nand U28252 (N_28252,N_26751,N_26691);
xor U28253 (N_28253,N_25807,N_25587);
or U28254 (N_28254,N_25581,N_25707);
and U28255 (N_28255,N_26826,N_25831);
or U28256 (N_28256,N_26617,N_26747);
nor U28257 (N_28257,N_26340,N_25505);
nor U28258 (N_28258,N_26127,N_26893);
nand U28259 (N_28259,N_26895,N_26849);
or U28260 (N_28260,N_26487,N_25863);
xnor U28261 (N_28261,N_26745,N_26772);
nor U28262 (N_28262,N_26752,N_26037);
nand U28263 (N_28263,N_26408,N_25798);
nor U28264 (N_28264,N_25915,N_25905);
or U28265 (N_28265,N_25673,N_26786);
xor U28266 (N_28266,N_26744,N_25736);
and U28267 (N_28267,N_25684,N_26496);
xnor U28268 (N_28268,N_25762,N_26734);
and U28269 (N_28269,N_25672,N_26942);
and U28270 (N_28270,N_25986,N_26150);
nor U28271 (N_28271,N_25617,N_26473);
nor U28272 (N_28272,N_26459,N_25578);
nand U28273 (N_28273,N_26183,N_26631);
and U28274 (N_28274,N_26642,N_26767);
xnor U28275 (N_28275,N_26661,N_26349);
xor U28276 (N_28276,N_26857,N_26629);
xnor U28277 (N_28277,N_26664,N_25959);
nor U28278 (N_28278,N_26426,N_26334);
nor U28279 (N_28279,N_26473,N_26339);
nand U28280 (N_28280,N_26131,N_26392);
xnor U28281 (N_28281,N_26716,N_26167);
xor U28282 (N_28282,N_26745,N_26372);
xor U28283 (N_28283,N_26196,N_25957);
nand U28284 (N_28284,N_25614,N_26066);
and U28285 (N_28285,N_26629,N_26862);
nor U28286 (N_28286,N_25539,N_25888);
nand U28287 (N_28287,N_25716,N_26180);
and U28288 (N_28288,N_25587,N_26505);
nor U28289 (N_28289,N_26623,N_26421);
nand U28290 (N_28290,N_26135,N_26937);
and U28291 (N_28291,N_25630,N_26078);
and U28292 (N_28292,N_26354,N_26660);
nand U28293 (N_28293,N_26346,N_26231);
and U28294 (N_28294,N_25986,N_25909);
nor U28295 (N_28295,N_25557,N_26392);
nor U28296 (N_28296,N_26523,N_26815);
nand U28297 (N_28297,N_26038,N_26691);
xor U28298 (N_28298,N_25665,N_25824);
nor U28299 (N_28299,N_25740,N_26538);
and U28300 (N_28300,N_26879,N_25551);
xor U28301 (N_28301,N_25783,N_25670);
and U28302 (N_28302,N_26904,N_26761);
nor U28303 (N_28303,N_26913,N_26832);
nor U28304 (N_28304,N_25816,N_25711);
nand U28305 (N_28305,N_26069,N_25730);
nand U28306 (N_28306,N_25830,N_25922);
and U28307 (N_28307,N_26094,N_26049);
or U28308 (N_28308,N_26434,N_26695);
nand U28309 (N_28309,N_25898,N_25741);
nor U28310 (N_28310,N_26127,N_26549);
xor U28311 (N_28311,N_26945,N_26661);
or U28312 (N_28312,N_26076,N_25788);
and U28313 (N_28313,N_26412,N_26402);
and U28314 (N_28314,N_25977,N_26582);
xor U28315 (N_28315,N_26312,N_26244);
xor U28316 (N_28316,N_26995,N_26542);
xor U28317 (N_28317,N_26469,N_26384);
nand U28318 (N_28318,N_25511,N_26629);
xnor U28319 (N_28319,N_26923,N_26672);
nand U28320 (N_28320,N_25814,N_26554);
nor U28321 (N_28321,N_26977,N_26177);
xnor U28322 (N_28322,N_26601,N_25535);
nand U28323 (N_28323,N_25659,N_25680);
xnor U28324 (N_28324,N_26477,N_25720);
nor U28325 (N_28325,N_25609,N_26952);
or U28326 (N_28326,N_25748,N_25800);
xnor U28327 (N_28327,N_26452,N_26532);
nor U28328 (N_28328,N_25905,N_26132);
nand U28329 (N_28329,N_26130,N_25892);
nand U28330 (N_28330,N_26649,N_26497);
nand U28331 (N_28331,N_26136,N_26507);
nand U28332 (N_28332,N_25804,N_26201);
nor U28333 (N_28333,N_26728,N_25845);
xor U28334 (N_28334,N_25854,N_26221);
nor U28335 (N_28335,N_25634,N_25848);
nand U28336 (N_28336,N_26657,N_26098);
nand U28337 (N_28337,N_26343,N_26564);
nor U28338 (N_28338,N_26682,N_26381);
and U28339 (N_28339,N_26040,N_25790);
and U28340 (N_28340,N_25767,N_25597);
nand U28341 (N_28341,N_26402,N_26877);
and U28342 (N_28342,N_26335,N_26414);
nand U28343 (N_28343,N_26847,N_26161);
or U28344 (N_28344,N_25686,N_25987);
nand U28345 (N_28345,N_25647,N_26502);
nor U28346 (N_28346,N_26145,N_25913);
nor U28347 (N_28347,N_25508,N_26627);
and U28348 (N_28348,N_26325,N_26372);
nor U28349 (N_28349,N_26554,N_26121);
or U28350 (N_28350,N_26807,N_26420);
and U28351 (N_28351,N_26919,N_26005);
and U28352 (N_28352,N_26310,N_25904);
nor U28353 (N_28353,N_25783,N_26995);
nand U28354 (N_28354,N_26147,N_25998);
nand U28355 (N_28355,N_26600,N_25594);
nor U28356 (N_28356,N_26355,N_26640);
xnor U28357 (N_28357,N_26651,N_26633);
or U28358 (N_28358,N_26530,N_26136);
nand U28359 (N_28359,N_26051,N_25572);
nand U28360 (N_28360,N_26361,N_26765);
and U28361 (N_28361,N_26698,N_26507);
nor U28362 (N_28362,N_26352,N_25634);
nand U28363 (N_28363,N_25810,N_26245);
and U28364 (N_28364,N_25593,N_26490);
nor U28365 (N_28365,N_25942,N_26296);
or U28366 (N_28366,N_26729,N_26642);
xnor U28367 (N_28367,N_26148,N_26963);
or U28368 (N_28368,N_26924,N_25633);
xor U28369 (N_28369,N_25898,N_26009);
xor U28370 (N_28370,N_26630,N_25500);
or U28371 (N_28371,N_26282,N_26157);
nand U28372 (N_28372,N_26588,N_26200);
xnor U28373 (N_28373,N_26693,N_25678);
and U28374 (N_28374,N_25733,N_26692);
or U28375 (N_28375,N_26463,N_26334);
nand U28376 (N_28376,N_26438,N_26102);
nor U28377 (N_28377,N_26391,N_25679);
nor U28378 (N_28378,N_25559,N_26234);
or U28379 (N_28379,N_26706,N_26485);
nand U28380 (N_28380,N_26962,N_26285);
xnor U28381 (N_28381,N_26556,N_26782);
nand U28382 (N_28382,N_26690,N_26348);
nor U28383 (N_28383,N_26746,N_26893);
nand U28384 (N_28384,N_26515,N_26403);
or U28385 (N_28385,N_25697,N_26147);
and U28386 (N_28386,N_26275,N_26276);
nand U28387 (N_28387,N_26774,N_26863);
xor U28388 (N_28388,N_26309,N_26520);
nand U28389 (N_28389,N_25981,N_26387);
xnor U28390 (N_28390,N_25562,N_25744);
xnor U28391 (N_28391,N_26713,N_26574);
and U28392 (N_28392,N_25767,N_26117);
or U28393 (N_28393,N_25666,N_26173);
and U28394 (N_28394,N_25559,N_26562);
or U28395 (N_28395,N_26305,N_25978);
and U28396 (N_28396,N_26338,N_26237);
nor U28397 (N_28397,N_26131,N_26045);
xor U28398 (N_28398,N_25838,N_26866);
and U28399 (N_28399,N_26350,N_26228);
or U28400 (N_28400,N_26403,N_26939);
nand U28401 (N_28401,N_26966,N_25803);
nor U28402 (N_28402,N_26255,N_25676);
nand U28403 (N_28403,N_26990,N_26533);
nand U28404 (N_28404,N_26700,N_25533);
xor U28405 (N_28405,N_25954,N_25573);
and U28406 (N_28406,N_26621,N_26047);
or U28407 (N_28407,N_25972,N_26510);
or U28408 (N_28408,N_26023,N_25798);
xor U28409 (N_28409,N_26471,N_26841);
or U28410 (N_28410,N_26547,N_26139);
or U28411 (N_28411,N_26822,N_26523);
nand U28412 (N_28412,N_26066,N_25689);
nand U28413 (N_28413,N_26804,N_26240);
xnor U28414 (N_28414,N_26200,N_25599);
nor U28415 (N_28415,N_25892,N_26122);
and U28416 (N_28416,N_26225,N_25888);
or U28417 (N_28417,N_26757,N_25754);
nor U28418 (N_28418,N_25538,N_26412);
and U28419 (N_28419,N_26386,N_26787);
nor U28420 (N_28420,N_26965,N_26772);
and U28421 (N_28421,N_25633,N_26671);
or U28422 (N_28422,N_26046,N_26478);
xnor U28423 (N_28423,N_25792,N_25501);
nor U28424 (N_28424,N_26627,N_25550);
nand U28425 (N_28425,N_26804,N_26781);
or U28426 (N_28426,N_26853,N_26077);
xor U28427 (N_28427,N_25856,N_26570);
nor U28428 (N_28428,N_25626,N_26340);
and U28429 (N_28429,N_25685,N_26094);
and U28430 (N_28430,N_26911,N_25536);
xnor U28431 (N_28431,N_26952,N_26249);
xor U28432 (N_28432,N_26975,N_26123);
or U28433 (N_28433,N_26464,N_26627);
nor U28434 (N_28434,N_26539,N_26299);
and U28435 (N_28435,N_25672,N_26269);
xor U28436 (N_28436,N_26582,N_25956);
or U28437 (N_28437,N_26809,N_26034);
nor U28438 (N_28438,N_26373,N_26679);
nand U28439 (N_28439,N_26502,N_26885);
nor U28440 (N_28440,N_25838,N_26527);
nand U28441 (N_28441,N_25987,N_26967);
nor U28442 (N_28442,N_26823,N_26625);
nor U28443 (N_28443,N_25721,N_26990);
xnor U28444 (N_28444,N_26150,N_26090);
xnor U28445 (N_28445,N_26641,N_25762);
and U28446 (N_28446,N_25795,N_26620);
xnor U28447 (N_28447,N_26783,N_26573);
nor U28448 (N_28448,N_25936,N_25620);
xor U28449 (N_28449,N_26969,N_26962);
nor U28450 (N_28450,N_26960,N_26070);
and U28451 (N_28451,N_26632,N_25718);
nand U28452 (N_28452,N_26576,N_25803);
nand U28453 (N_28453,N_26067,N_26969);
xor U28454 (N_28454,N_25853,N_26755);
nand U28455 (N_28455,N_26803,N_26660);
xnor U28456 (N_28456,N_25904,N_26464);
xor U28457 (N_28457,N_26174,N_25801);
and U28458 (N_28458,N_26459,N_25757);
and U28459 (N_28459,N_26055,N_25618);
or U28460 (N_28460,N_25807,N_26957);
nor U28461 (N_28461,N_26577,N_26250);
and U28462 (N_28462,N_26824,N_25915);
nand U28463 (N_28463,N_26412,N_26555);
and U28464 (N_28464,N_26891,N_26524);
xor U28465 (N_28465,N_26914,N_26027);
and U28466 (N_28466,N_26094,N_26257);
and U28467 (N_28467,N_25821,N_26466);
xnor U28468 (N_28468,N_25765,N_26559);
nor U28469 (N_28469,N_26214,N_25858);
or U28470 (N_28470,N_25721,N_25757);
or U28471 (N_28471,N_26201,N_25941);
nor U28472 (N_28472,N_25673,N_25941);
nand U28473 (N_28473,N_26436,N_25829);
nand U28474 (N_28474,N_25999,N_25637);
nand U28475 (N_28475,N_26037,N_26624);
nor U28476 (N_28476,N_26478,N_25759);
nand U28477 (N_28477,N_26353,N_26925);
nand U28478 (N_28478,N_25858,N_26719);
nand U28479 (N_28479,N_25577,N_26407);
or U28480 (N_28480,N_25782,N_26161);
nand U28481 (N_28481,N_25701,N_26547);
nor U28482 (N_28482,N_26455,N_25819);
xnor U28483 (N_28483,N_26481,N_26157);
xor U28484 (N_28484,N_26569,N_26338);
xor U28485 (N_28485,N_26229,N_26432);
xnor U28486 (N_28486,N_26691,N_26231);
or U28487 (N_28487,N_26095,N_26027);
nor U28488 (N_28488,N_25943,N_25995);
and U28489 (N_28489,N_26397,N_26132);
and U28490 (N_28490,N_25821,N_26486);
and U28491 (N_28491,N_26935,N_26250);
and U28492 (N_28492,N_26513,N_26226);
nor U28493 (N_28493,N_26396,N_25750);
nor U28494 (N_28494,N_25824,N_26811);
nand U28495 (N_28495,N_26005,N_26428);
or U28496 (N_28496,N_26390,N_25775);
and U28497 (N_28497,N_25587,N_26763);
nand U28498 (N_28498,N_26934,N_26901);
and U28499 (N_28499,N_25743,N_26773);
nor U28500 (N_28500,N_27148,N_27055);
nor U28501 (N_28501,N_27930,N_28045);
nor U28502 (N_28502,N_27184,N_27793);
or U28503 (N_28503,N_27418,N_27261);
nor U28504 (N_28504,N_28451,N_27673);
or U28505 (N_28505,N_27284,N_27658);
and U28506 (N_28506,N_27698,N_28154);
xor U28507 (N_28507,N_27295,N_27033);
or U28508 (N_28508,N_27165,N_27052);
nor U28509 (N_28509,N_27066,N_27922);
or U28510 (N_28510,N_28215,N_27512);
nand U28511 (N_28511,N_27123,N_28453);
and U28512 (N_28512,N_27352,N_28335);
xor U28513 (N_28513,N_27025,N_27902);
nor U28514 (N_28514,N_27924,N_28290);
and U28515 (N_28515,N_27207,N_27034);
and U28516 (N_28516,N_28002,N_28433);
xor U28517 (N_28517,N_28465,N_27278);
nand U28518 (N_28518,N_27600,N_28308);
or U28519 (N_28519,N_27592,N_28437);
nor U28520 (N_28520,N_28177,N_27120);
and U28521 (N_28521,N_28275,N_28157);
xnor U28522 (N_28522,N_28189,N_27577);
xnor U28523 (N_28523,N_27520,N_28051);
or U28524 (N_28524,N_27555,N_27450);
or U28525 (N_28525,N_28168,N_27378);
and U28526 (N_28526,N_27551,N_28474);
nor U28527 (N_28527,N_28210,N_27508);
nand U28528 (N_28528,N_27903,N_28193);
and U28529 (N_28529,N_27607,N_27294);
nor U28530 (N_28530,N_27029,N_28489);
nand U28531 (N_28531,N_27486,N_27744);
nand U28532 (N_28532,N_28363,N_27259);
nor U28533 (N_28533,N_27711,N_27767);
xnor U28534 (N_28534,N_27832,N_27884);
xor U28535 (N_28535,N_27626,N_27590);
nor U28536 (N_28536,N_27453,N_28485);
xnor U28537 (N_28537,N_28076,N_28438);
or U28538 (N_28538,N_27852,N_27897);
nor U28539 (N_28539,N_27572,N_28120);
xor U28540 (N_28540,N_28225,N_27208);
nand U28541 (N_28541,N_27335,N_27700);
xor U28542 (N_28542,N_27847,N_28094);
xor U28543 (N_28543,N_27712,N_28404);
nor U28544 (N_28544,N_27828,N_27384);
nor U28545 (N_28545,N_27099,N_28414);
nor U28546 (N_28546,N_27297,N_27398);
and U28547 (N_28547,N_28192,N_28163);
xnor U28548 (N_28548,N_27765,N_27763);
nor U28549 (N_28549,N_27535,N_27469);
xnor U28550 (N_28550,N_28462,N_27137);
or U28551 (N_28551,N_27833,N_27826);
nor U28552 (N_28552,N_28080,N_28318);
or U28553 (N_28553,N_27063,N_27468);
nor U28554 (N_28554,N_27650,N_27316);
nor U28555 (N_28555,N_27383,N_28392);
xor U28556 (N_28556,N_27699,N_27608);
and U28557 (N_28557,N_28203,N_28066);
nand U28558 (N_28558,N_28069,N_27532);
and U28559 (N_28559,N_27224,N_27204);
xor U28560 (N_28560,N_28204,N_27357);
nand U28561 (N_28561,N_27989,N_27427);
xor U28562 (N_28562,N_27941,N_27211);
xnor U28563 (N_28563,N_27701,N_27172);
nor U28564 (N_28564,N_28087,N_27812);
nand U28565 (N_28565,N_27946,N_27272);
or U28566 (N_28566,N_27426,N_27642);
nand U28567 (N_28567,N_28181,N_28178);
and U28568 (N_28568,N_27082,N_27027);
or U28569 (N_28569,N_27130,N_27057);
and U28570 (N_28570,N_28315,N_27495);
and U28571 (N_28571,N_27452,N_27973);
and U28572 (N_28572,N_27359,N_28039);
and U28573 (N_28573,N_27474,N_28011);
xor U28574 (N_28574,N_27375,N_27686);
xnor U28575 (N_28575,N_28243,N_27132);
nand U28576 (N_28576,N_27169,N_27938);
xnor U28577 (N_28577,N_27678,N_28387);
xor U28578 (N_28578,N_27872,N_28446);
nand U28579 (N_28579,N_27346,N_27965);
and U28580 (N_28580,N_27787,N_27436);
nor U28581 (N_28581,N_28077,N_27374);
or U28582 (N_28582,N_27772,N_28361);
nand U28583 (N_28583,N_27522,N_28072);
or U28584 (N_28584,N_27283,N_27933);
nor U28585 (N_28585,N_27843,N_27669);
or U28586 (N_28586,N_27153,N_27684);
nand U28587 (N_28587,N_27781,N_28382);
nor U28588 (N_28588,N_27963,N_27260);
xnor U28589 (N_28589,N_28369,N_27079);
or U28590 (N_28590,N_28434,N_28420);
nand U28591 (N_28591,N_27918,N_27072);
or U28592 (N_28592,N_28262,N_28377);
and U28593 (N_28593,N_28264,N_28050);
or U28594 (N_28594,N_27019,N_27271);
nand U28595 (N_28595,N_27596,N_28075);
nor U28596 (N_28596,N_28013,N_27156);
nor U28597 (N_28597,N_27853,N_28353);
or U28598 (N_28598,N_28017,N_27603);
or U28599 (N_28599,N_28313,N_27007);
and U28600 (N_28600,N_27097,N_27824);
nor U28601 (N_28601,N_28358,N_27906);
xnor U28602 (N_28602,N_27149,N_27714);
and U28603 (N_28603,N_28143,N_27205);
or U28604 (N_28604,N_27125,N_27320);
and U28605 (N_28605,N_28411,N_27877);
xor U28606 (N_28606,N_28252,N_28003);
xnor U28607 (N_28607,N_27147,N_27430);
xor U28608 (N_28608,N_27764,N_28067);
xor U28609 (N_28609,N_27223,N_28199);
nor U28610 (N_28610,N_27249,N_28498);
xnor U28611 (N_28611,N_27966,N_28138);
nor U28612 (N_28612,N_27410,N_28037);
xnor U28613 (N_28613,N_27245,N_28319);
nor U28614 (N_28614,N_28195,N_27371);
and U28615 (N_28615,N_27301,N_28398);
nand U28616 (N_28616,N_27862,N_27408);
nand U28617 (N_28617,N_27431,N_27662);
and U28618 (N_28618,N_27655,N_27598);
or U28619 (N_28619,N_27361,N_27492);
xor U28620 (N_28620,N_28025,N_27228);
or U28621 (N_28621,N_28337,N_27671);
xor U28622 (N_28622,N_28183,N_28468);
nor U28623 (N_28623,N_27717,N_28062);
xnor U28624 (N_28624,N_28359,N_27256);
or U28625 (N_28625,N_28022,N_27067);
xor U28626 (N_28626,N_27370,N_27854);
nor U28627 (N_28627,N_28108,N_28090);
and U28628 (N_28628,N_28127,N_27660);
xor U28629 (N_28629,N_27144,N_27885);
xor U28630 (N_28630,N_27643,N_28493);
xnor U28631 (N_28631,N_27730,N_27031);
nor U28632 (N_28632,N_28431,N_27974);
nand U28633 (N_28633,N_27285,N_28015);
nor U28634 (N_28634,N_27194,N_27244);
xor U28635 (N_28635,N_28009,N_28081);
or U28636 (N_28636,N_27951,N_27849);
nand U28637 (N_28637,N_27950,N_27338);
nand U28638 (N_28638,N_27788,N_27177);
nor U28639 (N_28639,N_27179,N_27612);
nor U28640 (N_28640,N_27387,N_28277);
or U28641 (N_28641,N_27583,N_27858);
and U28642 (N_28642,N_28299,N_27518);
and U28643 (N_28643,N_27102,N_27242);
or U28644 (N_28644,N_27571,N_27980);
xnor U28645 (N_28645,N_27866,N_28164);
and U28646 (N_28646,N_28055,N_27813);
nand U28647 (N_28647,N_27026,N_27108);
nand U28648 (N_28648,N_27775,N_27073);
nand U28649 (N_28649,N_27329,N_27797);
nand U28650 (N_28650,N_27065,N_27308);
nor U28651 (N_28651,N_27332,N_27106);
and U28652 (N_28652,N_27564,N_27936);
nor U28653 (N_28653,N_28410,N_27731);
xor U28654 (N_28654,N_27913,N_28146);
xor U28655 (N_28655,N_27038,N_27821);
nor U28656 (N_28656,N_27054,N_27347);
nand U28657 (N_28657,N_28091,N_27488);
xor U28658 (N_28658,N_27747,N_28294);
nor U28659 (N_28659,N_27243,N_27185);
nand U28660 (N_28660,N_27210,N_27089);
nor U28661 (N_28661,N_27039,N_27188);
xnor U28662 (N_28662,N_27085,N_27251);
and U28663 (N_28663,N_28245,N_27083);
nor U28664 (N_28664,N_28071,N_28479);
xnor U28665 (N_28665,N_27823,N_27511);
nor U28666 (N_28666,N_28060,N_28461);
nor U28667 (N_28667,N_27349,N_27726);
and U28668 (N_28668,N_27263,N_27516);
or U28669 (N_28669,N_27388,N_27032);
or U28670 (N_28670,N_27392,N_27127);
nand U28671 (N_28671,N_27619,N_27424);
xnor U28672 (N_28672,N_27562,N_27266);
or U28673 (N_28673,N_28208,N_27888);
and U28674 (N_28674,N_27623,N_28028);
or U28675 (N_28675,N_27136,N_27984);
xnor U28676 (N_28676,N_27445,N_27118);
and U28677 (N_28677,N_28267,N_28268);
nand U28678 (N_28678,N_27000,N_27735);
or U28679 (N_28679,N_28351,N_28161);
nand U28680 (N_28680,N_28310,N_28448);
nor U28681 (N_28681,N_27462,N_28038);
or U28682 (N_28682,N_28046,N_27561);
and U28683 (N_28683,N_28234,N_27479);
or U28684 (N_28684,N_27504,N_27956);
and U28685 (N_28685,N_28360,N_27088);
xnor U28686 (N_28686,N_27459,N_27501);
and U28687 (N_28687,N_28006,N_27454);
nor U28688 (N_28688,N_27421,N_28001);
or U28689 (N_28689,N_28226,N_27934);
and U28690 (N_28690,N_27287,N_27560);
nor U28691 (N_28691,N_28248,N_27901);
nand U28692 (N_28692,N_28336,N_28439);
nor U28693 (N_28693,N_27992,N_28324);
xnor U28694 (N_28694,N_28117,N_27203);
nor U28695 (N_28695,N_28463,N_28396);
and U28696 (N_28696,N_27931,N_27928);
and U28697 (N_28697,N_28135,N_28292);
nor U28698 (N_28698,N_28271,N_27745);
and U28699 (N_28699,N_27559,N_27354);
nor U28700 (N_28700,N_27896,N_27386);
nor U28701 (N_28701,N_27815,N_28171);
or U28702 (N_28702,N_28004,N_28123);
xnor U28703 (N_28703,N_28249,N_27799);
nand U28704 (N_28704,N_27939,N_27690);
and U28705 (N_28705,N_27145,N_27706);
nor U28706 (N_28706,N_28085,N_28409);
nor U28707 (N_28707,N_27523,N_28469);
nor U28708 (N_28708,N_27311,N_28442);
xor U28709 (N_28709,N_27809,N_27363);
or U28710 (N_28710,N_27013,N_27860);
nand U28711 (N_28711,N_27659,N_28147);
xnor U28712 (N_28712,N_27570,N_28390);
xor U28713 (N_28713,N_27192,N_27962);
nand U28714 (N_28714,N_28137,N_27566);
nand U28715 (N_28715,N_28429,N_28124);
nand U28716 (N_28716,N_27330,N_28356);
and U28717 (N_28717,N_27811,N_27327);
nor U28718 (N_28718,N_28238,N_28481);
xor U28719 (N_28719,N_28052,N_28441);
nand U28720 (N_28720,N_27369,N_27389);
xor U28721 (N_28721,N_28088,N_27954);
and U28722 (N_28722,N_28179,N_28328);
xnor U28723 (N_28723,N_27306,N_28298);
and U28724 (N_28724,N_27538,N_27317);
nor U28725 (N_28725,N_27176,N_27126);
nor U28726 (N_28726,N_28174,N_27842);
or U28727 (N_28727,N_27546,N_28029);
nand U28728 (N_28728,N_28343,N_27634);
xor U28729 (N_28729,N_27151,N_27554);
nand U28730 (N_28730,N_27796,N_28136);
xnor U28731 (N_28731,N_28272,N_27845);
or U28732 (N_28732,N_27423,N_27611);
or U28733 (N_28733,N_27952,N_27157);
or U28734 (N_28734,N_28340,N_27978);
nand U28735 (N_28735,N_27890,N_28338);
nor U28736 (N_28736,N_27653,N_27798);
xor U28737 (N_28737,N_27140,N_28300);
xnor U28738 (N_28738,N_28227,N_27968);
nand U28739 (N_28739,N_27290,N_27752);
or U28740 (N_28740,N_27233,N_28033);
or U28741 (N_28741,N_28084,N_27128);
xor U28742 (N_28742,N_28365,N_28008);
xnor U28743 (N_28743,N_27979,N_27892);
nand U28744 (N_28744,N_28099,N_28421);
and U28745 (N_28745,N_28016,N_27616);
nor U28746 (N_28746,N_27725,N_27983);
and U28747 (N_28747,N_27355,N_27341);
nand U28748 (N_28748,N_27475,N_27161);
or U28749 (N_28749,N_27344,N_27806);
and U28750 (N_28750,N_27414,N_27925);
and U28751 (N_28751,N_27870,N_28413);
xnor U28752 (N_28752,N_27691,N_28191);
and U28753 (N_28753,N_28041,N_27433);
xnor U28754 (N_28754,N_27785,N_28371);
nor U28755 (N_28755,N_27158,N_27171);
xor U28756 (N_28756,N_27834,N_28184);
and U28757 (N_28757,N_28422,N_27792);
nor U28758 (N_28758,N_27882,N_27718);
and U28759 (N_28759,N_27293,N_27040);
xor U28760 (N_28760,N_27539,N_27986);
and U28761 (N_28761,N_27489,N_28366);
nor U28762 (N_28762,N_28348,N_27621);
nor U28763 (N_28763,N_27578,N_27377);
nand U28764 (N_28764,N_27281,N_28381);
and U28765 (N_28765,N_28296,N_28027);
nor U28766 (N_28766,N_27343,N_27222);
nand U28767 (N_28767,N_27961,N_28142);
nor U28768 (N_28768,N_27439,N_27337);
nor U28769 (N_28769,N_28251,N_27837);
or U28770 (N_28770,N_27919,N_28211);
nand U28771 (N_28771,N_27982,N_28048);
xnor U28772 (N_28772,N_27345,N_28187);
nand U28773 (N_28773,N_27782,N_27446);
and U28774 (N_28774,N_28201,N_27498);
and U28775 (N_28775,N_28059,N_27248);
and U28776 (N_28776,N_28301,N_27727);
xnor U28777 (N_28777,N_27060,N_28418);
nor U28778 (N_28778,N_27456,N_28326);
nand U28779 (N_28779,N_27051,N_27746);
or U28780 (N_28780,N_28276,N_28070);
nor U28781 (N_28781,N_27069,N_27519);
xnor U28782 (N_28782,N_27753,N_28098);
or U28783 (N_28783,N_28162,N_27693);
nor U28784 (N_28784,N_28035,N_28477);
and U28785 (N_28785,N_28334,N_27117);
xnor U28786 (N_28786,N_28349,N_28018);
nor U28787 (N_28787,N_27661,N_28406);
and U28788 (N_28788,N_27995,N_28408);
and U28789 (N_28789,N_27390,N_27976);
nor U28790 (N_28790,N_28456,N_27993);
xnor U28791 (N_28791,N_28188,N_27315);
xnor U28792 (N_28792,N_28110,N_27307);
or U28793 (N_28793,N_28424,N_27556);
xnor U28794 (N_28794,N_27460,N_28233);
xor U28795 (N_28795,N_28492,N_28190);
and U28796 (N_28796,N_27422,N_27231);
nor U28797 (N_28797,N_28374,N_27086);
nand U28798 (N_28798,N_28364,N_27526);
xnor U28799 (N_28799,N_27981,N_27373);
or U28800 (N_28800,N_28128,N_27850);
nor U28801 (N_28801,N_27791,N_28295);
or U28802 (N_28802,N_28383,N_28397);
nor U28803 (N_28803,N_27865,N_27720);
nand U28804 (N_28804,N_27017,N_27757);
nand U28805 (N_28805,N_27124,N_28219);
xnor U28806 (N_28806,N_27841,N_27942);
nand U28807 (N_28807,N_28430,N_28362);
and U28808 (N_28808,N_28169,N_27937);
and U28809 (N_28809,N_28395,N_27304);
nor U28810 (N_28810,N_27232,N_27401);
nor U28811 (N_28811,N_28288,N_27601);
nand U28812 (N_28812,N_27904,N_28172);
and U28813 (N_28813,N_27816,N_27152);
or U28814 (N_28814,N_28475,N_28165);
xnor U28815 (N_28815,N_27695,N_27071);
nand U28816 (N_28816,N_27531,N_28419);
or U28817 (N_28817,N_27759,N_27114);
nand U28818 (N_28818,N_28176,N_27298);
nand U28819 (N_28819,N_28394,N_28281);
or U28820 (N_28820,N_28079,N_27497);
xor U28821 (N_28821,N_28255,N_28471);
nor U28822 (N_28822,N_27943,N_28487);
xnor U28823 (N_28823,N_28155,N_28043);
and U28824 (N_28824,N_27874,N_28266);
nand U28825 (N_28825,N_27372,N_27536);
or U28826 (N_28826,N_27397,N_27366);
xor U28827 (N_28827,N_27226,N_27457);
or U28828 (N_28828,N_27473,N_28150);
or U28829 (N_28829,N_27719,N_28068);
and U28830 (N_28830,N_27513,N_28236);
nand U28831 (N_28831,N_27585,N_27776);
and U28832 (N_28832,N_27328,N_28415);
or U28833 (N_28833,N_28218,N_27737);
or U28834 (N_28834,N_27042,N_28170);
nor U28835 (N_28835,N_27676,N_27987);
or U28836 (N_28836,N_27738,N_28024);
and U28837 (N_28837,N_27289,N_27217);
and U28838 (N_28838,N_28488,N_27070);
nand U28839 (N_28839,N_27638,N_27324);
and U28840 (N_28840,N_28105,N_27923);
xor U28841 (N_28841,N_28270,N_28283);
xnor U28842 (N_28842,N_27325,N_27133);
nor U28843 (N_28843,N_28460,N_27291);
and U28844 (N_28844,N_27444,N_28258);
nor U28845 (N_28845,N_28242,N_28486);
xnor U28846 (N_28846,N_27202,N_27722);
or U28847 (N_28847,N_27407,N_27964);
xor U28848 (N_28848,N_27754,N_27893);
nand U28849 (N_28849,N_28054,N_28470);
and U28850 (N_28850,N_27170,N_27021);
and U28851 (N_28851,N_27863,N_27053);
or U28852 (N_28852,N_28092,N_27356);
nor U28853 (N_28853,N_27182,N_27552);
xor U28854 (N_28854,N_28432,N_27958);
and U28855 (N_28855,N_27098,N_27008);
nor U28856 (N_28856,N_27247,N_27620);
and U28857 (N_28857,N_28257,N_27895);
nand U28858 (N_28858,N_27802,N_27351);
nand U28859 (N_28859,N_27804,N_27685);
and U28860 (N_28860,N_27898,N_28194);
or U28861 (N_28861,N_27005,N_27563);
nand U28862 (N_28862,N_28400,N_28244);
or U28863 (N_28863,N_27191,N_27020);
and U28864 (N_28864,N_28156,N_27379);
and U28865 (N_28865,N_28320,N_27448);
or U28866 (N_28866,N_27610,N_27449);
nand U28867 (N_28867,N_27839,N_27265);
xor U28868 (N_28868,N_27141,N_27829);
nand U28869 (N_28869,N_27894,N_27011);
and U28870 (N_28870,N_28153,N_28376);
and U28871 (N_28871,N_28274,N_27167);
and U28872 (N_28872,N_27920,N_27437);
nor U28873 (N_28873,N_27393,N_27309);
or U28874 (N_28874,N_27944,N_28223);
and U28875 (N_28875,N_27879,N_27689);
nand U28876 (N_28876,N_28206,N_27269);
nand U28877 (N_28877,N_27527,N_28370);
xor U28878 (N_28878,N_27368,N_27221);
xnor U28879 (N_28879,N_27971,N_27499);
and U28880 (N_28880,N_28316,N_27514);
xor U28881 (N_28881,N_27640,N_27047);
xnor U28882 (N_28882,N_27274,N_27030);
and U28883 (N_28883,N_27576,N_27945);
nor U28884 (N_28884,N_27183,N_28061);
xnor U28885 (N_28885,N_27783,N_28480);
or U28886 (N_28886,N_27012,N_27164);
nor U28887 (N_28887,N_27899,N_27641);
nand U28888 (N_28888,N_27035,N_27087);
xnor U28889 (N_28889,N_28247,N_28232);
xnor U28890 (N_28890,N_28435,N_27569);
nor U28891 (N_28891,N_28209,N_27955);
xor U28892 (N_28892,N_27908,N_27014);
xnor U28893 (N_28893,N_28005,N_27743);
or U28894 (N_28894,N_28352,N_28265);
xnor U28895 (N_28895,N_27022,N_28286);
and U28896 (N_28896,N_27517,N_28454);
xor U28897 (N_28897,N_27728,N_27400);
or U28898 (N_28898,N_27624,N_28014);
nand U28899 (N_28899,N_28472,N_27680);
nand U28900 (N_28900,N_27502,N_27557);
and U28901 (N_28901,N_28386,N_28333);
xnor U28902 (N_28902,N_27362,N_27413);
xor U28903 (N_28903,N_28200,N_27645);
nor U28904 (N_28904,N_27786,N_27595);
nor U28905 (N_28905,N_27059,N_28101);
and U28906 (N_28906,N_28484,N_27886);
or U28907 (N_28907,N_28303,N_27580);
nor U28908 (N_28908,N_28196,N_27957);
and U28909 (N_28909,N_28350,N_28132);
nor U28910 (N_28910,N_28134,N_27822);
nand U28911 (N_28911,N_27268,N_27048);
xnor U28912 (N_28912,N_28102,N_27139);
or U28913 (N_28913,N_27003,N_27288);
nor U28914 (N_28914,N_27058,N_28354);
nand U28915 (N_28915,N_27541,N_27314);
and U28916 (N_28916,N_28263,N_28185);
xor U28917 (N_28917,N_28259,N_27105);
and U28918 (N_28918,N_28086,N_27827);
nand U28919 (N_28919,N_27679,N_27104);
xor U28920 (N_28920,N_27166,N_28254);
or U28921 (N_28921,N_27323,N_28007);
nor U28922 (N_28922,N_28133,N_27675);
or U28923 (N_28923,N_27713,N_27458);
xnor U28924 (N_28924,N_28246,N_28447);
and U28925 (N_28925,N_27146,N_27322);
xor U28926 (N_28926,N_27415,N_27509);
nor U28927 (N_28927,N_27246,N_28260);
and U28928 (N_28928,N_27733,N_27932);
and U28929 (N_28929,N_28104,N_27927);
nand U28930 (N_28930,N_27991,N_28329);
nor U28931 (N_28931,N_27235,N_27574);
xor U28932 (N_28932,N_28000,N_27113);
nor U28933 (N_28933,N_27049,N_28455);
nand U28934 (N_28934,N_27360,N_27867);
and U28935 (N_28935,N_28314,N_27190);
xor U28936 (N_28936,N_27078,N_28368);
xnor U28937 (N_28937,N_27443,N_27209);
nand U28938 (N_28938,N_27900,N_27773);
nand U28939 (N_28939,N_28482,N_27681);
nand U28940 (N_28940,N_28113,N_27622);
or U28941 (N_28941,N_27455,N_27084);
and U28942 (N_28942,N_28149,N_27544);
nand U28943 (N_28943,N_28309,N_27573);
and U28944 (N_28944,N_27740,N_28040);
xnor U28945 (N_28945,N_28180,N_27947);
xor U28946 (N_28946,N_27302,N_27218);
nand U28947 (N_28947,N_27061,N_28426);
and U28948 (N_28948,N_27736,N_28097);
nor U28949 (N_28949,N_28483,N_27334);
xor U28950 (N_28950,N_27588,N_27214);
nand U28951 (N_28951,N_27134,N_28031);
and U28952 (N_28952,N_27748,N_27672);
nor U28953 (N_28953,N_28273,N_28116);
or U28954 (N_28954,N_27004,N_27817);
xnor U28955 (N_28955,N_27568,N_27006);
nand U28956 (N_28956,N_27694,N_27227);
xor U28957 (N_28957,N_27461,N_27476);
or U28958 (N_28958,N_27724,N_28457);
nand U28959 (N_28959,N_28373,N_27688);
nand U28960 (N_28960,N_27530,N_27162);
and U28961 (N_28961,N_27257,N_27887);
and U28962 (N_28962,N_27500,N_27254);
or U28963 (N_28963,N_27609,N_27666);
or U28964 (N_28964,N_27805,N_27239);
nor U28965 (N_28965,N_28466,N_27844);
xnor U28966 (N_28966,N_28095,N_27131);
nor U28967 (N_28967,N_27447,N_27432);
nand U28968 (N_28968,N_28427,N_28393);
nand U28969 (N_28969,N_27674,N_27216);
and U28970 (N_28970,N_27875,N_28220);
nand U28971 (N_28971,N_27312,N_27471);
nor U28972 (N_28972,N_27094,N_27543);
or U28973 (N_28973,N_27339,N_28034);
nand U28974 (N_28974,N_28239,N_27808);
xor U28975 (N_28975,N_27403,N_28384);
nor U28976 (N_28976,N_27093,N_27545);
xnor U28977 (N_28977,N_28312,N_27037);
nand U28978 (N_28978,N_28074,N_28036);
and U28979 (N_28979,N_28221,N_27091);
xor U28980 (N_28980,N_28083,N_28473);
or U28981 (N_28981,N_27173,N_27534);
nor U28982 (N_28982,N_27163,N_27593);
nor U28983 (N_28983,N_28152,N_27800);
nor U28984 (N_28984,N_28436,N_27604);
and U28985 (N_28985,N_28224,N_28240);
nand U28986 (N_28986,N_27646,N_27507);
nand U28987 (N_28987,N_27972,N_28096);
and U28988 (N_28988,N_27493,N_27252);
and U28989 (N_28989,N_27967,N_28205);
nand U28990 (N_28990,N_27766,N_27883);
nor U28991 (N_28991,N_27665,N_27487);
xnor U28992 (N_28992,N_27648,N_28444);
xor U28993 (N_28993,N_27081,N_27734);
or U28994 (N_28994,N_27451,N_28339);
or U28995 (N_28995,N_28425,N_27491);
or U28996 (N_28996,N_27442,N_28216);
xnor U28997 (N_28997,N_28388,N_28304);
or U28998 (N_28998,N_27411,N_28241);
nand U28999 (N_28999,N_27599,N_27174);
nor U29000 (N_29000,N_28023,N_27286);
or U29001 (N_29001,N_27770,N_28228);
or U29002 (N_29002,N_27705,N_27365);
xor U29003 (N_29003,N_27280,N_27825);
or U29004 (N_29004,N_27579,N_27396);
xor U29005 (N_29005,N_28082,N_28144);
or U29006 (N_29006,N_28341,N_27318);
nor U29007 (N_29007,N_28121,N_28499);
xnor U29008 (N_29008,N_28278,N_28167);
xnor U29009 (N_29009,N_28063,N_27189);
nor U29010 (N_29010,N_28412,N_27382);
xor U29011 (N_29011,N_27510,N_27756);
nand U29012 (N_29012,N_27855,N_27168);
xor U29013 (N_29013,N_28126,N_27614);
xor U29014 (N_29014,N_27505,N_27321);
and U29015 (N_29015,N_28139,N_28158);
or U29016 (N_29016,N_27417,N_28237);
or U29017 (N_29017,N_28151,N_28385);
nor U29018 (N_29018,N_28464,N_27819);
nor U29019 (N_29019,N_27631,N_28399);
and U29020 (N_29020,N_27279,N_27116);
nor U29021 (N_29021,N_28289,N_27840);
nand U29022 (N_29022,N_27016,N_28458);
nor U29023 (N_29023,N_28159,N_28428);
nand U29024 (N_29024,N_27046,N_28306);
nor U29025 (N_29025,N_27404,N_28450);
and U29026 (N_29026,N_28214,N_27969);
nor U29027 (N_29027,N_28020,N_28285);
or U29028 (N_29028,N_28182,N_27250);
and U29029 (N_29029,N_27213,N_27768);
nor U29030 (N_29030,N_28122,N_27594);
nand U29031 (N_29031,N_27441,N_28064);
or U29032 (N_29032,N_28322,N_27703);
nor U29033 (N_29033,N_27138,N_27529);
xnor U29034 (N_29034,N_27024,N_28287);
or U29035 (N_29035,N_27935,N_27692);
nor U29036 (N_29036,N_27336,N_27652);
nor U29037 (N_29037,N_27683,N_27319);
or U29038 (N_29038,N_27219,N_27112);
nor U29039 (N_29039,N_28297,N_28284);
or U29040 (N_29040,N_27632,N_27515);
xor U29041 (N_29041,N_27225,N_27466);
nand U29042 (N_29042,N_27023,N_27528);
xor U29043 (N_29043,N_27220,N_27409);
and U29044 (N_29044,N_27873,N_27953);
xnor U29045 (N_29045,N_28405,N_27831);
and U29046 (N_29046,N_28119,N_28131);
or U29047 (N_29047,N_27416,N_27434);
nand U29048 (N_29048,N_27670,N_28357);
nand U29049 (N_29049,N_27630,N_28261);
and U29050 (N_29050,N_27790,N_28230);
and U29051 (N_29051,N_27716,N_28129);
xor U29052 (N_29052,N_27615,N_27503);
or U29053 (N_29053,N_27095,N_27778);
xor U29054 (N_29054,N_27708,N_27236);
nand U29055 (N_29055,N_27869,N_27876);
and U29056 (N_29056,N_27150,N_27878);
xor U29057 (N_29057,N_27779,N_28056);
nor U29058 (N_29058,N_27197,N_27077);
xnor U29059 (N_29059,N_28323,N_27582);
xnor U29060 (N_29060,N_28445,N_27749);
nand U29061 (N_29061,N_27575,N_28293);
nor U29062 (N_29062,N_28440,N_28111);
or U29063 (N_29063,N_28291,N_27677);
and U29064 (N_29064,N_28073,N_28217);
nand U29065 (N_29065,N_28166,N_28311);
or U29066 (N_29066,N_27477,N_28375);
nor U29067 (N_29067,N_27997,N_27709);
xor U29068 (N_29068,N_28402,N_27143);
and U29069 (N_29069,N_28279,N_28417);
or U29070 (N_29070,N_27107,N_27122);
or U29071 (N_29071,N_28269,N_27056);
or U29072 (N_29072,N_27741,N_27277);
and U29073 (N_29073,N_27729,N_27540);
or U29074 (N_29074,N_28331,N_27348);
nor U29075 (N_29075,N_27696,N_27649);
nand U29076 (N_29076,N_28250,N_27267);
nor U29077 (N_29077,N_28367,N_27109);
nor U29078 (N_29078,N_28103,N_27342);
xor U29079 (N_29079,N_28186,N_27484);
or U29080 (N_29080,N_27292,N_27912);
nor U29081 (N_29081,N_27960,N_27230);
and U29082 (N_29082,N_27795,N_27350);
xnor U29083 (N_29083,N_27784,N_27542);
and U29084 (N_29084,N_27975,N_27206);
and U29085 (N_29085,N_27394,N_27506);
xor U29086 (N_29086,N_28112,N_28065);
or U29087 (N_29087,N_27110,N_27181);
and U29088 (N_29088,N_28021,N_27399);
xnor U29089 (N_29089,N_28235,N_27241);
nor U29090 (N_29090,N_27429,N_27999);
and U29091 (N_29091,N_27115,N_27533);
nor U29092 (N_29092,N_27159,N_27627);
and U29093 (N_29093,N_28459,N_28495);
xnor U29094 (N_29094,N_27076,N_28089);
xor U29095 (N_29095,N_27597,N_27949);
or U29096 (N_29096,N_27589,N_27618);
and U29097 (N_29097,N_27376,N_28449);
nand U29098 (N_29098,N_28231,N_27915);
and U29099 (N_29099,N_27009,N_27521);
nor U29100 (N_29100,N_27440,N_28042);
and U29101 (N_29101,N_27914,N_28130);
nand U29102 (N_29102,N_27358,N_27485);
nor U29103 (N_29103,N_27910,N_27856);
or U29104 (N_29104,N_27818,N_28141);
nand U29105 (N_29105,N_27155,N_27300);
nand U29106 (N_29106,N_27402,N_28280);
xor U29107 (N_29107,N_27036,N_27657);
xor U29108 (N_29108,N_28019,N_28145);
nand U29109 (N_29109,N_27663,N_27810);
or U29110 (N_29110,N_28403,N_28491);
nor U29111 (N_29111,N_27111,N_28452);
and U29112 (N_29112,N_27723,N_27715);
nor U29113 (N_29113,N_27835,N_27881);
nand U29114 (N_29114,N_27135,N_28494);
xnor U29115 (N_29115,N_28478,N_27212);
or U29116 (N_29116,N_28173,N_27606);
xnor U29117 (N_29117,N_27644,N_28253);
nand U29118 (N_29118,N_28327,N_27326);
or U29119 (N_29119,N_27435,N_27917);
xor U29120 (N_29120,N_28213,N_27175);
or U29121 (N_29121,N_27353,N_27121);
or U29122 (N_29122,N_28355,N_28305);
and U29123 (N_29123,N_27907,N_27229);
and U29124 (N_29124,N_27142,N_27921);
or U29125 (N_29125,N_27481,N_27187);
nor U29126 (N_29126,N_28378,N_27438);
or U29127 (N_29127,N_27769,N_27463);
nor U29128 (N_29128,N_27959,N_28125);
and U29129 (N_29129,N_27732,N_27483);
or U29130 (N_29130,N_27103,N_27010);
xor U29131 (N_29131,N_28148,N_27820);
or U29132 (N_29132,N_28391,N_27758);
nand U29133 (N_29133,N_27742,N_27859);
or U29134 (N_29134,N_27186,N_27668);
xor U29135 (N_29135,N_28078,N_27864);
nor U29136 (N_29136,N_27687,N_27180);
nor U29137 (N_29137,N_28332,N_27380);
or U29138 (N_29138,N_27196,N_27237);
or U29139 (N_29139,N_27567,N_27584);
and U29140 (N_29140,N_28053,N_28302);
and U29141 (N_29141,N_27721,N_27664);
nor U29142 (N_29142,N_27751,N_27857);
nor U29143 (N_29143,N_27525,N_27871);
nor U29144 (N_29144,N_27760,N_27780);
xor U29145 (N_29145,N_27215,N_27296);
nor U29146 (N_29146,N_27651,N_27761);
nand U29147 (N_29147,N_27200,N_27234);
nor U29148 (N_29148,N_27050,N_27639);
or U29149 (N_29149,N_28010,N_27710);
or U29150 (N_29150,N_27848,N_27762);
xnor U29151 (N_29151,N_27553,N_27015);
or U29152 (N_29152,N_28321,N_27926);
nor U29153 (N_29153,N_28049,N_27198);
or U29154 (N_29154,N_27275,N_27028);
or U29155 (N_29155,N_27494,N_27001);
nor U29156 (N_29156,N_28317,N_27524);
or U29157 (N_29157,N_28118,N_27154);
or U29158 (N_29158,N_27605,N_27405);
and U29159 (N_29159,N_27075,N_27909);
xor U29160 (N_29160,N_27880,N_27273);
and U29161 (N_29161,N_27064,N_27201);
and U29162 (N_29162,N_27395,N_27591);
or U29163 (N_29163,N_27419,N_27412);
nand U29164 (N_29164,N_27656,N_28467);
nor U29165 (N_29165,N_28330,N_27480);
xnor U29166 (N_29166,N_28342,N_27002);
xor U29167 (N_29167,N_27467,N_27774);
nand U29168 (N_29168,N_27385,N_27647);
nand U29169 (N_29169,N_28012,N_27282);
xnor U29170 (N_29170,N_27807,N_27240);
nor U29171 (N_29171,N_27940,N_27264);
or U29172 (N_29172,N_28380,N_28401);
and U29173 (N_29173,N_27303,N_27331);
nor U29174 (N_29174,N_28407,N_27637);
and U29175 (N_29175,N_27406,N_27310);
nand U29176 (N_29176,N_28443,N_28345);
xnor U29177 (N_29177,N_27367,N_27988);
and U29178 (N_29178,N_27090,N_27333);
xnor U29179 (N_29179,N_27096,N_27381);
or U29180 (N_29180,N_27199,N_27018);
nand U29181 (N_29181,N_27851,N_27998);
or U29182 (N_29182,N_28423,N_28497);
or U29183 (N_29183,N_28347,N_27482);
xor U29184 (N_29184,N_27635,N_28229);
and U29185 (N_29185,N_27628,N_28372);
and U29186 (N_29186,N_27565,N_27092);
nor U29187 (N_29187,N_28115,N_27490);
nand U29188 (N_29188,N_27868,N_27636);
nand U29189 (N_29189,N_27836,N_27100);
xor U29190 (N_29190,N_27587,N_27276);
nor U29191 (N_29191,N_27625,N_27581);
or U29192 (N_29192,N_27702,N_27238);
or U29193 (N_29193,N_27771,N_27464);
or U29194 (N_29194,N_27101,N_27041);
nand U29195 (N_29195,N_27043,N_28379);
nor U29196 (N_29196,N_27891,N_28058);
or U29197 (N_29197,N_27478,N_28197);
nand U29198 (N_29198,N_27299,N_27750);
nor U29199 (N_29199,N_27586,N_28490);
nand U29200 (N_29200,N_27602,N_27129);
and U29201 (N_29201,N_27861,N_28207);
xnor U29202 (N_29202,N_27905,N_27990);
nor U29203 (N_29203,N_27068,N_27777);
or U29204 (N_29204,N_27160,N_27548);
xnor U29205 (N_29205,N_28389,N_27846);
nand U29206 (N_29206,N_28026,N_28476);
nand U29207 (N_29207,N_28114,N_27074);
nand U29208 (N_29208,N_28202,N_27470);
and U29209 (N_29209,N_27549,N_27654);
nor U29210 (N_29210,N_27253,N_27313);
nand U29211 (N_29211,N_27970,N_27305);
nor U29212 (N_29212,N_28282,N_28307);
or U29213 (N_29213,N_27996,N_27558);
xor U29214 (N_29214,N_27270,N_27633);
and U29215 (N_29215,N_28212,N_27080);
or U29216 (N_29216,N_27547,N_27707);
and U29217 (N_29217,N_27948,N_28107);
nand U29218 (N_29218,N_27178,N_27195);
xnor U29219 (N_29219,N_27977,N_27258);
or U29220 (N_29220,N_27929,N_28222);
nor U29221 (N_29221,N_27062,N_27465);
or U29222 (N_29222,N_27550,N_27985);
nand U29223 (N_29223,N_27739,N_28044);
xnor U29224 (N_29224,N_27629,N_27814);
nor U29225 (N_29225,N_27193,N_27364);
and U29226 (N_29226,N_27262,N_27682);
nor U29227 (N_29227,N_27994,N_27916);
nand U29228 (N_29228,N_28175,N_27613);
or U29229 (N_29229,N_28093,N_27045);
nor U29230 (N_29230,N_27838,N_28496);
nand U29231 (N_29231,N_28416,N_27044);
and U29232 (N_29232,N_28140,N_28057);
nand U29233 (N_29233,N_27697,N_28030);
xor U29234 (N_29234,N_28106,N_28346);
nor U29235 (N_29235,N_27496,N_27911);
nand U29236 (N_29236,N_27830,N_28198);
xnor U29237 (N_29237,N_27428,N_28109);
nor U29238 (N_29238,N_27889,N_28344);
nand U29239 (N_29239,N_27340,N_28100);
or U29240 (N_29240,N_27789,N_27803);
xor U29241 (N_29241,N_27537,N_27755);
xnor U29242 (N_29242,N_27472,N_28032);
and U29243 (N_29243,N_27420,N_27667);
and U29244 (N_29244,N_28160,N_28047);
and U29245 (N_29245,N_27425,N_27119);
xor U29246 (N_29246,N_28325,N_27794);
or U29247 (N_29247,N_27704,N_27391);
and U29248 (N_29248,N_27617,N_27801);
nand U29249 (N_29249,N_28256,N_27255);
nand U29250 (N_29250,N_28459,N_27165);
nand U29251 (N_29251,N_27279,N_28114);
and U29252 (N_29252,N_27552,N_27342);
and U29253 (N_29253,N_27581,N_27401);
nor U29254 (N_29254,N_28425,N_27818);
nor U29255 (N_29255,N_27228,N_27734);
or U29256 (N_29256,N_27650,N_27061);
nor U29257 (N_29257,N_28465,N_27229);
and U29258 (N_29258,N_28022,N_28491);
nand U29259 (N_29259,N_27995,N_27005);
nand U29260 (N_29260,N_27187,N_28387);
nor U29261 (N_29261,N_28060,N_27016);
or U29262 (N_29262,N_28339,N_28133);
and U29263 (N_29263,N_27695,N_27593);
xnor U29264 (N_29264,N_28107,N_27851);
xnor U29265 (N_29265,N_28277,N_28327);
nor U29266 (N_29266,N_28056,N_27518);
and U29267 (N_29267,N_27718,N_28310);
nor U29268 (N_29268,N_27386,N_27832);
or U29269 (N_29269,N_27188,N_28365);
and U29270 (N_29270,N_27926,N_27663);
nor U29271 (N_29271,N_27207,N_28036);
nor U29272 (N_29272,N_27138,N_28360);
nor U29273 (N_29273,N_28266,N_27442);
xnor U29274 (N_29274,N_27668,N_27435);
or U29275 (N_29275,N_27348,N_28007);
nor U29276 (N_29276,N_28436,N_28238);
nor U29277 (N_29277,N_27114,N_28407);
nand U29278 (N_29278,N_27090,N_27457);
or U29279 (N_29279,N_27363,N_27476);
and U29280 (N_29280,N_27577,N_27764);
nor U29281 (N_29281,N_27044,N_27518);
xor U29282 (N_29282,N_27677,N_27629);
nand U29283 (N_29283,N_27934,N_27632);
nand U29284 (N_29284,N_27811,N_27779);
nand U29285 (N_29285,N_28165,N_27981);
nand U29286 (N_29286,N_27749,N_27100);
xnor U29287 (N_29287,N_27590,N_27395);
xor U29288 (N_29288,N_27569,N_27500);
nand U29289 (N_29289,N_27445,N_27402);
nand U29290 (N_29290,N_27054,N_27142);
and U29291 (N_29291,N_27481,N_27574);
nor U29292 (N_29292,N_27048,N_27152);
xor U29293 (N_29293,N_27130,N_27946);
or U29294 (N_29294,N_27067,N_27738);
nand U29295 (N_29295,N_27307,N_28315);
nand U29296 (N_29296,N_27413,N_28455);
and U29297 (N_29297,N_27954,N_27118);
nor U29298 (N_29298,N_27614,N_27218);
nor U29299 (N_29299,N_28018,N_27749);
nor U29300 (N_29300,N_27350,N_27125);
and U29301 (N_29301,N_27563,N_27660);
nor U29302 (N_29302,N_27539,N_27767);
nand U29303 (N_29303,N_27497,N_27194);
nand U29304 (N_29304,N_27923,N_27928);
xnor U29305 (N_29305,N_27435,N_28130);
or U29306 (N_29306,N_28264,N_27015);
xor U29307 (N_29307,N_28264,N_27369);
nor U29308 (N_29308,N_27752,N_28329);
nand U29309 (N_29309,N_27191,N_27420);
nor U29310 (N_29310,N_28252,N_27084);
or U29311 (N_29311,N_27779,N_27487);
nand U29312 (N_29312,N_27883,N_27044);
and U29313 (N_29313,N_27784,N_27147);
nor U29314 (N_29314,N_27081,N_28319);
and U29315 (N_29315,N_27291,N_27343);
nor U29316 (N_29316,N_27846,N_28165);
and U29317 (N_29317,N_27704,N_27730);
and U29318 (N_29318,N_28184,N_28244);
and U29319 (N_29319,N_28273,N_28033);
nand U29320 (N_29320,N_28246,N_27619);
and U29321 (N_29321,N_28163,N_27583);
xor U29322 (N_29322,N_27434,N_27436);
or U29323 (N_29323,N_27571,N_27709);
and U29324 (N_29324,N_27969,N_28177);
and U29325 (N_29325,N_27874,N_27610);
xnor U29326 (N_29326,N_27968,N_27185);
nor U29327 (N_29327,N_27800,N_27977);
nand U29328 (N_29328,N_27100,N_28233);
or U29329 (N_29329,N_28402,N_28016);
nor U29330 (N_29330,N_27301,N_27363);
nor U29331 (N_29331,N_28082,N_28110);
nand U29332 (N_29332,N_28274,N_27137);
or U29333 (N_29333,N_27198,N_27669);
nand U29334 (N_29334,N_27125,N_28487);
or U29335 (N_29335,N_27788,N_27520);
or U29336 (N_29336,N_27622,N_28392);
and U29337 (N_29337,N_27807,N_28205);
and U29338 (N_29338,N_28266,N_27559);
nor U29339 (N_29339,N_27471,N_27150);
xor U29340 (N_29340,N_27012,N_28095);
or U29341 (N_29341,N_27895,N_27740);
nand U29342 (N_29342,N_27633,N_27252);
and U29343 (N_29343,N_27542,N_27568);
xor U29344 (N_29344,N_27247,N_28003);
nand U29345 (N_29345,N_27189,N_27384);
and U29346 (N_29346,N_27932,N_28425);
nor U29347 (N_29347,N_28441,N_27167);
and U29348 (N_29348,N_27256,N_27328);
xor U29349 (N_29349,N_28102,N_27816);
nand U29350 (N_29350,N_28309,N_27247);
or U29351 (N_29351,N_27503,N_27939);
nand U29352 (N_29352,N_28324,N_27159);
and U29353 (N_29353,N_27943,N_27242);
nor U29354 (N_29354,N_27123,N_27421);
or U29355 (N_29355,N_27861,N_27554);
nand U29356 (N_29356,N_28125,N_27477);
and U29357 (N_29357,N_28059,N_28194);
nor U29358 (N_29358,N_27168,N_27875);
xnor U29359 (N_29359,N_27738,N_27325);
nand U29360 (N_29360,N_28420,N_28296);
nor U29361 (N_29361,N_27712,N_28234);
nor U29362 (N_29362,N_27653,N_28028);
xor U29363 (N_29363,N_27670,N_27058);
xnor U29364 (N_29364,N_28430,N_27773);
nor U29365 (N_29365,N_27285,N_28094);
or U29366 (N_29366,N_27159,N_28294);
nand U29367 (N_29367,N_27609,N_28143);
or U29368 (N_29368,N_28125,N_27170);
xnor U29369 (N_29369,N_28232,N_28128);
nor U29370 (N_29370,N_27831,N_27670);
or U29371 (N_29371,N_27708,N_28450);
and U29372 (N_29372,N_28473,N_28215);
nor U29373 (N_29373,N_27561,N_27788);
nor U29374 (N_29374,N_28056,N_27848);
nor U29375 (N_29375,N_27653,N_28408);
nand U29376 (N_29376,N_27483,N_28131);
and U29377 (N_29377,N_27461,N_28185);
and U29378 (N_29378,N_27376,N_28225);
nor U29379 (N_29379,N_27235,N_28272);
or U29380 (N_29380,N_27994,N_27398);
nor U29381 (N_29381,N_28386,N_28258);
nand U29382 (N_29382,N_27560,N_27309);
and U29383 (N_29383,N_28148,N_27198);
xnor U29384 (N_29384,N_27626,N_28132);
and U29385 (N_29385,N_28429,N_27812);
and U29386 (N_29386,N_27568,N_28245);
nor U29387 (N_29387,N_27001,N_27277);
and U29388 (N_29388,N_27819,N_27707);
nand U29389 (N_29389,N_28308,N_27599);
nor U29390 (N_29390,N_28175,N_27053);
xnor U29391 (N_29391,N_27086,N_28404);
nor U29392 (N_29392,N_28419,N_27522);
or U29393 (N_29393,N_27919,N_27725);
nand U29394 (N_29394,N_28436,N_27670);
nand U29395 (N_29395,N_28386,N_27131);
nand U29396 (N_29396,N_27316,N_27354);
or U29397 (N_29397,N_27490,N_27618);
or U29398 (N_29398,N_27054,N_27560);
nand U29399 (N_29399,N_27024,N_27237);
xor U29400 (N_29400,N_28322,N_28414);
nor U29401 (N_29401,N_27035,N_27494);
xor U29402 (N_29402,N_27494,N_27865);
nor U29403 (N_29403,N_27297,N_27038);
and U29404 (N_29404,N_28390,N_27575);
and U29405 (N_29405,N_28288,N_27090);
nand U29406 (N_29406,N_27397,N_27038);
nand U29407 (N_29407,N_27651,N_28174);
and U29408 (N_29408,N_27820,N_28209);
xor U29409 (N_29409,N_27505,N_27786);
or U29410 (N_29410,N_27124,N_28056);
or U29411 (N_29411,N_27563,N_27645);
xnor U29412 (N_29412,N_28236,N_27388);
nor U29413 (N_29413,N_28473,N_28163);
and U29414 (N_29414,N_28388,N_28209);
xnor U29415 (N_29415,N_27118,N_27237);
or U29416 (N_29416,N_28199,N_28387);
nand U29417 (N_29417,N_27640,N_28097);
nor U29418 (N_29418,N_28363,N_27303);
nor U29419 (N_29419,N_27872,N_28319);
nor U29420 (N_29420,N_28433,N_27053);
xor U29421 (N_29421,N_27212,N_27364);
and U29422 (N_29422,N_28332,N_27906);
nor U29423 (N_29423,N_27953,N_27840);
nor U29424 (N_29424,N_27579,N_27709);
nor U29425 (N_29425,N_27504,N_27961);
or U29426 (N_29426,N_27198,N_28022);
and U29427 (N_29427,N_28037,N_28233);
and U29428 (N_29428,N_28384,N_27762);
xnor U29429 (N_29429,N_27520,N_28164);
xnor U29430 (N_29430,N_27463,N_27032);
nor U29431 (N_29431,N_27847,N_27815);
and U29432 (N_29432,N_27192,N_27694);
and U29433 (N_29433,N_28204,N_28487);
nor U29434 (N_29434,N_27332,N_27248);
xnor U29435 (N_29435,N_28310,N_28202);
or U29436 (N_29436,N_28229,N_27697);
or U29437 (N_29437,N_27546,N_28134);
xnor U29438 (N_29438,N_27914,N_27626);
and U29439 (N_29439,N_28376,N_27745);
nor U29440 (N_29440,N_27828,N_27498);
nor U29441 (N_29441,N_27268,N_27219);
nand U29442 (N_29442,N_27812,N_27218);
nand U29443 (N_29443,N_27594,N_27461);
nand U29444 (N_29444,N_27237,N_27768);
or U29445 (N_29445,N_27292,N_27493);
xnor U29446 (N_29446,N_27550,N_27318);
nor U29447 (N_29447,N_28209,N_27201);
nor U29448 (N_29448,N_27400,N_27311);
nand U29449 (N_29449,N_27149,N_28229);
nor U29450 (N_29450,N_28132,N_27818);
nand U29451 (N_29451,N_27112,N_28194);
nor U29452 (N_29452,N_27825,N_27714);
and U29453 (N_29453,N_27967,N_27158);
nand U29454 (N_29454,N_28176,N_27107);
xnor U29455 (N_29455,N_28343,N_27608);
nor U29456 (N_29456,N_27812,N_27182);
and U29457 (N_29457,N_28405,N_27277);
and U29458 (N_29458,N_27599,N_27991);
and U29459 (N_29459,N_28335,N_28068);
or U29460 (N_29460,N_27000,N_27156);
or U29461 (N_29461,N_27347,N_28495);
nand U29462 (N_29462,N_27690,N_28044);
and U29463 (N_29463,N_28455,N_27551);
or U29464 (N_29464,N_27471,N_27217);
or U29465 (N_29465,N_27610,N_27648);
nor U29466 (N_29466,N_27426,N_28155);
nor U29467 (N_29467,N_27112,N_27795);
xor U29468 (N_29468,N_28066,N_27448);
or U29469 (N_29469,N_27196,N_27567);
and U29470 (N_29470,N_27761,N_28155);
nor U29471 (N_29471,N_28221,N_27249);
nand U29472 (N_29472,N_27060,N_27769);
xnor U29473 (N_29473,N_28346,N_27052);
xor U29474 (N_29474,N_27544,N_27580);
nor U29475 (N_29475,N_27862,N_28240);
nor U29476 (N_29476,N_27829,N_27293);
or U29477 (N_29477,N_27291,N_28207);
xor U29478 (N_29478,N_27687,N_27875);
xor U29479 (N_29479,N_27793,N_28248);
or U29480 (N_29480,N_27973,N_27204);
xnor U29481 (N_29481,N_28406,N_28125);
nor U29482 (N_29482,N_28451,N_27072);
and U29483 (N_29483,N_28206,N_27909);
nand U29484 (N_29484,N_27324,N_27883);
nor U29485 (N_29485,N_28267,N_27543);
or U29486 (N_29486,N_27633,N_28369);
nand U29487 (N_29487,N_27285,N_27664);
and U29488 (N_29488,N_27622,N_27707);
or U29489 (N_29489,N_27355,N_28277);
nor U29490 (N_29490,N_28487,N_27289);
or U29491 (N_29491,N_28368,N_27808);
xnor U29492 (N_29492,N_28383,N_27397);
or U29493 (N_29493,N_27301,N_27190);
nand U29494 (N_29494,N_28385,N_28023);
xnor U29495 (N_29495,N_27437,N_27758);
and U29496 (N_29496,N_27298,N_27733);
nand U29497 (N_29497,N_27673,N_27003);
xnor U29498 (N_29498,N_27646,N_27368);
and U29499 (N_29499,N_27324,N_28349);
xnor U29500 (N_29500,N_27491,N_28127);
xnor U29501 (N_29501,N_28044,N_27990);
nand U29502 (N_29502,N_28469,N_27364);
and U29503 (N_29503,N_28332,N_27537);
or U29504 (N_29504,N_28164,N_27861);
xor U29505 (N_29505,N_28403,N_27835);
nand U29506 (N_29506,N_28004,N_27249);
nand U29507 (N_29507,N_28278,N_27985);
or U29508 (N_29508,N_27314,N_27372);
xnor U29509 (N_29509,N_27986,N_27100);
and U29510 (N_29510,N_27128,N_28077);
or U29511 (N_29511,N_27841,N_27729);
or U29512 (N_29512,N_27144,N_28076);
and U29513 (N_29513,N_27821,N_27355);
nand U29514 (N_29514,N_28381,N_27048);
xor U29515 (N_29515,N_27813,N_28365);
nor U29516 (N_29516,N_28332,N_27957);
nand U29517 (N_29517,N_28394,N_28280);
and U29518 (N_29518,N_27027,N_28347);
nand U29519 (N_29519,N_28414,N_27643);
and U29520 (N_29520,N_27837,N_27162);
nand U29521 (N_29521,N_27834,N_27791);
nand U29522 (N_29522,N_27269,N_27002);
nand U29523 (N_29523,N_28490,N_27762);
nor U29524 (N_29524,N_27590,N_27944);
nand U29525 (N_29525,N_27292,N_28102);
and U29526 (N_29526,N_28484,N_27571);
or U29527 (N_29527,N_28270,N_27693);
and U29528 (N_29528,N_27105,N_27477);
or U29529 (N_29529,N_27845,N_28123);
nand U29530 (N_29530,N_27202,N_27927);
and U29531 (N_29531,N_28232,N_27494);
nand U29532 (N_29532,N_27375,N_27767);
and U29533 (N_29533,N_28070,N_27904);
xor U29534 (N_29534,N_27884,N_27889);
or U29535 (N_29535,N_28166,N_27243);
or U29536 (N_29536,N_27391,N_28172);
and U29537 (N_29537,N_27232,N_28410);
xor U29538 (N_29538,N_27026,N_27875);
nor U29539 (N_29539,N_27866,N_27439);
nor U29540 (N_29540,N_27665,N_27211);
nand U29541 (N_29541,N_28312,N_27783);
nor U29542 (N_29542,N_28217,N_27982);
nand U29543 (N_29543,N_28190,N_27952);
and U29544 (N_29544,N_28341,N_27009);
or U29545 (N_29545,N_28386,N_27460);
or U29546 (N_29546,N_28333,N_27614);
and U29547 (N_29547,N_27000,N_28328);
and U29548 (N_29548,N_27687,N_27803);
or U29549 (N_29549,N_28386,N_28446);
or U29550 (N_29550,N_28072,N_28242);
nand U29551 (N_29551,N_28305,N_27389);
or U29552 (N_29552,N_28093,N_27576);
and U29553 (N_29553,N_27159,N_28136);
xnor U29554 (N_29554,N_28235,N_27594);
nor U29555 (N_29555,N_27227,N_28439);
or U29556 (N_29556,N_28257,N_28200);
nor U29557 (N_29557,N_27922,N_27484);
or U29558 (N_29558,N_27177,N_28269);
xnor U29559 (N_29559,N_27188,N_27717);
nand U29560 (N_29560,N_28284,N_27479);
xnor U29561 (N_29561,N_27355,N_27128);
xnor U29562 (N_29562,N_27206,N_27353);
or U29563 (N_29563,N_27165,N_27945);
nor U29564 (N_29564,N_27528,N_28463);
xor U29565 (N_29565,N_28172,N_27373);
or U29566 (N_29566,N_28040,N_27313);
xor U29567 (N_29567,N_27926,N_28037);
or U29568 (N_29568,N_27095,N_27473);
or U29569 (N_29569,N_28039,N_27120);
or U29570 (N_29570,N_28436,N_28312);
or U29571 (N_29571,N_27534,N_28059);
nand U29572 (N_29572,N_28302,N_27578);
or U29573 (N_29573,N_27618,N_27271);
and U29574 (N_29574,N_27349,N_27436);
nor U29575 (N_29575,N_27538,N_28189);
xor U29576 (N_29576,N_28153,N_27271);
nand U29577 (N_29577,N_27969,N_27946);
nand U29578 (N_29578,N_27371,N_28131);
nor U29579 (N_29579,N_28131,N_28354);
and U29580 (N_29580,N_27434,N_27781);
nor U29581 (N_29581,N_27017,N_28494);
and U29582 (N_29582,N_28190,N_27034);
xnor U29583 (N_29583,N_28005,N_27244);
xnor U29584 (N_29584,N_28051,N_27876);
nor U29585 (N_29585,N_27412,N_28326);
xnor U29586 (N_29586,N_27592,N_27444);
nor U29587 (N_29587,N_27638,N_27837);
nor U29588 (N_29588,N_27010,N_28273);
nand U29589 (N_29589,N_27387,N_27461);
or U29590 (N_29590,N_27427,N_28363);
or U29591 (N_29591,N_27664,N_27562);
xor U29592 (N_29592,N_28212,N_27798);
or U29593 (N_29593,N_27847,N_27192);
xor U29594 (N_29594,N_28393,N_27926);
nor U29595 (N_29595,N_27358,N_27734);
xnor U29596 (N_29596,N_28057,N_27418);
nand U29597 (N_29597,N_27250,N_27261);
nand U29598 (N_29598,N_27272,N_27197);
and U29599 (N_29599,N_27402,N_27658);
nor U29600 (N_29600,N_27244,N_27884);
or U29601 (N_29601,N_27326,N_27852);
nand U29602 (N_29602,N_28485,N_27931);
and U29603 (N_29603,N_27985,N_28201);
nor U29604 (N_29604,N_28237,N_27204);
and U29605 (N_29605,N_27650,N_27903);
nand U29606 (N_29606,N_27247,N_27536);
and U29607 (N_29607,N_27808,N_27059);
or U29608 (N_29608,N_27748,N_27073);
or U29609 (N_29609,N_27306,N_28079);
or U29610 (N_29610,N_28491,N_27450);
nor U29611 (N_29611,N_27367,N_28038);
and U29612 (N_29612,N_28328,N_27714);
nor U29613 (N_29613,N_27590,N_27143);
nand U29614 (N_29614,N_27128,N_28053);
or U29615 (N_29615,N_27647,N_27869);
or U29616 (N_29616,N_27095,N_27335);
xor U29617 (N_29617,N_27149,N_27006);
or U29618 (N_29618,N_27091,N_27313);
or U29619 (N_29619,N_27929,N_27718);
or U29620 (N_29620,N_27252,N_27976);
nor U29621 (N_29621,N_28097,N_28203);
and U29622 (N_29622,N_27957,N_28082);
nand U29623 (N_29623,N_27475,N_27196);
nand U29624 (N_29624,N_27528,N_28484);
and U29625 (N_29625,N_27861,N_27571);
nor U29626 (N_29626,N_28490,N_27426);
nor U29627 (N_29627,N_27995,N_27562);
xnor U29628 (N_29628,N_27235,N_28233);
nand U29629 (N_29629,N_27644,N_27412);
xor U29630 (N_29630,N_28066,N_27621);
nand U29631 (N_29631,N_27804,N_28398);
and U29632 (N_29632,N_27569,N_27623);
and U29633 (N_29633,N_28404,N_28016);
nor U29634 (N_29634,N_28365,N_27956);
nor U29635 (N_29635,N_27586,N_27806);
nand U29636 (N_29636,N_28478,N_27610);
nand U29637 (N_29637,N_27697,N_28335);
xor U29638 (N_29638,N_27901,N_27045);
nand U29639 (N_29639,N_27875,N_27904);
or U29640 (N_29640,N_27839,N_28402);
or U29641 (N_29641,N_28266,N_27330);
and U29642 (N_29642,N_28271,N_28372);
or U29643 (N_29643,N_27774,N_27657);
nor U29644 (N_29644,N_27490,N_27464);
nand U29645 (N_29645,N_27979,N_27076);
nand U29646 (N_29646,N_27704,N_28340);
nor U29647 (N_29647,N_27074,N_27059);
or U29648 (N_29648,N_28006,N_27978);
xor U29649 (N_29649,N_28235,N_27523);
xnor U29650 (N_29650,N_28224,N_27269);
nand U29651 (N_29651,N_28166,N_27014);
or U29652 (N_29652,N_28321,N_27287);
xnor U29653 (N_29653,N_27427,N_27114);
nor U29654 (N_29654,N_27480,N_27753);
nor U29655 (N_29655,N_28384,N_27389);
or U29656 (N_29656,N_27402,N_28429);
or U29657 (N_29657,N_28084,N_27534);
or U29658 (N_29658,N_27870,N_28294);
or U29659 (N_29659,N_28419,N_27497);
nand U29660 (N_29660,N_27884,N_28143);
or U29661 (N_29661,N_27765,N_28135);
xor U29662 (N_29662,N_28019,N_27032);
and U29663 (N_29663,N_27139,N_27467);
xor U29664 (N_29664,N_28442,N_27752);
xnor U29665 (N_29665,N_27406,N_27963);
xor U29666 (N_29666,N_27414,N_28194);
and U29667 (N_29667,N_28120,N_27982);
nand U29668 (N_29668,N_27309,N_27340);
and U29669 (N_29669,N_27275,N_28396);
xor U29670 (N_29670,N_28071,N_27038);
nand U29671 (N_29671,N_27190,N_27468);
xor U29672 (N_29672,N_27853,N_28059);
xor U29673 (N_29673,N_28205,N_27680);
nor U29674 (N_29674,N_28292,N_27994);
xor U29675 (N_29675,N_28380,N_27498);
and U29676 (N_29676,N_28462,N_28107);
nor U29677 (N_29677,N_28131,N_28369);
or U29678 (N_29678,N_28008,N_27809);
nor U29679 (N_29679,N_27745,N_27776);
and U29680 (N_29680,N_27644,N_28229);
xor U29681 (N_29681,N_27844,N_27912);
xor U29682 (N_29682,N_28316,N_27493);
or U29683 (N_29683,N_27898,N_27829);
or U29684 (N_29684,N_27493,N_28410);
xnor U29685 (N_29685,N_27697,N_27645);
xnor U29686 (N_29686,N_27538,N_27402);
nor U29687 (N_29687,N_28296,N_27133);
or U29688 (N_29688,N_27727,N_28217);
or U29689 (N_29689,N_27114,N_27778);
or U29690 (N_29690,N_27418,N_28295);
and U29691 (N_29691,N_27816,N_28118);
or U29692 (N_29692,N_27176,N_28079);
and U29693 (N_29693,N_27779,N_27236);
and U29694 (N_29694,N_27575,N_28177);
nor U29695 (N_29695,N_27137,N_27379);
and U29696 (N_29696,N_27435,N_28206);
xnor U29697 (N_29697,N_28468,N_28352);
nand U29698 (N_29698,N_27031,N_28212);
xnor U29699 (N_29699,N_28132,N_27241);
or U29700 (N_29700,N_28282,N_27321);
xnor U29701 (N_29701,N_27086,N_27835);
or U29702 (N_29702,N_27062,N_27798);
nor U29703 (N_29703,N_27693,N_27491);
nand U29704 (N_29704,N_28059,N_27452);
or U29705 (N_29705,N_27437,N_28237);
nand U29706 (N_29706,N_28206,N_28363);
and U29707 (N_29707,N_27760,N_28128);
nor U29708 (N_29708,N_28369,N_28478);
or U29709 (N_29709,N_27120,N_27061);
and U29710 (N_29710,N_28465,N_27014);
or U29711 (N_29711,N_27466,N_28210);
or U29712 (N_29712,N_28152,N_28025);
and U29713 (N_29713,N_27063,N_28227);
nor U29714 (N_29714,N_27521,N_27676);
nand U29715 (N_29715,N_28447,N_28451);
nor U29716 (N_29716,N_27712,N_27090);
nor U29717 (N_29717,N_27450,N_27289);
nor U29718 (N_29718,N_28332,N_27614);
nand U29719 (N_29719,N_27893,N_27487);
nand U29720 (N_29720,N_27109,N_28042);
or U29721 (N_29721,N_28065,N_27352);
xnor U29722 (N_29722,N_28042,N_28347);
nor U29723 (N_29723,N_28017,N_27809);
xnor U29724 (N_29724,N_28347,N_27684);
nand U29725 (N_29725,N_27388,N_28334);
nand U29726 (N_29726,N_27276,N_28488);
nor U29727 (N_29727,N_27488,N_28046);
nor U29728 (N_29728,N_27379,N_27262);
xor U29729 (N_29729,N_28459,N_27674);
nor U29730 (N_29730,N_27140,N_27450);
or U29731 (N_29731,N_28151,N_28179);
nor U29732 (N_29732,N_28082,N_27395);
nor U29733 (N_29733,N_28281,N_27755);
nand U29734 (N_29734,N_27420,N_28289);
nor U29735 (N_29735,N_27630,N_27720);
nor U29736 (N_29736,N_27055,N_27969);
xnor U29737 (N_29737,N_27702,N_27289);
or U29738 (N_29738,N_28477,N_27795);
xor U29739 (N_29739,N_27666,N_28052);
nand U29740 (N_29740,N_27295,N_27631);
nor U29741 (N_29741,N_27783,N_27996);
nand U29742 (N_29742,N_27132,N_27945);
or U29743 (N_29743,N_28224,N_28312);
nor U29744 (N_29744,N_27234,N_27117);
xor U29745 (N_29745,N_28137,N_27192);
nand U29746 (N_29746,N_28273,N_27319);
and U29747 (N_29747,N_28067,N_27588);
nand U29748 (N_29748,N_28053,N_27744);
and U29749 (N_29749,N_28281,N_28390);
nand U29750 (N_29750,N_28308,N_27092);
or U29751 (N_29751,N_27921,N_27576);
and U29752 (N_29752,N_27535,N_28229);
or U29753 (N_29753,N_28414,N_27853);
nand U29754 (N_29754,N_27420,N_27997);
or U29755 (N_29755,N_27456,N_27098);
xor U29756 (N_29756,N_27321,N_27436);
and U29757 (N_29757,N_28298,N_27334);
or U29758 (N_29758,N_27300,N_28319);
or U29759 (N_29759,N_27780,N_27248);
and U29760 (N_29760,N_28447,N_27792);
nand U29761 (N_29761,N_27828,N_27051);
or U29762 (N_29762,N_27448,N_28100);
nor U29763 (N_29763,N_27249,N_27657);
nor U29764 (N_29764,N_27671,N_27526);
nor U29765 (N_29765,N_27874,N_27466);
nor U29766 (N_29766,N_27745,N_27598);
or U29767 (N_29767,N_27560,N_28349);
xor U29768 (N_29768,N_27065,N_27412);
and U29769 (N_29769,N_27196,N_27303);
nand U29770 (N_29770,N_27238,N_27294);
xnor U29771 (N_29771,N_27395,N_27073);
nand U29772 (N_29772,N_28306,N_28132);
or U29773 (N_29773,N_27476,N_28396);
or U29774 (N_29774,N_27381,N_27104);
nor U29775 (N_29775,N_28229,N_27915);
nand U29776 (N_29776,N_27542,N_27657);
or U29777 (N_29777,N_28446,N_28071);
xor U29778 (N_29778,N_27532,N_27290);
or U29779 (N_29779,N_27066,N_27734);
and U29780 (N_29780,N_27927,N_28035);
xnor U29781 (N_29781,N_27583,N_28266);
or U29782 (N_29782,N_27433,N_27795);
or U29783 (N_29783,N_28260,N_27144);
xnor U29784 (N_29784,N_27318,N_27448);
xnor U29785 (N_29785,N_28252,N_27429);
nand U29786 (N_29786,N_27525,N_27896);
and U29787 (N_29787,N_27148,N_28125);
xnor U29788 (N_29788,N_27687,N_27588);
nand U29789 (N_29789,N_27991,N_27629);
and U29790 (N_29790,N_27907,N_27215);
nor U29791 (N_29791,N_27265,N_27123);
nor U29792 (N_29792,N_27396,N_28205);
nand U29793 (N_29793,N_27478,N_27361);
or U29794 (N_29794,N_27628,N_27475);
or U29795 (N_29795,N_27279,N_27925);
or U29796 (N_29796,N_28305,N_27785);
nor U29797 (N_29797,N_27805,N_28439);
xnor U29798 (N_29798,N_27418,N_27950);
or U29799 (N_29799,N_28390,N_27988);
nor U29800 (N_29800,N_27030,N_27589);
xnor U29801 (N_29801,N_27529,N_27503);
nor U29802 (N_29802,N_27615,N_28431);
nor U29803 (N_29803,N_28407,N_27698);
or U29804 (N_29804,N_27382,N_28132);
or U29805 (N_29805,N_28402,N_28356);
xor U29806 (N_29806,N_27688,N_27160);
nand U29807 (N_29807,N_28138,N_27866);
and U29808 (N_29808,N_28215,N_27116);
or U29809 (N_29809,N_28127,N_28293);
nor U29810 (N_29810,N_27129,N_27547);
nor U29811 (N_29811,N_28367,N_27900);
xor U29812 (N_29812,N_27339,N_27180);
xnor U29813 (N_29813,N_28404,N_27704);
nor U29814 (N_29814,N_27523,N_28468);
xnor U29815 (N_29815,N_28154,N_28468);
nand U29816 (N_29816,N_27596,N_28270);
and U29817 (N_29817,N_28208,N_28289);
xnor U29818 (N_29818,N_27762,N_27730);
xnor U29819 (N_29819,N_27201,N_27683);
nor U29820 (N_29820,N_27868,N_27702);
or U29821 (N_29821,N_28031,N_27416);
and U29822 (N_29822,N_28348,N_28002);
nor U29823 (N_29823,N_28481,N_28113);
nand U29824 (N_29824,N_27614,N_27148);
xor U29825 (N_29825,N_27450,N_28018);
and U29826 (N_29826,N_28021,N_27112);
nand U29827 (N_29827,N_28037,N_27611);
nor U29828 (N_29828,N_27175,N_28478);
nand U29829 (N_29829,N_28446,N_28445);
or U29830 (N_29830,N_28231,N_27707);
nand U29831 (N_29831,N_27819,N_27333);
and U29832 (N_29832,N_28334,N_27795);
or U29833 (N_29833,N_28197,N_27632);
xor U29834 (N_29834,N_28114,N_27753);
nand U29835 (N_29835,N_27187,N_27080);
nand U29836 (N_29836,N_27992,N_27580);
nand U29837 (N_29837,N_28415,N_27169);
xor U29838 (N_29838,N_27630,N_27356);
nand U29839 (N_29839,N_27778,N_28269);
nor U29840 (N_29840,N_28266,N_27232);
nor U29841 (N_29841,N_27946,N_27952);
nor U29842 (N_29842,N_28326,N_27384);
nor U29843 (N_29843,N_27921,N_27093);
nor U29844 (N_29844,N_27013,N_27665);
xor U29845 (N_29845,N_27714,N_27268);
nor U29846 (N_29846,N_28045,N_27429);
xor U29847 (N_29847,N_27377,N_27674);
xnor U29848 (N_29848,N_27115,N_27205);
nand U29849 (N_29849,N_27986,N_28293);
nand U29850 (N_29850,N_27227,N_27515);
or U29851 (N_29851,N_28381,N_27087);
or U29852 (N_29852,N_27758,N_27290);
and U29853 (N_29853,N_27421,N_27278);
or U29854 (N_29854,N_28012,N_27986);
or U29855 (N_29855,N_28484,N_28462);
and U29856 (N_29856,N_27910,N_27813);
and U29857 (N_29857,N_28379,N_27388);
xnor U29858 (N_29858,N_27383,N_27387);
nand U29859 (N_29859,N_27825,N_27907);
and U29860 (N_29860,N_28119,N_27936);
and U29861 (N_29861,N_28358,N_27967);
or U29862 (N_29862,N_27393,N_28459);
and U29863 (N_29863,N_27571,N_28039);
nor U29864 (N_29864,N_27838,N_27788);
xor U29865 (N_29865,N_27621,N_27714);
nand U29866 (N_29866,N_27084,N_27173);
nand U29867 (N_29867,N_27152,N_27087);
and U29868 (N_29868,N_27114,N_28360);
nor U29869 (N_29869,N_27581,N_27990);
and U29870 (N_29870,N_27015,N_28351);
or U29871 (N_29871,N_27688,N_27578);
nand U29872 (N_29872,N_27136,N_27073);
or U29873 (N_29873,N_27453,N_27858);
and U29874 (N_29874,N_27649,N_27306);
or U29875 (N_29875,N_28131,N_27143);
and U29876 (N_29876,N_27873,N_27205);
nor U29877 (N_29877,N_27578,N_28415);
nand U29878 (N_29878,N_28418,N_27103);
nand U29879 (N_29879,N_28063,N_27538);
xor U29880 (N_29880,N_28027,N_27379);
nand U29881 (N_29881,N_28370,N_27612);
xor U29882 (N_29882,N_27533,N_27511);
and U29883 (N_29883,N_27277,N_28062);
or U29884 (N_29884,N_27634,N_27837);
or U29885 (N_29885,N_27369,N_28331);
nand U29886 (N_29886,N_27706,N_27508);
and U29887 (N_29887,N_28413,N_28375);
nand U29888 (N_29888,N_28248,N_27385);
nand U29889 (N_29889,N_28044,N_28372);
and U29890 (N_29890,N_27715,N_27666);
nor U29891 (N_29891,N_27110,N_28448);
or U29892 (N_29892,N_27554,N_27353);
and U29893 (N_29893,N_28096,N_28031);
nor U29894 (N_29894,N_27185,N_27604);
nand U29895 (N_29895,N_28330,N_28303);
or U29896 (N_29896,N_28321,N_27340);
nand U29897 (N_29897,N_27132,N_28414);
nor U29898 (N_29898,N_28187,N_27719);
xor U29899 (N_29899,N_28004,N_28252);
nor U29900 (N_29900,N_27561,N_27506);
nand U29901 (N_29901,N_27386,N_27722);
and U29902 (N_29902,N_27456,N_27208);
nand U29903 (N_29903,N_27498,N_27597);
or U29904 (N_29904,N_27147,N_27129);
and U29905 (N_29905,N_28059,N_28219);
xor U29906 (N_29906,N_27021,N_27987);
and U29907 (N_29907,N_27468,N_27011);
and U29908 (N_29908,N_27580,N_27978);
and U29909 (N_29909,N_27865,N_27847);
xor U29910 (N_29910,N_27884,N_28006);
nand U29911 (N_29911,N_28152,N_28130);
nor U29912 (N_29912,N_27484,N_27067);
nor U29913 (N_29913,N_28293,N_28401);
nand U29914 (N_29914,N_27726,N_28015);
nor U29915 (N_29915,N_27298,N_27222);
and U29916 (N_29916,N_28113,N_27132);
xor U29917 (N_29917,N_27426,N_27766);
xnor U29918 (N_29918,N_27032,N_27153);
nor U29919 (N_29919,N_28010,N_27738);
nor U29920 (N_29920,N_27642,N_27982);
xor U29921 (N_29921,N_28357,N_27529);
and U29922 (N_29922,N_27300,N_27103);
and U29923 (N_29923,N_28431,N_27105);
xor U29924 (N_29924,N_27546,N_28033);
nand U29925 (N_29925,N_27119,N_27571);
nor U29926 (N_29926,N_28417,N_27336);
nand U29927 (N_29927,N_27809,N_27577);
nor U29928 (N_29928,N_27613,N_28444);
nand U29929 (N_29929,N_27245,N_27517);
or U29930 (N_29930,N_27156,N_28447);
xor U29931 (N_29931,N_28019,N_27728);
or U29932 (N_29932,N_27159,N_28201);
or U29933 (N_29933,N_28418,N_27447);
xnor U29934 (N_29934,N_27973,N_27893);
xnor U29935 (N_29935,N_27522,N_27666);
xnor U29936 (N_29936,N_27559,N_27420);
and U29937 (N_29937,N_27204,N_28172);
nor U29938 (N_29938,N_27791,N_28073);
and U29939 (N_29939,N_27293,N_27282);
and U29940 (N_29940,N_27281,N_27001);
nor U29941 (N_29941,N_27400,N_28342);
nor U29942 (N_29942,N_28163,N_27412);
nor U29943 (N_29943,N_27050,N_28052);
and U29944 (N_29944,N_27423,N_27897);
nor U29945 (N_29945,N_27603,N_27795);
nand U29946 (N_29946,N_27585,N_28476);
nor U29947 (N_29947,N_27238,N_27131);
xnor U29948 (N_29948,N_27983,N_28248);
or U29949 (N_29949,N_27916,N_28358);
nor U29950 (N_29950,N_27164,N_27308);
nand U29951 (N_29951,N_27043,N_27391);
nand U29952 (N_29952,N_27139,N_28480);
nor U29953 (N_29953,N_27608,N_27239);
nor U29954 (N_29954,N_28310,N_27765);
and U29955 (N_29955,N_27574,N_27684);
or U29956 (N_29956,N_27533,N_27318);
and U29957 (N_29957,N_27194,N_27027);
xnor U29958 (N_29958,N_28338,N_28369);
and U29959 (N_29959,N_27938,N_28038);
and U29960 (N_29960,N_28425,N_27550);
nor U29961 (N_29961,N_27569,N_27536);
nand U29962 (N_29962,N_27040,N_28062);
or U29963 (N_29963,N_27356,N_27026);
xor U29964 (N_29964,N_27734,N_28088);
xnor U29965 (N_29965,N_28084,N_28338);
nor U29966 (N_29966,N_27812,N_28201);
nor U29967 (N_29967,N_27762,N_27075);
xnor U29968 (N_29968,N_28205,N_27728);
and U29969 (N_29969,N_27690,N_28495);
nor U29970 (N_29970,N_28479,N_28279);
xnor U29971 (N_29971,N_27260,N_27113);
and U29972 (N_29972,N_27364,N_27339);
and U29973 (N_29973,N_27181,N_27658);
xnor U29974 (N_29974,N_27873,N_28262);
xnor U29975 (N_29975,N_27717,N_28354);
and U29976 (N_29976,N_27653,N_27886);
nand U29977 (N_29977,N_28009,N_28434);
and U29978 (N_29978,N_27450,N_28029);
xnor U29979 (N_29979,N_28451,N_27059);
xnor U29980 (N_29980,N_27945,N_27335);
nor U29981 (N_29981,N_28286,N_27221);
and U29982 (N_29982,N_27971,N_27758);
nor U29983 (N_29983,N_27625,N_27769);
or U29984 (N_29984,N_28118,N_27033);
xnor U29985 (N_29985,N_28276,N_27613);
or U29986 (N_29986,N_28109,N_27411);
and U29987 (N_29987,N_28152,N_28047);
xor U29988 (N_29988,N_27106,N_27103);
nor U29989 (N_29989,N_28346,N_27345);
or U29990 (N_29990,N_28354,N_28037);
and U29991 (N_29991,N_28475,N_28053);
nand U29992 (N_29992,N_27950,N_28203);
nor U29993 (N_29993,N_27962,N_28382);
nand U29994 (N_29994,N_27300,N_28301);
and U29995 (N_29995,N_28441,N_27528);
or U29996 (N_29996,N_27423,N_27047);
xor U29997 (N_29997,N_28256,N_27831);
nand U29998 (N_29998,N_27892,N_27986);
and U29999 (N_29999,N_28249,N_28143);
xnor UO_0 (O_0,N_29212,N_29893);
nand UO_1 (O_1,N_29736,N_29780);
or UO_2 (O_2,N_29841,N_29294);
nor UO_3 (O_3,N_28626,N_29503);
or UO_4 (O_4,N_29013,N_28630);
and UO_5 (O_5,N_28503,N_28907);
nor UO_6 (O_6,N_29650,N_28903);
xor UO_7 (O_7,N_28874,N_29050);
nor UO_8 (O_8,N_29399,N_28863);
and UO_9 (O_9,N_28536,N_28752);
xnor UO_10 (O_10,N_29104,N_28582);
and UO_11 (O_11,N_29626,N_29540);
xor UO_12 (O_12,N_28706,N_29533);
and UO_13 (O_13,N_29357,N_29710);
and UO_14 (O_14,N_29960,N_29846);
and UO_15 (O_15,N_28543,N_28914);
nor UO_16 (O_16,N_29924,N_29674);
nor UO_17 (O_17,N_29567,N_29191);
nand UO_18 (O_18,N_29279,N_28856);
xor UO_19 (O_19,N_28820,N_29694);
nor UO_20 (O_20,N_29224,N_29946);
and UO_21 (O_21,N_28773,N_28768);
xor UO_22 (O_22,N_29782,N_29255);
nand UO_23 (O_23,N_29098,N_29119);
xnor UO_24 (O_24,N_29428,N_29022);
and UO_25 (O_25,N_28921,N_29851);
nor UO_26 (O_26,N_29882,N_29322);
or UO_27 (O_27,N_29200,N_29602);
or UO_28 (O_28,N_29732,N_29744);
or UO_29 (O_29,N_29048,N_29395);
nor UO_30 (O_30,N_29547,N_29296);
nand UO_31 (O_31,N_28806,N_29149);
nor UO_32 (O_32,N_29947,N_28590);
or UO_33 (O_33,N_29252,N_28682);
or UO_34 (O_34,N_29394,N_28584);
or UO_35 (O_35,N_29508,N_28559);
or UO_36 (O_36,N_28850,N_29730);
nand UO_37 (O_37,N_29570,N_28915);
and UO_38 (O_38,N_29774,N_29727);
and UO_39 (O_39,N_28946,N_29617);
xor UO_40 (O_40,N_29790,N_28765);
and UO_41 (O_41,N_28614,N_29784);
xor UO_42 (O_42,N_28848,N_29998);
xnor UO_43 (O_43,N_29226,N_29091);
or UO_44 (O_44,N_28668,N_29776);
nand UO_45 (O_45,N_29747,N_29138);
and UO_46 (O_46,N_28884,N_29114);
and UO_47 (O_47,N_28818,N_28955);
or UO_48 (O_48,N_29970,N_29686);
and UO_49 (O_49,N_29576,N_29654);
or UO_50 (O_50,N_28574,N_29139);
nor UO_51 (O_51,N_29342,N_29810);
and UO_52 (O_52,N_29573,N_29618);
xnor UO_53 (O_53,N_28697,N_28568);
nor UO_54 (O_54,N_28941,N_29315);
nand UO_55 (O_55,N_29684,N_29598);
xor UO_56 (O_56,N_29007,N_28645);
and UO_57 (O_57,N_29568,N_29645);
nand UO_58 (O_58,N_29661,N_28508);
and UO_59 (O_59,N_28809,N_28933);
nor UO_60 (O_60,N_29457,N_29140);
or UO_61 (O_61,N_29624,N_28663);
nor UO_62 (O_62,N_28545,N_29679);
xnor UO_63 (O_63,N_29872,N_28680);
or UO_64 (O_64,N_29109,N_28631);
or UO_65 (O_65,N_29858,N_28960);
or UO_66 (O_66,N_29484,N_29016);
or UO_67 (O_67,N_29943,N_29787);
and UO_68 (O_68,N_28742,N_28540);
xor UO_69 (O_69,N_29373,N_29170);
nand UO_70 (O_70,N_29830,N_28691);
or UO_71 (O_71,N_28635,N_28550);
xor UO_72 (O_72,N_29379,N_29623);
nand UO_73 (O_73,N_28887,N_29689);
nand UO_74 (O_74,N_29353,N_29037);
nand UO_75 (O_75,N_29116,N_29899);
xor UO_76 (O_76,N_28552,N_29932);
or UO_77 (O_77,N_29157,N_29417);
nand UO_78 (O_78,N_28846,N_29569);
nor UO_79 (O_79,N_28995,N_28959);
or UO_80 (O_80,N_29676,N_29409);
and UO_81 (O_81,N_29898,N_28815);
or UO_82 (O_82,N_29182,N_29390);
or UO_83 (O_83,N_29891,N_29148);
xor UO_84 (O_84,N_28601,N_28731);
nand UO_85 (O_85,N_29771,N_29431);
nor UO_86 (O_86,N_29311,N_28813);
xor UO_87 (O_87,N_29534,N_29589);
and UO_88 (O_88,N_29257,N_28716);
nor UO_89 (O_89,N_29752,N_29615);
and UO_90 (O_90,N_29997,N_29096);
or UO_91 (O_91,N_29376,N_29401);
nand UO_92 (O_92,N_28589,N_29788);
nor UO_93 (O_93,N_28902,N_29341);
or UO_94 (O_94,N_29942,N_29146);
and UO_95 (O_95,N_29672,N_28976);
or UO_96 (O_96,N_29528,N_28875);
nand UO_97 (O_97,N_29836,N_29829);
and UO_98 (O_98,N_29443,N_29078);
xor UO_99 (O_99,N_29772,N_29210);
and UO_100 (O_100,N_29607,N_28996);
nor UO_101 (O_101,N_28661,N_29205);
nor UO_102 (O_102,N_28934,N_28893);
and UO_103 (O_103,N_29495,N_28938);
nor UO_104 (O_104,N_28954,N_29886);
nor UO_105 (O_105,N_28533,N_29993);
nor UO_106 (O_106,N_29703,N_28586);
or UO_107 (O_107,N_28563,N_29388);
or UO_108 (O_108,N_29045,N_29444);
or UO_109 (O_109,N_29876,N_29693);
and UO_110 (O_110,N_28833,N_29913);
nor UO_111 (O_111,N_29826,N_29934);
xor UO_112 (O_112,N_28525,N_28736);
nand UO_113 (O_113,N_29208,N_29158);
nor UO_114 (O_114,N_29961,N_28708);
xor UO_115 (O_115,N_29980,N_29558);
nor UO_116 (O_116,N_29144,N_29462);
or UO_117 (O_117,N_29825,N_29290);
nand UO_118 (O_118,N_29364,N_29628);
or UO_119 (O_119,N_29377,N_28949);
and UO_120 (O_120,N_29209,N_28616);
xnor UO_121 (O_121,N_28511,N_29179);
xnor UO_122 (O_122,N_28862,N_28591);
nor UO_123 (O_123,N_29512,N_29214);
xor UO_124 (O_124,N_28615,N_28982);
nand UO_125 (O_125,N_29337,N_29099);
xnor UO_126 (O_126,N_29375,N_29845);
nand UO_127 (O_127,N_29954,N_29466);
and UO_128 (O_128,N_29621,N_28730);
nand UO_129 (O_129,N_28930,N_29967);
nand UO_130 (O_130,N_28623,N_29996);
or UO_131 (O_131,N_29593,N_28758);
or UO_132 (O_132,N_28764,N_29838);
xnor UO_133 (O_133,N_28627,N_28796);
xnor UO_134 (O_134,N_29759,N_29413);
nor UO_135 (O_135,N_29806,N_29966);
and UO_136 (O_136,N_29692,N_29956);
or UO_137 (O_137,N_29030,N_28883);
nor UO_138 (O_138,N_28712,N_29054);
nor UO_139 (O_139,N_28757,N_29344);
xor UO_140 (O_140,N_29268,N_29665);
xor UO_141 (O_141,N_29588,N_29392);
xor UO_142 (O_142,N_28531,N_28989);
and UO_143 (O_143,N_29218,N_29698);
nor UO_144 (O_144,N_29040,N_29374);
and UO_145 (O_145,N_28789,N_29012);
or UO_146 (O_146,N_28908,N_29737);
nor UO_147 (O_147,N_29516,N_28700);
nor UO_148 (O_148,N_29060,N_28876);
xnor UO_149 (O_149,N_28565,N_29683);
and UO_150 (O_150,N_28707,N_29133);
and UO_151 (O_151,N_28861,N_28767);
and UO_152 (O_152,N_29239,N_28807);
nor UO_153 (O_153,N_28926,N_29339);
nand UO_154 (O_154,N_29174,N_28541);
and UO_155 (O_155,N_29890,N_29843);
nor UO_156 (O_156,N_29137,N_29088);
nor UO_157 (O_157,N_29055,N_28664);
xor UO_158 (O_158,N_28561,N_29775);
or UO_159 (O_159,N_28958,N_29673);
nand UO_160 (O_160,N_29230,N_29396);
nor UO_161 (O_161,N_29561,N_29371);
nand UO_162 (O_162,N_28993,N_29193);
xor UO_163 (O_163,N_29253,N_29324);
nor UO_164 (O_164,N_29405,N_28797);
nor UO_165 (O_165,N_29637,N_29100);
or UO_166 (O_166,N_28885,N_29955);
and UO_167 (O_167,N_29892,N_28822);
or UO_168 (O_168,N_28642,N_29519);
or UO_169 (O_169,N_29307,N_28759);
nand UO_170 (O_170,N_29705,N_29172);
nand UO_171 (O_171,N_29385,N_28500);
xor UO_172 (O_172,N_29735,N_28608);
or UO_173 (O_173,N_29243,N_29948);
nand UO_174 (O_174,N_28978,N_29856);
and UO_175 (O_175,N_28944,N_28922);
nor UO_176 (O_176,N_29411,N_29192);
nand UO_177 (O_177,N_29128,N_29090);
xor UO_178 (O_178,N_29748,N_29629);
or UO_179 (O_179,N_29647,N_28782);
xor UO_180 (O_180,N_28769,N_29984);
and UO_181 (O_181,N_29949,N_28799);
nand UO_182 (O_182,N_28751,N_29605);
or UO_183 (O_183,N_29896,N_28667);
or UO_184 (O_184,N_29130,N_29450);
xnor UO_185 (O_185,N_28649,N_28805);
nor UO_186 (O_186,N_29087,N_29491);
xnor UO_187 (O_187,N_29909,N_28723);
and UO_188 (O_188,N_29802,N_29009);
nor UO_189 (O_189,N_28562,N_29143);
and UO_190 (O_190,N_28763,N_29750);
nor UO_191 (O_191,N_28841,N_29542);
or UO_192 (O_192,N_28600,N_29842);
nor UO_193 (O_193,N_29789,N_29520);
or UO_194 (O_194,N_29011,N_28880);
and UO_195 (O_195,N_29755,N_28629);
and UO_196 (O_196,N_29021,N_29778);
nor UO_197 (O_197,N_29820,N_29704);
and UO_198 (O_198,N_29719,N_29560);
or UO_199 (O_199,N_29577,N_29473);
or UO_200 (O_200,N_28928,N_29237);
nor UO_201 (O_201,N_29940,N_29887);
and UO_202 (O_202,N_28519,N_28690);
xnor UO_203 (O_203,N_29173,N_29132);
or UO_204 (O_204,N_28522,N_28913);
nand UO_205 (O_205,N_29599,N_29544);
xor UO_206 (O_206,N_28587,N_29840);
and UO_207 (O_207,N_29425,N_29490);
xnor UO_208 (O_208,N_29010,N_29415);
nor UO_209 (O_209,N_29420,N_29236);
xnor UO_210 (O_210,N_29131,N_29202);
and UO_211 (O_211,N_29517,N_29454);
xnor UO_212 (O_212,N_29223,N_29640);
and UO_213 (O_213,N_29059,N_29465);
or UO_214 (O_214,N_29112,N_28595);
xor UO_215 (O_215,N_29662,N_29766);
or UO_216 (O_216,N_29455,N_29039);
nand UO_217 (O_217,N_29077,N_29211);
and UO_218 (O_218,N_28739,N_29656);
or UO_219 (O_219,N_29436,N_29287);
nand UO_220 (O_220,N_29933,N_28747);
and UO_221 (O_221,N_29976,N_28842);
nor UO_222 (O_222,N_28577,N_29981);
and UO_223 (O_223,N_29270,N_29452);
or UO_224 (O_224,N_28640,N_28795);
nand UO_225 (O_225,N_29483,N_29975);
or UO_226 (O_226,N_28564,N_28572);
xor UO_227 (O_227,N_29908,N_29768);
or UO_228 (O_228,N_29584,N_29477);
nand UO_229 (O_229,N_28925,N_29278);
xnor UO_230 (O_230,N_29583,N_28968);
and UO_231 (O_231,N_29325,N_29818);
xor UO_232 (O_232,N_29219,N_29501);
or UO_233 (O_233,N_29809,N_28991);
or UO_234 (O_234,N_29485,N_28634);
and UO_235 (O_235,N_29220,N_29084);
nor UO_236 (O_236,N_29811,N_29515);
or UO_237 (O_237,N_28660,N_28865);
nand UO_238 (O_238,N_29958,N_29945);
xor UO_239 (O_239,N_29121,N_28713);
or UO_240 (O_240,N_28785,N_29176);
xor UO_241 (O_241,N_28953,N_29368);
and UO_242 (O_242,N_29824,N_29275);
nand UO_243 (O_243,N_29741,N_29707);
xor UO_244 (O_244,N_28814,N_29327);
nand UO_245 (O_245,N_29286,N_28872);
and UO_246 (O_246,N_29930,N_29075);
nand UO_247 (O_247,N_29482,N_28983);
or UO_248 (O_248,N_29715,N_28969);
and UO_249 (O_249,N_29742,N_29507);
and UO_250 (O_250,N_28720,N_29860);
and UO_251 (O_251,N_28844,N_28967);
nand UO_252 (O_252,N_29957,N_28684);
nor UO_253 (O_253,N_29292,N_29499);
and UO_254 (O_254,N_28864,N_29739);
nand UO_255 (O_255,N_29445,N_29827);
xor UO_256 (O_256,N_29797,N_29604);
nor UO_257 (O_257,N_29002,N_29563);
nand UO_258 (O_258,N_28659,N_29245);
or UO_259 (O_259,N_28892,N_29770);
xor UO_260 (O_260,N_29302,N_29639);
xnor UO_261 (O_261,N_28670,N_29232);
nor UO_262 (O_262,N_29690,N_28819);
and UO_263 (O_263,N_29289,N_29190);
or UO_264 (O_264,N_28897,N_29773);
nor UO_265 (O_265,N_29034,N_29105);
xnor UO_266 (O_266,N_29728,N_28936);
xor UO_267 (O_267,N_28620,N_29555);
nand UO_268 (O_268,N_28788,N_28639);
or UO_269 (O_269,N_29630,N_29823);
and UO_270 (O_270,N_28966,N_29785);
xor UO_271 (O_271,N_29983,N_29688);
and UO_272 (O_272,N_28579,N_29467);
or UO_273 (O_273,N_29545,N_29917);
xnor UO_274 (O_274,N_29271,N_29310);
and UO_275 (O_275,N_28553,N_29330);
or UO_276 (O_276,N_28625,N_29298);
nand UO_277 (O_277,N_29878,N_29763);
xor UO_278 (O_278,N_28889,N_28899);
and UO_279 (O_279,N_29633,N_29076);
or UO_280 (O_280,N_29986,N_29697);
or UO_281 (O_281,N_29102,N_29175);
or UO_282 (O_282,N_29888,N_29536);
or UO_283 (O_283,N_29726,N_28513);
nor UO_284 (O_284,N_29387,N_29221);
xnor UO_285 (O_285,N_29509,N_29026);
or UO_286 (O_286,N_28900,N_29803);
nor UO_287 (O_287,N_29063,N_29796);
and UO_288 (O_288,N_29521,N_29080);
nand UO_289 (O_289,N_29681,N_28858);
nor UO_290 (O_290,N_28517,N_28555);
and UO_291 (O_291,N_29594,N_29488);
xor UO_292 (O_292,N_28912,N_28650);
or UO_293 (O_293,N_29168,N_29541);
nand UO_294 (O_294,N_28962,N_29928);
xor UO_295 (O_295,N_29638,N_28811);
or UO_296 (O_296,N_29154,N_29999);
nand UO_297 (O_297,N_29862,N_29300);
xnor UO_298 (O_298,N_29769,N_29556);
nor UO_299 (O_299,N_29259,N_28749);
and UO_300 (O_300,N_29574,N_29419);
nand UO_301 (O_301,N_29000,N_29358);
or UO_302 (O_302,N_29525,N_29496);
and UO_303 (O_303,N_28950,N_28588);
nand UO_304 (O_304,N_29655,N_29895);
and UO_305 (O_305,N_28549,N_29181);
or UO_306 (O_306,N_29794,N_28607);
nor UO_307 (O_307,N_29038,N_28973);
xnor UO_308 (O_308,N_28853,N_28596);
and UO_309 (O_309,N_29498,N_29422);
or UO_310 (O_310,N_28802,N_28673);
and UO_311 (O_311,N_29108,N_28604);
or UO_312 (O_312,N_29288,N_29901);
xor UO_313 (O_313,N_29061,N_29363);
nand UO_314 (O_314,N_29651,N_29167);
xnor UO_315 (O_315,N_29006,N_29854);
or UO_316 (O_316,N_29894,N_29258);
or UO_317 (O_317,N_29240,N_29150);
nor UO_318 (O_318,N_29217,N_29147);
xnor UO_319 (O_319,N_29753,N_28677);
and UO_320 (O_320,N_29391,N_29326);
xnor UO_321 (O_321,N_29372,N_29792);
xnor UO_322 (O_322,N_28599,N_29267);
and UO_323 (O_323,N_29367,N_29834);
xnor UO_324 (O_324,N_29303,N_28877);
nand UO_325 (O_325,N_28942,N_29897);
xnor UO_326 (O_326,N_29625,N_29359);
or UO_327 (O_327,N_29733,N_29281);
nand UO_328 (O_328,N_29015,N_29106);
nor UO_329 (O_329,N_28857,N_29319);
and UO_330 (O_330,N_28952,N_29712);
or UO_331 (O_331,N_28729,N_29432);
and UO_332 (O_332,N_29049,N_29079);
and UO_333 (O_333,N_28648,N_29553);
and UO_334 (O_334,N_28910,N_29965);
nand UO_335 (O_335,N_29348,N_29642);
nand UO_336 (O_336,N_29458,N_29852);
nand UO_337 (O_337,N_28671,N_29156);
nor UO_338 (O_338,N_28994,N_28733);
or UO_339 (O_339,N_29643,N_29486);
or UO_340 (O_340,N_29867,N_29328);
or UO_341 (O_341,N_29713,N_29837);
or UO_342 (O_342,N_29864,N_29282);
and UO_343 (O_343,N_28837,N_29189);
nand UO_344 (O_344,N_28710,N_29043);
or UO_345 (O_345,N_29603,N_29821);
nor UO_346 (O_346,N_29875,N_28585);
nor UO_347 (O_347,N_29291,N_29201);
nor UO_348 (O_348,N_29922,N_28526);
xnor UO_349 (O_349,N_29863,N_29929);
xor UO_350 (O_350,N_28611,N_28836);
xor UO_351 (O_351,N_28786,N_29317);
or UO_352 (O_352,N_29722,N_28744);
and UO_353 (O_353,N_29398,N_29427);
and UO_354 (O_354,N_29127,N_29044);
or UO_355 (O_355,N_29849,N_29668);
xnor UO_356 (O_356,N_29366,N_28824);
or UO_357 (O_357,N_28534,N_29974);
nand UO_358 (O_358,N_28847,N_29350);
nand UO_359 (O_359,N_28605,N_28931);
nor UO_360 (O_360,N_29003,N_29118);
or UO_361 (O_361,N_29653,N_29437);
or UO_362 (O_362,N_28725,N_29447);
nand UO_363 (O_363,N_28834,N_29032);
nor UO_364 (O_364,N_28665,N_28935);
or UO_365 (O_365,N_29407,N_29180);
or UO_366 (O_366,N_29721,N_28547);
or UO_367 (O_367,N_28624,N_29720);
or UO_368 (O_368,N_28939,N_29426);
nand UO_369 (O_369,N_28686,N_29110);
or UO_370 (O_370,N_29497,N_29611);
or UO_371 (O_371,N_28560,N_28929);
nor UO_372 (O_372,N_29164,N_28669);
nand UO_373 (O_373,N_28637,N_29754);
xnor UO_374 (O_374,N_29155,N_29058);
or UO_375 (O_375,N_28554,N_29644);
nor UO_376 (O_376,N_29423,N_29559);
nor UO_377 (O_377,N_29786,N_29123);
nand UO_378 (O_378,N_29254,N_29227);
or UO_379 (O_379,N_29979,N_28558);
or UO_380 (O_380,N_29206,N_28835);
and UO_381 (O_381,N_29874,N_28803);
xor UO_382 (O_382,N_29765,N_28945);
and UO_383 (O_383,N_28571,N_29008);
xnor UO_384 (O_384,N_28636,N_29381);
nand UO_385 (O_385,N_29095,N_28878);
nand UO_386 (O_386,N_29001,N_29481);
xnor UO_387 (O_387,N_29360,N_29994);
nand UO_388 (O_388,N_29416,N_29471);
nor UO_389 (O_389,N_28521,N_29631);
xor UO_390 (O_390,N_29652,N_29273);
or UO_391 (O_391,N_29336,N_29831);
and UO_392 (O_392,N_28711,N_29429);
and UO_393 (O_393,N_29433,N_28658);
and UO_394 (O_394,N_29659,N_29758);
or UO_395 (O_395,N_29160,N_29613);
nand UO_396 (O_396,N_29906,N_29591);
and UO_397 (O_397,N_29814,N_28970);
or UO_398 (O_398,N_29808,N_28546);
xor UO_399 (O_399,N_29912,N_29596);
or UO_400 (O_400,N_29518,N_28685);
and UO_401 (O_401,N_29658,N_29262);
or UO_402 (O_402,N_29346,N_28651);
or UO_403 (O_403,N_29320,N_29163);
or UO_404 (O_404,N_28918,N_29522);
nand UO_405 (O_405,N_28990,N_28975);
or UO_406 (O_406,N_29269,N_29389);
or UO_407 (O_407,N_28548,N_29523);
xor UO_408 (O_408,N_28652,N_29985);
and UO_409 (O_409,N_28714,N_29169);
nor UO_410 (O_410,N_28812,N_28808);
nand UO_411 (O_411,N_29729,N_28515);
nor UO_412 (O_412,N_28632,N_29101);
or UO_413 (O_413,N_29071,N_29552);
or UO_414 (O_414,N_29141,N_29313);
nand UO_415 (O_415,N_29990,N_28871);
nor UO_416 (O_416,N_29592,N_29526);
xor UO_417 (O_417,N_29266,N_29068);
and UO_418 (O_418,N_29403,N_28501);
or UO_419 (O_419,N_28520,N_29691);
nand UO_420 (O_420,N_29085,N_29550);
or UO_421 (O_421,N_29578,N_29434);
and UO_422 (O_422,N_28746,N_28843);
nor UO_423 (O_423,N_28527,N_29274);
or UO_424 (O_424,N_29587,N_29261);
or UO_425 (O_425,N_28696,N_29988);
nor UO_426 (O_426,N_29365,N_29666);
nor UO_427 (O_427,N_29777,N_28672);
and UO_428 (O_428,N_29612,N_29460);
and UO_429 (O_429,N_28937,N_29277);
or UO_430 (O_430,N_29056,N_29046);
xor UO_431 (O_431,N_28704,N_29280);
or UO_432 (O_432,N_29815,N_28963);
and UO_433 (O_433,N_29935,N_28832);
xor UO_434 (O_434,N_28901,N_28575);
or UO_435 (O_435,N_29321,N_29461);
and UO_436 (O_436,N_28576,N_28556);
nor UO_437 (O_437,N_29514,N_29256);
nand UO_438 (O_438,N_28831,N_29023);
xor UO_439 (O_439,N_28699,N_29601);
nand UO_440 (O_440,N_28754,N_29585);
nand UO_441 (O_441,N_28916,N_29053);
and UO_442 (O_442,N_28766,N_29197);
xor UO_443 (O_443,N_28633,N_28826);
nor UO_444 (O_444,N_28947,N_29504);
xor UO_445 (O_445,N_28581,N_28728);
nor UO_446 (O_446,N_29557,N_28793);
nand UO_447 (O_447,N_29309,N_29885);
or UO_448 (O_448,N_28598,N_28886);
nor UO_449 (O_449,N_28781,N_29115);
nand UO_450 (O_450,N_29725,N_29474);
or UO_451 (O_451,N_28840,N_29500);
or UO_452 (O_452,N_29968,N_29332);
xnor UO_453 (O_453,N_29356,N_28743);
and UO_454 (O_454,N_29648,N_29805);
or UO_455 (O_455,N_28724,N_29472);
xnor UO_456 (O_456,N_29779,N_29590);
or UO_457 (O_457,N_29151,N_28722);
nor UO_458 (O_458,N_29196,N_28778);
nor UO_459 (O_459,N_29362,N_29546);
nand UO_460 (O_460,N_28726,N_29323);
xor UO_461 (O_461,N_29370,N_28999);
nor UO_462 (O_462,N_28692,N_29696);
nor UO_463 (O_463,N_29764,N_29687);
nor UO_464 (O_464,N_29036,N_28727);
nor UO_465 (O_465,N_29538,N_29072);
nand UO_466 (O_466,N_29793,N_29305);
or UO_467 (O_467,N_28800,N_28985);
and UO_468 (O_468,N_28719,N_28755);
nor UO_469 (O_469,N_28740,N_28641);
nor UO_470 (O_470,N_29795,N_29134);
and UO_471 (O_471,N_29616,N_29866);
and UO_472 (O_472,N_28617,N_28783);
nor UO_473 (O_473,N_29677,N_29952);
nand UO_474 (O_474,N_29680,N_29249);
nor UO_475 (O_475,N_28984,N_29216);
nand UO_476 (O_476,N_28679,N_29537);
xor UO_477 (O_477,N_28830,N_29921);
or UO_478 (O_478,N_29004,N_28644);
nor UO_479 (O_479,N_28867,N_28881);
nor UO_480 (O_480,N_28845,N_29920);
or UO_481 (O_481,N_29937,N_29340);
or UO_482 (O_482,N_29524,N_29925);
nor UO_483 (O_483,N_28851,N_28956);
nor UO_484 (O_484,N_29418,N_28906);
nand UO_485 (O_485,N_29847,N_29657);
and UO_486 (O_486,N_28655,N_29903);
nand UO_487 (O_487,N_29005,N_29028);
xor UO_488 (O_488,N_29551,N_28734);
xnor UO_489 (O_489,N_29186,N_29404);
nor UO_490 (O_490,N_29870,N_28890);
nor UO_491 (O_491,N_29740,N_28578);
nor UO_492 (O_492,N_28718,N_29745);
or UO_493 (O_493,N_29716,N_29632);
or UO_494 (O_494,N_29129,N_29865);
nor UO_495 (O_495,N_29708,N_29767);
nor UO_496 (O_496,N_29675,N_28957);
xor UO_497 (O_497,N_29347,N_28817);
xor UO_498 (O_498,N_29231,N_29178);
or UO_499 (O_499,N_29734,N_29978);
nand UO_500 (O_500,N_28610,N_29798);
nand UO_501 (O_501,N_29031,N_29812);
and UO_502 (O_502,N_29670,N_28948);
nand UO_503 (O_503,N_29738,N_28675);
or UO_504 (O_504,N_29660,N_29900);
or UO_505 (O_505,N_28762,N_29861);
nand UO_506 (O_506,N_29459,N_28810);
or UO_507 (O_507,N_29995,N_29065);
or UO_508 (O_508,N_29963,N_29857);
and UO_509 (O_509,N_29969,N_28512);
nand UO_510 (O_510,N_28971,N_29889);
nand UO_511 (O_511,N_28715,N_28666);
xnor UO_512 (O_512,N_28603,N_29614);
or UO_513 (O_513,N_28924,N_28551);
and UO_514 (O_514,N_29195,N_29017);
or UO_515 (O_515,N_29421,N_29844);
and UO_516 (O_516,N_29664,N_28904);
nor UO_517 (O_517,N_29620,N_28647);
xnor UO_518 (O_518,N_29799,N_28506);
nor UO_519 (O_519,N_29035,N_29489);
nand UO_520 (O_520,N_29487,N_29682);
nor UO_521 (O_521,N_29235,N_29361);
xnor UO_522 (O_522,N_29304,N_29318);
or UO_523 (O_523,N_29333,N_29597);
nor UO_524 (O_524,N_28839,N_29944);
or UO_525 (O_525,N_28567,N_29475);
xor UO_526 (O_526,N_29103,N_29018);
xor UO_527 (O_527,N_29505,N_29962);
or UO_528 (O_528,N_29800,N_29126);
nand UO_529 (O_529,N_29246,N_29746);
xnor UO_530 (O_530,N_29464,N_29081);
or UO_531 (O_531,N_29092,N_28544);
nand UO_532 (O_532,N_28750,N_29832);
nand UO_533 (O_533,N_28709,N_28701);
or UO_534 (O_534,N_28569,N_28693);
nor UO_535 (O_535,N_28787,N_28869);
or UO_536 (O_536,N_29272,N_29113);
nor UO_537 (O_537,N_29717,N_28980);
nand UO_538 (O_538,N_29177,N_28612);
nand UO_539 (O_539,N_29439,N_28594);
nor UO_540 (O_540,N_29159,N_28891);
nand UO_541 (O_541,N_28518,N_28986);
xnor UO_542 (O_542,N_29165,N_29723);
or UO_543 (O_543,N_29204,N_29393);
xor UO_544 (O_544,N_29402,N_29562);
nor UO_545 (O_545,N_29586,N_29873);
nor UO_546 (O_546,N_28741,N_29349);
xnor UO_547 (O_547,N_29188,N_28502);
xor UO_548 (O_548,N_29669,N_29222);
and UO_549 (O_549,N_29608,N_28997);
xor UO_550 (O_550,N_28852,N_29233);
or UO_551 (O_551,N_29355,N_29566);
xnor UO_552 (O_552,N_29369,N_28738);
nand UO_553 (O_553,N_29781,N_28529);
or UO_554 (O_554,N_28609,N_29083);
nor UO_555 (O_555,N_29636,N_28979);
nand UO_556 (O_556,N_29595,N_29911);
or UO_557 (O_557,N_28717,N_29510);
or UO_558 (O_558,N_28523,N_29627);
nor UO_559 (O_559,N_29136,N_29649);
or UO_560 (O_560,N_29724,N_29386);
nor UO_561 (O_561,N_28911,N_29153);
xor UO_562 (O_562,N_29706,N_29073);
or UO_563 (O_563,N_29819,N_29991);
or UO_564 (O_564,N_29869,N_29880);
and UO_565 (O_565,N_29316,N_28703);
nand UO_566 (O_566,N_28606,N_29822);
or UO_567 (O_567,N_28898,N_28849);
and UO_568 (O_568,N_28998,N_28961);
xnor UO_569 (O_569,N_28698,N_29067);
nand UO_570 (O_570,N_28917,N_28882);
or UO_571 (O_571,N_29228,N_29927);
nand UO_572 (O_572,N_28504,N_28771);
or UO_573 (O_573,N_29051,N_29959);
or UO_574 (O_574,N_28972,N_28974);
and UO_575 (O_575,N_29950,N_29695);
nand UO_576 (O_576,N_28735,N_29783);
nor UO_577 (O_577,N_28681,N_29916);
and UO_578 (O_578,N_29064,N_28619);
or UO_579 (O_579,N_29506,N_29992);
nor UO_580 (O_580,N_29410,N_29914);
nor UO_581 (O_581,N_29382,N_29334);
or UO_582 (O_582,N_28792,N_29502);
or UO_583 (O_583,N_29476,N_29380);
and UO_584 (O_584,N_28674,N_29066);
xor UO_585 (O_585,N_28532,N_29700);
and UO_586 (O_586,N_29234,N_28618);
nand UO_587 (O_587,N_29479,N_29301);
xnor UO_588 (O_588,N_28866,N_29276);
nand UO_589 (O_589,N_29314,N_28694);
or UO_590 (O_590,N_28873,N_29435);
xnor UO_591 (O_591,N_29671,N_29424);
and UO_592 (O_592,N_29329,N_28756);
or UO_593 (O_593,N_29828,N_29622);
nor UO_594 (O_594,N_28761,N_29879);
and UO_595 (O_595,N_29939,N_28638);
nor UO_596 (O_596,N_28530,N_29025);
or UO_597 (O_597,N_29299,N_28538);
xnor UO_598 (O_598,N_29250,N_28977);
xor UO_599 (O_599,N_29057,N_29702);
nand UO_600 (O_600,N_29029,N_28592);
and UO_601 (O_601,N_29312,N_28628);
xnor UO_602 (O_602,N_28987,N_29718);
or UO_603 (O_603,N_28909,N_28516);
xor UO_604 (O_604,N_29111,N_29699);
xor UO_605 (O_605,N_29242,N_29027);
and UO_606 (O_606,N_28919,N_28613);
and UO_607 (O_607,N_29199,N_28816);
nor UO_608 (O_608,N_28791,N_28524);
or UO_609 (O_609,N_29352,N_29213);
or UO_610 (O_610,N_29816,N_29548);
and UO_611 (O_611,N_29492,N_29469);
xnor UO_612 (O_612,N_28859,N_28542);
nand UO_613 (O_613,N_29971,N_29641);
or UO_614 (O_614,N_29171,N_28621);
nand UO_615 (O_615,N_29678,N_28932);
and UO_616 (O_616,N_29440,N_28528);
nand UO_617 (O_617,N_28829,N_29575);
or UO_618 (O_618,N_29194,N_29701);
nand UO_619 (O_619,N_28821,N_28745);
nand UO_620 (O_620,N_28894,N_29451);
nand UO_621 (O_621,N_29549,N_29033);
nand UO_622 (O_622,N_28779,N_28687);
nand UO_623 (O_623,N_29042,N_29283);
xor UO_624 (O_624,N_29511,N_28772);
nand UO_625 (O_625,N_29850,N_29964);
or UO_626 (O_626,N_28654,N_28964);
xor UO_627 (O_627,N_29070,N_28737);
nand UO_628 (O_628,N_29801,N_28776);
and UO_629 (O_629,N_29905,N_29791);
xor UO_630 (O_630,N_29019,N_28854);
nor UO_631 (O_631,N_28940,N_29378);
nand UO_632 (O_632,N_28823,N_29936);
xnor UO_633 (O_633,N_28870,N_29579);
nor UO_634 (O_634,N_29438,N_29807);
and UO_635 (O_635,N_29756,N_28790);
and UO_636 (O_636,N_29531,N_28537);
nand UO_637 (O_637,N_29835,N_28583);
nor UO_638 (O_638,N_29047,N_29014);
and UO_639 (O_639,N_28760,N_28535);
or UO_640 (O_640,N_28923,N_29762);
xnor UO_641 (O_641,N_29074,N_29839);
and UO_642 (O_642,N_29107,N_28905);
or UO_643 (O_643,N_29902,N_28676);
nand UO_644 (O_644,N_29125,N_29248);
nand UO_645 (O_645,N_28888,N_28965);
nor UO_646 (O_646,N_29709,N_28943);
nor UO_647 (O_647,N_29751,N_28732);
nand UO_648 (O_648,N_29412,N_29931);
xnor UO_649 (O_649,N_29089,N_29203);
and UO_650 (O_650,N_29804,N_29989);
nor UO_651 (O_651,N_28780,N_29020);
and UO_652 (O_652,N_29571,N_29910);
xnor UO_653 (O_653,N_28662,N_29198);
or UO_654 (O_654,N_29229,N_28896);
and UO_655 (O_655,N_29093,N_28868);
and UO_656 (O_656,N_28860,N_28580);
and UO_657 (O_657,N_29453,N_28678);
xnor UO_658 (O_658,N_29972,N_29264);
and UO_659 (O_659,N_29610,N_28825);
and UO_660 (O_660,N_28570,N_28702);
xor UO_661 (O_661,N_28566,N_28951);
nor UO_662 (O_662,N_29572,N_28657);
xnor UO_663 (O_663,N_29351,N_29430);
nor UO_664 (O_664,N_29535,N_29354);
nor UO_665 (O_665,N_29565,N_29973);
xor UO_666 (O_666,N_29494,N_29145);
nor UO_667 (O_667,N_29532,N_29414);
and UO_668 (O_668,N_29446,N_29600);
nor UO_669 (O_669,N_29187,N_29883);
and UO_670 (O_670,N_29926,N_28573);
xnor UO_671 (O_671,N_29853,N_29086);
or UO_672 (O_672,N_29124,N_28683);
and UO_673 (O_673,N_28981,N_29938);
xor UO_674 (O_674,N_29442,N_29448);
nand UO_675 (O_675,N_29345,N_29646);
xor UO_676 (O_676,N_28827,N_28895);
and UO_677 (O_677,N_29923,N_29166);
and UO_678 (O_678,N_28656,N_29918);
or UO_679 (O_679,N_29749,N_29244);
or UO_680 (O_680,N_28505,N_29919);
xnor UO_681 (O_681,N_29907,N_28770);
xnor UO_682 (O_682,N_28643,N_28557);
or UO_683 (O_683,N_29977,N_29135);
nor UO_684 (O_684,N_29609,N_29859);
nand UO_685 (O_685,N_28539,N_29855);
and UO_686 (O_686,N_29215,N_29953);
and UO_687 (O_687,N_28695,N_29635);
nor UO_688 (O_688,N_29062,N_29871);
xor UO_689 (O_689,N_28646,N_29343);
xnor UO_690 (O_690,N_28920,N_29247);
nor UO_691 (O_691,N_28988,N_29760);
or UO_692 (O_692,N_29606,N_28828);
nor UO_693 (O_693,N_29877,N_29530);
xnor UO_694 (O_694,N_29449,N_29293);
nand UO_695 (O_695,N_29580,N_29408);
nor UO_696 (O_696,N_28507,N_29982);
and UO_697 (O_697,N_28804,N_29120);
and UO_698 (O_698,N_29529,N_28992);
nand UO_699 (O_699,N_29543,N_28777);
or UO_700 (O_700,N_29743,N_29207);
xnor UO_701 (O_701,N_29731,N_29335);
xnor UO_702 (O_702,N_29241,N_29265);
and UO_703 (O_703,N_29295,N_29297);
or UO_704 (O_704,N_29564,N_29941);
nand UO_705 (O_705,N_29493,N_29634);
nand UO_706 (O_706,N_29757,N_28597);
xor UO_707 (O_707,N_29185,N_29397);
and UO_708 (O_708,N_29478,N_28775);
nand UO_709 (O_709,N_29225,N_29400);
nor UO_710 (O_710,N_29251,N_28602);
nand UO_711 (O_711,N_29761,N_29868);
or UO_712 (O_712,N_29383,N_29527);
nand UO_713 (O_713,N_29463,N_29513);
and UO_714 (O_714,N_29480,N_29714);
nor UO_715 (O_715,N_29581,N_28855);
and UO_716 (O_716,N_29619,N_29456);
or UO_717 (O_717,N_29284,N_29162);
xnor UO_718 (O_718,N_29041,N_28688);
or UO_719 (O_719,N_29184,N_29097);
or UO_720 (O_720,N_29338,N_28748);
or UO_721 (O_721,N_29122,N_29915);
or UO_722 (O_722,N_28509,N_29539);
nand UO_723 (O_723,N_28753,N_29667);
or UO_724 (O_724,N_29406,N_29082);
nand UO_725 (O_725,N_28510,N_29470);
nor UO_726 (O_726,N_29052,N_29468);
nor UO_727 (O_727,N_28774,N_29663);
and UO_728 (O_728,N_28705,N_28798);
nor UO_729 (O_729,N_29848,N_28838);
and UO_730 (O_730,N_29161,N_29987);
and UO_731 (O_731,N_29582,N_29069);
nor UO_732 (O_732,N_28593,N_29884);
nor UO_733 (O_733,N_29306,N_29881);
nor UO_734 (O_734,N_29238,N_29142);
and UO_735 (O_735,N_29331,N_29094);
nor UO_736 (O_736,N_29951,N_29117);
xor UO_737 (O_737,N_29308,N_29183);
and UO_738 (O_738,N_29260,N_29711);
or UO_739 (O_739,N_29817,N_28514);
nor UO_740 (O_740,N_29441,N_28801);
or UO_741 (O_741,N_28927,N_28794);
or UO_742 (O_742,N_29384,N_29833);
and UO_743 (O_743,N_28879,N_29685);
or UO_744 (O_744,N_29554,N_29152);
nand UO_745 (O_745,N_28721,N_28653);
xor UO_746 (O_746,N_28689,N_29024);
nand UO_747 (O_747,N_28622,N_29285);
nand UO_748 (O_748,N_29904,N_29263);
nor UO_749 (O_749,N_28784,N_29813);
nand UO_750 (O_750,N_28912,N_29662);
xnor UO_751 (O_751,N_29784,N_29128);
xnor UO_752 (O_752,N_29692,N_28672);
nand UO_753 (O_753,N_29831,N_29671);
xnor UO_754 (O_754,N_29280,N_28706);
nor UO_755 (O_755,N_29915,N_29782);
xor UO_756 (O_756,N_29525,N_29350);
nand UO_757 (O_757,N_29665,N_28514);
and UO_758 (O_758,N_28537,N_29443);
nor UO_759 (O_759,N_29375,N_29772);
or UO_760 (O_760,N_29588,N_29201);
xnor UO_761 (O_761,N_28666,N_29301);
nand UO_762 (O_762,N_29132,N_29881);
nand UO_763 (O_763,N_29707,N_29210);
and UO_764 (O_764,N_29959,N_29041);
nand UO_765 (O_765,N_29493,N_29857);
and UO_766 (O_766,N_29437,N_29217);
nand UO_767 (O_767,N_29264,N_29080);
and UO_768 (O_768,N_29629,N_29756);
and UO_769 (O_769,N_28593,N_28637);
nand UO_770 (O_770,N_29536,N_28718);
and UO_771 (O_771,N_29710,N_29347);
nor UO_772 (O_772,N_28825,N_29807);
nor UO_773 (O_773,N_28782,N_28687);
xnor UO_774 (O_774,N_29509,N_28700);
xor UO_775 (O_775,N_29615,N_29329);
nor UO_776 (O_776,N_28569,N_29690);
or UO_777 (O_777,N_28633,N_28738);
or UO_778 (O_778,N_29474,N_29440);
nor UO_779 (O_779,N_29865,N_29537);
nand UO_780 (O_780,N_29659,N_29835);
nor UO_781 (O_781,N_29098,N_29451);
nor UO_782 (O_782,N_28843,N_28928);
nand UO_783 (O_783,N_29376,N_29219);
nand UO_784 (O_784,N_28563,N_28863);
nand UO_785 (O_785,N_28796,N_28967);
nor UO_786 (O_786,N_29467,N_29942);
nand UO_787 (O_787,N_28925,N_28555);
nand UO_788 (O_788,N_28763,N_28979);
xor UO_789 (O_789,N_29437,N_28669);
nand UO_790 (O_790,N_28745,N_29552);
xor UO_791 (O_791,N_28538,N_29500);
or UO_792 (O_792,N_29284,N_29332);
or UO_793 (O_793,N_29947,N_29388);
nand UO_794 (O_794,N_28718,N_29756);
or UO_795 (O_795,N_29556,N_28835);
and UO_796 (O_796,N_28920,N_29885);
and UO_797 (O_797,N_28559,N_28906);
xnor UO_798 (O_798,N_28703,N_28898);
xor UO_799 (O_799,N_29140,N_29943);
nand UO_800 (O_800,N_29941,N_28682);
xnor UO_801 (O_801,N_29185,N_29837);
and UO_802 (O_802,N_29563,N_28769);
or UO_803 (O_803,N_28818,N_28757);
nand UO_804 (O_804,N_29426,N_29685);
or UO_805 (O_805,N_29154,N_29325);
xor UO_806 (O_806,N_28969,N_29197);
and UO_807 (O_807,N_29299,N_28554);
xnor UO_808 (O_808,N_29812,N_29250);
and UO_809 (O_809,N_29739,N_28909);
and UO_810 (O_810,N_29855,N_29682);
nand UO_811 (O_811,N_29613,N_29601);
and UO_812 (O_812,N_29696,N_29122);
xnor UO_813 (O_813,N_29852,N_29926);
nand UO_814 (O_814,N_28521,N_28631);
xnor UO_815 (O_815,N_28796,N_28885);
xnor UO_816 (O_816,N_29504,N_28973);
or UO_817 (O_817,N_29393,N_29963);
and UO_818 (O_818,N_29427,N_28538);
nor UO_819 (O_819,N_29158,N_29500);
nor UO_820 (O_820,N_29072,N_29027);
and UO_821 (O_821,N_29925,N_29534);
nand UO_822 (O_822,N_29185,N_29502);
nand UO_823 (O_823,N_29581,N_29895);
xor UO_824 (O_824,N_29379,N_29555);
and UO_825 (O_825,N_29790,N_29133);
nor UO_826 (O_826,N_28677,N_28935);
or UO_827 (O_827,N_28804,N_29469);
nor UO_828 (O_828,N_28916,N_29178);
nand UO_829 (O_829,N_29893,N_28901);
nand UO_830 (O_830,N_29168,N_28629);
xor UO_831 (O_831,N_28629,N_29680);
nand UO_832 (O_832,N_29608,N_29668);
or UO_833 (O_833,N_28934,N_29108);
or UO_834 (O_834,N_29799,N_29056);
and UO_835 (O_835,N_29915,N_29804);
nor UO_836 (O_836,N_29779,N_28836);
nand UO_837 (O_837,N_29150,N_29999);
xnor UO_838 (O_838,N_29008,N_28739);
nor UO_839 (O_839,N_28937,N_29539);
nor UO_840 (O_840,N_29618,N_28799);
or UO_841 (O_841,N_28503,N_29016);
and UO_842 (O_842,N_29858,N_29184);
xnor UO_843 (O_843,N_28996,N_29078);
xnor UO_844 (O_844,N_28505,N_29894);
xor UO_845 (O_845,N_29889,N_29597);
or UO_846 (O_846,N_29219,N_28522);
xnor UO_847 (O_847,N_29235,N_29421);
and UO_848 (O_848,N_28797,N_28503);
nor UO_849 (O_849,N_29087,N_28904);
and UO_850 (O_850,N_29774,N_28984);
and UO_851 (O_851,N_29829,N_29508);
nand UO_852 (O_852,N_29218,N_28792);
or UO_853 (O_853,N_28729,N_28744);
nor UO_854 (O_854,N_28580,N_28838);
xor UO_855 (O_855,N_28787,N_29049);
or UO_856 (O_856,N_29231,N_29073);
nor UO_857 (O_857,N_29466,N_29825);
xnor UO_858 (O_858,N_28836,N_28730);
nand UO_859 (O_859,N_29018,N_29447);
nor UO_860 (O_860,N_29851,N_29601);
and UO_861 (O_861,N_29011,N_28954);
nand UO_862 (O_862,N_28539,N_29823);
nor UO_863 (O_863,N_29102,N_29886);
and UO_864 (O_864,N_29321,N_28853);
nor UO_865 (O_865,N_29805,N_29453);
and UO_866 (O_866,N_28875,N_28979);
or UO_867 (O_867,N_28594,N_28509);
nand UO_868 (O_868,N_28556,N_28803);
xnor UO_869 (O_869,N_28511,N_28862);
nand UO_870 (O_870,N_28852,N_28960);
xnor UO_871 (O_871,N_29782,N_28932);
xnor UO_872 (O_872,N_28519,N_29123);
or UO_873 (O_873,N_29828,N_29135);
or UO_874 (O_874,N_29000,N_29304);
nand UO_875 (O_875,N_28752,N_28521);
and UO_876 (O_876,N_28811,N_29800);
and UO_877 (O_877,N_29776,N_29818);
nand UO_878 (O_878,N_29319,N_29154);
and UO_879 (O_879,N_28973,N_29298);
and UO_880 (O_880,N_29896,N_29088);
xor UO_881 (O_881,N_29558,N_29653);
nor UO_882 (O_882,N_29018,N_29165);
and UO_883 (O_883,N_28964,N_29429);
and UO_884 (O_884,N_28654,N_28677);
xor UO_885 (O_885,N_29119,N_28643);
or UO_886 (O_886,N_28945,N_29647);
nor UO_887 (O_887,N_29692,N_28955);
nor UO_888 (O_888,N_29650,N_28629);
or UO_889 (O_889,N_29176,N_29587);
nor UO_890 (O_890,N_29433,N_29134);
and UO_891 (O_891,N_28877,N_29438);
and UO_892 (O_892,N_29481,N_29475);
xor UO_893 (O_893,N_28500,N_29986);
and UO_894 (O_894,N_29319,N_29914);
and UO_895 (O_895,N_29840,N_28660);
nand UO_896 (O_896,N_29127,N_29312);
nand UO_897 (O_897,N_29291,N_28574);
nand UO_898 (O_898,N_29159,N_28524);
nor UO_899 (O_899,N_29703,N_28992);
and UO_900 (O_900,N_28967,N_29645);
nor UO_901 (O_901,N_28717,N_29140);
xnor UO_902 (O_902,N_29725,N_29852);
and UO_903 (O_903,N_29153,N_29793);
nor UO_904 (O_904,N_28581,N_29807);
nor UO_905 (O_905,N_29057,N_29431);
xnor UO_906 (O_906,N_28814,N_29084);
nor UO_907 (O_907,N_28881,N_28839);
and UO_908 (O_908,N_28612,N_29568);
or UO_909 (O_909,N_29496,N_29138);
and UO_910 (O_910,N_29841,N_28832);
xnor UO_911 (O_911,N_29713,N_29226);
nor UO_912 (O_912,N_29158,N_29684);
and UO_913 (O_913,N_29583,N_29167);
or UO_914 (O_914,N_28533,N_29108);
and UO_915 (O_915,N_28563,N_28700);
nor UO_916 (O_916,N_28530,N_29716);
xor UO_917 (O_917,N_29028,N_28794);
xnor UO_918 (O_918,N_28725,N_29366);
and UO_919 (O_919,N_28771,N_29302);
or UO_920 (O_920,N_28570,N_28875);
and UO_921 (O_921,N_28569,N_29520);
and UO_922 (O_922,N_29778,N_29230);
xnor UO_923 (O_923,N_28701,N_29787);
nand UO_924 (O_924,N_29832,N_28753);
and UO_925 (O_925,N_29301,N_28900);
xnor UO_926 (O_926,N_28714,N_28503);
nand UO_927 (O_927,N_29232,N_28568);
nand UO_928 (O_928,N_29694,N_28975);
nand UO_929 (O_929,N_29513,N_29257);
nand UO_930 (O_930,N_29627,N_29831);
nor UO_931 (O_931,N_29821,N_29767);
or UO_932 (O_932,N_29218,N_29389);
nand UO_933 (O_933,N_29997,N_29235);
nor UO_934 (O_934,N_29217,N_28569);
and UO_935 (O_935,N_29305,N_29201);
xnor UO_936 (O_936,N_29319,N_29758);
nand UO_937 (O_937,N_29518,N_29393);
and UO_938 (O_938,N_28689,N_29107);
or UO_939 (O_939,N_28516,N_29090);
or UO_940 (O_940,N_28803,N_29580);
or UO_941 (O_941,N_28928,N_29426);
or UO_942 (O_942,N_29317,N_28849);
or UO_943 (O_943,N_29598,N_28699);
nand UO_944 (O_944,N_29930,N_28942);
and UO_945 (O_945,N_29255,N_29277);
xnor UO_946 (O_946,N_29411,N_29382);
and UO_947 (O_947,N_29029,N_28961);
and UO_948 (O_948,N_28777,N_29898);
and UO_949 (O_949,N_29752,N_29548);
nor UO_950 (O_950,N_28775,N_29524);
nor UO_951 (O_951,N_29309,N_29008);
and UO_952 (O_952,N_29606,N_29885);
nor UO_953 (O_953,N_29454,N_28818);
xnor UO_954 (O_954,N_28722,N_29148);
or UO_955 (O_955,N_29143,N_29518);
xnor UO_956 (O_956,N_29896,N_28608);
nand UO_957 (O_957,N_29830,N_29903);
or UO_958 (O_958,N_29964,N_28537);
nor UO_959 (O_959,N_29186,N_29469);
and UO_960 (O_960,N_29572,N_28781);
nor UO_961 (O_961,N_29136,N_28807);
and UO_962 (O_962,N_29718,N_28555);
and UO_963 (O_963,N_29872,N_28853);
and UO_964 (O_964,N_29429,N_29576);
or UO_965 (O_965,N_28665,N_29013);
and UO_966 (O_966,N_29103,N_28984);
nor UO_967 (O_967,N_28646,N_29587);
nor UO_968 (O_968,N_28546,N_28926);
nor UO_969 (O_969,N_29283,N_28585);
or UO_970 (O_970,N_29236,N_29844);
nor UO_971 (O_971,N_28843,N_28912);
xnor UO_972 (O_972,N_29203,N_29841);
xnor UO_973 (O_973,N_29439,N_29829);
nor UO_974 (O_974,N_28990,N_29516);
xor UO_975 (O_975,N_28678,N_29915);
xor UO_976 (O_976,N_29676,N_28650);
xnor UO_977 (O_977,N_28866,N_28874);
xor UO_978 (O_978,N_29688,N_29426);
and UO_979 (O_979,N_28870,N_29345);
or UO_980 (O_980,N_28755,N_29917);
nand UO_981 (O_981,N_28724,N_29706);
and UO_982 (O_982,N_29108,N_29116);
nand UO_983 (O_983,N_29610,N_28574);
nor UO_984 (O_984,N_29682,N_29055);
nand UO_985 (O_985,N_28924,N_28688);
and UO_986 (O_986,N_29027,N_29879);
or UO_987 (O_987,N_29472,N_28633);
or UO_988 (O_988,N_29434,N_29888);
or UO_989 (O_989,N_29106,N_29344);
or UO_990 (O_990,N_29777,N_28627);
and UO_991 (O_991,N_28903,N_29611);
or UO_992 (O_992,N_28741,N_29320);
or UO_993 (O_993,N_29671,N_28859);
xnor UO_994 (O_994,N_29416,N_29271);
and UO_995 (O_995,N_29180,N_29800);
nor UO_996 (O_996,N_29369,N_28971);
nor UO_997 (O_997,N_28724,N_29878);
nor UO_998 (O_998,N_29755,N_29983);
nand UO_999 (O_999,N_29145,N_29488);
xor UO_1000 (O_1000,N_28973,N_29583);
nand UO_1001 (O_1001,N_28530,N_29003);
nand UO_1002 (O_1002,N_29563,N_28815);
or UO_1003 (O_1003,N_29254,N_29393);
xnor UO_1004 (O_1004,N_29854,N_29123);
xor UO_1005 (O_1005,N_28788,N_29780);
nand UO_1006 (O_1006,N_28649,N_28954);
xor UO_1007 (O_1007,N_29727,N_29624);
or UO_1008 (O_1008,N_28811,N_29723);
xor UO_1009 (O_1009,N_28992,N_28842);
nand UO_1010 (O_1010,N_29539,N_29995);
xor UO_1011 (O_1011,N_28862,N_29271);
nor UO_1012 (O_1012,N_29660,N_28684);
xnor UO_1013 (O_1013,N_29675,N_29063);
or UO_1014 (O_1014,N_29218,N_29410);
or UO_1015 (O_1015,N_29503,N_28847);
nor UO_1016 (O_1016,N_28736,N_28726);
xnor UO_1017 (O_1017,N_28541,N_29496);
nor UO_1018 (O_1018,N_28882,N_28557);
or UO_1019 (O_1019,N_29135,N_29988);
xnor UO_1020 (O_1020,N_29921,N_29404);
or UO_1021 (O_1021,N_29190,N_29415);
nor UO_1022 (O_1022,N_29578,N_28723);
xnor UO_1023 (O_1023,N_28974,N_29714);
or UO_1024 (O_1024,N_29515,N_29454);
and UO_1025 (O_1025,N_29717,N_28516);
nor UO_1026 (O_1026,N_29110,N_29269);
and UO_1027 (O_1027,N_28829,N_29068);
or UO_1028 (O_1028,N_28627,N_29401);
nor UO_1029 (O_1029,N_29777,N_29674);
nor UO_1030 (O_1030,N_29361,N_29902);
nor UO_1031 (O_1031,N_28625,N_29680);
and UO_1032 (O_1032,N_29388,N_29515);
or UO_1033 (O_1033,N_29712,N_28778);
or UO_1034 (O_1034,N_29978,N_29119);
nor UO_1035 (O_1035,N_29143,N_29340);
or UO_1036 (O_1036,N_29674,N_28638);
or UO_1037 (O_1037,N_28759,N_29231);
xor UO_1038 (O_1038,N_29723,N_28798);
nand UO_1039 (O_1039,N_29471,N_28789);
or UO_1040 (O_1040,N_29104,N_28954);
xnor UO_1041 (O_1041,N_28500,N_29106);
nor UO_1042 (O_1042,N_28922,N_29193);
and UO_1043 (O_1043,N_28696,N_29424);
nor UO_1044 (O_1044,N_29671,N_29213);
xor UO_1045 (O_1045,N_29707,N_29764);
or UO_1046 (O_1046,N_29239,N_29045);
and UO_1047 (O_1047,N_29413,N_28548);
nand UO_1048 (O_1048,N_29895,N_29978);
and UO_1049 (O_1049,N_29669,N_29923);
xor UO_1050 (O_1050,N_28702,N_29266);
and UO_1051 (O_1051,N_29205,N_28921);
or UO_1052 (O_1052,N_29427,N_29088);
nor UO_1053 (O_1053,N_29591,N_29056);
or UO_1054 (O_1054,N_29913,N_29849);
or UO_1055 (O_1055,N_29785,N_28530);
xor UO_1056 (O_1056,N_29285,N_29846);
and UO_1057 (O_1057,N_28667,N_29405);
nand UO_1058 (O_1058,N_28619,N_28513);
xor UO_1059 (O_1059,N_29314,N_29414);
or UO_1060 (O_1060,N_28814,N_29710);
nand UO_1061 (O_1061,N_29539,N_29692);
nand UO_1062 (O_1062,N_28679,N_28844);
nor UO_1063 (O_1063,N_29540,N_29439);
or UO_1064 (O_1064,N_29786,N_29105);
xor UO_1065 (O_1065,N_28635,N_28933);
or UO_1066 (O_1066,N_28601,N_28796);
nor UO_1067 (O_1067,N_29676,N_29825);
nor UO_1068 (O_1068,N_29390,N_28888);
xor UO_1069 (O_1069,N_28734,N_29337);
xor UO_1070 (O_1070,N_29905,N_29748);
nor UO_1071 (O_1071,N_28741,N_29246);
xor UO_1072 (O_1072,N_28844,N_29521);
nand UO_1073 (O_1073,N_28845,N_29286);
or UO_1074 (O_1074,N_29730,N_29868);
or UO_1075 (O_1075,N_29305,N_29784);
xnor UO_1076 (O_1076,N_28816,N_28582);
xor UO_1077 (O_1077,N_28726,N_29602);
and UO_1078 (O_1078,N_29001,N_29781);
and UO_1079 (O_1079,N_29911,N_29318);
and UO_1080 (O_1080,N_29631,N_29119);
or UO_1081 (O_1081,N_29587,N_29184);
and UO_1082 (O_1082,N_29203,N_29714);
xor UO_1083 (O_1083,N_29059,N_29140);
xnor UO_1084 (O_1084,N_29873,N_28659);
and UO_1085 (O_1085,N_29619,N_29069);
nand UO_1086 (O_1086,N_29109,N_29157);
nand UO_1087 (O_1087,N_28988,N_29919);
or UO_1088 (O_1088,N_29374,N_29931);
xnor UO_1089 (O_1089,N_28742,N_28908);
or UO_1090 (O_1090,N_28931,N_29441);
nor UO_1091 (O_1091,N_28760,N_28814);
and UO_1092 (O_1092,N_28804,N_29850);
or UO_1093 (O_1093,N_28517,N_28730);
nand UO_1094 (O_1094,N_28866,N_29986);
nand UO_1095 (O_1095,N_28548,N_29341);
nor UO_1096 (O_1096,N_29566,N_29034);
or UO_1097 (O_1097,N_28502,N_29881);
or UO_1098 (O_1098,N_29484,N_28690);
xor UO_1099 (O_1099,N_28945,N_29294);
and UO_1100 (O_1100,N_29476,N_29394);
nand UO_1101 (O_1101,N_28993,N_28938);
and UO_1102 (O_1102,N_29941,N_28693);
and UO_1103 (O_1103,N_29637,N_29318);
nand UO_1104 (O_1104,N_29847,N_28788);
or UO_1105 (O_1105,N_28522,N_29656);
xnor UO_1106 (O_1106,N_28503,N_29125);
or UO_1107 (O_1107,N_29313,N_29788);
xnor UO_1108 (O_1108,N_29631,N_29189);
xor UO_1109 (O_1109,N_29460,N_28675);
xnor UO_1110 (O_1110,N_28926,N_29130);
and UO_1111 (O_1111,N_29730,N_28986);
xor UO_1112 (O_1112,N_28821,N_29664);
or UO_1113 (O_1113,N_29558,N_29320);
nor UO_1114 (O_1114,N_28609,N_28685);
and UO_1115 (O_1115,N_28520,N_28688);
xnor UO_1116 (O_1116,N_29267,N_28961);
nor UO_1117 (O_1117,N_29285,N_29323);
or UO_1118 (O_1118,N_29859,N_28527);
nand UO_1119 (O_1119,N_28906,N_29505);
nand UO_1120 (O_1120,N_29814,N_29083);
nor UO_1121 (O_1121,N_29785,N_29331);
or UO_1122 (O_1122,N_28768,N_28621);
xnor UO_1123 (O_1123,N_28570,N_29685);
and UO_1124 (O_1124,N_29177,N_28906);
and UO_1125 (O_1125,N_29488,N_29892);
or UO_1126 (O_1126,N_28656,N_29114);
and UO_1127 (O_1127,N_29647,N_28698);
or UO_1128 (O_1128,N_28942,N_28759);
nand UO_1129 (O_1129,N_29494,N_28800);
xnor UO_1130 (O_1130,N_29079,N_29659);
nor UO_1131 (O_1131,N_29681,N_28623);
or UO_1132 (O_1132,N_29411,N_29541);
nor UO_1133 (O_1133,N_29870,N_29034);
and UO_1134 (O_1134,N_29779,N_29006);
and UO_1135 (O_1135,N_28500,N_29079);
nor UO_1136 (O_1136,N_28634,N_29538);
nor UO_1137 (O_1137,N_29964,N_28632);
and UO_1138 (O_1138,N_28802,N_29078);
nor UO_1139 (O_1139,N_28785,N_29132);
and UO_1140 (O_1140,N_29794,N_29439);
and UO_1141 (O_1141,N_29524,N_29160);
nand UO_1142 (O_1142,N_28736,N_28724);
xnor UO_1143 (O_1143,N_29365,N_29683);
nor UO_1144 (O_1144,N_29621,N_29609);
xor UO_1145 (O_1145,N_29695,N_28770);
xor UO_1146 (O_1146,N_28576,N_29353);
or UO_1147 (O_1147,N_29223,N_29135);
nor UO_1148 (O_1148,N_29963,N_29919);
nand UO_1149 (O_1149,N_29920,N_29280);
or UO_1150 (O_1150,N_28706,N_29515);
xnor UO_1151 (O_1151,N_29575,N_29451);
nand UO_1152 (O_1152,N_29759,N_28713);
and UO_1153 (O_1153,N_29509,N_29520);
xor UO_1154 (O_1154,N_28850,N_29712);
nor UO_1155 (O_1155,N_28594,N_28600);
xnor UO_1156 (O_1156,N_29488,N_29890);
nand UO_1157 (O_1157,N_28564,N_29723);
nand UO_1158 (O_1158,N_29197,N_29672);
and UO_1159 (O_1159,N_29967,N_29423);
or UO_1160 (O_1160,N_29161,N_28558);
nand UO_1161 (O_1161,N_29119,N_28687);
and UO_1162 (O_1162,N_29974,N_29287);
nand UO_1163 (O_1163,N_29365,N_29222);
and UO_1164 (O_1164,N_29773,N_29860);
nor UO_1165 (O_1165,N_29957,N_28510);
nand UO_1166 (O_1166,N_28592,N_28579);
nand UO_1167 (O_1167,N_28718,N_28858);
nand UO_1168 (O_1168,N_29434,N_28812);
and UO_1169 (O_1169,N_29307,N_28661);
xor UO_1170 (O_1170,N_28543,N_28529);
and UO_1171 (O_1171,N_29270,N_28894);
and UO_1172 (O_1172,N_29916,N_29597);
nand UO_1173 (O_1173,N_29691,N_28959);
xnor UO_1174 (O_1174,N_29964,N_29179);
nand UO_1175 (O_1175,N_29707,N_29637);
xnor UO_1176 (O_1176,N_29090,N_28940);
nand UO_1177 (O_1177,N_28535,N_29354);
nor UO_1178 (O_1178,N_29712,N_29744);
or UO_1179 (O_1179,N_29884,N_28518);
xnor UO_1180 (O_1180,N_29408,N_29722);
nor UO_1181 (O_1181,N_29092,N_29752);
nand UO_1182 (O_1182,N_29851,N_29792);
and UO_1183 (O_1183,N_28770,N_28932);
xnor UO_1184 (O_1184,N_29199,N_29338);
and UO_1185 (O_1185,N_29104,N_29782);
nand UO_1186 (O_1186,N_28965,N_29697);
or UO_1187 (O_1187,N_29094,N_29036);
or UO_1188 (O_1188,N_29178,N_28509);
and UO_1189 (O_1189,N_28787,N_28655);
nor UO_1190 (O_1190,N_29294,N_28580);
nand UO_1191 (O_1191,N_28794,N_29725);
xnor UO_1192 (O_1192,N_28969,N_29738);
or UO_1193 (O_1193,N_29419,N_29878);
nor UO_1194 (O_1194,N_28778,N_29380);
nor UO_1195 (O_1195,N_29802,N_29005);
nor UO_1196 (O_1196,N_29494,N_28956);
nand UO_1197 (O_1197,N_28615,N_29849);
nand UO_1198 (O_1198,N_29299,N_29363);
nor UO_1199 (O_1199,N_29540,N_29415);
nand UO_1200 (O_1200,N_29026,N_29324);
nor UO_1201 (O_1201,N_28588,N_28517);
nor UO_1202 (O_1202,N_29033,N_28800);
and UO_1203 (O_1203,N_29105,N_28891);
nand UO_1204 (O_1204,N_29786,N_29856);
or UO_1205 (O_1205,N_29091,N_29272);
xnor UO_1206 (O_1206,N_28634,N_29675);
and UO_1207 (O_1207,N_29310,N_29379);
nand UO_1208 (O_1208,N_29329,N_29428);
and UO_1209 (O_1209,N_28948,N_29924);
nor UO_1210 (O_1210,N_28966,N_28908);
and UO_1211 (O_1211,N_29927,N_29300);
xnor UO_1212 (O_1212,N_29338,N_29119);
and UO_1213 (O_1213,N_29534,N_28600);
nand UO_1214 (O_1214,N_28690,N_29605);
nor UO_1215 (O_1215,N_29619,N_29180);
nor UO_1216 (O_1216,N_28871,N_29511);
nor UO_1217 (O_1217,N_28777,N_28554);
and UO_1218 (O_1218,N_29172,N_29742);
and UO_1219 (O_1219,N_29464,N_28567);
and UO_1220 (O_1220,N_29455,N_28610);
nand UO_1221 (O_1221,N_28792,N_29882);
or UO_1222 (O_1222,N_29216,N_28585);
xor UO_1223 (O_1223,N_29250,N_29847);
xor UO_1224 (O_1224,N_29363,N_29423);
or UO_1225 (O_1225,N_29770,N_29806);
xnor UO_1226 (O_1226,N_29280,N_28527);
and UO_1227 (O_1227,N_29077,N_29720);
nor UO_1228 (O_1228,N_28596,N_29984);
xnor UO_1229 (O_1229,N_29396,N_28581);
or UO_1230 (O_1230,N_29432,N_28894);
or UO_1231 (O_1231,N_28750,N_28862);
xor UO_1232 (O_1232,N_28802,N_28701);
or UO_1233 (O_1233,N_29191,N_29858);
nor UO_1234 (O_1234,N_28557,N_29970);
xor UO_1235 (O_1235,N_29869,N_28917);
and UO_1236 (O_1236,N_28813,N_28852);
xnor UO_1237 (O_1237,N_29507,N_28661);
nand UO_1238 (O_1238,N_28565,N_28850);
nand UO_1239 (O_1239,N_28741,N_29210);
and UO_1240 (O_1240,N_28513,N_29715);
nand UO_1241 (O_1241,N_28870,N_28770);
nand UO_1242 (O_1242,N_29631,N_28846);
xnor UO_1243 (O_1243,N_29766,N_29956);
nor UO_1244 (O_1244,N_28689,N_28939);
or UO_1245 (O_1245,N_29916,N_29918);
or UO_1246 (O_1246,N_28674,N_28920);
xor UO_1247 (O_1247,N_29919,N_29566);
nand UO_1248 (O_1248,N_28913,N_29084);
nand UO_1249 (O_1249,N_29104,N_28827);
or UO_1250 (O_1250,N_29204,N_28927);
nand UO_1251 (O_1251,N_29148,N_28835);
nor UO_1252 (O_1252,N_28799,N_28540);
xor UO_1253 (O_1253,N_28728,N_29189);
xor UO_1254 (O_1254,N_29076,N_29948);
nor UO_1255 (O_1255,N_28616,N_28918);
and UO_1256 (O_1256,N_29584,N_28518);
nor UO_1257 (O_1257,N_29975,N_29789);
nor UO_1258 (O_1258,N_29641,N_29657);
nor UO_1259 (O_1259,N_29273,N_29565);
xor UO_1260 (O_1260,N_29017,N_29099);
xnor UO_1261 (O_1261,N_29057,N_29347);
nand UO_1262 (O_1262,N_28502,N_29070);
nand UO_1263 (O_1263,N_29705,N_29629);
and UO_1264 (O_1264,N_29021,N_29315);
xor UO_1265 (O_1265,N_28806,N_29985);
nor UO_1266 (O_1266,N_29354,N_28761);
nor UO_1267 (O_1267,N_29619,N_29534);
nand UO_1268 (O_1268,N_29876,N_29642);
nand UO_1269 (O_1269,N_29211,N_28789);
nor UO_1270 (O_1270,N_29089,N_29787);
xnor UO_1271 (O_1271,N_29163,N_28624);
nor UO_1272 (O_1272,N_28756,N_28563);
nor UO_1273 (O_1273,N_29355,N_29738);
nand UO_1274 (O_1274,N_28969,N_29564);
xor UO_1275 (O_1275,N_29296,N_29353);
or UO_1276 (O_1276,N_28891,N_28903);
xor UO_1277 (O_1277,N_29104,N_28956);
nor UO_1278 (O_1278,N_28768,N_28911);
and UO_1279 (O_1279,N_28670,N_29710);
and UO_1280 (O_1280,N_29287,N_28725);
xor UO_1281 (O_1281,N_29228,N_29977);
nand UO_1282 (O_1282,N_29387,N_29084);
nor UO_1283 (O_1283,N_28935,N_28771);
xor UO_1284 (O_1284,N_29249,N_29299);
nand UO_1285 (O_1285,N_28535,N_29513);
and UO_1286 (O_1286,N_29872,N_29117);
nor UO_1287 (O_1287,N_29891,N_28733);
nor UO_1288 (O_1288,N_29317,N_28774);
xnor UO_1289 (O_1289,N_29439,N_29176);
xnor UO_1290 (O_1290,N_29841,N_28720);
and UO_1291 (O_1291,N_29011,N_28649);
or UO_1292 (O_1292,N_29178,N_29843);
nor UO_1293 (O_1293,N_29703,N_29002);
nand UO_1294 (O_1294,N_29737,N_29022);
or UO_1295 (O_1295,N_28711,N_29971);
nand UO_1296 (O_1296,N_28777,N_29718);
xnor UO_1297 (O_1297,N_29120,N_29459);
xor UO_1298 (O_1298,N_29025,N_29365);
nand UO_1299 (O_1299,N_29190,N_29201);
or UO_1300 (O_1300,N_28595,N_28747);
and UO_1301 (O_1301,N_29657,N_29782);
nor UO_1302 (O_1302,N_29654,N_29313);
xnor UO_1303 (O_1303,N_29888,N_29372);
and UO_1304 (O_1304,N_29776,N_29369);
xnor UO_1305 (O_1305,N_29386,N_29208);
nor UO_1306 (O_1306,N_28707,N_29261);
nor UO_1307 (O_1307,N_29805,N_28738);
nand UO_1308 (O_1308,N_29760,N_29665);
and UO_1309 (O_1309,N_29270,N_29439);
xnor UO_1310 (O_1310,N_29964,N_29892);
xnor UO_1311 (O_1311,N_29233,N_29206);
and UO_1312 (O_1312,N_29697,N_29740);
xor UO_1313 (O_1313,N_29816,N_29798);
xor UO_1314 (O_1314,N_29997,N_28947);
and UO_1315 (O_1315,N_29863,N_29806);
nand UO_1316 (O_1316,N_29589,N_29196);
nand UO_1317 (O_1317,N_28608,N_28677);
xnor UO_1318 (O_1318,N_29635,N_29233);
nand UO_1319 (O_1319,N_28590,N_29492);
or UO_1320 (O_1320,N_29997,N_29355);
xor UO_1321 (O_1321,N_28802,N_29853);
nand UO_1322 (O_1322,N_28982,N_29769);
nor UO_1323 (O_1323,N_28838,N_29768);
xor UO_1324 (O_1324,N_28866,N_28554);
xnor UO_1325 (O_1325,N_29009,N_29016);
or UO_1326 (O_1326,N_29202,N_28779);
xor UO_1327 (O_1327,N_28654,N_28811);
or UO_1328 (O_1328,N_28937,N_29760);
nor UO_1329 (O_1329,N_29693,N_28589);
nand UO_1330 (O_1330,N_28732,N_28947);
nor UO_1331 (O_1331,N_28515,N_29087);
and UO_1332 (O_1332,N_28997,N_28814);
xnor UO_1333 (O_1333,N_29150,N_29056);
and UO_1334 (O_1334,N_29702,N_29843);
nor UO_1335 (O_1335,N_29558,N_29702);
nor UO_1336 (O_1336,N_29815,N_29131);
nand UO_1337 (O_1337,N_29311,N_29431);
or UO_1338 (O_1338,N_29628,N_29246);
and UO_1339 (O_1339,N_29704,N_29455);
and UO_1340 (O_1340,N_29960,N_29942);
or UO_1341 (O_1341,N_29403,N_29971);
xor UO_1342 (O_1342,N_29789,N_29381);
nand UO_1343 (O_1343,N_28678,N_29568);
or UO_1344 (O_1344,N_29167,N_28516);
and UO_1345 (O_1345,N_29658,N_29564);
nor UO_1346 (O_1346,N_29194,N_28863);
nor UO_1347 (O_1347,N_29207,N_29399);
nand UO_1348 (O_1348,N_29585,N_29507);
and UO_1349 (O_1349,N_29567,N_28851);
xor UO_1350 (O_1350,N_29514,N_28640);
and UO_1351 (O_1351,N_29487,N_29361);
or UO_1352 (O_1352,N_29713,N_29448);
and UO_1353 (O_1353,N_28720,N_29410);
nor UO_1354 (O_1354,N_29178,N_29601);
nor UO_1355 (O_1355,N_29708,N_28536);
nor UO_1356 (O_1356,N_29726,N_29665);
or UO_1357 (O_1357,N_29746,N_29753);
xor UO_1358 (O_1358,N_28746,N_29236);
and UO_1359 (O_1359,N_28601,N_29418);
nand UO_1360 (O_1360,N_29470,N_28846);
xor UO_1361 (O_1361,N_28923,N_29206);
or UO_1362 (O_1362,N_29365,N_28617);
nand UO_1363 (O_1363,N_29001,N_29807);
nand UO_1364 (O_1364,N_29767,N_28946);
or UO_1365 (O_1365,N_29652,N_29919);
and UO_1366 (O_1366,N_29988,N_29387);
xor UO_1367 (O_1367,N_28983,N_29630);
or UO_1368 (O_1368,N_29624,N_29633);
and UO_1369 (O_1369,N_29108,N_28813);
and UO_1370 (O_1370,N_28684,N_29045);
and UO_1371 (O_1371,N_29897,N_29108);
xnor UO_1372 (O_1372,N_28584,N_29855);
nand UO_1373 (O_1373,N_29661,N_29051);
and UO_1374 (O_1374,N_29409,N_29291);
and UO_1375 (O_1375,N_29626,N_29462);
xor UO_1376 (O_1376,N_29778,N_29135);
xnor UO_1377 (O_1377,N_28790,N_29935);
xor UO_1378 (O_1378,N_29256,N_29102);
nor UO_1379 (O_1379,N_28554,N_29118);
xor UO_1380 (O_1380,N_28747,N_29355);
and UO_1381 (O_1381,N_29058,N_29188);
xnor UO_1382 (O_1382,N_29813,N_29164);
or UO_1383 (O_1383,N_29099,N_28949);
nand UO_1384 (O_1384,N_29626,N_28659);
xor UO_1385 (O_1385,N_28757,N_29435);
nand UO_1386 (O_1386,N_28532,N_28920);
xnor UO_1387 (O_1387,N_29590,N_29484);
or UO_1388 (O_1388,N_29633,N_28979);
nand UO_1389 (O_1389,N_29702,N_28502);
nor UO_1390 (O_1390,N_29714,N_29703);
or UO_1391 (O_1391,N_28580,N_28695);
nand UO_1392 (O_1392,N_29991,N_29319);
nor UO_1393 (O_1393,N_29226,N_29214);
and UO_1394 (O_1394,N_29350,N_29853);
and UO_1395 (O_1395,N_28776,N_29221);
nand UO_1396 (O_1396,N_28920,N_29835);
or UO_1397 (O_1397,N_29682,N_29111);
nor UO_1398 (O_1398,N_28757,N_28572);
nand UO_1399 (O_1399,N_28581,N_29634);
nor UO_1400 (O_1400,N_29578,N_29673);
and UO_1401 (O_1401,N_29976,N_29376);
nand UO_1402 (O_1402,N_29052,N_29389);
nand UO_1403 (O_1403,N_29622,N_28534);
or UO_1404 (O_1404,N_28979,N_29088);
nand UO_1405 (O_1405,N_29753,N_28733);
nand UO_1406 (O_1406,N_29614,N_29212);
or UO_1407 (O_1407,N_29647,N_29862);
nor UO_1408 (O_1408,N_29780,N_28828);
nor UO_1409 (O_1409,N_29961,N_29741);
nor UO_1410 (O_1410,N_29057,N_28842);
nor UO_1411 (O_1411,N_29296,N_28622);
nand UO_1412 (O_1412,N_28726,N_29892);
xnor UO_1413 (O_1413,N_29641,N_28606);
and UO_1414 (O_1414,N_29833,N_29469);
nand UO_1415 (O_1415,N_29048,N_29952);
and UO_1416 (O_1416,N_29449,N_29292);
or UO_1417 (O_1417,N_28823,N_28935);
nor UO_1418 (O_1418,N_29899,N_28502);
nor UO_1419 (O_1419,N_28895,N_29871);
nor UO_1420 (O_1420,N_29064,N_28721);
nor UO_1421 (O_1421,N_29602,N_29303);
nand UO_1422 (O_1422,N_28575,N_29456);
nand UO_1423 (O_1423,N_28918,N_29037);
nand UO_1424 (O_1424,N_29667,N_28732);
xnor UO_1425 (O_1425,N_29330,N_29595);
and UO_1426 (O_1426,N_29242,N_29256);
nand UO_1427 (O_1427,N_29004,N_29731);
xor UO_1428 (O_1428,N_29172,N_29917);
nand UO_1429 (O_1429,N_29518,N_29103);
nand UO_1430 (O_1430,N_28650,N_29401);
and UO_1431 (O_1431,N_28886,N_29427);
or UO_1432 (O_1432,N_28584,N_29340);
nor UO_1433 (O_1433,N_28617,N_29796);
nand UO_1434 (O_1434,N_29328,N_29050);
or UO_1435 (O_1435,N_29639,N_28870);
nor UO_1436 (O_1436,N_29175,N_28651);
nor UO_1437 (O_1437,N_29330,N_28787);
nor UO_1438 (O_1438,N_29411,N_28705);
or UO_1439 (O_1439,N_28984,N_29472);
nand UO_1440 (O_1440,N_28555,N_28582);
or UO_1441 (O_1441,N_28730,N_28985);
and UO_1442 (O_1442,N_29752,N_28953);
nor UO_1443 (O_1443,N_29711,N_29457);
xnor UO_1444 (O_1444,N_28866,N_29958);
nand UO_1445 (O_1445,N_29794,N_28562);
nor UO_1446 (O_1446,N_29299,N_29211);
xor UO_1447 (O_1447,N_29454,N_29125);
xor UO_1448 (O_1448,N_28984,N_28936);
and UO_1449 (O_1449,N_29070,N_29032);
or UO_1450 (O_1450,N_29148,N_29834);
nand UO_1451 (O_1451,N_29380,N_28594);
and UO_1452 (O_1452,N_29573,N_29316);
and UO_1453 (O_1453,N_29767,N_29659);
or UO_1454 (O_1454,N_29701,N_28563);
nand UO_1455 (O_1455,N_28743,N_29980);
nor UO_1456 (O_1456,N_29023,N_29076);
and UO_1457 (O_1457,N_29887,N_29924);
or UO_1458 (O_1458,N_29083,N_29638);
nor UO_1459 (O_1459,N_29036,N_28561);
nand UO_1460 (O_1460,N_28701,N_29500);
nand UO_1461 (O_1461,N_29796,N_28608);
xnor UO_1462 (O_1462,N_29663,N_28568);
and UO_1463 (O_1463,N_28764,N_28849);
xnor UO_1464 (O_1464,N_28702,N_29773);
or UO_1465 (O_1465,N_28696,N_29642);
and UO_1466 (O_1466,N_28986,N_29277);
nand UO_1467 (O_1467,N_28673,N_29772);
and UO_1468 (O_1468,N_29822,N_29783);
or UO_1469 (O_1469,N_28833,N_29133);
nand UO_1470 (O_1470,N_29330,N_28867);
nor UO_1471 (O_1471,N_28541,N_29360);
nand UO_1472 (O_1472,N_28596,N_29623);
xnor UO_1473 (O_1473,N_29231,N_28855);
nand UO_1474 (O_1474,N_29833,N_29979);
and UO_1475 (O_1475,N_29568,N_28520);
nand UO_1476 (O_1476,N_29275,N_28690);
nand UO_1477 (O_1477,N_29310,N_29627);
xor UO_1478 (O_1478,N_28551,N_29794);
and UO_1479 (O_1479,N_28990,N_28916);
xor UO_1480 (O_1480,N_29655,N_29263);
xor UO_1481 (O_1481,N_29140,N_29449);
nor UO_1482 (O_1482,N_28843,N_29821);
nor UO_1483 (O_1483,N_29292,N_29852);
nor UO_1484 (O_1484,N_29674,N_28974);
or UO_1485 (O_1485,N_29979,N_28962);
and UO_1486 (O_1486,N_28980,N_29250);
or UO_1487 (O_1487,N_28685,N_29300);
and UO_1488 (O_1488,N_29243,N_29234);
nand UO_1489 (O_1489,N_29184,N_29829);
xor UO_1490 (O_1490,N_29303,N_28566);
xnor UO_1491 (O_1491,N_29053,N_29534);
nor UO_1492 (O_1492,N_28999,N_28551);
or UO_1493 (O_1493,N_28939,N_29715);
nand UO_1494 (O_1494,N_28943,N_29942);
xnor UO_1495 (O_1495,N_28543,N_29881);
and UO_1496 (O_1496,N_28502,N_28668);
nand UO_1497 (O_1497,N_29423,N_29817);
nand UO_1498 (O_1498,N_28654,N_29526);
or UO_1499 (O_1499,N_29978,N_29821);
nor UO_1500 (O_1500,N_29841,N_29704);
xnor UO_1501 (O_1501,N_29225,N_29449);
nor UO_1502 (O_1502,N_29327,N_29954);
and UO_1503 (O_1503,N_28913,N_28730);
and UO_1504 (O_1504,N_28919,N_29710);
nand UO_1505 (O_1505,N_28867,N_29523);
nand UO_1506 (O_1506,N_29721,N_29835);
nor UO_1507 (O_1507,N_29684,N_28555);
xor UO_1508 (O_1508,N_29632,N_28681);
or UO_1509 (O_1509,N_28508,N_28913);
nor UO_1510 (O_1510,N_29488,N_29371);
nor UO_1511 (O_1511,N_29106,N_29876);
nand UO_1512 (O_1512,N_29316,N_28884);
or UO_1513 (O_1513,N_29498,N_29434);
nor UO_1514 (O_1514,N_28577,N_29811);
nor UO_1515 (O_1515,N_28522,N_28551);
or UO_1516 (O_1516,N_28866,N_29815);
xor UO_1517 (O_1517,N_29983,N_29262);
and UO_1518 (O_1518,N_28923,N_28671);
and UO_1519 (O_1519,N_28973,N_29696);
nor UO_1520 (O_1520,N_29059,N_28543);
xor UO_1521 (O_1521,N_29043,N_28566);
xnor UO_1522 (O_1522,N_29979,N_28879);
nand UO_1523 (O_1523,N_29379,N_29407);
xnor UO_1524 (O_1524,N_28920,N_29101);
xnor UO_1525 (O_1525,N_29800,N_29845);
nand UO_1526 (O_1526,N_29311,N_29736);
nor UO_1527 (O_1527,N_29913,N_29271);
xor UO_1528 (O_1528,N_28843,N_29895);
nand UO_1529 (O_1529,N_28822,N_28626);
xnor UO_1530 (O_1530,N_28836,N_29233);
xor UO_1531 (O_1531,N_28649,N_28903);
nor UO_1532 (O_1532,N_29976,N_29701);
nor UO_1533 (O_1533,N_29505,N_29429);
nand UO_1534 (O_1534,N_29465,N_28966);
or UO_1535 (O_1535,N_28819,N_29058);
and UO_1536 (O_1536,N_29210,N_29829);
nand UO_1537 (O_1537,N_28767,N_29581);
nand UO_1538 (O_1538,N_28689,N_29066);
or UO_1539 (O_1539,N_29983,N_28714);
xnor UO_1540 (O_1540,N_29384,N_29153);
nor UO_1541 (O_1541,N_29061,N_29580);
xor UO_1542 (O_1542,N_28648,N_29096);
nand UO_1543 (O_1543,N_29852,N_29551);
nor UO_1544 (O_1544,N_29314,N_29731);
or UO_1545 (O_1545,N_29633,N_28776);
nor UO_1546 (O_1546,N_29471,N_28577);
nor UO_1547 (O_1547,N_28567,N_29287);
nand UO_1548 (O_1548,N_29148,N_29150);
nand UO_1549 (O_1549,N_29347,N_29350);
nor UO_1550 (O_1550,N_29888,N_29488);
and UO_1551 (O_1551,N_29711,N_29429);
nand UO_1552 (O_1552,N_29898,N_29873);
xnor UO_1553 (O_1553,N_28533,N_29390);
and UO_1554 (O_1554,N_29126,N_29331);
or UO_1555 (O_1555,N_28860,N_29445);
xor UO_1556 (O_1556,N_29791,N_29318);
or UO_1557 (O_1557,N_29480,N_29035);
and UO_1558 (O_1558,N_29564,N_28703);
or UO_1559 (O_1559,N_29174,N_29278);
nand UO_1560 (O_1560,N_28586,N_29114);
nand UO_1561 (O_1561,N_29448,N_28685);
xor UO_1562 (O_1562,N_28676,N_29851);
and UO_1563 (O_1563,N_29871,N_28939);
nor UO_1564 (O_1564,N_29785,N_29406);
or UO_1565 (O_1565,N_28691,N_29779);
nor UO_1566 (O_1566,N_28801,N_28972);
nand UO_1567 (O_1567,N_28954,N_29929);
or UO_1568 (O_1568,N_29469,N_29533);
nor UO_1569 (O_1569,N_28764,N_29120);
xnor UO_1570 (O_1570,N_29309,N_28640);
nand UO_1571 (O_1571,N_29951,N_28850);
and UO_1572 (O_1572,N_29877,N_29645);
xor UO_1573 (O_1573,N_29724,N_29984);
and UO_1574 (O_1574,N_28964,N_29378);
nand UO_1575 (O_1575,N_29546,N_28531);
or UO_1576 (O_1576,N_28508,N_29983);
nor UO_1577 (O_1577,N_28946,N_29910);
or UO_1578 (O_1578,N_29166,N_28849);
xnor UO_1579 (O_1579,N_28702,N_29352);
and UO_1580 (O_1580,N_29889,N_29580);
and UO_1581 (O_1581,N_28623,N_28849);
nor UO_1582 (O_1582,N_29335,N_28507);
xor UO_1583 (O_1583,N_29874,N_29623);
nor UO_1584 (O_1584,N_29785,N_28507);
nor UO_1585 (O_1585,N_29048,N_28938);
and UO_1586 (O_1586,N_28502,N_28741);
nand UO_1587 (O_1587,N_29055,N_29824);
nand UO_1588 (O_1588,N_28895,N_28929);
nor UO_1589 (O_1589,N_28748,N_28560);
nor UO_1590 (O_1590,N_28653,N_29269);
or UO_1591 (O_1591,N_29594,N_29754);
xnor UO_1592 (O_1592,N_29489,N_28635);
nand UO_1593 (O_1593,N_29913,N_29687);
xor UO_1594 (O_1594,N_29646,N_28763);
nor UO_1595 (O_1595,N_28787,N_29898);
xnor UO_1596 (O_1596,N_29198,N_28678);
nor UO_1597 (O_1597,N_29114,N_29437);
nand UO_1598 (O_1598,N_29699,N_28988);
xnor UO_1599 (O_1599,N_29786,N_28706);
nand UO_1600 (O_1600,N_28518,N_29520);
nor UO_1601 (O_1601,N_28840,N_29059);
or UO_1602 (O_1602,N_29143,N_29233);
and UO_1603 (O_1603,N_29932,N_29520);
or UO_1604 (O_1604,N_28948,N_28528);
nor UO_1605 (O_1605,N_28773,N_28599);
nor UO_1606 (O_1606,N_28959,N_29979);
xnor UO_1607 (O_1607,N_29689,N_28855);
nor UO_1608 (O_1608,N_29200,N_29742);
or UO_1609 (O_1609,N_29206,N_28794);
xnor UO_1610 (O_1610,N_28524,N_28611);
nand UO_1611 (O_1611,N_29346,N_29058);
xor UO_1612 (O_1612,N_28947,N_29552);
nand UO_1613 (O_1613,N_29212,N_28972);
xnor UO_1614 (O_1614,N_28963,N_28557);
nor UO_1615 (O_1615,N_29520,N_29957);
nand UO_1616 (O_1616,N_29904,N_29290);
nand UO_1617 (O_1617,N_28877,N_29739);
nand UO_1618 (O_1618,N_29286,N_28558);
and UO_1619 (O_1619,N_28976,N_28545);
nand UO_1620 (O_1620,N_29174,N_29565);
nand UO_1621 (O_1621,N_28803,N_29679);
and UO_1622 (O_1622,N_29815,N_29303);
nor UO_1623 (O_1623,N_29616,N_29408);
or UO_1624 (O_1624,N_29175,N_29248);
nand UO_1625 (O_1625,N_29634,N_29404);
xnor UO_1626 (O_1626,N_28974,N_28964);
or UO_1627 (O_1627,N_29828,N_28660);
xor UO_1628 (O_1628,N_29813,N_28892);
nand UO_1629 (O_1629,N_28812,N_28731);
xor UO_1630 (O_1630,N_28715,N_28926);
and UO_1631 (O_1631,N_29933,N_28808);
or UO_1632 (O_1632,N_28687,N_29789);
or UO_1633 (O_1633,N_29839,N_29561);
or UO_1634 (O_1634,N_29833,N_29879);
xor UO_1635 (O_1635,N_28756,N_28890);
and UO_1636 (O_1636,N_29632,N_28638);
nand UO_1637 (O_1637,N_28796,N_29764);
nand UO_1638 (O_1638,N_29336,N_29999);
and UO_1639 (O_1639,N_29337,N_28561);
nor UO_1640 (O_1640,N_28745,N_29312);
or UO_1641 (O_1641,N_29684,N_29977);
and UO_1642 (O_1642,N_28616,N_29973);
nor UO_1643 (O_1643,N_28546,N_29570);
nor UO_1644 (O_1644,N_28851,N_29799);
xor UO_1645 (O_1645,N_29437,N_29899);
xor UO_1646 (O_1646,N_28688,N_28678);
nor UO_1647 (O_1647,N_29748,N_29792);
nor UO_1648 (O_1648,N_28618,N_28653);
and UO_1649 (O_1649,N_29140,N_29835);
and UO_1650 (O_1650,N_29953,N_28856);
and UO_1651 (O_1651,N_28994,N_28935);
xor UO_1652 (O_1652,N_29325,N_28983);
nand UO_1653 (O_1653,N_29249,N_29076);
and UO_1654 (O_1654,N_28773,N_28891);
xor UO_1655 (O_1655,N_29462,N_29255);
xnor UO_1656 (O_1656,N_28545,N_29240);
nor UO_1657 (O_1657,N_29586,N_28809);
nand UO_1658 (O_1658,N_29820,N_29406);
nand UO_1659 (O_1659,N_29079,N_29889);
or UO_1660 (O_1660,N_29858,N_29501);
or UO_1661 (O_1661,N_28675,N_28760);
xnor UO_1662 (O_1662,N_29457,N_29454);
nor UO_1663 (O_1663,N_29119,N_28842);
or UO_1664 (O_1664,N_28732,N_29949);
xor UO_1665 (O_1665,N_29181,N_28866);
and UO_1666 (O_1666,N_28825,N_29204);
nand UO_1667 (O_1667,N_28823,N_29487);
nor UO_1668 (O_1668,N_29290,N_29481);
xnor UO_1669 (O_1669,N_29479,N_29309);
and UO_1670 (O_1670,N_29692,N_29568);
nor UO_1671 (O_1671,N_29718,N_29102);
nor UO_1672 (O_1672,N_29026,N_29572);
nor UO_1673 (O_1673,N_29001,N_29586);
and UO_1674 (O_1674,N_29149,N_28939);
or UO_1675 (O_1675,N_28516,N_29702);
xor UO_1676 (O_1676,N_29238,N_28664);
nor UO_1677 (O_1677,N_29739,N_28882);
xor UO_1678 (O_1678,N_29811,N_28599);
and UO_1679 (O_1679,N_28927,N_28985);
or UO_1680 (O_1680,N_28950,N_29766);
nand UO_1681 (O_1681,N_29446,N_29316);
nand UO_1682 (O_1682,N_28708,N_29397);
nand UO_1683 (O_1683,N_28580,N_28709);
or UO_1684 (O_1684,N_28776,N_29318);
xor UO_1685 (O_1685,N_29630,N_28801);
or UO_1686 (O_1686,N_29606,N_28787);
or UO_1687 (O_1687,N_29583,N_29759);
xnor UO_1688 (O_1688,N_28800,N_29841);
and UO_1689 (O_1689,N_29947,N_29829);
nand UO_1690 (O_1690,N_29765,N_28721);
xor UO_1691 (O_1691,N_29492,N_28547);
and UO_1692 (O_1692,N_29255,N_29764);
or UO_1693 (O_1693,N_29994,N_28552);
nand UO_1694 (O_1694,N_28784,N_29244);
nand UO_1695 (O_1695,N_29579,N_29158);
and UO_1696 (O_1696,N_29321,N_29535);
nand UO_1697 (O_1697,N_29810,N_29245);
nand UO_1698 (O_1698,N_29157,N_28787);
nor UO_1699 (O_1699,N_29247,N_28645);
nand UO_1700 (O_1700,N_29971,N_29076);
or UO_1701 (O_1701,N_28934,N_29165);
nor UO_1702 (O_1702,N_29373,N_28933);
nor UO_1703 (O_1703,N_29593,N_28538);
xor UO_1704 (O_1704,N_29506,N_29381);
or UO_1705 (O_1705,N_28541,N_28583);
or UO_1706 (O_1706,N_28684,N_28631);
or UO_1707 (O_1707,N_29286,N_28534);
xor UO_1708 (O_1708,N_28878,N_29719);
nand UO_1709 (O_1709,N_29295,N_28639);
nand UO_1710 (O_1710,N_29608,N_29152);
xor UO_1711 (O_1711,N_29179,N_29524);
nand UO_1712 (O_1712,N_29390,N_29879);
nand UO_1713 (O_1713,N_29227,N_29322);
nand UO_1714 (O_1714,N_29429,N_28720);
xor UO_1715 (O_1715,N_29749,N_28942);
and UO_1716 (O_1716,N_29921,N_29177);
xnor UO_1717 (O_1717,N_29649,N_29728);
and UO_1718 (O_1718,N_29273,N_28795);
and UO_1719 (O_1719,N_29841,N_29304);
nand UO_1720 (O_1720,N_28524,N_29348);
xnor UO_1721 (O_1721,N_29819,N_28606);
or UO_1722 (O_1722,N_28624,N_28752);
xor UO_1723 (O_1723,N_29884,N_28813);
or UO_1724 (O_1724,N_28781,N_29564);
and UO_1725 (O_1725,N_29222,N_29763);
xnor UO_1726 (O_1726,N_29654,N_28741);
nor UO_1727 (O_1727,N_29663,N_28911);
nand UO_1728 (O_1728,N_28757,N_28672);
nand UO_1729 (O_1729,N_29975,N_29324);
or UO_1730 (O_1730,N_29466,N_29577);
and UO_1731 (O_1731,N_29532,N_28842);
and UO_1732 (O_1732,N_28599,N_29712);
nor UO_1733 (O_1733,N_29927,N_28613);
or UO_1734 (O_1734,N_29801,N_29217);
and UO_1735 (O_1735,N_29044,N_29265);
or UO_1736 (O_1736,N_29895,N_29924);
or UO_1737 (O_1737,N_29458,N_29050);
nor UO_1738 (O_1738,N_28741,N_29665);
or UO_1739 (O_1739,N_29983,N_29461);
nor UO_1740 (O_1740,N_29145,N_28950);
nor UO_1741 (O_1741,N_28768,N_28871);
and UO_1742 (O_1742,N_29049,N_29441);
and UO_1743 (O_1743,N_28712,N_28536);
or UO_1744 (O_1744,N_28751,N_28780);
xnor UO_1745 (O_1745,N_28601,N_28802);
xor UO_1746 (O_1746,N_28918,N_29494);
nor UO_1747 (O_1747,N_29588,N_29904);
nor UO_1748 (O_1748,N_29457,N_28563);
nor UO_1749 (O_1749,N_29417,N_29464);
and UO_1750 (O_1750,N_29643,N_28876);
nor UO_1751 (O_1751,N_29150,N_29160);
or UO_1752 (O_1752,N_29660,N_29497);
and UO_1753 (O_1753,N_29165,N_29843);
or UO_1754 (O_1754,N_29266,N_29993);
and UO_1755 (O_1755,N_28732,N_29402);
nand UO_1756 (O_1756,N_29511,N_29680);
nor UO_1757 (O_1757,N_29842,N_29201);
and UO_1758 (O_1758,N_29807,N_28529);
nor UO_1759 (O_1759,N_29695,N_29641);
and UO_1760 (O_1760,N_28596,N_28907);
or UO_1761 (O_1761,N_28570,N_29162);
xor UO_1762 (O_1762,N_29019,N_28627);
nor UO_1763 (O_1763,N_28633,N_29397);
nor UO_1764 (O_1764,N_29277,N_28550);
or UO_1765 (O_1765,N_29570,N_28648);
xor UO_1766 (O_1766,N_29293,N_29754);
xnor UO_1767 (O_1767,N_29078,N_28518);
xor UO_1768 (O_1768,N_29960,N_29713);
nand UO_1769 (O_1769,N_29708,N_29490);
xnor UO_1770 (O_1770,N_28523,N_29964);
and UO_1771 (O_1771,N_29020,N_29583);
nor UO_1772 (O_1772,N_28899,N_29283);
nor UO_1773 (O_1773,N_29548,N_29915);
nor UO_1774 (O_1774,N_29832,N_28547);
or UO_1775 (O_1775,N_28864,N_28849);
nor UO_1776 (O_1776,N_29214,N_28851);
and UO_1777 (O_1777,N_29205,N_28613);
or UO_1778 (O_1778,N_28542,N_28698);
nand UO_1779 (O_1779,N_29128,N_29693);
xnor UO_1780 (O_1780,N_29566,N_28976);
nand UO_1781 (O_1781,N_29476,N_28994);
and UO_1782 (O_1782,N_28700,N_29189);
nand UO_1783 (O_1783,N_28696,N_28899);
or UO_1784 (O_1784,N_28974,N_29597);
or UO_1785 (O_1785,N_29755,N_28768);
and UO_1786 (O_1786,N_29293,N_28547);
xor UO_1787 (O_1787,N_29420,N_29205);
xor UO_1788 (O_1788,N_28625,N_29612);
and UO_1789 (O_1789,N_29078,N_29450);
nand UO_1790 (O_1790,N_29779,N_28513);
and UO_1791 (O_1791,N_29812,N_29545);
nor UO_1792 (O_1792,N_29797,N_29566);
xnor UO_1793 (O_1793,N_28823,N_29510);
or UO_1794 (O_1794,N_29886,N_29928);
nand UO_1795 (O_1795,N_29784,N_29249);
xnor UO_1796 (O_1796,N_29168,N_29990);
xnor UO_1797 (O_1797,N_28719,N_29172);
nand UO_1798 (O_1798,N_29175,N_29091);
nand UO_1799 (O_1799,N_29187,N_29969);
or UO_1800 (O_1800,N_28664,N_29696);
nand UO_1801 (O_1801,N_29250,N_29698);
nor UO_1802 (O_1802,N_28805,N_29077);
xnor UO_1803 (O_1803,N_29445,N_29118);
nand UO_1804 (O_1804,N_28606,N_29682);
nand UO_1805 (O_1805,N_29138,N_29212);
and UO_1806 (O_1806,N_29532,N_28731);
or UO_1807 (O_1807,N_28678,N_29376);
nor UO_1808 (O_1808,N_28785,N_28879);
nand UO_1809 (O_1809,N_28694,N_29995);
nand UO_1810 (O_1810,N_29536,N_29257);
xor UO_1811 (O_1811,N_29419,N_28532);
or UO_1812 (O_1812,N_29194,N_29135);
xnor UO_1813 (O_1813,N_28764,N_29693);
nor UO_1814 (O_1814,N_28706,N_28837);
xor UO_1815 (O_1815,N_29012,N_29274);
and UO_1816 (O_1816,N_29945,N_28878);
nand UO_1817 (O_1817,N_29416,N_28831);
nand UO_1818 (O_1818,N_28670,N_28576);
xnor UO_1819 (O_1819,N_29205,N_29811);
and UO_1820 (O_1820,N_29396,N_29132);
xor UO_1821 (O_1821,N_29063,N_29515);
nor UO_1822 (O_1822,N_29841,N_29074);
nand UO_1823 (O_1823,N_29311,N_29532);
or UO_1824 (O_1824,N_29535,N_29088);
and UO_1825 (O_1825,N_29531,N_29412);
nor UO_1826 (O_1826,N_28552,N_29235);
xnor UO_1827 (O_1827,N_29824,N_29747);
nand UO_1828 (O_1828,N_29854,N_28963);
nor UO_1829 (O_1829,N_29208,N_28980);
and UO_1830 (O_1830,N_29366,N_29872);
nand UO_1831 (O_1831,N_28811,N_29456);
or UO_1832 (O_1832,N_29593,N_29184);
and UO_1833 (O_1833,N_29218,N_28831);
nor UO_1834 (O_1834,N_28750,N_29844);
xnor UO_1835 (O_1835,N_29554,N_29188);
and UO_1836 (O_1836,N_29817,N_29766);
nand UO_1837 (O_1837,N_29036,N_29153);
nor UO_1838 (O_1838,N_28803,N_29333);
nor UO_1839 (O_1839,N_29430,N_28659);
and UO_1840 (O_1840,N_29350,N_29399);
nand UO_1841 (O_1841,N_28621,N_29551);
nand UO_1842 (O_1842,N_29733,N_29113);
nor UO_1843 (O_1843,N_29843,N_29692);
xnor UO_1844 (O_1844,N_29040,N_29966);
nor UO_1845 (O_1845,N_29937,N_29238);
and UO_1846 (O_1846,N_29391,N_29290);
or UO_1847 (O_1847,N_29615,N_29977);
or UO_1848 (O_1848,N_29210,N_29294);
nand UO_1849 (O_1849,N_29757,N_28633);
and UO_1850 (O_1850,N_29344,N_28601);
or UO_1851 (O_1851,N_29123,N_29679);
nor UO_1852 (O_1852,N_29184,N_28630);
and UO_1853 (O_1853,N_29618,N_29281);
and UO_1854 (O_1854,N_29161,N_28943);
xnor UO_1855 (O_1855,N_29678,N_29713);
and UO_1856 (O_1856,N_29281,N_29362);
nor UO_1857 (O_1857,N_29694,N_29030);
and UO_1858 (O_1858,N_28906,N_29983);
nand UO_1859 (O_1859,N_29552,N_29736);
xnor UO_1860 (O_1860,N_28957,N_29829);
nor UO_1861 (O_1861,N_28654,N_28749);
nor UO_1862 (O_1862,N_28835,N_29976);
xor UO_1863 (O_1863,N_29165,N_29529);
or UO_1864 (O_1864,N_29388,N_28988);
or UO_1865 (O_1865,N_29253,N_29725);
nor UO_1866 (O_1866,N_28506,N_28557);
or UO_1867 (O_1867,N_29966,N_29721);
nor UO_1868 (O_1868,N_28737,N_28641);
xor UO_1869 (O_1869,N_29343,N_29764);
xor UO_1870 (O_1870,N_28935,N_29544);
nor UO_1871 (O_1871,N_29960,N_28885);
nand UO_1872 (O_1872,N_29228,N_29514);
nor UO_1873 (O_1873,N_29011,N_28625);
and UO_1874 (O_1874,N_29217,N_29643);
and UO_1875 (O_1875,N_28659,N_29220);
and UO_1876 (O_1876,N_29573,N_28733);
and UO_1877 (O_1877,N_28585,N_29982);
or UO_1878 (O_1878,N_29942,N_28607);
nand UO_1879 (O_1879,N_28638,N_29324);
or UO_1880 (O_1880,N_29466,N_29925);
nor UO_1881 (O_1881,N_28932,N_29778);
nor UO_1882 (O_1882,N_29272,N_28598);
nor UO_1883 (O_1883,N_28701,N_28630);
nor UO_1884 (O_1884,N_28889,N_29962);
or UO_1885 (O_1885,N_28875,N_28623);
or UO_1886 (O_1886,N_29537,N_29611);
or UO_1887 (O_1887,N_29854,N_28560);
nor UO_1888 (O_1888,N_29706,N_28670);
and UO_1889 (O_1889,N_29049,N_28608);
nand UO_1890 (O_1890,N_29825,N_29666);
or UO_1891 (O_1891,N_29174,N_29896);
nor UO_1892 (O_1892,N_29233,N_29307);
xnor UO_1893 (O_1893,N_29083,N_29260);
nor UO_1894 (O_1894,N_29398,N_29161);
or UO_1895 (O_1895,N_29867,N_29111);
or UO_1896 (O_1896,N_29980,N_29101);
nand UO_1897 (O_1897,N_29606,N_29692);
and UO_1898 (O_1898,N_29215,N_28833);
nand UO_1899 (O_1899,N_29968,N_29577);
xor UO_1900 (O_1900,N_29790,N_28960);
nand UO_1901 (O_1901,N_28739,N_29871);
and UO_1902 (O_1902,N_28517,N_29929);
nor UO_1903 (O_1903,N_29770,N_29369);
and UO_1904 (O_1904,N_29779,N_29213);
or UO_1905 (O_1905,N_29551,N_29449);
nor UO_1906 (O_1906,N_29687,N_29583);
and UO_1907 (O_1907,N_29789,N_28874);
nand UO_1908 (O_1908,N_29506,N_29187);
nand UO_1909 (O_1909,N_28642,N_29956);
xor UO_1910 (O_1910,N_29175,N_29697);
nand UO_1911 (O_1911,N_29707,N_29059);
and UO_1912 (O_1912,N_29436,N_29110);
or UO_1913 (O_1913,N_29721,N_29949);
nand UO_1914 (O_1914,N_29871,N_29458);
or UO_1915 (O_1915,N_28600,N_29011);
or UO_1916 (O_1916,N_29121,N_29466);
and UO_1917 (O_1917,N_28881,N_29186);
xnor UO_1918 (O_1918,N_28596,N_28806);
and UO_1919 (O_1919,N_29012,N_28673);
nand UO_1920 (O_1920,N_29843,N_29509);
nor UO_1921 (O_1921,N_29401,N_29048);
or UO_1922 (O_1922,N_29424,N_29514);
nand UO_1923 (O_1923,N_29169,N_29346);
nor UO_1924 (O_1924,N_29896,N_28525);
nor UO_1925 (O_1925,N_29308,N_28691);
nor UO_1926 (O_1926,N_29934,N_29433);
or UO_1927 (O_1927,N_28952,N_28565);
xnor UO_1928 (O_1928,N_29906,N_29656);
or UO_1929 (O_1929,N_29222,N_29414);
xor UO_1930 (O_1930,N_28858,N_28634);
nand UO_1931 (O_1931,N_29311,N_29235);
and UO_1932 (O_1932,N_29887,N_28798);
nor UO_1933 (O_1933,N_28836,N_28604);
nand UO_1934 (O_1934,N_29901,N_29981);
nor UO_1935 (O_1935,N_28910,N_29543);
nand UO_1936 (O_1936,N_28865,N_29060);
and UO_1937 (O_1937,N_29403,N_29529);
or UO_1938 (O_1938,N_29434,N_28555);
or UO_1939 (O_1939,N_28834,N_28763);
xnor UO_1940 (O_1940,N_29562,N_28623);
nand UO_1941 (O_1941,N_29617,N_29460);
xor UO_1942 (O_1942,N_29228,N_28520);
and UO_1943 (O_1943,N_29392,N_28559);
nand UO_1944 (O_1944,N_28562,N_29868);
or UO_1945 (O_1945,N_29398,N_28573);
nor UO_1946 (O_1946,N_29516,N_29265);
xor UO_1947 (O_1947,N_29921,N_28821);
or UO_1948 (O_1948,N_29880,N_29302);
or UO_1949 (O_1949,N_28671,N_29493);
xnor UO_1950 (O_1950,N_29779,N_29791);
nand UO_1951 (O_1951,N_28656,N_28547);
xnor UO_1952 (O_1952,N_29284,N_29222);
xor UO_1953 (O_1953,N_29674,N_29313);
or UO_1954 (O_1954,N_28819,N_29553);
or UO_1955 (O_1955,N_28828,N_28733);
nor UO_1956 (O_1956,N_29699,N_29859);
nor UO_1957 (O_1957,N_29828,N_29841);
nand UO_1958 (O_1958,N_29652,N_29611);
and UO_1959 (O_1959,N_28961,N_28773);
nor UO_1960 (O_1960,N_29870,N_29820);
nor UO_1961 (O_1961,N_28953,N_29099);
nor UO_1962 (O_1962,N_28592,N_29078);
and UO_1963 (O_1963,N_29128,N_28995);
nor UO_1964 (O_1964,N_29291,N_29463);
or UO_1965 (O_1965,N_29943,N_29766);
or UO_1966 (O_1966,N_29602,N_29715);
nand UO_1967 (O_1967,N_28844,N_29066);
nand UO_1968 (O_1968,N_29081,N_29676);
and UO_1969 (O_1969,N_28579,N_29150);
xor UO_1970 (O_1970,N_28565,N_28819);
xor UO_1971 (O_1971,N_29504,N_29645);
or UO_1972 (O_1972,N_29223,N_29634);
or UO_1973 (O_1973,N_28892,N_29625);
nand UO_1974 (O_1974,N_28720,N_28504);
xor UO_1975 (O_1975,N_29226,N_28812);
nand UO_1976 (O_1976,N_28760,N_29916);
and UO_1977 (O_1977,N_29054,N_28816);
xnor UO_1978 (O_1978,N_29623,N_28715);
and UO_1979 (O_1979,N_28777,N_29444);
xnor UO_1980 (O_1980,N_28927,N_28598);
and UO_1981 (O_1981,N_29386,N_29584);
or UO_1982 (O_1982,N_28753,N_29524);
or UO_1983 (O_1983,N_29174,N_28683);
nor UO_1984 (O_1984,N_29361,N_29834);
nand UO_1985 (O_1985,N_29740,N_28506);
nor UO_1986 (O_1986,N_29268,N_29839);
nor UO_1987 (O_1987,N_28869,N_28582);
nand UO_1988 (O_1988,N_29222,N_29608);
or UO_1989 (O_1989,N_29015,N_29115);
nand UO_1990 (O_1990,N_29040,N_28812);
nor UO_1991 (O_1991,N_29009,N_29271);
xnor UO_1992 (O_1992,N_29853,N_29430);
nand UO_1993 (O_1993,N_28620,N_28827);
xnor UO_1994 (O_1994,N_29653,N_29576);
xor UO_1995 (O_1995,N_29155,N_28804);
or UO_1996 (O_1996,N_29987,N_28806);
xnor UO_1997 (O_1997,N_28843,N_29431);
or UO_1998 (O_1998,N_29833,N_29088);
and UO_1999 (O_1999,N_28626,N_29488);
xor UO_2000 (O_2000,N_28939,N_29935);
nand UO_2001 (O_2001,N_28740,N_29272);
nor UO_2002 (O_2002,N_28617,N_28893);
nand UO_2003 (O_2003,N_28978,N_29316);
nor UO_2004 (O_2004,N_29038,N_28704);
xor UO_2005 (O_2005,N_28800,N_28590);
xnor UO_2006 (O_2006,N_29708,N_28943);
or UO_2007 (O_2007,N_28633,N_28525);
nand UO_2008 (O_2008,N_29707,N_29462);
or UO_2009 (O_2009,N_29968,N_29721);
nand UO_2010 (O_2010,N_28557,N_29106);
nand UO_2011 (O_2011,N_29701,N_29196);
nand UO_2012 (O_2012,N_29354,N_29412);
nand UO_2013 (O_2013,N_28713,N_29955);
nand UO_2014 (O_2014,N_28813,N_29665);
nand UO_2015 (O_2015,N_29044,N_28845);
or UO_2016 (O_2016,N_29756,N_29594);
or UO_2017 (O_2017,N_29194,N_28854);
xor UO_2018 (O_2018,N_29096,N_28584);
or UO_2019 (O_2019,N_28623,N_29182);
and UO_2020 (O_2020,N_29448,N_29438);
nand UO_2021 (O_2021,N_29801,N_29694);
and UO_2022 (O_2022,N_28536,N_28754);
and UO_2023 (O_2023,N_28766,N_29625);
nand UO_2024 (O_2024,N_29378,N_29587);
or UO_2025 (O_2025,N_29626,N_29190);
xor UO_2026 (O_2026,N_29572,N_29966);
nand UO_2027 (O_2027,N_28960,N_28988);
nand UO_2028 (O_2028,N_28539,N_29153);
and UO_2029 (O_2029,N_29024,N_29975);
or UO_2030 (O_2030,N_28619,N_29320);
xnor UO_2031 (O_2031,N_28851,N_29860);
nor UO_2032 (O_2032,N_29695,N_29211);
or UO_2033 (O_2033,N_29594,N_29860);
nand UO_2034 (O_2034,N_29351,N_29518);
nand UO_2035 (O_2035,N_28831,N_28649);
and UO_2036 (O_2036,N_29562,N_29753);
nor UO_2037 (O_2037,N_29373,N_29542);
and UO_2038 (O_2038,N_29123,N_28588);
nand UO_2039 (O_2039,N_29074,N_29405);
nand UO_2040 (O_2040,N_29844,N_29249);
xnor UO_2041 (O_2041,N_29660,N_28761);
and UO_2042 (O_2042,N_29082,N_28860);
and UO_2043 (O_2043,N_29268,N_29485);
or UO_2044 (O_2044,N_29407,N_29296);
nor UO_2045 (O_2045,N_29320,N_29166);
nor UO_2046 (O_2046,N_28746,N_29245);
xnor UO_2047 (O_2047,N_28505,N_28857);
nand UO_2048 (O_2048,N_28673,N_29080);
and UO_2049 (O_2049,N_29587,N_28736);
nor UO_2050 (O_2050,N_28930,N_29497);
and UO_2051 (O_2051,N_29482,N_29799);
nand UO_2052 (O_2052,N_29862,N_29408);
xor UO_2053 (O_2053,N_29794,N_29823);
nor UO_2054 (O_2054,N_28611,N_28722);
nand UO_2055 (O_2055,N_28665,N_28544);
nor UO_2056 (O_2056,N_29422,N_28536);
xor UO_2057 (O_2057,N_28795,N_28698);
or UO_2058 (O_2058,N_29963,N_29343);
xnor UO_2059 (O_2059,N_29146,N_28853);
nand UO_2060 (O_2060,N_29370,N_29944);
and UO_2061 (O_2061,N_28812,N_29760);
and UO_2062 (O_2062,N_28880,N_28502);
or UO_2063 (O_2063,N_29036,N_29489);
or UO_2064 (O_2064,N_29941,N_29773);
nor UO_2065 (O_2065,N_29822,N_29545);
or UO_2066 (O_2066,N_29133,N_29738);
nor UO_2067 (O_2067,N_29262,N_29822);
xor UO_2068 (O_2068,N_29890,N_29340);
or UO_2069 (O_2069,N_28727,N_28946);
nor UO_2070 (O_2070,N_28728,N_29719);
xnor UO_2071 (O_2071,N_29769,N_28554);
and UO_2072 (O_2072,N_28526,N_29492);
nor UO_2073 (O_2073,N_29224,N_28796);
and UO_2074 (O_2074,N_29282,N_28829);
xor UO_2075 (O_2075,N_29332,N_29393);
nand UO_2076 (O_2076,N_29631,N_29670);
nor UO_2077 (O_2077,N_29909,N_29260);
nor UO_2078 (O_2078,N_28845,N_28788);
xor UO_2079 (O_2079,N_28528,N_28522);
or UO_2080 (O_2080,N_29299,N_28653);
nor UO_2081 (O_2081,N_29075,N_28746);
xor UO_2082 (O_2082,N_29973,N_28983);
xor UO_2083 (O_2083,N_29914,N_29161);
or UO_2084 (O_2084,N_29487,N_28883);
or UO_2085 (O_2085,N_29517,N_29448);
or UO_2086 (O_2086,N_28632,N_29915);
nand UO_2087 (O_2087,N_28832,N_29499);
or UO_2088 (O_2088,N_29715,N_28519);
and UO_2089 (O_2089,N_29973,N_28574);
or UO_2090 (O_2090,N_29738,N_29992);
xor UO_2091 (O_2091,N_29193,N_29461);
xor UO_2092 (O_2092,N_29651,N_29120);
nor UO_2093 (O_2093,N_29193,N_29047);
nand UO_2094 (O_2094,N_28720,N_28936);
and UO_2095 (O_2095,N_28528,N_28960);
xor UO_2096 (O_2096,N_29223,N_29101);
nor UO_2097 (O_2097,N_29485,N_29126);
or UO_2098 (O_2098,N_29619,N_29340);
nand UO_2099 (O_2099,N_29842,N_29506);
nor UO_2100 (O_2100,N_28882,N_28685);
xnor UO_2101 (O_2101,N_29498,N_29342);
nor UO_2102 (O_2102,N_29314,N_29776);
nand UO_2103 (O_2103,N_29664,N_29352);
nor UO_2104 (O_2104,N_28981,N_29682);
or UO_2105 (O_2105,N_28537,N_29527);
nand UO_2106 (O_2106,N_28718,N_29467);
and UO_2107 (O_2107,N_28684,N_29127);
nor UO_2108 (O_2108,N_29054,N_29055);
nand UO_2109 (O_2109,N_28856,N_29822);
or UO_2110 (O_2110,N_29798,N_29049);
nand UO_2111 (O_2111,N_28900,N_29809);
nor UO_2112 (O_2112,N_29162,N_29383);
nand UO_2113 (O_2113,N_29476,N_29416);
and UO_2114 (O_2114,N_28504,N_29814);
nor UO_2115 (O_2115,N_29124,N_29006);
nand UO_2116 (O_2116,N_29463,N_28649);
xor UO_2117 (O_2117,N_29794,N_29610);
or UO_2118 (O_2118,N_28546,N_28977);
and UO_2119 (O_2119,N_29269,N_29888);
and UO_2120 (O_2120,N_29798,N_28714);
nor UO_2121 (O_2121,N_29737,N_29336);
or UO_2122 (O_2122,N_28983,N_29684);
nor UO_2123 (O_2123,N_29445,N_28725);
or UO_2124 (O_2124,N_28982,N_29557);
nor UO_2125 (O_2125,N_28740,N_29836);
nand UO_2126 (O_2126,N_29418,N_28613);
or UO_2127 (O_2127,N_28647,N_29874);
nor UO_2128 (O_2128,N_29789,N_29449);
nor UO_2129 (O_2129,N_28565,N_29573);
xor UO_2130 (O_2130,N_29663,N_29958);
and UO_2131 (O_2131,N_29744,N_29511);
nand UO_2132 (O_2132,N_28989,N_29576);
nor UO_2133 (O_2133,N_29773,N_29609);
nand UO_2134 (O_2134,N_29364,N_29287);
nor UO_2135 (O_2135,N_29694,N_28749);
nand UO_2136 (O_2136,N_29057,N_28578);
or UO_2137 (O_2137,N_28996,N_29984);
and UO_2138 (O_2138,N_29761,N_29052);
nand UO_2139 (O_2139,N_28838,N_29273);
and UO_2140 (O_2140,N_29906,N_28903);
nor UO_2141 (O_2141,N_28849,N_29856);
or UO_2142 (O_2142,N_29041,N_29667);
or UO_2143 (O_2143,N_29789,N_29608);
and UO_2144 (O_2144,N_29699,N_29778);
and UO_2145 (O_2145,N_29878,N_29666);
xor UO_2146 (O_2146,N_29817,N_29574);
or UO_2147 (O_2147,N_28935,N_29921);
xor UO_2148 (O_2148,N_29176,N_28750);
nand UO_2149 (O_2149,N_29745,N_28864);
xor UO_2150 (O_2150,N_29752,N_29113);
xnor UO_2151 (O_2151,N_29661,N_29281);
nand UO_2152 (O_2152,N_29386,N_28701);
and UO_2153 (O_2153,N_29504,N_29616);
or UO_2154 (O_2154,N_29567,N_28893);
nand UO_2155 (O_2155,N_29459,N_29073);
nand UO_2156 (O_2156,N_29498,N_28817);
nor UO_2157 (O_2157,N_28589,N_29226);
nor UO_2158 (O_2158,N_28989,N_29408);
or UO_2159 (O_2159,N_28850,N_29393);
nand UO_2160 (O_2160,N_29943,N_29250);
xnor UO_2161 (O_2161,N_29156,N_29277);
nor UO_2162 (O_2162,N_29847,N_29855);
nor UO_2163 (O_2163,N_28759,N_29563);
xor UO_2164 (O_2164,N_29588,N_28630);
nand UO_2165 (O_2165,N_29037,N_29439);
xor UO_2166 (O_2166,N_29234,N_29352);
nor UO_2167 (O_2167,N_29890,N_28953);
and UO_2168 (O_2168,N_29023,N_29520);
xnor UO_2169 (O_2169,N_29891,N_29873);
xor UO_2170 (O_2170,N_28727,N_29117);
or UO_2171 (O_2171,N_29509,N_29335);
nand UO_2172 (O_2172,N_29098,N_28714);
nor UO_2173 (O_2173,N_28931,N_29139);
xnor UO_2174 (O_2174,N_28570,N_29373);
and UO_2175 (O_2175,N_29382,N_28632);
nand UO_2176 (O_2176,N_28798,N_28958);
and UO_2177 (O_2177,N_29159,N_29728);
nor UO_2178 (O_2178,N_28919,N_28952);
xnor UO_2179 (O_2179,N_29826,N_28899);
nand UO_2180 (O_2180,N_29499,N_29263);
or UO_2181 (O_2181,N_28561,N_29989);
or UO_2182 (O_2182,N_29068,N_28588);
nor UO_2183 (O_2183,N_29896,N_28960);
nor UO_2184 (O_2184,N_29996,N_29434);
nand UO_2185 (O_2185,N_28752,N_29611);
or UO_2186 (O_2186,N_29353,N_28540);
or UO_2187 (O_2187,N_29622,N_29282);
xor UO_2188 (O_2188,N_28943,N_29812);
nand UO_2189 (O_2189,N_28782,N_29093);
and UO_2190 (O_2190,N_29043,N_29834);
and UO_2191 (O_2191,N_29695,N_28547);
xor UO_2192 (O_2192,N_28807,N_28569);
and UO_2193 (O_2193,N_29926,N_29288);
nor UO_2194 (O_2194,N_29121,N_29135);
nand UO_2195 (O_2195,N_28981,N_29768);
nor UO_2196 (O_2196,N_29731,N_29209);
or UO_2197 (O_2197,N_28836,N_29114);
xor UO_2198 (O_2198,N_29548,N_29742);
or UO_2199 (O_2199,N_29315,N_29663);
xor UO_2200 (O_2200,N_28505,N_28915);
and UO_2201 (O_2201,N_29668,N_28713);
nand UO_2202 (O_2202,N_29468,N_28978);
and UO_2203 (O_2203,N_29918,N_28998);
xnor UO_2204 (O_2204,N_29264,N_29740);
or UO_2205 (O_2205,N_29738,N_29152);
or UO_2206 (O_2206,N_29729,N_29505);
nand UO_2207 (O_2207,N_29439,N_29635);
xnor UO_2208 (O_2208,N_29414,N_29112);
and UO_2209 (O_2209,N_28801,N_29875);
and UO_2210 (O_2210,N_29670,N_29200);
or UO_2211 (O_2211,N_28660,N_29977);
nand UO_2212 (O_2212,N_29726,N_29038);
and UO_2213 (O_2213,N_29428,N_29586);
xor UO_2214 (O_2214,N_29194,N_29971);
nor UO_2215 (O_2215,N_29172,N_29867);
nand UO_2216 (O_2216,N_29890,N_29572);
and UO_2217 (O_2217,N_28773,N_29439);
nor UO_2218 (O_2218,N_29987,N_29148);
xnor UO_2219 (O_2219,N_29058,N_29415);
nand UO_2220 (O_2220,N_29556,N_29580);
xnor UO_2221 (O_2221,N_28948,N_29838);
nand UO_2222 (O_2222,N_28684,N_29080);
or UO_2223 (O_2223,N_29278,N_29609);
nor UO_2224 (O_2224,N_29028,N_28965);
xor UO_2225 (O_2225,N_29153,N_29166);
xnor UO_2226 (O_2226,N_29391,N_29648);
and UO_2227 (O_2227,N_28883,N_29402);
nor UO_2228 (O_2228,N_28723,N_29716);
nand UO_2229 (O_2229,N_28994,N_29252);
nor UO_2230 (O_2230,N_28943,N_29746);
xor UO_2231 (O_2231,N_28971,N_28815);
nand UO_2232 (O_2232,N_29134,N_28829);
nand UO_2233 (O_2233,N_29009,N_29918);
and UO_2234 (O_2234,N_29607,N_29198);
or UO_2235 (O_2235,N_28762,N_28966);
nand UO_2236 (O_2236,N_29390,N_29344);
nand UO_2237 (O_2237,N_29274,N_28661);
nor UO_2238 (O_2238,N_28598,N_29245);
and UO_2239 (O_2239,N_29738,N_29434);
nand UO_2240 (O_2240,N_28944,N_29804);
nor UO_2241 (O_2241,N_28552,N_28560);
nor UO_2242 (O_2242,N_29492,N_29105);
xor UO_2243 (O_2243,N_29878,N_29110);
nor UO_2244 (O_2244,N_28929,N_29718);
xor UO_2245 (O_2245,N_29432,N_28618);
nor UO_2246 (O_2246,N_29628,N_29516);
nand UO_2247 (O_2247,N_28663,N_28799);
and UO_2248 (O_2248,N_29615,N_29784);
or UO_2249 (O_2249,N_28747,N_29786);
or UO_2250 (O_2250,N_29772,N_29321);
and UO_2251 (O_2251,N_29243,N_29984);
or UO_2252 (O_2252,N_29553,N_29693);
nor UO_2253 (O_2253,N_28905,N_28771);
and UO_2254 (O_2254,N_29402,N_28657);
nor UO_2255 (O_2255,N_28585,N_28667);
xnor UO_2256 (O_2256,N_29338,N_28795);
and UO_2257 (O_2257,N_29474,N_28516);
or UO_2258 (O_2258,N_28826,N_29845);
and UO_2259 (O_2259,N_28904,N_28582);
xnor UO_2260 (O_2260,N_29539,N_28752);
nor UO_2261 (O_2261,N_28728,N_29212);
nand UO_2262 (O_2262,N_28921,N_29781);
xor UO_2263 (O_2263,N_28954,N_28975);
nor UO_2264 (O_2264,N_28634,N_29483);
and UO_2265 (O_2265,N_29369,N_28861);
nand UO_2266 (O_2266,N_29717,N_28962);
or UO_2267 (O_2267,N_28697,N_29025);
nand UO_2268 (O_2268,N_29951,N_29550);
xor UO_2269 (O_2269,N_29018,N_29227);
xor UO_2270 (O_2270,N_28891,N_29583);
xor UO_2271 (O_2271,N_29531,N_29882);
nand UO_2272 (O_2272,N_29543,N_29255);
nor UO_2273 (O_2273,N_29992,N_29384);
xor UO_2274 (O_2274,N_29283,N_29336);
xor UO_2275 (O_2275,N_29675,N_29378);
nand UO_2276 (O_2276,N_28868,N_29199);
nor UO_2277 (O_2277,N_29459,N_29937);
and UO_2278 (O_2278,N_28918,N_29336);
nor UO_2279 (O_2279,N_28738,N_29896);
nand UO_2280 (O_2280,N_29646,N_28770);
and UO_2281 (O_2281,N_29854,N_29463);
xor UO_2282 (O_2282,N_28837,N_28534);
xor UO_2283 (O_2283,N_29191,N_28725);
or UO_2284 (O_2284,N_29349,N_28969);
nand UO_2285 (O_2285,N_28675,N_29319);
and UO_2286 (O_2286,N_28715,N_29603);
or UO_2287 (O_2287,N_29943,N_29503);
nor UO_2288 (O_2288,N_28689,N_29014);
nor UO_2289 (O_2289,N_28688,N_29597);
nor UO_2290 (O_2290,N_29909,N_29065);
and UO_2291 (O_2291,N_28714,N_29573);
and UO_2292 (O_2292,N_29206,N_28971);
xnor UO_2293 (O_2293,N_29298,N_29423);
or UO_2294 (O_2294,N_28768,N_29191);
nand UO_2295 (O_2295,N_28620,N_29850);
xnor UO_2296 (O_2296,N_29355,N_29699);
and UO_2297 (O_2297,N_28760,N_29268);
nor UO_2298 (O_2298,N_29546,N_28824);
nor UO_2299 (O_2299,N_29626,N_28913);
or UO_2300 (O_2300,N_29882,N_28941);
xor UO_2301 (O_2301,N_29685,N_29687);
or UO_2302 (O_2302,N_28577,N_29639);
xnor UO_2303 (O_2303,N_29281,N_29946);
and UO_2304 (O_2304,N_29844,N_29717);
nand UO_2305 (O_2305,N_28894,N_29188);
xor UO_2306 (O_2306,N_29024,N_29514);
xnor UO_2307 (O_2307,N_28530,N_29486);
nand UO_2308 (O_2308,N_29751,N_29132);
nand UO_2309 (O_2309,N_28712,N_28891);
or UO_2310 (O_2310,N_29495,N_29936);
and UO_2311 (O_2311,N_28747,N_29605);
or UO_2312 (O_2312,N_29027,N_28750);
or UO_2313 (O_2313,N_28983,N_28507);
nand UO_2314 (O_2314,N_29789,N_29711);
nand UO_2315 (O_2315,N_29353,N_29316);
nor UO_2316 (O_2316,N_28800,N_28820);
nand UO_2317 (O_2317,N_29649,N_28684);
nor UO_2318 (O_2318,N_29624,N_28764);
xor UO_2319 (O_2319,N_28783,N_28624);
and UO_2320 (O_2320,N_29616,N_28816);
nand UO_2321 (O_2321,N_29624,N_28614);
xor UO_2322 (O_2322,N_29365,N_28903);
or UO_2323 (O_2323,N_29557,N_28946);
nor UO_2324 (O_2324,N_28756,N_29210);
nor UO_2325 (O_2325,N_29810,N_29375);
and UO_2326 (O_2326,N_29203,N_29880);
nand UO_2327 (O_2327,N_29385,N_29829);
or UO_2328 (O_2328,N_29875,N_29448);
and UO_2329 (O_2329,N_29722,N_29050);
nor UO_2330 (O_2330,N_29072,N_28606);
or UO_2331 (O_2331,N_29783,N_28904);
nand UO_2332 (O_2332,N_29755,N_29222);
nand UO_2333 (O_2333,N_29979,N_28747);
xor UO_2334 (O_2334,N_29222,N_28732);
nor UO_2335 (O_2335,N_28517,N_29345);
or UO_2336 (O_2336,N_29563,N_29230);
nor UO_2337 (O_2337,N_29538,N_29603);
or UO_2338 (O_2338,N_29662,N_28922);
and UO_2339 (O_2339,N_28803,N_29202);
and UO_2340 (O_2340,N_28619,N_29750);
nand UO_2341 (O_2341,N_29966,N_29918);
nor UO_2342 (O_2342,N_28991,N_28724);
or UO_2343 (O_2343,N_29267,N_29533);
nand UO_2344 (O_2344,N_28699,N_29360);
and UO_2345 (O_2345,N_29050,N_28927);
nor UO_2346 (O_2346,N_29870,N_29351);
and UO_2347 (O_2347,N_29969,N_28818);
xnor UO_2348 (O_2348,N_28580,N_29411);
xnor UO_2349 (O_2349,N_29963,N_29091);
or UO_2350 (O_2350,N_28941,N_29937);
and UO_2351 (O_2351,N_29997,N_29330);
xnor UO_2352 (O_2352,N_29235,N_29784);
nor UO_2353 (O_2353,N_29006,N_29547);
or UO_2354 (O_2354,N_29075,N_28813);
and UO_2355 (O_2355,N_29491,N_29298);
nor UO_2356 (O_2356,N_28937,N_28990);
and UO_2357 (O_2357,N_29532,N_28883);
nor UO_2358 (O_2358,N_28738,N_29709);
xor UO_2359 (O_2359,N_29445,N_29392);
xor UO_2360 (O_2360,N_29769,N_29514);
nand UO_2361 (O_2361,N_29769,N_29935);
or UO_2362 (O_2362,N_29382,N_29620);
nor UO_2363 (O_2363,N_29790,N_29941);
nand UO_2364 (O_2364,N_28967,N_29724);
nor UO_2365 (O_2365,N_29318,N_29873);
and UO_2366 (O_2366,N_29225,N_28652);
nor UO_2367 (O_2367,N_29190,N_28517);
nand UO_2368 (O_2368,N_29549,N_29094);
nand UO_2369 (O_2369,N_29738,N_28590);
nor UO_2370 (O_2370,N_29125,N_29974);
nor UO_2371 (O_2371,N_28948,N_28997);
nor UO_2372 (O_2372,N_29667,N_29228);
and UO_2373 (O_2373,N_28570,N_29883);
nand UO_2374 (O_2374,N_29082,N_29116);
and UO_2375 (O_2375,N_28617,N_29972);
nor UO_2376 (O_2376,N_28995,N_29994);
and UO_2377 (O_2377,N_29999,N_28999);
nor UO_2378 (O_2378,N_29134,N_28552);
nand UO_2379 (O_2379,N_29576,N_28805);
nor UO_2380 (O_2380,N_29858,N_29809);
xnor UO_2381 (O_2381,N_28756,N_28609);
nand UO_2382 (O_2382,N_29870,N_28557);
nor UO_2383 (O_2383,N_29894,N_29498);
xnor UO_2384 (O_2384,N_28923,N_28736);
and UO_2385 (O_2385,N_29719,N_29749);
nand UO_2386 (O_2386,N_28609,N_29894);
and UO_2387 (O_2387,N_29991,N_28889);
nand UO_2388 (O_2388,N_28589,N_28840);
nand UO_2389 (O_2389,N_29850,N_28564);
nor UO_2390 (O_2390,N_29616,N_29212);
and UO_2391 (O_2391,N_28747,N_28994);
and UO_2392 (O_2392,N_29339,N_28681);
and UO_2393 (O_2393,N_29330,N_29088);
xor UO_2394 (O_2394,N_28814,N_29256);
and UO_2395 (O_2395,N_29873,N_29243);
nor UO_2396 (O_2396,N_28791,N_29066);
or UO_2397 (O_2397,N_29946,N_29576);
nand UO_2398 (O_2398,N_29266,N_29279);
or UO_2399 (O_2399,N_28745,N_29438);
xnor UO_2400 (O_2400,N_28641,N_29354);
or UO_2401 (O_2401,N_29518,N_29583);
nor UO_2402 (O_2402,N_28971,N_29554);
xor UO_2403 (O_2403,N_28509,N_28607);
xor UO_2404 (O_2404,N_28517,N_29404);
or UO_2405 (O_2405,N_29022,N_29989);
nor UO_2406 (O_2406,N_29770,N_29651);
xor UO_2407 (O_2407,N_29358,N_28617);
and UO_2408 (O_2408,N_28943,N_29416);
xnor UO_2409 (O_2409,N_28884,N_29217);
xnor UO_2410 (O_2410,N_29886,N_29387);
nor UO_2411 (O_2411,N_29085,N_29461);
or UO_2412 (O_2412,N_28826,N_29874);
xor UO_2413 (O_2413,N_28516,N_29118);
nand UO_2414 (O_2414,N_29403,N_29839);
nand UO_2415 (O_2415,N_29918,N_28803);
xnor UO_2416 (O_2416,N_29906,N_28515);
xnor UO_2417 (O_2417,N_29685,N_29944);
nand UO_2418 (O_2418,N_28561,N_29654);
xnor UO_2419 (O_2419,N_29648,N_29999);
or UO_2420 (O_2420,N_29989,N_29042);
nor UO_2421 (O_2421,N_29348,N_29891);
nor UO_2422 (O_2422,N_28689,N_29704);
xnor UO_2423 (O_2423,N_29237,N_28700);
and UO_2424 (O_2424,N_29571,N_28760);
and UO_2425 (O_2425,N_29260,N_28592);
nand UO_2426 (O_2426,N_29672,N_28557);
nor UO_2427 (O_2427,N_28887,N_29675);
or UO_2428 (O_2428,N_29094,N_29099);
nand UO_2429 (O_2429,N_29473,N_29514);
nor UO_2430 (O_2430,N_29545,N_28900);
xnor UO_2431 (O_2431,N_29423,N_28585);
or UO_2432 (O_2432,N_29202,N_29319);
and UO_2433 (O_2433,N_29880,N_29689);
or UO_2434 (O_2434,N_29522,N_28604);
nand UO_2435 (O_2435,N_29429,N_29033);
nor UO_2436 (O_2436,N_29381,N_28713);
nand UO_2437 (O_2437,N_29552,N_29963);
xnor UO_2438 (O_2438,N_29114,N_28926);
xor UO_2439 (O_2439,N_29293,N_29187);
xor UO_2440 (O_2440,N_29085,N_29067);
and UO_2441 (O_2441,N_28637,N_29612);
or UO_2442 (O_2442,N_28897,N_29095);
or UO_2443 (O_2443,N_28565,N_28540);
and UO_2444 (O_2444,N_29140,N_28696);
and UO_2445 (O_2445,N_28551,N_29860);
xor UO_2446 (O_2446,N_29785,N_29809);
xor UO_2447 (O_2447,N_28816,N_29180);
or UO_2448 (O_2448,N_28827,N_29160);
nor UO_2449 (O_2449,N_29429,N_28618);
and UO_2450 (O_2450,N_29653,N_28803);
nand UO_2451 (O_2451,N_29552,N_29869);
nand UO_2452 (O_2452,N_28690,N_29460);
nor UO_2453 (O_2453,N_29472,N_29064);
and UO_2454 (O_2454,N_29359,N_29351);
and UO_2455 (O_2455,N_29760,N_29474);
nand UO_2456 (O_2456,N_29305,N_29709);
or UO_2457 (O_2457,N_29017,N_28578);
and UO_2458 (O_2458,N_28840,N_28547);
or UO_2459 (O_2459,N_28769,N_29132);
xnor UO_2460 (O_2460,N_29410,N_28642);
nor UO_2461 (O_2461,N_29076,N_28513);
nor UO_2462 (O_2462,N_29707,N_29257);
and UO_2463 (O_2463,N_28741,N_28653);
nor UO_2464 (O_2464,N_29918,N_29435);
nor UO_2465 (O_2465,N_28688,N_28681);
nand UO_2466 (O_2466,N_28572,N_29159);
xor UO_2467 (O_2467,N_28957,N_29034);
nand UO_2468 (O_2468,N_29039,N_28537);
and UO_2469 (O_2469,N_29004,N_28808);
xnor UO_2470 (O_2470,N_29695,N_29880);
and UO_2471 (O_2471,N_28692,N_28537);
and UO_2472 (O_2472,N_29231,N_28882);
nand UO_2473 (O_2473,N_29324,N_28942);
or UO_2474 (O_2474,N_29662,N_29890);
nor UO_2475 (O_2475,N_29249,N_29361);
xnor UO_2476 (O_2476,N_29698,N_29898);
nand UO_2477 (O_2477,N_28711,N_29450);
or UO_2478 (O_2478,N_28717,N_29193);
nor UO_2479 (O_2479,N_29881,N_28631);
nand UO_2480 (O_2480,N_28932,N_28807);
nand UO_2481 (O_2481,N_29239,N_28625);
xnor UO_2482 (O_2482,N_29623,N_29267);
nand UO_2483 (O_2483,N_29345,N_29669);
nand UO_2484 (O_2484,N_29119,N_29650);
and UO_2485 (O_2485,N_29041,N_29337);
xor UO_2486 (O_2486,N_29876,N_28849);
and UO_2487 (O_2487,N_29669,N_29325);
nand UO_2488 (O_2488,N_29470,N_28872);
and UO_2489 (O_2489,N_29765,N_29162);
or UO_2490 (O_2490,N_29900,N_29282);
nor UO_2491 (O_2491,N_28555,N_28915);
or UO_2492 (O_2492,N_29886,N_29221);
nand UO_2493 (O_2493,N_29672,N_28731);
or UO_2494 (O_2494,N_28927,N_29917);
and UO_2495 (O_2495,N_28854,N_29363);
xnor UO_2496 (O_2496,N_29868,N_29957);
nor UO_2497 (O_2497,N_29922,N_29843);
nor UO_2498 (O_2498,N_29502,N_28605);
nor UO_2499 (O_2499,N_28502,N_29973);
and UO_2500 (O_2500,N_29024,N_29799);
and UO_2501 (O_2501,N_28629,N_29995);
xor UO_2502 (O_2502,N_28784,N_29657);
nand UO_2503 (O_2503,N_28865,N_29877);
nor UO_2504 (O_2504,N_28711,N_29520);
and UO_2505 (O_2505,N_29829,N_29803);
and UO_2506 (O_2506,N_29947,N_28944);
and UO_2507 (O_2507,N_29079,N_29684);
or UO_2508 (O_2508,N_29497,N_29556);
or UO_2509 (O_2509,N_28746,N_28908);
and UO_2510 (O_2510,N_29945,N_29222);
xnor UO_2511 (O_2511,N_29558,N_29795);
xnor UO_2512 (O_2512,N_29803,N_29602);
and UO_2513 (O_2513,N_28718,N_29490);
or UO_2514 (O_2514,N_28790,N_29334);
and UO_2515 (O_2515,N_29598,N_28834);
or UO_2516 (O_2516,N_29246,N_29181);
or UO_2517 (O_2517,N_29670,N_29974);
xnor UO_2518 (O_2518,N_29866,N_28908);
nand UO_2519 (O_2519,N_29556,N_29777);
nor UO_2520 (O_2520,N_29518,N_29229);
xor UO_2521 (O_2521,N_29395,N_29016);
xnor UO_2522 (O_2522,N_29539,N_29150);
nor UO_2523 (O_2523,N_29010,N_29748);
xnor UO_2524 (O_2524,N_29607,N_29766);
xnor UO_2525 (O_2525,N_29267,N_29559);
and UO_2526 (O_2526,N_29111,N_29235);
and UO_2527 (O_2527,N_28714,N_29150);
xor UO_2528 (O_2528,N_29833,N_29645);
xor UO_2529 (O_2529,N_29064,N_29518);
and UO_2530 (O_2530,N_29944,N_28681);
and UO_2531 (O_2531,N_29574,N_29157);
nand UO_2532 (O_2532,N_29833,N_29433);
and UO_2533 (O_2533,N_29266,N_28929);
xnor UO_2534 (O_2534,N_29569,N_29929);
and UO_2535 (O_2535,N_28614,N_29408);
nand UO_2536 (O_2536,N_29104,N_28845);
and UO_2537 (O_2537,N_28506,N_29558);
nor UO_2538 (O_2538,N_29187,N_28512);
nor UO_2539 (O_2539,N_29826,N_29266);
nor UO_2540 (O_2540,N_29821,N_29135);
nand UO_2541 (O_2541,N_29495,N_29379);
nor UO_2542 (O_2542,N_28972,N_28919);
nor UO_2543 (O_2543,N_29111,N_29020);
and UO_2544 (O_2544,N_28948,N_29539);
and UO_2545 (O_2545,N_28785,N_28601);
and UO_2546 (O_2546,N_29020,N_28655);
or UO_2547 (O_2547,N_29968,N_29829);
or UO_2548 (O_2548,N_28563,N_29255);
and UO_2549 (O_2549,N_29283,N_28602);
and UO_2550 (O_2550,N_29561,N_28625);
nor UO_2551 (O_2551,N_29225,N_28752);
nor UO_2552 (O_2552,N_28697,N_29083);
xor UO_2553 (O_2553,N_29537,N_29595);
xnor UO_2554 (O_2554,N_29416,N_28880);
or UO_2555 (O_2555,N_29480,N_28947);
xnor UO_2556 (O_2556,N_29412,N_29001);
nor UO_2557 (O_2557,N_29912,N_29336);
nor UO_2558 (O_2558,N_28925,N_28666);
and UO_2559 (O_2559,N_29958,N_29186);
nand UO_2560 (O_2560,N_29119,N_28700);
or UO_2561 (O_2561,N_29125,N_28809);
or UO_2562 (O_2562,N_29940,N_28977);
nand UO_2563 (O_2563,N_29134,N_29336);
nor UO_2564 (O_2564,N_28542,N_29565);
and UO_2565 (O_2565,N_28765,N_28694);
nor UO_2566 (O_2566,N_29437,N_29610);
nor UO_2567 (O_2567,N_29198,N_28771);
nand UO_2568 (O_2568,N_29828,N_28621);
nor UO_2569 (O_2569,N_29424,N_29622);
xor UO_2570 (O_2570,N_29047,N_28780);
and UO_2571 (O_2571,N_28735,N_29821);
and UO_2572 (O_2572,N_29936,N_28722);
xnor UO_2573 (O_2573,N_28789,N_29084);
nand UO_2574 (O_2574,N_29249,N_29913);
nor UO_2575 (O_2575,N_28577,N_29006);
or UO_2576 (O_2576,N_28920,N_29283);
nand UO_2577 (O_2577,N_29240,N_28778);
nand UO_2578 (O_2578,N_29555,N_29258);
or UO_2579 (O_2579,N_29874,N_28862);
nor UO_2580 (O_2580,N_29588,N_28804);
xor UO_2581 (O_2581,N_29652,N_29564);
or UO_2582 (O_2582,N_28593,N_29928);
xnor UO_2583 (O_2583,N_29529,N_28625);
nor UO_2584 (O_2584,N_29825,N_28795);
nand UO_2585 (O_2585,N_29953,N_29078);
or UO_2586 (O_2586,N_28727,N_29594);
xor UO_2587 (O_2587,N_28778,N_28519);
nand UO_2588 (O_2588,N_28711,N_29643);
and UO_2589 (O_2589,N_29882,N_29588);
xnor UO_2590 (O_2590,N_29960,N_29865);
and UO_2591 (O_2591,N_29579,N_28889);
or UO_2592 (O_2592,N_29469,N_28982);
and UO_2593 (O_2593,N_28854,N_28752);
and UO_2594 (O_2594,N_28524,N_29481);
or UO_2595 (O_2595,N_28614,N_28806);
or UO_2596 (O_2596,N_29945,N_29173);
or UO_2597 (O_2597,N_29181,N_28850);
xnor UO_2598 (O_2598,N_28584,N_28587);
xor UO_2599 (O_2599,N_29887,N_28526);
xor UO_2600 (O_2600,N_29064,N_28629);
nand UO_2601 (O_2601,N_29178,N_29221);
nand UO_2602 (O_2602,N_28970,N_29666);
and UO_2603 (O_2603,N_29847,N_29391);
nor UO_2604 (O_2604,N_29585,N_29242);
or UO_2605 (O_2605,N_28965,N_29471);
and UO_2606 (O_2606,N_28888,N_29197);
nor UO_2607 (O_2607,N_29501,N_28875);
or UO_2608 (O_2608,N_29349,N_29852);
or UO_2609 (O_2609,N_29589,N_29867);
or UO_2610 (O_2610,N_29071,N_29290);
nor UO_2611 (O_2611,N_28585,N_28969);
nand UO_2612 (O_2612,N_28511,N_29812);
xor UO_2613 (O_2613,N_29037,N_28808);
and UO_2614 (O_2614,N_29801,N_29233);
xor UO_2615 (O_2615,N_29772,N_29265);
nand UO_2616 (O_2616,N_29120,N_29452);
xnor UO_2617 (O_2617,N_29396,N_29368);
xor UO_2618 (O_2618,N_29610,N_29040);
or UO_2619 (O_2619,N_29970,N_29946);
or UO_2620 (O_2620,N_29937,N_28968);
xnor UO_2621 (O_2621,N_29526,N_29258);
nand UO_2622 (O_2622,N_29996,N_29418);
or UO_2623 (O_2623,N_29308,N_29773);
or UO_2624 (O_2624,N_28842,N_29656);
nand UO_2625 (O_2625,N_29442,N_29363);
and UO_2626 (O_2626,N_29938,N_28697);
xnor UO_2627 (O_2627,N_29117,N_29181);
nor UO_2628 (O_2628,N_28586,N_29002);
nor UO_2629 (O_2629,N_29341,N_29875);
or UO_2630 (O_2630,N_29144,N_29274);
nand UO_2631 (O_2631,N_29989,N_29292);
nor UO_2632 (O_2632,N_29185,N_29977);
nor UO_2633 (O_2633,N_28927,N_28676);
nand UO_2634 (O_2634,N_28886,N_28727);
xor UO_2635 (O_2635,N_29371,N_28999);
nor UO_2636 (O_2636,N_29056,N_29037);
and UO_2637 (O_2637,N_29326,N_28539);
nor UO_2638 (O_2638,N_29891,N_28504);
nand UO_2639 (O_2639,N_29144,N_28809);
xnor UO_2640 (O_2640,N_28806,N_29516);
or UO_2641 (O_2641,N_29454,N_29885);
xor UO_2642 (O_2642,N_29257,N_29799);
or UO_2643 (O_2643,N_29154,N_29720);
nand UO_2644 (O_2644,N_29523,N_28551);
nand UO_2645 (O_2645,N_29556,N_29893);
nand UO_2646 (O_2646,N_29952,N_28890);
nand UO_2647 (O_2647,N_29500,N_28565);
nor UO_2648 (O_2648,N_29312,N_29466);
xor UO_2649 (O_2649,N_29726,N_28807);
nor UO_2650 (O_2650,N_29381,N_29890);
and UO_2651 (O_2651,N_28571,N_29641);
or UO_2652 (O_2652,N_28628,N_28828);
or UO_2653 (O_2653,N_29115,N_28616);
nand UO_2654 (O_2654,N_29147,N_29326);
nand UO_2655 (O_2655,N_28584,N_29547);
nor UO_2656 (O_2656,N_28983,N_29784);
or UO_2657 (O_2657,N_29620,N_29806);
nand UO_2658 (O_2658,N_28818,N_29963);
xor UO_2659 (O_2659,N_28627,N_29028);
xor UO_2660 (O_2660,N_28804,N_29009);
nand UO_2661 (O_2661,N_29142,N_28910);
nand UO_2662 (O_2662,N_29920,N_29940);
nand UO_2663 (O_2663,N_28820,N_29392);
nand UO_2664 (O_2664,N_29503,N_28798);
xnor UO_2665 (O_2665,N_29755,N_29288);
and UO_2666 (O_2666,N_29401,N_29031);
nand UO_2667 (O_2667,N_29244,N_29754);
and UO_2668 (O_2668,N_29263,N_29047);
or UO_2669 (O_2669,N_29788,N_29284);
xor UO_2670 (O_2670,N_29029,N_29971);
nor UO_2671 (O_2671,N_28733,N_29716);
xnor UO_2672 (O_2672,N_29847,N_28566);
and UO_2673 (O_2673,N_28765,N_29357);
nand UO_2674 (O_2674,N_29942,N_28501);
nand UO_2675 (O_2675,N_29635,N_29720);
and UO_2676 (O_2676,N_29818,N_28869);
nor UO_2677 (O_2677,N_29207,N_28876);
and UO_2678 (O_2678,N_29384,N_29528);
or UO_2679 (O_2679,N_28987,N_29969);
and UO_2680 (O_2680,N_29274,N_29425);
nand UO_2681 (O_2681,N_28595,N_29930);
or UO_2682 (O_2682,N_29708,N_28729);
nand UO_2683 (O_2683,N_29273,N_28925);
xnor UO_2684 (O_2684,N_28914,N_28932);
and UO_2685 (O_2685,N_29503,N_29295);
and UO_2686 (O_2686,N_29816,N_29703);
xnor UO_2687 (O_2687,N_29938,N_29728);
xor UO_2688 (O_2688,N_29187,N_28953);
and UO_2689 (O_2689,N_29237,N_28625);
and UO_2690 (O_2690,N_29384,N_29020);
nand UO_2691 (O_2691,N_29280,N_28698);
xnor UO_2692 (O_2692,N_29876,N_29669);
xnor UO_2693 (O_2693,N_28851,N_28518);
nor UO_2694 (O_2694,N_29150,N_29768);
and UO_2695 (O_2695,N_29551,N_29584);
xnor UO_2696 (O_2696,N_29787,N_28539);
and UO_2697 (O_2697,N_29898,N_29540);
nor UO_2698 (O_2698,N_28881,N_29495);
or UO_2699 (O_2699,N_29663,N_29076);
or UO_2700 (O_2700,N_28807,N_29962);
nor UO_2701 (O_2701,N_29512,N_29648);
nor UO_2702 (O_2702,N_29234,N_29332);
xnor UO_2703 (O_2703,N_29468,N_29345);
xor UO_2704 (O_2704,N_28630,N_29291);
and UO_2705 (O_2705,N_29082,N_29660);
nor UO_2706 (O_2706,N_28555,N_28683);
nor UO_2707 (O_2707,N_29796,N_29347);
nand UO_2708 (O_2708,N_29036,N_29167);
nor UO_2709 (O_2709,N_28976,N_29084);
xnor UO_2710 (O_2710,N_28664,N_29511);
nand UO_2711 (O_2711,N_28923,N_29645);
xnor UO_2712 (O_2712,N_28810,N_29816);
nand UO_2713 (O_2713,N_29239,N_29184);
nand UO_2714 (O_2714,N_29607,N_29102);
nand UO_2715 (O_2715,N_29591,N_28939);
xor UO_2716 (O_2716,N_28961,N_28920);
or UO_2717 (O_2717,N_29968,N_28931);
nor UO_2718 (O_2718,N_28965,N_28870);
nand UO_2719 (O_2719,N_29383,N_29346);
nor UO_2720 (O_2720,N_29264,N_28600);
or UO_2721 (O_2721,N_28689,N_28619);
nand UO_2722 (O_2722,N_28711,N_29130);
nor UO_2723 (O_2723,N_29320,N_29869);
xnor UO_2724 (O_2724,N_29206,N_29167);
xnor UO_2725 (O_2725,N_29552,N_29596);
nand UO_2726 (O_2726,N_29873,N_28795);
and UO_2727 (O_2727,N_29809,N_29465);
nand UO_2728 (O_2728,N_29171,N_29008);
or UO_2729 (O_2729,N_29317,N_29206);
and UO_2730 (O_2730,N_29971,N_28667);
nand UO_2731 (O_2731,N_28810,N_29682);
nor UO_2732 (O_2732,N_29544,N_28660);
nand UO_2733 (O_2733,N_29582,N_28743);
nand UO_2734 (O_2734,N_28553,N_29236);
or UO_2735 (O_2735,N_29691,N_29521);
nand UO_2736 (O_2736,N_29081,N_28698);
nor UO_2737 (O_2737,N_28743,N_28976);
xnor UO_2738 (O_2738,N_28744,N_29388);
nand UO_2739 (O_2739,N_29677,N_29046);
or UO_2740 (O_2740,N_28567,N_29719);
xnor UO_2741 (O_2741,N_29662,N_29399);
xnor UO_2742 (O_2742,N_29579,N_29651);
and UO_2743 (O_2743,N_29123,N_29554);
xor UO_2744 (O_2744,N_29503,N_28728);
nand UO_2745 (O_2745,N_29137,N_29669);
nand UO_2746 (O_2746,N_29125,N_29863);
nor UO_2747 (O_2747,N_28910,N_29606);
or UO_2748 (O_2748,N_29867,N_28506);
nand UO_2749 (O_2749,N_28915,N_29897);
or UO_2750 (O_2750,N_29656,N_28889);
and UO_2751 (O_2751,N_29919,N_29435);
nor UO_2752 (O_2752,N_28599,N_28891);
and UO_2753 (O_2753,N_29896,N_28985);
nor UO_2754 (O_2754,N_29459,N_29111);
or UO_2755 (O_2755,N_28599,N_28518);
nor UO_2756 (O_2756,N_29106,N_29769);
xnor UO_2757 (O_2757,N_28604,N_29712);
and UO_2758 (O_2758,N_29050,N_29936);
xnor UO_2759 (O_2759,N_29293,N_29614);
and UO_2760 (O_2760,N_29008,N_29088);
or UO_2761 (O_2761,N_28843,N_29587);
xnor UO_2762 (O_2762,N_29625,N_29108);
xor UO_2763 (O_2763,N_29885,N_29572);
and UO_2764 (O_2764,N_29965,N_29262);
and UO_2765 (O_2765,N_28549,N_29602);
or UO_2766 (O_2766,N_29715,N_28919);
or UO_2767 (O_2767,N_29825,N_28791);
nand UO_2768 (O_2768,N_28735,N_29028);
or UO_2769 (O_2769,N_29988,N_29807);
nand UO_2770 (O_2770,N_29397,N_28617);
nor UO_2771 (O_2771,N_29201,N_29138);
or UO_2772 (O_2772,N_28615,N_28897);
or UO_2773 (O_2773,N_28697,N_29099);
xor UO_2774 (O_2774,N_28872,N_29712);
or UO_2775 (O_2775,N_29933,N_29029);
nor UO_2776 (O_2776,N_29952,N_29403);
nor UO_2777 (O_2777,N_29560,N_29921);
nand UO_2778 (O_2778,N_29635,N_29426);
and UO_2779 (O_2779,N_28707,N_29481);
nand UO_2780 (O_2780,N_29860,N_29903);
xnor UO_2781 (O_2781,N_29708,N_28786);
xnor UO_2782 (O_2782,N_29400,N_28732);
xnor UO_2783 (O_2783,N_29652,N_29783);
and UO_2784 (O_2784,N_29689,N_29406);
and UO_2785 (O_2785,N_28817,N_29207);
and UO_2786 (O_2786,N_29917,N_29743);
and UO_2787 (O_2787,N_29502,N_28512);
xnor UO_2788 (O_2788,N_28978,N_28857);
nand UO_2789 (O_2789,N_29241,N_29100);
or UO_2790 (O_2790,N_29383,N_29663);
xnor UO_2791 (O_2791,N_28681,N_29865);
xor UO_2792 (O_2792,N_29610,N_29240);
nand UO_2793 (O_2793,N_28691,N_28980);
and UO_2794 (O_2794,N_29389,N_28689);
xor UO_2795 (O_2795,N_29466,N_29820);
xnor UO_2796 (O_2796,N_28972,N_28920);
nor UO_2797 (O_2797,N_29429,N_29188);
and UO_2798 (O_2798,N_28623,N_29995);
and UO_2799 (O_2799,N_29010,N_29576);
nand UO_2800 (O_2800,N_29742,N_29265);
nor UO_2801 (O_2801,N_29799,N_29426);
and UO_2802 (O_2802,N_28727,N_29271);
nand UO_2803 (O_2803,N_29815,N_29788);
or UO_2804 (O_2804,N_29124,N_29348);
and UO_2805 (O_2805,N_29320,N_29851);
xor UO_2806 (O_2806,N_28667,N_29073);
and UO_2807 (O_2807,N_28990,N_29255);
or UO_2808 (O_2808,N_28750,N_28895);
and UO_2809 (O_2809,N_29857,N_29764);
xnor UO_2810 (O_2810,N_28986,N_29784);
nor UO_2811 (O_2811,N_29682,N_29582);
nor UO_2812 (O_2812,N_29795,N_29456);
nor UO_2813 (O_2813,N_28554,N_28923);
or UO_2814 (O_2814,N_28849,N_28673);
and UO_2815 (O_2815,N_29232,N_28564);
nor UO_2816 (O_2816,N_29378,N_28804);
xnor UO_2817 (O_2817,N_29532,N_29047);
xnor UO_2818 (O_2818,N_29441,N_29916);
nand UO_2819 (O_2819,N_29156,N_29516);
nand UO_2820 (O_2820,N_29163,N_29343);
nand UO_2821 (O_2821,N_28620,N_28674);
nor UO_2822 (O_2822,N_28828,N_29851);
and UO_2823 (O_2823,N_28515,N_28989);
xnor UO_2824 (O_2824,N_29146,N_29296);
and UO_2825 (O_2825,N_28528,N_28772);
and UO_2826 (O_2826,N_29640,N_29000);
nand UO_2827 (O_2827,N_29868,N_28793);
xnor UO_2828 (O_2828,N_29002,N_29004);
and UO_2829 (O_2829,N_28991,N_29638);
or UO_2830 (O_2830,N_29836,N_28647);
or UO_2831 (O_2831,N_29294,N_29616);
nand UO_2832 (O_2832,N_29835,N_29983);
and UO_2833 (O_2833,N_28613,N_29390);
xnor UO_2834 (O_2834,N_29990,N_28621);
and UO_2835 (O_2835,N_29143,N_29348);
nand UO_2836 (O_2836,N_29855,N_29347);
xor UO_2837 (O_2837,N_28949,N_29001);
nand UO_2838 (O_2838,N_28503,N_29035);
xnor UO_2839 (O_2839,N_29058,N_28590);
nand UO_2840 (O_2840,N_29346,N_29563);
nor UO_2841 (O_2841,N_28873,N_29859);
xnor UO_2842 (O_2842,N_28530,N_29511);
xnor UO_2843 (O_2843,N_29508,N_29738);
nand UO_2844 (O_2844,N_29908,N_29952);
nand UO_2845 (O_2845,N_28946,N_29958);
or UO_2846 (O_2846,N_28828,N_29256);
xnor UO_2847 (O_2847,N_29088,N_28942);
and UO_2848 (O_2848,N_29320,N_29259);
nand UO_2849 (O_2849,N_29222,N_28992);
or UO_2850 (O_2850,N_29422,N_29604);
or UO_2851 (O_2851,N_29124,N_29274);
nand UO_2852 (O_2852,N_28719,N_28637);
or UO_2853 (O_2853,N_29827,N_29321);
xnor UO_2854 (O_2854,N_29463,N_29150);
xor UO_2855 (O_2855,N_28601,N_29438);
nand UO_2856 (O_2856,N_28868,N_29559);
or UO_2857 (O_2857,N_29994,N_28820);
nand UO_2858 (O_2858,N_29169,N_29010);
and UO_2859 (O_2859,N_28871,N_29179);
xnor UO_2860 (O_2860,N_29599,N_29991);
nand UO_2861 (O_2861,N_29222,N_29563);
nand UO_2862 (O_2862,N_29360,N_28825);
xnor UO_2863 (O_2863,N_28938,N_29989);
and UO_2864 (O_2864,N_29327,N_29491);
or UO_2865 (O_2865,N_29365,N_28846);
nor UO_2866 (O_2866,N_29661,N_29779);
nand UO_2867 (O_2867,N_29241,N_28975);
and UO_2868 (O_2868,N_29603,N_29652);
and UO_2869 (O_2869,N_29999,N_29237);
nand UO_2870 (O_2870,N_28966,N_28561);
nor UO_2871 (O_2871,N_29884,N_28687);
xnor UO_2872 (O_2872,N_29271,N_29966);
nor UO_2873 (O_2873,N_29587,N_29461);
xor UO_2874 (O_2874,N_29720,N_28880);
xor UO_2875 (O_2875,N_29306,N_29796);
and UO_2876 (O_2876,N_29351,N_29747);
and UO_2877 (O_2877,N_29205,N_28871);
nor UO_2878 (O_2878,N_29977,N_29309);
nand UO_2879 (O_2879,N_29560,N_29929);
nor UO_2880 (O_2880,N_29497,N_29191);
xor UO_2881 (O_2881,N_29575,N_29365);
nor UO_2882 (O_2882,N_28857,N_29711);
nand UO_2883 (O_2883,N_29049,N_28578);
and UO_2884 (O_2884,N_28570,N_29954);
xor UO_2885 (O_2885,N_28877,N_28698);
or UO_2886 (O_2886,N_29714,N_29015);
nand UO_2887 (O_2887,N_29839,N_29017);
nand UO_2888 (O_2888,N_29357,N_29183);
nand UO_2889 (O_2889,N_29326,N_28937);
xnor UO_2890 (O_2890,N_29364,N_29606);
or UO_2891 (O_2891,N_28879,N_28867);
nand UO_2892 (O_2892,N_28522,N_29713);
and UO_2893 (O_2893,N_29282,N_29088);
xor UO_2894 (O_2894,N_29796,N_29275);
xor UO_2895 (O_2895,N_28890,N_28539);
nor UO_2896 (O_2896,N_28932,N_29009);
nor UO_2897 (O_2897,N_29737,N_28982);
nand UO_2898 (O_2898,N_28932,N_29661);
xnor UO_2899 (O_2899,N_29414,N_29257);
xnor UO_2900 (O_2900,N_29955,N_28807);
nand UO_2901 (O_2901,N_29392,N_29998);
or UO_2902 (O_2902,N_29216,N_29879);
nor UO_2903 (O_2903,N_28742,N_29135);
nand UO_2904 (O_2904,N_29643,N_29030);
and UO_2905 (O_2905,N_29139,N_28845);
nand UO_2906 (O_2906,N_29925,N_29971);
xor UO_2907 (O_2907,N_28676,N_28508);
nand UO_2908 (O_2908,N_29479,N_29882);
and UO_2909 (O_2909,N_28908,N_28872);
or UO_2910 (O_2910,N_28629,N_29673);
or UO_2911 (O_2911,N_29366,N_29783);
nand UO_2912 (O_2912,N_29590,N_29071);
xnor UO_2913 (O_2913,N_29911,N_28601);
or UO_2914 (O_2914,N_29311,N_28940);
or UO_2915 (O_2915,N_29006,N_29564);
xor UO_2916 (O_2916,N_29612,N_29164);
xnor UO_2917 (O_2917,N_29142,N_29136);
nor UO_2918 (O_2918,N_29255,N_29058);
and UO_2919 (O_2919,N_28579,N_29461);
nand UO_2920 (O_2920,N_28831,N_29480);
or UO_2921 (O_2921,N_29410,N_29203);
and UO_2922 (O_2922,N_29330,N_28556);
nor UO_2923 (O_2923,N_29569,N_29208);
nand UO_2924 (O_2924,N_29401,N_28980);
nand UO_2925 (O_2925,N_29414,N_29026);
nor UO_2926 (O_2926,N_29845,N_28968);
or UO_2927 (O_2927,N_29723,N_29199);
nand UO_2928 (O_2928,N_28740,N_28788);
nor UO_2929 (O_2929,N_28500,N_29555);
nor UO_2930 (O_2930,N_28938,N_29371);
nor UO_2931 (O_2931,N_29821,N_29349);
nand UO_2932 (O_2932,N_29891,N_28900);
and UO_2933 (O_2933,N_29880,N_29117);
nor UO_2934 (O_2934,N_29095,N_28726);
nor UO_2935 (O_2935,N_28758,N_29350);
nand UO_2936 (O_2936,N_29129,N_29942);
nand UO_2937 (O_2937,N_29038,N_29971);
xor UO_2938 (O_2938,N_29136,N_28532);
nor UO_2939 (O_2939,N_29383,N_29322);
and UO_2940 (O_2940,N_29891,N_28839);
xnor UO_2941 (O_2941,N_29655,N_29114);
and UO_2942 (O_2942,N_29006,N_29958);
nand UO_2943 (O_2943,N_29834,N_29730);
xnor UO_2944 (O_2944,N_29257,N_29917);
or UO_2945 (O_2945,N_28742,N_29957);
nand UO_2946 (O_2946,N_29583,N_29678);
and UO_2947 (O_2947,N_28670,N_29637);
nand UO_2948 (O_2948,N_28523,N_29505);
xnor UO_2949 (O_2949,N_29913,N_29183);
nand UO_2950 (O_2950,N_29897,N_29307);
and UO_2951 (O_2951,N_28513,N_29083);
xnor UO_2952 (O_2952,N_29822,N_28989);
and UO_2953 (O_2953,N_28638,N_29466);
nand UO_2954 (O_2954,N_29311,N_28546);
nor UO_2955 (O_2955,N_29851,N_29627);
nor UO_2956 (O_2956,N_29734,N_28975);
and UO_2957 (O_2957,N_28943,N_28987);
nand UO_2958 (O_2958,N_29488,N_29276);
nor UO_2959 (O_2959,N_29122,N_28924);
xor UO_2960 (O_2960,N_29258,N_28836);
or UO_2961 (O_2961,N_29322,N_28636);
xor UO_2962 (O_2962,N_29371,N_29588);
xnor UO_2963 (O_2963,N_29006,N_29913);
or UO_2964 (O_2964,N_29360,N_28786);
xor UO_2965 (O_2965,N_29558,N_28907);
and UO_2966 (O_2966,N_29866,N_29606);
nand UO_2967 (O_2967,N_28981,N_28980);
or UO_2968 (O_2968,N_29862,N_28976);
xor UO_2969 (O_2969,N_29175,N_29144);
nor UO_2970 (O_2970,N_29891,N_29749);
nand UO_2971 (O_2971,N_28950,N_29632);
nor UO_2972 (O_2972,N_28912,N_29438);
xor UO_2973 (O_2973,N_29293,N_29581);
or UO_2974 (O_2974,N_29509,N_29571);
nor UO_2975 (O_2975,N_29412,N_29081);
and UO_2976 (O_2976,N_29374,N_29220);
nor UO_2977 (O_2977,N_29086,N_28576);
xor UO_2978 (O_2978,N_28731,N_29430);
nand UO_2979 (O_2979,N_28693,N_29490);
nand UO_2980 (O_2980,N_29142,N_29211);
nand UO_2981 (O_2981,N_29766,N_29793);
nand UO_2982 (O_2982,N_28945,N_28993);
nand UO_2983 (O_2983,N_28777,N_28806);
nor UO_2984 (O_2984,N_29170,N_28800);
xnor UO_2985 (O_2985,N_29269,N_29712);
and UO_2986 (O_2986,N_29341,N_29071);
nand UO_2987 (O_2987,N_29255,N_29818);
xor UO_2988 (O_2988,N_28711,N_29111);
nand UO_2989 (O_2989,N_28535,N_29468);
xnor UO_2990 (O_2990,N_29708,N_29845);
nor UO_2991 (O_2991,N_29145,N_28612);
nand UO_2992 (O_2992,N_29437,N_29793);
xnor UO_2993 (O_2993,N_28663,N_29440);
nand UO_2994 (O_2994,N_29618,N_29143);
and UO_2995 (O_2995,N_29549,N_29808);
nand UO_2996 (O_2996,N_28806,N_29552);
or UO_2997 (O_2997,N_29823,N_29527);
nor UO_2998 (O_2998,N_29829,N_29790);
or UO_2999 (O_2999,N_28835,N_28993);
xnor UO_3000 (O_3000,N_28559,N_29569);
nor UO_3001 (O_3001,N_29771,N_29567);
nand UO_3002 (O_3002,N_28647,N_29247);
or UO_3003 (O_3003,N_29258,N_29912);
nor UO_3004 (O_3004,N_28594,N_28910);
nor UO_3005 (O_3005,N_29512,N_28591);
nand UO_3006 (O_3006,N_29804,N_29482);
nor UO_3007 (O_3007,N_29543,N_29420);
and UO_3008 (O_3008,N_28900,N_29632);
and UO_3009 (O_3009,N_29081,N_29847);
and UO_3010 (O_3010,N_29570,N_28965);
and UO_3011 (O_3011,N_29124,N_28766);
xor UO_3012 (O_3012,N_29910,N_29768);
or UO_3013 (O_3013,N_29134,N_28927);
xnor UO_3014 (O_3014,N_29349,N_28557);
and UO_3015 (O_3015,N_29638,N_29848);
nor UO_3016 (O_3016,N_28796,N_28523);
or UO_3017 (O_3017,N_28694,N_28798);
and UO_3018 (O_3018,N_29665,N_29038);
or UO_3019 (O_3019,N_28902,N_29060);
and UO_3020 (O_3020,N_29146,N_29751);
xnor UO_3021 (O_3021,N_29693,N_29771);
xnor UO_3022 (O_3022,N_29631,N_29727);
nand UO_3023 (O_3023,N_28868,N_29060);
and UO_3024 (O_3024,N_29076,N_29243);
xnor UO_3025 (O_3025,N_29762,N_29363);
xnor UO_3026 (O_3026,N_28906,N_29507);
or UO_3027 (O_3027,N_28925,N_28545);
and UO_3028 (O_3028,N_28836,N_29349);
xor UO_3029 (O_3029,N_28517,N_29728);
xnor UO_3030 (O_3030,N_28779,N_28992);
nand UO_3031 (O_3031,N_29669,N_29617);
xnor UO_3032 (O_3032,N_28929,N_28806);
or UO_3033 (O_3033,N_29929,N_29378);
or UO_3034 (O_3034,N_29909,N_29009);
nand UO_3035 (O_3035,N_28539,N_29382);
nand UO_3036 (O_3036,N_28967,N_28919);
nor UO_3037 (O_3037,N_29591,N_28895);
and UO_3038 (O_3038,N_29358,N_28555);
nand UO_3039 (O_3039,N_28740,N_28911);
nand UO_3040 (O_3040,N_29528,N_29770);
nand UO_3041 (O_3041,N_29506,N_29452);
or UO_3042 (O_3042,N_28946,N_28669);
xor UO_3043 (O_3043,N_29886,N_28864);
nor UO_3044 (O_3044,N_29031,N_29353);
nor UO_3045 (O_3045,N_28629,N_29876);
nor UO_3046 (O_3046,N_29772,N_28524);
xor UO_3047 (O_3047,N_28699,N_29967);
xnor UO_3048 (O_3048,N_29511,N_28715);
xnor UO_3049 (O_3049,N_28760,N_29651);
nand UO_3050 (O_3050,N_29483,N_29219);
xor UO_3051 (O_3051,N_29200,N_29387);
xor UO_3052 (O_3052,N_29715,N_29936);
and UO_3053 (O_3053,N_29328,N_29179);
or UO_3054 (O_3054,N_29946,N_28506);
nand UO_3055 (O_3055,N_29737,N_29699);
nor UO_3056 (O_3056,N_29660,N_29693);
xor UO_3057 (O_3057,N_29037,N_29978);
nand UO_3058 (O_3058,N_28985,N_28849);
and UO_3059 (O_3059,N_28588,N_28944);
and UO_3060 (O_3060,N_29208,N_29402);
xnor UO_3061 (O_3061,N_28565,N_28527);
nand UO_3062 (O_3062,N_28585,N_28714);
or UO_3063 (O_3063,N_29691,N_29944);
nor UO_3064 (O_3064,N_29167,N_29669);
nand UO_3065 (O_3065,N_28539,N_29924);
or UO_3066 (O_3066,N_29687,N_28708);
nor UO_3067 (O_3067,N_29276,N_29884);
and UO_3068 (O_3068,N_29200,N_28803);
nand UO_3069 (O_3069,N_29190,N_29615);
nor UO_3070 (O_3070,N_29448,N_29970);
or UO_3071 (O_3071,N_29970,N_29152);
nand UO_3072 (O_3072,N_29577,N_28853);
xor UO_3073 (O_3073,N_29701,N_29011);
and UO_3074 (O_3074,N_29684,N_28533);
nor UO_3075 (O_3075,N_29151,N_28660);
or UO_3076 (O_3076,N_28799,N_28737);
or UO_3077 (O_3077,N_28611,N_29785);
and UO_3078 (O_3078,N_29309,N_28747);
xor UO_3079 (O_3079,N_29121,N_29646);
xnor UO_3080 (O_3080,N_29373,N_29438);
and UO_3081 (O_3081,N_29514,N_29455);
nor UO_3082 (O_3082,N_29355,N_29425);
nand UO_3083 (O_3083,N_29806,N_29783);
and UO_3084 (O_3084,N_29690,N_29316);
nor UO_3085 (O_3085,N_29446,N_28561);
xor UO_3086 (O_3086,N_29558,N_29118);
or UO_3087 (O_3087,N_29489,N_28598);
xor UO_3088 (O_3088,N_29524,N_29558);
xnor UO_3089 (O_3089,N_28600,N_28553);
nor UO_3090 (O_3090,N_29050,N_28808);
nand UO_3091 (O_3091,N_29658,N_29312);
nand UO_3092 (O_3092,N_29239,N_28972);
nor UO_3093 (O_3093,N_28989,N_28828);
or UO_3094 (O_3094,N_28627,N_28838);
or UO_3095 (O_3095,N_29006,N_29235);
or UO_3096 (O_3096,N_28537,N_28727);
xor UO_3097 (O_3097,N_28660,N_29799);
xnor UO_3098 (O_3098,N_29571,N_29209);
and UO_3099 (O_3099,N_29778,N_29467);
xor UO_3100 (O_3100,N_29623,N_29915);
nand UO_3101 (O_3101,N_28837,N_28923);
nor UO_3102 (O_3102,N_29010,N_28981);
nand UO_3103 (O_3103,N_29302,N_29906);
and UO_3104 (O_3104,N_28647,N_28782);
and UO_3105 (O_3105,N_29479,N_28965);
and UO_3106 (O_3106,N_29094,N_28911);
nand UO_3107 (O_3107,N_29715,N_29437);
nor UO_3108 (O_3108,N_28859,N_29605);
or UO_3109 (O_3109,N_29222,N_29257);
nand UO_3110 (O_3110,N_28621,N_29983);
xor UO_3111 (O_3111,N_29603,N_29217);
nand UO_3112 (O_3112,N_29747,N_29180);
and UO_3113 (O_3113,N_28765,N_29431);
or UO_3114 (O_3114,N_28946,N_29028);
or UO_3115 (O_3115,N_29286,N_29479);
or UO_3116 (O_3116,N_28669,N_28606);
and UO_3117 (O_3117,N_28579,N_29582);
xor UO_3118 (O_3118,N_29680,N_29628);
and UO_3119 (O_3119,N_28983,N_28671);
or UO_3120 (O_3120,N_28896,N_29425);
xor UO_3121 (O_3121,N_29834,N_29099);
and UO_3122 (O_3122,N_29080,N_29702);
or UO_3123 (O_3123,N_28931,N_29463);
nor UO_3124 (O_3124,N_28984,N_29149);
and UO_3125 (O_3125,N_28522,N_28889);
or UO_3126 (O_3126,N_28614,N_29518);
nor UO_3127 (O_3127,N_29938,N_28920);
nand UO_3128 (O_3128,N_29248,N_28983);
xnor UO_3129 (O_3129,N_29744,N_29851);
nand UO_3130 (O_3130,N_29722,N_28578);
nor UO_3131 (O_3131,N_29629,N_29882);
nand UO_3132 (O_3132,N_28564,N_29009);
xor UO_3133 (O_3133,N_29461,N_29428);
or UO_3134 (O_3134,N_29999,N_29777);
xor UO_3135 (O_3135,N_29520,N_29504);
nand UO_3136 (O_3136,N_29189,N_29924);
nor UO_3137 (O_3137,N_29915,N_28843);
or UO_3138 (O_3138,N_29333,N_29385);
and UO_3139 (O_3139,N_29071,N_29450);
xor UO_3140 (O_3140,N_28739,N_29279);
nor UO_3141 (O_3141,N_28954,N_29690);
nand UO_3142 (O_3142,N_29046,N_28968);
and UO_3143 (O_3143,N_28818,N_29275);
xnor UO_3144 (O_3144,N_28748,N_29545);
nand UO_3145 (O_3145,N_29974,N_28682);
or UO_3146 (O_3146,N_28608,N_29528);
and UO_3147 (O_3147,N_29731,N_29816);
nand UO_3148 (O_3148,N_29849,N_29315);
and UO_3149 (O_3149,N_29426,N_29460);
or UO_3150 (O_3150,N_29034,N_29587);
or UO_3151 (O_3151,N_28960,N_29549);
or UO_3152 (O_3152,N_29337,N_29688);
xnor UO_3153 (O_3153,N_29436,N_29058);
xor UO_3154 (O_3154,N_28840,N_28926);
xor UO_3155 (O_3155,N_29324,N_28643);
or UO_3156 (O_3156,N_29011,N_29735);
or UO_3157 (O_3157,N_28623,N_29735);
nand UO_3158 (O_3158,N_29716,N_28667);
nor UO_3159 (O_3159,N_29044,N_28963);
and UO_3160 (O_3160,N_28735,N_28936);
or UO_3161 (O_3161,N_28926,N_29268);
or UO_3162 (O_3162,N_28518,N_28860);
nor UO_3163 (O_3163,N_29423,N_29564);
or UO_3164 (O_3164,N_28755,N_29027);
xnor UO_3165 (O_3165,N_28676,N_29763);
or UO_3166 (O_3166,N_29549,N_29851);
or UO_3167 (O_3167,N_29366,N_28871);
or UO_3168 (O_3168,N_29581,N_29654);
xnor UO_3169 (O_3169,N_28544,N_29265);
nand UO_3170 (O_3170,N_28907,N_29987);
and UO_3171 (O_3171,N_29854,N_29112);
or UO_3172 (O_3172,N_29441,N_29848);
and UO_3173 (O_3173,N_29141,N_29931);
or UO_3174 (O_3174,N_29093,N_29857);
nand UO_3175 (O_3175,N_29967,N_28939);
or UO_3176 (O_3176,N_29970,N_28566);
and UO_3177 (O_3177,N_29613,N_29464);
nand UO_3178 (O_3178,N_29667,N_28954);
xnor UO_3179 (O_3179,N_29758,N_29862);
nor UO_3180 (O_3180,N_29381,N_29826);
nand UO_3181 (O_3181,N_28552,N_28919);
xnor UO_3182 (O_3182,N_28924,N_29839);
nor UO_3183 (O_3183,N_29330,N_28863);
and UO_3184 (O_3184,N_29835,N_28575);
or UO_3185 (O_3185,N_29219,N_28683);
and UO_3186 (O_3186,N_29944,N_29635);
xor UO_3187 (O_3187,N_28772,N_29015);
or UO_3188 (O_3188,N_29597,N_28903);
xor UO_3189 (O_3189,N_29009,N_29059);
xnor UO_3190 (O_3190,N_29064,N_28848);
xor UO_3191 (O_3191,N_29898,N_29469);
xor UO_3192 (O_3192,N_28781,N_29349);
nor UO_3193 (O_3193,N_28855,N_28993);
nor UO_3194 (O_3194,N_29061,N_28512);
nor UO_3195 (O_3195,N_29527,N_28715);
nor UO_3196 (O_3196,N_29446,N_28819);
xnor UO_3197 (O_3197,N_29202,N_29656);
nand UO_3198 (O_3198,N_28881,N_29762);
nand UO_3199 (O_3199,N_29767,N_28926);
or UO_3200 (O_3200,N_29598,N_29321);
xnor UO_3201 (O_3201,N_29567,N_29658);
nor UO_3202 (O_3202,N_29830,N_29494);
or UO_3203 (O_3203,N_29201,N_28887);
nand UO_3204 (O_3204,N_29039,N_28552);
and UO_3205 (O_3205,N_29896,N_28513);
nand UO_3206 (O_3206,N_29487,N_29087);
or UO_3207 (O_3207,N_28540,N_29182);
nor UO_3208 (O_3208,N_28530,N_28688);
nand UO_3209 (O_3209,N_29656,N_29851);
or UO_3210 (O_3210,N_29565,N_28804);
or UO_3211 (O_3211,N_28895,N_29925);
or UO_3212 (O_3212,N_28895,N_29133);
xor UO_3213 (O_3213,N_28952,N_29862);
nor UO_3214 (O_3214,N_29460,N_29958);
and UO_3215 (O_3215,N_29172,N_29528);
nand UO_3216 (O_3216,N_29063,N_28988);
and UO_3217 (O_3217,N_29604,N_28512);
or UO_3218 (O_3218,N_28652,N_28943);
and UO_3219 (O_3219,N_29362,N_28675);
nor UO_3220 (O_3220,N_29699,N_28598);
or UO_3221 (O_3221,N_29792,N_29031);
xnor UO_3222 (O_3222,N_29360,N_29625);
nand UO_3223 (O_3223,N_29252,N_29530);
nor UO_3224 (O_3224,N_29442,N_29256);
nor UO_3225 (O_3225,N_28516,N_29583);
or UO_3226 (O_3226,N_28836,N_29505);
and UO_3227 (O_3227,N_29680,N_29678);
xnor UO_3228 (O_3228,N_29844,N_29363);
xor UO_3229 (O_3229,N_29262,N_28982);
nand UO_3230 (O_3230,N_28893,N_28802);
or UO_3231 (O_3231,N_29534,N_29798);
xnor UO_3232 (O_3232,N_29714,N_29065);
xor UO_3233 (O_3233,N_29471,N_29793);
or UO_3234 (O_3234,N_28990,N_29732);
and UO_3235 (O_3235,N_29094,N_29424);
xor UO_3236 (O_3236,N_29525,N_29388);
xnor UO_3237 (O_3237,N_29071,N_29067);
or UO_3238 (O_3238,N_29181,N_29921);
nand UO_3239 (O_3239,N_29924,N_28548);
xnor UO_3240 (O_3240,N_29206,N_29458);
and UO_3241 (O_3241,N_29796,N_29774);
and UO_3242 (O_3242,N_28501,N_29149);
xnor UO_3243 (O_3243,N_28973,N_29639);
nand UO_3244 (O_3244,N_28959,N_29660);
nand UO_3245 (O_3245,N_29428,N_29245);
and UO_3246 (O_3246,N_29891,N_29448);
nand UO_3247 (O_3247,N_29967,N_28692);
xnor UO_3248 (O_3248,N_29060,N_29606);
nand UO_3249 (O_3249,N_28643,N_28702);
and UO_3250 (O_3250,N_28592,N_28764);
or UO_3251 (O_3251,N_29168,N_29281);
nand UO_3252 (O_3252,N_29311,N_28947);
or UO_3253 (O_3253,N_29093,N_28704);
xor UO_3254 (O_3254,N_29838,N_29872);
nor UO_3255 (O_3255,N_29358,N_29008);
nor UO_3256 (O_3256,N_28619,N_29767);
nor UO_3257 (O_3257,N_29379,N_29016);
nand UO_3258 (O_3258,N_28876,N_29049);
nor UO_3259 (O_3259,N_29504,N_28975);
nand UO_3260 (O_3260,N_28791,N_29000);
xor UO_3261 (O_3261,N_28778,N_29259);
xor UO_3262 (O_3262,N_29310,N_29555);
nor UO_3263 (O_3263,N_29167,N_28690);
or UO_3264 (O_3264,N_29897,N_29447);
and UO_3265 (O_3265,N_29183,N_29596);
nand UO_3266 (O_3266,N_29715,N_29196);
nand UO_3267 (O_3267,N_28815,N_29036);
or UO_3268 (O_3268,N_28957,N_29584);
and UO_3269 (O_3269,N_29094,N_29372);
nand UO_3270 (O_3270,N_29996,N_29500);
nand UO_3271 (O_3271,N_29878,N_29439);
or UO_3272 (O_3272,N_29820,N_28848);
nand UO_3273 (O_3273,N_29522,N_28704);
and UO_3274 (O_3274,N_28920,N_29099);
xor UO_3275 (O_3275,N_29304,N_29979);
and UO_3276 (O_3276,N_29511,N_29500);
xor UO_3277 (O_3277,N_28676,N_29307);
and UO_3278 (O_3278,N_29868,N_29519);
nand UO_3279 (O_3279,N_28866,N_29348);
xor UO_3280 (O_3280,N_29622,N_28824);
xor UO_3281 (O_3281,N_29400,N_28736);
nand UO_3282 (O_3282,N_29607,N_28664);
nand UO_3283 (O_3283,N_29759,N_29805);
and UO_3284 (O_3284,N_28654,N_29872);
or UO_3285 (O_3285,N_28573,N_28649);
nand UO_3286 (O_3286,N_29396,N_29524);
and UO_3287 (O_3287,N_29697,N_28752);
or UO_3288 (O_3288,N_28580,N_28684);
nand UO_3289 (O_3289,N_28993,N_29206);
nand UO_3290 (O_3290,N_29327,N_29453);
xor UO_3291 (O_3291,N_29479,N_29172);
xnor UO_3292 (O_3292,N_29048,N_28803);
nand UO_3293 (O_3293,N_28690,N_29175);
or UO_3294 (O_3294,N_28752,N_29635);
and UO_3295 (O_3295,N_29191,N_29066);
nor UO_3296 (O_3296,N_28888,N_29969);
or UO_3297 (O_3297,N_29190,N_29137);
and UO_3298 (O_3298,N_28765,N_28746);
xor UO_3299 (O_3299,N_28727,N_29979);
xnor UO_3300 (O_3300,N_29724,N_29695);
nor UO_3301 (O_3301,N_28836,N_29806);
xnor UO_3302 (O_3302,N_28567,N_29259);
and UO_3303 (O_3303,N_28945,N_29640);
and UO_3304 (O_3304,N_28885,N_29507);
nand UO_3305 (O_3305,N_29950,N_29219);
nand UO_3306 (O_3306,N_29398,N_29013);
and UO_3307 (O_3307,N_29924,N_29178);
nor UO_3308 (O_3308,N_29949,N_29506);
or UO_3309 (O_3309,N_28982,N_29211);
xnor UO_3310 (O_3310,N_29373,N_29583);
or UO_3311 (O_3311,N_29633,N_29454);
nor UO_3312 (O_3312,N_28724,N_29633);
or UO_3313 (O_3313,N_29913,N_28588);
nor UO_3314 (O_3314,N_29917,N_29932);
nand UO_3315 (O_3315,N_29862,N_29791);
xor UO_3316 (O_3316,N_29991,N_28544);
and UO_3317 (O_3317,N_28737,N_29689);
xnor UO_3318 (O_3318,N_28884,N_29275);
or UO_3319 (O_3319,N_29045,N_29057);
nand UO_3320 (O_3320,N_28519,N_28641);
xor UO_3321 (O_3321,N_29055,N_29523);
and UO_3322 (O_3322,N_29169,N_29472);
xor UO_3323 (O_3323,N_29672,N_29019);
nor UO_3324 (O_3324,N_29316,N_28651);
or UO_3325 (O_3325,N_29323,N_29232);
nand UO_3326 (O_3326,N_28889,N_29325);
nor UO_3327 (O_3327,N_29047,N_29205);
or UO_3328 (O_3328,N_28703,N_29005);
xnor UO_3329 (O_3329,N_28523,N_29434);
nor UO_3330 (O_3330,N_29807,N_29624);
and UO_3331 (O_3331,N_28654,N_29657);
or UO_3332 (O_3332,N_29449,N_29569);
nor UO_3333 (O_3333,N_29527,N_29254);
nand UO_3334 (O_3334,N_29602,N_29269);
nand UO_3335 (O_3335,N_28851,N_29704);
nand UO_3336 (O_3336,N_28768,N_28950);
nand UO_3337 (O_3337,N_28764,N_29234);
or UO_3338 (O_3338,N_29793,N_29957);
and UO_3339 (O_3339,N_28945,N_29695);
nor UO_3340 (O_3340,N_28534,N_28585);
or UO_3341 (O_3341,N_28517,N_29066);
and UO_3342 (O_3342,N_29116,N_29611);
or UO_3343 (O_3343,N_28532,N_29583);
or UO_3344 (O_3344,N_29220,N_29680);
nor UO_3345 (O_3345,N_29520,N_29471);
nand UO_3346 (O_3346,N_28884,N_29579);
nor UO_3347 (O_3347,N_28654,N_28962);
nand UO_3348 (O_3348,N_29333,N_28672);
xnor UO_3349 (O_3349,N_29098,N_28985);
and UO_3350 (O_3350,N_29834,N_29654);
xnor UO_3351 (O_3351,N_29569,N_28723);
and UO_3352 (O_3352,N_29696,N_29675);
nand UO_3353 (O_3353,N_29487,N_28775);
or UO_3354 (O_3354,N_29081,N_29696);
and UO_3355 (O_3355,N_29453,N_29983);
nor UO_3356 (O_3356,N_29484,N_29185);
xor UO_3357 (O_3357,N_29934,N_28726);
and UO_3358 (O_3358,N_29599,N_28964);
nand UO_3359 (O_3359,N_28586,N_29936);
xnor UO_3360 (O_3360,N_29811,N_29007);
nor UO_3361 (O_3361,N_29030,N_29545);
nand UO_3362 (O_3362,N_28517,N_29150);
nor UO_3363 (O_3363,N_29547,N_29134);
nand UO_3364 (O_3364,N_29971,N_28855);
nor UO_3365 (O_3365,N_29401,N_29124);
nor UO_3366 (O_3366,N_29822,N_28729);
or UO_3367 (O_3367,N_29724,N_29964);
nor UO_3368 (O_3368,N_29841,N_29506);
xor UO_3369 (O_3369,N_29841,N_29840);
or UO_3370 (O_3370,N_28569,N_29914);
nor UO_3371 (O_3371,N_29219,N_29258);
xnor UO_3372 (O_3372,N_28648,N_28804);
xnor UO_3373 (O_3373,N_29254,N_29543);
nand UO_3374 (O_3374,N_29953,N_28802);
nor UO_3375 (O_3375,N_29125,N_28878);
or UO_3376 (O_3376,N_29393,N_29079);
nand UO_3377 (O_3377,N_29342,N_29465);
nor UO_3378 (O_3378,N_29003,N_28769);
or UO_3379 (O_3379,N_29212,N_29792);
and UO_3380 (O_3380,N_29725,N_28611);
or UO_3381 (O_3381,N_29048,N_29285);
nor UO_3382 (O_3382,N_28790,N_28786);
and UO_3383 (O_3383,N_29486,N_28533);
and UO_3384 (O_3384,N_29754,N_28504);
nor UO_3385 (O_3385,N_29868,N_29259);
and UO_3386 (O_3386,N_29386,N_29980);
and UO_3387 (O_3387,N_29476,N_28591);
xnor UO_3388 (O_3388,N_28702,N_29051);
and UO_3389 (O_3389,N_29676,N_29006);
or UO_3390 (O_3390,N_29573,N_29960);
nor UO_3391 (O_3391,N_29248,N_29017);
or UO_3392 (O_3392,N_28815,N_28899);
nor UO_3393 (O_3393,N_29523,N_28539);
or UO_3394 (O_3394,N_29581,N_29919);
xor UO_3395 (O_3395,N_29975,N_29011);
xnor UO_3396 (O_3396,N_29143,N_29130);
and UO_3397 (O_3397,N_29251,N_28773);
nand UO_3398 (O_3398,N_29977,N_29890);
xor UO_3399 (O_3399,N_28897,N_28563);
nand UO_3400 (O_3400,N_29824,N_28673);
or UO_3401 (O_3401,N_29708,N_29209);
nor UO_3402 (O_3402,N_29297,N_29844);
xor UO_3403 (O_3403,N_28704,N_29888);
xnor UO_3404 (O_3404,N_29770,N_28823);
nand UO_3405 (O_3405,N_29035,N_29577);
xnor UO_3406 (O_3406,N_29474,N_29339);
or UO_3407 (O_3407,N_28687,N_29885);
or UO_3408 (O_3408,N_29168,N_29392);
nand UO_3409 (O_3409,N_29653,N_29618);
xor UO_3410 (O_3410,N_29922,N_29686);
or UO_3411 (O_3411,N_28712,N_29911);
or UO_3412 (O_3412,N_29262,N_28752);
nand UO_3413 (O_3413,N_29289,N_29458);
xnor UO_3414 (O_3414,N_29988,N_29409);
or UO_3415 (O_3415,N_28553,N_28833);
nand UO_3416 (O_3416,N_29660,N_29232);
nor UO_3417 (O_3417,N_29831,N_28513);
nand UO_3418 (O_3418,N_29602,N_29473);
or UO_3419 (O_3419,N_29640,N_28864);
nand UO_3420 (O_3420,N_29023,N_29028);
or UO_3421 (O_3421,N_29197,N_28836);
xnor UO_3422 (O_3422,N_29002,N_28518);
and UO_3423 (O_3423,N_29536,N_29639);
nor UO_3424 (O_3424,N_29652,N_29742);
nor UO_3425 (O_3425,N_29295,N_29162);
and UO_3426 (O_3426,N_29450,N_29100);
nand UO_3427 (O_3427,N_28722,N_29517);
and UO_3428 (O_3428,N_28647,N_29399);
nand UO_3429 (O_3429,N_29805,N_28787);
xor UO_3430 (O_3430,N_29902,N_28737);
or UO_3431 (O_3431,N_29454,N_29248);
and UO_3432 (O_3432,N_29556,N_29142);
nor UO_3433 (O_3433,N_29608,N_29968);
or UO_3434 (O_3434,N_29962,N_29619);
nor UO_3435 (O_3435,N_28505,N_29023);
nor UO_3436 (O_3436,N_29104,N_29357);
xnor UO_3437 (O_3437,N_29214,N_29014);
or UO_3438 (O_3438,N_29381,N_28875);
nand UO_3439 (O_3439,N_29429,N_29780);
xor UO_3440 (O_3440,N_28714,N_29623);
and UO_3441 (O_3441,N_29184,N_29954);
nand UO_3442 (O_3442,N_29125,N_28576);
nor UO_3443 (O_3443,N_28634,N_29092);
and UO_3444 (O_3444,N_29827,N_29295);
xor UO_3445 (O_3445,N_29529,N_29498);
nor UO_3446 (O_3446,N_29337,N_29834);
nand UO_3447 (O_3447,N_29939,N_29367);
or UO_3448 (O_3448,N_29280,N_29771);
and UO_3449 (O_3449,N_28672,N_29462);
xor UO_3450 (O_3450,N_28867,N_29484);
and UO_3451 (O_3451,N_29184,N_28638);
nand UO_3452 (O_3452,N_28889,N_29367);
nor UO_3453 (O_3453,N_28967,N_29890);
xor UO_3454 (O_3454,N_28748,N_28950);
xnor UO_3455 (O_3455,N_29354,N_29621);
or UO_3456 (O_3456,N_28736,N_28603);
or UO_3457 (O_3457,N_29227,N_28977);
nand UO_3458 (O_3458,N_29187,N_29259);
and UO_3459 (O_3459,N_28889,N_29576);
and UO_3460 (O_3460,N_29044,N_29238);
nand UO_3461 (O_3461,N_29088,N_28500);
or UO_3462 (O_3462,N_28880,N_28820);
nor UO_3463 (O_3463,N_28804,N_28939);
nor UO_3464 (O_3464,N_29299,N_28740);
or UO_3465 (O_3465,N_29151,N_29748);
and UO_3466 (O_3466,N_29938,N_29007);
or UO_3467 (O_3467,N_29718,N_29625);
nor UO_3468 (O_3468,N_29226,N_29490);
and UO_3469 (O_3469,N_29985,N_29798);
or UO_3470 (O_3470,N_28829,N_28911);
nor UO_3471 (O_3471,N_29610,N_28643);
or UO_3472 (O_3472,N_29655,N_29154);
xnor UO_3473 (O_3473,N_28526,N_28912);
or UO_3474 (O_3474,N_28731,N_28700);
or UO_3475 (O_3475,N_29318,N_29486);
or UO_3476 (O_3476,N_28789,N_29771);
or UO_3477 (O_3477,N_29203,N_29168);
nand UO_3478 (O_3478,N_29555,N_28661);
xnor UO_3479 (O_3479,N_29773,N_29442);
and UO_3480 (O_3480,N_29380,N_29736);
xnor UO_3481 (O_3481,N_28741,N_29908);
nor UO_3482 (O_3482,N_29555,N_28933);
or UO_3483 (O_3483,N_28962,N_28792);
xor UO_3484 (O_3484,N_29174,N_29594);
nand UO_3485 (O_3485,N_29862,N_29528);
or UO_3486 (O_3486,N_29964,N_29937);
or UO_3487 (O_3487,N_29412,N_28725);
and UO_3488 (O_3488,N_29912,N_29449);
or UO_3489 (O_3489,N_29702,N_29229);
nand UO_3490 (O_3490,N_29099,N_29158);
nor UO_3491 (O_3491,N_29925,N_29996);
nand UO_3492 (O_3492,N_28591,N_29781);
xor UO_3493 (O_3493,N_28744,N_29751);
xor UO_3494 (O_3494,N_28836,N_29421);
xor UO_3495 (O_3495,N_29608,N_29392);
or UO_3496 (O_3496,N_28711,N_29167);
xor UO_3497 (O_3497,N_29377,N_29478);
nor UO_3498 (O_3498,N_29832,N_28502);
nor UO_3499 (O_3499,N_28864,N_28768);
endmodule