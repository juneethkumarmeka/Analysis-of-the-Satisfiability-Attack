module basic_750_5000_1000_25_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
or U0 (N_0,In_39,In_51);
nor U1 (N_1,In_613,In_479);
nor U2 (N_2,In_300,In_387);
or U3 (N_3,In_656,In_440);
xor U4 (N_4,In_181,In_580);
and U5 (N_5,In_225,In_735);
and U6 (N_6,In_354,In_342);
xnor U7 (N_7,In_22,In_411);
and U8 (N_8,In_66,In_657);
nor U9 (N_9,In_89,In_467);
nand U10 (N_10,In_168,In_159);
xnor U11 (N_11,In_235,In_299);
or U12 (N_12,In_289,In_645);
nand U13 (N_13,In_267,In_612);
nor U14 (N_14,In_582,In_686);
and U15 (N_15,In_359,In_595);
xor U16 (N_16,In_394,In_196);
xnor U17 (N_17,In_527,In_661);
nand U18 (N_18,In_130,In_632);
xor U19 (N_19,In_373,In_55);
xnor U20 (N_20,In_386,In_471);
nand U21 (N_21,In_677,In_81);
xnor U22 (N_22,In_207,In_624);
xnor U23 (N_23,In_572,In_364);
or U24 (N_24,In_2,In_366);
and U25 (N_25,In_586,In_301);
nor U26 (N_26,In_112,In_244);
nand U27 (N_27,In_665,In_331);
nor U28 (N_28,In_108,In_74);
xor U29 (N_29,In_293,In_230);
xor U30 (N_30,In_675,In_737);
and U31 (N_31,In_34,In_623);
xor U32 (N_32,In_5,In_454);
nand U33 (N_33,In_187,In_369);
and U34 (N_34,In_689,In_337);
nand U35 (N_35,In_578,In_120);
xor U36 (N_36,In_738,In_189);
nand U37 (N_37,In_642,In_643);
and U38 (N_38,In_637,In_336);
nor U39 (N_39,In_118,In_156);
or U40 (N_40,In_177,In_715);
or U41 (N_41,In_102,In_93);
nand U42 (N_42,In_104,In_127);
or U43 (N_43,In_721,In_88);
xnor U44 (N_44,In_135,In_536);
nor U45 (N_45,In_636,In_325);
xnor U46 (N_46,In_353,In_182);
xor U47 (N_47,In_310,In_631);
or U48 (N_48,In_234,In_24);
nand U49 (N_49,In_427,In_634);
nor U50 (N_50,In_397,In_483);
nand U51 (N_51,In_286,In_101);
nor U52 (N_52,In_734,In_589);
nor U53 (N_53,In_407,In_747);
and U54 (N_54,In_72,In_152);
and U55 (N_55,In_423,In_206);
nor U56 (N_56,In_324,In_662);
nand U57 (N_57,In_518,In_224);
nor U58 (N_58,In_746,In_257);
and U59 (N_59,In_504,In_131);
nor U60 (N_60,In_659,In_258);
xor U61 (N_61,In_450,In_14);
and U62 (N_62,In_683,In_568);
xnor U63 (N_63,In_283,In_320);
xor U64 (N_64,In_98,In_158);
xnor U65 (N_65,In_178,In_604);
nor U66 (N_66,In_113,In_501);
or U67 (N_67,In_462,In_195);
and U68 (N_68,In_626,In_87);
or U69 (N_69,In_71,In_555);
xor U70 (N_70,In_546,In_363);
xnor U71 (N_71,In_539,In_512);
nand U72 (N_72,In_139,In_345);
or U73 (N_73,In_273,In_498);
and U74 (N_74,In_640,In_576);
or U75 (N_75,In_429,In_264);
and U76 (N_76,In_202,In_605);
or U77 (N_77,In_648,In_185);
and U78 (N_78,In_415,In_153);
or U79 (N_79,In_263,In_560);
or U80 (N_80,In_193,In_302);
and U81 (N_81,In_630,In_327);
nand U82 (N_82,In_489,In_682);
nand U83 (N_83,In_166,In_692);
and U84 (N_84,In_426,In_729);
nor U85 (N_85,In_314,In_708);
nor U86 (N_86,In_585,In_36);
and U87 (N_87,In_664,In_140);
xnor U88 (N_88,In_651,In_649);
nand U89 (N_89,In_164,In_250);
nand U90 (N_90,In_94,In_162);
nor U91 (N_91,In_514,In_10);
and U92 (N_92,In_468,In_491);
or U93 (N_93,In_610,In_639);
xnor U94 (N_94,In_124,In_487);
nor U95 (N_95,In_368,In_295);
and U96 (N_96,In_376,In_571);
or U97 (N_97,In_396,In_303);
nand U98 (N_98,In_259,In_236);
or U99 (N_99,In_183,In_305);
or U100 (N_100,In_97,In_384);
or U101 (N_101,In_609,In_70);
or U102 (N_102,In_69,In_211);
nor U103 (N_103,In_524,In_277);
nand U104 (N_104,In_220,In_41);
or U105 (N_105,In_528,In_134);
nand U106 (N_106,In_272,In_451);
nand U107 (N_107,In_247,In_122);
nor U108 (N_108,In_511,In_591);
nand U109 (N_109,In_281,In_237);
xor U110 (N_110,In_219,In_175);
nand U111 (N_111,In_35,In_606);
nor U112 (N_112,In_575,In_274);
nand U113 (N_113,In_222,In_92);
nor U114 (N_114,In_298,In_275);
and U115 (N_115,In_502,In_532);
or U116 (N_116,In_684,In_388);
xor U117 (N_117,In_76,In_495);
nand U118 (N_118,In_562,In_420);
nand U119 (N_119,In_367,In_21);
and U120 (N_120,In_456,In_566);
or U121 (N_121,In_461,In_103);
and U122 (N_122,In_343,In_748);
nand U123 (N_123,In_592,In_442);
nor U124 (N_124,In_297,In_121);
xor U125 (N_125,In_599,In_111);
xor U126 (N_126,In_728,In_523);
nand U127 (N_127,In_490,In_16);
nor U128 (N_128,In_169,In_745);
xor U129 (N_129,In_284,In_484);
and U130 (N_130,In_198,In_658);
or U131 (N_131,In_702,In_319);
and U132 (N_132,In_554,In_339);
nor U133 (N_133,In_64,In_254);
nor U134 (N_134,In_570,In_433);
xnor U135 (N_135,In_688,In_401);
xor U136 (N_136,In_186,In_614);
and U137 (N_137,In_438,In_465);
and U138 (N_138,In_463,In_707);
and U139 (N_139,In_378,In_425);
nor U140 (N_140,In_223,In_507);
xor U141 (N_141,In_232,In_603);
or U142 (N_142,In_650,In_154);
xnor U143 (N_143,In_553,In_63);
nand U144 (N_144,In_44,In_443);
or U145 (N_145,In_672,In_133);
and U146 (N_146,In_473,In_448);
xor U147 (N_147,In_598,In_667);
nor U148 (N_148,In_749,In_204);
nand U149 (N_149,In_482,In_360);
and U150 (N_150,In_216,In_80);
nand U151 (N_151,In_23,In_341);
and U152 (N_152,In_711,In_252);
xor U153 (N_153,In_9,In_392);
xnor U154 (N_154,In_290,In_556);
and U155 (N_155,In_654,In_79);
xor U156 (N_156,In_530,In_497);
and U157 (N_157,In_478,In_73);
nor U158 (N_158,In_188,In_285);
nor U159 (N_159,In_531,In_418);
or U160 (N_160,In_57,In_709);
xor U161 (N_161,In_557,In_26);
xnor U162 (N_162,In_633,In_240);
and U163 (N_163,In_375,In_516);
nand U164 (N_164,In_307,In_99);
nand U165 (N_165,In_48,In_311);
and U166 (N_166,In_458,In_344);
nor U167 (N_167,In_646,In_262);
or U168 (N_168,In_493,In_62);
xnor U169 (N_169,In_100,In_242);
and U170 (N_170,In_663,In_340);
xor U171 (N_171,In_318,In_710);
nor U172 (N_172,In_357,In_733);
nand U173 (N_173,In_409,In_165);
xnor U174 (N_174,In_544,In_243);
nand U175 (N_175,In_472,In_45);
and U176 (N_176,In_282,In_726);
nand U177 (N_177,In_541,In_453);
nor U178 (N_178,In_404,In_671);
nor U179 (N_179,In_703,In_308);
nor U180 (N_180,In_736,In_226);
xor U181 (N_181,In_410,In_65);
and U182 (N_182,In_573,In_229);
nor U183 (N_183,In_115,In_291);
and U184 (N_184,In_678,In_540);
or U185 (N_185,In_545,In_374);
and U186 (N_186,In_408,In_137);
xor U187 (N_187,In_25,In_447);
nor U188 (N_188,In_668,In_417);
and U189 (N_189,In_190,In_33);
and U190 (N_190,In_402,In_61);
nand U191 (N_191,In_564,In_1);
nor U192 (N_192,In_525,In_727);
xor U193 (N_193,In_329,In_379);
xor U194 (N_194,In_53,In_246);
xnor U195 (N_195,In_414,In_322);
nand U196 (N_196,In_171,In_563);
nand U197 (N_197,In_611,In_647);
nand U198 (N_198,In_519,In_693);
xor U199 (N_199,In_132,In_348);
xnor U200 (N_200,N_143,N_9);
nand U201 (N_201,In_77,N_182);
and U202 (N_202,In_338,In_559);
nor U203 (N_203,N_149,N_129);
and U204 (N_204,In_205,In_551);
nor U205 (N_205,In_255,N_39);
nand U206 (N_206,N_37,In_160);
nand U207 (N_207,In_15,In_607);
or U208 (N_208,In_385,In_296);
or U209 (N_209,In_270,In_136);
nand U210 (N_210,In_214,N_61);
xor U211 (N_211,N_191,In_174);
and U212 (N_212,In_597,In_248);
xor U213 (N_213,N_180,In_644);
nand U214 (N_214,N_159,In_577);
xor U215 (N_215,N_19,N_36);
or U216 (N_216,In_722,In_146);
nand U217 (N_217,N_87,In_29);
nor U218 (N_218,In_54,In_155);
and U219 (N_219,In_123,In_352);
xnor U220 (N_220,N_77,N_68);
xor U221 (N_221,N_130,In_725);
or U222 (N_222,In_355,In_260);
nor U223 (N_223,N_32,In_655);
and U224 (N_224,N_13,In_506);
xor U225 (N_225,N_83,In_8);
and U226 (N_226,In_616,In_526);
nand U227 (N_227,N_128,N_80);
and U228 (N_228,N_1,In_625);
or U229 (N_229,In_587,In_362);
and U230 (N_230,N_66,In_43);
nand U231 (N_231,In_201,In_334);
xnor U232 (N_232,In_278,N_194);
and U233 (N_233,In_517,In_670);
nand U234 (N_234,In_543,In_622);
or U235 (N_235,N_85,In_717);
xnor U236 (N_236,In_380,In_86);
xor U237 (N_237,In_27,In_91);
and U238 (N_238,In_485,In_513);
xnor U239 (N_239,N_16,N_124);
nor U240 (N_240,In_125,In_312);
xor U241 (N_241,N_98,N_99);
or U242 (N_242,In_534,In_569);
xnor U243 (N_243,In_617,N_151);
nand U244 (N_244,N_100,In_515);
xnor U245 (N_245,In_107,In_50);
xor U246 (N_246,In_698,N_23);
nand U247 (N_247,N_4,N_119);
nor U248 (N_248,N_164,In_391);
and U249 (N_249,N_190,In_480);
nor U250 (N_250,In_475,In_313);
nand U251 (N_251,In_95,N_29);
or U252 (N_252,In_184,In_31);
nand U253 (N_253,In_691,N_81);
and U254 (N_254,N_75,In_430);
xor U255 (N_255,In_567,In_12);
nor U256 (N_256,N_35,In_681);
xor U257 (N_257,N_101,In_78);
or U258 (N_258,In_84,In_161);
xnor U259 (N_259,In_720,In_744);
or U260 (N_260,In_588,N_7);
nor U261 (N_261,N_148,N_156);
nor U262 (N_262,N_42,N_186);
and U263 (N_263,In_83,In_492);
nand U264 (N_264,N_86,In_280);
or U265 (N_265,N_8,N_104);
or U266 (N_266,N_34,N_97);
or U267 (N_267,In_694,In_434);
and U268 (N_268,In_537,N_125);
or U269 (N_269,In_444,In_581);
xnor U270 (N_270,In_416,In_138);
nor U271 (N_271,In_615,N_198);
nor U272 (N_272,In_696,In_256);
xor U273 (N_273,N_135,N_132);
nor U274 (N_274,N_90,In_227);
nand U275 (N_275,N_31,In_317);
nand U276 (N_276,In_446,N_138);
nand U277 (N_277,N_92,In_105);
xor U278 (N_278,In_574,N_115);
nor U279 (N_279,In_157,N_78);
nand U280 (N_280,N_175,In_584);
nand U281 (N_281,N_172,N_154);
nor U282 (N_282,In_333,In_436);
nor U283 (N_283,In_538,N_165);
nand U284 (N_284,In_629,In_316);
xor U285 (N_285,In_549,In_590);
or U286 (N_286,N_88,N_163);
or U287 (N_287,In_172,N_93);
nor U288 (N_288,N_57,In_579);
and U289 (N_289,In_180,In_740);
nor U290 (N_290,N_157,In_212);
and U291 (N_291,N_91,In_253);
xor U292 (N_292,N_54,In_608);
nand U293 (N_293,N_111,N_176);
xnor U294 (N_294,N_178,In_266);
xnor U295 (N_295,In_638,N_199);
xnor U296 (N_296,In_142,In_129);
xnor U297 (N_297,N_142,N_47);
or U298 (N_298,In_390,N_64);
nand U299 (N_299,N_74,In_149);
xnor U300 (N_300,In_508,In_346);
or U301 (N_301,N_105,N_137);
nor U302 (N_302,In_221,In_405);
nand U303 (N_303,In_494,N_118);
nand U304 (N_304,N_3,N_177);
or U305 (N_305,In_412,In_238);
xnor U306 (N_306,N_43,In_0);
and U307 (N_307,N_179,N_63);
nand U308 (N_308,N_50,In_690);
nand U309 (N_309,In_49,In_268);
nand U310 (N_310,In_419,In_231);
xnor U311 (N_311,In_383,N_51);
and U312 (N_312,In_32,In_18);
xor U313 (N_313,In_449,In_676);
nand U314 (N_314,N_123,In_209);
nor U315 (N_315,In_469,N_24);
or U316 (N_316,In_697,N_45);
and U317 (N_317,In_38,In_561);
or U318 (N_318,N_40,N_11);
nor U319 (N_319,In_424,N_120);
nand U320 (N_320,In_326,In_403);
nor U321 (N_321,N_65,N_62);
nand U322 (N_322,In_474,N_153);
or U323 (N_323,N_5,N_136);
nor U324 (N_324,In_110,In_347);
and U325 (N_325,In_685,In_128);
and U326 (N_326,In_712,In_718);
nor U327 (N_327,In_328,In_673);
or U328 (N_328,In_371,In_109);
nor U329 (N_329,In_635,In_47);
xor U330 (N_330,In_558,N_6);
xnor U331 (N_331,N_181,N_79);
or U332 (N_332,In_428,In_547);
and U333 (N_333,N_113,In_28);
nand U334 (N_334,In_56,In_723);
xor U335 (N_335,In_421,N_107);
xor U336 (N_336,In_509,In_332);
and U337 (N_337,In_321,N_150);
or U338 (N_338,In_208,In_413);
and U339 (N_339,N_158,In_217);
nor U340 (N_340,In_309,In_276);
or U341 (N_341,In_170,In_67);
nor U342 (N_342,In_452,N_127);
and U343 (N_343,In_601,N_20);
nand U344 (N_344,N_140,In_239);
nor U345 (N_345,In_457,In_372);
or U346 (N_346,In_533,In_304);
or U347 (N_347,In_116,In_481);
nor U348 (N_348,In_4,In_143);
and U349 (N_349,In_288,N_144);
nor U350 (N_350,In_739,N_49);
or U351 (N_351,In_151,In_695);
or U352 (N_352,In_147,In_521);
and U353 (N_353,In_741,In_594);
xor U354 (N_354,In_618,In_389);
nor U355 (N_355,N_170,N_12);
nand U356 (N_356,In_701,In_652);
nor U357 (N_357,In_395,In_215);
or U358 (N_358,N_121,In_7);
and U359 (N_359,In_213,In_641);
nor U360 (N_360,In_510,In_30);
and U361 (N_361,N_134,In_435);
nor U362 (N_362,N_46,N_72);
xor U363 (N_363,In_68,In_176);
and U364 (N_364,N_84,In_400);
nor U365 (N_365,In_716,In_505);
and U366 (N_366,N_59,In_3);
nor U367 (N_367,N_196,N_44);
xor U368 (N_368,In_653,N_168);
xnor U369 (N_369,N_116,N_162);
nor U370 (N_370,N_94,N_112);
nor U371 (N_371,N_21,In_459);
nand U372 (N_372,In_439,N_58);
xnor U373 (N_373,N_0,In_292);
xor U374 (N_374,In_552,In_705);
nand U375 (N_375,In_370,In_382);
or U376 (N_376,In_218,In_503);
nand U377 (N_377,N_52,N_155);
or U378 (N_378,In_596,In_315);
nor U379 (N_379,In_251,N_145);
or U380 (N_380,In_550,In_265);
xor U381 (N_381,In_713,In_548);
xor U382 (N_382,In_687,N_14);
xnor U383 (N_383,N_139,In_680);
nand U384 (N_384,N_167,In_279);
nand U385 (N_385,In_361,In_488);
and U386 (N_386,In_117,N_187);
nor U387 (N_387,N_95,In_496);
xor U388 (N_388,In_730,In_714);
and U389 (N_389,N_141,In_706);
or U390 (N_390,In_200,In_666);
nor U391 (N_391,In_59,In_58);
xnor U392 (N_392,In_704,In_85);
xnor U393 (N_393,N_25,N_161);
nand U394 (N_394,N_192,N_33);
nand U395 (N_395,N_110,N_55);
nor U396 (N_396,N_27,In_583);
nand U397 (N_397,In_294,In_60);
and U398 (N_398,In_192,In_306);
nand U399 (N_399,In_627,N_106);
xnor U400 (N_400,N_285,N_269);
or U401 (N_401,In_106,N_232);
or U402 (N_402,N_336,N_56);
or U403 (N_403,N_357,In_406);
and U404 (N_404,N_73,N_207);
xor U405 (N_405,N_389,N_274);
xnor U406 (N_406,In_529,N_321);
and U407 (N_407,In_441,N_327);
and U408 (N_408,In_228,N_287);
and U409 (N_409,N_331,N_386);
nand U410 (N_410,In_179,N_275);
xnor U411 (N_411,In_731,In_323);
nor U412 (N_412,N_218,N_356);
xnor U413 (N_413,N_394,N_302);
nand U414 (N_414,N_249,In_620);
xor U415 (N_415,N_184,N_365);
and U416 (N_416,In_399,N_307);
or U417 (N_417,N_234,In_75);
and U418 (N_418,In_40,N_208);
nand U419 (N_419,In_37,N_313);
xnor U420 (N_420,N_322,In_13);
or U421 (N_421,N_265,N_343);
xor U422 (N_422,In_351,N_366);
xnor U423 (N_423,N_303,N_205);
nand U424 (N_424,N_335,N_38);
nand U425 (N_425,N_383,N_297);
and U426 (N_426,N_26,N_253);
nand U427 (N_427,N_237,In_350);
nor U428 (N_428,N_195,N_290);
nand U429 (N_429,N_244,N_223);
xnor U430 (N_430,N_255,N_277);
xor U431 (N_431,In_669,N_131);
nand U432 (N_432,N_377,N_18);
or U433 (N_433,N_71,N_264);
and U434 (N_434,N_340,In_42);
or U435 (N_435,In_144,In_19);
or U436 (N_436,N_375,In_287);
xor U437 (N_437,N_318,N_283);
and U438 (N_438,In_520,In_621);
or U439 (N_439,N_82,N_399);
xnor U440 (N_440,N_299,N_296);
and U441 (N_441,N_384,N_222);
or U442 (N_442,N_319,N_270);
nor U443 (N_443,In_163,N_22);
or U444 (N_444,N_330,N_203);
xor U445 (N_445,N_267,N_373);
and U446 (N_446,N_53,N_272);
nand U447 (N_447,In_422,N_273);
nor U448 (N_448,N_368,N_263);
nand U449 (N_449,In_365,In_199);
nor U450 (N_450,In_119,N_395);
nor U451 (N_451,N_126,N_388);
or U452 (N_452,N_108,N_183);
nor U453 (N_453,N_189,N_236);
and U454 (N_454,In_173,In_464);
and U455 (N_455,In_126,N_268);
xnor U456 (N_456,N_28,In_46);
nand U457 (N_457,In_167,N_60);
nand U458 (N_458,In_679,N_213);
or U459 (N_459,In_114,N_2);
xnor U460 (N_460,N_235,N_344);
or U461 (N_461,N_256,N_233);
and U462 (N_462,N_133,N_245);
and U463 (N_463,N_292,In_245);
and U464 (N_464,N_355,N_333);
nand U465 (N_465,In_271,N_240);
or U466 (N_466,N_298,N_238);
or U467 (N_467,In_6,In_460);
nor U468 (N_468,N_257,N_122);
or U469 (N_469,N_193,N_341);
and U470 (N_470,N_239,N_315);
or U471 (N_471,N_241,N_173);
and U472 (N_472,In_699,N_361);
nor U473 (N_473,N_70,N_109);
and U474 (N_474,In_330,N_246);
or U475 (N_475,N_247,N_204);
nor U476 (N_476,N_248,In_486);
or U477 (N_477,N_306,N_278);
or U478 (N_478,In_477,N_300);
or U479 (N_479,N_374,N_291);
and U480 (N_480,N_259,N_15);
nor U481 (N_481,N_230,N_358);
or U482 (N_482,In_600,N_174);
xor U483 (N_483,N_202,N_390);
or U484 (N_484,In_96,In_393);
nor U485 (N_485,N_220,N_188);
and U486 (N_486,N_169,N_201);
nand U487 (N_487,N_279,N_258);
xor U488 (N_488,In_732,N_387);
xnor U489 (N_489,In_377,N_301);
or U490 (N_490,N_229,In_565);
and U491 (N_491,N_282,N_362);
xor U492 (N_492,In_674,N_295);
nor U493 (N_493,N_242,In_535);
xnor U494 (N_494,In_145,N_206);
xnor U495 (N_495,In_269,N_304);
xor U496 (N_496,N_117,N_380);
and U497 (N_497,N_243,N_324);
xor U498 (N_498,N_379,N_227);
and U499 (N_499,N_76,N_312);
nand U500 (N_500,In_602,N_41);
nand U501 (N_501,N_211,N_381);
or U502 (N_502,N_147,In_52);
or U503 (N_503,N_171,In_148);
nand U504 (N_504,In_358,N_337);
nor U505 (N_505,In_141,In_724);
or U506 (N_506,In_700,N_328);
xor U507 (N_507,In_660,In_466);
nor U508 (N_508,N_281,N_360);
or U509 (N_509,N_215,In_17);
nor U510 (N_510,In_261,In_194);
or U511 (N_511,N_276,In_593);
nor U512 (N_512,N_288,N_316);
or U513 (N_513,In_432,N_294);
and U514 (N_514,N_216,N_228);
or U515 (N_515,In_455,N_103);
nand U516 (N_516,N_293,N_250);
nor U517 (N_517,N_221,N_369);
or U518 (N_518,N_345,N_309);
and U519 (N_519,N_376,In_437);
nand U520 (N_520,N_351,N_354);
and U521 (N_521,In_191,N_348);
xnor U522 (N_522,N_363,N_310);
and U523 (N_523,N_160,N_210);
xor U524 (N_524,N_329,N_308);
nand U525 (N_525,N_48,In_249);
nand U526 (N_526,In_82,N_209);
and U527 (N_527,In_431,N_334);
or U528 (N_528,N_152,N_305);
and U529 (N_529,N_260,N_67);
xor U530 (N_530,N_10,N_385);
and U531 (N_531,N_367,In_499);
and U532 (N_532,In_241,N_350);
nand U533 (N_533,N_317,N_185);
or U534 (N_534,N_96,N_325);
xnor U535 (N_535,In_210,In_11);
nor U536 (N_536,N_396,N_371);
nor U537 (N_537,N_364,N_114);
nor U538 (N_538,N_346,N_197);
xor U539 (N_539,In_500,N_224);
or U540 (N_540,In_349,N_266);
nand U541 (N_541,N_30,N_326);
or U542 (N_542,N_212,In_90);
nand U543 (N_543,In_150,In_445);
nor U544 (N_544,In_203,N_217);
nor U545 (N_545,N_146,In_476);
nor U546 (N_546,N_352,N_231);
and U547 (N_547,N_214,N_393);
xnor U548 (N_548,N_397,N_102);
nor U549 (N_549,N_261,In_719);
nor U550 (N_550,N_17,N_280);
nor U551 (N_551,N_353,In_743);
xor U552 (N_552,In_522,N_254);
nor U553 (N_553,N_200,N_347);
nand U554 (N_554,In_628,In_335);
and U555 (N_555,In_20,In_197);
nand U556 (N_556,N_320,N_225);
xnor U557 (N_557,In_381,N_398);
xnor U558 (N_558,N_219,N_349);
nor U559 (N_559,In_470,N_311);
xor U560 (N_560,N_392,N_286);
or U561 (N_561,In_619,N_370);
nor U562 (N_562,N_372,N_251);
xnor U563 (N_563,N_262,In_356);
or U564 (N_564,N_359,N_166);
and U565 (N_565,N_69,N_271);
xnor U566 (N_566,N_342,N_391);
xnor U567 (N_567,N_89,In_233);
nor U568 (N_568,N_314,N_226);
xnor U569 (N_569,N_338,N_378);
nand U570 (N_570,In_542,N_382);
nor U571 (N_571,In_398,In_742);
and U572 (N_572,N_339,N_252);
or U573 (N_573,N_332,N_323);
nor U574 (N_574,N_289,N_284);
and U575 (N_575,N_292,N_152);
or U576 (N_576,N_342,N_275);
nand U577 (N_577,N_369,N_242);
and U578 (N_578,N_146,N_231);
nand U579 (N_579,N_213,In_228);
nor U580 (N_580,N_236,N_221);
nand U581 (N_581,N_216,In_20);
or U582 (N_582,N_317,N_221);
nor U583 (N_583,In_476,N_251);
nand U584 (N_584,N_246,N_22);
or U585 (N_585,N_362,N_256);
nor U586 (N_586,In_441,In_245);
nand U587 (N_587,N_381,N_320);
or U588 (N_588,In_700,N_373);
xnor U589 (N_589,N_225,N_355);
and U590 (N_590,N_38,In_432);
and U591 (N_591,N_236,N_358);
nand U592 (N_592,In_399,N_26);
nand U593 (N_593,N_278,N_332);
or U594 (N_594,In_191,N_344);
xnor U595 (N_595,N_341,N_305);
xnor U596 (N_596,N_152,N_224);
and U597 (N_597,N_380,N_241);
and U598 (N_598,N_249,N_260);
nor U599 (N_599,In_323,In_179);
and U600 (N_600,N_402,N_404);
and U601 (N_601,N_492,N_517);
nor U602 (N_602,N_452,N_465);
or U603 (N_603,N_496,N_558);
xor U604 (N_604,N_549,N_563);
nor U605 (N_605,N_444,N_420);
xnor U606 (N_606,N_490,N_596);
nand U607 (N_607,N_488,N_590);
nor U608 (N_608,N_501,N_483);
nor U609 (N_609,N_526,N_578);
xnor U610 (N_610,N_564,N_557);
or U611 (N_611,N_500,N_507);
and U612 (N_612,N_512,N_516);
and U613 (N_613,N_560,N_595);
and U614 (N_614,N_427,N_550);
or U615 (N_615,N_541,N_570);
or U616 (N_616,N_469,N_450);
xnor U617 (N_617,N_518,N_553);
and U618 (N_618,N_588,N_457);
nand U619 (N_619,N_476,N_555);
nand U620 (N_620,N_439,N_508);
or U621 (N_621,N_477,N_568);
and U622 (N_622,N_432,N_414);
nor U623 (N_623,N_587,N_535);
or U624 (N_624,N_413,N_544);
or U625 (N_625,N_429,N_593);
nor U626 (N_626,N_505,N_581);
xnor U627 (N_627,N_461,N_425);
nand U628 (N_628,N_575,N_491);
or U629 (N_629,N_407,N_435);
xor U630 (N_630,N_521,N_442);
nand U631 (N_631,N_585,N_424);
xor U632 (N_632,N_576,N_479);
or U633 (N_633,N_511,N_470);
or U634 (N_634,N_494,N_498);
xnor U635 (N_635,N_583,N_484);
or U636 (N_636,N_542,N_466);
and U637 (N_637,N_562,N_421);
and U638 (N_638,N_504,N_572);
or U639 (N_639,N_403,N_410);
nor U640 (N_640,N_559,N_536);
or U641 (N_641,N_474,N_592);
nand U642 (N_642,N_497,N_556);
or U643 (N_643,N_565,N_577);
nor U644 (N_644,N_486,N_487);
nand U645 (N_645,N_561,N_408);
nor U646 (N_646,N_417,N_552);
nand U647 (N_647,N_456,N_545);
nand U648 (N_648,N_419,N_423);
nor U649 (N_649,N_449,N_416);
xor U650 (N_650,N_597,N_400);
nor U651 (N_651,N_509,N_527);
nand U652 (N_652,N_589,N_510);
or U653 (N_653,N_548,N_471);
or U654 (N_654,N_514,N_438);
or U655 (N_655,N_431,N_415);
xor U656 (N_656,N_513,N_478);
nor U657 (N_657,N_537,N_454);
and U658 (N_658,N_547,N_463);
or U659 (N_659,N_554,N_401);
nor U660 (N_660,N_418,N_571);
and U661 (N_661,N_443,N_428);
nand U662 (N_662,N_499,N_502);
or U663 (N_663,N_566,N_495);
nand U664 (N_664,N_412,N_409);
and U665 (N_665,N_472,N_598);
nor U666 (N_666,N_522,N_532);
nor U667 (N_667,N_586,N_426);
and U668 (N_668,N_519,N_460);
nand U669 (N_669,N_482,N_434);
or U670 (N_670,N_475,N_473);
nand U671 (N_671,N_567,N_533);
or U672 (N_672,N_515,N_448);
nor U673 (N_673,N_437,N_422);
and U674 (N_674,N_481,N_530);
and U675 (N_675,N_540,N_445);
xor U676 (N_676,N_430,N_546);
nor U677 (N_677,N_579,N_584);
nand U678 (N_678,N_433,N_447);
and U679 (N_679,N_520,N_485);
nand U680 (N_680,N_506,N_539);
and U681 (N_681,N_464,N_436);
or U682 (N_682,N_524,N_455);
and U683 (N_683,N_441,N_405);
nor U684 (N_684,N_458,N_582);
and U685 (N_685,N_440,N_580);
nor U686 (N_686,N_523,N_569);
nor U687 (N_687,N_574,N_406);
and U688 (N_688,N_573,N_538);
xor U689 (N_689,N_459,N_551);
nor U690 (N_690,N_468,N_489);
nand U691 (N_691,N_543,N_503);
nor U692 (N_692,N_528,N_462);
xnor U693 (N_693,N_467,N_594);
and U694 (N_694,N_534,N_599);
nor U695 (N_695,N_446,N_451);
nand U696 (N_696,N_480,N_411);
xnor U697 (N_697,N_531,N_453);
or U698 (N_698,N_493,N_591);
xor U699 (N_699,N_525,N_529);
nor U700 (N_700,N_529,N_555);
and U701 (N_701,N_503,N_544);
or U702 (N_702,N_552,N_509);
or U703 (N_703,N_572,N_401);
or U704 (N_704,N_481,N_576);
nand U705 (N_705,N_430,N_487);
nand U706 (N_706,N_595,N_538);
and U707 (N_707,N_531,N_467);
nand U708 (N_708,N_464,N_566);
and U709 (N_709,N_535,N_513);
and U710 (N_710,N_490,N_410);
and U711 (N_711,N_517,N_539);
nand U712 (N_712,N_515,N_558);
nor U713 (N_713,N_489,N_595);
nor U714 (N_714,N_525,N_573);
or U715 (N_715,N_435,N_420);
or U716 (N_716,N_489,N_549);
and U717 (N_717,N_441,N_478);
and U718 (N_718,N_559,N_455);
nand U719 (N_719,N_504,N_416);
nand U720 (N_720,N_598,N_596);
nor U721 (N_721,N_453,N_581);
or U722 (N_722,N_475,N_575);
nand U723 (N_723,N_583,N_571);
nor U724 (N_724,N_468,N_536);
and U725 (N_725,N_516,N_465);
nand U726 (N_726,N_515,N_574);
and U727 (N_727,N_429,N_561);
and U728 (N_728,N_579,N_453);
and U729 (N_729,N_402,N_539);
and U730 (N_730,N_459,N_401);
or U731 (N_731,N_479,N_419);
nor U732 (N_732,N_440,N_459);
and U733 (N_733,N_523,N_547);
or U734 (N_734,N_558,N_444);
nand U735 (N_735,N_418,N_578);
and U736 (N_736,N_554,N_455);
or U737 (N_737,N_581,N_510);
nand U738 (N_738,N_435,N_489);
or U739 (N_739,N_440,N_497);
xnor U740 (N_740,N_519,N_525);
nor U741 (N_741,N_497,N_402);
nand U742 (N_742,N_525,N_415);
nor U743 (N_743,N_453,N_451);
nand U744 (N_744,N_467,N_510);
nor U745 (N_745,N_510,N_410);
or U746 (N_746,N_597,N_572);
xor U747 (N_747,N_546,N_569);
nand U748 (N_748,N_556,N_469);
xnor U749 (N_749,N_524,N_440);
nand U750 (N_750,N_549,N_477);
or U751 (N_751,N_571,N_440);
nand U752 (N_752,N_573,N_586);
nor U753 (N_753,N_506,N_578);
nor U754 (N_754,N_417,N_550);
nand U755 (N_755,N_410,N_533);
or U756 (N_756,N_416,N_581);
and U757 (N_757,N_575,N_510);
or U758 (N_758,N_554,N_446);
and U759 (N_759,N_579,N_541);
nand U760 (N_760,N_431,N_490);
and U761 (N_761,N_401,N_439);
and U762 (N_762,N_472,N_564);
nand U763 (N_763,N_580,N_543);
or U764 (N_764,N_566,N_445);
nand U765 (N_765,N_495,N_475);
nor U766 (N_766,N_427,N_498);
and U767 (N_767,N_419,N_487);
xor U768 (N_768,N_467,N_522);
nor U769 (N_769,N_586,N_554);
xor U770 (N_770,N_491,N_589);
xnor U771 (N_771,N_532,N_573);
xnor U772 (N_772,N_419,N_410);
nor U773 (N_773,N_590,N_589);
or U774 (N_774,N_454,N_556);
or U775 (N_775,N_483,N_446);
and U776 (N_776,N_471,N_567);
xor U777 (N_777,N_443,N_595);
xnor U778 (N_778,N_443,N_447);
xnor U779 (N_779,N_435,N_563);
xor U780 (N_780,N_508,N_592);
nand U781 (N_781,N_472,N_477);
nor U782 (N_782,N_588,N_433);
xnor U783 (N_783,N_494,N_552);
nand U784 (N_784,N_538,N_491);
or U785 (N_785,N_458,N_585);
and U786 (N_786,N_406,N_529);
nor U787 (N_787,N_440,N_506);
or U788 (N_788,N_557,N_435);
xnor U789 (N_789,N_581,N_455);
or U790 (N_790,N_486,N_501);
nor U791 (N_791,N_596,N_577);
or U792 (N_792,N_464,N_486);
xnor U793 (N_793,N_579,N_527);
nand U794 (N_794,N_502,N_411);
nor U795 (N_795,N_550,N_436);
xnor U796 (N_796,N_433,N_514);
xnor U797 (N_797,N_417,N_547);
or U798 (N_798,N_431,N_481);
nand U799 (N_799,N_586,N_455);
nor U800 (N_800,N_668,N_721);
xnor U801 (N_801,N_726,N_622);
xor U802 (N_802,N_629,N_713);
xnor U803 (N_803,N_723,N_683);
nor U804 (N_804,N_787,N_605);
nor U805 (N_805,N_711,N_670);
nand U806 (N_806,N_748,N_732);
xnor U807 (N_807,N_740,N_798);
or U808 (N_808,N_655,N_776);
nor U809 (N_809,N_648,N_615);
xnor U810 (N_810,N_734,N_606);
xnor U811 (N_811,N_651,N_628);
xnor U812 (N_812,N_632,N_686);
xnor U813 (N_813,N_757,N_669);
xnor U814 (N_814,N_642,N_637);
nand U815 (N_815,N_645,N_631);
nand U816 (N_816,N_613,N_735);
or U817 (N_817,N_792,N_659);
and U818 (N_818,N_638,N_603);
xnor U819 (N_819,N_728,N_633);
nor U820 (N_820,N_676,N_783);
xnor U821 (N_821,N_724,N_799);
nor U822 (N_822,N_601,N_649);
xnor U823 (N_823,N_795,N_785);
xor U824 (N_824,N_718,N_781);
or U825 (N_825,N_607,N_709);
xnor U826 (N_826,N_667,N_652);
nand U827 (N_827,N_674,N_727);
and U828 (N_828,N_707,N_763);
and U829 (N_829,N_744,N_710);
or U830 (N_830,N_762,N_664);
or U831 (N_831,N_758,N_616);
nor U832 (N_832,N_730,N_600);
or U833 (N_833,N_729,N_775);
nand U834 (N_834,N_630,N_706);
xor U835 (N_835,N_754,N_746);
and U836 (N_836,N_764,N_656);
and U837 (N_837,N_786,N_793);
nor U838 (N_838,N_789,N_759);
xor U839 (N_839,N_647,N_643);
xnor U840 (N_840,N_620,N_722);
or U841 (N_841,N_691,N_719);
nor U842 (N_842,N_708,N_665);
nand U843 (N_843,N_703,N_687);
or U844 (N_844,N_773,N_769);
nand U845 (N_845,N_702,N_612);
xor U846 (N_846,N_602,N_611);
and U847 (N_847,N_767,N_662);
nor U848 (N_848,N_696,N_690);
xor U849 (N_849,N_716,N_742);
or U850 (N_850,N_692,N_747);
nor U851 (N_851,N_743,N_680);
or U852 (N_852,N_624,N_644);
nor U853 (N_853,N_617,N_663);
nand U854 (N_854,N_698,N_766);
xor U855 (N_855,N_768,N_650);
nand U856 (N_856,N_635,N_756);
and U857 (N_857,N_797,N_782);
xor U858 (N_858,N_604,N_614);
or U859 (N_859,N_788,N_639);
xnor U860 (N_860,N_646,N_666);
or U861 (N_861,N_731,N_741);
or U862 (N_862,N_694,N_771);
nor U863 (N_863,N_755,N_688);
or U864 (N_864,N_753,N_653);
nor U865 (N_865,N_761,N_658);
xnor U866 (N_866,N_699,N_749);
and U867 (N_867,N_750,N_794);
xor U868 (N_868,N_790,N_610);
nor U869 (N_869,N_752,N_791);
xnor U870 (N_870,N_720,N_751);
and U871 (N_871,N_736,N_704);
nand U872 (N_872,N_671,N_717);
or U873 (N_873,N_725,N_677);
or U874 (N_874,N_701,N_693);
nor U875 (N_875,N_654,N_619);
nand U876 (N_876,N_774,N_626);
xor U877 (N_877,N_796,N_661);
nor U878 (N_878,N_672,N_623);
nand U879 (N_879,N_609,N_678);
or U880 (N_880,N_737,N_679);
nor U881 (N_881,N_778,N_673);
and U882 (N_882,N_760,N_634);
nand U883 (N_883,N_784,N_608);
nand U884 (N_884,N_780,N_770);
and U885 (N_885,N_697,N_745);
xnor U886 (N_886,N_682,N_660);
nand U887 (N_887,N_636,N_695);
nand U888 (N_888,N_689,N_712);
and U889 (N_889,N_621,N_739);
xnor U890 (N_890,N_714,N_625);
and U891 (N_891,N_618,N_681);
or U892 (N_892,N_715,N_684);
xor U893 (N_893,N_705,N_772);
xor U894 (N_894,N_627,N_640);
and U895 (N_895,N_779,N_777);
nand U896 (N_896,N_641,N_675);
or U897 (N_897,N_738,N_700);
nor U898 (N_898,N_685,N_733);
or U899 (N_899,N_765,N_657);
and U900 (N_900,N_673,N_600);
nand U901 (N_901,N_727,N_601);
and U902 (N_902,N_694,N_763);
nand U903 (N_903,N_743,N_753);
nor U904 (N_904,N_667,N_635);
or U905 (N_905,N_707,N_765);
nor U906 (N_906,N_670,N_665);
nor U907 (N_907,N_678,N_657);
and U908 (N_908,N_728,N_740);
or U909 (N_909,N_600,N_651);
xnor U910 (N_910,N_638,N_755);
xor U911 (N_911,N_719,N_613);
and U912 (N_912,N_709,N_744);
nor U913 (N_913,N_777,N_739);
or U914 (N_914,N_689,N_725);
nand U915 (N_915,N_626,N_696);
nor U916 (N_916,N_770,N_658);
and U917 (N_917,N_713,N_778);
nand U918 (N_918,N_608,N_703);
nor U919 (N_919,N_766,N_760);
nand U920 (N_920,N_667,N_648);
nor U921 (N_921,N_623,N_615);
nor U922 (N_922,N_707,N_775);
or U923 (N_923,N_696,N_680);
nand U924 (N_924,N_737,N_624);
nor U925 (N_925,N_717,N_763);
xnor U926 (N_926,N_714,N_636);
xnor U927 (N_927,N_759,N_736);
or U928 (N_928,N_732,N_782);
nor U929 (N_929,N_611,N_688);
or U930 (N_930,N_751,N_765);
nand U931 (N_931,N_791,N_786);
nor U932 (N_932,N_647,N_640);
nor U933 (N_933,N_633,N_717);
nor U934 (N_934,N_731,N_798);
nand U935 (N_935,N_617,N_735);
and U936 (N_936,N_744,N_624);
nor U937 (N_937,N_648,N_729);
nand U938 (N_938,N_795,N_693);
nand U939 (N_939,N_659,N_650);
or U940 (N_940,N_683,N_759);
xor U941 (N_941,N_769,N_612);
or U942 (N_942,N_793,N_795);
and U943 (N_943,N_703,N_735);
and U944 (N_944,N_686,N_640);
nand U945 (N_945,N_680,N_734);
and U946 (N_946,N_749,N_645);
or U947 (N_947,N_668,N_662);
xnor U948 (N_948,N_747,N_768);
nor U949 (N_949,N_683,N_748);
nor U950 (N_950,N_745,N_620);
xor U951 (N_951,N_760,N_709);
nor U952 (N_952,N_691,N_739);
and U953 (N_953,N_748,N_636);
nand U954 (N_954,N_619,N_757);
and U955 (N_955,N_752,N_632);
nor U956 (N_956,N_604,N_741);
and U957 (N_957,N_673,N_712);
or U958 (N_958,N_677,N_689);
nor U959 (N_959,N_681,N_716);
or U960 (N_960,N_655,N_690);
nor U961 (N_961,N_684,N_763);
or U962 (N_962,N_696,N_656);
nor U963 (N_963,N_755,N_730);
nor U964 (N_964,N_736,N_617);
nor U965 (N_965,N_745,N_621);
nor U966 (N_966,N_761,N_669);
xnor U967 (N_967,N_676,N_613);
or U968 (N_968,N_741,N_656);
xnor U969 (N_969,N_678,N_618);
or U970 (N_970,N_653,N_647);
and U971 (N_971,N_749,N_680);
or U972 (N_972,N_752,N_766);
or U973 (N_973,N_732,N_760);
nor U974 (N_974,N_780,N_667);
or U975 (N_975,N_779,N_797);
nor U976 (N_976,N_758,N_780);
or U977 (N_977,N_635,N_708);
nor U978 (N_978,N_758,N_635);
nand U979 (N_979,N_778,N_604);
nor U980 (N_980,N_727,N_793);
or U981 (N_981,N_621,N_712);
nor U982 (N_982,N_657,N_704);
nand U983 (N_983,N_634,N_642);
or U984 (N_984,N_786,N_736);
and U985 (N_985,N_791,N_629);
and U986 (N_986,N_781,N_607);
nand U987 (N_987,N_757,N_618);
or U988 (N_988,N_623,N_663);
or U989 (N_989,N_753,N_728);
or U990 (N_990,N_779,N_766);
nand U991 (N_991,N_670,N_692);
xor U992 (N_992,N_664,N_783);
nand U993 (N_993,N_744,N_615);
and U994 (N_994,N_665,N_662);
xor U995 (N_995,N_727,N_747);
nor U996 (N_996,N_746,N_794);
nand U997 (N_997,N_681,N_707);
and U998 (N_998,N_778,N_684);
nor U999 (N_999,N_611,N_779);
xor U1000 (N_1000,N_833,N_867);
or U1001 (N_1001,N_970,N_848);
xnor U1002 (N_1002,N_850,N_870);
nor U1003 (N_1003,N_847,N_901);
xor U1004 (N_1004,N_990,N_812);
nor U1005 (N_1005,N_924,N_932);
nor U1006 (N_1006,N_974,N_834);
and U1007 (N_1007,N_895,N_839);
or U1008 (N_1008,N_897,N_816);
or U1009 (N_1009,N_982,N_918);
nand U1010 (N_1010,N_852,N_824);
nand U1011 (N_1011,N_937,N_800);
or U1012 (N_1012,N_960,N_996);
and U1013 (N_1013,N_920,N_963);
or U1014 (N_1014,N_859,N_994);
nor U1015 (N_1015,N_896,N_868);
xnor U1016 (N_1016,N_945,N_957);
and U1017 (N_1017,N_806,N_854);
nand U1018 (N_1018,N_909,N_843);
nor U1019 (N_1019,N_931,N_907);
xnor U1020 (N_1020,N_911,N_904);
nor U1021 (N_1021,N_878,N_899);
or U1022 (N_1022,N_876,N_914);
xnor U1023 (N_1023,N_978,N_803);
nor U1024 (N_1024,N_922,N_849);
nand U1025 (N_1025,N_884,N_823);
xnor U1026 (N_1026,N_998,N_964);
nor U1027 (N_1027,N_934,N_939);
and U1028 (N_1028,N_820,N_969);
or U1029 (N_1029,N_921,N_988);
and U1030 (N_1030,N_827,N_837);
xor U1031 (N_1031,N_925,N_866);
nor U1032 (N_1032,N_940,N_917);
and U1033 (N_1033,N_908,N_973);
and U1034 (N_1034,N_912,N_936);
xor U1035 (N_1035,N_900,N_822);
and U1036 (N_1036,N_976,N_802);
or U1037 (N_1037,N_894,N_818);
nand U1038 (N_1038,N_984,N_942);
xor U1039 (N_1039,N_814,N_983);
xnor U1040 (N_1040,N_811,N_910);
nand U1041 (N_1041,N_805,N_948);
nor U1042 (N_1042,N_966,N_882);
nand U1043 (N_1043,N_880,N_840);
or U1044 (N_1044,N_893,N_889);
or U1045 (N_1045,N_916,N_831);
xnor U1046 (N_1046,N_986,N_943);
nor U1047 (N_1047,N_951,N_846);
or U1048 (N_1048,N_863,N_985);
xnor U1049 (N_1049,N_875,N_980);
or U1050 (N_1050,N_926,N_923);
and U1051 (N_1051,N_828,N_968);
nor U1052 (N_1052,N_946,N_930);
and U1053 (N_1053,N_858,N_883);
nor U1054 (N_1054,N_887,N_913);
xor U1055 (N_1055,N_997,N_987);
or U1056 (N_1056,N_952,N_874);
xor U1057 (N_1057,N_941,N_979);
or U1058 (N_1058,N_993,N_999);
nor U1059 (N_1059,N_869,N_989);
nor U1060 (N_1060,N_864,N_872);
xor U1061 (N_1061,N_809,N_861);
xor U1062 (N_1062,N_873,N_842);
nor U1063 (N_1063,N_906,N_838);
nor U1064 (N_1064,N_845,N_959);
nand U1065 (N_1065,N_958,N_933);
nand U1066 (N_1066,N_905,N_855);
and U1067 (N_1067,N_857,N_881);
xnor U1068 (N_1068,N_832,N_836);
and U1069 (N_1069,N_853,N_808);
and U1070 (N_1070,N_991,N_927);
nand U1071 (N_1071,N_804,N_992);
and U1072 (N_1072,N_915,N_928);
and U1073 (N_1073,N_944,N_891);
nor U1074 (N_1074,N_947,N_871);
nor U1075 (N_1075,N_885,N_965);
and U1076 (N_1076,N_961,N_813);
nand U1077 (N_1077,N_844,N_971);
nand U1078 (N_1078,N_886,N_956);
xnor U1079 (N_1079,N_972,N_817);
nand U1080 (N_1080,N_877,N_954);
and U1081 (N_1081,N_967,N_856);
xor U1082 (N_1082,N_953,N_929);
nor U1083 (N_1083,N_950,N_801);
and U1084 (N_1084,N_865,N_995);
xor U1085 (N_1085,N_835,N_902);
and U1086 (N_1086,N_879,N_903);
or U1087 (N_1087,N_815,N_810);
nor U1088 (N_1088,N_888,N_935);
nand U1089 (N_1089,N_892,N_898);
and U1090 (N_1090,N_975,N_962);
nand U1091 (N_1091,N_819,N_841);
or U1092 (N_1092,N_829,N_919);
xnor U1093 (N_1093,N_890,N_807);
nand U1094 (N_1094,N_825,N_938);
nand U1095 (N_1095,N_821,N_981);
nor U1096 (N_1096,N_862,N_851);
nand U1097 (N_1097,N_826,N_955);
xnor U1098 (N_1098,N_949,N_977);
nand U1099 (N_1099,N_860,N_830);
nand U1100 (N_1100,N_925,N_847);
and U1101 (N_1101,N_819,N_822);
or U1102 (N_1102,N_886,N_974);
xnor U1103 (N_1103,N_897,N_920);
nor U1104 (N_1104,N_819,N_999);
nor U1105 (N_1105,N_961,N_898);
xor U1106 (N_1106,N_946,N_941);
or U1107 (N_1107,N_890,N_809);
nor U1108 (N_1108,N_859,N_979);
xor U1109 (N_1109,N_874,N_908);
nor U1110 (N_1110,N_835,N_953);
nor U1111 (N_1111,N_931,N_962);
nand U1112 (N_1112,N_831,N_942);
nor U1113 (N_1113,N_825,N_839);
and U1114 (N_1114,N_852,N_958);
and U1115 (N_1115,N_826,N_887);
nand U1116 (N_1116,N_823,N_855);
nor U1117 (N_1117,N_938,N_847);
xor U1118 (N_1118,N_815,N_820);
and U1119 (N_1119,N_992,N_934);
nand U1120 (N_1120,N_904,N_884);
nor U1121 (N_1121,N_919,N_941);
nand U1122 (N_1122,N_961,N_959);
or U1123 (N_1123,N_993,N_883);
nor U1124 (N_1124,N_809,N_883);
and U1125 (N_1125,N_922,N_927);
and U1126 (N_1126,N_870,N_845);
or U1127 (N_1127,N_996,N_864);
and U1128 (N_1128,N_934,N_962);
xor U1129 (N_1129,N_897,N_867);
xor U1130 (N_1130,N_964,N_819);
and U1131 (N_1131,N_814,N_876);
and U1132 (N_1132,N_910,N_838);
nand U1133 (N_1133,N_968,N_883);
xor U1134 (N_1134,N_914,N_857);
xnor U1135 (N_1135,N_843,N_903);
and U1136 (N_1136,N_873,N_809);
and U1137 (N_1137,N_956,N_969);
nor U1138 (N_1138,N_832,N_838);
or U1139 (N_1139,N_824,N_823);
nand U1140 (N_1140,N_860,N_925);
nor U1141 (N_1141,N_829,N_800);
or U1142 (N_1142,N_833,N_886);
or U1143 (N_1143,N_912,N_851);
nor U1144 (N_1144,N_983,N_957);
or U1145 (N_1145,N_941,N_976);
nor U1146 (N_1146,N_891,N_873);
nor U1147 (N_1147,N_897,N_850);
xor U1148 (N_1148,N_815,N_843);
and U1149 (N_1149,N_845,N_990);
nor U1150 (N_1150,N_995,N_821);
or U1151 (N_1151,N_963,N_885);
and U1152 (N_1152,N_987,N_866);
nand U1153 (N_1153,N_963,N_838);
xnor U1154 (N_1154,N_918,N_810);
xnor U1155 (N_1155,N_949,N_902);
or U1156 (N_1156,N_851,N_949);
or U1157 (N_1157,N_858,N_978);
nand U1158 (N_1158,N_892,N_895);
nor U1159 (N_1159,N_915,N_807);
nand U1160 (N_1160,N_807,N_878);
and U1161 (N_1161,N_912,N_940);
or U1162 (N_1162,N_854,N_851);
or U1163 (N_1163,N_932,N_975);
and U1164 (N_1164,N_978,N_906);
xor U1165 (N_1165,N_865,N_839);
nand U1166 (N_1166,N_879,N_845);
nor U1167 (N_1167,N_832,N_878);
xor U1168 (N_1168,N_953,N_821);
and U1169 (N_1169,N_936,N_910);
and U1170 (N_1170,N_823,N_896);
nand U1171 (N_1171,N_950,N_989);
or U1172 (N_1172,N_959,N_806);
nor U1173 (N_1173,N_915,N_835);
nand U1174 (N_1174,N_930,N_931);
xnor U1175 (N_1175,N_879,N_841);
nand U1176 (N_1176,N_999,N_871);
nand U1177 (N_1177,N_917,N_909);
nand U1178 (N_1178,N_988,N_832);
nand U1179 (N_1179,N_816,N_948);
or U1180 (N_1180,N_973,N_826);
nand U1181 (N_1181,N_938,N_827);
xnor U1182 (N_1182,N_903,N_815);
nand U1183 (N_1183,N_960,N_989);
and U1184 (N_1184,N_934,N_846);
nor U1185 (N_1185,N_933,N_812);
nand U1186 (N_1186,N_874,N_979);
xor U1187 (N_1187,N_880,N_895);
nor U1188 (N_1188,N_953,N_989);
xor U1189 (N_1189,N_929,N_974);
and U1190 (N_1190,N_966,N_845);
nor U1191 (N_1191,N_918,N_802);
nor U1192 (N_1192,N_918,N_938);
or U1193 (N_1193,N_807,N_838);
nand U1194 (N_1194,N_830,N_865);
or U1195 (N_1195,N_812,N_970);
nor U1196 (N_1196,N_878,N_846);
nor U1197 (N_1197,N_818,N_968);
and U1198 (N_1198,N_868,N_923);
xnor U1199 (N_1199,N_905,N_837);
and U1200 (N_1200,N_1189,N_1002);
or U1201 (N_1201,N_1158,N_1100);
and U1202 (N_1202,N_1043,N_1077);
or U1203 (N_1203,N_1029,N_1178);
nor U1204 (N_1204,N_1163,N_1152);
xnor U1205 (N_1205,N_1110,N_1062);
or U1206 (N_1206,N_1119,N_1056);
nor U1207 (N_1207,N_1097,N_1160);
and U1208 (N_1208,N_1113,N_1041);
nand U1209 (N_1209,N_1085,N_1096);
nand U1210 (N_1210,N_1023,N_1080);
xor U1211 (N_1211,N_1188,N_1084);
xor U1212 (N_1212,N_1187,N_1009);
and U1213 (N_1213,N_1014,N_1017);
or U1214 (N_1214,N_1156,N_1021);
xor U1215 (N_1215,N_1065,N_1054);
nor U1216 (N_1216,N_1185,N_1164);
xnor U1217 (N_1217,N_1015,N_1153);
nor U1218 (N_1218,N_1154,N_1000);
nor U1219 (N_1219,N_1073,N_1167);
and U1220 (N_1220,N_1070,N_1010);
xor U1221 (N_1221,N_1131,N_1087);
nand U1222 (N_1222,N_1127,N_1045);
and U1223 (N_1223,N_1033,N_1016);
nor U1224 (N_1224,N_1179,N_1137);
or U1225 (N_1225,N_1134,N_1012);
xnor U1226 (N_1226,N_1174,N_1061);
and U1227 (N_1227,N_1108,N_1175);
xnor U1228 (N_1228,N_1165,N_1025);
nor U1229 (N_1229,N_1095,N_1176);
nand U1230 (N_1230,N_1072,N_1150);
or U1231 (N_1231,N_1067,N_1183);
or U1232 (N_1232,N_1122,N_1120);
or U1233 (N_1233,N_1155,N_1032);
and U1234 (N_1234,N_1112,N_1143);
xor U1235 (N_1235,N_1079,N_1046);
xnor U1236 (N_1236,N_1173,N_1193);
xnor U1237 (N_1237,N_1049,N_1132);
nor U1238 (N_1238,N_1055,N_1138);
xnor U1239 (N_1239,N_1184,N_1081);
nand U1240 (N_1240,N_1013,N_1038);
xnor U1241 (N_1241,N_1007,N_1109);
and U1242 (N_1242,N_1166,N_1129);
or U1243 (N_1243,N_1196,N_1069);
and U1244 (N_1244,N_1036,N_1197);
nor U1245 (N_1245,N_1071,N_1181);
nor U1246 (N_1246,N_1058,N_1005);
and U1247 (N_1247,N_1082,N_1086);
nand U1248 (N_1248,N_1123,N_1111);
and U1249 (N_1249,N_1136,N_1141);
or U1250 (N_1250,N_1044,N_1116);
nand U1251 (N_1251,N_1075,N_1161);
xor U1252 (N_1252,N_1018,N_1117);
and U1253 (N_1253,N_1126,N_1028);
xor U1254 (N_1254,N_1140,N_1020);
xnor U1255 (N_1255,N_1051,N_1114);
nor U1256 (N_1256,N_1170,N_1064);
or U1257 (N_1257,N_1125,N_1074);
xor U1258 (N_1258,N_1001,N_1121);
or U1259 (N_1259,N_1004,N_1133);
or U1260 (N_1260,N_1130,N_1091);
xnor U1261 (N_1261,N_1157,N_1144);
or U1262 (N_1262,N_1052,N_1030);
and U1263 (N_1263,N_1198,N_1151);
xor U1264 (N_1264,N_1159,N_1146);
nor U1265 (N_1265,N_1078,N_1094);
or U1266 (N_1266,N_1019,N_1191);
xor U1267 (N_1267,N_1060,N_1171);
and U1268 (N_1268,N_1124,N_1008);
and U1269 (N_1269,N_1149,N_1059);
or U1270 (N_1270,N_1106,N_1148);
nor U1271 (N_1271,N_1199,N_1092);
or U1272 (N_1272,N_1022,N_1047);
or U1273 (N_1273,N_1195,N_1066);
xor U1274 (N_1274,N_1006,N_1050);
or U1275 (N_1275,N_1168,N_1105);
or U1276 (N_1276,N_1090,N_1135);
nand U1277 (N_1277,N_1169,N_1011);
and U1278 (N_1278,N_1180,N_1088);
or U1279 (N_1279,N_1039,N_1031);
nand U1280 (N_1280,N_1142,N_1040);
nor U1281 (N_1281,N_1093,N_1177);
and U1282 (N_1282,N_1103,N_1076);
xor U1283 (N_1283,N_1063,N_1102);
nor U1284 (N_1284,N_1034,N_1068);
nor U1285 (N_1285,N_1037,N_1147);
nand U1286 (N_1286,N_1190,N_1053);
nor U1287 (N_1287,N_1118,N_1057);
xor U1288 (N_1288,N_1182,N_1098);
or U1289 (N_1289,N_1048,N_1162);
nor U1290 (N_1290,N_1128,N_1107);
and U1291 (N_1291,N_1035,N_1083);
nor U1292 (N_1292,N_1027,N_1115);
xor U1293 (N_1293,N_1194,N_1145);
or U1294 (N_1294,N_1186,N_1104);
nand U1295 (N_1295,N_1192,N_1026);
or U1296 (N_1296,N_1172,N_1024);
or U1297 (N_1297,N_1101,N_1003);
and U1298 (N_1298,N_1042,N_1139);
nor U1299 (N_1299,N_1089,N_1099);
and U1300 (N_1300,N_1113,N_1138);
xnor U1301 (N_1301,N_1061,N_1074);
nand U1302 (N_1302,N_1017,N_1169);
nand U1303 (N_1303,N_1183,N_1078);
nand U1304 (N_1304,N_1008,N_1180);
xor U1305 (N_1305,N_1100,N_1174);
xor U1306 (N_1306,N_1012,N_1049);
nand U1307 (N_1307,N_1094,N_1150);
and U1308 (N_1308,N_1058,N_1191);
or U1309 (N_1309,N_1073,N_1197);
nand U1310 (N_1310,N_1064,N_1159);
and U1311 (N_1311,N_1057,N_1131);
or U1312 (N_1312,N_1113,N_1124);
nor U1313 (N_1313,N_1109,N_1079);
nand U1314 (N_1314,N_1196,N_1003);
and U1315 (N_1315,N_1193,N_1145);
or U1316 (N_1316,N_1190,N_1116);
or U1317 (N_1317,N_1107,N_1062);
and U1318 (N_1318,N_1156,N_1100);
nand U1319 (N_1319,N_1184,N_1082);
nor U1320 (N_1320,N_1158,N_1077);
nand U1321 (N_1321,N_1009,N_1132);
xnor U1322 (N_1322,N_1161,N_1097);
and U1323 (N_1323,N_1002,N_1102);
and U1324 (N_1324,N_1028,N_1189);
xor U1325 (N_1325,N_1192,N_1070);
xnor U1326 (N_1326,N_1003,N_1042);
nor U1327 (N_1327,N_1074,N_1154);
and U1328 (N_1328,N_1158,N_1018);
or U1329 (N_1329,N_1170,N_1115);
or U1330 (N_1330,N_1071,N_1120);
nand U1331 (N_1331,N_1129,N_1050);
xnor U1332 (N_1332,N_1128,N_1041);
nand U1333 (N_1333,N_1115,N_1089);
nand U1334 (N_1334,N_1178,N_1165);
xnor U1335 (N_1335,N_1101,N_1087);
or U1336 (N_1336,N_1079,N_1106);
nand U1337 (N_1337,N_1039,N_1102);
or U1338 (N_1338,N_1059,N_1062);
nand U1339 (N_1339,N_1014,N_1153);
xnor U1340 (N_1340,N_1086,N_1000);
nand U1341 (N_1341,N_1121,N_1107);
xnor U1342 (N_1342,N_1138,N_1141);
or U1343 (N_1343,N_1109,N_1158);
nand U1344 (N_1344,N_1138,N_1002);
xor U1345 (N_1345,N_1197,N_1138);
and U1346 (N_1346,N_1043,N_1186);
nor U1347 (N_1347,N_1023,N_1090);
and U1348 (N_1348,N_1011,N_1100);
and U1349 (N_1349,N_1088,N_1198);
and U1350 (N_1350,N_1184,N_1131);
nand U1351 (N_1351,N_1127,N_1001);
nand U1352 (N_1352,N_1193,N_1023);
nand U1353 (N_1353,N_1027,N_1158);
or U1354 (N_1354,N_1036,N_1034);
xnor U1355 (N_1355,N_1189,N_1172);
and U1356 (N_1356,N_1157,N_1194);
xnor U1357 (N_1357,N_1187,N_1074);
nor U1358 (N_1358,N_1195,N_1122);
and U1359 (N_1359,N_1029,N_1163);
nor U1360 (N_1360,N_1149,N_1063);
nor U1361 (N_1361,N_1029,N_1019);
xnor U1362 (N_1362,N_1124,N_1012);
xnor U1363 (N_1363,N_1045,N_1172);
or U1364 (N_1364,N_1138,N_1067);
and U1365 (N_1365,N_1088,N_1172);
xnor U1366 (N_1366,N_1182,N_1194);
xor U1367 (N_1367,N_1070,N_1182);
nor U1368 (N_1368,N_1024,N_1170);
and U1369 (N_1369,N_1172,N_1128);
or U1370 (N_1370,N_1033,N_1154);
nand U1371 (N_1371,N_1042,N_1121);
xnor U1372 (N_1372,N_1155,N_1092);
and U1373 (N_1373,N_1008,N_1138);
xor U1374 (N_1374,N_1171,N_1152);
and U1375 (N_1375,N_1002,N_1146);
and U1376 (N_1376,N_1166,N_1080);
and U1377 (N_1377,N_1188,N_1135);
or U1378 (N_1378,N_1094,N_1025);
nor U1379 (N_1379,N_1063,N_1002);
or U1380 (N_1380,N_1027,N_1061);
and U1381 (N_1381,N_1054,N_1038);
nand U1382 (N_1382,N_1090,N_1032);
or U1383 (N_1383,N_1128,N_1188);
and U1384 (N_1384,N_1012,N_1110);
and U1385 (N_1385,N_1162,N_1039);
nor U1386 (N_1386,N_1187,N_1068);
and U1387 (N_1387,N_1031,N_1118);
nor U1388 (N_1388,N_1189,N_1084);
and U1389 (N_1389,N_1133,N_1015);
or U1390 (N_1390,N_1025,N_1133);
xnor U1391 (N_1391,N_1095,N_1022);
nor U1392 (N_1392,N_1081,N_1025);
and U1393 (N_1393,N_1127,N_1003);
and U1394 (N_1394,N_1096,N_1041);
and U1395 (N_1395,N_1198,N_1180);
or U1396 (N_1396,N_1145,N_1153);
and U1397 (N_1397,N_1094,N_1031);
and U1398 (N_1398,N_1080,N_1132);
xnor U1399 (N_1399,N_1183,N_1006);
or U1400 (N_1400,N_1234,N_1320);
and U1401 (N_1401,N_1392,N_1307);
nor U1402 (N_1402,N_1325,N_1338);
and U1403 (N_1403,N_1237,N_1354);
xnor U1404 (N_1404,N_1309,N_1371);
and U1405 (N_1405,N_1351,N_1229);
nand U1406 (N_1406,N_1274,N_1321);
or U1407 (N_1407,N_1296,N_1258);
and U1408 (N_1408,N_1323,N_1376);
nor U1409 (N_1409,N_1260,N_1275);
or U1410 (N_1410,N_1399,N_1250);
and U1411 (N_1411,N_1304,N_1340);
or U1412 (N_1412,N_1339,N_1386);
or U1413 (N_1413,N_1330,N_1231);
and U1414 (N_1414,N_1252,N_1383);
nand U1415 (N_1415,N_1389,N_1302);
nand U1416 (N_1416,N_1397,N_1335);
or U1417 (N_1417,N_1380,N_1227);
nor U1418 (N_1418,N_1262,N_1295);
xnor U1419 (N_1419,N_1347,N_1301);
nor U1420 (N_1420,N_1255,N_1271);
nor U1421 (N_1421,N_1220,N_1328);
and U1422 (N_1422,N_1310,N_1205);
or U1423 (N_1423,N_1344,N_1261);
or U1424 (N_1424,N_1221,N_1239);
nand U1425 (N_1425,N_1379,N_1242);
nor U1426 (N_1426,N_1342,N_1305);
xnor U1427 (N_1427,N_1289,N_1358);
xnor U1428 (N_1428,N_1228,N_1348);
or U1429 (N_1429,N_1212,N_1312);
and U1430 (N_1430,N_1286,N_1284);
xor U1431 (N_1431,N_1355,N_1254);
and U1432 (N_1432,N_1230,N_1269);
or U1433 (N_1433,N_1246,N_1277);
or U1434 (N_1434,N_1243,N_1236);
nand U1435 (N_1435,N_1224,N_1327);
xnor U1436 (N_1436,N_1353,N_1385);
xnor U1437 (N_1437,N_1217,N_1247);
or U1438 (N_1438,N_1341,N_1244);
nand U1439 (N_1439,N_1362,N_1281);
nand U1440 (N_1440,N_1334,N_1349);
nand U1441 (N_1441,N_1282,N_1293);
nor U1442 (N_1442,N_1387,N_1273);
or U1443 (N_1443,N_1360,N_1209);
or U1444 (N_1444,N_1369,N_1241);
or U1445 (N_1445,N_1300,N_1337);
nor U1446 (N_1446,N_1366,N_1216);
nand U1447 (N_1447,N_1226,N_1265);
xnor U1448 (N_1448,N_1336,N_1288);
and U1449 (N_1449,N_1391,N_1257);
and U1450 (N_1450,N_1393,N_1390);
xnor U1451 (N_1451,N_1382,N_1233);
xnor U1452 (N_1452,N_1331,N_1316);
and U1453 (N_1453,N_1238,N_1395);
and U1454 (N_1454,N_1364,N_1333);
nor U1455 (N_1455,N_1245,N_1291);
nand U1456 (N_1456,N_1368,N_1365);
nand U1457 (N_1457,N_1378,N_1235);
or U1458 (N_1458,N_1208,N_1232);
nor U1459 (N_1459,N_1319,N_1279);
nand U1460 (N_1460,N_1346,N_1259);
nand U1461 (N_1461,N_1329,N_1350);
nor U1462 (N_1462,N_1213,N_1200);
nor U1463 (N_1463,N_1357,N_1314);
nand U1464 (N_1464,N_1240,N_1270);
nand U1465 (N_1465,N_1370,N_1207);
or U1466 (N_1466,N_1278,N_1372);
or U1467 (N_1467,N_1377,N_1367);
xor U1468 (N_1468,N_1266,N_1373);
nor U1469 (N_1469,N_1253,N_1332);
nor U1470 (N_1470,N_1214,N_1363);
nand U1471 (N_1471,N_1287,N_1272);
or U1472 (N_1472,N_1361,N_1264);
or U1473 (N_1473,N_1326,N_1268);
xor U1474 (N_1474,N_1248,N_1203);
xnor U1475 (N_1475,N_1317,N_1294);
and U1476 (N_1476,N_1204,N_1315);
nor U1477 (N_1477,N_1218,N_1345);
or U1478 (N_1478,N_1256,N_1299);
nor U1479 (N_1479,N_1343,N_1306);
or U1480 (N_1480,N_1381,N_1313);
nand U1481 (N_1481,N_1374,N_1311);
nor U1482 (N_1482,N_1276,N_1303);
nand U1483 (N_1483,N_1225,N_1388);
nand U1484 (N_1484,N_1280,N_1285);
and U1485 (N_1485,N_1298,N_1202);
nand U1486 (N_1486,N_1283,N_1297);
xor U1487 (N_1487,N_1267,N_1206);
nor U1488 (N_1488,N_1396,N_1211);
xnor U1489 (N_1489,N_1251,N_1263);
and U1490 (N_1490,N_1219,N_1394);
and U1491 (N_1491,N_1215,N_1308);
nand U1492 (N_1492,N_1384,N_1201);
or U1493 (N_1493,N_1375,N_1356);
nor U1494 (N_1494,N_1318,N_1398);
and U1495 (N_1495,N_1324,N_1290);
xor U1496 (N_1496,N_1222,N_1359);
or U1497 (N_1497,N_1249,N_1352);
and U1498 (N_1498,N_1322,N_1210);
or U1499 (N_1499,N_1223,N_1292);
and U1500 (N_1500,N_1202,N_1223);
or U1501 (N_1501,N_1341,N_1305);
nor U1502 (N_1502,N_1366,N_1331);
nor U1503 (N_1503,N_1389,N_1232);
nor U1504 (N_1504,N_1356,N_1352);
nand U1505 (N_1505,N_1396,N_1375);
xor U1506 (N_1506,N_1284,N_1264);
or U1507 (N_1507,N_1371,N_1249);
nor U1508 (N_1508,N_1320,N_1289);
xor U1509 (N_1509,N_1352,N_1247);
or U1510 (N_1510,N_1325,N_1219);
or U1511 (N_1511,N_1238,N_1281);
or U1512 (N_1512,N_1379,N_1228);
nand U1513 (N_1513,N_1225,N_1236);
or U1514 (N_1514,N_1288,N_1308);
or U1515 (N_1515,N_1366,N_1286);
and U1516 (N_1516,N_1214,N_1302);
and U1517 (N_1517,N_1212,N_1356);
nor U1518 (N_1518,N_1369,N_1367);
xnor U1519 (N_1519,N_1248,N_1285);
nor U1520 (N_1520,N_1236,N_1253);
or U1521 (N_1521,N_1206,N_1341);
or U1522 (N_1522,N_1265,N_1231);
nand U1523 (N_1523,N_1354,N_1378);
and U1524 (N_1524,N_1330,N_1317);
or U1525 (N_1525,N_1377,N_1343);
nor U1526 (N_1526,N_1291,N_1369);
nand U1527 (N_1527,N_1338,N_1342);
or U1528 (N_1528,N_1309,N_1295);
and U1529 (N_1529,N_1229,N_1360);
nor U1530 (N_1530,N_1393,N_1327);
nor U1531 (N_1531,N_1240,N_1283);
nand U1532 (N_1532,N_1345,N_1334);
or U1533 (N_1533,N_1379,N_1357);
nand U1534 (N_1534,N_1254,N_1273);
or U1535 (N_1535,N_1233,N_1345);
or U1536 (N_1536,N_1377,N_1355);
nor U1537 (N_1537,N_1248,N_1284);
xor U1538 (N_1538,N_1349,N_1270);
nand U1539 (N_1539,N_1294,N_1309);
nor U1540 (N_1540,N_1275,N_1299);
and U1541 (N_1541,N_1310,N_1295);
or U1542 (N_1542,N_1218,N_1324);
nand U1543 (N_1543,N_1369,N_1330);
nand U1544 (N_1544,N_1238,N_1394);
or U1545 (N_1545,N_1304,N_1249);
nor U1546 (N_1546,N_1252,N_1382);
nand U1547 (N_1547,N_1297,N_1230);
and U1548 (N_1548,N_1206,N_1228);
or U1549 (N_1549,N_1362,N_1349);
and U1550 (N_1550,N_1390,N_1290);
nand U1551 (N_1551,N_1387,N_1260);
and U1552 (N_1552,N_1284,N_1204);
nand U1553 (N_1553,N_1272,N_1267);
or U1554 (N_1554,N_1397,N_1280);
nand U1555 (N_1555,N_1268,N_1229);
xnor U1556 (N_1556,N_1294,N_1301);
or U1557 (N_1557,N_1222,N_1347);
nor U1558 (N_1558,N_1378,N_1310);
or U1559 (N_1559,N_1347,N_1371);
nor U1560 (N_1560,N_1210,N_1378);
nand U1561 (N_1561,N_1232,N_1260);
nor U1562 (N_1562,N_1217,N_1209);
and U1563 (N_1563,N_1367,N_1327);
or U1564 (N_1564,N_1290,N_1391);
nand U1565 (N_1565,N_1331,N_1280);
nor U1566 (N_1566,N_1328,N_1259);
or U1567 (N_1567,N_1283,N_1222);
nor U1568 (N_1568,N_1204,N_1385);
nor U1569 (N_1569,N_1304,N_1225);
nand U1570 (N_1570,N_1355,N_1262);
and U1571 (N_1571,N_1382,N_1211);
xnor U1572 (N_1572,N_1278,N_1218);
nor U1573 (N_1573,N_1398,N_1334);
or U1574 (N_1574,N_1358,N_1200);
xnor U1575 (N_1575,N_1397,N_1330);
nor U1576 (N_1576,N_1246,N_1240);
and U1577 (N_1577,N_1222,N_1345);
nand U1578 (N_1578,N_1348,N_1235);
nor U1579 (N_1579,N_1332,N_1315);
or U1580 (N_1580,N_1351,N_1303);
and U1581 (N_1581,N_1300,N_1265);
or U1582 (N_1582,N_1319,N_1293);
and U1583 (N_1583,N_1310,N_1252);
and U1584 (N_1584,N_1229,N_1236);
and U1585 (N_1585,N_1283,N_1301);
nor U1586 (N_1586,N_1244,N_1309);
or U1587 (N_1587,N_1329,N_1253);
nor U1588 (N_1588,N_1253,N_1375);
xor U1589 (N_1589,N_1327,N_1380);
xor U1590 (N_1590,N_1370,N_1267);
nor U1591 (N_1591,N_1346,N_1351);
or U1592 (N_1592,N_1375,N_1385);
or U1593 (N_1593,N_1301,N_1303);
nor U1594 (N_1594,N_1318,N_1200);
and U1595 (N_1595,N_1371,N_1294);
xnor U1596 (N_1596,N_1305,N_1217);
xor U1597 (N_1597,N_1297,N_1236);
nand U1598 (N_1598,N_1289,N_1375);
xor U1599 (N_1599,N_1253,N_1255);
and U1600 (N_1600,N_1578,N_1505);
xor U1601 (N_1601,N_1510,N_1575);
xor U1602 (N_1602,N_1560,N_1572);
and U1603 (N_1603,N_1412,N_1467);
or U1604 (N_1604,N_1498,N_1537);
nor U1605 (N_1605,N_1503,N_1546);
or U1606 (N_1606,N_1594,N_1584);
nand U1607 (N_1607,N_1490,N_1436);
xor U1608 (N_1608,N_1532,N_1434);
nand U1609 (N_1609,N_1554,N_1448);
and U1610 (N_1610,N_1471,N_1564);
nand U1611 (N_1611,N_1568,N_1496);
nand U1612 (N_1612,N_1463,N_1414);
xnor U1613 (N_1613,N_1542,N_1550);
xnor U1614 (N_1614,N_1566,N_1509);
or U1615 (N_1615,N_1459,N_1426);
xor U1616 (N_1616,N_1598,N_1423);
or U1617 (N_1617,N_1461,N_1494);
nand U1618 (N_1618,N_1438,N_1526);
nand U1619 (N_1619,N_1429,N_1403);
xnor U1620 (N_1620,N_1504,N_1480);
xnor U1621 (N_1621,N_1474,N_1535);
nand U1622 (N_1622,N_1472,N_1432);
nor U1623 (N_1623,N_1405,N_1430);
nand U1624 (N_1624,N_1497,N_1457);
or U1625 (N_1625,N_1588,N_1541);
or U1626 (N_1626,N_1417,N_1529);
and U1627 (N_1627,N_1407,N_1402);
nor U1628 (N_1628,N_1516,N_1593);
nor U1629 (N_1629,N_1525,N_1439);
and U1630 (N_1630,N_1443,N_1538);
and U1631 (N_1631,N_1431,N_1413);
or U1632 (N_1632,N_1507,N_1482);
nor U1633 (N_1633,N_1419,N_1580);
and U1634 (N_1634,N_1454,N_1552);
nor U1635 (N_1635,N_1523,N_1577);
nand U1636 (N_1636,N_1519,N_1492);
nand U1637 (N_1637,N_1437,N_1478);
or U1638 (N_1638,N_1597,N_1487);
nor U1639 (N_1639,N_1565,N_1420);
nand U1640 (N_1640,N_1585,N_1514);
nor U1641 (N_1641,N_1473,N_1571);
xnor U1642 (N_1642,N_1469,N_1530);
or U1643 (N_1643,N_1488,N_1421);
or U1644 (N_1644,N_1485,N_1524);
and U1645 (N_1645,N_1415,N_1460);
and U1646 (N_1646,N_1586,N_1531);
nor U1647 (N_1647,N_1547,N_1567);
and U1648 (N_1648,N_1518,N_1579);
nand U1649 (N_1649,N_1596,N_1553);
nand U1650 (N_1650,N_1528,N_1455);
and U1651 (N_1651,N_1587,N_1483);
nor U1652 (N_1652,N_1540,N_1477);
nor U1653 (N_1653,N_1447,N_1555);
xnor U1654 (N_1654,N_1539,N_1549);
nor U1655 (N_1655,N_1570,N_1410);
nor U1656 (N_1656,N_1446,N_1449);
and U1657 (N_1657,N_1453,N_1557);
xor U1658 (N_1658,N_1527,N_1464);
xnor U1659 (N_1659,N_1515,N_1562);
xor U1660 (N_1660,N_1573,N_1559);
nand U1661 (N_1661,N_1400,N_1409);
and U1662 (N_1662,N_1468,N_1501);
and U1663 (N_1663,N_1445,N_1581);
nand U1664 (N_1664,N_1408,N_1563);
or U1665 (N_1665,N_1479,N_1574);
or U1666 (N_1666,N_1545,N_1595);
nor U1667 (N_1667,N_1544,N_1591);
or U1668 (N_1668,N_1416,N_1489);
nand U1669 (N_1669,N_1599,N_1442);
or U1670 (N_1670,N_1592,N_1561);
xnor U1671 (N_1671,N_1558,N_1536);
nor U1672 (N_1672,N_1456,N_1458);
xnor U1673 (N_1673,N_1441,N_1401);
xnor U1674 (N_1674,N_1590,N_1404);
or U1675 (N_1675,N_1521,N_1534);
nand U1676 (N_1676,N_1440,N_1517);
or U1677 (N_1677,N_1502,N_1486);
and U1678 (N_1678,N_1425,N_1452);
or U1679 (N_1679,N_1499,N_1511);
or U1680 (N_1680,N_1556,N_1533);
nand U1681 (N_1681,N_1481,N_1424);
nor U1682 (N_1682,N_1495,N_1422);
nand U1683 (N_1683,N_1428,N_1548);
xor U1684 (N_1684,N_1513,N_1520);
or U1685 (N_1685,N_1476,N_1444);
or U1686 (N_1686,N_1522,N_1465);
and U1687 (N_1687,N_1450,N_1475);
xnor U1688 (N_1688,N_1411,N_1493);
xnor U1689 (N_1689,N_1582,N_1569);
and U1690 (N_1690,N_1500,N_1470);
and U1691 (N_1691,N_1543,N_1491);
nand U1692 (N_1692,N_1418,N_1466);
nand U1693 (N_1693,N_1484,N_1451);
nor U1694 (N_1694,N_1435,N_1551);
and U1695 (N_1695,N_1406,N_1583);
xnor U1696 (N_1696,N_1433,N_1506);
nand U1697 (N_1697,N_1462,N_1589);
xor U1698 (N_1698,N_1427,N_1576);
and U1699 (N_1699,N_1512,N_1508);
nor U1700 (N_1700,N_1560,N_1422);
xor U1701 (N_1701,N_1517,N_1472);
nand U1702 (N_1702,N_1415,N_1502);
nor U1703 (N_1703,N_1559,N_1532);
nor U1704 (N_1704,N_1495,N_1413);
xnor U1705 (N_1705,N_1458,N_1479);
xor U1706 (N_1706,N_1557,N_1420);
nor U1707 (N_1707,N_1563,N_1501);
and U1708 (N_1708,N_1410,N_1428);
nor U1709 (N_1709,N_1556,N_1559);
nand U1710 (N_1710,N_1424,N_1579);
nand U1711 (N_1711,N_1498,N_1597);
or U1712 (N_1712,N_1413,N_1566);
or U1713 (N_1713,N_1499,N_1402);
nor U1714 (N_1714,N_1481,N_1578);
and U1715 (N_1715,N_1409,N_1401);
or U1716 (N_1716,N_1432,N_1493);
or U1717 (N_1717,N_1430,N_1435);
nand U1718 (N_1718,N_1464,N_1558);
xor U1719 (N_1719,N_1486,N_1573);
nand U1720 (N_1720,N_1417,N_1557);
or U1721 (N_1721,N_1443,N_1529);
nand U1722 (N_1722,N_1477,N_1518);
nand U1723 (N_1723,N_1560,N_1577);
and U1724 (N_1724,N_1540,N_1515);
and U1725 (N_1725,N_1590,N_1501);
nand U1726 (N_1726,N_1499,N_1559);
nor U1727 (N_1727,N_1522,N_1448);
xor U1728 (N_1728,N_1527,N_1433);
or U1729 (N_1729,N_1420,N_1418);
or U1730 (N_1730,N_1413,N_1461);
nor U1731 (N_1731,N_1578,N_1533);
nor U1732 (N_1732,N_1455,N_1428);
and U1733 (N_1733,N_1504,N_1458);
or U1734 (N_1734,N_1538,N_1426);
or U1735 (N_1735,N_1467,N_1462);
nor U1736 (N_1736,N_1546,N_1417);
nand U1737 (N_1737,N_1482,N_1486);
and U1738 (N_1738,N_1599,N_1456);
and U1739 (N_1739,N_1553,N_1505);
or U1740 (N_1740,N_1427,N_1549);
and U1741 (N_1741,N_1417,N_1523);
or U1742 (N_1742,N_1478,N_1534);
or U1743 (N_1743,N_1407,N_1541);
nand U1744 (N_1744,N_1472,N_1582);
or U1745 (N_1745,N_1441,N_1428);
or U1746 (N_1746,N_1544,N_1469);
or U1747 (N_1747,N_1525,N_1588);
or U1748 (N_1748,N_1561,N_1535);
and U1749 (N_1749,N_1585,N_1483);
or U1750 (N_1750,N_1546,N_1493);
nand U1751 (N_1751,N_1532,N_1444);
and U1752 (N_1752,N_1508,N_1591);
nand U1753 (N_1753,N_1453,N_1579);
nand U1754 (N_1754,N_1482,N_1516);
xnor U1755 (N_1755,N_1503,N_1574);
nor U1756 (N_1756,N_1430,N_1540);
xnor U1757 (N_1757,N_1556,N_1560);
and U1758 (N_1758,N_1412,N_1583);
or U1759 (N_1759,N_1583,N_1519);
xor U1760 (N_1760,N_1442,N_1520);
and U1761 (N_1761,N_1534,N_1567);
or U1762 (N_1762,N_1458,N_1525);
nor U1763 (N_1763,N_1559,N_1512);
xor U1764 (N_1764,N_1506,N_1451);
or U1765 (N_1765,N_1567,N_1423);
and U1766 (N_1766,N_1499,N_1532);
nor U1767 (N_1767,N_1479,N_1514);
nand U1768 (N_1768,N_1510,N_1468);
nor U1769 (N_1769,N_1490,N_1466);
xnor U1770 (N_1770,N_1509,N_1513);
or U1771 (N_1771,N_1451,N_1548);
nor U1772 (N_1772,N_1462,N_1503);
xor U1773 (N_1773,N_1464,N_1576);
xor U1774 (N_1774,N_1433,N_1574);
nor U1775 (N_1775,N_1443,N_1503);
or U1776 (N_1776,N_1523,N_1427);
and U1777 (N_1777,N_1401,N_1538);
nand U1778 (N_1778,N_1501,N_1409);
and U1779 (N_1779,N_1477,N_1501);
or U1780 (N_1780,N_1422,N_1528);
nor U1781 (N_1781,N_1569,N_1545);
or U1782 (N_1782,N_1556,N_1439);
nand U1783 (N_1783,N_1493,N_1491);
xor U1784 (N_1784,N_1451,N_1592);
and U1785 (N_1785,N_1545,N_1556);
nand U1786 (N_1786,N_1400,N_1421);
xnor U1787 (N_1787,N_1492,N_1437);
or U1788 (N_1788,N_1431,N_1555);
nand U1789 (N_1789,N_1565,N_1522);
or U1790 (N_1790,N_1468,N_1401);
or U1791 (N_1791,N_1452,N_1418);
nor U1792 (N_1792,N_1544,N_1503);
nand U1793 (N_1793,N_1568,N_1514);
nand U1794 (N_1794,N_1564,N_1557);
or U1795 (N_1795,N_1437,N_1587);
or U1796 (N_1796,N_1582,N_1508);
xnor U1797 (N_1797,N_1407,N_1424);
nand U1798 (N_1798,N_1463,N_1522);
and U1799 (N_1799,N_1545,N_1439);
or U1800 (N_1800,N_1727,N_1706);
and U1801 (N_1801,N_1742,N_1689);
nand U1802 (N_1802,N_1781,N_1693);
and U1803 (N_1803,N_1739,N_1671);
and U1804 (N_1804,N_1798,N_1780);
nor U1805 (N_1805,N_1684,N_1743);
nand U1806 (N_1806,N_1772,N_1711);
and U1807 (N_1807,N_1606,N_1696);
and U1808 (N_1808,N_1767,N_1650);
and U1809 (N_1809,N_1732,N_1627);
xor U1810 (N_1810,N_1701,N_1687);
or U1811 (N_1811,N_1611,N_1628);
xnor U1812 (N_1812,N_1635,N_1709);
and U1813 (N_1813,N_1786,N_1640);
nand U1814 (N_1814,N_1788,N_1753);
or U1815 (N_1815,N_1631,N_1661);
nor U1816 (N_1816,N_1641,N_1700);
and U1817 (N_1817,N_1707,N_1715);
or U1818 (N_1818,N_1737,N_1769);
or U1819 (N_1819,N_1785,N_1666);
and U1820 (N_1820,N_1698,N_1680);
xor U1821 (N_1821,N_1756,N_1676);
and U1822 (N_1822,N_1605,N_1622);
xor U1823 (N_1823,N_1674,N_1642);
nor U1824 (N_1824,N_1738,N_1757);
nand U1825 (N_1825,N_1765,N_1665);
nand U1826 (N_1826,N_1751,N_1600);
nor U1827 (N_1827,N_1710,N_1621);
xor U1828 (N_1828,N_1691,N_1759);
nor U1829 (N_1829,N_1662,N_1784);
nor U1830 (N_1830,N_1720,N_1673);
or U1831 (N_1831,N_1768,N_1690);
nand U1832 (N_1832,N_1633,N_1758);
and U1833 (N_1833,N_1754,N_1744);
nand U1834 (N_1834,N_1668,N_1736);
or U1835 (N_1835,N_1723,N_1764);
or U1836 (N_1836,N_1649,N_1774);
nand U1837 (N_1837,N_1614,N_1638);
and U1838 (N_1838,N_1797,N_1799);
xor U1839 (N_1839,N_1770,N_1783);
and U1840 (N_1840,N_1603,N_1717);
nand U1841 (N_1841,N_1672,N_1714);
and U1842 (N_1842,N_1705,N_1771);
nand U1843 (N_1843,N_1669,N_1643);
nand U1844 (N_1844,N_1636,N_1791);
nor U1845 (N_1845,N_1721,N_1664);
or U1846 (N_1846,N_1763,N_1745);
nand U1847 (N_1847,N_1708,N_1777);
and U1848 (N_1848,N_1703,N_1761);
nand U1849 (N_1849,N_1694,N_1681);
or U1850 (N_1850,N_1660,N_1652);
xnor U1851 (N_1851,N_1655,N_1794);
nand U1852 (N_1852,N_1644,N_1733);
xnor U1853 (N_1853,N_1702,N_1778);
or U1854 (N_1854,N_1730,N_1601);
nor U1855 (N_1855,N_1697,N_1752);
nand U1856 (N_1856,N_1716,N_1724);
and U1857 (N_1857,N_1740,N_1729);
xnor U1858 (N_1858,N_1648,N_1760);
or U1859 (N_1859,N_1677,N_1735);
xnor U1860 (N_1860,N_1773,N_1670);
or U1861 (N_1861,N_1625,N_1645);
or U1862 (N_1862,N_1747,N_1615);
or U1863 (N_1863,N_1675,N_1748);
nor U1864 (N_1864,N_1719,N_1775);
and U1865 (N_1865,N_1617,N_1604);
and U1866 (N_1866,N_1779,N_1612);
and U1867 (N_1867,N_1679,N_1699);
and U1868 (N_1868,N_1790,N_1678);
xor U1869 (N_1869,N_1792,N_1646);
and U1870 (N_1870,N_1731,N_1782);
nand U1871 (N_1871,N_1762,N_1616);
or U1872 (N_1872,N_1629,N_1634);
nor U1873 (N_1873,N_1658,N_1607);
or U1874 (N_1874,N_1657,N_1750);
nand U1875 (N_1875,N_1695,N_1647);
and U1876 (N_1876,N_1682,N_1632);
and U1877 (N_1877,N_1722,N_1776);
nor U1878 (N_1878,N_1718,N_1725);
or U1879 (N_1879,N_1796,N_1686);
xor U1880 (N_1880,N_1626,N_1746);
nand U1881 (N_1881,N_1704,N_1624);
nand U1882 (N_1882,N_1630,N_1712);
xnor U1883 (N_1883,N_1659,N_1602);
and U1884 (N_1884,N_1637,N_1749);
and U1885 (N_1885,N_1713,N_1610);
or U1886 (N_1886,N_1618,N_1728);
nor U1887 (N_1887,N_1741,N_1688);
or U1888 (N_1888,N_1608,N_1726);
or U1889 (N_1889,N_1623,N_1656);
nand U1890 (N_1890,N_1653,N_1734);
nand U1891 (N_1891,N_1620,N_1692);
and U1892 (N_1892,N_1793,N_1639);
or U1893 (N_1893,N_1683,N_1613);
or U1894 (N_1894,N_1651,N_1667);
or U1895 (N_1895,N_1787,N_1685);
nand U1896 (N_1896,N_1609,N_1654);
nor U1897 (N_1897,N_1619,N_1663);
and U1898 (N_1898,N_1789,N_1795);
or U1899 (N_1899,N_1755,N_1766);
nand U1900 (N_1900,N_1613,N_1647);
nand U1901 (N_1901,N_1601,N_1606);
nor U1902 (N_1902,N_1643,N_1778);
nand U1903 (N_1903,N_1746,N_1682);
and U1904 (N_1904,N_1798,N_1678);
or U1905 (N_1905,N_1740,N_1701);
or U1906 (N_1906,N_1642,N_1710);
or U1907 (N_1907,N_1738,N_1717);
or U1908 (N_1908,N_1693,N_1703);
nand U1909 (N_1909,N_1787,N_1660);
and U1910 (N_1910,N_1645,N_1633);
or U1911 (N_1911,N_1679,N_1696);
or U1912 (N_1912,N_1731,N_1715);
and U1913 (N_1913,N_1761,N_1747);
or U1914 (N_1914,N_1666,N_1761);
nor U1915 (N_1915,N_1633,N_1639);
and U1916 (N_1916,N_1682,N_1736);
and U1917 (N_1917,N_1787,N_1669);
nand U1918 (N_1918,N_1709,N_1641);
or U1919 (N_1919,N_1798,N_1683);
and U1920 (N_1920,N_1712,N_1612);
nor U1921 (N_1921,N_1783,N_1707);
xnor U1922 (N_1922,N_1783,N_1650);
and U1923 (N_1923,N_1796,N_1642);
nand U1924 (N_1924,N_1695,N_1632);
nor U1925 (N_1925,N_1622,N_1695);
nand U1926 (N_1926,N_1771,N_1746);
nand U1927 (N_1927,N_1611,N_1700);
nand U1928 (N_1928,N_1753,N_1734);
nor U1929 (N_1929,N_1687,N_1648);
or U1930 (N_1930,N_1740,N_1736);
or U1931 (N_1931,N_1752,N_1793);
nand U1932 (N_1932,N_1753,N_1714);
nor U1933 (N_1933,N_1678,N_1696);
or U1934 (N_1934,N_1662,N_1695);
nand U1935 (N_1935,N_1675,N_1614);
or U1936 (N_1936,N_1639,N_1794);
xor U1937 (N_1937,N_1686,N_1781);
nor U1938 (N_1938,N_1739,N_1784);
nand U1939 (N_1939,N_1671,N_1686);
and U1940 (N_1940,N_1793,N_1612);
or U1941 (N_1941,N_1759,N_1618);
or U1942 (N_1942,N_1783,N_1675);
nor U1943 (N_1943,N_1647,N_1697);
nand U1944 (N_1944,N_1750,N_1632);
and U1945 (N_1945,N_1653,N_1776);
nand U1946 (N_1946,N_1660,N_1641);
nor U1947 (N_1947,N_1611,N_1723);
nand U1948 (N_1948,N_1799,N_1698);
xnor U1949 (N_1949,N_1670,N_1674);
nor U1950 (N_1950,N_1656,N_1798);
and U1951 (N_1951,N_1688,N_1622);
nor U1952 (N_1952,N_1741,N_1744);
xnor U1953 (N_1953,N_1693,N_1637);
nor U1954 (N_1954,N_1680,N_1648);
xnor U1955 (N_1955,N_1663,N_1680);
xnor U1956 (N_1956,N_1668,N_1700);
or U1957 (N_1957,N_1651,N_1718);
nand U1958 (N_1958,N_1699,N_1664);
or U1959 (N_1959,N_1620,N_1742);
or U1960 (N_1960,N_1793,N_1655);
nor U1961 (N_1961,N_1772,N_1630);
or U1962 (N_1962,N_1687,N_1754);
nand U1963 (N_1963,N_1741,N_1754);
or U1964 (N_1964,N_1645,N_1690);
xnor U1965 (N_1965,N_1795,N_1603);
nor U1966 (N_1966,N_1624,N_1617);
nand U1967 (N_1967,N_1664,N_1668);
xor U1968 (N_1968,N_1773,N_1769);
xor U1969 (N_1969,N_1624,N_1681);
xor U1970 (N_1970,N_1611,N_1648);
nand U1971 (N_1971,N_1702,N_1699);
and U1972 (N_1972,N_1758,N_1731);
or U1973 (N_1973,N_1615,N_1735);
nor U1974 (N_1974,N_1769,N_1605);
nor U1975 (N_1975,N_1600,N_1687);
nor U1976 (N_1976,N_1685,N_1707);
nand U1977 (N_1977,N_1752,N_1651);
nand U1978 (N_1978,N_1680,N_1600);
nor U1979 (N_1979,N_1633,N_1713);
or U1980 (N_1980,N_1741,N_1703);
and U1981 (N_1981,N_1689,N_1614);
or U1982 (N_1982,N_1713,N_1705);
nand U1983 (N_1983,N_1605,N_1669);
or U1984 (N_1984,N_1751,N_1706);
and U1985 (N_1985,N_1753,N_1603);
nor U1986 (N_1986,N_1706,N_1795);
nor U1987 (N_1987,N_1600,N_1632);
or U1988 (N_1988,N_1668,N_1714);
nor U1989 (N_1989,N_1749,N_1770);
or U1990 (N_1990,N_1771,N_1739);
or U1991 (N_1991,N_1606,N_1719);
or U1992 (N_1992,N_1739,N_1787);
or U1993 (N_1993,N_1644,N_1616);
or U1994 (N_1994,N_1677,N_1608);
or U1995 (N_1995,N_1681,N_1788);
or U1996 (N_1996,N_1770,N_1649);
and U1997 (N_1997,N_1724,N_1770);
or U1998 (N_1998,N_1656,N_1653);
and U1999 (N_1999,N_1672,N_1730);
nand U2000 (N_2000,N_1856,N_1929);
nand U2001 (N_2001,N_1928,N_1802);
xnor U2002 (N_2002,N_1917,N_1860);
or U2003 (N_2003,N_1813,N_1957);
nor U2004 (N_2004,N_1948,N_1939);
xor U2005 (N_2005,N_1967,N_1958);
or U2006 (N_2006,N_1830,N_1940);
and U2007 (N_2007,N_1851,N_1991);
and U2008 (N_2008,N_1823,N_1885);
nand U2009 (N_2009,N_1960,N_1808);
nor U2010 (N_2010,N_1945,N_1911);
nor U2011 (N_2011,N_1882,N_1873);
nand U2012 (N_2012,N_1903,N_1867);
nand U2013 (N_2013,N_1891,N_1861);
and U2014 (N_2014,N_1952,N_1923);
and U2015 (N_2015,N_1820,N_1838);
or U2016 (N_2016,N_1825,N_1970);
nand U2017 (N_2017,N_1998,N_1919);
and U2018 (N_2018,N_1961,N_1826);
nor U2019 (N_2019,N_1857,N_1978);
nor U2020 (N_2020,N_1976,N_1890);
and U2021 (N_2021,N_1966,N_1990);
nor U2022 (N_2022,N_1827,N_1997);
xor U2023 (N_2023,N_1931,N_1921);
nand U2024 (N_2024,N_1979,N_1992);
nand U2025 (N_2025,N_1924,N_1804);
nand U2026 (N_2026,N_1853,N_1995);
or U2027 (N_2027,N_1902,N_1855);
or U2028 (N_2028,N_1810,N_1892);
nor U2029 (N_2029,N_1932,N_1816);
or U2030 (N_2030,N_1974,N_1878);
or U2031 (N_2031,N_1847,N_1844);
nor U2032 (N_2032,N_1865,N_1800);
nand U2033 (N_2033,N_1982,N_1840);
nand U2034 (N_2034,N_1963,N_1984);
nor U2035 (N_2035,N_1941,N_1875);
nor U2036 (N_2036,N_1845,N_1905);
and U2037 (N_2037,N_1883,N_1812);
nand U2038 (N_2038,N_1811,N_1887);
xnor U2039 (N_2039,N_1869,N_1909);
and U2040 (N_2040,N_1834,N_1946);
and U2041 (N_2041,N_1950,N_1849);
nor U2042 (N_2042,N_1870,N_1968);
nand U2043 (N_2043,N_1988,N_1925);
and U2044 (N_2044,N_1858,N_1897);
nor U2045 (N_2045,N_1955,N_1951);
nand U2046 (N_2046,N_1837,N_1803);
nor U2047 (N_2047,N_1913,N_1895);
xor U2048 (N_2048,N_1972,N_1815);
and U2049 (N_2049,N_1859,N_1971);
and U2050 (N_2050,N_1912,N_1835);
or U2051 (N_2051,N_1836,N_1977);
and U2052 (N_2052,N_1936,N_1801);
xor U2053 (N_2053,N_1954,N_1818);
xor U2054 (N_2054,N_1985,N_1852);
nor U2055 (N_2055,N_1839,N_1888);
xnor U2056 (N_2056,N_1807,N_1898);
xnor U2057 (N_2057,N_1841,N_1994);
or U2058 (N_2058,N_1962,N_1908);
or U2059 (N_2059,N_1880,N_1822);
xor U2060 (N_2060,N_1894,N_1956);
nor U2061 (N_2061,N_1964,N_1876);
nand U2062 (N_2062,N_1805,N_1886);
xnor U2063 (N_2063,N_1863,N_1907);
and U2064 (N_2064,N_1874,N_1914);
nand U2065 (N_2065,N_1901,N_1893);
xnor U2066 (N_2066,N_1831,N_1983);
and U2067 (N_2067,N_1809,N_1942);
nor U2068 (N_2068,N_1934,N_1993);
xor U2069 (N_2069,N_1899,N_1949);
and U2070 (N_2070,N_1930,N_1922);
nand U2071 (N_2071,N_1848,N_1937);
and U2072 (N_2072,N_1889,N_1969);
nand U2073 (N_2073,N_1904,N_1829);
xor U2074 (N_2074,N_1866,N_1871);
and U2075 (N_2075,N_1935,N_1806);
or U2076 (N_2076,N_1943,N_1959);
nor U2077 (N_2077,N_1900,N_1918);
or U2078 (N_2078,N_1965,N_1864);
nor U2079 (N_2079,N_1833,N_1842);
xnor U2080 (N_2080,N_1846,N_1896);
or U2081 (N_2081,N_1879,N_1915);
xor U2082 (N_2082,N_1884,N_1916);
and U2083 (N_2083,N_1927,N_1980);
xor U2084 (N_2084,N_1987,N_1920);
nand U2085 (N_2085,N_1843,N_1989);
xnor U2086 (N_2086,N_1819,N_1906);
xnor U2087 (N_2087,N_1975,N_1850);
nor U2088 (N_2088,N_1824,N_1973);
and U2089 (N_2089,N_1926,N_1933);
or U2090 (N_2090,N_1868,N_1862);
or U2091 (N_2091,N_1832,N_1996);
nand U2092 (N_2092,N_1877,N_1817);
xor U2093 (N_2093,N_1981,N_1814);
and U2094 (N_2094,N_1944,N_1910);
nor U2095 (N_2095,N_1938,N_1986);
or U2096 (N_2096,N_1828,N_1953);
nor U2097 (N_2097,N_1947,N_1881);
and U2098 (N_2098,N_1872,N_1854);
nand U2099 (N_2099,N_1999,N_1821);
or U2100 (N_2100,N_1928,N_1888);
xnor U2101 (N_2101,N_1922,N_1979);
or U2102 (N_2102,N_1969,N_1832);
xor U2103 (N_2103,N_1977,N_1949);
nand U2104 (N_2104,N_1841,N_1982);
xor U2105 (N_2105,N_1971,N_1957);
xnor U2106 (N_2106,N_1807,N_1809);
and U2107 (N_2107,N_1877,N_1816);
nand U2108 (N_2108,N_1850,N_1875);
or U2109 (N_2109,N_1843,N_1833);
nand U2110 (N_2110,N_1976,N_1936);
and U2111 (N_2111,N_1892,N_1903);
or U2112 (N_2112,N_1842,N_1885);
or U2113 (N_2113,N_1961,N_1893);
or U2114 (N_2114,N_1947,N_1902);
and U2115 (N_2115,N_1859,N_1978);
or U2116 (N_2116,N_1847,N_1858);
and U2117 (N_2117,N_1880,N_1808);
or U2118 (N_2118,N_1813,N_1853);
and U2119 (N_2119,N_1824,N_1985);
nand U2120 (N_2120,N_1827,N_1941);
or U2121 (N_2121,N_1817,N_1828);
or U2122 (N_2122,N_1922,N_1957);
nor U2123 (N_2123,N_1868,N_1957);
xor U2124 (N_2124,N_1967,N_1846);
and U2125 (N_2125,N_1999,N_1938);
nand U2126 (N_2126,N_1874,N_1958);
nor U2127 (N_2127,N_1860,N_1896);
or U2128 (N_2128,N_1815,N_1960);
and U2129 (N_2129,N_1886,N_1939);
and U2130 (N_2130,N_1905,N_1997);
nor U2131 (N_2131,N_1938,N_1975);
nor U2132 (N_2132,N_1892,N_1924);
xnor U2133 (N_2133,N_1933,N_1989);
or U2134 (N_2134,N_1998,N_1921);
nor U2135 (N_2135,N_1983,N_1905);
xor U2136 (N_2136,N_1885,N_1994);
nand U2137 (N_2137,N_1841,N_1950);
nand U2138 (N_2138,N_1968,N_1868);
or U2139 (N_2139,N_1911,N_1889);
and U2140 (N_2140,N_1943,N_1926);
or U2141 (N_2141,N_1976,N_1993);
nand U2142 (N_2142,N_1870,N_1924);
nor U2143 (N_2143,N_1875,N_1903);
nor U2144 (N_2144,N_1907,N_1830);
nand U2145 (N_2145,N_1904,N_1937);
or U2146 (N_2146,N_1885,N_1926);
and U2147 (N_2147,N_1920,N_1854);
nor U2148 (N_2148,N_1830,N_1816);
nor U2149 (N_2149,N_1983,N_1898);
or U2150 (N_2150,N_1967,N_1968);
and U2151 (N_2151,N_1874,N_1919);
nor U2152 (N_2152,N_1866,N_1839);
and U2153 (N_2153,N_1905,N_1808);
nand U2154 (N_2154,N_1882,N_1819);
and U2155 (N_2155,N_1880,N_1891);
or U2156 (N_2156,N_1994,N_1955);
and U2157 (N_2157,N_1965,N_1962);
xor U2158 (N_2158,N_1911,N_1873);
xor U2159 (N_2159,N_1825,N_1901);
and U2160 (N_2160,N_1921,N_1929);
or U2161 (N_2161,N_1914,N_1877);
nand U2162 (N_2162,N_1865,N_1948);
xnor U2163 (N_2163,N_1852,N_1811);
nor U2164 (N_2164,N_1945,N_1986);
nor U2165 (N_2165,N_1861,N_1905);
nand U2166 (N_2166,N_1831,N_1968);
and U2167 (N_2167,N_1834,N_1843);
xor U2168 (N_2168,N_1835,N_1869);
nor U2169 (N_2169,N_1875,N_1854);
or U2170 (N_2170,N_1802,N_1988);
or U2171 (N_2171,N_1895,N_1921);
nand U2172 (N_2172,N_1959,N_1877);
xnor U2173 (N_2173,N_1872,N_1847);
and U2174 (N_2174,N_1891,N_1842);
nand U2175 (N_2175,N_1879,N_1802);
nand U2176 (N_2176,N_1941,N_1959);
or U2177 (N_2177,N_1881,N_1904);
nor U2178 (N_2178,N_1996,N_1936);
or U2179 (N_2179,N_1909,N_1867);
xor U2180 (N_2180,N_1978,N_1954);
nor U2181 (N_2181,N_1998,N_1800);
and U2182 (N_2182,N_1898,N_1818);
xnor U2183 (N_2183,N_1952,N_1912);
or U2184 (N_2184,N_1826,N_1882);
nor U2185 (N_2185,N_1914,N_1876);
or U2186 (N_2186,N_1925,N_1951);
nor U2187 (N_2187,N_1830,N_1984);
xnor U2188 (N_2188,N_1955,N_1869);
nor U2189 (N_2189,N_1846,N_1806);
and U2190 (N_2190,N_1868,N_1814);
xnor U2191 (N_2191,N_1999,N_1937);
xnor U2192 (N_2192,N_1904,N_1965);
nand U2193 (N_2193,N_1892,N_1935);
xor U2194 (N_2194,N_1854,N_1912);
nand U2195 (N_2195,N_1912,N_1838);
and U2196 (N_2196,N_1851,N_1973);
nor U2197 (N_2197,N_1829,N_1822);
and U2198 (N_2198,N_1938,N_1853);
and U2199 (N_2199,N_1865,N_1854);
nor U2200 (N_2200,N_2122,N_2109);
nor U2201 (N_2201,N_2084,N_2181);
nor U2202 (N_2202,N_2119,N_2150);
nor U2203 (N_2203,N_2158,N_2094);
or U2204 (N_2204,N_2170,N_2117);
nor U2205 (N_2205,N_2161,N_2176);
xor U2206 (N_2206,N_2155,N_2057);
nor U2207 (N_2207,N_2187,N_2003);
nor U2208 (N_2208,N_2001,N_2036);
xor U2209 (N_2209,N_2163,N_2103);
and U2210 (N_2210,N_2125,N_2016);
xnor U2211 (N_2211,N_2090,N_2083);
nand U2212 (N_2212,N_2132,N_2086);
nand U2213 (N_2213,N_2139,N_2008);
or U2214 (N_2214,N_2178,N_2006);
and U2215 (N_2215,N_2040,N_2118);
and U2216 (N_2216,N_2157,N_2093);
xnor U2217 (N_2217,N_2049,N_2110);
nand U2218 (N_2218,N_2112,N_2046);
and U2219 (N_2219,N_2026,N_2194);
or U2220 (N_2220,N_2153,N_2022);
and U2221 (N_2221,N_2072,N_2114);
or U2222 (N_2222,N_2159,N_2149);
xnor U2223 (N_2223,N_2073,N_2120);
xor U2224 (N_2224,N_2175,N_2104);
nor U2225 (N_2225,N_2140,N_2146);
nand U2226 (N_2226,N_2031,N_2071);
nor U2227 (N_2227,N_2043,N_2076);
or U2228 (N_2228,N_2052,N_2018);
xor U2229 (N_2229,N_2130,N_2169);
xnor U2230 (N_2230,N_2033,N_2079);
nor U2231 (N_2231,N_2065,N_2037);
nor U2232 (N_2232,N_2095,N_2106);
xor U2233 (N_2233,N_2053,N_2180);
or U2234 (N_2234,N_2188,N_2190);
or U2235 (N_2235,N_2099,N_2168);
or U2236 (N_2236,N_2183,N_2074);
or U2237 (N_2237,N_2034,N_2056);
or U2238 (N_2238,N_2167,N_2010);
and U2239 (N_2239,N_2038,N_2129);
xnor U2240 (N_2240,N_2151,N_2013);
nor U2241 (N_2241,N_2024,N_2067);
nand U2242 (N_2242,N_2039,N_2060);
xnor U2243 (N_2243,N_2032,N_2023);
nor U2244 (N_2244,N_2126,N_2124);
nor U2245 (N_2245,N_2198,N_2135);
and U2246 (N_2246,N_2195,N_2004);
nand U2247 (N_2247,N_2047,N_2179);
nor U2248 (N_2248,N_2171,N_2091);
xor U2249 (N_2249,N_2160,N_2045);
xor U2250 (N_2250,N_2154,N_2182);
and U2251 (N_2251,N_2185,N_2141);
and U2252 (N_2252,N_2152,N_2044);
or U2253 (N_2253,N_2005,N_2051);
nand U2254 (N_2254,N_2059,N_2189);
nor U2255 (N_2255,N_2142,N_2148);
or U2256 (N_2256,N_2029,N_2173);
nand U2257 (N_2257,N_2098,N_2042);
nor U2258 (N_2258,N_2105,N_2102);
or U2259 (N_2259,N_2144,N_2111);
xor U2260 (N_2260,N_2156,N_2002);
xnor U2261 (N_2261,N_2186,N_2066);
and U2262 (N_2262,N_2162,N_2075);
or U2263 (N_2263,N_2035,N_2192);
nand U2264 (N_2264,N_2021,N_2070);
or U2265 (N_2265,N_2143,N_2041);
and U2266 (N_2266,N_2089,N_2048);
nor U2267 (N_2267,N_2115,N_2080);
nand U2268 (N_2268,N_2197,N_2088);
and U2269 (N_2269,N_2009,N_2134);
and U2270 (N_2270,N_2131,N_2191);
nand U2271 (N_2271,N_2078,N_2165);
nor U2272 (N_2272,N_2127,N_2121);
xnor U2273 (N_2273,N_2087,N_2054);
nand U2274 (N_2274,N_2164,N_2014);
xor U2275 (N_2275,N_2017,N_2123);
xnor U2276 (N_2276,N_2113,N_2068);
or U2277 (N_2277,N_2199,N_2020);
nand U2278 (N_2278,N_2145,N_2172);
xnor U2279 (N_2279,N_2108,N_2092);
nand U2280 (N_2280,N_2166,N_2136);
nand U2281 (N_2281,N_2027,N_2055);
nor U2282 (N_2282,N_2107,N_2050);
and U2283 (N_2283,N_2184,N_2063);
nor U2284 (N_2284,N_2147,N_2082);
xnor U2285 (N_2285,N_2064,N_2096);
nand U2286 (N_2286,N_2019,N_2077);
xnor U2287 (N_2287,N_2012,N_2028);
or U2288 (N_2288,N_2138,N_2025);
or U2289 (N_2289,N_2177,N_2116);
xor U2290 (N_2290,N_2174,N_2133);
or U2291 (N_2291,N_2011,N_2061);
or U2292 (N_2292,N_2193,N_2081);
or U2293 (N_2293,N_2030,N_2015);
nor U2294 (N_2294,N_2058,N_2007);
and U2295 (N_2295,N_2000,N_2196);
and U2296 (N_2296,N_2128,N_2137);
and U2297 (N_2297,N_2069,N_2100);
xnor U2298 (N_2298,N_2062,N_2101);
or U2299 (N_2299,N_2097,N_2085);
nand U2300 (N_2300,N_2043,N_2168);
or U2301 (N_2301,N_2100,N_2115);
xor U2302 (N_2302,N_2179,N_2081);
and U2303 (N_2303,N_2194,N_2085);
xor U2304 (N_2304,N_2097,N_2176);
or U2305 (N_2305,N_2001,N_2108);
xor U2306 (N_2306,N_2088,N_2067);
xnor U2307 (N_2307,N_2029,N_2121);
xor U2308 (N_2308,N_2148,N_2167);
nand U2309 (N_2309,N_2135,N_2103);
nor U2310 (N_2310,N_2041,N_2116);
or U2311 (N_2311,N_2046,N_2014);
nor U2312 (N_2312,N_2044,N_2145);
or U2313 (N_2313,N_2080,N_2155);
and U2314 (N_2314,N_2068,N_2098);
nand U2315 (N_2315,N_2055,N_2079);
xnor U2316 (N_2316,N_2172,N_2011);
or U2317 (N_2317,N_2055,N_2182);
xor U2318 (N_2318,N_2169,N_2004);
nand U2319 (N_2319,N_2126,N_2051);
nand U2320 (N_2320,N_2093,N_2061);
xor U2321 (N_2321,N_2027,N_2093);
nand U2322 (N_2322,N_2105,N_2008);
xnor U2323 (N_2323,N_2149,N_2035);
and U2324 (N_2324,N_2166,N_2190);
nand U2325 (N_2325,N_2179,N_2045);
or U2326 (N_2326,N_2060,N_2038);
nor U2327 (N_2327,N_2167,N_2184);
and U2328 (N_2328,N_2164,N_2082);
or U2329 (N_2329,N_2125,N_2168);
xnor U2330 (N_2330,N_2052,N_2031);
and U2331 (N_2331,N_2150,N_2087);
and U2332 (N_2332,N_2154,N_2198);
nor U2333 (N_2333,N_2121,N_2140);
xnor U2334 (N_2334,N_2159,N_2164);
and U2335 (N_2335,N_2023,N_2095);
nand U2336 (N_2336,N_2087,N_2069);
xnor U2337 (N_2337,N_2163,N_2083);
nand U2338 (N_2338,N_2046,N_2015);
nand U2339 (N_2339,N_2190,N_2081);
nor U2340 (N_2340,N_2141,N_2010);
xor U2341 (N_2341,N_2149,N_2185);
and U2342 (N_2342,N_2019,N_2025);
nand U2343 (N_2343,N_2034,N_2164);
nor U2344 (N_2344,N_2030,N_2174);
xnor U2345 (N_2345,N_2138,N_2071);
nand U2346 (N_2346,N_2078,N_2068);
nand U2347 (N_2347,N_2025,N_2128);
or U2348 (N_2348,N_2123,N_2082);
or U2349 (N_2349,N_2188,N_2191);
and U2350 (N_2350,N_2065,N_2146);
or U2351 (N_2351,N_2010,N_2011);
nand U2352 (N_2352,N_2099,N_2174);
nor U2353 (N_2353,N_2112,N_2135);
nand U2354 (N_2354,N_2162,N_2019);
and U2355 (N_2355,N_2027,N_2061);
nand U2356 (N_2356,N_2199,N_2065);
or U2357 (N_2357,N_2117,N_2144);
and U2358 (N_2358,N_2007,N_2026);
or U2359 (N_2359,N_2102,N_2029);
nor U2360 (N_2360,N_2028,N_2010);
xor U2361 (N_2361,N_2078,N_2199);
or U2362 (N_2362,N_2036,N_2197);
nand U2363 (N_2363,N_2176,N_2109);
xnor U2364 (N_2364,N_2002,N_2143);
and U2365 (N_2365,N_2025,N_2095);
and U2366 (N_2366,N_2037,N_2085);
nor U2367 (N_2367,N_2175,N_2036);
nand U2368 (N_2368,N_2075,N_2181);
or U2369 (N_2369,N_2102,N_2065);
nand U2370 (N_2370,N_2158,N_2033);
xnor U2371 (N_2371,N_2197,N_2186);
or U2372 (N_2372,N_2029,N_2000);
or U2373 (N_2373,N_2162,N_2155);
nor U2374 (N_2374,N_2114,N_2161);
xnor U2375 (N_2375,N_2104,N_2076);
nand U2376 (N_2376,N_2136,N_2151);
nor U2377 (N_2377,N_2097,N_2161);
or U2378 (N_2378,N_2191,N_2092);
or U2379 (N_2379,N_2150,N_2070);
or U2380 (N_2380,N_2196,N_2169);
xor U2381 (N_2381,N_2017,N_2020);
and U2382 (N_2382,N_2068,N_2058);
nand U2383 (N_2383,N_2114,N_2041);
or U2384 (N_2384,N_2119,N_2040);
nand U2385 (N_2385,N_2168,N_2069);
and U2386 (N_2386,N_2038,N_2020);
or U2387 (N_2387,N_2148,N_2004);
and U2388 (N_2388,N_2160,N_2102);
nor U2389 (N_2389,N_2175,N_2183);
and U2390 (N_2390,N_2175,N_2162);
and U2391 (N_2391,N_2193,N_2087);
and U2392 (N_2392,N_2003,N_2008);
xor U2393 (N_2393,N_2189,N_2007);
nor U2394 (N_2394,N_2014,N_2036);
xnor U2395 (N_2395,N_2027,N_2010);
and U2396 (N_2396,N_2072,N_2100);
nor U2397 (N_2397,N_2102,N_2190);
or U2398 (N_2398,N_2084,N_2039);
or U2399 (N_2399,N_2001,N_2041);
nor U2400 (N_2400,N_2264,N_2272);
and U2401 (N_2401,N_2365,N_2302);
or U2402 (N_2402,N_2243,N_2318);
nand U2403 (N_2403,N_2290,N_2269);
or U2404 (N_2404,N_2330,N_2287);
and U2405 (N_2405,N_2210,N_2329);
nand U2406 (N_2406,N_2308,N_2256);
nor U2407 (N_2407,N_2212,N_2366);
nand U2408 (N_2408,N_2320,N_2386);
nor U2409 (N_2409,N_2231,N_2216);
nand U2410 (N_2410,N_2339,N_2217);
and U2411 (N_2411,N_2208,N_2346);
nor U2412 (N_2412,N_2313,N_2332);
and U2413 (N_2413,N_2393,N_2340);
nand U2414 (N_2414,N_2286,N_2224);
or U2415 (N_2415,N_2271,N_2301);
or U2416 (N_2416,N_2259,N_2277);
or U2417 (N_2417,N_2295,N_2384);
xnor U2418 (N_2418,N_2334,N_2294);
nand U2419 (N_2419,N_2336,N_2250);
xor U2420 (N_2420,N_2267,N_2317);
nor U2421 (N_2421,N_2283,N_2222);
nor U2422 (N_2422,N_2394,N_2335);
xnor U2423 (N_2423,N_2344,N_2253);
and U2424 (N_2424,N_2363,N_2281);
and U2425 (N_2425,N_2296,N_2205);
nand U2426 (N_2426,N_2331,N_2399);
and U2427 (N_2427,N_2280,N_2227);
and U2428 (N_2428,N_2263,N_2323);
nand U2429 (N_2429,N_2390,N_2225);
nor U2430 (N_2430,N_2369,N_2378);
nor U2431 (N_2431,N_2388,N_2273);
nand U2432 (N_2432,N_2262,N_2315);
nand U2433 (N_2433,N_2252,N_2314);
nor U2434 (N_2434,N_2300,N_2348);
xor U2435 (N_2435,N_2357,N_2321);
nand U2436 (N_2436,N_2345,N_2247);
nor U2437 (N_2437,N_2333,N_2209);
nand U2438 (N_2438,N_2355,N_2228);
nand U2439 (N_2439,N_2245,N_2239);
or U2440 (N_2440,N_2251,N_2299);
nand U2441 (N_2441,N_2398,N_2254);
xnor U2442 (N_2442,N_2235,N_2322);
and U2443 (N_2443,N_2337,N_2350);
and U2444 (N_2444,N_2328,N_2376);
nor U2445 (N_2445,N_2229,N_2242);
and U2446 (N_2446,N_2391,N_2289);
and U2447 (N_2447,N_2358,N_2232);
or U2448 (N_2448,N_2327,N_2375);
or U2449 (N_2449,N_2237,N_2361);
or U2450 (N_2450,N_2260,N_2324);
nand U2451 (N_2451,N_2382,N_2213);
nand U2452 (N_2452,N_2354,N_2219);
nand U2453 (N_2453,N_2373,N_2265);
xor U2454 (N_2454,N_2274,N_2293);
and U2455 (N_2455,N_2367,N_2288);
or U2456 (N_2456,N_2372,N_2352);
nand U2457 (N_2457,N_2223,N_2364);
or U2458 (N_2458,N_2220,N_2349);
or U2459 (N_2459,N_2310,N_2215);
and U2460 (N_2460,N_2207,N_2309);
or U2461 (N_2461,N_2374,N_2279);
nor U2462 (N_2462,N_2278,N_2284);
nand U2463 (N_2463,N_2204,N_2285);
nand U2464 (N_2464,N_2351,N_2396);
nor U2465 (N_2465,N_2203,N_2246);
and U2466 (N_2466,N_2275,N_2240);
or U2467 (N_2467,N_2362,N_2206);
nor U2468 (N_2468,N_2257,N_2325);
nand U2469 (N_2469,N_2266,N_2241);
nand U2470 (N_2470,N_2291,N_2201);
or U2471 (N_2471,N_2236,N_2311);
nor U2472 (N_2472,N_2326,N_2233);
nand U2473 (N_2473,N_2297,N_2395);
nand U2474 (N_2474,N_2316,N_2381);
xor U2475 (N_2475,N_2214,N_2276);
nor U2476 (N_2476,N_2303,N_2249);
nor U2477 (N_2477,N_2338,N_2255);
or U2478 (N_2478,N_2200,N_2305);
and U2479 (N_2479,N_2379,N_2377);
nand U2480 (N_2480,N_2226,N_2202);
or U2481 (N_2481,N_2298,N_2307);
and U2482 (N_2482,N_2234,N_2383);
nor U2483 (N_2483,N_2270,N_2221);
xnor U2484 (N_2484,N_2343,N_2258);
nand U2485 (N_2485,N_2268,N_2282);
nand U2486 (N_2486,N_2370,N_2371);
xnor U2487 (N_2487,N_2261,N_2218);
xor U2488 (N_2488,N_2387,N_2342);
xnor U2489 (N_2489,N_2359,N_2385);
and U2490 (N_2490,N_2360,N_2248);
xnor U2491 (N_2491,N_2392,N_2356);
nand U2492 (N_2492,N_2347,N_2389);
and U2493 (N_2493,N_2238,N_2244);
and U2494 (N_2494,N_2292,N_2397);
nor U2495 (N_2495,N_2304,N_2319);
nor U2496 (N_2496,N_2380,N_2341);
xnor U2497 (N_2497,N_2230,N_2353);
or U2498 (N_2498,N_2306,N_2312);
or U2499 (N_2499,N_2368,N_2211);
and U2500 (N_2500,N_2320,N_2219);
nor U2501 (N_2501,N_2335,N_2333);
nor U2502 (N_2502,N_2377,N_2333);
nor U2503 (N_2503,N_2223,N_2354);
or U2504 (N_2504,N_2220,N_2213);
or U2505 (N_2505,N_2285,N_2221);
or U2506 (N_2506,N_2356,N_2224);
xor U2507 (N_2507,N_2390,N_2322);
or U2508 (N_2508,N_2336,N_2260);
or U2509 (N_2509,N_2385,N_2288);
xnor U2510 (N_2510,N_2215,N_2394);
nand U2511 (N_2511,N_2231,N_2296);
nand U2512 (N_2512,N_2247,N_2279);
xor U2513 (N_2513,N_2249,N_2229);
xor U2514 (N_2514,N_2215,N_2365);
and U2515 (N_2515,N_2368,N_2261);
nand U2516 (N_2516,N_2243,N_2398);
and U2517 (N_2517,N_2279,N_2253);
and U2518 (N_2518,N_2224,N_2223);
xor U2519 (N_2519,N_2374,N_2222);
nand U2520 (N_2520,N_2311,N_2256);
or U2521 (N_2521,N_2340,N_2254);
or U2522 (N_2522,N_2235,N_2333);
nand U2523 (N_2523,N_2206,N_2319);
and U2524 (N_2524,N_2240,N_2373);
nor U2525 (N_2525,N_2368,N_2326);
nand U2526 (N_2526,N_2224,N_2387);
and U2527 (N_2527,N_2205,N_2369);
nand U2528 (N_2528,N_2329,N_2336);
nor U2529 (N_2529,N_2304,N_2338);
nor U2530 (N_2530,N_2331,N_2251);
or U2531 (N_2531,N_2264,N_2394);
or U2532 (N_2532,N_2202,N_2371);
and U2533 (N_2533,N_2273,N_2367);
or U2534 (N_2534,N_2317,N_2324);
and U2535 (N_2535,N_2299,N_2376);
nor U2536 (N_2536,N_2375,N_2305);
xnor U2537 (N_2537,N_2327,N_2207);
xor U2538 (N_2538,N_2316,N_2322);
and U2539 (N_2539,N_2341,N_2279);
nand U2540 (N_2540,N_2236,N_2278);
nand U2541 (N_2541,N_2272,N_2310);
nor U2542 (N_2542,N_2343,N_2363);
nand U2543 (N_2543,N_2361,N_2239);
nor U2544 (N_2544,N_2242,N_2393);
or U2545 (N_2545,N_2333,N_2325);
and U2546 (N_2546,N_2388,N_2243);
and U2547 (N_2547,N_2340,N_2217);
or U2548 (N_2548,N_2361,N_2211);
and U2549 (N_2549,N_2202,N_2300);
and U2550 (N_2550,N_2338,N_2286);
and U2551 (N_2551,N_2267,N_2333);
nor U2552 (N_2552,N_2217,N_2232);
xnor U2553 (N_2553,N_2257,N_2391);
nor U2554 (N_2554,N_2246,N_2394);
or U2555 (N_2555,N_2364,N_2320);
or U2556 (N_2556,N_2268,N_2249);
and U2557 (N_2557,N_2359,N_2270);
and U2558 (N_2558,N_2306,N_2292);
nand U2559 (N_2559,N_2202,N_2246);
and U2560 (N_2560,N_2334,N_2218);
nand U2561 (N_2561,N_2393,N_2354);
or U2562 (N_2562,N_2297,N_2373);
nand U2563 (N_2563,N_2395,N_2372);
xnor U2564 (N_2564,N_2319,N_2208);
and U2565 (N_2565,N_2385,N_2388);
xor U2566 (N_2566,N_2215,N_2348);
nand U2567 (N_2567,N_2270,N_2237);
nand U2568 (N_2568,N_2245,N_2367);
xor U2569 (N_2569,N_2363,N_2242);
or U2570 (N_2570,N_2340,N_2284);
nor U2571 (N_2571,N_2253,N_2273);
or U2572 (N_2572,N_2247,N_2384);
and U2573 (N_2573,N_2329,N_2218);
and U2574 (N_2574,N_2256,N_2260);
xor U2575 (N_2575,N_2285,N_2283);
nand U2576 (N_2576,N_2332,N_2319);
or U2577 (N_2577,N_2251,N_2212);
xnor U2578 (N_2578,N_2232,N_2285);
and U2579 (N_2579,N_2378,N_2360);
xnor U2580 (N_2580,N_2262,N_2225);
nor U2581 (N_2581,N_2329,N_2300);
nor U2582 (N_2582,N_2311,N_2228);
nand U2583 (N_2583,N_2252,N_2290);
nand U2584 (N_2584,N_2308,N_2210);
xnor U2585 (N_2585,N_2319,N_2378);
or U2586 (N_2586,N_2208,N_2222);
nand U2587 (N_2587,N_2356,N_2380);
nand U2588 (N_2588,N_2214,N_2290);
or U2589 (N_2589,N_2384,N_2373);
xor U2590 (N_2590,N_2307,N_2283);
nand U2591 (N_2591,N_2394,N_2237);
nand U2592 (N_2592,N_2216,N_2233);
nand U2593 (N_2593,N_2303,N_2324);
nand U2594 (N_2594,N_2357,N_2212);
or U2595 (N_2595,N_2347,N_2330);
or U2596 (N_2596,N_2216,N_2264);
and U2597 (N_2597,N_2284,N_2367);
nor U2598 (N_2598,N_2277,N_2223);
or U2599 (N_2599,N_2227,N_2338);
nor U2600 (N_2600,N_2453,N_2505);
and U2601 (N_2601,N_2474,N_2443);
or U2602 (N_2602,N_2492,N_2510);
nand U2603 (N_2603,N_2403,N_2545);
and U2604 (N_2604,N_2495,N_2573);
xor U2605 (N_2605,N_2419,N_2460);
and U2606 (N_2606,N_2524,N_2559);
or U2607 (N_2607,N_2572,N_2449);
and U2608 (N_2608,N_2469,N_2409);
nand U2609 (N_2609,N_2480,N_2564);
xnor U2610 (N_2610,N_2478,N_2597);
nand U2611 (N_2611,N_2520,N_2535);
nand U2612 (N_2612,N_2570,N_2551);
or U2613 (N_2613,N_2549,N_2422);
and U2614 (N_2614,N_2404,N_2569);
xnor U2615 (N_2615,N_2499,N_2424);
or U2616 (N_2616,N_2596,N_2405);
xor U2617 (N_2617,N_2582,N_2482);
nand U2618 (N_2618,N_2555,N_2437);
nand U2619 (N_2619,N_2531,N_2455);
xor U2620 (N_2620,N_2457,N_2518);
or U2621 (N_2621,N_2546,N_2477);
and U2622 (N_2622,N_2500,N_2466);
nor U2623 (N_2623,N_2538,N_2463);
nand U2624 (N_2624,N_2542,N_2561);
or U2625 (N_2625,N_2446,N_2451);
xnor U2626 (N_2626,N_2454,N_2571);
nor U2627 (N_2627,N_2515,N_2441);
and U2628 (N_2628,N_2563,N_2503);
and U2629 (N_2629,N_2496,N_2498);
nand U2630 (N_2630,N_2523,N_2445);
nor U2631 (N_2631,N_2416,N_2593);
or U2632 (N_2632,N_2444,N_2565);
xor U2633 (N_2633,N_2588,N_2430);
xor U2634 (N_2634,N_2487,N_2586);
and U2635 (N_2635,N_2472,N_2526);
and U2636 (N_2636,N_2567,N_2591);
xnor U2637 (N_2637,N_2458,N_2556);
or U2638 (N_2638,N_2512,N_2506);
nor U2639 (N_2639,N_2576,N_2410);
nand U2640 (N_2640,N_2401,N_2544);
nand U2641 (N_2641,N_2516,N_2452);
nand U2642 (N_2642,N_2522,N_2429);
xor U2643 (N_2643,N_2461,N_2427);
xor U2644 (N_2644,N_2585,N_2552);
nand U2645 (N_2645,N_2468,N_2470);
xnor U2646 (N_2646,N_2558,N_2583);
or U2647 (N_2647,N_2511,N_2548);
nor U2648 (N_2648,N_2432,N_2581);
nand U2649 (N_2649,N_2434,N_2431);
and U2650 (N_2650,N_2473,N_2527);
xor U2651 (N_2651,N_2486,N_2528);
and U2652 (N_2652,N_2568,N_2465);
xor U2653 (N_2653,N_2436,N_2519);
xnor U2654 (N_2654,N_2536,N_2580);
or U2655 (N_2655,N_2464,N_2423);
xnor U2656 (N_2656,N_2442,N_2440);
nor U2657 (N_2657,N_2476,N_2598);
and U2658 (N_2658,N_2514,N_2507);
and U2659 (N_2659,N_2493,N_2533);
xnor U2660 (N_2660,N_2578,N_2584);
or U2661 (N_2661,N_2575,N_2537);
and U2662 (N_2662,N_2557,N_2553);
or U2663 (N_2663,N_2574,N_2554);
nor U2664 (N_2664,N_2543,N_2412);
xnor U2665 (N_2665,N_2566,N_2433);
xor U2666 (N_2666,N_2481,N_2428);
nor U2667 (N_2667,N_2489,N_2530);
or U2668 (N_2668,N_2456,N_2508);
or U2669 (N_2669,N_2501,N_2579);
and U2670 (N_2670,N_2550,N_2414);
xnor U2671 (N_2671,N_2491,N_2447);
nand U2672 (N_2672,N_2521,N_2594);
xnor U2673 (N_2673,N_2411,N_2539);
nand U2674 (N_2674,N_2599,N_2494);
or U2675 (N_2675,N_2459,N_2450);
nor U2676 (N_2676,N_2587,N_2438);
nor U2677 (N_2677,N_2407,N_2488);
or U2678 (N_2678,N_2483,N_2417);
or U2679 (N_2679,N_2534,N_2595);
xor U2680 (N_2680,N_2540,N_2418);
nor U2681 (N_2681,N_2406,N_2467);
xor U2682 (N_2682,N_2497,N_2562);
or U2683 (N_2683,N_2426,N_2425);
xnor U2684 (N_2684,N_2421,N_2517);
nand U2685 (N_2685,N_2547,N_2415);
nand U2686 (N_2686,N_2400,N_2509);
xor U2687 (N_2687,N_2435,N_2532);
nor U2688 (N_2688,N_2471,N_2402);
nand U2689 (N_2689,N_2560,N_2479);
nand U2690 (N_2690,N_2577,N_2408);
and U2691 (N_2691,N_2462,N_2504);
nor U2692 (N_2692,N_2485,N_2589);
or U2693 (N_2693,N_2439,N_2541);
or U2694 (N_2694,N_2490,N_2513);
and U2695 (N_2695,N_2592,N_2420);
or U2696 (N_2696,N_2525,N_2590);
nor U2697 (N_2697,N_2502,N_2413);
nand U2698 (N_2698,N_2484,N_2448);
or U2699 (N_2699,N_2475,N_2529);
xor U2700 (N_2700,N_2429,N_2509);
or U2701 (N_2701,N_2472,N_2594);
and U2702 (N_2702,N_2526,N_2507);
or U2703 (N_2703,N_2470,N_2568);
and U2704 (N_2704,N_2544,N_2551);
or U2705 (N_2705,N_2488,N_2434);
nor U2706 (N_2706,N_2468,N_2547);
and U2707 (N_2707,N_2472,N_2444);
nand U2708 (N_2708,N_2495,N_2411);
nor U2709 (N_2709,N_2459,N_2516);
nor U2710 (N_2710,N_2501,N_2421);
nor U2711 (N_2711,N_2564,N_2478);
xnor U2712 (N_2712,N_2401,N_2594);
nand U2713 (N_2713,N_2594,N_2450);
nand U2714 (N_2714,N_2483,N_2557);
and U2715 (N_2715,N_2450,N_2544);
or U2716 (N_2716,N_2520,N_2420);
and U2717 (N_2717,N_2587,N_2413);
and U2718 (N_2718,N_2520,N_2481);
nor U2719 (N_2719,N_2512,N_2598);
nand U2720 (N_2720,N_2459,N_2512);
xnor U2721 (N_2721,N_2501,N_2473);
nand U2722 (N_2722,N_2473,N_2444);
xor U2723 (N_2723,N_2405,N_2548);
nor U2724 (N_2724,N_2450,N_2409);
and U2725 (N_2725,N_2501,N_2534);
nor U2726 (N_2726,N_2514,N_2497);
and U2727 (N_2727,N_2429,N_2434);
and U2728 (N_2728,N_2582,N_2492);
nand U2729 (N_2729,N_2560,N_2423);
nor U2730 (N_2730,N_2534,N_2594);
and U2731 (N_2731,N_2474,N_2551);
nor U2732 (N_2732,N_2421,N_2457);
nand U2733 (N_2733,N_2526,N_2540);
xor U2734 (N_2734,N_2555,N_2424);
or U2735 (N_2735,N_2445,N_2475);
or U2736 (N_2736,N_2562,N_2526);
and U2737 (N_2737,N_2580,N_2456);
xnor U2738 (N_2738,N_2582,N_2462);
nand U2739 (N_2739,N_2515,N_2526);
and U2740 (N_2740,N_2447,N_2532);
nor U2741 (N_2741,N_2471,N_2475);
xor U2742 (N_2742,N_2574,N_2576);
or U2743 (N_2743,N_2587,N_2440);
nor U2744 (N_2744,N_2437,N_2520);
or U2745 (N_2745,N_2425,N_2457);
nor U2746 (N_2746,N_2575,N_2427);
or U2747 (N_2747,N_2422,N_2510);
xnor U2748 (N_2748,N_2518,N_2571);
nor U2749 (N_2749,N_2421,N_2416);
nand U2750 (N_2750,N_2402,N_2407);
or U2751 (N_2751,N_2469,N_2425);
xor U2752 (N_2752,N_2577,N_2555);
nor U2753 (N_2753,N_2486,N_2491);
and U2754 (N_2754,N_2487,N_2567);
xor U2755 (N_2755,N_2466,N_2485);
nand U2756 (N_2756,N_2568,N_2553);
or U2757 (N_2757,N_2565,N_2508);
or U2758 (N_2758,N_2462,N_2505);
nand U2759 (N_2759,N_2401,N_2443);
or U2760 (N_2760,N_2449,N_2476);
or U2761 (N_2761,N_2432,N_2591);
nand U2762 (N_2762,N_2448,N_2557);
xor U2763 (N_2763,N_2438,N_2460);
nor U2764 (N_2764,N_2503,N_2429);
xnor U2765 (N_2765,N_2499,N_2537);
and U2766 (N_2766,N_2560,N_2572);
nor U2767 (N_2767,N_2473,N_2541);
nor U2768 (N_2768,N_2408,N_2569);
xnor U2769 (N_2769,N_2481,N_2410);
nand U2770 (N_2770,N_2412,N_2535);
nand U2771 (N_2771,N_2492,N_2563);
xor U2772 (N_2772,N_2544,N_2516);
and U2773 (N_2773,N_2548,N_2567);
and U2774 (N_2774,N_2463,N_2464);
or U2775 (N_2775,N_2444,N_2540);
nand U2776 (N_2776,N_2567,N_2474);
nand U2777 (N_2777,N_2485,N_2511);
xnor U2778 (N_2778,N_2550,N_2430);
and U2779 (N_2779,N_2589,N_2541);
nand U2780 (N_2780,N_2445,N_2549);
nor U2781 (N_2781,N_2425,N_2554);
and U2782 (N_2782,N_2467,N_2543);
or U2783 (N_2783,N_2587,N_2414);
and U2784 (N_2784,N_2413,N_2404);
and U2785 (N_2785,N_2594,N_2478);
nor U2786 (N_2786,N_2417,N_2429);
and U2787 (N_2787,N_2585,N_2458);
nand U2788 (N_2788,N_2561,N_2435);
and U2789 (N_2789,N_2486,N_2575);
or U2790 (N_2790,N_2559,N_2480);
nor U2791 (N_2791,N_2491,N_2409);
nor U2792 (N_2792,N_2588,N_2533);
or U2793 (N_2793,N_2404,N_2550);
or U2794 (N_2794,N_2525,N_2439);
nor U2795 (N_2795,N_2536,N_2492);
xor U2796 (N_2796,N_2506,N_2466);
or U2797 (N_2797,N_2579,N_2566);
nor U2798 (N_2798,N_2505,N_2572);
xnor U2799 (N_2799,N_2470,N_2526);
or U2800 (N_2800,N_2761,N_2615);
nand U2801 (N_2801,N_2714,N_2716);
nor U2802 (N_2802,N_2609,N_2725);
xnor U2803 (N_2803,N_2684,N_2629);
nor U2804 (N_2804,N_2666,N_2766);
nor U2805 (N_2805,N_2775,N_2641);
nor U2806 (N_2806,N_2763,N_2786);
xnor U2807 (N_2807,N_2648,N_2784);
xor U2808 (N_2808,N_2650,N_2799);
xor U2809 (N_2809,N_2633,N_2652);
or U2810 (N_2810,N_2721,N_2625);
and U2811 (N_2811,N_2793,N_2731);
or U2812 (N_2812,N_2690,N_2760);
nor U2813 (N_2813,N_2749,N_2751);
nor U2814 (N_2814,N_2737,N_2774);
or U2815 (N_2815,N_2767,N_2722);
or U2816 (N_2816,N_2671,N_2602);
or U2817 (N_2817,N_2733,N_2709);
and U2818 (N_2818,N_2619,N_2742);
nor U2819 (N_2819,N_2655,N_2768);
and U2820 (N_2820,N_2620,N_2656);
nand U2821 (N_2821,N_2753,N_2704);
and U2822 (N_2822,N_2638,N_2682);
nand U2823 (N_2823,N_2632,N_2739);
or U2824 (N_2824,N_2715,N_2644);
or U2825 (N_2825,N_2667,N_2796);
or U2826 (N_2826,N_2747,N_2734);
nand U2827 (N_2827,N_2635,N_2788);
xor U2828 (N_2828,N_2705,N_2643);
and U2829 (N_2829,N_2701,N_2732);
or U2830 (N_2830,N_2678,N_2694);
xnor U2831 (N_2831,N_2614,N_2745);
xnor U2832 (N_2832,N_2624,N_2675);
or U2833 (N_2833,N_2706,N_2683);
xnor U2834 (N_2834,N_2617,N_2670);
or U2835 (N_2835,N_2627,N_2699);
or U2836 (N_2836,N_2639,N_2673);
nand U2837 (N_2837,N_2770,N_2718);
and U2838 (N_2838,N_2657,N_2728);
and U2839 (N_2839,N_2622,N_2794);
nand U2840 (N_2840,N_2750,N_2634);
nor U2841 (N_2841,N_2758,N_2748);
xnor U2842 (N_2842,N_2792,N_2754);
and U2843 (N_2843,N_2689,N_2752);
nand U2844 (N_2844,N_2736,N_2623);
and U2845 (N_2845,N_2746,N_2759);
or U2846 (N_2846,N_2695,N_2698);
nor U2847 (N_2847,N_2646,N_2783);
and U2848 (N_2848,N_2631,N_2727);
nor U2849 (N_2849,N_2743,N_2703);
and U2850 (N_2850,N_2755,N_2658);
or U2851 (N_2851,N_2654,N_2661);
xnor U2852 (N_2852,N_2708,N_2659);
nor U2853 (N_2853,N_2756,N_2691);
nand U2854 (N_2854,N_2710,N_2687);
xor U2855 (N_2855,N_2744,N_2681);
or U2856 (N_2856,N_2712,N_2740);
xnor U2857 (N_2857,N_2613,N_2647);
or U2858 (N_2858,N_2677,N_2789);
and U2859 (N_2859,N_2771,N_2669);
or U2860 (N_2860,N_2676,N_2610);
xor U2861 (N_2861,N_2779,N_2680);
nand U2862 (N_2862,N_2757,N_2780);
or U2863 (N_2863,N_2685,N_2713);
nand U2864 (N_2864,N_2664,N_2640);
xor U2865 (N_2865,N_2787,N_2662);
xor U2866 (N_2866,N_2621,N_2636);
nand U2867 (N_2867,N_2618,N_2711);
and U2868 (N_2868,N_2653,N_2762);
and U2869 (N_2869,N_2605,N_2791);
and U2870 (N_2870,N_2637,N_2798);
nor U2871 (N_2871,N_2692,N_2778);
xnor U2872 (N_2872,N_2723,N_2628);
nand U2873 (N_2873,N_2608,N_2773);
and U2874 (N_2874,N_2741,N_2612);
and U2875 (N_2875,N_2630,N_2688);
nand U2876 (N_2876,N_2679,N_2672);
xnor U2877 (N_2877,N_2797,N_2642);
or U2878 (N_2878,N_2772,N_2665);
nand U2879 (N_2879,N_2781,N_2776);
nor U2880 (N_2880,N_2611,N_2702);
and U2881 (N_2881,N_2645,N_2600);
nand U2882 (N_2882,N_2663,N_2730);
or U2883 (N_2883,N_2777,N_2651);
xnor U2884 (N_2884,N_2795,N_2604);
nor U2885 (N_2885,N_2790,N_2693);
and U2886 (N_2886,N_2717,N_2735);
or U2887 (N_2887,N_2707,N_2785);
xor U2888 (N_2888,N_2782,N_2649);
or U2889 (N_2889,N_2720,N_2686);
nor U2890 (N_2890,N_2626,N_2660);
and U2891 (N_2891,N_2726,N_2769);
nand U2892 (N_2892,N_2601,N_2607);
and U2893 (N_2893,N_2603,N_2674);
and U2894 (N_2894,N_2738,N_2729);
or U2895 (N_2895,N_2696,N_2616);
nand U2896 (N_2896,N_2697,N_2724);
nand U2897 (N_2897,N_2668,N_2700);
or U2898 (N_2898,N_2764,N_2719);
nand U2899 (N_2899,N_2765,N_2606);
nor U2900 (N_2900,N_2620,N_2627);
or U2901 (N_2901,N_2702,N_2712);
nor U2902 (N_2902,N_2664,N_2632);
xor U2903 (N_2903,N_2731,N_2735);
or U2904 (N_2904,N_2734,N_2667);
and U2905 (N_2905,N_2720,N_2791);
or U2906 (N_2906,N_2659,N_2648);
or U2907 (N_2907,N_2603,N_2737);
and U2908 (N_2908,N_2660,N_2798);
nand U2909 (N_2909,N_2764,N_2691);
nand U2910 (N_2910,N_2774,N_2700);
nor U2911 (N_2911,N_2659,N_2764);
xnor U2912 (N_2912,N_2740,N_2748);
xor U2913 (N_2913,N_2663,N_2705);
xnor U2914 (N_2914,N_2601,N_2750);
nand U2915 (N_2915,N_2725,N_2745);
xnor U2916 (N_2916,N_2651,N_2739);
or U2917 (N_2917,N_2680,N_2619);
nand U2918 (N_2918,N_2695,N_2667);
or U2919 (N_2919,N_2642,N_2774);
and U2920 (N_2920,N_2786,N_2743);
xnor U2921 (N_2921,N_2701,N_2687);
or U2922 (N_2922,N_2614,N_2749);
and U2923 (N_2923,N_2634,N_2658);
and U2924 (N_2924,N_2766,N_2772);
nor U2925 (N_2925,N_2776,N_2614);
or U2926 (N_2926,N_2636,N_2654);
nand U2927 (N_2927,N_2679,N_2661);
and U2928 (N_2928,N_2678,N_2746);
or U2929 (N_2929,N_2778,N_2726);
or U2930 (N_2930,N_2713,N_2632);
xnor U2931 (N_2931,N_2608,N_2776);
nand U2932 (N_2932,N_2606,N_2799);
or U2933 (N_2933,N_2767,N_2708);
xor U2934 (N_2934,N_2604,N_2718);
nand U2935 (N_2935,N_2669,N_2759);
xor U2936 (N_2936,N_2724,N_2619);
xnor U2937 (N_2937,N_2764,N_2755);
or U2938 (N_2938,N_2644,N_2714);
nand U2939 (N_2939,N_2604,N_2683);
or U2940 (N_2940,N_2746,N_2758);
nor U2941 (N_2941,N_2690,N_2608);
or U2942 (N_2942,N_2789,N_2746);
or U2943 (N_2943,N_2648,N_2600);
nand U2944 (N_2944,N_2639,N_2700);
nand U2945 (N_2945,N_2789,N_2665);
and U2946 (N_2946,N_2710,N_2664);
or U2947 (N_2947,N_2785,N_2655);
nor U2948 (N_2948,N_2695,N_2656);
and U2949 (N_2949,N_2792,N_2633);
nor U2950 (N_2950,N_2636,N_2780);
nand U2951 (N_2951,N_2766,N_2613);
nand U2952 (N_2952,N_2793,N_2603);
nor U2953 (N_2953,N_2741,N_2678);
or U2954 (N_2954,N_2785,N_2609);
or U2955 (N_2955,N_2795,N_2654);
and U2956 (N_2956,N_2766,N_2693);
and U2957 (N_2957,N_2682,N_2743);
nand U2958 (N_2958,N_2735,N_2743);
nor U2959 (N_2959,N_2742,N_2766);
nand U2960 (N_2960,N_2651,N_2755);
or U2961 (N_2961,N_2612,N_2755);
xor U2962 (N_2962,N_2604,N_2730);
xnor U2963 (N_2963,N_2642,N_2777);
nand U2964 (N_2964,N_2772,N_2637);
nor U2965 (N_2965,N_2709,N_2756);
or U2966 (N_2966,N_2653,N_2716);
nand U2967 (N_2967,N_2605,N_2660);
xnor U2968 (N_2968,N_2635,N_2747);
xor U2969 (N_2969,N_2697,N_2600);
or U2970 (N_2970,N_2656,N_2680);
xor U2971 (N_2971,N_2709,N_2779);
or U2972 (N_2972,N_2712,N_2757);
or U2973 (N_2973,N_2624,N_2782);
nand U2974 (N_2974,N_2709,N_2623);
nor U2975 (N_2975,N_2736,N_2690);
nor U2976 (N_2976,N_2742,N_2688);
or U2977 (N_2977,N_2781,N_2702);
and U2978 (N_2978,N_2665,N_2643);
nand U2979 (N_2979,N_2656,N_2676);
or U2980 (N_2980,N_2709,N_2715);
or U2981 (N_2981,N_2748,N_2714);
xor U2982 (N_2982,N_2618,N_2714);
or U2983 (N_2983,N_2675,N_2656);
nand U2984 (N_2984,N_2750,N_2633);
and U2985 (N_2985,N_2671,N_2785);
nor U2986 (N_2986,N_2761,N_2716);
xor U2987 (N_2987,N_2652,N_2710);
nand U2988 (N_2988,N_2714,N_2624);
and U2989 (N_2989,N_2693,N_2763);
xor U2990 (N_2990,N_2783,N_2638);
nand U2991 (N_2991,N_2741,N_2666);
or U2992 (N_2992,N_2698,N_2700);
nor U2993 (N_2993,N_2644,N_2787);
or U2994 (N_2994,N_2626,N_2649);
and U2995 (N_2995,N_2754,N_2610);
nand U2996 (N_2996,N_2698,N_2626);
and U2997 (N_2997,N_2779,N_2696);
or U2998 (N_2998,N_2606,N_2701);
xnor U2999 (N_2999,N_2719,N_2771);
and U3000 (N_3000,N_2974,N_2973);
nand U3001 (N_3001,N_2955,N_2909);
or U3002 (N_3002,N_2906,N_2837);
xnor U3003 (N_3003,N_2954,N_2975);
and U3004 (N_3004,N_2825,N_2891);
xnor U3005 (N_3005,N_2811,N_2856);
nor U3006 (N_3006,N_2927,N_2847);
xnor U3007 (N_3007,N_2858,N_2862);
xor U3008 (N_3008,N_2816,N_2870);
or U3009 (N_3009,N_2941,N_2923);
or U3010 (N_3010,N_2874,N_2890);
xor U3011 (N_3011,N_2866,N_2828);
xnor U3012 (N_3012,N_2972,N_2822);
nand U3013 (N_3013,N_2885,N_2841);
nand U3014 (N_3014,N_2865,N_2814);
or U3015 (N_3015,N_2996,N_2873);
or U3016 (N_3016,N_2881,N_2971);
or U3017 (N_3017,N_2989,N_2898);
and U3018 (N_3018,N_2809,N_2976);
and U3019 (N_3019,N_2857,N_2838);
nand U3020 (N_3020,N_2805,N_2995);
or U3021 (N_3021,N_2854,N_2876);
or U3022 (N_3022,N_2926,N_2820);
nand U3023 (N_3023,N_2978,N_2803);
nand U3024 (N_3024,N_2907,N_2864);
or U3025 (N_3025,N_2892,N_2932);
nand U3026 (N_3026,N_2986,N_2928);
xnor U3027 (N_3027,N_2846,N_2819);
xnor U3028 (N_3028,N_2908,N_2951);
xnor U3029 (N_3029,N_2880,N_2912);
nand U3030 (N_3030,N_2813,N_2947);
and U3031 (N_3031,N_2879,N_2990);
nand U3032 (N_3032,N_2903,N_2897);
or U3033 (N_3033,N_2987,N_2829);
nor U3034 (N_3034,N_2935,N_2861);
xor U3035 (N_3035,N_2920,N_2895);
xor U3036 (N_3036,N_2807,N_2888);
nor U3037 (N_3037,N_2969,N_2868);
xor U3038 (N_3038,N_2872,N_2843);
nand U3039 (N_3039,N_2842,N_2966);
nand U3040 (N_3040,N_2802,N_2899);
nor U3041 (N_3041,N_2877,N_2934);
and U3042 (N_3042,N_2961,N_2806);
xor U3043 (N_3043,N_2939,N_2942);
nor U3044 (N_3044,N_2833,N_2921);
nand U3045 (N_3045,N_2911,N_2937);
and U3046 (N_3046,N_2882,N_2998);
and U3047 (N_3047,N_2982,N_2808);
and U3048 (N_3048,N_2924,N_2992);
or U3049 (N_3049,N_2867,N_2844);
nor U3050 (N_3050,N_2860,N_2940);
nor U3051 (N_3051,N_2889,N_2810);
or U3052 (N_3052,N_2804,N_2917);
nor U3053 (N_3053,N_2950,N_2958);
nand U3054 (N_3054,N_2902,N_2968);
nand U3055 (N_3055,N_2994,N_2945);
nor U3056 (N_3056,N_2904,N_2981);
xor U3057 (N_3057,N_2824,N_2812);
or U3058 (N_3058,N_2970,N_2884);
xnor U3059 (N_3059,N_2993,N_2896);
nand U3060 (N_3060,N_2850,N_2848);
and U3061 (N_3061,N_2869,N_2997);
or U3062 (N_3062,N_2916,N_2988);
or U3063 (N_3063,N_2979,N_2913);
nor U3064 (N_3064,N_2963,N_2894);
and U3065 (N_3065,N_2818,N_2823);
nand U3066 (N_3066,N_2977,N_2827);
or U3067 (N_3067,N_2836,N_2956);
and U3068 (N_3068,N_2815,N_2914);
nor U3069 (N_3069,N_2871,N_2826);
or U3070 (N_3070,N_2938,N_2964);
nand U3071 (N_3071,N_2946,N_2817);
xor U3072 (N_3072,N_2830,N_2952);
nor U3073 (N_3073,N_2915,N_2943);
or U3074 (N_3074,N_2863,N_2859);
or U3075 (N_3075,N_2984,N_2851);
xor U3076 (N_3076,N_2983,N_2801);
xor U3077 (N_3077,N_2919,N_2834);
or U3078 (N_3078,N_2900,N_2901);
or U3079 (N_3079,N_2887,N_2960);
and U3080 (N_3080,N_2929,N_2883);
nor U3081 (N_3081,N_2849,N_2832);
xnor U3082 (N_3082,N_2953,N_2949);
xnor U3083 (N_3083,N_2980,N_2922);
nand U3084 (N_3084,N_2991,N_2831);
xor U3085 (N_3085,N_2839,N_2936);
and U3086 (N_3086,N_2878,N_2845);
nor U3087 (N_3087,N_2835,N_2840);
nand U3088 (N_3088,N_2875,N_2800);
xor U3089 (N_3089,N_2930,N_2910);
and U3090 (N_3090,N_2886,N_2957);
and U3091 (N_3091,N_2925,N_2999);
or U3092 (N_3092,N_2855,N_2962);
xor U3093 (N_3093,N_2905,N_2965);
and U3094 (N_3094,N_2931,N_2918);
nand U3095 (N_3095,N_2967,N_2933);
nor U3096 (N_3096,N_2853,N_2959);
xor U3097 (N_3097,N_2985,N_2821);
xor U3098 (N_3098,N_2948,N_2893);
or U3099 (N_3099,N_2944,N_2852);
xnor U3100 (N_3100,N_2966,N_2902);
nor U3101 (N_3101,N_2857,N_2997);
nand U3102 (N_3102,N_2835,N_2924);
or U3103 (N_3103,N_2801,N_2963);
xor U3104 (N_3104,N_2934,N_2947);
or U3105 (N_3105,N_2880,N_2983);
and U3106 (N_3106,N_2860,N_2831);
or U3107 (N_3107,N_2822,N_2826);
xnor U3108 (N_3108,N_2816,N_2914);
or U3109 (N_3109,N_2893,N_2875);
xor U3110 (N_3110,N_2809,N_2956);
nand U3111 (N_3111,N_2960,N_2953);
or U3112 (N_3112,N_2866,N_2881);
nor U3113 (N_3113,N_2895,N_2822);
xnor U3114 (N_3114,N_2814,N_2935);
nor U3115 (N_3115,N_2937,N_2899);
or U3116 (N_3116,N_2816,N_2819);
nand U3117 (N_3117,N_2995,N_2821);
and U3118 (N_3118,N_2836,N_2820);
xor U3119 (N_3119,N_2842,N_2965);
or U3120 (N_3120,N_2839,N_2969);
nand U3121 (N_3121,N_2924,N_2930);
and U3122 (N_3122,N_2927,N_2875);
nor U3123 (N_3123,N_2841,N_2832);
and U3124 (N_3124,N_2807,N_2810);
nor U3125 (N_3125,N_2920,N_2914);
xor U3126 (N_3126,N_2976,N_2924);
or U3127 (N_3127,N_2957,N_2800);
and U3128 (N_3128,N_2885,N_2831);
and U3129 (N_3129,N_2801,N_2816);
and U3130 (N_3130,N_2922,N_2822);
or U3131 (N_3131,N_2978,N_2825);
or U3132 (N_3132,N_2955,N_2917);
xor U3133 (N_3133,N_2864,N_2832);
or U3134 (N_3134,N_2981,N_2986);
xnor U3135 (N_3135,N_2825,N_2801);
xnor U3136 (N_3136,N_2997,N_2853);
or U3137 (N_3137,N_2998,N_2918);
or U3138 (N_3138,N_2832,N_2946);
nor U3139 (N_3139,N_2830,N_2987);
nand U3140 (N_3140,N_2874,N_2845);
xnor U3141 (N_3141,N_2887,N_2828);
xor U3142 (N_3142,N_2802,N_2902);
nand U3143 (N_3143,N_2874,N_2964);
xor U3144 (N_3144,N_2843,N_2904);
nand U3145 (N_3145,N_2893,N_2998);
nor U3146 (N_3146,N_2836,N_2973);
or U3147 (N_3147,N_2946,N_2969);
nand U3148 (N_3148,N_2869,N_2802);
xnor U3149 (N_3149,N_2817,N_2975);
or U3150 (N_3150,N_2903,N_2822);
nor U3151 (N_3151,N_2866,N_2923);
nor U3152 (N_3152,N_2866,N_2933);
or U3153 (N_3153,N_2853,N_2812);
nand U3154 (N_3154,N_2881,N_2931);
and U3155 (N_3155,N_2928,N_2810);
nand U3156 (N_3156,N_2887,N_2800);
xor U3157 (N_3157,N_2844,N_2897);
and U3158 (N_3158,N_2934,N_2924);
xor U3159 (N_3159,N_2935,N_2894);
nor U3160 (N_3160,N_2887,N_2944);
xnor U3161 (N_3161,N_2864,N_2892);
xor U3162 (N_3162,N_2852,N_2983);
xor U3163 (N_3163,N_2942,N_2902);
nor U3164 (N_3164,N_2845,N_2946);
and U3165 (N_3165,N_2909,N_2805);
nand U3166 (N_3166,N_2934,N_2992);
nor U3167 (N_3167,N_2808,N_2833);
nor U3168 (N_3168,N_2976,N_2918);
or U3169 (N_3169,N_2822,N_2831);
or U3170 (N_3170,N_2848,N_2962);
or U3171 (N_3171,N_2970,N_2922);
nand U3172 (N_3172,N_2865,N_2822);
xnor U3173 (N_3173,N_2803,N_2931);
nand U3174 (N_3174,N_2996,N_2979);
xor U3175 (N_3175,N_2821,N_2815);
nor U3176 (N_3176,N_2871,N_2938);
or U3177 (N_3177,N_2963,N_2989);
or U3178 (N_3178,N_2834,N_2822);
nor U3179 (N_3179,N_2984,N_2802);
nor U3180 (N_3180,N_2973,N_2995);
nor U3181 (N_3181,N_2890,N_2818);
and U3182 (N_3182,N_2865,N_2886);
nor U3183 (N_3183,N_2839,N_2872);
nor U3184 (N_3184,N_2852,N_2899);
nand U3185 (N_3185,N_2873,N_2859);
and U3186 (N_3186,N_2961,N_2954);
xor U3187 (N_3187,N_2926,N_2849);
nand U3188 (N_3188,N_2866,N_2947);
nor U3189 (N_3189,N_2826,N_2945);
or U3190 (N_3190,N_2837,N_2962);
and U3191 (N_3191,N_2831,N_2982);
and U3192 (N_3192,N_2989,N_2975);
nand U3193 (N_3193,N_2882,N_2805);
nand U3194 (N_3194,N_2978,N_2935);
xnor U3195 (N_3195,N_2832,N_2979);
xor U3196 (N_3196,N_2826,N_2861);
or U3197 (N_3197,N_2906,N_2905);
or U3198 (N_3198,N_2930,N_2805);
xor U3199 (N_3199,N_2846,N_2996);
xnor U3200 (N_3200,N_3070,N_3122);
nor U3201 (N_3201,N_3099,N_3081);
xnor U3202 (N_3202,N_3075,N_3023);
nor U3203 (N_3203,N_3160,N_3130);
nor U3204 (N_3204,N_3091,N_3012);
xor U3205 (N_3205,N_3129,N_3008);
or U3206 (N_3206,N_3123,N_3180);
nand U3207 (N_3207,N_3127,N_3197);
and U3208 (N_3208,N_3189,N_3108);
nand U3209 (N_3209,N_3114,N_3131);
nand U3210 (N_3210,N_3198,N_3051);
nor U3211 (N_3211,N_3097,N_3034);
and U3212 (N_3212,N_3046,N_3173);
xor U3213 (N_3213,N_3086,N_3104);
xnor U3214 (N_3214,N_3025,N_3192);
nor U3215 (N_3215,N_3052,N_3098);
and U3216 (N_3216,N_3026,N_3067);
and U3217 (N_3217,N_3037,N_3007);
xnor U3218 (N_3218,N_3177,N_3141);
and U3219 (N_3219,N_3056,N_3065);
and U3220 (N_3220,N_3027,N_3121);
and U3221 (N_3221,N_3041,N_3149);
and U3222 (N_3222,N_3009,N_3029);
or U3223 (N_3223,N_3186,N_3115);
nor U3224 (N_3224,N_3182,N_3014);
nand U3225 (N_3225,N_3080,N_3001);
nor U3226 (N_3226,N_3168,N_3040);
or U3227 (N_3227,N_3054,N_3132);
nand U3228 (N_3228,N_3015,N_3120);
and U3229 (N_3229,N_3083,N_3154);
or U3230 (N_3230,N_3107,N_3110);
xnor U3231 (N_3231,N_3077,N_3092);
and U3232 (N_3232,N_3150,N_3148);
xor U3233 (N_3233,N_3116,N_3044);
nand U3234 (N_3234,N_3109,N_3060);
xor U3235 (N_3235,N_3159,N_3050);
or U3236 (N_3236,N_3006,N_3024);
and U3237 (N_3237,N_3158,N_3066);
xor U3238 (N_3238,N_3035,N_3011);
nand U3239 (N_3239,N_3094,N_3128);
nor U3240 (N_3240,N_3076,N_3117);
nor U3241 (N_3241,N_3181,N_3157);
nand U3242 (N_3242,N_3093,N_3048);
xnor U3243 (N_3243,N_3096,N_3018);
or U3244 (N_3244,N_3195,N_3085);
xor U3245 (N_3245,N_3119,N_3071);
or U3246 (N_3246,N_3161,N_3118);
nand U3247 (N_3247,N_3072,N_3064);
or U3248 (N_3248,N_3038,N_3171);
and U3249 (N_3249,N_3089,N_3095);
or U3250 (N_3250,N_3021,N_3191);
nand U3251 (N_3251,N_3088,N_3151);
nor U3252 (N_3252,N_3004,N_3084);
or U3253 (N_3253,N_3111,N_3152);
xor U3254 (N_3254,N_3124,N_3045);
or U3255 (N_3255,N_3000,N_3153);
nor U3256 (N_3256,N_3100,N_3178);
nor U3257 (N_3257,N_3169,N_3032);
nor U3258 (N_3258,N_3142,N_3135);
or U3259 (N_3259,N_3090,N_3101);
xor U3260 (N_3260,N_3112,N_3069);
xor U3261 (N_3261,N_3106,N_3126);
or U3262 (N_3262,N_3176,N_3047);
and U3263 (N_3263,N_3102,N_3188);
and U3264 (N_3264,N_3031,N_3033);
nor U3265 (N_3265,N_3162,N_3183);
nand U3266 (N_3266,N_3010,N_3113);
and U3267 (N_3267,N_3194,N_3184);
or U3268 (N_3268,N_3030,N_3147);
or U3269 (N_3269,N_3187,N_3042);
and U3270 (N_3270,N_3053,N_3059);
xor U3271 (N_3271,N_3156,N_3002);
or U3272 (N_3272,N_3016,N_3179);
nor U3273 (N_3273,N_3105,N_3172);
and U3274 (N_3274,N_3125,N_3199);
and U3275 (N_3275,N_3013,N_3166);
nand U3276 (N_3276,N_3165,N_3028);
and U3277 (N_3277,N_3140,N_3138);
and U3278 (N_3278,N_3163,N_3145);
nand U3279 (N_3279,N_3022,N_3079);
nand U3280 (N_3280,N_3057,N_3136);
nor U3281 (N_3281,N_3068,N_3103);
nand U3282 (N_3282,N_3144,N_3193);
nand U3283 (N_3283,N_3055,N_3134);
or U3284 (N_3284,N_3146,N_3164);
or U3285 (N_3285,N_3175,N_3143);
xor U3286 (N_3286,N_3174,N_3036);
or U3287 (N_3287,N_3082,N_3003);
or U3288 (N_3288,N_3137,N_3019);
and U3289 (N_3289,N_3074,N_3058);
and U3290 (N_3290,N_3049,N_3170);
xor U3291 (N_3291,N_3039,N_3190);
or U3292 (N_3292,N_3062,N_3043);
and U3293 (N_3293,N_3185,N_3005);
xnor U3294 (N_3294,N_3061,N_3073);
nor U3295 (N_3295,N_3087,N_3078);
nand U3296 (N_3296,N_3020,N_3196);
nand U3297 (N_3297,N_3139,N_3063);
and U3298 (N_3298,N_3017,N_3167);
and U3299 (N_3299,N_3155,N_3133);
and U3300 (N_3300,N_3045,N_3185);
xnor U3301 (N_3301,N_3029,N_3086);
nor U3302 (N_3302,N_3085,N_3194);
nor U3303 (N_3303,N_3152,N_3190);
xor U3304 (N_3304,N_3172,N_3083);
and U3305 (N_3305,N_3168,N_3193);
nand U3306 (N_3306,N_3054,N_3112);
and U3307 (N_3307,N_3028,N_3053);
or U3308 (N_3308,N_3091,N_3020);
nand U3309 (N_3309,N_3111,N_3100);
and U3310 (N_3310,N_3180,N_3177);
xnor U3311 (N_3311,N_3192,N_3078);
or U3312 (N_3312,N_3169,N_3021);
and U3313 (N_3313,N_3033,N_3004);
nor U3314 (N_3314,N_3017,N_3082);
nor U3315 (N_3315,N_3019,N_3136);
nand U3316 (N_3316,N_3113,N_3174);
or U3317 (N_3317,N_3012,N_3054);
or U3318 (N_3318,N_3028,N_3188);
nor U3319 (N_3319,N_3178,N_3034);
and U3320 (N_3320,N_3071,N_3193);
nor U3321 (N_3321,N_3180,N_3157);
or U3322 (N_3322,N_3037,N_3137);
and U3323 (N_3323,N_3176,N_3072);
or U3324 (N_3324,N_3094,N_3181);
or U3325 (N_3325,N_3078,N_3015);
xor U3326 (N_3326,N_3022,N_3187);
nand U3327 (N_3327,N_3053,N_3049);
or U3328 (N_3328,N_3147,N_3102);
nand U3329 (N_3329,N_3133,N_3152);
or U3330 (N_3330,N_3169,N_3137);
nand U3331 (N_3331,N_3151,N_3021);
xor U3332 (N_3332,N_3039,N_3056);
and U3333 (N_3333,N_3100,N_3078);
nor U3334 (N_3334,N_3018,N_3102);
and U3335 (N_3335,N_3147,N_3068);
nand U3336 (N_3336,N_3093,N_3094);
and U3337 (N_3337,N_3160,N_3036);
nand U3338 (N_3338,N_3124,N_3080);
xor U3339 (N_3339,N_3161,N_3057);
xnor U3340 (N_3340,N_3151,N_3142);
nor U3341 (N_3341,N_3076,N_3118);
xor U3342 (N_3342,N_3137,N_3171);
nor U3343 (N_3343,N_3030,N_3024);
or U3344 (N_3344,N_3048,N_3108);
and U3345 (N_3345,N_3192,N_3165);
and U3346 (N_3346,N_3148,N_3063);
xor U3347 (N_3347,N_3161,N_3018);
and U3348 (N_3348,N_3025,N_3035);
xor U3349 (N_3349,N_3147,N_3088);
or U3350 (N_3350,N_3122,N_3185);
nand U3351 (N_3351,N_3149,N_3166);
nor U3352 (N_3352,N_3121,N_3143);
nand U3353 (N_3353,N_3124,N_3048);
or U3354 (N_3354,N_3168,N_3161);
or U3355 (N_3355,N_3017,N_3050);
nor U3356 (N_3356,N_3068,N_3156);
nand U3357 (N_3357,N_3084,N_3047);
or U3358 (N_3358,N_3067,N_3190);
and U3359 (N_3359,N_3135,N_3189);
or U3360 (N_3360,N_3052,N_3075);
or U3361 (N_3361,N_3186,N_3062);
nor U3362 (N_3362,N_3133,N_3174);
nor U3363 (N_3363,N_3098,N_3034);
and U3364 (N_3364,N_3176,N_3196);
and U3365 (N_3365,N_3029,N_3142);
nand U3366 (N_3366,N_3028,N_3065);
xor U3367 (N_3367,N_3164,N_3079);
nand U3368 (N_3368,N_3167,N_3113);
nand U3369 (N_3369,N_3020,N_3186);
or U3370 (N_3370,N_3107,N_3083);
nand U3371 (N_3371,N_3040,N_3116);
and U3372 (N_3372,N_3193,N_3009);
nand U3373 (N_3373,N_3146,N_3121);
and U3374 (N_3374,N_3159,N_3106);
nand U3375 (N_3375,N_3077,N_3090);
nand U3376 (N_3376,N_3126,N_3043);
xor U3377 (N_3377,N_3152,N_3047);
nor U3378 (N_3378,N_3173,N_3195);
and U3379 (N_3379,N_3005,N_3077);
nor U3380 (N_3380,N_3006,N_3017);
nor U3381 (N_3381,N_3083,N_3141);
or U3382 (N_3382,N_3154,N_3109);
nor U3383 (N_3383,N_3000,N_3143);
xnor U3384 (N_3384,N_3016,N_3037);
or U3385 (N_3385,N_3012,N_3093);
xnor U3386 (N_3386,N_3140,N_3125);
nor U3387 (N_3387,N_3020,N_3034);
nor U3388 (N_3388,N_3069,N_3059);
and U3389 (N_3389,N_3056,N_3016);
nand U3390 (N_3390,N_3064,N_3183);
and U3391 (N_3391,N_3024,N_3051);
and U3392 (N_3392,N_3140,N_3108);
nor U3393 (N_3393,N_3131,N_3142);
nand U3394 (N_3394,N_3199,N_3083);
or U3395 (N_3395,N_3109,N_3110);
or U3396 (N_3396,N_3119,N_3171);
nor U3397 (N_3397,N_3151,N_3198);
nor U3398 (N_3398,N_3043,N_3187);
nor U3399 (N_3399,N_3078,N_3072);
xnor U3400 (N_3400,N_3316,N_3334);
nand U3401 (N_3401,N_3232,N_3359);
and U3402 (N_3402,N_3395,N_3312);
xor U3403 (N_3403,N_3385,N_3336);
nand U3404 (N_3404,N_3324,N_3358);
and U3405 (N_3405,N_3218,N_3235);
nand U3406 (N_3406,N_3289,N_3343);
or U3407 (N_3407,N_3331,N_3352);
nor U3408 (N_3408,N_3306,N_3217);
nand U3409 (N_3409,N_3221,N_3297);
nor U3410 (N_3410,N_3227,N_3208);
or U3411 (N_3411,N_3398,N_3247);
nand U3412 (N_3412,N_3240,N_3201);
and U3413 (N_3413,N_3371,N_3292);
or U3414 (N_3414,N_3392,N_3287);
and U3415 (N_3415,N_3216,N_3268);
or U3416 (N_3416,N_3384,N_3285);
and U3417 (N_3417,N_3250,N_3367);
nand U3418 (N_3418,N_3326,N_3283);
nor U3419 (N_3419,N_3238,N_3323);
or U3420 (N_3420,N_3328,N_3222);
or U3421 (N_3421,N_3304,N_3231);
xor U3422 (N_3422,N_3209,N_3315);
and U3423 (N_3423,N_3399,N_3275);
nor U3424 (N_3424,N_3258,N_3303);
and U3425 (N_3425,N_3281,N_3291);
nand U3426 (N_3426,N_3251,N_3294);
or U3427 (N_3427,N_3362,N_3223);
and U3428 (N_3428,N_3338,N_3350);
nand U3429 (N_3429,N_3288,N_3224);
and U3430 (N_3430,N_3376,N_3284);
and U3431 (N_3431,N_3295,N_3205);
xor U3432 (N_3432,N_3301,N_3347);
nand U3433 (N_3433,N_3394,N_3229);
nand U3434 (N_3434,N_3349,N_3225);
and U3435 (N_3435,N_3259,N_3272);
and U3436 (N_3436,N_3299,N_3228);
or U3437 (N_3437,N_3356,N_3375);
or U3438 (N_3438,N_3345,N_3354);
and U3439 (N_3439,N_3280,N_3346);
and U3440 (N_3440,N_3246,N_3317);
and U3441 (N_3441,N_3242,N_3322);
or U3442 (N_3442,N_3339,N_3374);
or U3443 (N_3443,N_3387,N_3265);
xnor U3444 (N_3444,N_3266,N_3220);
or U3445 (N_3445,N_3377,N_3274);
or U3446 (N_3446,N_3381,N_3373);
nand U3447 (N_3447,N_3300,N_3293);
and U3448 (N_3448,N_3244,N_3340);
xor U3449 (N_3449,N_3278,N_3200);
nor U3450 (N_3450,N_3202,N_3389);
nand U3451 (N_3451,N_3363,N_3256);
and U3452 (N_3452,N_3378,N_3388);
and U3453 (N_3453,N_3310,N_3311);
nand U3454 (N_3454,N_3271,N_3397);
or U3455 (N_3455,N_3210,N_3357);
nor U3456 (N_3456,N_3333,N_3255);
nor U3457 (N_3457,N_3273,N_3369);
nor U3458 (N_3458,N_3254,N_3213);
nand U3459 (N_3459,N_3321,N_3348);
xor U3460 (N_3460,N_3344,N_3361);
xnor U3461 (N_3461,N_3267,N_3261);
xor U3462 (N_3462,N_3330,N_3342);
and U3463 (N_3463,N_3262,N_3309);
nand U3464 (N_3464,N_3351,N_3329);
and U3465 (N_3465,N_3390,N_3364);
or U3466 (N_3466,N_3263,N_3243);
or U3467 (N_3467,N_3206,N_3270);
nor U3468 (N_3468,N_3332,N_3325);
nand U3469 (N_3469,N_3365,N_3277);
nor U3470 (N_3470,N_3253,N_3234);
and U3471 (N_3471,N_3382,N_3302);
nor U3472 (N_3472,N_3319,N_3282);
xnor U3473 (N_3473,N_3236,N_3318);
nor U3474 (N_3474,N_3245,N_3298);
nor U3475 (N_3475,N_3207,N_3396);
xnor U3476 (N_3476,N_3237,N_3355);
xnor U3477 (N_3477,N_3249,N_3233);
and U3478 (N_3478,N_3214,N_3204);
nand U3479 (N_3479,N_3386,N_3335);
nand U3480 (N_3480,N_3215,N_3380);
nor U3481 (N_3481,N_3383,N_3252);
xnor U3482 (N_3482,N_3203,N_3269);
xor U3483 (N_3483,N_3230,N_3366);
or U3484 (N_3484,N_3370,N_3307);
nand U3485 (N_3485,N_3241,N_3239);
nor U3486 (N_3486,N_3212,N_3226);
xnor U3487 (N_3487,N_3391,N_3296);
nand U3488 (N_3488,N_3341,N_3286);
or U3489 (N_3489,N_3308,N_3305);
nand U3490 (N_3490,N_3279,N_3260);
nand U3491 (N_3491,N_3314,N_3372);
or U3492 (N_3492,N_3360,N_3290);
xor U3493 (N_3493,N_3257,N_3248);
nand U3494 (N_3494,N_3264,N_3393);
xnor U3495 (N_3495,N_3320,N_3379);
xnor U3496 (N_3496,N_3353,N_3327);
and U3497 (N_3497,N_3337,N_3219);
nand U3498 (N_3498,N_3313,N_3276);
or U3499 (N_3499,N_3211,N_3368);
or U3500 (N_3500,N_3327,N_3344);
nor U3501 (N_3501,N_3269,N_3353);
or U3502 (N_3502,N_3360,N_3369);
or U3503 (N_3503,N_3378,N_3299);
nand U3504 (N_3504,N_3212,N_3308);
and U3505 (N_3505,N_3280,N_3223);
nor U3506 (N_3506,N_3313,N_3219);
nor U3507 (N_3507,N_3224,N_3302);
xnor U3508 (N_3508,N_3244,N_3321);
or U3509 (N_3509,N_3342,N_3209);
and U3510 (N_3510,N_3371,N_3392);
xnor U3511 (N_3511,N_3330,N_3309);
xnor U3512 (N_3512,N_3209,N_3286);
nor U3513 (N_3513,N_3279,N_3376);
or U3514 (N_3514,N_3299,N_3200);
xnor U3515 (N_3515,N_3378,N_3385);
and U3516 (N_3516,N_3363,N_3349);
and U3517 (N_3517,N_3321,N_3223);
nand U3518 (N_3518,N_3327,N_3316);
nand U3519 (N_3519,N_3311,N_3390);
nand U3520 (N_3520,N_3394,N_3300);
nor U3521 (N_3521,N_3344,N_3223);
nand U3522 (N_3522,N_3337,N_3233);
xnor U3523 (N_3523,N_3225,N_3338);
nor U3524 (N_3524,N_3333,N_3328);
nor U3525 (N_3525,N_3394,N_3309);
nor U3526 (N_3526,N_3336,N_3397);
and U3527 (N_3527,N_3289,N_3258);
nor U3528 (N_3528,N_3389,N_3364);
nand U3529 (N_3529,N_3212,N_3310);
or U3530 (N_3530,N_3388,N_3395);
xnor U3531 (N_3531,N_3201,N_3256);
or U3532 (N_3532,N_3223,N_3380);
nand U3533 (N_3533,N_3326,N_3371);
or U3534 (N_3534,N_3287,N_3296);
or U3535 (N_3535,N_3213,N_3370);
nor U3536 (N_3536,N_3234,N_3288);
nand U3537 (N_3537,N_3393,N_3332);
nor U3538 (N_3538,N_3241,N_3249);
or U3539 (N_3539,N_3275,N_3249);
xnor U3540 (N_3540,N_3202,N_3279);
nand U3541 (N_3541,N_3349,N_3361);
nand U3542 (N_3542,N_3365,N_3208);
nor U3543 (N_3543,N_3211,N_3275);
nand U3544 (N_3544,N_3256,N_3260);
nor U3545 (N_3545,N_3201,N_3209);
nor U3546 (N_3546,N_3210,N_3231);
xor U3547 (N_3547,N_3327,N_3358);
and U3548 (N_3548,N_3352,N_3379);
xnor U3549 (N_3549,N_3210,N_3350);
nor U3550 (N_3550,N_3353,N_3392);
nor U3551 (N_3551,N_3305,N_3325);
or U3552 (N_3552,N_3216,N_3303);
xnor U3553 (N_3553,N_3375,N_3298);
nor U3554 (N_3554,N_3255,N_3320);
or U3555 (N_3555,N_3212,N_3394);
or U3556 (N_3556,N_3264,N_3288);
nand U3557 (N_3557,N_3311,N_3268);
nand U3558 (N_3558,N_3392,N_3331);
or U3559 (N_3559,N_3351,N_3206);
and U3560 (N_3560,N_3267,N_3255);
nor U3561 (N_3561,N_3272,N_3215);
nand U3562 (N_3562,N_3295,N_3392);
xnor U3563 (N_3563,N_3352,N_3369);
and U3564 (N_3564,N_3399,N_3216);
nand U3565 (N_3565,N_3328,N_3347);
xnor U3566 (N_3566,N_3316,N_3271);
nor U3567 (N_3567,N_3373,N_3310);
nand U3568 (N_3568,N_3378,N_3312);
xor U3569 (N_3569,N_3301,N_3236);
or U3570 (N_3570,N_3278,N_3207);
nand U3571 (N_3571,N_3317,N_3372);
and U3572 (N_3572,N_3288,N_3368);
nand U3573 (N_3573,N_3257,N_3389);
nor U3574 (N_3574,N_3269,N_3376);
nor U3575 (N_3575,N_3393,N_3279);
and U3576 (N_3576,N_3364,N_3363);
xnor U3577 (N_3577,N_3371,N_3234);
xor U3578 (N_3578,N_3205,N_3323);
and U3579 (N_3579,N_3319,N_3217);
nor U3580 (N_3580,N_3289,N_3287);
and U3581 (N_3581,N_3335,N_3296);
xor U3582 (N_3582,N_3236,N_3257);
and U3583 (N_3583,N_3201,N_3339);
nor U3584 (N_3584,N_3336,N_3206);
nand U3585 (N_3585,N_3278,N_3325);
xnor U3586 (N_3586,N_3295,N_3381);
nand U3587 (N_3587,N_3237,N_3232);
or U3588 (N_3588,N_3265,N_3398);
xnor U3589 (N_3589,N_3268,N_3331);
nand U3590 (N_3590,N_3272,N_3310);
or U3591 (N_3591,N_3263,N_3295);
and U3592 (N_3592,N_3346,N_3216);
xor U3593 (N_3593,N_3351,N_3216);
nor U3594 (N_3594,N_3267,N_3389);
and U3595 (N_3595,N_3236,N_3267);
xnor U3596 (N_3596,N_3350,N_3382);
or U3597 (N_3597,N_3352,N_3313);
and U3598 (N_3598,N_3266,N_3365);
nor U3599 (N_3599,N_3230,N_3206);
and U3600 (N_3600,N_3482,N_3534);
nor U3601 (N_3601,N_3540,N_3558);
nor U3602 (N_3602,N_3599,N_3524);
nor U3603 (N_3603,N_3541,N_3401);
and U3604 (N_3604,N_3598,N_3466);
xnor U3605 (N_3605,N_3458,N_3530);
xnor U3606 (N_3606,N_3441,N_3418);
nor U3607 (N_3607,N_3561,N_3456);
nor U3608 (N_3608,N_3461,N_3450);
or U3609 (N_3609,N_3426,N_3568);
xnor U3610 (N_3610,N_3517,N_3416);
nand U3611 (N_3611,N_3449,N_3547);
or U3612 (N_3612,N_3504,N_3486);
xor U3613 (N_3613,N_3481,N_3510);
and U3614 (N_3614,N_3439,N_3436);
and U3615 (N_3615,N_3538,N_3408);
or U3616 (N_3616,N_3499,N_3583);
xor U3617 (N_3617,N_3548,N_3576);
nand U3618 (N_3618,N_3485,N_3593);
nand U3619 (N_3619,N_3569,N_3406);
nand U3620 (N_3620,N_3545,N_3597);
nand U3621 (N_3621,N_3577,N_3596);
nand U3622 (N_3622,N_3529,N_3484);
xnor U3623 (N_3623,N_3442,N_3532);
xor U3624 (N_3624,N_3460,N_3565);
nand U3625 (N_3625,N_3453,N_3405);
xnor U3626 (N_3626,N_3516,N_3518);
and U3627 (N_3627,N_3472,N_3434);
nor U3628 (N_3628,N_3411,N_3417);
nand U3629 (N_3629,N_3476,N_3490);
xor U3630 (N_3630,N_3556,N_3489);
and U3631 (N_3631,N_3425,N_3457);
and U3632 (N_3632,N_3463,N_3432);
or U3633 (N_3633,N_3400,N_3559);
or U3634 (N_3634,N_3522,N_3474);
nand U3635 (N_3635,N_3551,N_3528);
xnor U3636 (N_3636,N_3487,N_3507);
and U3637 (N_3637,N_3465,N_3563);
and U3638 (N_3638,N_3550,N_3586);
nor U3639 (N_3639,N_3501,N_3494);
or U3640 (N_3640,N_3580,N_3478);
or U3641 (N_3641,N_3578,N_3575);
and U3642 (N_3642,N_3520,N_3468);
xnor U3643 (N_3643,N_3462,N_3433);
nand U3644 (N_3644,N_3536,N_3448);
nand U3645 (N_3645,N_3573,N_3553);
xor U3646 (N_3646,N_3446,N_3570);
nor U3647 (N_3647,N_3495,N_3493);
xor U3648 (N_3648,N_3506,N_3554);
nor U3649 (N_3649,N_3566,N_3491);
xnor U3650 (N_3650,N_3531,N_3475);
and U3651 (N_3651,N_3469,N_3574);
or U3652 (N_3652,N_3582,N_3473);
xor U3653 (N_3653,N_3455,N_3492);
nor U3654 (N_3654,N_3431,N_3526);
or U3655 (N_3655,N_3591,N_3527);
and U3656 (N_3656,N_3572,N_3454);
nand U3657 (N_3657,N_3423,N_3584);
nor U3658 (N_3658,N_3421,N_3430);
nor U3659 (N_3659,N_3424,N_3537);
nand U3660 (N_3660,N_3410,N_3525);
and U3661 (N_3661,N_3579,N_3543);
nor U3662 (N_3662,N_3443,N_3585);
xnor U3663 (N_3663,N_3444,N_3451);
nand U3664 (N_3664,N_3594,N_3587);
or U3665 (N_3665,N_3519,N_3503);
or U3666 (N_3666,N_3515,N_3452);
or U3667 (N_3667,N_3477,N_3514);
nand U3668 (N_3668,N_3505,N_3523);
nand U3669 (N_3669,N_3445,N_3404);
and U3670 (N_3670,N_3483,N_3459);
xnor U3671 (N_3671,N_3480,N_3564);
and U3672 (N_3672,N_3428,N_3562);
nand U3673 (N_3673,N_3511,N_3595);
nand U3674 (N_3674,N_3412,N_3414);
nand U3675 (N_3675,N_3513,N_3555);
xor U3676 (N_3676,N_3542,N_3470);
or U3677 (N_3677,N_3498,N_3438);
nand U3678 (N_3678,N_3409,N_3581);
nand U3679 (N_3679,N_3557,N_3535);
xor U3680 (N_3680,N_3509,N_3533);
or U3681 (N_3681,N_3415,N_3549);
nor U3682 (N_3682,N_3403,N_3539);
and U3683 (N_3683,N_3571,N_3521);
nand U3684 (N_3684,N_3427,N_3544);
and U3685 (N_3685,N_3502,N_3440);
or U3686 (N_3686,N_3512,N_3497);
or U3687 (N_3687,N_3592,N_3479);
or U3688 (N_3688,N_3500,N_3546);
xnor U3689 (N_3689,N_3467,N_3419);
xor U3690 (N_3690,N_3447,N_3471);
xnor U3691 (N_3691,N_3407,N_3508);
and U3692 (N_3692,N_3588,N_3464);
nand U3693 (N_3693,N_3437,N_3422);
and U3694 (N_3694,N_3590,N_3560);
xor U3695 (N_3695,N_3429,N_3552);
or U3696 (N_3696,N_3435,N_3496);
nor U3697 (N_3697,N_3589,N_3402);
nor U3698 (N_3698,N_3488,N_3413);
nor U3699 (N_3699,N_3567,N_3420);
nand U3700 (N_3700,N_3466,N_3481);
nand U3701 (N_3701,N_3442,N_3434);
nor U3702 (N_3702,N_3465,N_3452);
xnor U3703 (N_3703,N_3417,N_3414);
or U3704 (N_3704,N_3572,N_3582);
or U3705 (N_3705,N_3555,N_3552);
nor U3706 (N_3706,N_3513,N_3559);
or U3707 (N_3707,N_3497,N_3436);
or U3708 (N_3708,N_3532,N_3569);
and U3709 (N_3709,N_3549,N_3451);
nor U3710 (N_3710,N_3407,N_3518);
and U3711 (N_3711,N_3517,N_3521);
nand U3712 (N_3712,N_3561,N_3446);
nor U3713 (N_3713,N_3530,N_3465);
or U3714 (N_3714,N_3435,N_3478);
nor U3715 (N_3715,N_3440,N_3472);
xor U3716 (N_3716,N_3559,N_3511);
xor U3717 (N_3717,N_3534,N_3417);
nor U3718 (N_3718,N_3492,N_3487);
nor U3719 (N_3719,N_3515,N_3507);
or U3720 (N_3720,N_3504,N_3415);
nor U3721 (N_3721,N_3457,N_3556);
and U3722 (N_3722,N_3599,N_3534);
nand U3723 (N_3723,N_3482,N_3502);
or U3724 (N_3724,N_3418,N_3424);
nand U3725 (N_3725,N_3579,N_3411);
or U3726 (N_3726,N_3440,N_3560);
nor U3727 (N_3727,N_3501,N_3592);
nor U3728 (N_3728,N_3517,N_3572);
nor U3729 (N_3729,N_3530,N_3474);
xnor U3730 (N_3730,N_3553,N_3407);
xnor U3731 (N_3731,N_3458,N_3439);
nand U3732 (N_3732,N_3481,N_3538);
or U3733 (N_3733,N_3516,N_3529);
nand U3734 (N_3734,N_3550,N_3421);
or U3735 (N_3735,N_3524,N_3402);
nor U3736 (N_3736,N_3547,N_3425);
nand U3737 (N_3737,N_3488,N_3467);
and U3738 (N_3738,N_3594,N_3457);
xor U3739 (N_3739,N_3570,N_3452);
and U3740 (N_3740,N_3406,N_3430);
nand U3741 (N_3741,N_3431,N_3452);
nor U3742 (N_3742,N_3421,N_3511);
nand U3743 (N_3743,N_3568,N_3554);
nor U3744 (N_3744,N_3454,N_3551);
or U3745 (N_3745,N_3431,N_3492);
nor U3746 (N_3746,N_3449,N_3475);
or U3747 (N_3747,N_3525,N_3545);
and U3748 (N_3748,N_3560,N_3577);
xnor U3749 (N_3749,N_3544,N_3476);
nand U3750 (N_3750,N_3501,N_3541);
or U3751 (N_3751,N_3588,N_3485);
xor U3752 (N_3752,N_3407,N_3488);
nor U3753 (N_3753,N_3573,N_3420);
or U3754 (N_3754,N_3558,N_3573);
nand U3755 (N_3755,N_3491,N_3538);
nand U3756 (N_3756,N_3441,N_3424);
and U3757 (N_3757,N_3429,N_3409);
nor U3758 (N_3758,N_3583,N_3406);
nand U3759 (N_3759,N_3422,N_3489);
nor U3760 (N_3760,N_3421,N_3483);
nor U3761 (N_3761,N_3452,N_3451);
nor U3762 (N_3762,N_3576,N_3526);
nor U3763 (N_3763,N_3450,N_3412);
nand U3764 (N_3764,N_3593,N_3405);
or U3765 (N_3765,N_3496,N_3440);
xnor U3766 (N_3766,N_3472,N_3439);
or U3767 (N_3767,N_3532,N_3424);
xnor U3768 (N_3768,N_3457,N_3407);
xor U3769 (N_3769,N_3529,N_3559);
and U3770 (N_3770,N_3412,N_3506);
xnor U3771 (N_3771,N_3546,N_3550);
nand U3772 (N_3772,N_3454,N_3443);
nor U3773 (N_3773,N_3586,N_3541);
xor U3774 (N_3774,N_3540,N_3550);
nor U3775 (N_3775,N_3431,N_3547);
nor U3776 (N_3776,N_3548,N_3502);
nor U3777 (N_3777,N_3544,N_3530);
xnor U3778 (N_3778,N_3482,N_3517);
nand U3779 (N_3779,N_3423,N_3532);
nor U3780 (N_3780,N_3541,N_3594);
nand U3781 (N_3781,N_3553,N_3462);
xnor U3782 (N_3782,N_3490,N_3593);
xnor U3783 (N_3783,N_3434,N_3537);
nand U3784 (N_3784,N_3501,N_3511);
or U3785 (N_3785,N_3589,N_3433);
xor U3786 (N_3786,N_3462,N_3533);
xnor U3787 (N_3787,N_3528,N_3572);
or U3788 (N_3788,N_3468,N_3416);
nor U3789 (N_3789,N_3460,N_3402);
and U3790 (N_3790,N_3474,N_3507);
or U3791 (N_3791,N_3532,N_3475);
xnor U3792 (N_3792,N_3536,N_3436);
or U3793 (N_3793,N_3504,N_3423);
xnor U3794 (N_3794,N_3410,N_3461);
nand U3795 (N_3795,N_3429,N_3500);
nor U3796 (N_3796,N_3435,N_3446);
nand U3797 (N_3797,N_3594,N_3401);
xnor U3798 (N_3798,N_3408,N_3568);
nand U3799 (N_3799,N_3545,N_3555);
and U3800 (N_3800,N_3621,N_3702);
nor U3801 (N_3801,N_3639,N_3737);
xor U3802 (N_3802,N_3766,N_3778);
xor U3803 (N_3803,N_3683,N_3690);
and U3804 (N_3804,N_3751,N_3672);
xor U3805 (N_3805,N_3636,N_3638);
or U3806 (N_3806,N_3600,N_3675);
and U3807 (N_3807,N_3742,N_3635);
nor U3808 (N_3808,N_3796,N_3748);
or U3809 (N_3809,N_3789,N_3700);
xnor U3810 (N_3810,N_3604,N_3694);
or U3811 (N_3811,N_3707,N_3723);
xnor U3812 (N_3812,N_3689,N_3659);
nand U3813 (N_3813,N_3761,N_3623);
and U3814 (N_3814,N_3767,N_3719);
and U3815 (N_3815,N_3769,N_3676);
nor U3816 (N_3816,N_3661,N_3648);
or U3817 (N_3817,N_3627,N_3653);
and U3818 (N_3818,N_3651,N_3601);
nor U3819 (N_3819,N_3711,N_3791);
nand U3820 (N_3820,N_3739,N_3770);
nand U3821 (N_3821,N_3725,N_3756);
and U3822 (N_3822,N_3797,N_3734);
nor U3823 (N_3823,N_3680,N_3745);
nor U3824 (N_3824,N_3727,N_3630);
xnor U3825 (N_3825,N_3671,N_3714);
xor U3826 (N_3826,N_3697,N_3765);
nand U3827 (N_3827,N_3781,N_3677);
xnor U3828 (N_3828,N_3721,N_3617);
and U3829 (N_3829,N_3664,N_3669);
xor U3830 (N_3830,N_3691,N_3762);
xnor U3831 (N_3831,N_3724,N_3631);
nand U3832 (N_3832,N_3649,N_3624);
xor U3833 (N_3833,N_3607,N_3759);
nor U3834 (N_3834,N_3720,N_3663);
or U3835 (N_3835,N_3611,N_3795);
or U3836 (N_3836,N_3792,N_3692);
nor U3837 (N_3837,N_3755,N_3660);
xnor U3838 (N_3838,N_3655,N_3674);
and U3839 (N_3839,N_3729,N_3608);
nor U3840 (N_3840,N_3763,N_3602);
or U3841 (N_3841,N_3798,N_3634);
and U3842 (N_3842,N_3696,N_3752);
nor U3843 (N_3843,N_3656,N_3657);
nor U3844 (N_3844,N_3790,N_3668);
or U3845 (N_3845,N_3612,N_3771);
and U3846 (N_3846,N_3787,N_3643);
or U3847 (N_3847,N_3750,N_3741);
and U3848 (N_3848,N_3686,N_3757);
nor U3849 (N_3849,N_3754,N_3747);
and U3850 (N_3850,N_3666,N_3736);
xor U3851 (N_3851,N_3642,N_3646);
nor U3852 (N_3852,N_3774,N_3654);
or U3853 (N_3853,N_3760,N_3710);
and U3854 (N_3854,N_3609,N_3626);
and U3855 (N_3855,N_3799,N_3738);
xnor U3856 (N_3856,N_3753,N_3768);
or U3857 (N_3857,N_3633,N_3773);
nor U3858 (N_3858,N_3632,N_3794);
xor U3859 (N_3859,N_3645,N_3640);
or U3860 (N_3860,N_3641,N_3780);
or U3861 (N_3861,N_3722,N_3732);
xnor U3862 (N_3862,N_3740,N_3749);
or U3863 (N_3863,N_3775,N_3678);
nor U3864 (N_3864,N_3699,N_3704);
or U3865 (N_3865,N_3744,N_3667);
or U3866 (N_3866,N_3628,N_3764);
or U3867 (N_3867,N_3715,N_3673);
or U3868 (N_3868,N_3665,N_3731);
or U3869 (N_3869,N_3629,N_3603);
nor U3870 (N_3870,N_3698,N_3650);
xor U3871 (N_3871,N_3610,N_3793);
and U3872 (N_3872,N_3705,N_3644);
nor U3873 (N_3873,N_3622,N_3713);
xnor U3874 (N_3874,N_3652,N_3701);
nor U3875 (N_3875,N_3788,N_3735);
and U3876 (N_3876,N_3647,N_3708);
nand U3877 (N_3877,N_3620,N_3777);
nand U3878 (N_3878,N_3679,N_3681);
or U3879 (N_3879,N_3682,N_3684);
nor U3880 (N_3880,N_3730,N_3784);
xor U3881 (N_3881,N_3779,N_3726);
and U3882 (N_3882,N_3637,N_3706);
or U3883 (N_3883,N_3785,N_3695);
nand U3884 (N_3884,N_3718,N_3782);
nor U3885 (N_3885,N_3717,N_3783);
nand U3886 (N_3886,N_3685,N_3786);
nand U3887 (N_3887,N_3743,N_3712);
or U3888 (N_3888,N_3605,N_3614);
and U3889 (N_3889,N_3670,N_3746);
xnor U3890 (N_3890,N_3613,N_3716);
or U3891 (N_3891,N_3728,N_3615);
nand U3892 (N_3892,N_3618,N_3758);
nor U3893 (N_3893,N_3776,N_3772);
xor U3894 (N_3894,N_3662,N_3688);
or U3895 (N_3895,N_3606,N_3625);
or U3896 (N_3896,N_3703,N_3687);
or U3897 (N_3897,N_3619,N_3658);
nand U3898 (N_3898,N_3733,N_3616);
or U3899 (N_3899,N_3709,N_3693);
nand U3900 (N_3900,N_3632,N_3610);
xor U3901 (N_3901,N_3730,N_3624);
nor U3902 (N_3902,N_3746,N_3766);
nor U3903 (N_3903,N_3703,N_3696);
xnor U3904 (N_3904,N_3712,N_3791);
nand U3905 (N_3905,N_3761,N_3775);
or U3906 (N_3906,N_3748,N_3725);
or U3907 (N_3907,N_3765,N_3708);
and U3908 (N_3908,N_3631,N_3715);
nor U3909 (N_3909,N_3710,N_3792);
nand U3910 (N_3910,N_3625,N_3681);
nor U3911 (N_3911,N_3763,N_3767);
xnor U3912 (N_3912,N_3719,N_3722);
xor U3913 (N_3913,N_3707,N_3643);
nand U3914 (N_3914,N_3632,N_3677);
or U3915 (N_3915,N_3793,N_3676);
and U3916 (N_3916,N_3753,N_3618);
or U3917 (N_3917,N_3635,N_3643);
or U3918 (N_3918,N_3648,N_3749);
nor U3919 (N_3919,N_3702,N_3631);
or U3920 (N_3920,N_3717,N_3706);
xnor U3921 (N_3921,N_3691,N_3791);
nand U3922 (N_3922,N_3637,N_3682);
nor U3923 (N_3923,N_3687,N_3781);
xor U3924 (N_3924,N_3739,N_3775);
xor U3925 (N_3925,N_3606,N_3705);
nor U3926 (N_3926,N_3694,N_3661);
or U3927 (N_3927,N_3672,N_3649);
and U3928 (N_3928,N_3673,N_3753);
nor U3929 (N_3929,N_3717,N_3648);
xnor U3930 (N_3930,N_3655,N_3688);
xor U3931 (N_3931,N_3676,N_3764);
xor U3932 (N_3932,N_3658,N_3776);
nand U3933 (N_3933,N_3697,N_3669);
nor U3934 (N_3934,N_3621,N_3610);
or U3935 (N_3935,N_3649,N_3611);
or U3936 (N_3936,N_3722,N_3648);
nor U3937 (N_3937,N_3746,N_3757);
nand U3938 (N_3938,N_3768,N_3609);
xnor U3939 (N_3939,N_3701,N_3676);
or U3940 (N_3940,N_3621,N_3690);
and U3941 (N_3941,N_3670,N_3728);
nor U3942 (N_3942,N_3619,N_3677);
nor U3943 (N_3943,N_3666,N_3600);
and U3944 (N_3944,N_3700,N_3779);
and U3945 (N_3945,N_3759,N_3748);
xnor U3946 (N_3946,N_3639,N_3677);
and U3947 (N_3947,N_3761,N_3726);
and U3948 (N_3948,N_3637,N_3772);
xor U3949 (N_3949,N_3605,N_3739);
and U3950 (N_3950,N_3682,N_3655);
or U3951 (N_3951,N_3626,N_3713);
nor U3952 (N_3952,N_3690,N_3600);
and U3953 (N_3953,N_3641,N_3722);
or U3954 (N_3954,N_3616,N_3725);
nor U3955 (N_3955,N_3721,N_3741);
or U3956 (N_3956,N_3635,N_3719);
or U3957 (N_3957,N_3680,N_3672);
xor U3958 (N_3958,N_3694,N_3792);
and U3959 (N_3959,N_3723,N_3606);
nor U3960 (N_3960,N_3763,N_3715);
and U3961 (N_3961,N_3733,N_3727);
nor U3962 (N_3962,N_3601,N_3704);
nor U3963 (N_3963,N_3759,N_3617);
nor U3964 (N_3964,N_3772,N_3782);
nor U3965 (N_3965,N_3640,N_3792);
and U3966 (N_3966,N_3624,N_3785);
xor U3967 (N_3967,N_3708,N_3651);
nand U3968 (N_3968,N_3762,N_3664);
and U3969 (N_3969,N_3645,N_3763);
or U3970 (N_3970,N_3625,N_3724);
nand U3971 (N_3971,N_3736,N_3610);
xnor U3972 (N_3972,N_3626,N_3615);
and U3973 (N_3973,N_3685,N_3607);
nand U3974 (N_3974,N_3645,N_3777);
or U3975 (N_3975,N_3659,N_3679);
nor U3976 (N_3976,N_3667,N_3607);
or U3977 (N_3977,N_3637,N_3640);
or U3978 (N_3978,N_3640,N_3619);
xnor U3979 (N_3979,N_3769,N_3725);
nand U3980 (N_3980,N_3664,N_3744);
or U3981 (N_3981,N_3682,N_3783);
nor U3982 (N_3982,N_3656,N_3658);
and U3983 (N_3983,N_3697,N_3611);
and U3984 (N_3984,N_3689,N_3669);
nor U3985 (N_3985,N_3720,N_3734);
or U3986 (N_3986,N_3699,N_3753);
nand U3987 (N_3987,N_3750,N_3726);
or U3988 (N_3988,N_3792,N_3659);
nor U3989 (N_3989,N_3784,N_3657);
nand U3990 (N_3990,N_3695,N_3643);
and U3991 (N_3991,N_3647,N_3613);
nor U3992 (N_3992,N_3639,N_3724);
or U3993 (N_3993,N_3679,N_3737);
or U3994 (N_3994,N_3763,N_3731);
xor U3995 (N_3995,N_3603,N_3783);
or U3996 (N_3996,N_3784,N_3736);
and U3997 (N_3997,N_3653,N_3635);
and U3998 (N_3998,N_3742,N_3624);
or U3999 (N_3999,N_3615,N_3633);
and U4000 (N_4000,N_3945,N_3833);
nand U4001 (N_4001,N_3994,N_3952);
xnor U4002 (N_4002,N_3973,N_3832);
xnor U4003 (N_4003,N_3817,N_3921);
xnor U4004 (N_4004,N_3909,N_3811);
or U4005 (N_4005,N_3871,N_3820);
nand U4006 (N_4006,N_3987,N_3948);
nand U4007 (N_4007,N_3883,N_3935);
or U4008 (N_4008,N_3849,N_3861);
nand U4009 (N_4009,N_3838,N_3895);
xnor U4010 (N_4010,N_3988,N_3951);
xnor U4011 (N_4011,N_3940,N_3876);
nor U4012 (N_4012,N_3828,N_3950);
or U4013 (N_4013,N_3971,N_3865);
xor U4014 (N_4014,N_3864,N_3844);
nand U4015 (N_4015,N_3941,N_3834);
xor U4016 (N_4016,N_3818,N_3852);
nand U4017 (N_4017,N_3919,N_3862);
xor U4018 (N_4018,N_3809,N_3930);
nand U4019 (N_4019,N_3867,N_3915);
or U4020 (N_4020,N_3880,N_3962);
xnor U4021 (N_4021,N_3899,N_3860);
nand U4022 (N_4022,N_3819,N_3824);
xor U4023 (N_4023,N_3808,N_3914);
or U4024 (N_4024,N_3850,N_3841);
nand U4025 (N_4025,N_3890,N_3939);
nand U4026 (N_4026,N_3918,N_3953);
and U4027 (N_4027,N_3884,N_3908);
xnor U4028 (N_4028,N_3858,N_3814);
xor U4029 (N_4029,N_3972,N_3803);
nor U4030 (N_4030,N_3916,N_3957);
nor U4031 (N_4031,N_3831,N_3936);
nor U4032 (N_4032,N_3882,N_3924);
nand U4033 (N_4033,N_3801,N_3857);
nand U4034 (N_4034,N_3846,N_3998);
nor U4035 (N_4035,N_3905,N_3896);
and U4036 (N_4036,N_3874,N_3949);
or U4037 (N_4037,N_3968,N_3989);
xnor U4038 (N_4038,N_3926,N_3917);
or U4039 (N_4039,N_3845,N_3901);
nand U4040 (N_4040,N_3863,N_3879);
nand U4041 (N_4041,N_3878,N_3955);
nor U4042 (N_4042,N_3859,N_3995);
xor U4043 (N_4043,N_3847,N_3985);
nand U4044 (N_4044,N_3868,N_3893);
nand U4045 (N_4045,N_3802,N_3958);
or U4046 (N_4046,N_3856,N_3830);
nand U4047 (N_4047,N_3923,N_3969);
nor U4048 (N_4048,N_3960,N_3894);
and U4049 (N_4049,N_3843,N_3877);
nand U4050 (N_4050,N_3813,N_3888);
xnor U4051 (N_4051,N_3854,N_3815);
nor U4052 (N_4052,N_3934,N_3977);
nor U4053 (N_4053,N_3990,N_3933);
nor U4054 (N_4054,N_3822,N_3966);
xor U4055 (N_4055,N_3805,N_3944);
or U4056 (N_4056,N_3932,N_3821);
or U4057 (N_4057,N_3992,N_3910);
nor U4058 (N_4058,N_3900,N_3997);
nand U4059 (N_4059,N_3853,N_3826);
nand U4060 (N_4060,N_3891,N_3903);
xor U4061 (N_4061,N_3970,N_3980);
nor U4062 (N_4062,N_3889,N_3993);
or U4063 (N_4063,N_3938,N_3946);
xnor U4064 (N_4064,N_3892,N_3807);
and U4065 (N_4065,N_3929,N_3996);
nand U4066 (N_4066,N_3912,N_3855);
xor U4067 (N_4067,N_3800,N_3978);
xnor U4068 (N_4068,N_3851,N_3967);
xor U4069 (N_4069,N_3837,N_3963);
xnor U4070 (N_4070,N_3991,N_3906);
or U4071 (N_4071,N_3928,N_3947);
xnor U4072 (N_4072,N_3954,N_3839);
xnor U4073 (N_4073,N_3979,N_3961);
nand U4074 (N_4074,N_3983,N_3823);
and U4075 (N_4075,N_3902,N_3897);
nor U4076 (N_4076,N_3870,N_3810);
nand U4077 (N_4077,N_3975,N_3904);
xor U4078 (N_4078,N_3881,N_3925);
or U4079 (N_4079,N_3920,N_3907);
and U4080 (N_4080,N_3872,N_3964);
nor U4081 (N_4081,N_3825,N_3827);
xor U4082 (N_4082,N_3887,N_3835);
nand U4083 (N_4083,N_3942,N_3937);
nand U4084 (N_4084,N_3984,N_3922);
or U4085 (N_4085,N_3959,N_3875);
xor U4086 (N_4086,N_3956,N_3885);
nand U4087 (N_4087,N_3982,N_3869);
or U4088 (N_4088,N_3931,N_3836);
nor U4089 (N_4089,N_3999,N_3913);
or U4090 (N_4090,N_3829,N_3812);
nand U4091 (N_4091,N_3943,N_3848);
nand U4092 (N_4092,N_3976,N_3886);
nand U4093 (N_4093,N_3898,N_3927);
and U4094 (N_4094,N_3866,N_3911);
xnor U4095 (N_4095,N_3806,N_3981);
nand U4096 (N_4096,N_3873,N_3804);
nand U4097 (N_4097,N_3842,N_3974);
xor U4098 (N_4098,N_3986,N_3840);
xor U4099 (N_4099,N_3965,N_3816);
or U4100 (N_4100,N_3808,N_3835);
and U4101 (N_4101,N_3901,N_3837);
and U4102 (N_4102,N_3959,N_3837);
nand U4103 (N_4103,N_3870,N_3860);
and U4104 (N_4104,N_3967,N_3894);
nor U4105 (N_4105,N_3895,N_3944);
xor U4106 (N_4106,N_3844,N_3852);
xnor U4107 (N_4107,N_3979,N_3938);
or U4108 (N_4108,N_3823,N_3933);
xnor U4109 (N_4109,N_3876,N_3878);
and U4110 (N_4110,N_3916,N_3884);
and U4111 (N_4111,N_3935,N_3954);
and U4112 (N_4112,N_3891,N_3854);
nor U4113 (N_4113,N_3825,N_3850);
nand U4114 (N_4114,N_3834,N_3879);
nor U4115 (N_4115,N_3856,N_3989);
nand U4116 (N_4116,N_3855,N_3849);
or U4117 (N_4117,N_3836,N_3940);
or U4118 (N_4118,N_3921,N_3947);
xor U4119 (N_4119,N_3884,N_3829);
and U4120 (N_4120,N_3840,N_3892);
or U4121 (N_4121,N_3916,N_3860);
nand U4122 (N_4122,N_3850,N_3901);
nor U4123 (N_4123,N_3836,N_3819);
and U4124 (N_4124,N_3947,N_3818);
or U4125 (N_4125,N_3942,N_3888);
nor U4126 (N_4126,N_3843,N_3965);
and U4127 (N_4127,N_3894,N_3957);
or U4128 (N_4128,N_3817,N_3937);
xnor U4129 (N_4129,N_3893,N_3864);
nor U4130 (N_4130,N_3958,N_3892);
and U4131 (N_4131,N_3960,N_3804);
nand U4132 (N_4132,N_3952,N_3991);
nand U4133 (N_4133,N_3878,N_3831);
nand U4134 (N_4134,N_3810,N_3896);
and U4135 (N_4135,N_3925,N_3968);
nand U4136 (N_4136,N_3813,N_3953);
nor U4137 (N_4137,N_3935,N_3907);
or U4138 (N_4138,N_3956,N_3848);
and U4139 (N_4139,N_3902,N_3990);
or U4140 (N_4140,N_3930,N_3899);
or U4141 (N_4141,N_3918,N_3829);
nor U4142 (N_4142,N_3942,N_3819);
nor U4143 (N_4143,N_3900,N_3899);
and U4144 (N_4144,N_3851,N_3868);
xor U4145 (N_4145,N_3887,N_3994);
or U4146 (N_4146,N_3867,N_3943);
nand U4147 (N_4147,N_3883,N_3877);
and U4148 (N_4148,N_3982,N_3849);
and U4149 (N_4149,N_3898,N_3924);
and U4150 (N_4150,N_3891,N_3884);
nor U4151 (N_4151,N_3877,N_3908);
xor U4152 (N_4152,N_3848,N_3985);
xnor U4153 (N_4153,N_3936,N_3929);
and U4154 (N_4154,N_3853,N_3981);
nand U4155 (N_4155,N_3868,N_3838);
xnor U4156 (N_4156,N_3965,N_3840);
xor U4157 (N_4157,N_3957,N_3819);
xnor U4158 (N_4158,N_3984,N_3871);
xnor U4159 (N_4159,N_3822,N_3876);
nor U4160 (N_4160,N_3833,N_3809);
and U4161 (N_4161,N_3983,N_3882);
nand U4162 (N_4162,N_3940,N_3881);
nor U4163 (N_4163,N_3922,N_3970);
or U4164 (N_4164,N_3971,N_3802);
nor U4165 (N_4165,N_3902,N_3915);
xnor U4166 (N_4166,N_3984,N_3844);
nand U4167 (N_4167,N_3827,N_3934);
or U4168 (N_4168,N_3877,N_3812);
nor U4169 (N_4169,N_3800,N_3995);
or U4170 (N_4170,N_3803,N_3954);
nor U4171 (N_4171,N_3847,N_3961);
nand U4172 (N_4172,N_3858,N_3879);
xor U4173 (N_4173,N_3989,N_3993);
xor U4174 (N_4174,N_3948,N_3839);
nand U4175 (N_4175,N_3965,N_3971);
and U4176 (N_4176,N_3876,N_3958);
and U4177 (N_4177,N_3865,N_3802);
xnor U4178 (N_4178,N_3901,N_3857);
nor U4179 (N_4179,N_3840,N_3803);
xor U4180 (N_4180,N_3846,N_3947);
xor U4181 (N_4181,N_3998,N_3930);
nand U4182 (N_4182,N_3872,N_3997);
nand U4183 (N_4183,N_3965,N_3906);
or U4184 (N_4184,N_3934,N_3998);
xor U4185 (N_4185,N_3854,N_3987);
or U4186 (N_4186,N_3983,N_3820);
nor U4187 (N_4187,N_3955,N_3833);
xor U4188 (N_4188,N_3882,N_3925);
nor U4189 (N_4189,N_3854,N_3911);
or U4190 (N_4190,N_3939,N_3819);
or U4191 (N_4191,N_3868,N_3884);
nand U4192 (N_4192,N_3868,N_3975);
and U4193 (N_4193,N_3850,N_3959);
or U4194 (N_4194,N_3929,N_3979);
xnor U4195 (N_4195,N_3898,N_3809);
nand U4196 (N_4196,N_3830,N_3966);
and U4197 (N_4197,N_3984,N_3896);
nor U4198 (N_4198,N_3982,N_3920);
xor U4199 (N_4199,N_3946,N_3911);
nand U4200 (N_4200,N_4012,N_4116);
nand U4201 (N_4201,N_4159,N_4189);
or U4202 (N_4202,N_4034,N_4117);
nor U4203 (N_4203,N_4047,N_4102);
or U4204 (N_4204,N_4065,N_4179);
xnor U4205 (N_4205,N_4042,N_4180);
nor U4206 (N_4206,N_4162,N_4135);
xnor U4207 (N_4207,N_4129,N_4027);
xor U4208 (N_4208,N_4196,N_4068);
nand U4209 (N_4209,N_4053,N_4173);
or U4210 (N_4210,N_4055,N_4130);
and U4211 (N_4211,N_4061,N_4045);
nor U4212 (N_4212,N_4084,N_4126);
nor U4213 (N_4213,N_4104,N_4132);
nor U4214 (N_4214,N_4066,N_4188);
xor U4215 (N_4215,N_4051,N_4150);
and U4216 (N_4216,N_4170,N_4146);
or U4217 (N_4217,N_4094,N_4103);
nand U4218 (N_4218,N_4165,N_4167);
nand U4219 (N_4219,N_4141,N_4058);
and U4220 (N_4220,N_4006,N_4015);
nand U4221 (N_4221,N_4046,N_4054);
and U4222 (N_4222,N_4067,N_4052);
nand U4223 (N_4223,N_4093,N_4002);
xnor U4224 (N_4224,N_4059,N_4030);
nor U4225 (N_4225,N_4044,N_4166);
xnor U4226 (N_4226,N_4151,N_4194);
nor U4227 (N_4227,N_4041,N_4005);
nand U4228 (N_4228,N_4082,N_4119);
nand U4229 (N_4229,N_4021,N_4195);
xor U4230 (N_4230,N_4143,N_4097);
or U4231 (N_4231,N_4001,N_4112);
nor U4232 (N_4232,N_4137,N_4062);
and U4233 (N_4233,N_4131,N_4168);
nor U4234 (N_4234,N_4086,N_4096);
nand U4235 (N_4235,N_4035,N_4175);
xor U4236 (N_4236,N_4163,N_4176);
nor U4237 (N_4237,N_4128,N_4120);
and U4238 (N_4238,N_4043,N_4157);
nor U4239 (N_4239,N_4014,N_4088);
nand U4240 (N_4240,N_4010,N_4193);
xor U4241 (N_4241,N_4029,N_4048);
xnor U4242 (N_4242,N_4106,N_4018);
nor U4243 (N_4243,N_4114,N_4020);
xor U4244 (N_4244,N_4145,N_4024);
nand U4245 (N_4245,N_4078,N_4095);
xor U4246 (N_4246,N_4172,N_4098);
or U4247 (N_4247,N_4123,N_4164);
nor U4248 (N_4248,N_4075,N_4009);
or U4249 (N_4249,N_4108,N_4031);
and U4250 (N_4250,N_4153,N_4142);
xnor U4251 (N_4251,N_4060,N_4064);
nor U4252 (N_4252,N_4063,N_4070);
and U4253 (N_4253,N_4100,N_4049);
and U4254 (N_4254,N_4154,N_4033);
and U4255 (N_4255,N_4085,N_4022);
or U4256 (N_4256,N_4122,N_4039);
and U4257 (N_4257,N_4185,N_4107);
and U4258 (N_4258,N_4110,N_4152);
or U4259 (N_4259,N_4008,N_4174);
xor U4260 (N_4260,N_4071,N_4139);
or U4261 (N_4261,N_4149,N_4040);
and U4262 (N_4262,N_4171,N_4025);
nor U4263 (N_4263,N_4081,N_4004);
nand U4264 (N_4264,N_4007,N_4133);
xnor U4265 (N_4265,N_4169,N_4080);
nor U4266 (N_4266,N_4109,N_4187);
nor U4267 (N_4267,N_4144,N_4192);
and U4268 (N_4268,N_4023,N_4083);
nor U4269 (N_4269,N_4101,N_4115);
or U4270 (N_4270,N_4077,N_4191);
nand U4271 (N_4271,N_4136,N_4019);
and U4272 (N_4272,N_4190,N_4124);
nor U4273 (N_4273,N_4155,N_4183);
nor U4274 (N_4274,N_4003,N_4032);
and U4275 (N_4275,N_4199,N_4134);
and U4276 (N_4276,N_4198,N_4091);
or U4277 (N_4277,N_4092,N_4182);
or U4278 (N_4278,N_4076,N_4089);
nand U4279 (N_4279,N_4016,N_4178);
and U4280 (N_4280,N_4161,N_4099);
or U4281 (N_4281,N_4013,N_4073);
nor U4282 (N_4282,N_4125,N_4181);
and U4283 (N_4283,N_4037,N_4113);
nor U4284 (N_4284,N_4074,N_4017);
nand U4285 (N_4285,N_4105,N_4121);
nand U4286 (N_4286,N_4127,N_4028);
or U4287 (N_4287,N_4038,N_4079);
xnor U4288 (N_4288,N_4087,N_4118);
nand U4289 (N_4289,N_4036,N_4069);
nand U4290 (N_4290,N_4050,N_4160);
nor U4291 (N_4291,N_4148,N_4186);
xor U4292 (N_4292,N_4090,N_4056);
and U4293 (N_4293,N_4026,N_4177);
nand U4294 (N_4294,N_4140,N_4156);
nand U4295 (N_4295,N_4158,N_4072);
nor U4296 (N_4296,N_4057,N_4000);
nor U4297 (N_4297,N_4111,N_4011);
or U4298 (N_4298,N_4184,N_4197);
xor U4299 (N_4299,N_4147,N_4138);
nor U4300 (N_4300,N_4137,N_4163);
nand U4301 (N_4301,N_4192,N_4183);
nand U4302 (N_4302,N_4029,N_4074);
nor U4303 (N_4303,N_4066,N_4096);
and U4304 (N_4304,N_4051,N_4054);
nand U4305 (N_4305,N_4071,N_4110);
nand U4306 (N_4306,N_4017,N_4037);
or U4307 (N_4307,N_4041,N_4191);
xor U4308 (N_4308,N_4030,N_4076);
or U4309 (N_4309,N_4115,N_4016);
nor U4310 (N_4310,N_4157,N_4176);
xnor U4311 (N_4311,N_4047,N_4125);
xor U4312 (N_4312,N_4028,N_4033);
nor U4313 (N_4313,N_4005,N_4093);
nand U4314 (N_4314,N_4041,N_4150);
nand U4315 (N_4315,N_4110,N_4086);
nand U4316 (N_4316,N_4055,N_4031);
and U4317 (N_4317,N_4138,N_4047);
or U4318 (N_4318,N_4132,N_4007);
or U4319 (N_4319,N_4170,N_4198);
nand U4320 (N_4320,N_4101,N_4032);
nand U4321 (N_4321,N_4143,N_4037);
xnor U4322 (N_4322,N_4118,N_4016);
nand U4323 (N_4323,N_4161,N_4152);
or U4324 (N_4324,N_4189,N_4198);
nand U4325 (N_4325,N_4157,N_4139);
nor U4326 (N_4326,N_4103,N_4077);
nor U4327 (N_4327,N_4144,N_4098);
xor U4328 (N_4328,N_4166,N_4160);
xor U4329 (N_4329,N_4020,N_4141);
nand U4330 (N_4330,N_4013,N_4126);
or U4331 (N_4331,N_4165,N_4106);
xor U4332 (N_4332,N_4171,N_4102);
xnor U4333 (N_4333,N_4107,N_4163);
or U4334 (N_4334,N_4014,N_4021);
nand U4335 (N_4335,N_4027,N_4108);
and U4336 (N_4336,N_4126,N_4079);
and U4337 (N_4337,N_4040,N_4104);
nand U4338 (N_4338,N_4153,N_4011);
nand U4339 (N_4339,N_4007,N_4185);
xor U4340 (N_4340,N_4011,N_4048);
xnor U4341 (N_4341,N_4106,N_4175);
and U4342 (N_4342,N_4136,N_4020);
or U4343 (N_4343,N_4048,N_4033);
and U4344 (N_4344,N_4185,N_4190);
nand U4345 (N_4345,N_4009,N_4089);
nor U4346 (N_4346,N_4106,N_4129);
nand U4347 (N_4347,N_4155,N_4083);
xnor U4348 (N_4348,N_4199,N_4090);
xor U4349 (N_4349,N_4009,N_4140);
nand U4350 (N_4350,N_4194,N_4153);
or U4351 (N_4351,N_4112,N_4183);
or U4352 (N_4352,N_4084,N_4083);
and U4353 (N_4353,N_4003,N_4005);
nand U4354 (N_4354,N_4053,N_4068);
nand U4355 (N_4355,N_4183,N_4181);
and U4356 (N_4356,N_4025,N_4014);
and U4357 (N_4357,N_4035,N_4122);
xor U4358 (N_4358,N_4081,N_4096);
nor U4359 (N_4359,N_4096,N_4049);
and U4360 (N_4360,N_4119,N_4019);
or U4361 (N_4361,N_4072,N_4136);
or U4362 (N_4362,N_4117,N_4164);
xnor U4363 (N_4363,N_4124,N_4079);
and U4364 (N_4364,N_4064,N_4094);
nor U4365 (N_4365,N_4057,N_4056);
xnor U4366 (N_4366,N_4145,N_4141);
nor U4367 (N_4367,N_4137,N_4140);
xor U4368 (N_4368,N_4185,N_4173);
nand U4369 (N_4369,N_4109,N_4158);
or U4370 (N_4370,N_4131,N_4048);
and U4371 (N_4371,N_4197,N_4081);
or U4372 (N_4372,N_4155,N_4135);
or U4373 (N_4373,N_4038,N_4081);
and U4374 (N_4374,N_4125,N_4061);
nand U4375 (N_4375,N_4174,N_4191);
nor U4376 (N_4376,N_4152,N_4108);
and U4377 (N_4377,N_4062,N_4123);
xor U4378 (N_4378,N_4068,N_4061);
or U4379 (N_4379,N_4158,N_4039);
nor U4380 (N_4380,N_4001,N_4147);
nand U4381 (N_4381,N_4014,N_4041);
nand U4382 (N_4382,N_4106,N_4131);
xnor U4383 (N_4383,N_4193,N_4156);
or U4384 (N_4384,N_4130,N_4177);
nand U4385 (N_4385,N_4011,N_4089);
or U4386 (N_4386,N_4179,N_4129);
nand U4387 (N_4387,N_4191,N_4020);
nor U4388 (N_4388,N_4054,N_4167);
or U4389 (N_4389,N_4114,N_4056);
nor U4390 (N_4390,N_4054,N_4060);
and U4391 (N_4391,N_4106,N_4113);
nor U4392 (N_4392,N_4196,N_4085);
nor U4393 (N_4393,N_4167,N_4023);
or U4394 (N_4394,N_4026,N_4044);
or U4395 (N_4395,N_4174,N_4018);
or U4396 (N_4396,N_4097,N_4016);
nor U4397 (N_4397,N_4128,N_4028);
nor U4398 (N_4398,N_4084,N_4196);
and U4399 (N_4399,N_4003,N_4118);
xnor U4400 (N_4400,N_4207,N_4206);
nand U4401 (N_4401,N_4249,N_4370);
xnor U4402 (N_4402,N_4326,N_4387);
and U4403 (N_4403,N_4311,N_4399);
nand U4404 (N_4404,N_4354,N_4313);
and U4405 (N_4405,N_4378,N_4367);
nand U4406 (N_4406,N_4369,N_4218);
and U4407 (N_4407,N_4352,N_4362);
nor U4408 (N_4408,N_4255,N_4364);
or U4409 (N_4409,N_4304,N_4295);
nor U4410 (N_4410,N_4355,N_4336);
nor U4411 (N_4411,N_4317,N_4358);
or U4412 (N_4412,N_4390,N_4333);
xor U4413 (N_4413,N_4238,N_4231);
nand U4414 (N_4414,N_4222,N_4217);
nor U4415 (N_4415,N_4240,N_4351);
and U4416 (N_4416,N_4323,N_4345);
nand U4417 (N_4417,N_4228,N_4381);
xor U4418 (N_4418,N_4346,N_4350);
xnor U4419 (N_4419,N_4303,N_4274);
nand U4420 (N_4420,N_4262,N_4359);
or U4421 (N_4421,N_4296,N_4357);
nor U4422 (N_4422,N_4300,N_4319);
or U4423 (N_4423,N_4276,N_4371);
nor U4424 (N_4424,N_4261,N_4325);
and U4425 (N_4425,N_4290,N_4223);
or U4426 (N_4426,N_4327,N_4385);
and U4427 (N_4427,N_4324,N_4334);
nor U4428 (N_4428,N_4375,N_4342);
xor U4429 (N_4429,N_4252,N_4271);
xnor U4430 (N_4430,N_4245,N_4329);
nand U4431 (N_4431,N_4281,N_4332);
and U4432 (N_4432,N_4353,N_4259);
and U4433 (N_4433,N_4395,N_4239);
xnor U4434 (N_4434,N_4205,N_4340);
nand U4435 (N_4435,N_4200,N_4339);
xnor U4436 (N_4436,N_4383,N_4384);
or U4437 (N_4437,N_4305,N_4224);
nor U4438 (N_4438,N_4308,N_4373);
nor U4439 (N_4439,N_4256,N_4212);
nor U4440 (N_4440,N_4275,N_4204);
or U4441 (N_4441,N_4368,N_4283);
or U4442 (N_4442,N_4363,N_4312);
nor U4443 (N_4443,N_4388,N_4232);
and U4444 (N_4444,N_4243,N_4341);
and U4445 (N_4445,N_4277,N_4233);
or U4446 (N_4446,N_4246,N_4316);
and U4447 (N_4447,N_4338,N_4251);
nand U4448 (N_4448,N_4309,N_4314);
or U4449 (N_4449,N_4310,N_4297);
or U4450 (N_4450,N_4210,N_4229);
and U4451 (N_4451,N_4285,N_4214);
or U4452 (N_4452,N_4216,N_4289);
nor U4453 (N_4453,N_4230,N_4299);
xor U4454 (N_4454,N_4237,N_4248);
or U4455 (N_4455,N_4382,N_4268);
xnor U4456 (N_4456,N_4272,N_4318);
or U4457 (N_4457,N_4202,N_4322);
nor U4458 (N_4458,N_4293,N_4306);
or U4459 (N_4459,N_4365,N_4220);
nor U4460 (N_4460,N_4307,N_4288);
nor U4461 (N_4461,N_4344,N_4227);
xnor U4462 (N_4462,N_4208,N_4267);
or U4463 (N_4463,N_4225,N_4349);
or U4464 (N_4464,N_4389,N_4392);
and U4465 (N_4465,N_4376,N_4221);
or U4466 (N_4466,N_4379,N_4377);
nor U4467 (N_4467,N_4247,N_4374);
nand U4468 (N_4468,N_4253,N_4291);
xnor U4469 (N_4469,N_4366,N_4279);
or U4470 (N_4470,N_4215,N_4337);
or U4471 (N_4471,N_4330,N_4254);
nor U4472 (N_4472,N_4282,N_4284);
xor U4473 (N_4473,N_4236,N_4328);
nor U4474 (N_4474,N_4396,N_4235);
xor U4475 (N_4475,N_4302,N_4294);
xor U4476 (N_4476,N_4356,N_4241);
or U4477 (N_4477,N_4391,N_4260);
xor U4478 (N_4478,N_4331,N_4360);
or U4479 (N_4479,N_4213,N_4372);
or U4480 (N_4480,N_4219,N_4301);
and U4481 (N_4481,N_4266,N_4386);
nor U4482 (N_4482,N_4263,N_4280);
xnor U4483 (N_4483,N_4380,N_4250);
nand U4484 (N_4484,N_4278,N_4394);
and U4485 (N_4485,N_4320,N_4201);
xor U4486 (N_4486,N_4286,N_4315);
nand U4487 (N_4487,N_4244,N_4211);
nor U4488 (N_4488,N_4203,N_4335);
xnor U4489 (N_4489,N_4257,N_4393);
nand U4490 (N_4490,N_4347,N_4398);
xor U4491 (N_4491,N_4361,N_4209);
nor U4492 (N_4492,N_4273,N_4397);
or U4493 (N_4493,N_4242,N_4265);
nor U4494 (N_4494,N_4321,N_4343);
or U4495 (N_4495,N_4258,N_4269);
and U4496 (N_4496,N_4292,N_4234);
xnor U4497 (N_4497,N_4348,N_4270);
or U4498 (N_4498,N_4264,N_4298);
xor U4499 (N_4499,N_4287,N_4226);
nor U4500 (N_4500,N_4315,N_4247);
xnor U4501 (N_4501,N_4254,N_4234);
xnor U4502 (N_4502,N_4361,N_4277);
nand U4503 (N_4503,N_4227,N_4210);
nand U4504 (N_4504,N_4345,N_4339);
nand U4505 (N_4505,N_4368,N_4371);
nand U4506 (N_4506,N_4269,N_4250);
and U4507 (N_4507,N_4302,N_4254);
and U4508 (N_4508,N_4345,N_4266);
and U4509 (N_4509,N_4262,N_4300);
nor U4510 (N_4510,N_4275,N_4216);
or U4511 (N_4511,N_4228,N_4336);
nand U4512 (N_4512,N_4309,N_4334);
nand U4513 (N_4513,N_4278,N_4384);
xor U4514 (N_4514,N_4204,N_4362);
nand U4515 (N_4515,N_4388,N_4375);
or U4516 (N_4516,N_4296,N_4333);
or U4517 (N_4517,N_4328,N_4343);
or U4518 (N_4518,N_4209,N_4232);
or U4519 (N_4519,N_4302,N_4390);
nor U4520 (N_4520,N_4209,N_4380);
xnor U4521 (N_4521,N_4256,N_4306);
and U4522 (N_4522,N_4382,N_4295);
nand U4523 (N_4523,N_4386,N_4247);
and U4524 (N_4524,N_4332,N_4322);
and U4525 (N_4525,N_4213,N_4308);
xnor U4526 (N_4526,N_4218,N_4265);
nand U4527 (N_4527,N_4314,N_4297);
nor U4528 (N_4528,N_4213,N_4361);
xor U4529 (N_4529,N_4274,N_4397);
nand U4530 (N_4530,N_4218,N_4296);
xor U4531 (N_4531,N_4299,N_4324);
and U4532 (N_4532,N_4244,N_4330);
nor U4533 (N_4533,N_4234,N_4219);
nor U4534 (N_4534,N_4271,N_4242);
and U4535 (N_4535,N_4218,N_4293);
nor U4536 (N_4536,N_4346,N_4223);
nor U4537 (N_4537,N_4246,N_4248);
nand U4538 (N_4538,N_4219,N_4286);
xor U4539 (N_4539,N_4325,N_4260);
nor U4540 (N_4540,N_4246,N_4380);
and U4541 (N_4541,N_4384,N_4271);
or U4542 (N_4542,N_4283,N_4265);
and U4543 (N_4543,N_4304,N_4307);
or U4544 (N_4544,N_4281,N_4354);
nand U4545 (N_4545,N_4377,N_4368);
nor U4546 (N_4546,N_4261,N_4397);
nand U4547 (N_4547,N_4359,N_4202);
nor U4548 (N_4548,N_4201,N_4306);
and U4549 (N_4549,N_4362,N_4294);
nand U4550 (N_4550,N_4374,N_4342);
nor U4551 (N_4551,N_4260,N_4266);
nand U4552 (N_4552,N_4250,N_4356);
nor U4553 (N_4553,N_4246,N_4313);
nand U4554 (N_4554,N_4292,N_4315);
and U4555 (N_4555,N_4267,N_4206);
nand U4556 (N_4556,N_4366,N_4313);
and U4557 (N_4557,N_4286,N_4221);
xor U4558 (N_4558,N_4242,N_4279);
and U4559 (N_4559,N_4311,N_4381);
xor U4560 (N_4560,N_4211,N_4376);
nor U4561 (N_4561,N_4373,N_4312);
xnor U4562 (N_4562,N_4315,N_4323);
nor U4563 (N_4563,N_4305,N_4207);
or U4564 (N_4564,N_4373,N_4387);
or U4565 (N_4565,N_4298,N_4220);
nor U4566 (N_4566,N_4247,N_4307);
or U4567 (N_4567,N_4322,N_4278);
nor U4568 (N_4568,N_4202,N_4366);
and U4569 (N_4569,N_4318,N_4235);
and U4570 (N_4570,N_4306,N_4228);
nand U4571 (N_4571,N_4392,N_4261);
and U4572 (N_4572,N_4387,N_4383);
nor U4573 (N_4573,N_4399,N_4273);
xnor U4574 (N_4574,N_4311,N_4284);
nor U4575 (N_4575,N_4393,N_4317);
or U4576 (N_4576,N_4362,N_4304);
and U4577 (N_4577,N_4307,N_4372);
nor U4578 (N_4578,N_4341,N_4330);
or U4579 (N_4579,N_4226,N_4288);
and U4580 (N_4580,N_4354,N_4330);
nor U4581 (N_4581,N_4310,N_4329);
or U4582 (N_4582,N_4254,N_4391);
nor U4583 (N_4583,N_4325,N_4359);
nand U4584 (N_4584,N_4245,N_4217);
and U4585 (N_4585,N_4397,N_4370);
or U4586 (N_4586,N_4297,N_4350);
nand U4587 (N_4587,N_4265,N_4353);
xor U4588 (N_4588,N_4237,N_4268);
and U4589 (N_4589,N_4230,N_4246);
nor U4590 (N_4590,N_4263,N_4264);
or U4591 (N_4591,N_4376,N_4329);
nor U4592 (N_4592,N_4311,N_4325);
xnor U4593 (N_4593,N_4253,N_4350);
nand U4594 (N_4594,N_4338,N_4325);
nand U4595 (N_4595,N_4357,N_4395);
and U4596 (N_4596,N_4291,N_4396);
nor U4597 (N_4597,N_4207,N_4297);
or U4598 (N_4598,N_4208,N_4399);
nand U4599 (N_4599,N_4233,N_4231);
nor U4600 (N_4600,N_4509,N_4491);
or U4601 (N_4601,N_4436,N_4589);
nor U4602 (N_4602,N_4561,N_4588);
and U4603 (N_4603,N_4575,N_4478);
nand U4604 (N_4604,N_4531,N_4407);
xor U4605 (N_4605,N_4424,N_4429);
nor U4606 (N_4606,N_4423,N_4455);
xnor U4607 (N_4607,N_4517,N_4581);
and U4608 (N_4608,N_4500,N_4524);
nand U4609 (N_4609,N_4578,N_4579);
xor U4610 (N_4610,N_4598,N_4415);
or U4611 (N_4611,N_4454,N_4456);
nor U4612 (N_4612,N_4545,N_4583);
or U4613 (N_4613,N_4433,N_4582);
nand U4614 (N_4614,N_4514,N_4551);
nand U4615 (N_4615,N_4483,N_4550);
and U4616 (N_4616,N_4472,N_4526);
nor U4617 (N_4617,N_4417,N_4449);
and U4618 (N_4618,N_4493,N_4492);
or U4619 (N_4619,N_4430,N_4494);
or U4620 (N_4620,N_4566,N_4549);
xor U4621 (N_4621,N_4554,N_4422);
or U4622 (N_4622,N_4595,N_4539);
nand U4623 (N_4623,N_4504,N_4489);
nand U4624 (N_4624,N_4507,N_4591);
xnor U4625 (N_4625,N_4568,N_4442);
and U4626 (N_4626,N_4497,N_4486);
xor U4627 (N_4627,N_4406,N_4419);
xnor U4628 (N_4628,N_4576,N_4401);
or U4629 (N_4629,N_4558,N_4488);
and U4630 (N_4630,N_4434,N_4470);
nand U4631 (N_4631,N_4599,N_4452);
xnor U4632 (N_4632,N_4428,N_4469);
or U4633 (N_4633,N_4503,N_4559);
or U4634 (N_4634,N_4577,N_4527);
or U4635 (N_4635,N_4462,N_4446);
or U4636 (N_4636,N_4404,N_4438);
xnor U4637 (N_4637,N_4521,N_4516);
nor U4638 (N_4638,N_4444,N_4465);
nor U4639 (N_4639,N_4510,N_4515);
nand U4640 (N_4640,N_4416,N_4587);
or U4641 (N_4641,N_4513,N_4410);
nor U4642 (N_4642,N_4480,N_4445);
nand U4643 (N_4643,N_4400,N_4467);
and U4644 (N_4644,N_4475,N_4567);
nand U4645 (N_4645,N_4443,N_4542);
nor U4646 (N_4646,N_4411,N_4511);
nand U4647 (N_4647,N_4448,N_4570);
and U4648 (N_4648,N_4490,N_4560);
and U4649 (N_4649,N_4530,N_4519);
nor U4650 (N_4650,N_4476,N_4590);
and U4651 (N_4651,N_4565,N_4474);
xnor U4652 (N_4652,N_4528,N_4569);
nor U4653 (N_4653,N_4414,N_4453);
nor U4654 (N_4654,N_4541,N_4537);
nand U4655 (N_4655,N_4440,N_4501);
or U4656 (N_4656,N_4502,N_4512);
or U4657 (N_4657,N_4425,N_4466);
nor U4658 (N_4658,N_4482,N_4518);
nand U4659 (N_4659,N_4538,N_4557);
nand U4660 (N_4660,N_4437,N_4413);
and U4661 (N_4661,N_4552,N_4457);
nand U4662 (N_4662,N_4555,N_4597);
nor U4663 (N_4663,N_4523,N_4572);
and U4664 (N_4664,N_4409,N_4594);
nand U4665 (N_4665,N_4471,N_4548);
nand U4666 (N_4666,N_4525,N_4468);
xor U4667 (N_4667,N_4562,N_4499);
nor U4668 (N_4668,N_4460,N_4584);
xor U4669 (N_4669,N_4459,N_4573);
or U4670 (N_4670,N_4431,N_4458);
and U4671 (N_4671,N_4418,N_4580);
nand U4672 (N_4672,N_4571,N_4403);
or U4673 (N_4673,N_4544,N_4479);
xnor U4674 (N_4674,N_4447,N_4574);
nand U4675 (N_4675,N_4427,N_4432);
nor U4676 (N_4676,N_4435,N_4543);
xnor U4677 (N_4677,N_4534,N_4596);
nand U4678 (N_4678,N_4451,N_4473);
or U4679 (N_4679,N_4498,N_4420);
and U4680 (N_4680,N_4464,N_4463);
xnor U4681 (N_4681,N_4495,N_4533);
nand U4682 (N_4682,N_4520,N_4535);
nand U4683 (N_4683,N_4402,N_4553);
and U4684 (N_4684,N_4484,N_4461);
and U4685 (N_4685,N_4506,N_4586);
xnor U4686 (N_4686,N_4405,N_4505);
and U4687 (N_4687,N_4546,N_4477);
or U4688 (N_4688,N_4485,N_4540);
and U4689 (N_4689,N_4585,N_4426);
xnor U4690 (N_4690,N_4564,N_4481);
nand U4691 (N_4691,N_4421,N_4496);
xor U4692 (N_4692,N_4439,N_4522);
or U4693 (N_4693,N_4529,N_4593);
or U4694 (N_4694,N_4563,N_4532);
xor U4695 (N_4695,N_4547,N_4508);
nand U4696 (N_4696,N_4487,N_4408);
nand U4697 (N_4697,N_4536,N_4556);
or U4698 (N_4698,N_4441,N_4592);
and U4699 (N_4699,N_4412,N_4450);
and U4700 (N_4700,N_4548,N_4404);
nand U4701 (N_4701,N_4558,N_4469);
or U4702 (N_4702,N_4431,N_4546);
xor U4703 (N_4703,N_4438,N_4502);
or U4704 (N_4704,N_4511,N_4499);
xnor U4705 (N_4705,N_4491,N_4413);
nor U4706 (N_4706,N_4422,N_4537);
nor U4707 (N_4707,N_4480,N_4494);
nand U4708 (N_4708,N_4583,N_4549);
nor U4709 (N_4709,N_4493,N_4418);
nand U4710 (N_4710,N_4474,N_4427);
nor U4711 (N_4711,N_4413,N_4532);
nor U4712 (N_4712,N_4431,N_4521);
xnor U4713 (N_4713,N_4575,N_4491);
and U4714 (N_4714,N_4460,N_4504);
nor U4715 (N_4715,N_4464,N_4527);
xnor U4716 (N_4716,N_4423,N_4404);
nor U4717 (N_4717,N_4404,N_4571);
and U4718 (N_4718,N_4528,N_4411);
and U4719 (N_4719,N_4480,N_4479);
and U4720 (N_4720,N_4479,N_4505);
xor U4721 (N_4721,N_4517,N_4441);
nand U4722 (N_4722,N_4485,N_4484);
xnor U4723 (N_4723,N_4534,N_4478);
xnor U4724 (N_4724,N_4487,N_4519);
xnor U4725 (N_4725,N_4499,N_4510);
nand U4726 (N_4726,N_4460,N_4593);
and U4727 (N_4727,N_4547,N_4451);
nand U4728 (N_4728,N_4577,N_4572);
xor U4729 (N_4729,N_4503,N_4419);
xnor U4730 (N_4730,N_4439,N_4571);
and U4731 (N_4731,N_4524,N_4481);
nor U4732 (N_4732,N_4498,N_4526);
nand U4733 (N_4733,N_4506,N_4548);
or U4734 (N_4734,N_4548,N_4421);
nor U4735 (N_4735,N_4548,N_4452);
nand U4736 (N_4736,N_4419,N_4570);
or U4737 (N_4737,N_4562,N_4418);
or U4738 (N_4738,N_4452,N_4514);
and U4739 (N_4739,N_4449,N_4409);
and U4740 (N_4740,N_4588,N_4568);
nor U4741 (N_4741,N_4572,N_4443);
or U4742 (N_4742,N_4572,N_4436);
nand U4743 (N_4743,N_4428,N_4453);
or U4744 (N_4744,N_4480,N_4450);
nand U4745 (N_4745,N_4460,N_4552);
nor U4746 (N_4746,N_4594,N_4599);
or U4747 (N_4747,N_4579,N_4511);
or U4748 (N_4748,N_4596,N_4468);
or U4749 (N_4749,N_4578,N_4525);
or U4750 (N_4750,N_4571,N_4460);
nor U4751 (N_4751,N_4439,N_4529);
nor U4752 (N_4752,N_4458,N_4401);
nand U4753 (N_4753,N_4458,N_4553);
or U4754 (N_4754,N_4595,N_4434);
or U4755 (N_4755,N_4517,N_4425);
xor U4756 (N_4756,N_4498,N_4408);
nand U4757 (N_4757,N_4463,N_4493);
or U4758 (N_4758,N_4411,N_4558);
nand U4759 (N_4759,N_4404,N_4541);
or U4760 (N_4760,N_4553,N_4534);
nor U4761 (N_4761,N_4440,N_4586);
xnor U4762 (N_4762,N_4475,N_4427);
nand U4763 (N_4763,N_4429,N_4577);
or U4764 (N_4764,N_4483,N_4553);
or U4765 (N_4765,N_4424,N_4413);
xnor U4766 (N_4766,N_4583,N_4547);
nor U4767 (N_4767,N_4435,N_4497);
or U4768 (N_4768,N_4570,N_4503);
xnor U4769 (N_4769,N_4477,N_4595);
and U4770 (N_4770,N_4429,N_4422);
and U4771 (N_4771,N_4558,N_4413);
nand U4772 (N_4772,N_4419,N_4444);
or U4773 (N_4773,N_4488,N_4469);
nand U4774 (N_4774,N_4457,N_4405);
or U4775 (N_4775,N_4432,N_4440);
nand U4776 (N_4776,N_4430,N_4464);
or U4777 (N_4777,N_4511,N_4557);
xor U4778 (N_4778,N_4511,N_4471);
and U4779 (N_4779,N_4452,N_4563);
or U4780 (N_4780,N_4465,N_4437);
nand U4781 (N_4781,N_4479,N_4489);
and U4782 (N_4782,N_4559,N_4501);
and U4783 (N_4783,N_4402,N_4480);
or U4784 (N_4784,N_4565,N_4514);
or U4785 (N_4785,N_4427,N_4454);
and U4786 (N_4786,N_4511,N_4596);
or U4787 (N_4787,N_4464,N_4461);
nand U4788 (N_4788,N_4480,N_4544);
nor U4789 (N_4789,N_4511,N_4419);
xnor U4790 (N_4790,N_4458,N_4413);
xnor U4791 (N_4791,N_4408,N_4476);
nand U4792 (N_4792,N_4497,N_4587);
or U4793 (N_4793,N_4528,N_4473);
nand U4794 (N_4794,N_4593,N_4530);
xor U4795 (N_4795,N_4520,N_4589);
and U4796 (N_4796,N_4472,N_4491);
xnor U4797 (N_4797,N_4404,N_4476);
or U4798 (N_4798,N_4450,N_4421);
xnor U4799 (N_4799,N_4410,N_4407);
and U4800 (N_4800,N_4618,N_4713);
nand U4801 (N_4801,N_4630,N_4660);
nand U4802 (N_4802,N_4700,N_4645);
and U4803 (N_4803,N_4730,N_4725);
xnor U4804 (N_4804,N_4624,N_4726);
and U4805 (N_4805,N_4667,N_4600);
xor U4806 (N_4806,N_4631,N_4751);
xnor U4807 (N_4807,N_4762,N_4737);
and U4808 (N_4808,N_4634,N_4721);
or U4809 (N_4809,N_4633,N_4680);
or U4810 (N_4810,N_4778,N_4642);
xnor U4811 (N_4811,N_4682,N_4668);
nand U4812 (N_4812,N_4761,N_4720);
nand U4813 (N_4813,N_4698,N_4678);
nor U4814 (N_4814,N_4671,N_4753);
xor U4815 (N_4815,N_4729,N_4641);
or U4816 (N_4816,N_4752,N_4677);
or U4817 (N_4817,N_4657,N_4654);
or U4818 (N_4818,N_4760,N_4676);
xor U4819 (N_4819,N_4664,N_4627);
nand U4820 (N_4820,N_4644,N_4786);
xnor U4821 (N_4821,N_4782,N_4665);
or U4822 (N_4822,N_4690,N_4775);
nor U4823 (N_4823,N_4614,N_4735);
nor U4824 (N_4824,N_4792,N_4767);
and U4825 (N_4825,N_4727,N_4679);
and U4826 (N_4826,N_4717,N_4758);
or U4827 (N_4827,N_4702,N_4647);
xor U4828 (N_4828,N_4691,N_4709);
xnor U4829 (N_4829,N_4621,N_4636);
and U4830 (N_4830,N_4773,N_4797);
nor U4831 (N_4831,N_4711,N_4777);
and U4832 (N_4832,N_4731,N_4639);
nand U4833 (N_4833,N_4609,N_4683);
nand U4834 (N_4834,N_4707,N_4756);
nor U4835 (N_4835,N_4620,N_4705);
nand U4836 (N_4836,N_4781,N_4744);
nor U4837 (N_4837,N_4776,N_4672);
and U4838 (N_4838,N_4670,N_4622);
and U4839 (N_4839,N_4673,N_4794);
and U4840 (N_4840,N_4694,N_4685);
or U4841 (N_4841,N_4712,N_4610);
xor U4842 (N_4842,N_4728,N_4750);
nor U4843 (N_4843,N_4789,N_4611);
xor U4844 (N_4844,N_4790,N_4669);
and U4845 (N_4845,N_4710,N_4708);
or U4846 (N_4846,N_4687,N_4653);
and U4847 (N_4847,N_4625,N_4798);
nand U4848 (N_4848,N_4719,N_4770);
or U4849 (N_4849,N_4604,N_4733);
or U4850 (N_4850,N_4732,N_4774);
and U4851 (N_4851,N_4605,N_4616);
and U4852 (N_4852,N_4745,N_4764);
xor U4853 (N_4853,N_4799,N_4615);
nor U4854 (N_4854,N_4619,N_4689);
nand U4855 (N_4855,N_4637,N_4638);
nor U4856 (N_4856,N_4701,N_4791);
nor U4857 (N_4857,N_4697,N_4628);
and U4858 (N_4858,N_4715,N_4606);
nor U4859 (N_4859,N_4743,N_4724);
nor U4860 (N_4860,N_4795,N_4649);
or U4861 (N_4861,N_4771,N_4612);
and U4862 (N_4862,N_4688,N_4646);
nand U4863 (N_4863,N_4716,N_4693);
nand U4864 (N_4864,N_4659,N_4740);
or U4865 (N_4865,N_4703,N_4662);
or U4866 (N_4866,N_4635,N_4632);
nor U4867 (N_4867,N_4757,N_4796);
or U4868 (N_4868,N_4656,N_4602);
and U4869 (N_4869,N_4759,N_4772);
nor U4870 (N_4870,N_4617,N_4755);
and U4871 (N_4871,N_4736,N_4648);
nand U4872 (N_4872,N_4746,N_4613);
nand U4873 (N_4873,N_4788,N_4629);
or U4874 (N_4874,N_4784,N_4748);
and U4875 (N_4875,N_4655,N_4658);
or U4876 (N_4876,N_4608,N_4674);
and U4877 (N_4877,N_4651,N_4692);
or U4878 (N_4878,N_4603,N_4706);
and U4879 (N_4879,N_4783,N_4779);
nor U4880 (N_4880,N_4763,N_4623);
and U4881 (N_4881,N_4686,N_4643);
xnor U4882 (N_4882,N_4765,N_4601);
nand U4883 (N_4883,N_4769,N_4704);
nor U4884 (N_4884,N_4661,N_4699);
and U4885 (N_4885,N_4734,N_4747);
nor U4886 (N_4886,N_4780,N_4766);
and U4887 (N_4887,N_4793,N_4607);
and U4888 (N_4888,N_4741,N_4768);
nor U4889 (N_4889,N_4754,N_4640);
nand U4890 (N_4890,N_4652,N_4675);
nor U4891 (N_4891,N_4684,N_4749);
or U4892 (N_4892,N_4787,N_4714);
xnor U4893 (N_4893,N_4666,N_4739);
xnor U4894 (N_4894,N_4663,N_4718);
nand U4895 (N_4895,N_4738,N_4723);
xnor U4896 (N_4896,N_4785,N_4696);
xor U4897 (N_4897,N_4681,N_4742);
nand U4898 (N_4898,N_4626,N_4650);
xnor U4899 (N_4899,N_4695,N_4722);
nand U4900 (N_4900,N_4701,N_4695);
nor U4901 (N_4901,N_4685,N_4710);
nand U4902 (N_4902,N_4639,N_4765);
and U4903 (N_4903,N_4793,N_4685);
or U4904 (N_4904,N_4673,N_4773);
nor U4905 (N_4905,N_4678,N_4663);
nand U4906 (N_4906,N_4608,N_4751);
and U4907 (N_4907,N_4692,N_4665);
and U4908 (N_4908,N_4643,N_4618);
nand U4909 (N_4909,N_4780,N_4773);
or U4910 (N_4910,N_4606,N_4662);
and U4911 (N_4911,N_4622,N_4665);
nor U4912 (N_4912,N_4730,N_4652);
and U4913 (N_4913,N_4671,N_4622);
or U4914 (N_4914,N_4716,N_4779);
nand U4915 (N_4915,N_4667,N_4657);
nand U4916 (N_4916,N_4679,N_4728);
nor U4917 (N_4917,N_4624,N_4707);
xnor U4918 (N_4918,N_4778,N_4789);
nand U4919 (N_4919,N_4650,N_4794);
xnor U4920 (N_4920,N_4707,N_4731);
nor U4921 (N_4921,N_4678,N_4649);
and U4922 (N_4922,N_4636,N_4617);
or U4923 (N_4923,N_4710,N_4729);
or U4924 (N_4924,N_4735,N_4771);
nor U4925 (N_4925,N_4793,N_4791);
xor U4926 (N_4926,N_4757,N_4635);
and U4927 (N_4927,N_4703,N_4645);
and U4928 (N_4928,N_4690,N_4606);
nand U4929 (N_4929,N_4727,N_4640);
xor U4930 (N_4930,N_4658,N_4742);
nand U4931 (N_4931,N_4749,N_4611);
nor U4932 (N_4932,N_4795,N_4762);
nand U4933 (N_4933,N_4760,N_4777);
nand U4934 (N_4934,N_4651,N_4789);
xor U4935 (N_4935,N_4786,N_4774);
and U4936 (N_4936,N_4712,N_4609);
xor U4937 (N_4937,N_4663,N_4632);
and U4938 (N_4938,N_4627,N_4656);
and U4939 (N_4939,N_4775,N_4790);
nor U4940 (N_4940,N_4750,N_4684);
nor U4941 (N_4941,N_4763,N_4667);
or U4942 (N_4942,N_4748,N_4680);
xor U4943 (N_4943,N_4648,N_4663);
nand U4944 (N_4944,N_4656,N_4703);
nand U4945 (N_4945,N_4606,N_4604);
xnor U4946 (N_4946,N_4774,N_4684);
or U4947 (N_4947,N_4702,N_4632);
nor U4948 (N_4948,N_4602,N_4743);
nor U4949 (N_4949,N_4796,N_4635);
or U4950 (N_4950,N_4785,N_4719);
and U4951 (N_4951,N_4607,N_4623);
nand U4952 (N_4952,N_4620,N_4689);
xor U4953 (N_4953,N_4647,N_4694);
xnor U4954 (N_4954,N_4791,N_4617);
xor U4955 (N_4955,N_4600,N_4627);
or U4956 (N_4956,N_4739,N_4660);
nor U4957 (N_4957,N_4760,N_4690);
nand U4958 (N_4958,N_4615,N_4722);
or U4959 (N_4959,N_4640,N_4621);
and U4960 (N_4960,N_4710,N_4622);
nand U4961 (N_4961,N_4767,N_4709);
nand U4962 (N_4962,N_4753,N_4746);
nand U4963 (N_4963,N_4648,N_4796);
nor U4964 (N_4964,N_4727,N_4623);
or U4965 (N_4965,N_4753,N_4787);
nor U4966 (N_4966,N_4673,N_4756);
xor U4967 (N_4967,N_4678,N_4780);
nor U4968 (N_4968,N_4615,N_4612);
nor U4969 (N_4969,N_4735,N_4794);
nor U4970 (N_4970,N_4675,N_4761);
xor U4971 (N_4971,N_4645,N_4760);
nand U4972 (N_4972,N_4772,N_4688);
and U4973 (N_4973,N_4703,N_4799);
xor U4974 (N_4974,N_4692,N_4608);
or U4975 (N_4975,N_4658,N_4657);
xor U4976 (N_4976,N_4727,N_4697);
xnor U4977 (N_4977,N_4685,N_4739);
nor U4978 (N_4978,N_4705,N_4612);
xor U4979 (N_4979,N_4760,N_4620);
xnor U4980 (N_4980,N_4789,N_4698);
or U4981 (N_4981,N_4772,N_4620);
or U4982 (N_4982,N_4778,N_4775);
nand U4983 (N_4983,N_4754,N_4783);
and U4984 (N_4984,N_4682,N_4761);
nor U4985 (N_4985,N_4653,N_4753);
nand U4986 (N_4986,N_4798,N_4715);
xor U4987 (N_4987,N_4604,N_4776);
xnor U4988 (N_4988,N_4700,N_4751);
xnor U4989 (N_4989,N_4629,N_4785);
xor U4990 (N_4990,N_4601,N_4738);
or U4991 (N_4991,N_4617,N_4734);
xor U4992 (N_4992,N_4642,N_4693);
and U4993 (N_4993,N_4641,N_4618);
nor U4994 (N_4994,N_4676,N_4652);
nor U4995 (N_4995,N_4660,N_4618);
nor U4996 (N_4996,N_4735,N_4799);
or U4997 (N_4997,N_4695,N_4625);
and U4998 (N_4998,N_4637,N_4625);
nor U4999 (N_4999,N_4655,N_4757);
and UO_0 (O_0,N_4942,N_4936);
xnor UO_1 (O_1,N_4940,N_4812);
xor UO_2 (O_2,N_4938,N_4918);
nand UO_3 (O_3,N_4872,N_4935);
xor UO_4 (O_4,N_4819,N_4976);
nor UO_5 (O_5,N_4882,N_4852);
and UO_6 (O_6,N_4966,N_4922);
and UO_7 (O_7,N_4848,N_4906);
nand UO_8 (O_8,N_4865,N_4818);
nand UO_9 (O_9,N_4822,N_4801);
nand UO_10 (O_10,N_4899,N_4989);
nor UO_11 (O_11,N_4866,N_4917);
and UO_12 (O_12,N_4894,N_4914);
nor UO_13 (O_13,N_4953,N_4971);
or UO_14 (O_14,N_4880,N_4910);
nand UO_15 (O_15,N_4999,N_4802);
or UO_16 (O_16,N_4877,N_4944);
nor UO_17 (O_17,N_4887,N_4920);
xor UO_18 (O_18,N_4932,N_4820);
nor UO_19 (O_19,N_4827,N_4842);
nor UO_20 (O_20,N_4916,N_4998);
xor UO_21 (O_21,N_4980,N_4851);
and UO_22 (O_22,N_4909,N_4832);
xor UO_23 (O_23,N_4839,N_4809);
nor UO_24 (O_24,N_4869,N_4881);
nand UO_25 (O_25,N_4965,N_4968);
nor UO_26 (O_26,N_4883,N_4833);
xor UO_27 (O_27,N_4817,N_4987);
or UO_28 (O_28,N_4943,N_4805);
nand UO_29 (O_29,N_4874,N_4908);
nand UO_30 (O_30,N_4905,N_4950);
and UO_31 (O_31,N_4859,N_4947);
xnor UO_32 (O_32,N_4836,N_4855);
nand UO_33 (O_33,N_4939,N_4838);
xnor UO_34 (O_34,N_4961,N_4853);
nand UO_35 (O_35,N_4896,N_4810);
nand UO_36 (O_36,N_4901,N_4867);
xnor UO_37 (O_37,N_4862,N_4983);
xor UO_38 (O_38,N_4902,N_4997);
nand UO_39 (O_39,N_4926,N_4927);
and UO_40 (O_40,N_4915,N_4956);
and UO_41 (O_41,N_4890,N_4856);
nand UO_42 (O_42,N_4973,N_4959);
nor UO_43 (O_43,N_4892,N_4904);
nor UO_44 (O_44,N_4990,N_4845);
or UO_45 (O_45,N_4975,N_4811);
nor UO_46 (O_46,N_4854,N_4834);
nor UO_47 (O_47,N_4807,N_4829);
xnor UO_48 (O_48,N_4945,N_4974);
nor UO_49 (O_49,N_4824,N_4954);
nand UO_50 (O_50,N_4982,N_4955);
or UO_51 (O_51,N_4925,N_4849);
or UO_52 (O_52,N_4930,N_4952);
xnor UO_53 (O_53,N_4913,N_4825);
xnor UO_54 (O_54,N_4841,N_4941);
xnor UO_55 (O_55,N_4995,N_4847);
nor UO_56 (O_56,N_4868,N_4876);
nand UO_57 (O_57,N_4803,N_4857);
nor UO_58 (O_58,N_4900,N_4804);
and UO_59 (O_59,N_4919,N_4814);
or UO_60 (O_60,N_4821,N_4889);
nor UO_61 (O_61,N_4994,N_4813);
or UO_62 (O_62,N_4957,N_4948);
and UO_63 (O_63,N_4937,N_4970);
and UO_64 (O_64,N_4873,N_4985);
xnor UO_65 (O_65,N_4823,N_4963);
nor UO_66 (O_66,N_4981,N_4806);
or UO_67 (O_67,N_4992,N_4893);
xnor UO_68 (O_68,N_4984,N_4891);
nand UO_69 (O_69,N_4993,N_4870);
and UO_70 (O_70,N_4960,N_4837);
xnor UO_71 (O_71,N_4949,N_4898);
or UO_72 (O_72,N_4986,N_4969);
or UO_73 (O_73,N_4991,N_4886);
or UO_74 (O_74,N_4929,N_4879);
xor UO_75 (O_75,N_4861,N_4967);
nor UO_76 (O_76,N_4988,N_4924);
and UO_77 (O_77,N_4828,N_4931);
nor UO_78 (O_78,N_4850,N_4885);
xnor UO_79 (O_79,N_4878,N_4831);
or UO_80 (O_80,N_4840,N_4815);
or UO_81 (O_81,N_4972,N_4912);
and UO_82 (O_82,N_4844,N_4977);
and UO_83 (O_83,N_4826,N_4903);
or UO_84 (O_84,N_4933,N_4934);
or UO_85 (O_85,N_4846,N_4962);
xor UO_86 (O_86,N_4907,N_4863);
nor UO_87 (O_87,N_4923,N_4808);
or UO_88 (O_88,N_4843,N_4816);
nand UO_89 (O_89,N_4858,N_4911);
nand UO_90 (O_90,N_4921,N_4875);
or UO_91 (O_91,N_4964,N_4884);
nand UO_92 (O_92,N_4996,N_4897);
nor UO_93 (O_93,N_4860,N_4800);
nand UO_94 (O_94,N_4864,N_4951);
nand UO_95 (O_95,N_4835,N_4946);
nand UO_96 (O_96,N_4978,N_4895);
and UO_97 (O_97,N_4958,N_4888);
or UO_98 (O_98,N_4871,N_4830);
and UO_99 (O_99,N_4928,N_4979);
xor UO_100 (O_100,N_4974,N_4802);
xnor UO_101 (O_101,N_4899,N_4856);
nand UO_102 (O_102,N_4864,N_4947);
or UO_103 (O_103,N_4882,N_4806);
or UO_104 (O_104,N_4821,N_4816);
nor UO_105 (O_105,N_4946,N_4878);
and UO_106 (O_106,N_4957,N_4908);
or UO_107 (O_107,N_4811,N_4852);
xor UO_108 (O_108,N_4908,N_4918);
xnor UO_109 (O_109,N_4935,N_4956);
xnor UO_110 (O_110,N_4820,N_4843);
or UO_111 (O_111,N_4922,N_4920);
xor UO_112 (O_112,N_4875,N_4977);
nand UO_113 (O_113,N_4968,N_4805);
nand UO_114 (O_114,N_4868,N_4950);
xnor UO_115 (O_115,N_4931,N_4803);
or UO_116 (O_116,N_4823,N_4881);
nor UO_117 (O_117,N_4924,N_4867);
or UO_118 (O_118,N_4873,N_4854);
nand UO_119 (O_119,N_4820,N_4819);
or UO_120 (O_120,N_4858,N_4959);
xnor UO_121 (O_121,N_4964,N_4934);
nand UO_122 (O_122,N_4912,N_4982);
xor UO_123 (O_123,N_4920,N_4878);
nand UO_124 (O_124,N_4867,N_4843);
xor UO_125 (O_125,N_4964,N_4863);
or UO_126 (O_126,N_4839,N_4992);
nor UO_127 (O_127,N_4848,N_4963);
xnor UO_128 (O_128,N_4913,N_4827);
or UO_129 (O_129,N_4877,N_4915);
nand UO_130 (O_130,N_4849,N_4964);
nor UO_131 (O_131,N_4914,N_4978);
nand UO_132 (O_132,N_4979,N_4943);
xor UO_133 (O_133,N_4817,N_4980);
xor UO_134 (O_134,N_4843,N_4991);
nand UO_135 (O_135,N_4832,N_4884);
nor UO_136 (O_136,N_4902,N_4848);
nand UO_137 (O_137,N_4853,N_4811);
and UO_138 (O_138,N_4803,N_4854);
or UO_139 (O_139,N_4867,N_4936);
xor UO_140 (O_140,N_4852,N_4851);
nand UO_141 (O_141,N_4932,N_4981);
xor UO_142 (O_142,N_4963,N_4810);
nor UO_143 (O_143,N_4823,N_4958);
nor UO_144 (O_144,N_4938,N_4975);
nand UO_145 (O_145,N_4986,N_4848);
xnor UO_146 (O_146,N_4897,N_4812);
xnor UO_147 (O_147,N_4947,N_4849);
nand UO_148 (O_148,N_4906,N_4902);
nand UO_149 (O_149,N_4982,N_4873);
nand UO_150 (O_150,N_4940,N_4998);
nand UO_151 (O_151,N_4862,N_4995);
or UO_152 (O_152,N_4828,N_4932);
xnor UO_153 (O_153,N_4880,N_4843);
nor UO_154 (O_154,N_4919,N_4833);
and UO_155 (O_155,N_4850,N_4809);
and UO_156 (O_156,N_4907,N_4801);
and UO_157 (O_157,N_4904,N_4964);
nand UO_158 (O_158,N_4817,N_4856);
nor UO_159 (O_159,N_4935,N_4998);
nand UO_160 (O_160,N_4820,N_4807);
and UO_161 (O_161,N_4937,N_4815);
or UO_162 (O_162,N_4917,N_4851);
and UO_163 (O_163,N_4831,N_4970);
and UO_164 (O_164,N_4932,N_4853);
xor UO_165 (O_165,N_4844,N_4813);
nor UO_166 (O_166,N_4889,N_4968);
nand UO_167 (O_167,N_4997,N_4842);
nand UO_168 (O_168,N_4845,N_4970);
xnor UO_169 (O_169,N_4878,N_4898);
or UO_170 (O_170,N_4837,N_4840);
nor UO_171 (O_171,N_4998,N_4992);
nor UO_172 (O_172,N_4913,N_4814);
or UO_173 (O_173,N_4952,N_4939);
xor UO_174 (O_174,N_4913,N_4844);
nor UO_175 (O_175,N_4967,N_4947);
nand UO_176 (O_176,N_4931,N_4865);
nand UO_177 (O_177,N_4964,N_4898);
and UO_178 (O_178,N_4958,N_4929);
nand UO_179 (O_179,N_4879,N_4808);
or UO_180 (O_180,N_4873,N_4924);
xnor UO_181 (O_181,N_4958,N_4963);
or UO_182 (O_182,N_4863,N_4870);
xor UO_183 (O_183,N_4921,N_4836);
or UO_184 (O_184,N_4998,N_4866);
and UO_185 (O_185,N_4979,N_4915);
nand UO_186 (O_186,N_4923,N_4961);
xor UO_187 (O_187,N_4836,N_4847);
nand UO_188 (O_188,N_4897,N_4963);
nor UO_189 (O_189,N_4924,N_4828);
or UO_190 (O_190,N_4971,N_4855);
nand UO_191 (O_191,N_4952,N_4979);
and UO_192 (O_192,N_4928,N_4872);
xnor UO_193 (O_193,N_4907,N_4920);
and UO_194 (O_194,N_4919,N_4921);
xnor UO_195 (O_195,N_4970,N_4841);
or UO_196 (O_196,N_4863,N_4899);
or UO_197 (O_197,N_4810,N_4859);
xnor UO_198 (O_198,N_4955,N_4864);
nor UO_199 (O_199,N_4951,N_4967);
and UO_200 (O_200,N_4803,N_4818);
nand UO_201 (O_201,N_4804,N_4816);
or UO_202 (O_202,N_4868,N_4872);
nand UO_203 (O_203,N_4825,N_4856);
xnor UO_204 (O_204,N_4870,N_4832);
xor UO_205 (O_205,N_4905,N_4846);
nor UO_206 (O_206,N_4954,N_4886);
nor UO_207 (O_207,N_4912,N_4842);
xnor UO_208 (O_208,N_4935,N_4919);
or UO_209 (O_209,N_4911,N_4835);
or UO_210 (O_210,N_4830,N_4966);
and UO_211 (O_211,N_4957,N_4998);
xnor UO_212 (O_212,N_4887,N_4846);
xor UO_213 (O_213,N_4907,N_4891);
nand UO_214 (O_214,N_4841,N_4839);
nand UO_215 (O_215,N_4997,N_4839);
nand UO_216 (O_216,N_4840,N_4873);
nand UO_217 (O_217,N_4870,N_4950);
xnor UO_218 (O_218,N_4909,N_4809);
or UO_219 (O_219,N_4979,N_4977);
nand UO_220 (O_220,N_4888,N_4900);
nand UO_221 (O_221,N_4860,N_4896);
and UO_222 (O_222,N_4986,N_4956);
xor UO_223 (O_223,N_4847,N_4913);
or UO_224 (O_224,N_4991,N_4806);
nand UO_225 (O_225,N_4986,N_4871);
nor UO_226 (O_226,N_4923,N_4996);
and UO_227 (O_227,N_4887,N_4991);
nand UO_228 (O_228,N_4898,N_4858);
nor UO_229 (O_229,N_4864,N_4932);
nand UO_230 (O_230,N_4815,N_4953);
nand UO_231 (O_231,N_4907,N_4889);
and UO_232 (O_232,N_4923,N_4937);
and UO_233 (O_233,N_4985,N_4961);
nor UO_234 (O_234,N_4870,N_4916);
nor UO_235 (O_235,N_4878,N_4948);
xnor UO_236 (O_236,N_4825,N_4823);
and UO_237 (O_237,N_4815,N_4865);
and UO_238 (O_238,N_4914,N_4970);
or UO_239 (O_239,N_4881,N_4845);
or UO_240 (O_240,N_4812,N_4804);
nand UO_241 (O_241,N_4935,N_4882);
nand UO_242 (O_242,N_4977,N_4931);
xor UO_243 (O_243,N_4869,N_4908);
xnor UO_244 (O_244,N_4893,N_4933);
nor UO_245 (O_245,N_4880,N_4830);
xnor UO_246 (O_246,N_4930,N_4872);
nand UO_247 (O_247,N_4904,N_4894);
nand UO_248 (O_248,N_4957,N_4968);
and UO_249 (O_249,N_4998,N_4826);
and UO_250 (O_250,N_4895,N_4956);
and UO_251 (O_251,N_4861,N_4942);
and UO_252 (O_252,N_4897,N_4814);
nor UO_253 (O_253,N_4967,N_4990);
nand UO_254 (O_254,N_4800,N_4825);
nor UO_255 (O_255,N_4819,N_4858);
nor UO_256 (O_256,N_4974,N_4844);
nand UO_257 (O_257,N_4833,N_4912);
nand UO_258 (O_258,N_4900,N_4907);
nand UO_259 (O_259,N_4934,N_4852);
nor UO_260 (O_260,N_4990,N_4892);
xnor UO_261 (O_261,N_4877,N_4815);
nand UO_262 (O_262,N_4884,N_4836);
nand UO_263 (O_263,N_4870,N_4839);
nand UO_264 (O_264,N_4958,N_4939);
nand UO_265 (O_265,N_4889,N_4954);
and UO_266 (O_266,N_4944,N_4941);
and UO_267 (O_267,N_4855,N_4984);
or UO_268 (O_268,N_4970,N_4887);
or UO_269 (O_269,N_4860,N_4956);
or UO_270 (O_270,N_4809,N_4851);
or UO_271 (O_271,N_4978,N_4846);
xor UO_272 (O_272,N_4955,N_4960);
or UO_273 (O_273,N_4818,N_4987);
or UO_274 (O_274,N_4811,N_4814);
xor UO_275 (O_275,N_4954,N_4908);
nor UO_276 (O_276,N_4914,N_4843);
nor UO_277 (O_277,N_4850,N_4862);
and UO_278 (O_278,N_4859,N_4878);
xor UO_279 (O_279,N_4930,N_4832);
xnor UO_280 (O_280,N_4936,N_4963);
nor UO_281 (O_281,N_4807,N_4909);
nor UO_282 (O_282,N_4915,N_4870);
nor UO_283 (O_283,N_4976,N_4801);
or UO_284 (O_284,N_4827,N_4980);
or UO_285 (O_285,N_4812,N_4872);
or UO_286 (O_286,N_4993,N_4905);
nor UO_287 (O_287,N_4876,N_4833);
or UO_288 (O_288,N_4950,N_4910);
nand UO_289 (O_289,N_4969,N_4835);
nor UO_290 (O_290,N_4836,N_4837);
xor UO_291 (O_291,N_4959,N_4924);
xor UO_292 (O_292,N_4871,N_4846);
and UO_293 (O_293,N_4892,N_4874);
or UO_294 (O_294,N_4988,N_4863);
and UO_295 (O_295,N_4878,N_4958);
and UO_296 (O_296,N_4855,N_4944);
xnor UO_297 (O_297,N_4995,N_4936);
xor UO_298 (O_298,N_4844,N_4988);
and UO_299 (O_299,N_4811,N_4982);
nand UO_300 (O_300,N_4826,N_4925);
and UO_301 (O_301,N_4836,N_4905);
nor UO_302 (O_302,N_4892,N_4827);
or UO_303 (O_303,N_4873,N_4909);
or UO_304 (O_304,N_4851,N_4925);
xor UO_305 (O_305,N_4837,N_4922);
or UO_306 (O_306,N_4966,N_4975);
nand UO_307 (O_307,N_4861,N_4854);
nor UO_308 (O_308,N_4996,N_4969);
or UO_309 (O_309,N_4925,N_4850);
xnor UO_310 (O_310,N_4954,N_4876);
or UO_311 (O_311,N_4890,N_4901);
and UO_312 (O_312,N_4979,N_4834);
nor UO_313 (O_313,N_4933,N_4821);
or UO_314 (O_314,N_4827,N_4938);
nand UO_315 (O_315,N_4968,N_4970);
nand UO_316 (O_316,N_4954,N_4958);
nor UO_317 (O_317,N_4994,N_4850);
or UO_318 (O_318,N_4834,N_4945);
nand UO_319 (O_319,N_4825,N_4872);
and UO_320 (O_320,N_4888,N_4893);
xor UO_321 (O_321,N_4983,N_4896);
xor UO_322 (O_322,N_4803,N_4920);
nor UO_323 (O_323,N_4965,N_4864);
nand UO_324 (O_324,N_4830,N_4926);
or UO_325 (O_325,N_4915,N_4991);
nor UO_326 (O_326,N_4986,N_4841);
xnor UO_327 (O_327,N_4931,N_4936);
nand UO_328 (O_328,N_4921,N_4891);
and UO_329 (O_329,N_4989,N_4828);
nand UO_330 (O_330,N_4961,N_4900);
xnor UO_331 (O_331,N_4905,N_4948);
nor UO_332 (O_332,N_4869,N_4888);
or UO_333 (O_333,N_4859,N_4855);
xnor UO_334 (O_334,N_4904,N_4898);
nand UO_335 (O_335,N_4905,N_4935);
nand UO_336 (O_336,N_4981,N_4849);
nand UO_337 (O_337,N_4803,N_4882);
xor UO_338 (O_338,N_4902,N_4931);
nor UO_339 (O_339,N_4962,N_4957);
nor UO_340 (O_340,N_4902,N_4834);
or UO_341 (O_341,N_4925,N_4838);
nor UO_342 (O_342,N_4906,N_4908);
xor UO_343 (O_343,N_4874,N_4831);
xnor UO_344 (O_344,N_4822,N_4850);
or UO_345 (O_345,N_4979,N_4844);
and UO_346 (O_346,N_4948,N_4898);
nor UO_347 (O_347,N_4949,N_4853);
and UO_348 (O_348,N_4857,N_4800);
xor UO_349 (O_349,N_4873,N_4933);
or UO_350 (O_350,N_4989,N_4864);
xnor UO_351 (O_351,N_4995,N_4808);
and UO_352 (O_352,N_4908,N_4942);
nand UO_353 (O_353,N_4878,N_4966);
nor UO_354 (O_354,N_4876,N_4866);
and UO_355 (O_355,N_4858,N_4940);
xnor UO_356 (O_356,N_4987,N_4979);
xnor UO_357 (O_357,N_4944,N_4839);
nor UO_358 (O_358,N_4953,N_4891);
or UO_359 (O_359,N_4914,N_4995);
nand UO_360 (O_360,N_4842,N_4864);
nand UO_361 (O_361,N_4889,N_4888);
and UO_362 (O_362,N_4898,N_4819);
nand UO_363 (O_363,N_4896,N_4991);
nand UO_364 (O_364,N_4924,N_4934);
or UO_365 (O_365,N_4858,N_4855);
nor UO_366 (O_366,N_4882,N_4836);
or UO_367 (O_367,N_4884,N_4893);
xnor UO_368 (O_368,N_4912,N_4966);
or UO_369 (O_369,N_4946,N_4822);
nand UO_370 (O_370,N_4872,N_4937);
or UO_371 (O_371,N_4897,N_4958);
nand UO_372 (O_372,N_4855,N_4885);
or UO_373 (O_373,N_4826,N_4827);
nand UO_374 (O_374,N_4926,N_4866);
nand UO_375 (O_375,N_4882,N_4828);
xnor UO_376 (O_376,N_4985,N_4912);
nand UO_377 (O_377,N_4834,N_4899);
nand UO_378 (O_378,N_4951,N_4986);
nand UO_379 (O_379,N_4928,N_4827);
xnor UO_380 (O_380,N_4956,N_4818);
xnor UO_381 (O_381,N_4831,N_4863);
nand UO_382 (O_382,N_4860,N_4967);
nor UO_383 (O_383,N_4966,N_4803);
nand UO_384 (O_384,N_4931,N_4894);
nand UO_385 (O_385,N_4901,N_4983);
or UO_386 (O_386,N_4838,N_4843);
nor UO_387 (O_387,N_4962,N_4813);
nand UO_388 (O_388,N_4919,N_4973);
nor UO_389 (O_389,N_4930,N_4889);
nand UO_390 (O_390,N_4843,N_4919);
xnor UO_391 (O_391,N_4889,N_4860);
and UO_392 (O_392,N_4961,N_4869);
nor UO_393 (O_393,N_4814,N_4801);
nor UO_394 (O_394,N_4973,N_4901);
nand UO_395 (O_395,N_4993,N_4868);
and UO_396 (O_396,N_4975,N_4989);
nor UO_397 (O_397,N_4889,N_4938);
or UO_398 (O_398,N_4940,N_4819);
or UO_399 (O_399,N_4817,N_4833);
xnor UO_400 (O_400,N_4947,N_4831);
nor UO_401 (O_401,N_4845,N_4870);
nand UO_402 (O_402,N_4875,N_4988);
nor UO_403 (O_403,N_4989,N_4998);
nand UO_404 (O_404,N_4957,N_4928);
or UO_405 (O_405,N_4926,N_4939);
nor UO_406 (O_406,N_4814,N_4954);
nand UO_407 (O_407,N_4828,N_4856);
nand UO_408 (O_408,N_4965,N_4967);
nor UO_409 (O_409,N_4872,N_4807);
nor UO_410 (O_410,N_4863,N_4868);
nand UO_411 (O_411,N_4974,N_4984);
and UO_412 (O_412,N_4973,N_4830);
and UO_413 (O_413,N_4805,N_4947);
xnor UO_414 (O_414,N_4833,N_4815);
or UO_415 (O_415,N_4976,N_4998);
or UO_416 (O_416,N_4917,N_4871);
nand UO_417 (O_417,N_4910,N_4848);
nand UO_418 (O_418,N_4866,N_4920);
xnor UO_419 (O_419,N_4885,N_4859);
or UO_420 (O_420,N_4990,N_4841);
or UO_421 (O_421,N_4840,N_4844);
nand UO_422 (O_422,N_4805,N_4803);
nand UO_423 (O_423,N_4810,N_4863);
nor UO_424 (O_424,N_4943,N_4987);
nor UO_425 (O_425,N_4894,N_4992);
nor UO_426 (O_426,N_4973,N_4823);
xor UO_427 (O_427,N_4856,N_4873);
and UO_428 (O_428,N_4823,N_4945);
or UO_429 (O_429,N_4950,N_4975);
nand UO_430 (O_430,N_4914,N_4941);
and UO_431 (O_431,N_4922,N_4989);
nor UO_432 (O_432,N_4923,N_4968);
xor UO_433 (O_433,N_4895,N_4972);
nand UO_434 (O_434,N_4827,N_4847);
xnor UO_435 (O_435,N_4887,N_4840);
xnor UO_436 (O_436,N_4895,N_4934);
or UO_437 (O_437,N_4938,N_4998);
nand UO_438 (O_438,N_4811,N_4919);
nand UO_439 (O_439,N_4992,N_4811);
and UO_440 (O_440,N_4886,N_4873);
nor UO_441 (O_441,N_4822,N_4959);
nand UO_442 (O_442,N_4988,N_4803);
nor UO_443 (O_443,N_4886,N_4801);
xor UO_444 (O_444,N_4811,N_4875);
or UO_445 (O_445,N_4906,N_4806);
nor UO_446 (O_446,N_4868,N_4833);
nor UO_447 (O_447,N_4831,N_4948);
nor UO_448 (O_448,N_4860,N_4827);
nand UO_449 (O_449,N_4923,N_4846);
xnor UO_450 (O_450,N_4910,N_4868);
nand UO_451 (O_451,N_4843,N_4933);
and UO_452 (O_452,N_4928,N_4944);
and UO_453 (O_453,N_4921,N_4927);
nor UO_454 (O_454,N_4820,N_4857);
nor UO_455 (O_455,N_4953,N_4898);
and UO_456 (O_456,N_4974,N_4817);
nor UO_457 (O_457,N_4983,N_4916);
nand UO_458 (O_458,N_4845,N_4937);
and UO_459 (O_459,N_4912,N_4801);
or UO_460 (O_460,N_4856,N_4946);
nor UO_461 (O_461,N_4888,N_4879);
xor UO_462 (O_462,N_4969,N_4935);
and UO_463 (O_463,N_4832,N_4869);
or UO_464 (O_464,N_4894,N_4812);
or UO_465 (O_465,N_4931,N_4862);
nand UO_466 (O_466,N_4827,N_4903);
xor UO_467 (O_467,N_4946,N_4898);
nand UO_468 (O_468,N_4888,N_4887);
xnor UO_469 (O_469,N_4807,N_4819);
nand UO_470 (O_470,N_4960,N_4990);
nor UO_471 (O_471,N_4948,N_4994);
nand UO_472 (O_472,N_4824,N_4971);
nand UO_473 (O_473,N_4883,N_4915);
nand UO_474 (O_474,N_4870,N_4999);
and UO_475 (O_475,N_4816,N_4844);
nor UO_476 (O_476,N_4806,N_4885);
xor UO_477 (O_477,N_4840,N_4934);
and UO_478 (O_478,N_4828,N_4830);
and UO_479 (O_479,N_4952,N_4967);
nor UO_480 (O_480,N_4981,N_4858);
or UO_481 (O_481,N_4893,N_4906);
nand UO_482 (O_482,N_4986,N_4820);
xnor UO_483 (O_483,N_4948,N_4918);
nor UO_484 (O_484,N_4875,N_4838);
or UO_485 (O_485,N_4969,N_4916);
nand UO_486 (O_486,N_4915,N_4849);
xnor UO_487 (O_487,N_4856,N_4880);
or UO_488 (O_488,N_4955,N_4973);
nand UO_489 (O_489,N_4940,N_4954);
and UO_490 (O_490,N_4863,N_4879);
nand UO_491 (O_491,N_4994,N_4844);
xnor UO_492 (O_492,N_4832,N_4835);
nand UO_493 (O_493,N_4995,N_4849);
nand UO_494 (O_494,N_4981,N_4870);
or UO_495 (O_495,N_4807,N_4893);
nand UO_496 (O_496,N_4889,N_4895);
xnor UO_497 (O_497,N_4918,N_4854);
nor UO_498 (O_498,N_4841,N_4939);
and UO_499 (O_499,N_4817,N_4979);
nor UO_500 (O_500,N_4860,N_4809);
or UO_501 (O_501,N_4828,N_4814);
and UO_502 (O_502,N_4852,N_4858);
or UO_503 (O_503,N_4967,N_4974);
xor UO_504 (O_504,N_4991,N_4889);
and UO_505 (O_505,N_4964,N_4826);
nor UO_506 (O_506,N_4807,N_4885);
nor UO_507 (O_507,N_4887,N_4881);
xor UO_508 (O_508,N_4892,N_4864);
nor UO_509 (O_509,N_4973,N_4962);
or UO_510 (O_510,N_4883,N_4922);
nor UO_511 (O_511,N_4892,N_4845);
nand UO_512 (O_512,N_4827,N_4874);
xnor UO_513 (O_513,N_4972,N_4918);
nand UO_514 (O_514,N_4944,N_4924);
nand UO_515 (O_515,N_4812,N_4956);
xnor UO_516 (O_516,N_4899,N_4967);
nor UO_517 (O_517,N_4872,N_4830);
nor UO_518 (O_518,N_4935,N_4804);
xnor UO_519 (O_519,N_4925,N_4922);
nand UO_520 (O_520,N_4983,N_4877);
and UO_521 (O_521,N_4865,N_4971);
or UO_522 (O_522,N_4918,N_4907);
xor UO_523 (O_523,N_4935,N_4826);
or UO_524 (O_524,N_4816,N_4953);
and UO_525 (O_525,N_4826,N_4874);
nand UO_526 (O_526,N_4831,N_4910);
nor UO_527 (O_527,N_4969,N_4948);
and UO_528 (O_528,N_4925,N_4869);
and UO_529 (O_529,N_4813,N_4834);
nor UO_530 (O_530,N_4970,N_4918);
or UO_531 (O_531,N_4852,N_4807);
or UO_532 (O_532,N_4849,N_4894);
or UO_533 (O_533,N_4876,N_4839);
nand UO_534 (O_534,N_4832,N_4926);
and UO_535 (O_535,N_4813,N_4850);
and UO_536 (O_536,N_4982,N_4890);
nor UO_537 (O_537,N_4944,N_4942);
or UO_538 (O_538,N_4985,N_4909);
nand UO_539 (O_539,N_4912,N_4820);
xnor UO_540 (O_540,N_4814,N_4860);
and UO_541 (O_541,N_4929,N_4817);
xor UO_542 (O_542,N_4921,N_4928);
nor UO_543 (O_543,N_4954,N_4950);
or UO_544 (O_544,N_4852,N_4949);
nand UO_545 (O_545,N_4970,N_4945);
nor UO_546 (O_546,N_4811,N_4954);
nor UO_547 (O_547,N_4919,N_4874);
xnor UO_548 (O_548,N_4854,N_4868);
nor UO_549 (O_549,N_4880,N_4873);
nand UO_550 (O_550,N_4919,N_4810);
or UO_551 (O_551,N_4980,N_4821);
nand UO_552 (O_552,N_4874,N_4904);
xor UO_553 (O_553,N_4924,N_4835);
or UO_554 (O_554,N_4822,N_4902);
nor UO_555 (O_555,N_4976,N_4957);
nand UO_556 (O_556,N_4882,N_4907);
nor UO_557 (O_557,N_4818,N_4953);
nor UO_558 (O_558,N_4923,N_4848);
or UO_559 (O_559,N_4906,N_4941);
and UO_560 (O_560,N_4816,N_4916);
nor UO_561 (O_561,N_4920,N_4836);
nand UO_562 (O_562,N_4897,N_4888);
or UO_563 (O_563,N_4803,N_4952);
or UO_564 (O_564,N_4931,N_4850);
or UO_565 (O_565,N_4945,N_4832);
xnor UO_566 (O_566,N_4906,N_4930);
xnor UO_567 (O_567,N_4940,N_4841);
nor UO_568 (O_568,N_4899,N_4825);
or UO_569 (O_569,N_4980,N_4930);
or UO_570 (O_570,N_4900,N_4993);
and UO_571 (O_571,N_4825,N_4971);
xor UO_572 (O_572,N_4964,N_4974);
or UO_573 (O_573,N_4985,N_4922);
nor UO_574 (O_574,N_4850,N_4910);
nand UO_575 (O_575,N_4899,N_4801);
and UO_576 (O_576,N_4922,N_4867);
or UO_577 (O_577,N_4824,N_4897);
nor UO_578 (O_578,N_4968,N_4802);
xnor UO_579 (O_579,N_4824,N_4854);
and UO_580 (O_580,N_4878,N_4921);
or UO_581 (O_581,N_4802,N_4990);
xnor UO_582 (O_582,N_4910,N_4865);
nor UO_583 (O_583,N_4916,N_4885);
nor UO_584 (O_584,N_4927,N_4974);
nor UO_585 (O_585,N_4928,N_4949);
and UO_586 (O_586,N_4935,N_4981);
and UO_587 (O_587,N_4800,N_4879);
nand UO_588 (O_588,N_4838,N_4954);
nand UO_589 (O_589,N_4952,N_4853);
or UO_590 (O_590,N_4884,N_4979);
xnor UO_591 (O_591,N_4834,N_4889);
nor UO_592 (O_592,N_4885,N_4945);
xor UO_593 (O_593,N_4891,N_4956);
nor UO_594 (O_594,N_4888,N_4875);
xor UO_595 (O_595,N_4840,N_4963);
nor UO_596 (O_596,N_4834,N_4839);
and UO_597 (O_597,N_4888,N_4967);
nor UO_598 (O_598,N_4858,N_4865);
nand UO_599 (O_599,N_4978,N_4905);
and UO_600 (O_600,N_4900,N_4926);
and UO_601 (O_601,N_4836,N_4901);
xnor UO_602 (O_602,N_4895,N_4940);
xor UO_603 (O_603,N_4823,N_4904);
nand UO_604 (O_604,N_4933,N_4850);
nor UO_605 (O_605,N_4800,N_4922);
or UO_606 (O_606,N_4815,N_4928);
and UO_607 (O_607,N_4972,N_4887);
and UO_608 (O_608,N_4962,N_4863);
and UO_609 (O_609,N_4941,N_4807);
or UO_610 (O_610,N_4995,N_4870);
xnor UO_611 (O_611,N_4829,N_4995);
nand UO_612 (O_612,N_4857,N_4969);
or UO_613 (O_613,N_4993,N_4949);
or UO_614 (O_614,N_4845,N_4890);
nand UO_615 (O_615,N_4822,N_4849);
nor UO_616 (O_616,N_4926,N_4904);
nand UO_617 (O_617,N_4969,N_4923);
nand UO_618 (O_618,N_4936,N_4895);
or UO_619 (O_619,N_4940,N_4991);
nand UO_620 (O_620,N_4934,N_4955);
nand UO_621 (O_621,N_4938,N_4806);
nor UO_622 (O_622,N_4958,N_4809);
and UO_623 (O_623,N_4911,N_4984);
and UO_624 (O_624,N_4945,N_4862);
or UO_625 (O_625,N_4986,N_4962);
or UO_626 (O_626,N_4911,N_4969);
or UO_627 (O_627,N_4856,N_4838);
nor UO_628 (O_628,N_4933,N_4876);
and UO_629 (O_629,N_4912,N_4832);
nor UO_630 (O_630,N_4804,N_4959);
nand UO_631 (O_631,N_4963,N_4931);
nand UO_632 (O_632,N_4850,N_4811);
or UO_633 (O_633,N_4912,N_4887);
xor UO_634 (O_634,N_4924,N_4931);
nor UO_635 (O_635,N_4946,N_4887);
or UO_636 (O_636,N_4817,N_4922);
nand UO_637 (O_637,N_4926,N_4822);
nor UO_638 (O_638,N_4843,N_4868);
nor UO_639 (O_639,N_4851,N_4990);
and UO_640 (O_640,N_4875,N_4851);
nand UO_641 (O_641,N_4870,N_4834);
nand UO_642 (O_642,N_4996,N_4938);
xnor UO_643 (O_643,N_4818,N_4864);
xnor UO_644 (O_644,N_4947,N_4907);
and UO_645 (O_645,N_4824,N_4834);
nor UO_646 (O_646,N_4953,N_4923);
nand UO_647 (O_647,N_4841,N_4943);
xnor UO_648 (O_648,N_4837,N_4809);
nor UO_649 (O_649,N_4932,N_4903);
nand UO_650 (O_650,N_4971,N_4982);
xor UO_651 (O_651,N_4937,N_4807);
nand UO_652 (O_652,N_4996,N_4805);
and UO_653 (O_653,N_4840,N_4808);
nand UO_654 (O_654,N_4946,N_4982);
nor UO_655 (O_655,N_4941,N_4836);
nand UO_656 (O_656,N_4864,N_4819);
xor UO_657 (O_657,N_4955,N_4943);
nand UO_658 (O_658,N_4885,N_4951);
nand UO_659 (O_659,N_4898,N_4848);
xnor UO_660 (O_660,N_4849,N_4815);
nor UO_661 (O_661,N_4890,N_4957);
nand UO_662 (O_662,N_4964,N_4801);
xor UO_663 (O_663,N_4873,N_4989);
nand UO_664 (O_664,N_4990,N_4939);
and UO_665 (O_665,N_4894,N_4869);
or UO_666 (O_666,N_4867,N_4815);
xnor UO_667 (O_667,N_4848,N_4913);
xnor UO_668 (O_668,N_4819,N_4818);
and UO_669 (O_669,N_4964,N_4948);
nor UO_670 (O_670,N_4893,N_4910);
nand UO_671 (O_671,N_4992,N_4907);
nand UO_672 (O_672,N_4975,N_4945);
nand UO_673 (O_673,N_4889,N_4822);
nand UO_674 (O_674,N_4808,N_4851);
nand UO_675 (O_675,N_4955,N_4967);
and UO_676 (O_676,N_4925,N_4919);
nand UO_677 (O_677,N_4883,N_4846);
xnor UO_678 (O_678,N_4857,N_4901);
xnor UO_679 (O_679,N_4854,N_4908);
nand UO_680 (O_680,N_4868,N_4893);
xor UO_681 (O_681,N_4935,N_4908);
and UO_682 (O_682,N_4984,N_4940);
or UO_683 (O_683,N_4890,N_4947);
and UO_684 (O_684,N_4812,N_4921);
and UO_685 (O_685,N_4861,N_4994);
nor UO_686 (O_686,N_4936,N_4880);
nand UO_687 (O_687,N_4850,N_4912);
nor UO_688 (O_688,N_4805,N_4992);
nand UO_689 (O_689,N_4972,N_4890);
nand UO_690 (O_690,N_4914,N_4819);
nand UO_691 (O_691,N_4807,N_4959);
and UO_692 (O_692,N_4930,N_4855);
or UO_693 (O_693,N_4866,N_4904);
nor UO_694 (O_694,N_4919,N_4932);
xor UO_695 (O_695,N_4893,N_4826);
nand UO_696 (O_696,N_4989,N_4870);
or UO_697 (O_697,N_4886,N_4895);
xor UO_698 (O_698,N_4905,N_4825);
or UO_699 (O_699,N_4988,N_4824);
and UO_700 (O_700,N_4800,N_4980);
xnor UO_701 (O_701,N_4875,N_4889);
xor UO_702 (O_702,N_4966,N_4897);
or UO_703 (O_703,N_4992,N_4829);
nand UO_704 (O_704,N_4955,N_4916);
nand UO_705 (O_705,N_4893,N_4955);
nand UO_706 (O_706,N_4919,N_4807);
xnor UO_707 (O_707,N_4893,N_4921);
nor UO_708 (O_708,N_4969,N_4945);
or UO_709 (O_709,N_4845,N_4843);
nand UO_710 (O_710,N_4900,N_4837);
or UO_711 (O_711,N_4878,N_4820);
or UO_712 (O_712,N_4958,N_4947);
xnor UO_713 (O_713,N_4965,N_4951);
and UO_714 (O_714,N_4904,N_4895);
or UO_715 (O_715,N_4899,N_4923);
nor UO_716 (O_716,N_4854,N_4874);
nor UO_717 (O_717,N_4835,N_4802);
nor UO_718 (O_718,N_4963,N_4802);
and UO_719 (O_719,N_4987,N_4881);
and UO_720 (O_720,N_4859,N_4970);
xor UO_721 (O_721,N_4963,N_4863);
nand UO_722 (O_722,N_4970,N_4879);
nor UO_723 (O_723,N_4955,N_4956);
and UO_724 (O_724,N_4878,N_4801);
or UO_725 (O_725,N_4828,N_4861);
nand UO_726 (O_726,N_4909,N_4802);
and UO_727 (O_727,N_4808,N_4807);
xor UO_728 (O_728,N_4809,N_4802);
or UO_729 (O_729,N_4865,N_4831);
xnor UO_730 (O_730,N_4824,N_4996);
and UO_731 (O_731,N_4880,N_4990);
nor UO_732 (O_732,N_4988,N_4869);
nand UO_733 (O_733,N_4938,N_4909);
nand UO_734 (O_734,N_4852,N_4834);
nand UO_735 (O_735,N_4965,N_4986);
nor UO_736 (O_736,N_4870,N_4830);
xnor UO_737 (O_737,N_4973,N_4984);
and UO_738 (O_738,N_4832,N_4811);
and UO_739 (O_739,N_4859,N_4960);
nand UO_740 (O_740,N_4972,N_4901);
nand UO_741 (O_741,N_4992,N_4957);
xor UO_742 (O_742,N_4993,N_4930);
nand UO_743 (O_743,N_4975,N_4916);
xor UO_744 (O_744,N_4889,N_4981);
nand UO_745 (O_745,N_4836,N_4971);
xor UO_746 (O_746,N_4947,N_4914);
nor UO_747 (O_747,N_4945,N_4986);
or UO_748 (O_748,N_4864,N_4858);
nand UO_749 (O_749,N_4859,N_4841);
nand UO_750 (O_750,N_4914,N_4961);
nand UO_751 (O_751,N_4824,N_4872);
xnor UO_752 (O_752,N_4801,N_4984);
nor UO_753 (O_753,N_4966,N_4943);
nand UO_754 (O_754,N_4895,N_4941);
and UO_755 (O_755,N_4833,N_4820);
and UO_756 (O_756,N_4914,N_4960);
nor UO_757 (O_757,N_4988,N_4877);
or UO_758 (O_758,N_4816,N_4845);
and UO_759 (O_759,N_4931,N_4835);
nand UO_760 (O_760,N_4834,N_4919);
nor UO_761 (O_761,N_4874,N_4915);
or UO_762 (O_762,N_4852,N_4862);
xnor UO_763 (O_763,N_4983,N_4850);
nand UO_764 (O_764,N_4947,N_4853);
nand UO_765 (O_765,N_4967,N_4921);
and UO_766 (O_766,N_4809,N_4881);
and UO_767 (O_767,N_4827,N_4941);
and UO_768 (O_768,N_4872,N_4948);
nor UO_769 (O_769,N_4817,N_4868);
nand UO_770 (O_770,N_4905,N_4866);
or UO_771 (O_771,N_4905,N_4850);
or UO_772 (O_772,N_4805,N_4980);
and UO_773 (O_773,N_4862,N_4849);
nand UO_774 (O_774,N_4845,N_4848);
or UO_775 (O_775,N_4889,N_4900);
and UO_776 (O_776,N_4914,N_4998);
and UO_777 (O_777,N_4869,N_4957);
xor UO_778 (O_778,N_4987,N_4854);
nor UO_779 (O_779,N_4977,N_4853);
xnor UO_780 (O_780,N_4843,N_4927);
nor UO_781 (O_781,N_4945,N_4825);
and UO_782 (O_782,N_4822,N_4998);
nor UO_783 (O_783,N_4864,N_4824);
or UO_784 (O_784,N_4937,N_4927);
or UO_785 (O_785,N_4854,N_4973);
or UO_786 (O_786,N_4868,N_4869);
xnor UO_787 (O_787,N_4943,N_4830);
xnor UO_788 (O_788,N_4926,N_4855);
nor UO_789 (O_789,N_4965,N_4985);
xnor UO_790 (O_790,N_4988,N_4849);
nor UO_791 (O_791,N_4936,N_4886);
xnor UO_792 (O_792,N_4888,N_4886);
or UO_793 (O_793,N_4984,N_4918);
nand UO_794 (O_794,N_4810,N_4959);
or UO_795 (O_795,N_4806,N_4816);
or UO_796 (O_796,N_4879,N_4973);
or UO_797 (O_797,N_4917,N_4981);
nor UO_798 (O_798,N_4951,N_4838);
nand UO_799 (O_799,N_4983,N_4882);
nor UO_800 (O_800,N_4992,N_4825);
xnor UO_801 (O_801,N_4828,N_4848);
xor UO_802 (O_802,N_4965,N_4879);
xnor UO_803 (O_803,N_4899,N_4816);
nand UO_804 (O_804,N_4955,N_4968);
xnor UO_805 (O_805,N_4963,N_4875);
nor UO_806 (O_806,N_4883,N_4902);
and UO_807 (O_807,N_4907,N_4850);
nor UO_808 (O_808,N_4954,N_4951);
xnor UO_809 (O_809,N_4951,N_4952);
nand UO_810 (O_810,N_4893,N_4860);
xor UO_811 (O_811,N_4987,N_4814);
nand UO_812 (O_812,N_4963,N_4834);
xor UO_813 (O_813,N_4812,N_4985);
or UO_814 (O_814,N_4869,N_4962);
and UO_815 (O_815,N_4801,N_4956);
nand UO_816 (O_816,N_4820,N_4930);
nor UO_817 (O_817,N_4969,N_4934);
or UO_818 (O_818,N_4945,N_4884);
xor UO_819 (O_819,N_4988,N_4936);
and UO_820 (O_820,N_4972,N_4806);
nand UO_821 (O_821,N_4837,N_4870);
or UO_822 (O_822,N_4959,N_4980);
nor UO_823 (O_823,N_4892,N_4989);
and UO_824 (O_824,N_4972,N_4897);
and UO_825 (O_825,N_4838,N_4921);
xor UO_826 (O_826,N_4911,N_4868);
nor UO_827 (O_827,N_4997,N_4862);
and UO_828 (O_828,N_4834,N_4805);
nand UO_829 (O_829,N_4935,N_4886);
xor UO_830 (O_830,N_4938,N_4937);
nand UO_831 (O_831,N_4999,N_4944);
or UO_832 (O_832,N_4976,N_4920);
nand UO_833 (O_833,N_4958,N_4826);
nor UO_834 (O_834,N_4956,N_4850);
or UO_835 (O_835,N_4879,N_4841);
or UO_836 (O_836,N_4837,N_4964);
or UO_837 (O_837,N_4860,N_4895);
or UO_838 (O_838,N_4993,N_4808);
and UO_839 (O_839,N_4990,N_4966);
xnor UO_840 (O_840,N_4837,N_4910);
xor UO_841 (O_841,N_4905,N_4992);
nor UO_842 (O_842,N_4856,N_4869);
xor UO_843 (O_843,N_4863,N_4905);
xnor UO_844 (O_844,N_4814,N_4842);
or UO_845 (O_845,N_4882,N_4888);
xor UO_846 (O_846,N_4915,N_4966);
xor UO_847 (O_847,N_4895,N_4933);
or UO_848 (O_848,N_4876,N_4803);
or UO_849 (O_849,N_4943,N_4838);
xnor UO_850 (O_850,N_4929,N_4978);
nor UO_851 (O_851,N_4862,N_4958);
and UO_852 (O_852,N_4826,N_4962);
and UO_853 (O_853,N_4810,N_4829);
or UO_854 (O_854,N_4977,N_4916);
or UO_855 (O_855,N_4927,N_4874);
or UO_856 (O_856,N_4846,N_4853);
and UO_857 (O_857,N_4818,N_4830);
and UO_858 (O_858,N_4889,N_4814);
nor UO_859 (O_859,N_4876,N_4843);
or UO_860 (O_860,N_4881,N_4936);
or UO_861 (O_861,N_4855,N_4950);
and UO_862 (O_862,N_4834,N_4843);
nand UO_863 (O_863,N_4879,N_4821);
and UO_864 (O_864,N_4869,N_4874);
or UO_865 (O_865,N_4952,N_4998);
nand UO_866 (O_866,N_4978,N_4898);
or UO_867 (O_867,N_4939,N_4949);
and UO_868 (O_868,N_4986,N_4952);
or UO_869 (O_869,N_4872,N_4953);
and UO_870 (O_870,N_4857,N_4822);
nor UO_871 (O_871,N_4834,N_4955);
xor UO_872 (O_872,N_4934,N_4842);
or UO_873 (O_873,N_4845,N_4980);
and UO_874 (O_874,N_4953,N_4878);
or UO_875 (O_875,N_4977,N_4968);
nand UO_876 (O_876,N_4981,N_4959);
nor UO_877 (O_877,N_4973,N_4898);
nor UO_878 (O_878,N_4850,N_4854);
xor UO_879 (O_879,N_4872,N_4884);
xnor UO_880 (O_880,N_4961,N_4941);
nand UO_881 (O_881,N_4940,N_4930);
nor UO_882 (O_882,N_4821,N_4934);
nand UO_883 (O_883,N_4817,N_4965);
nand UO_884 (O_884,N_4851,N_4955);
xor UO_885 (O_885,N_4913,N_4824);
and UO_886 (O_886,N_4900,N_4821);
nor UO_887 (O_887,N_4823,N_4866);
and UO_888 (O_888,N_4882,N_4802);
or UO_889 (O_889,N_4870,N_4923);
or UO_890 (O_890,N_4983,N_4957);
and UO_891 (O_891,N_4905,N_4995);
nand UO_892 (O_892,N_4838,N_4859);
xnor UO_893 (O_893,N_4893,N_4827);
and UO_894 (O_894,N_4988,N_4881);
or UO_895 (O_895,N_4908,N_4800);
nand UO_896 (O_896,N_4903,N_4937);
nand UO_897 (O_897,N_4822,N_4813);
nand UO_898 (O_898,N_4943,N_4808);
xnor UO_899 (O_899,N_4881,N_4934);
nand UO_900 (O_900,N_4839,N_4984);
and UO_901 (O_901,N_4890,N_4927);
nor UO_902 (O_902,N_4960,N_4856);
nor UO_903 (O_903,N_4816,N_4975);
and UO_904 (O_904,N_4863,N_4816);
nor UO_905 (O_905,N_4917,N_4966);
and UO_906 (O_906,N_4836,N_4987);
and UO_907 (O_907,N_4814,N_4957);
and UO_908 (O_908,N_4927,N_4873);
and UO_909 (O_909,N_4916,N_4900);
or UO_910 (O_910,N_4943,N_4894);
or UO_911 (O_911,N_4897,N_4908);
xor UO_912 (O_912,N_4891,N_4955);
xnor UO_913 (O_913,N_4975,N_4895);
and UO_914 (O_914,N_4968,N_4824);
and UO_915 (O_915,N_4942,N_4901);
xor UO_916 (O_916,N_4927,N_4980);
or UO_917 (O_917,N_4832,N_4981);
nand UO_918 (O_918,N_4878,N_4854);
nand UO_919 (O_919,N_4857,N_4861);
and UO_920 (O_920,N_4954,N_4820);
and UO_921 (O_921,N_4985,N_4926);
and UO_922 (O_922,N_4884,N_4821);
xor UO_923 (O_923,N_4840,N_4952);
and UO_924 (O_924,N_4899,N_4941);
and UO_925 (O_925,N_4950,N_4820);
nor UO_926 (O_926,N_4990,N_4807);
nand UO_927 (O_927,N_4874,N_4825);
nand UO_928 (O_928,N_4934,N_4948);
nand UO_929 (O_929,N_4951,N_4835);
nor UO_930 (O_930,N_4869,N_4972);
or UO_931 (O_931,N_4883,N_4937);
nor UO_932 (O_932,N_4946,N_4842);
nor UO_933 (O_933,N_4806,N_4916);
nor UO_934 (O_934,N_4857,N_4841);
nand UO_935 (O_935,N_4854,N_4927);
nand UO_936 (O_936,N_4862,N_4888);
xnor UO_937 (O_937,N_4873,N_4938);
or UO_938 (O_938,N_4922,N_4993);
or UO_939 (O_939,N_4873,N_4891);
or UO_940 (O_940,N_4918,N_4814);
or UO_941 (O_941,N_4859,N_4903);
or UO_942 (O_942,N_4946,N_4872);
or UO_943 (O_943,N_4951,N_4918);
xnor UO_944 (O_944,N_4802,N_4806);
nor UO_945 (O_945,N_4813,N_4837);
nand UO_946 (O_946,N_4931,N_4809);
xor UO_947 (O_947,N_4976,N_4973);
nand UO_948 (O_948,N_4934,N_4827);
and UO_949 (O_949,N_4871,N_4937);
and UO_950 (O_950,N_4891,N_4844);
and UO_951 (O_951,N_4931,N_4824);
nor UO_952 (O_952,N_4982,N_4923);
or UO_953 (O_953,N_4872,N_4840);
nor UO_954 (O_954,N_4900,N_4938);
or UO_955 (O_955,N_4829,N_4827);
and UO_956 (O_956,N_4810,N_4908);
or UO_957 (O_957,N_4962,N_4945);
or UO_958 (O_958,N_4911,N_4816);
nand UO_959 (O_959,N_4904,N_4961);
or UO_960 (O_960,N_4805,N_4838);
xnor UO_961 (O_961,N_4813,N_4990);
or UO_962 (O_962,N_4917,N_4838);
or UO_963 (O_963,N_4930,N_4884);
nor UO_964 (O_964,N_4906,N_4839);
nand UO_965 (O_965,N_4855,N_4821);
or UO_966 (O_966,N_4889,N_4964);
or UO_967 (O_967,N_4993,N_4971);
nor UO_968 (O_968,N_4801,N_4887);
nor UO_969 (O_969,N_4968,N_4893);
nor UO_970 (O_970,N_4993,N_4939);
xor UO_971 (O_971,N_4872,N_4837);
xor UO_972 (O_972,N_4846,N_4986);
nor UO_973 (O_973,N_4986,N_4891);
and UO_974 (O_974,N_4939,N_4999);
nand UO_975 (O_975,N_4923,N_4926);
nor UO_976 (O_976,N_4935,N_4842);
and UO_977 (O_977,N_4895,N_4865);
xor UO_978 (O_978,N_4905,N_4889);
or UO_979 (O_979,N_4920,N_4996);
nor UO_980 (O_980,N_4948,N_4876);
or UO_981 (O_981,N_4975,N_4866);
xor UO_982 (O_982,N_4957,N_4913);
and UO_983 (O_983,N_4986,N_4813);
and UO_984 (O_984,N_4850,N_4903);
nor UO_985 (O_985,N_4897,N_4949);
or UO_986 (O_986,N_4828,N_4916);
xor UO_987 (O_987,N_4995,N_4908);
xnor UO_988 (O_988,N_4924,N_4851);
and UO_989 (O_989,N_4855,N_4904);
nand UO_990 (O_990,N_4828,N_4843);
nor UO_991 (O_991,N_4844,N_4982);
nor UO_992 (O_992,N_4822,N_4922);
xnor UO_993 (O_993,N_4966,N_4827);
nand UO_994 (O_994,N_4957,N_4805);
and UO_995 (O_995,N_4949,N_4869);
xnor UO_996 (O_996,N_4942,N_4962);
nand UO_997 (O_997,N_4913,N_4833);
nor UO_998 (O_998,N_4876,N_4951);
xor UO_999 (O_999,N_4827,N_4843);
endmodule