module basic_500_3000_500_60_levels_2xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_296,In_286);
nor U1 (N_1,In_191,In_7);
and U2 (N_2,In_164,In_358);
nor U3 (N_3,In_400,In_74);
or U4 (N_4,In_349,In_421);
and U5 (N_5,In_390,In_226);
nor U6 (N_6,In_347,In_50);
nor U7 (N_7,In_489,In_172);
and U8 (N_8,In_289,In_426);
nor U9 (N_9,In_395,In_352);
or U10 (N_10,In_449,In_469);
nor U11 (N_11,In_423,In_133);
nor U12 (N_12,In_419,In_236);
or U13 (N_13,In_47,In_63);
nand U14 (N_14,In_486,In_44);
or U15 (N_15,In_269,In_313);
nand U16 (N_16,In_430,In_276);
nand U17 (N_17,In_16,In_314);
nor U18 (N_18,In_285,In_483);
or U19 (N_19,In_246,In_362);
and U20 (N_20,In_279,In_363);
or U21 (N_21,In_413,In_273);
nor U22 (N_22,In_447,In_141);
nor U23 (N_23,In_379,In_482);
nor U24 (N_24,In_192,In_374);
or U25 (N_25,In_368,In_4);
nand U26 (N_26,In_18,In_163);
nand U27 (N_27,In_101,In_54);
and U28 (N_28,In_418,In_306);
or U29 (N_29,In_341,In_458);
nand U30 (N_30,In_278,In_144);
nand U31 (N_31,In_274,In_28);
and U32 (N_32,In_224,In_179);
nor U33 (N_33,In_340,In_478);
nand U34 (N_34,In_221,In_20);
or U35 (N_35,In_206,In_99);
nand U36 (N_36,In_290,In_348);
nor U37 (N_37,In_175,In_403);
and U38 (N_38,In_176,In_309);
nor U39 (N_39,In_51,In_448);
nor U40 (N_40,In_250,In_337);
or U41 (N_41,In_304,In_117);
or U42 (N_42,In_152,In_215);
nand U43 (N_43,In_312,In_109);
nor U44 (N_44,In_477,In_254);
and U45 (N_45,In_231,In_267);
nand U46 (N_46,In_9,In_135);
nand U47 (N_47,In_451,In_414);
nor U48 (N_48,In_234,In_339);
nor U49 (N_49,In_405,In_329);
or U50 (N_50,In_190,In_387);
nor U51 (N_51,In_444,In_456);
xor U52 (N_52,In_38,In_394);
and U53 (N_53,In_480,In_169);
nand U54 (N_54,In_216,N_0);
nor U55 (N_55,In_31,In_167);
nand U56 (N_56,In_159,In_33);
nor U57 (N_57,In_199,In_377);
nand U58 (N_58,In_454,In_407);
nor U59 (N_59,In_61,In_62);
and U60 (N_60,In_131,In_177);
or U61 (N_61,In_212,In_227);
and U62 (N_62,In_432,In_265);
and U63 (N_63,In_208,In_459);
or U64 (N_64,In_137,In_282);
nand U65 (N_65,In_154,In_55);
or U66 (N_66,In_409,In_326);
nand U67 (N_67,In_126,In_41);
and U68 (N_68,In_168,In_283);
or U69 (N_69,In_263,N_15);
and U70 (N_70,In_485,N_4);
nor U71 (N_71,In_183,In_331);
nor U72 (N_72,In_196,In_261);
and U73 (N_73,In_219,In_357);
nor U74 (N_74,In_19,N_21);
xor U75 (N_75,In_58,In_123);
nor U76 (N_76,In_284,In_66);
nand U77 (N_77,In_27,In_270);
nand U78 (N_78,In_130,In_12);
and U79 (N_79,In_193,In_499);
or U80 (N_80,In_411,In_264);
nand U81 (N_81,In_355,In_60);
and U82 (N_82,In_287,N_5);
and U83 (N_83,In_0,In_452);
nand U84 (N_84,In_369,In_136);
or U85 (N_85,In_497,In_84);
nor U86 (N_86,In_392,In_437);
nor U87 (N_87,In_461,In_67);
xnor U88 (N_88,In_83,In_210);
nor U89 (N_89,In_460,In_440);
or U90 (N_90,In_380,In_52);
nor U91 (N_91,In_376,In_338);
or U92 (N_92,In_149,In_57);
xnor U93 (N_93,In_217,In_324);
or U94 (N_94,In_23,In_156);
nand U95 (N_95,N_24,In_92);
nor U96 (N_96,In_252,In_373);
or U97 (N_97,In_463,In_297);
and U98 (N_98,In_105,In_147);
or U99 (N_99,In_481,In_434);
and U100 (N_100,In_402,In_132);
nand U101 (N_101,In_360,In_361);
nor U102 (N_102,In_239,In_351);
and U103 (N_103,N_18,In_86);
and U104 (N_104,In_404,In_325);
and U105 (N_105,In_140,In_96);
or U106 (N_106,In_195,N_86);
nor U107 (N_107,In_40,In_128);
and U108 (N_108,In_198,In_32);
nand U109 (N_109,In_476,In_435);
or U110 (N_110,In_81,In_238);
or U111 (N_111,In_155,In_300);
nor U112 (N_112,In_13,In_39);
or U113 (N_113,In_307,In_294);
nor U114 (N_114,In_272,In_124);
xnor U115 (N_115,In_364,In_315);
nor U116 (N_116,In_120,N_3);
or U117 (N_117,In_366,In_11);
nor U118 (N_118,In_108,In_420);
and U119 (N_119,In_77,N_6);
nor U120 (N_120,In_470,N_77);
xnor U121 (N_121,In_194,In_88);
or U122 (N_122,In_327,In_429);
and U123 (N_123,N_91,In_310);
nand U124 (N_124,N_31,In_153);
or U125 (N_125,In_111,In_253);
nand U126 (N_126,N_52,In_122);
or U127 (N_127,In_229,N_96);
nand U128 (N_128,N_20,N_60);
nor U129 (N_129,N_67,In_268);
nand U130 (N_130,In_431,In_75);
nand U131 (N_131,In_71,In_383);
nor U132 (N_132,In_473,N_69);
and U133 (N_133,In_334,In_491);
nor U134 (N_134,In_112,In_100);
or U135 (N_135,In_415,In_30);
nand U136 (N_136,In_378,In_359);
nor U137 (N_137,In_174,In_249);
and U138 (N_138,In_43,In_1);
and U139 (N_139,In_445,N_89);
nor U140 (N_140,In_76,N_29);
nor U141 (N_141,In_433,N_37);
nor U142 (N_142,In_46,In_271);
nor U143 (N_143,In_259,In_382);
nor U144 (N_144,In_145,In_406);
or U145 (N_145,In_25,In_479);
and U146 (N_146,N_66,In_391);
and U147 (N_147,N_34,N_85);
or U148 (N_148,In_298,In_370);
nor U149 (N_149,In_350,In_484);
nand U150 (N_150,N_90,In_53);
or U151 (N_151,In_464,In_35);
nor U152 (N_152,In_427,In_34);
or U153 (N_153,In_346,In_488);
nor U154 (N_154,In_15,N_8);
nand U155 (N_155,N_125,N_87);
or U156 (N_156,N_83,N_43);
nor U157 (N_157,In_213,N_142);
and U158 (N_158,N_147,In_320);
and U159 (N_159,N_27,In_98);
or U160 (N_160,N_120,N_106);
and U161 (N_161,N_97,In_322);
nor U162 (N_162,N_98,In_142);
nand U163 (N_163,In_260,N_101);
nand U164 (N_164,In_93,In_173);
nand U165 (N_165,N_51,N_107);
nor U166 (N_166,N_65,In_24);
and U167 (N_167,N_70,In_328);
and U168 (N_168,N_109,N_133);
or U169 (N_169,In_48,N_123);
or U170 (N_170,In_365,In_59);
nor U171 (N_171,N_61,In_89);
or U172 (N_172,In_318,In_416);
and U173 (N_173,In_281,In_220);
and U174 (N_174,N_23,N_1);
or U175 (N_175,In_330,In_425);
and U176 (N_176,In_182,In_422);
and U177 (N_177,N_148,In_233);
or U178 (N_178,In_319,N_54);
or U179 (N_179,In_295,In_14);
or U180 (N_180,N_88,In_222);
nor U181 (N_181,In_180,In_257);
nand U182 (N_182,In_336,N_141);
and U183 (N_183,N_30,In_299);
or U184 (N_184,In_397,N_48);
and U185 (N_185,In_321,N_127);
nor U186 (N_186,N_33,In_389);
and U187 (N_187,In_243,N_14);
and U188 (N_188,In_80,In_251);
nor U189 (N_189,In_496,In_171);
nor U190 (N_190,N_38,N_62);
nor U191 (N_191,In_288,In_201);
nor U192 (N_192,N_25,In_443);
nand U193 (N_193,N_146,In_146);
nor U194 (N_194,In_308,In_367);
or U195 (N_195,N_100,In_230);
nor U196 (N_196,In_85,In_178);
nor U197 (N_197,In_26,In_200);
or U198 (N_198,In_138,In_446);
nand U199 (N_199,N_40,N_75);
and U200 (N_200,N_49,In_490);
and U201 (N_201,N_144,N_199);
nor U202 (N_202,N_103,In_56);
or U203 (N_203,In_205,In_121);
nand U204 (N_204,N_39,In_428);
nand U205 (N_205,In_170,N_81);
nor U206 (N_206,In_36,N_16);
nor U207 (N_207,N_50,In_211);
nor U208 (N_208,N_130,In_293);
nand U209 (N_209,N_155,N_64);
nand U210 (N_210,N_189,In_166);
and U211 (N_211,N_129,N_116);
and U212 (N_212,In_204,In_277);
or U213 (N_213,N_131,In_453);
nand U214 (N_214,N_159,In_468);
nor U215 (N_215,N_173,In_119);
nand U216 (N_216,N_138,N_151);
nor U217 (N_217,N_119,N_92);
nand U218 (N_218,In_457,N_198);
and U219 (N_219,In_244,N_197);
and U220 (N_220,In_255,N_84);
nand U221 (N_221,In_22,In_223);
or U222 (N_222,In_45,In_256);
and U223 (N_223,In_129,N_134);
nor U224 (N_224,In_393,In_303);
and U225 (N_225,N_58,N_145);
xnor U226 (N_226,N_187,In_301);
nor U227 (N_227,In_372,In_69);
or U228 (N_228,N_121,In_371);
nand U229 (N_229,In_197,N_175);
and U230 (N_230,N_172,N_19);
and U231 (N_231,In_381,In_386);
and U232 (N_232,In_90,N_111);
or U233 (N_233,N_17,N_152);
or U234 (N_234,In_401,N_170);
and U235 (N_235,In_73,N_42);
nor U236 (N_236,In_266,N_186);
and U237 (N_237,N_140,In_187);
nor U238 (N_238,N_56,N_35);
and U239 (N_239,In_462,N_105);
nand U240 (N_240,In_110,N_63);
or U241 (N_241,N_79,In_248);
and U242 (N_242,In_291,N_157);
and U243 (N_243,N_41,N_28);
or U244 (N_244,In_343,In_412);
nand U245 (N_245,In_94,In_436);
nor U246 (N_246,In_424,In_65);
nand U247 (N_247,In_218,In_127);
nor U248 (N_248,N_10,N_160);
nand U249 (N_249,In_202,In_64);
nor U250 (N_250,N_9,N_213);
nor U251 (N_251,In_157,N_158);
or U252 (N_252,In_207,In_114);
and U253 (N_253,N_22,N_214);
and U254 (N_254,In_385,In_134);
nor U255 (N_255,In_465,In_356);
nand U256 (N_256,N_193,In_118);
or U257 (N_257,N_222,In_185);
nand U258 (N_258,N_240,In_472);
nand U259 (N_259,In_72,N_71);
or U260 (N_260,In_292,N_241);
nor U261 (N_261,N_249,N_166);
and U262 (N_262,In_42,N_149);
or U263 (N_263,N_212,N_95);
nor U264 (N_264,In_165,N_154);
nor U265 (N_265,N_196,N_80);
nand U266 (N_266,In_29,N_112);
nand U267 (N_267,N_190,In_209);
and U268 (N_268,N_183,N_174);
and U269 (N_269,N_244,N_167);
nor U270 (N_270,In_245,In_162);
or U271 (N_271,N_46,N_223);
nor U272 (N_272,N_2,N_245);
xor U273 (N_273,In_189,In_408);
nand U274 (N_274,N_55,N_194);
nand U275 (N_275,N_72,In_113);
or U276 (N_276,In_450,In_242);
nor U277 (N_277,N_118,N_68);
or U278 (N_278,In_467,N_150);
and U279 (N_279,In_87,N_169);
or U280 (N_280,In_214,N_132);
nor U281 (N_281,N_45,In_21);
nand U282 (N_282,N_182,N_82);
nand U283 (N_283,In_150,N_234);
nor U284 (N_284,In_8,In_280);
or U285 (N_285,In_2,N_117);
and U286 (N_286,In_10,N_229);
nor U287 (N_287,In_487,In_237);
and U288 (N_288,In_228,N_200);
nor U289 (N_289,N_237,N_153);
nor U290 (N_290,In_353,In_116);
nand U291 (N_291,In_49,N_243);
nor U292 (N_292,N_115,N_238);
and U293 (N_293,N_248,N_74);
nand U294 (N_294,N_94,In_262);
nand U295 (N_295,In_442,In_3);
nand U296 (N_296,N_192,N_114);
nor U297 (N_297,N_235,N_206);
or U298 (N_298,N_239,N_178);
or U299 (N_299,In_275,In_115);
nor U300 (N_300,In_79,N_108);
or U301 (N_301,N_204,In_439);
nor U302 (N_302,N_44,N_215);
or U303 (N_303,N_288,In_332);
and U304 (N_304,In_5,In_235);
and U305 (N_305,In_78,In_354);
nand U306 (N_306,N_12,N_278);
and U307 (N_307,N_208,N_162);
or U308 (N_308,In_37,In_151);
or U309 (N_309,In_396,N_221);
nor U310 (N_310,In_17,N_287);
and U311 (N_311,N_217,N_36);
nor U312 (N_312,In_399,N_277);
nor U313 (N_313,N_293,N_180);
nor U314 (N_314,In_388,N_78);
nor U315 (N_315,N_104,In_95);
nor U316 (N_316,N_281,N_225);
and U317 (N_317,N_224,N_26);
or U318 (N_318,N_252,N_126);
and U319 (N_319,In_186,N_282);
nor U320 (N_320,N_139,In_240);
or U321 (N_321,In_475,N_210);
nor U322 (N_322,N_143,In_311);
or U323 (N_323,N_279,N_191);
or U324 (N_324,N_299,N_220);
nand U325 (N_325,In_102,In_384);
or U326 (N_326,N_271,N_102);
nand U327 (N_327,N_272,N_247);
or U328 (N_328,In_302,N_289);
nand U329 (N_329,N_254,N_230);
nand U330 (N_330,In_455,N_216);
nand U331 (N_331,N_47,N_269);
nor U332 (N_332,N_262,In_70);
and U333 (N_333,N_202,N_135);
and U334 (N_334,N_264,N_246);
nand U335 (N_335,In_91,N_207);
and U336 (N_336,N_176,In_342);
nor U337 (N_337,In_438,In_161);
or U338 (N_338,N_179,N_242);
nand U339 (N_339,In_148,In_474);
or U340 (N_340,N_53,N_168);
or U341 (N_341,N_283,N_263);
and U342 (N_342,N_253,N_231);
or U343 (N_343,N_292,In_323);
or U344 (N_344,N_261,In_225);
or U345 (N_345,N_99,N_291);
nand U346 (N_346,N_274,N_171);
and U347 (N_347,In_103,In_184);
or U348 (N_348,In_232,In_106);
nand U349 (N_349,In_344,N_11);
nand U350 (N_350,In_258,N_236);
nor U351 (N_351,In_375,N_270);
nand U352 (N_352,N_285,N_218);
nand U353 (N_353,N_284,N_290);
nand U354 (N_354,N_309,N_205);
nor U355 (N_355,In_181,N_347);
or U356 (N_356,In_493,N_300);
nor U357 (N_357,In_6,N_306);
or U358 (N_358,In_317,N_76);
and U359 (N_359,In_495,In_316);
nand U360 (N_360,N_335,N_346);
or U361 (N_361,N_345,N_294);
or U362 (N_362,N_320,In_125);
nand U363 (N_363,N_73,N_165);
or U364 (N_364,N_336,N_255);
nor U365 (N_365,N_341,In_398);
and U366 (N_366,N_273,N_295);
and U367 (N_367,N_156,N_227);
or U368 (N_368,N_317,In_143);
and U369 (N_369,N_310,In_68);
or U370 (N_370,N_177,N_276);
or U371 (N_371,N_93,N_296);
or U372 (N_372,In_471,N_298);
nand U373 (N_373,N_137,N_203);
and U374 (N_374,In_417,In_335);
or U375 (N_375,N_188,N_59);
and U376 (N_376,N_7,N_342);
nand U377 (N_377,In_104,N_260);
nand U378 (N_378,In_203,N_301);
or U379 (N_379,N_297,N_251);
nor U380 (N_380,N_316,N_313);
nor U381 (N_381,N_329,N_331);
nor U382 (N_382,In_241,N_185);
nor U383 (N_383,N_315,N_307);
and U384 (N_384,N_267,N_330);
or U385 (N_385,In_139,N_311);
nor U386 (N_386,N_163,N_136);
nor U387 (N_387,N_337,N_184);
and U388 (N_388,N_124,N_195);
and U389 (N_389,N_339,N_256);
xor U390 (N_390,In_247,In_492);
and U391 (N_391,N_319,N_303);
or U392 (N_392,In_345,N_258);
nor U393 (N_393,N_209,N_164);
or U394 (N_394,N_250,N_226);
nor U395 (N_395,N_304,N_275);
nand U396 (N_396,N_328,N_327);
nor U397 (N_397,N_181,N_325);
nor U398 (N_398,N_110,N_305);
and U399 (N_399,N_265,N_340);
and U400 (N_400,N_113,N_377);
nand U401 (N_401,N_383,In_158);
and U402 (N_402,N_369,In_410);
nor U403 (N_403,N_392,N_384);
and U404 (N_404,N_378,In_441);
nand U405 (N_405,N_232,N_302);
nand U406 (N_406,N_366,N_380);
and U407 (N_407,In_188,N_390);
or U408 (N_408,N_374,N_322);
or U409 (N_409,N_333,N_259);
or U410 (N_410,N_350,N_338);
nand U411 (N_411,N_372,N_13);
nand U412 (N_412,N_352,N_360);
nand U413 (N_413,N_375,In_494);
nor U414 (N_414,N_318,N_353);
xor U415 (N_415,N_394,N_228);
nand U416 (N_416,N_128,N_363);
and U417 (N_417,N_57,N_397);
or U418 (N_418,N_348,N_362);
xnor U419 (N_419,N_386,N_356);
or U420 (N_420,N_398,N_381);
nand U421 (N_421,N_365,N_268);
xnor U422 (N_422,N_389,N_326);
nand U423 (N_423,N_391,N_344);
and U424 (N_424,N_349,N_395);
and U425 (N_425,N_393,N_379);
or U426 (N_426,N_388,N_233);
nand U427 (N_427,N_368,In_160);
and U428 (N_428,N_357,N_332);
nand U429 (N_429,In_305,In_107);
nor U430 (N_430,N_364,N_359);
or U431 (N_431,N_373,N_396);
or U432 (N_432,N_385,N_351);
xor U433 (N_433,N_321,N_32);
nand U434 (N_434,N_201,N_355);
and U435 (N_435,N_122,N_219);
and U436 (N_436,N_161,N_370);
nand U437 (N_437,N_387,N_367);
nand U438 (N_438,In_498,N_280);
nand U439 (N_439,N_286,N_358);
and U440 (N_440,N_376,N_361);
and U441 (N_441,N_354,N_371);
and U442 (N_442,N_323,In_82);
nand U443 (N_443,In_97,N_343);
or U444 (N_444,N_324,N_382);
or U445 (N_445,N_314,N_308);
nor U446 (N_446,N_266,N_312);
xnor U447 (N_447,In_466,N_257);
nor U448 (N_448,N_334,N_399);
and U449 (N_449,N_211,In_333);
or U450 (N_450,N_443,N_449);
nor U451 (N_451,N_427,N_407);
or U452 (N_452,N_416,N_428);
or U453 (N_453,N_418,N_431);
and U454 (N_454,N_406,N_442);
nor U455 (N_455,N_435,N_441);
nor U456 (N_456,N_439,N_409);
or U457 (N_457,N_448,N_400);
nor U458 (N_458,N_447,N_417);
xor U459 (N_459,N_433,N_426);
nand U460 (N_460,N_425,N_429);
nor U461 (N_461,N_436,N_445);
and U462 (N_462,N_432,N_415);
nor U463 (N_463,N_413,N_414);
nand U464 (N_464,N_444,N_410);
and U465 (N_465,N_405,N_430);
nand U466 (N_466,N_422,N_423);
or U467 (N_467,N_420,N_440);
or U468 (N_468,N_401,N_411);
and U469 (N_469,N_424,N_402);
or U470 (N_470,N_437,N_412);
or U471 (N_471,N_434,N_438);
or U472 (N_472,N_404,N_421);
and U473 (N_473,N_419,N_446);
nor U474 (N_474,N_408,N_403);
and U475 (N_475,N_432,N_442);
nor U476 (N_476,N_424,N_433);
or U477 (N_477,N_443,N_417);
or U478 (N_478,N_432,N_445);
nand U479 (N_479,N_401,N_400);
or U480 (N_480,N_443,N_414);
or U481 (N_481,N_438,N_410);
nand U482 (N_482,N_402,N_401);
nand U483 (N_483,N_401,N_404);
or U484 (N_484,N_425,N_414);
or U485 (N_485,N_431,N_429);
or U486 (N_486,N_401,N_449);
nor U487 (N_487,N_402,N_437);
nor U488 (N_488,N_405,N_416);
nand U489 (N_489,N_447,N_403);
and U490 (N_490,N_433,N_420);
nor U491 (N_491,N_415,N_401);
or U492 (N_492,N_416,N_436);
nand U493 (N_493,N_421,N_436);
or U494 (N_494,N_438,N_443);
or U495 (N_495,N_427,N_408);
nor U496 (N_496,N_425,N_441);
or U497 (N_497,N_427,N_412);
and U498 (N_498,N_424,N_430);
nand U499 (N_499,N_434,N_442);
nor U500 (N_500,N_470,N_462);
and U501 (N_501,N_473,N_475);
or U502 (N_502,N_457,N_460);
or U503 (N_503,N_497,N_468);
and U504 (N_504,N_499,N_489);
nor U505 (N_505,N_471,N_461);
nand U506 (N_506,N_485,N_459);
and U507 (N_507,N_456,N_480);
nor U508 (N_508,N_454,N_492);
and U509 (N_509,N_491,N_479);
or U510 (N_510,N_477,N_464);
nor U511 (N_511,N_469,N_481);
nor U512 (N_512,N_494,N_474);
and U513 (N_513,N_458,N_467);
xor U514 (N_514,N_498,N_487);
and U515 (N_515,N_472,N_484);
and U516 (N_516,N_495,N_450);
nand U517 (N_517,N_483,N_463);
nor U518 (N_518,N_488,N_465);
nand U519 (N_519,N_490,N_452);
nand U520 (N_520,N_486,N_451);
nor U521 (N_521,N_466,N_496);
or U522 (N_522,N_478,N_493);
nor U523 (N_523,N_455,N_476);
or U524 (N_524,N_453,N_482);
or U525 (N_525,N_477,N_469);
or U526 (N_526,N_492,N_495);
and U527 (N_527,N_464,N_456);
xor U528 (N_528,N_493,N_459);
nand U529 (N_529,N_454,N_450);
nor U530 (N_530,N_494,N_475);
nor U531 (N_531,N_458,N_456);
nor U532 (N_532,N_458,N_486);
or U533 (N_533,N_470,N_476);
or U534 (N_534,N_450,N_482);
and U535 (N_535,N_469,N_499);
nand U536 (N_536,N_498,N_482);
nor U537 (N_537,N_492,N_469);
or U538 (N_538,N_453,N_481);
and U539 (N_539,N_453,N_451);
nor U540 (N_540,N_461,N_496);
or U541 (N_541,N_469,N_453);
nor U542 (N_542,N_461,N_476);
or U543 (N_543,N_495,N_474);
nor U544 (N_544,N_486,N_460);
nand U545 (N_545,N_499,N_456);
nand U546 (N_546,N_473,N_479);
nand U547 (N_547,N_458,N_451);
or U548 (N_548,N_475,N_477);
nor U549 (N_549,N_474,N_465);
nor U550 (N_550,N_501,N_529);
and U551 (N_551,N_505,N_538);
nand U552 (N_552,N_520,N_543);
or U553 (N_553,N_542,N_527);
and U554 (N_554,N_526,N_506);
nor U555 (N_555,N_544,N_546);
nand U556 (N_556,N_533,N_509);
nor U557 (N_557,N_502,N_504);
nor U558 (N_558,N_511,N_531);
or U559 (N_559,N_540,N_534);
nand U560 (N_560,N_525,N_548);
or U561 (N_561,N_512,N_541);
and U562 (N_562,N_539,N_530);
nand U563 (N_563,N_537,N_507);
nor U564 (N_564,N_514,N_522);
nor U565 (N_565,N_508,N_503);
and U566 (N_566,N_513,N_516);
and U567 (N_567,N_519,N_523);
or U568 (N_568,N_536,N_524);
nor U569 (N_569,N_528,N_532);
nor U570 (N_570,N_549,N_500);
nand U571 (N_571,N_515,N_518);
or U572 (N_572,N_545,N_521);
xor U573 (N_573,N_547,N_510);
xnor U574 (N_574,N_535,N_517);
or U575 (N_575,N_512,N_503);
or U576 (N_576,N_510,N_520);
nor U577 (N_577,N_521,N_514);
and U578 (N_578,N_500,N_545);
nand U579 (N_579,N_528,N_539);
nor U580 (N_580,N_541,N_532);
nand U581 (N_581,N_546,N_533);
and U582 (N_582,N_506,N_516);
or U583 (N_583,N_515,N_516);
nand U584 (N_584,N_522,N_515);
nand U585 (N_585,N_509,N_519);
or U586 (N_586,N_501,N_520);
or U587 (N_587,N_537,N_536);
or U588 (N_588,N_533,N_541);
or U589 (N_589,N_509,N_543);
and U590 (N_590,N_513,N_520);
and U591 (N_591,N_523,N_522);
and U592 (N_592,N_505,N_512);
and U593 (N_593,N_526,N_516);
or U594 (N_594,N_530,N_537);
or U595 (N_595,N_544,N_507);
or U596 (N_596,N_535,N_540);
nor U597 (N_597,N_539,N_531);
and U598 (N_598,N_540,N_523);
nor U599 (N_599,N_508,N_516);
xor U600 (N_600,N_553,N_599);
and U601 (N_601,N_597,N_573);
nor U602 (N_602,N_578,N_565);
nand U603 (N_603,N_576,N_592);
nor U604 (N_604,N_588,N_585);
xor U605 (N_605,N_567,N_550);
nor U606 (N_606,N_561,N_584);
nor U607 (N_607,N_580,N_563);
and U608 (N_608,N_569,N_555);
or U609 (N_609,N_568,N_590);
nor U610 (N_610,N_586,N_562);
and U611 (N_611,N_566,N_572);
nand U612 (N_612,N_552,N_559);
nand U613 (N_613,N_595,N_594);
or U614 (N_614,N_558,N_596);
or U615 (N_615,N_581,N_591);
or U616 (N_616,N_570,N_589);
and U617 (N_617,N_556,N_575);
nand U618 (N_618,N_554,N_593);
nand U619 (N_619,N_557,N_598);
nand U620 (N_620,N_571,N_587);
nor U621 (N_621,N_579,N_564);
nand U622 (N_622,N_583,N_577);
nor U623 (N_623,N_551,N_582);
and U624 (N_624,N_560,N_574);
nor U625 (N_625,N_564,N_572);
and U626 (N_626,N_558,N_585);
and U627 (N_627,N_575,N_597);
nor U628 (N_628,N_573,N_550);
nand U629 (N_629,N_588,N_555);
nand U630 (N_630,N_590,N_588);
nor U631 (N_631,N_569,N_595);
or U632 (N_632,N_592,N_559);
or U633 (N_633,N_568,N_586);
or U634 (N_634,N_595,N_563);
nand U635 (N_635,N_594,N_560);
nor U636 (N_636,N_588,N_589);
nor U637 (N_637,N_592,N_562);
nand U638 (N_638,N_554,N_596);
or U639 (N_639,N_557,N_589);
or U640 (N_640,N_568,N_588);
nor U641 (N_641,N_567,N_581);
and U642 (N_642,N_559,N_598);
or U643 (N_643,N_598,N_560);
or U644 (N_644,N_579,N_555);
nand U645 (N_645,N_556,N_585);
and U646 (N_646,N_570,N_579);
or U647 (N_647,N_596,N_598);
or U648 (N_648,N_589,N_592);
or U649 (N_649,N_559,N_554);
or U650 (N_650,N_612,N_615);
or U651 (N_651,N_614,N_600);
or U652 (N_652,N_627,N_605);
nand U653 (N_653,N_639,N_622);
nor U654 (N_654,N_624,N_608);
or U655 (N_655,N_632,N_619);
or U656 (N_656,N_629,N_643);
or U657 (N_657,N_628,N_630);
nor U658 (N_658,N_631,N_626);
xor U659 (N_659,N_621,N_647);
nand U660 (N_660,N_611,N_613);
nand U661 (N_661,N_603,N_649);
or U662 (N_662,N_618,N_602);
and U663 (N_663,N_620,N_601);
or U664 (N_664,N_640,N_606);
or U665 (N_665,N_636,N_642);
nand U666 (N_666,N_623,N_641);
nand U667 (N_667,N_644,N_625);
nor U668 (N_668,N_604,N_648);
or U669 (N_669,N_646,N_610);
nand U670 (N_670,N_607,N_617);
nand U671 (N_671,N_634,N_633);
and U672 (N_672,N_645,N_638);
and U673 (N_673,N_616,N_609);
or U674 (N_674,N_637,N_635);
and U675 (N_675,N_617,N_626);
nand U676 (N_676,N_609,N_608);
and U677 (N_677,N_621,N_633);
or U678 (N_678,N_641,N_646);
and U679 (N_679,N_634,N_606);
nand U680 (N_680,N_647,N_611);
nand U681 (N_681,N_617,N_613);
nor U682 (N_682,N_614,N_639);
and U683 (N_683,N_605,N_648);
nand U684 (N_684,N_619,N_613);
nand U685 (N_685,N_629,N_608);
or U686 (N_686,N_626,N_648);
and U687 (N_687,N_641,N_615);
or U688 (N_688,N_649,N_624);
or U689 (N_689,N_610,N_643);
and U690 (N_690,N_646,N_633);
nand U691 (N_691,N_624,N_615);
nand U692 (N_692,N_607,N_635);
and U693 (N_693,N_633,N_607);
nand U694 (N_694,N_632,N_621);
and U695 (N_695,N_618,N_644);
nor U696 (N_696,N_639,N_644);
or U697 (N_697,N_647,N_641);
and U698 (N_698,N_638,N_632);
nor U699 (N_699,N_632,N_620);
or U700 (N_700,N_665,N_676);
or U701 (N_701,N_670,N_663);
or U702 (N_702,N_679,N_692);
nand U703 (N_703,N_659,N_654);
or U704 (N_704,N_660,N_667);
nor U705 (N_705,N_671,N_682);
and U706 (N_706,N_661,N_672);
or U707 (N_707,N_664,N_688);
and U708 (N_708,N_698,N_695);
nand U709 (N_709,N_653,N_656);
or U710 (N_710,N_655,N_669);
nand U711 (N_711,N_684,N_658);
and U712 (N_712,N_673,N_687);
nor U713 (N_713,N_677,N_683);
and U714 (N_714,N_691,N_662);
or U715 (N_715,N_675,N_652);
or U716 (N_716,N_678,N_680);
nand U717 (N_717,N_666,N_685);
nand U718 (N_718,N_697,N_674);
and U719 (N_719,N_681,N_668);
nand U720 (N_720,N_650,N_699);
or U721 (N_721,N_690,N_686);
nand U722 (N_722,N_651,N_693);
or U723 (N_723,N_657,N_696);
nand U724 (N_724,N_689,N_694);
nor U725 (N_725,N_680,N_679);
nand U726 (N_726,N_651,N_660);
and U727 (N_727,N_677,N_653);
or U728 (N_728,N_692,N_653);
or U729 (N_729,N_667,N_653);
or U730 (N_730,N_658,N_678);
nor U731 (N_731,N_688,N_692);
nor U732 (N_732,N_677,N_690);
and U733 (N_733,N_656,N_698);
nor U734 (N_734,N_653,N_689);
and U735 (N_735,N_660,N_692);
or U736 (N_736,N_653,N_661);
and U737 (N_737,N_699,N_690);
and U738 (N_738,N_689,N_666);
or U739 (N_739,N_665,N_688);
and U740 (N_740,N_668,N_673);
or U741 (N_741,N_652,N_673);
nand U742 (N_742,N_661,N_662);
nand U743 (N_743,N_652,N_660);
nor U744 (N_744,N_653,N_658);
nor U745 (N_745,N_671,N_664);
nor U746 (N_746,N_673,N_677);
or U747 (N_747,N_664,N_662);
and U748 (N_748,N_696,N_659);
and U749 (N_749,N_675,N_660);
nand U750 (N_750,N_747,N_709);
and U751 (N_751,N_727,N_713);
and U752 (N_752,N_728,N_732);
nor U753 (N_753,N_703,N_731);
nor U754 (N_754,N_741,N_723);
nor U755 (N_755,N_717,N_705);
or U756 (N_756,N_706,N_722);
or U757 (N_757,N_725,N_746);
and U758 (N_758,N_735,N_737);
nand U759 (N_759,N_738,N_724);
and U760 (N_760,N_700,N_745);
or U761 (N_761,N_730,N_721);
nand U762 (N_762,N_707,N_742);
nand U763 (N_763,N_736,N_743);
or U764 (N_764,N_749,N_716);
and U765 (N_765,N_744,N_704);
nor U766 (N_766,N_702,N_726);
nand U767 (N_767,N_729,N_708);
or U768 (N_768,N_733,N_715);
and U769 (N_769,N_718,N_714);
and U770 (N_770,N_740,N_719);
and U771 (N_771,N_720,N_739);
nor U772 (N_772,N_712,N_734);
or U773 (N_773,N_711,N_748);
and U774 (N_774,N_701,N_710);
xor U775 (N_775,N_717,N_709);
xor U776 (N_776,N_736,N_710);
nand U777 (N_777,N_701,N_740);
or U778 (N_778,N_743,N_716);
xor U779 (N_779,N_726,N_743);
nand U780 (N_780,N_724,N_710);
nand U781 (N_781,N_746,N_719);
nor U782 (N_782,N_727,N_719);
xor U783 (N_783,N_710,N_717);
nand U784 (N_784,N_731,N_715);
nor U785 (N_785,N_729,N_746);
and U786 (N_786,N_742,N_740);
nor U787 (N_787,N_716,N_746);
nor U788 (N_788,N_749,N_738);
nand U789 (N_789,N_748,N_720);
and U790 (N_790,N_725,N_712);
xnor U791 (N_791,N_703,N_706);
or U792 (N_792,N_737,N_721);
nand U793 (N_793,N_723,N_707);
nor U794 (N_794,N_728,N_713);
nand U795 (N_795,N_727,N_722);
or U796 (N_796,N_733,N_722);
nand U797 (N_797,N_728,N_722);
and U798 (N_798,N_749,N_723);
nand U799 (N_799,N_720,N_746);
or U800 (N_800,N_764,N_779);
and U801 (N_801,N_799,N_759);
or U802 (N_802,N_777,N_780);
or U803 (N_803,N_758,N_762);
and U804 (N_804,N_763,N_765);
and U805 (N_805,N_786,N_756);
nand U806 (N_806,N_794,N_751);
and U807 (N_807,N_769,N_792);
nand U808 (N_808,N_775,N_768);
nor U809 (N_809,N_789,N_793);
and U810 (N_810,N_767,N_760);
and U811 (N_811,N_788,N_784);
nand U812 (N_812,N_782,N_754);
or U813 (N_813,N_752,N_755);
and U814 (N_814,N_797,N_783);
and U815 (N_815,N_790,N_761);
and U816 (N_816,N_795,N_750);
nor U817 (N_817,N_771,N_785);
nor U818 (N_818,N_778,N_773);
nand U819 (N_819,N_796,N_772);
nand U820 (N_820,N_787,N_791);
or U821 (N_821,N_757,N_766);
nor U822 (N_822,N_776,N_798);
or U823 (N_823,N_770,N_753);
and U824 (N_824,N_781,N_774);
or U825 (N_825,N_768,N_785);
nor U826 (N_826,N_751,N_793);
nand U827 (N_827,N_785,N_786);
nor U828 (N_828,N_795,N_754);
or U829 (N_829,N_782,N_757);
nand U830 (N_830,N_798,N_783);
and U831 (N_831,N_750,N_796);
nand U832 (N_832,N_790,N_788);
nand U833 (N_833,N_770,N_791);
nor U834 (N_834,N_799,N_751);
nor U835 (N_835,N_762,N_768);
and U836 (N_836,N_780,N_765);
nand U837 (N_837,N_794,N_785);
or U838 (N_838,N_797,N_785);
nor U839 (N_839,N_792,N_752);
nand U840 (N_840,N_779,N_758);
nor U841 (N_841,N_751,N_784);
nand U842 (N_842,N_799,N_783);
or U843 (N_843,N_753,N_778);
nand U844 (N_844,N_770,N_780);
nand U845 (N_845,N_773,N_754);
or U846 (N_846,N_798,N_785);
nor U847 (N_847,N_788,N_769);
nor U848 (N_848,N_795,N_774);
nand U849 (N_849,N_795,N_764);
nor U850 (N_850,N_803,N_824);
nand U851 (N_851,N_809,N_834);
nand U852 (N_852,N_833,N_801);
and U853 (N_853,N_823,N_827);
nand U854 (N_854,N_811,N_817);
nand U855 (N_855,N_847,N_829);
nand U856 (N_856,N_846,N_818);
nor U857 (N_857,N_838,N_815);
or U858 (N_858,N_810,N_842);
nor U859 (N_859,N_844,N_819);
or U860 (N_860,N_802,N_804);
and U861 (N_861,N_835,N_826);
nor U862 (N_862,N_841,N_814);
nand U863 (N_863,N_843,N_805);
xor U864 (N_864,N_816,N_836);
or U865 (N_865,N_830,N_828);
nor U866 (N_866,N_808,N_831);
or U867 (N_867,N_812,N_848);
and U868 (N_868,N_825,N_820);
nor U869 (N_869,N_806,N_822);
or U870 (N_870,N_840,N_845);
nand U871 (N_871,N_807,N_821);
or U872 (N_872,N_832,N_813);
or U873 (N_873,N_800,N_837);
nor U874 (N_874,N_839,N_849);
xor U875 (N_875,N_836,N_846);
nor U876 (N_876,N_830,N_838);
or U877 (N_877,N_839,N_815);
and U878 (N_878,N_835,N_848);
or U879 (N_879,N_848,N_833);
nor U880 (N_880,N_831,N_832);
and U881 (N_881,N_833,N_840);
nand U882 (N_882,N_821,N_814);
nor U883 (N_883,N_832,N_804);
nand U884 (N_884,N_835,N_815);
nor U885 (N_885,N_833,N_829);
nand U886 (N_886,N_832,N_846);
and U887 (N_887,N_830,N_825);
or U888 (N_888,N_837,N_831);
and U889 (N_889,N_834,N_831);
nand U890 (N_890,N_813,N_829);
nand U891 (N_891,N_806,N_828);
and U892 (N_892,N_805,N_845);
xnor U893 (N_893,N_811,N_827);
or U894 (N_894,N_804,N_837);
and U895 (N_895,N_812,N_816);
and U896 (N_896,N_801,N_823);
nand U897 (N_897,N_825,N_803);
or U898 (N_898,N_840,N_808);
nor U899 (N_899,N_835,N_828);
nor U900 (N_900,N_872,N_860);
xnor U901 (N_901,N_867,N_857);
and U902 (N_902,N_882,N_884);
xnor U903 (N_903,N_873,N_878);
nand U904 (N_904,N_861,N_887);
and U905 (N_905,N_885,N_853);
nand U906 (N_906,N_856,N_854);
or U907 (N_907,N_863,N_877);
nor U908 (N_908,N_869,N_880);
and U909 (N_909,N_896,N_862);
or U910 (N_910,N_895,N_875);
or U911 (N_911,N_881,N_866);
nand U912 (N_912,N_893,N_876);
and U913 (N_913,N_889,N_858);
nand U914 (N_914,N_898,N_894);
nor U915 (N_915,N_851,N_859);
or U916 (N_916,N_891,N_883);
xnor U917 (N_917,N_850,N_864);
nand U918 (N_918,N_888,N_892);
nand U919 (N_919,N_870,N_879);
xor U920 (N_920,N_871,N_852);
or U921 (N_921,N_874,N_868);
and U922 (N_922,N_886,N_865);
nor U923 (N_923,N_897,N_899);
and U924 (N_924,N_890,N_855);
and U925 (N_925,N_897,N_863);
nand U926 (N_926,N_866,N_885);
nor U927 (N_927,N_884,N_887);
nor U928 (N_928,N_884,N_872);
nor U929 (N_929,N_899,N_872);
nor U930 (N_930,N_856,N_874);
nor U931 (N_931,N_850,N_894);
and U932 (N_932,N_865,N_882);
nor U933 (N_933,N_889,N_898);
nand U934 (N_934,N_864,N_897);
and U935 (N_935,N_852,N_859);
xnor U936 (N_936,N_854,N_893);
nand U937 (N_937,N_858,N_894);
and U938 (N_938,N_867,N_866);
xor U939 (N_939,N_897,N_898);
nand U940 (N_940,N_893,N_855);
and U941 (N_941,N_888,N_890);
or U942 (N_942,N_862,N_861);
or U943 (N_943,N_869,N_872);
xor U944 (N_944,N_884,N_879);
nand U945 (N_945,N_892,N_896);
and U946 (N_946,N_855,N_894);
and U947 (N_947,N_887,N_865);
or U948 (N_948,N_878,N_882);
or U949 (N_949,N_875,N_899);
xnor U950 (N_950,N_945,N_915);
nand U951 (N_951,N_949,N_916);
nand U952 (N_952,N_914,N_912);
or U953 (N_953,N_921,N_929);
nand U954 (N_954,N_942,N_941);
and U955 (N_955,N_908,N_905);
or U956 (N_956,N_906,N_901);
and U957 (N_957,N_922,N_931);
nand U958 (N_958,N_902,N_903);
xor U959 (N_959,N_932,N_940);
nor U960 (N_960,N_930,N_936);
and U961 (N_961,N_927,N_935);
or U962 (N_962,N_944,N_917);
nand U963 (N_963,N_928,N_919);
nor U964 (N_964,N_926,N_933);
xor U965 (N_965,N_910,N_943);
or U966 (N_966,N_911,N_923);
and U967 (N_967,N_907,N_937);
or U968 (N_968,N_946,N_920);
and U969 (N_969,N_938,N_948);
nor U970 (N_970,N_934,N_918);
and U971 (N_971,N_913,N_900);
or U972 (N_972,N_909,N_947);
and U973 (N_973,N_939,N_925);
and U974 (N_974,N_924,N_904);
nand U975 (N_975,N_910,N_934);
nand U976 (N_976,N_921,N_941);
or U977 (N_977,N_935,N_933);
and U978 (N_978,N_922,N_912);
xor U979 (N_979,N_924,N_914);
nor U980 (N_980,N_922,N_918);
or U981 (N_981,N_934,N_920);
and U982 (N_982,N_914,N_928);
and U983 (N_983,N_900,N_938);
and U984 (N_984,N_923,N_946);
xor U985 (N_985,N_907,N_941);
xnor U986 (N_986,N_913,N_948);
nand U987 (N_987,N_929,N_926);
nor U988 (N_988,N_923,N_919);
nor U989 (N_989,N_916,N_914);
nor U990 (N_990,N_930,N_918);
or U991 (N_991,N_925,N_948);
or U992 (N_992,N_941,N_928);
nand U993 (N_993,N_920,N_909);
nand U994 (N_994,N_948,N_904);
nor U995 (N_995,N_947,N_934);
nor U996 (N_996,N_924,N_902);
nand U997 (N_997,N_930,N_935);
nor U998 (N_998,N_930,N_904);
nor U999 (N_999,N_925,N_947);
nor U1000 (N_1000,N_968,N_984);
nand U1001 (N_1001,N_951,N_985);
or U1002 (N_1002,N_960,N_979);
nor U1003 (N_1003,N_976,N_950);
nand U1004 (N_1004,N_970,N_982);
nand U1005 (N_1005,N_994,N_953);
nand U1006 (N_1006,N_978,N_959);
nand U1007 (N_1007,N_992,N_964);
and U1008 (N_1008,N_969,N_987);
or U1009 (N_1009,N_958,N_961);
or U1010 (N_1010,N_952,N_999);
or U1011 (N_1011,N_972,N_991);
nand U1012 (N_1012,N_990,N_993);
nand U1013 (N_1013,N_986,N_965);
xnor U1014 (N_1014,N_975,N_957);
nand U1015 (N_1015,N_981,N_988);
nand U1016 (N_1016,N_983,N_980);
or U1017 (N_1017,N_996,N_998);
or U1018 (N_1018,N_971,N_974);
nand U1019 (N_1019,N_977,N_997);
nor U1020 (N_1020,N_962,N_973);
xnor U1021 (N_1021,N_995,N_955);
or U1022 (N_1022,N_963,N_956);
and U1023 (N_1023,N_989,N_954);
nor U1024 (N_1024,N_966,N_967);
or U1025 (N_1025,N_980,N_956);
nand U1026 (N_1026,N_979,N_955);
and U1027 (N_1027,N_997,N_996);
nor U1028 (N_1028,N_995,N_982);
and U1029 (N_1029,N_984,N_964);
and U1030 (N_1030,N_992,N_957);
and U1031 (N_1031,N_997,N_979);
and U1032 (N_1032,N_980,N_979);
or U1033 (N_1033,N_978,N_997);
and U1034 (N_1034,N_971,N_992);
or U1035 (N_1035,N_977,N_987);
or U1036 (N_1036,N_992,N_955);
nor U1037 (N_1037,N_987,N_986);
or U1038 (N_1038,N_960,N_964);
or U1039 (N_1039,N_972,N_981);
nor U1040 (N_1040,N_958,N_966);
nor U1041 (N_1041,N_975,N_981);
and U1042 (N_1042,N_964,N_991);
nand U1043 (N_1043,N_978,N_991);
nand U1044 (N_1044,N_984,N_951);
xor U1045 (N_1045,N_989,N_998);
nand U1046 (N_1046,N_968,N_958);
and U1047 (N_1047,N_998,N_963);
nand U1048 (N_1048,N_974,N_972);
nor U1049 (N_1049,N_981,N_950);
or U1050 (N_1050,N_1047,N_1021);
nand U1051 (N_1051,N_1017,N_1044);
nand U1052 (N_1052,N_1004,N_1002);
nand U1053 (N_1053,N_1032,N_1012);
nor U1054 (N_1054,N_1034,N_1046);
or U1055 (N_1055,N_1022,N_1041);
or U1056 (N_1056,N_1031,N_1033);
or U1057 (N_1057,N_1000,N_1018);
and U1058 (N_1058,N_1042,N_1048);
nand U1059 (N_1059,N_1015,N_1005);
and U1060 (N_1060,N_1026,N_1049);
nor U1061 (N_1061,N_1006,N_1008);
and U1062 (N_1062,N_1009,N_1013);
nor U1063 (N_1063,N_1037,N_1003);
nor U1064 (N_1064,N_1027,N_1011);
or U1065 (N_1065,N_1001,N_1024);
and U1066 (N_1066,N_1028,N_1040);
and U1067 (N_1067,N_1043,N_1025);
or U1068 (N_1068,N_1019,N_1020);
nor U1069 (N_1069,N_1036,N_1016);
nor U1070 (N_1070,N_1023,N_1038);
or U1071 (N_1071,N_1039,N_1035);
or U1072 (N_1072,N_1007,N_1014);
nor U1073 (N_1073,N_1030,N_1045);
or U1074 (N_1074,N_1029,N_1010);
or U1075 (N_1075,N_1028,N_1021);
xor U1076 (N_1076,N_1042,N_1000);
xor U1077 (N_1077,N_1025,N_1034);
nor U1078 (N_1078,N_1044,N_1047);
nand U1079 (N_1079,N_1034,N_1006);
nand U1080 (N_1080,N_1001,N_1007);
nor U1081 (N_1081,N_1010,N_1040);
or U1082 (N_1082,N_1010,N_1020);
and U1083 (N_1083,N_1024,N_1049);
nor U1084 (N_1084,N_1034,N_1041);
nor U1085 (N_1085,N_1049,N_1015);
nor U1086 (N_1086,N_1014,N_1042);
and U1087 (N_1087,N_1041,N_1002);
or U1088 (N_1088,N_1026,N_1039);
nor U1089 (N_1089,N_1011,N_1001);
or U1090 (N_1090,N_1043,N_1001);
or U1091 (N_1091,N_1029,N_1037);
and U1092 (N_1092,N_1013,N_1029);
or U1093 (N_1093,N_1035,N_1041);
and U1094 (N_1094,N_1005,N_1023);
nand U1095 (N_1095,N_1018,N_1038);
and U1096 (N_1096,N_1007,N_1021);
and U1097 (N_1097,N_1047,N_1032);
and U1098 (N_1098,N_1016,N_1010);
or U1099 (N_1099,N_1020,N_1048);
or U1100 (N_1100,N_1069,N_1092);
nand U1101 (N_1101,N_1084,N_1074);
nand U1102 (N_1102,N_1055,N_1053);
nand U1103 (N_1103,N_1082,N_1056);
nand U1104 (N_1104,N_1064,N_1081);
and U1105 (N_1105,N_1088,N_1091);
and U1106 (N_1106,N_1051,N_1054);
and U1107 (N_1107,N_1073,N_1099);
nand U1108 (N_1108,N_1080,N_1086);
nand U1109 (N_1109,N_1059,N_1066);
nor U1110 (N_1110,N_1095,N_1052);
or U1111 (N_1111,N_1057,N_1070);
nand U1112 (N_1112,N_1050,N_1079);
nand U1113 (N_1113,N_1058,N_1085);
nor U1114 (N_1114,N_1071,N_1089);
or U1115 (N_1115,N_1062,N_1083);
nor U1116 (N_1116,N_1090,N_1093);
nand U1117 (N_1117,N_1072,N_1068);
or U1118 (N_1118,N_1077,N_1075);
nand U1119 (N_1119,N_1078,N_1065);
nor U1120 (N_1120,N_1087,N_1063);
or U1121 (N_1121,N_1096,N_1067);
and U1122 (N_1122,N_1098,N_1097);
nor U1123 (N_1123,N_1076,N_1094);
nand U1124 (N_1124,N_1061,N_1060);
or U1125 (N_1125,N_1066,N_1099);
nor U1126 (N_1126,N_1055,N_1073);
nand U1127 (N_1127,N_1055,N_1089);
or U1128 (N_1128,N_1076,N_1095);
nand U1129 (N_1129,N_1053,N_1076);
and U1130 (N_1130,N_1071,N_1088);
and U1131 (N_1131,N_1081,N_1060);
nand U1132 (N_1132,N_1068,N_1073);
and U1133 (N_1133,N_1078,N_1060);
and U1134 (N_1134,N_1079,N_1072);
nor U1135 (N_1135,N_1092,N_1096);
and U1136 (N_1136,N_1092,N_1099);
nand U1137 (N_1137,N_1094,N_1077);
and U1138 (N_1138,N_1070,N_1093);
and U1139 (N_1139,N_1081,N_1082);
nor U1140 (N_1140,N_1084,N_1099);
nor U1141 (N_1141,N_1093,N_1055);
and U1142 (N_1142,N_1056,N_1067);
nand U1143 (N_1143,N_1053,N_1087);
or U1144 (N_1144,N_1098,N_1072);
nor U1145 (N_1145,N_1087,N_1093);
nand U1146 (N_1146,N_1094,N_1057);
or U1147 (N_1147,N_1091,N_1055);
and U1148 (N_1148,N_1075,N_1083);
nand U1149 (N_1149,N_1083,N_1096);
or U1150 (N_1150,N_1125,N_1134);
nor U1151 (N_1151,N_1101,N_1105);
nand U1152 (N_1152,N_1104,N_1142);
or U1153 (N_1153,N_1127,N_1141);
and U1154 (N_1154,N_1122,N_1123);
xnor U1155 (N_1155,N_1136,N_1111);
nand U1156 (N_1156,N_1118,N_1124);
and U1157 (N_1157,N_1139,N_1148);
nand U1158 (N_1158,N_1138,N_1106);
nand U1159 (N_1159,N_1113,N_1147);
and U1160 (N_1160,N_1137,N_1112);
or U1161 (N_1161,N_1110,N_1145);
nor U1162 (N_1162,N_1117,N_1130);
and U1163 (N_1163,N_1100,N_1131);
or U1164 (N_1164,N_1133,N_1109);
nor U1165 (N_1165,N_1103,N_1108);
and U1166 (N_1166,N_1149,N_1132);
nand U1167 (N_1167,N_1126,N_1135);
or U1168 (N_1168,N_1116,N_1144);
or U1169 (N_1169,N_1140,N_1119);
xnor U1170 (N_1170,N_1107,N_1102);
nor U1171 (N_1171,N_1143,N_1120);
or U1172 (N_1172,N_1146,N_1121);
nand U1173 (N_1173,N_1115,N_1114);
or U1174 (N_1174,N_1129,N_1128);
and U1175 (N_1175,N_1136,N_1145);
nor U1176 (N_1176,N_1114,N_1118);
nand U1177 (N_1177,N_1131,N_1139);
nand U1178 (N_1178,N_1117,N_1118);
nand U1179 (N_1179,N_1126,N_1129);
nand U1180 (N_1180,N_1126,N_1112);
or U1181 (N_1181,N_1103,N_1136);
xor U1182 (N_1182,N_1113,N_1145);
or U1183 (N_1183,N_1136,N_1143);
or U1184 (N_1184,N_1116,N_1122);
and U1185 (N_1185,N_1141,N_1147);
and U1186 (N_1186,N_1108,N_1133);
or U1187 (N_1187,N_1131,N_1130);
nand U1188 (N_1188,N_1121,N_1136);
nand U1189 (N_1189,N_1118,N_1109);
and U1190 (N_1190,N_1104,N_1145);
nand U1191 (N_1191,N_1101,N_1113);
and U1192 (N_1192,N_1115,N_1112);
and U1193 (N_1193,N_1113,N_1120);
nor U1194 (N_1194,N_1105,N_1114);
nor U1195 (N_1195,N_1122,N_1110);
or U1196 (N_1196,N_1136,N_1114);
or U1197 (N_1197,N_1133,N_1104);
nor U1198 (N_1198,N_1133,N_1129);
and U1199 (N_1199,N_1122,N_1143);
and U1200 (N_1200,N_1199,N_1184);
or U1201 (N_1201,N_1155,N_1179);
nand U1202 (N_1202,N_1187,N_1167);
or U1203 (N_1203,N_1168,N_1174);
or U1204 (N_1204,N_1152,N_1151);
nand U1205 (N_1205,N_1176,N_1177);
nor U1206 (N_1206,N_1185,N_1169);
nand U1207 (N_1207,N_1191,N_1183);
or U1208 (N_1208,N_1165,N_1156);
or U1209 (N_1209,N_1162,N_1186);
nand U1210 (N_1210,N_1159,N_1195);
or U1211 (N_1211,N_1161,N_1175);
nand U1212 (N_1212,N_1150,N_1189);
and U1213 (N_1213,N_1154,N_1178);
nor U1214 (N_1214,N_1158,N_1194);
nand U1215 (N_1215,N_1164,N_1180);
nand U1216 (N_1216,N_1198,N_1170);
and U1217 (N_1217,N_1153,N_1163);
nor U1218 (N_1218,N_1166,N_1196);
nor U1219 (N_1219,N_1193,N_1190);
and U1220 (N_1220,N_1182,N_1171);
nand U1221 (N_1221,N_1192,N_1173);
or U1222 (N_1222,N_1188,N_1157);
nand U1223 (N_1223,N_1172,N_1197);
nor U1224 (N_1224,N_1181,N_1160);
nand U1225 (N_1225,N_1191,N_1162);
or U1226 (N_1226,N_1199,N_1154);
nor U1227 (N_1227,N_1189,N_1191);
nand U1228 (N_1228,N_1181,N_1195);
nand U1229 (N_1229,N_1198,N_1195);
nor U1230 (N_1230,N_1185,N_1191);
xor U1231 (N_1231,N_1199,N_1163);
and U1232 (N_1232,N_1199,N_1194);
nand U1233 (N_1233,N_1161,N_1151);
or U1234 (N_1234,N_1190,N_1154);
or U1235 (N_1235,N_1183,N_1190);
or U1236 (N_1236,N_1158,N_1182);
and U1237 (N_1237,N_1185,N_1194);
and U1238 (N_1238,N_1151,N_1191);
nand U1239 (N_1239,N_1154,N_1157);
and U1240 (N_1240,N_1167,N_1170);
or U1241 (N_1241,N_1169,N_1184);
or U1242 (N_1242,N_1174,N_1171);
nor U1243 (N_1243,N_1167,N_1190);
or U1244 (N_1244,N_1155,N_1189);
nand U1245 (N_1245,N_1157,N_1160);
nor U1246 (N_1246,N_1182,N_1154);
nand U1247 (N_1247,N_1194,N_1157);
nor U1248 (N_1248,N_1168,N_1158);
nand U1249 (N_1249,N_1171,N_1195);
nand U1250 (N_1250,N_1228,N_1241);
and U1251 (N_1251,N_1232,N_1222);
nand U1252 (N_1252,N_1248,N_1242);
and U1253 (N_1253,N_1245,N_1244);
nor U1254 (N_1254,N_1230,N_1219);
nor U1255 (N_1255,N_1247,N_1240);
nand U1256 (N_1256,N_1220,N_1202);
and U1257 (N_1257,N_1238,N_1249);
nor U1258 (N_1258,N_1205,N_1208);
nor U1259 (N_1259,N_1211,N_1215);
and U1260 (N_1260,N_1233,N_1204);
nand U1261 (N_1261,N_1223,N_1212);
or U1262 (N_1262,N_1237,N_1246);
or U1263 (N_1263,N_1226,N_1214);
and U1264 (N_1264,N_1224,N_1234);
or U1265 (N_1265,N_1221,N_1200);
nand U1266 (N_1266,N_1206,N_1229);
xor U1267 (N_1267,N_1218,N_1227);
nand U1268 (N_1268,N_1217,N_1243);
nor U1269 (N_1269,N_1236,N_1225);
and U1270 (N_1270,N_1207,N_1239);
xnor U1271 (N_1271,N_1203,N_1213);
or U1272 (N_1272,N_1210,N_1231);
or U1273 (N_1273,N_1235,N_1209);
and U1274 (N_1274,N_1201,N_1216);
or U1275 (N_1275,N_1231,N_1219);
nand U1276 (N_1276,N_1213,N_1244);
nand U1277 (N_1277,N_1248,N_1236);
xor U1278 (N_1278,N_1211,N_1235);
nor U1279 (N_1279,N_1205,N_1227);
and U1280 (N_1280,N_1230,N_1234);
or U1281 (N_1281,N_1229,N_1223);
nand U1282 (N_1282,N_1202,N_1227);
nor U1283 (N_1283,N_1217,N_1207);
and U1284 (N_1284,N_1210,N_1211);
and U1285 (N_1285,N_1221,N_1222);
or U1286 (N_1286,N_1213,N_1237);
nor U1287 (N_1287,N_1245,N_1242);
nor U1288 (N_1288,N_1244,N_1205);
and U1289 (N_1289,N_1239,N_1242);
or U1290 (N_1290,N_1248,N_1233);
nand U1291 (N_1291,N_1248,N_1246);
and U1292 (N_1292,N_1229,N_1212);
or U1293 (N_1293,N_1230,N_1216);
and U1294 (N_1294,N_1234,N_1239);
nand U1295 (N_1295,N_1208,N_1241);
and U1296 (N_1296,N_1237,N_1206);
or U1297 (N_1297,N_1225,N_1237);
nor U1298 (N_1298,N_1233,N_1215);
xnor U1299 (N_1299,N_1228,N_1205);
and U1300 (N_1300,N_1282,N_1275);
xnor U1301 (N_1301,N_1296,N_1266);
and U1302 (N_1302,N_1265,N_1289);
or U1303 (N_1303,N_1270,N_1292);
and U1304 (N_1304,N_1263,N_1252);
or U1305 (N_1305,N_1253,N_1268);
nor U1306 (N_1306,N_1280,N_1278);
or U1307 (N_1307,N_1269,N_1264);
nand U1308 (N_1308,N_1288,N_1290);
nor U1309 (N_1309,N_1261,N_1294);
and U1310 (N_1310,N_1274,N_1258);
nand U1311 (N_1311,N_1254,N_1257);
nand U1312 (N_1312,N_1297,N_1281);
nor U1313 (N_1313,N_1276,N_1251);
or U1314 (N_1314,N_1260,N_1285);
and U1315 (N_1315,N_1291,N_1271);
xnor U1316 (N_1316,N_1273,N_1284);
nor U1317 (N_1317,N_1256,N_1255);
nor U1318 (N_1318,N_1267,N_1250);
or U1319 (N_1319,N_1277,N_1262);
and U1320 (N_1320,N_1299,N_1293);
and U1321 (N_1321,N_1287,N_1286);
and U1322 (N_1322,N_1272,N_1283);
and U1323 (N_1323,N_1295,N_1298);
and U1324 (N_1324,N_1279,N_1259);
nand U1325 (N_1325,N_1289,N_1282);
nor U1326 (N_1326,N_1279,N_1258);
nand U1327 (N_1327,N_1257,N_1295);
nand U1328 (N_1328,N_1273,N_1264);
and U1329 (N_1329,N_1268,N_1287);
xnor U1330 (N_1330,N_1281,N_1266);
nor U1331 (N_1331,N_1280,N_1275);
and U1332 (N_1332,N_1258,N_1295);
nand U1333 (N_1333,N_1274,N_1275);
or U1334 (N_1334,N_1266,N_1282);
nor U1335 (N_1335,N_1269,N_1261);
nor U1336 (N_1336,N_1288,N_1274);
nor U1337 (N_1337,N_1282,N_1267);
nand U1338 (N_1338,N_1271,N_1263);
xor U1339 (N_1339,N_1262,N_1251);
or U1340 (N_1340,N_1277,N_1294);
nand U1341 (N_1341,N_1296,N_1289);
nor U1342 (N_1342,N_1299,N_1263);
or U1343 (N_1343,N_1298,N_1274);
nor U1344 (N_1344,N_1279,N_1268);
or U1345 (N_1345,N_1291,N_1254);
nor U1346 (N_1346,N_1267,N_1288);
and U1347 (N_1347,N_1273,N_1280);
nor U1348 (N_1348,N_1283,N_1293);
and U1349 (N_1349,N_1294,N_1286);
nor U1350 (N_1350,N_1332,N_1330);
or U1351 (N_1351,N_1304,N_1327);
or U1352 (N_1352,N_1325,N_1334);
nand U1353 (N_1353,N_1326,N_1349);
and U1354 (N_1354,N_1348,N_1307);
xor U1355 (N_1355,N_1306,N_1303);
nor U1356 (N_1356,N_1347,N_1342);
nand U1357 (N_1357,N_1329,N_1343);
nor U1358 (N_1358,N_1320,N_1339);
xor U1359 (N_1359,N_1322,N_1316);
nand U1360 (N_1360,N_1344,N_1319);
nand U1361 (N_1361,N_1308,N_1337);
or U1362 (N_1362,N_1328,N_1310);
or U1363 (N_1363,N_1314,N_1333);
nand U1364 (N_1364,N_1341,N_1317);
and U1365 (N_1365,N_1302,N_1318);
or U1366 (N_1366,N_1340,N_1311);
and U1367 (N_1367,N_1301,N_1305);
nor U1368 (N_1368,N_1335,N_1331);
nor U1369 (N_1369,N_1345,N_1315);
and U1370 (N_1370,N_1313,N_1346);
or U1371 (N_1371,N_1336,N_1338);
and U1372 (N_1372,N_1324,N_1323);
nor U1373 (N_1373,N_1309,N_1300);
nand U1374 (N_1374,N_1312,N_1321);
nor U1375 (N_1375,N_1310,N_1326);
nand U1376 (N_1376,N_1308,N_1330);
nor U1377 (N_1377,N_1342,N_1346);
and U1378 (N_1378,N_1321,N_1338);
or U1379 (N_1379,N_1329,N_1341);
or U1380 (N_1380,N_1319,N_1337);
and U1381 (N_1381,N_1324,N_1327);
nand U1382 (N_1382,N_1339,N_1301);
or U1383 (N_1383,N_1335,N_1346);
or U1384 (N_1384,N_1308,N_1346);
and U1385 (N_1385,N_1308,N_1341);
and U1386 (N_1386,N_1300,N_1306);
and U1387 (N_1387,N_1326,N_1344);
nor U1388 (N_1388,N_1340,N_1319);
nand U1389 (N_1389,N_1339,N_1311);
nor U1390 (N_1390,N_1324,N_1341);
nand U1391 (N_1391,N_1340,N_1327);
nor U1392 (N_1392,N_1309,N_1304);
and U1393 (N_1393,N_1337,N_1313);
nor U1394 (N_1394,N_1304,N_1303);
nand U1395 (N_1395,N_1320,N_1337);
or U1396 (N_1396,N_1334,N_1326);
or U1397 (N_1397,N_1307,N_1303);
and U1398 (N_1398,N_1301,N_1348);
and U1399 (N_1399,N_1328,N_1326);
nor U1400 (N_1400,N_1364,N_1360);
nand U1401 (N_1401,N_1355,N_1362);
xnor U1402 (N_1402,N_1359,N_1386);
or U1403 (N_1403,N_1369,N_1356);
nand U1404 (N_1404,N_1393,N_1354);
or U1405 (N_1405,N_1370,N_1389);
nor U1406 (N_1406,N_1366,N_1368);
and U1407 (N_1407,N_1371,N_1361);
or U1408 (N_1408,N_1392,N_1374);
nand U1409 (N_1409,N_1373,N_1353);
nand U1410 (N_1410,N_1372,N_1378);
nand U1411 (N_1411,N_1398,N_1357);
nand U1412 (N_1412,N_1377,N_1375);
nand U1413 (N_1413,N_1391,N_1351);
nor U1414 (N_1414,N_1383,N_1376);
and U1415 (N_1415,N_1397,N_1384);
nor U1416 (N_1416,N_1381,N_1350);
or U1417 (N_1417,N_1388,N_1396);
nor U1418 (N_1418,N_1390,N_1387);
nand U1419 (N_1419,N_1363,N_1394);
or U1420 (N_1420,N_1352,N_1358);
nand U1421 (N_1421,N_1395,N_1379);
and U1422 (N_1422,N_1382,N_1365);
xnor U1423 (N_1423,N_1367,N_1385);
nand U1424 (N_1424,N_1380,N_1399);
nor U1425 (N_1425,N_1352,N_1398);
or U1426 (N_1426,N_1394,N_1377);
or U1427 (N_1427,N_1391,N_1397);
nand U1428 (N_1428,N_1359,N_1394);
or U1429 (N_1429,N_1395,N_1354);
nor U1430 (N_1430,N_1375,N_1398);
nor U1431 (N_1431,N_1388,N_1384);
and U1432 (N_1432,N_1378,N_1398);
nor U1433 (N_1433,N_1364,N_1357);
nand U1434 (N_1434,N_1356,N_1360);
nor U1435 (N_1435,N_1363,N_1395);
and U1436 (N_1436,N_1397,N_1369);
or U1437 (N_1437,N_1384,N_1369);
nor U1438 (N_1438,N_1370,N_1372);
and U1439 (N_1439,N_1393,N_1377);
or U1440 (N_1440,N_1387,N_1353);
or U1441 (N_1441,N_1381,N_1387);
and U1442 (N_1442,N_1359,N_1398);
and U1443 (N_1443,N_1351,N_1359);
or U1444 (N_1444,N_1376,N_1357);
nand U1445 (N_1445,N_1363,N_1376);
nor U1446 (N_1446,N_1396,N_1362);
and U1447 (N_1447,N_1366,N_1395);
nand U1448 (N_1448,N_1378,N_1356);
or U1449 (N_1449,N_1368,N_1396);
and U1450 (N_1450,N_1424,N_1447);
or U1451 (N_1451,N_1410,N_1427);
and U1452 (N_1452,N_1443,N_1404);
nand U1453 (N_1453,N_1445,N_1436);
and U1454 (N_1454,N_1416,N_1423);
or U1455 (N_1455,N_1432,N_1444);
and U1456 (N_1456,N_1421,N_1411);
or U1457 (N_1457,N_1446,N_1403);
and U1458 (N_1458,N_1429,N_1438);
and U1459 (N_1459,N_1435,N_1400);
or U1460 (N_1460,N_1406,N_1434);
or U1461 (N_1461,N_1431,N_1409);
and U1462 (N_1462,N_1442,N_1437);
nand U1463 (N_1463,N_1402,N_1426);
nand U1464 (N_1464,N_1439,N_1405);
and U1465 (N_1465,N_1407,N_1433);
nor U1466 (N_1466,N_1428,N_1413);
and U1467 (N_1467,N_1415,N_1408);
nand U1468 (N_1468,N_1420,N_1414);
xnor U1469 (N_1469,N_1430,N_1440);
nor U1470 (N_1470,N_1418,N_1449);
and U1471 (N_1471,N_1425,N_1419);
and U1472 (N_1472,N_1448,N_1417);
or U1473 (N_1473,N_1422,N_1412);
or U1474 (N_1474,N_1401,N_1441);
nor U1475 (N_1475,N_1446,N_1434);
or U1476 (N_1476,N_1431,N_1403);
or U1477 (N_1477,N_1442,N_1413);
nand U1478 (N_1478,N_1431,N_1444);
xor U1479 (N_1479,N_1433,N_1400);
nor U1480 (N_1480,N_1415,N_1431);
nor U1481 (N_1481,N_1406,N_1432);
nor U1482 (N_1482,N_1444,N_1425);
nand U1483 (N_1483,N_1406,N_1447);
or U1484 (N_1484,N_1417,N_1436);
or U1485 (N_1485,N_1420,N_1440);
nand U1486 (N_1486,N_1446,N_1431);
xnor U1487 (N_1487,N_1403,N_1408);
or U1488 (N_1488,N_1446,N_1436);
or U1489 (N_1489,N_1426,N_1401);
or U1490 (N_1490,N_1414,N_1416);
or U1491 (N_1491,N_1438,N_1449);
and U1492 (N_1492,N_1403,N_1438);
nor U1493 (N_1493,N_1429,N_1443);
nand U1494 (N_1494,N_1421,N_1416);
and U1495 (N_1495,N_1430,N_1442);
or U1496 (N_1496,N_1417,N_1443);
nand U1497 (N_1497,N_1409,N_1402);
nor U1498 (N_1498,N_1430,N_1416);
nand U1499 (N_1499,N_1440,N_1432);
or U1500 (N_1500,N_1457,N_1494);
and U1501 (N_1501,N_1497,N_1486);
nand U1502 (N_1502,N_1454,N_1481);
and U1503 (N_1503,N_1477,N_1480);
or U1504 (N_1504,N_1492,N_1484);
and U1505 (N_1505,N_1475,N_1471);
nand U1506 (N_1506,N_1487,N_1491);
and U1507 (N_1507,N_1455,N_1452);
or U1508 (N_1508,N_1482,N_1462);
and U1509 (N_1509,N_1451,N_1466);
and U1510 (N_1510,N_1461,N_1450);
or U1511 (N_1511,N_1460,N_1483);
nand U1512 (N_1512,N_1467,N_1468);
nand U1513 (N_1513,N_1453,N_1472);
nor U1514 (N_1514,N_1469,N_1465);
nor U1515 (N_1515,N_1485,N_1489);
and U1516 (N_1516,N_1490,N_1479);
nand U1517 (N_1517,N_1498,N_1476);
and U1518 (N_1518,N_1463,N_1499);
nand U1519 (N_1519,N_1464,N_1459);
nand U1520 (N_1520,N_1478,N_1474);
nor U1521 (N_1521,N_1496,N_1470);
nor U1522 (N_1522,N_1458,N_1456);
and U1523 (N_1523,N_1493,N_1495);
and U1524 (N_1524,N_1473,N_1488);
and U1525 (N_1525,N_1474,N_1461);
or U1526 (N_1526,N_1473,N_1467);
nand U1527 (N_1527,N_1476,N_1479);
nand U1528 (N_1528,N_1466,N_1472);
nor U1529 (N_1529,N_1464,N_1474);
nand U1530 (N_1530,N_1478,N_1464);
or U1531 (N_1531,N_1496,N_1450);
and U1532 (N_1532,N_1460,N_1478);
and U1533 (N_1533,N_1452,N_1467);
nand U1534 (N_1534,N_1483,N_1463);
nand U1535 (N_1535,N_1460,N_1493);
or U1536 (N_1536,N_1487,N_1479);
or U1537 (N_1537,N_1497,N_1453);
or U1538 (N_1538,N_1463,N_1465);
or U1539 (N_1539,N_1498,N_1495);
and U1540 (N_1540,N_1450,N_1485);
or U1541 (N_1541,N_1488,N_1466);
and U1542 (N_1542,N_1482,N_1468);
or U1543 (N_1543,N_1459,N_1450);
nor U1544 (N_1544,N_1453,N_1454);
and U1545 (N_1545,N_1490,N_1467);
nor U1546 (N_1546,N_1467,N_1474);
nor U1547 (N_1547,N_1490,N_1496);
and U1548 (N_1548,N_1459,N_1472);
and U1549 (N_1549,N_1481,N_1456);
and U1550 (N_1550,N_1547,N_1516);
or U1551 (N_1551,N_1512,N_1545);
or U1552 (N_1552,N_1532,N_1528);
and U1553 (N_1553,N_1524,N_1506);
or U1554 (N_1554,N_1505,N_1548);
or U1555 (N_1555,N_1507,N_1543);
and U1556 (N_1556,N_1536,N_1518);
xor U1557 (N_1557,N_1531,N_1525);
and U1558 (N_1558,N_1510,N_1541);
and U1559 (N_1559,N_1521,N_1515);
and U1560 (N_1560,N_1519,N_1514);
or U1561 (N_1561,N_1509,N_1535);
nor U1562 (N_1562,N_1530,N_1539);
nor U1563 (N_1563,N_1546,N_1529);
nor U1564 (N_1564,N_1533,N_1502);
or U1565 (N_1565,N_1513,N_1523);
and U1566 (N_1566,N_1527,N_1503);
nor U1567 (N_1567,N_1526,N_1508);
and U1568 (N_1568,N_1544,N_1538);
or U1569 (N_1569,N_1540,N_1542);
or U1570 (N_1570,N_1522,N_1517);
or U1571 (N_1571,N_1534,N_1501);
and U1572 (N_1572,N_1500,N_1549);
nor U1573 (N_1573,N_1511,N_1537);
and U1574 (N_1574,N_1520,N_1504);
or U1575 (N_1575,N_1520,N_1542);
and U1576 (N_1576,N_1510,N_1521);
xor U1577 (N_1577,N_1525,N_1548);
nor U1578 (N_1578,N_1517,N_1502);
nor U1579 (N_1579,N_1520,N_1522);
or U1580 (N_1580,N_1530,N_1538);
and U1581 (N_1581,N_1546,N_1528);
nor U1582 (N_1582,N_1521,N_1548);
nor U1583 (N_1583,N_1511,N_1528);
xor U1584 (N_1584,N_1517,N_1542);
nand U1585 (N_1585,N_1507,N_1538);
nand U1586 (N_1586,N_1535,N_1541);
nand U1587 (N_1587,N_1527,N_1538);
or U1588 (N_1588,N_1549,N_1524);
nor U1589 (N_1589,N_1546,N_1549);
nor U1590 (N_1590,N_1511,N_1533);
nand U1591 (N_1591,N_1528,N_1502);
nor U1592 (N_1592,N_1546,N_1544);
nand U1593 (N_1593,N_1520,N_1501);
or U1594 (N_1594,N_1540,N_1518);
nor U1595 (N_1595,N_1517,N_1540);
and U1596 (N_1596,N_1547,N_1528);
nor U1597 (N_1597,N_1502,N_1531);
or U1598 (N_1598,N_1513,N_1516);
or U1599 (N_1599,N_1516,N_1530);
nor U1600 (N_1600,N_1598,N_1591);
nand U1601 (N_1601,N_1577,N_1580);
nand U1602 (N_1602,N_1573,N_1585);
and U1603 (N_1603,N_1581,N_1578);
or U1604 (N_1604,N_1589,N_1595);
nor U1605 (N_1605,N_1567,N_1568);
nor U1606 (N_1606,N_1586,N_1592);
or U1607 (N_1607,N_1566,N_1559);
or U1608 (N_1608,N_1575,N_1570);
nor U1609 (N_1609,N_1555,N_1571);
or U1610 (N_1610,N_1561,N_1556);
and U1611 (N_1611,N_1554,N_1564);
nand U1612 (N_1612,N_1594,N_1569);
and U1613 (N_1613,N_1599,N_1552);
nand U1614 (N_1614,N_1579,N_1597);
or U1615 (N_1615,N_1584,N_1558);
and U1616 (N_1616,N_1565,N_1587);
nand U1617 (N_1617,N_1582,N_1563);
and U1618 (N_1618,N_1593,N_1576);
nand U1619 (N_1619,N_1550,N_1562);
and U1620 (N_1620,N_1590,N_1551);
or U1621 (N_1621,N_1583,N_1560);
nor U1622 (N_1622,N_1557,N_1588);
nand U1623 (N_1623,N_1574,N_1553);
or U1624 (N_1624,N_1572,N_1596);
and U1625 (N_1625,N_1585,N_1555);
and U1626 (N_1626,N_1574,N_1598);
nand U1627 (N_1627,N_1556,N_1555);
nand U1628 (N_1628,N_1570,N_1593);
and U1629 (N_1629,N_1590,N_1568);
nor U1630 (N_1630,N_1583,N_1561);
nand U1631 (N_1631,N_1584,N_1587);
nand U1632 (N_1632,N_1559,N_1560);
nor U1633 (N_1633,N_1587,N_1593);
nand U1634 (N_1634,N_1563,N_1559);
nand U1635 (N_1635,N_1569,N_1573);
nor U1636 (N_1636,N_1562,N_1580);
or U1637 (N_1637,N_1565,N_1588);
nor U1638 (N_1638,N_1595,N_1555);
and U1639 (N_1639,N_1559,N_1555);
nor U1640 (N_1640,N_1568,N_1574);
or U1641 (N_1641,N_1593,N_1582);
or U1642 (N_1642,N_1596,N_1570);
or U1643 (N_1643,N_1566,N_1591);
nand U1644 (N_1644,N_1596,N_1590);
nor U1645 (N_1645,N_1560,N_1565);
nand U1646 (N_1646,N_1566,N_1550);
nor U1647 (N_1647,N_1599,N_1562);
nor U1648 (N_1648,N_1551,N_1555);
or U1649 (N_1649,N_1589,N_1590);
nor U1650 (N_1650,N_1616,N_1641);
nand U1651 (N_1651,N_1615,N_1633);
or U1652 (N_1652,N_1643,N_1636);
nand U1653 (N_1653,N_1638,N_1604);
nor U1654 (N_1654,N_1648,N_1629);
or U1655 (N_1655,N_1649,N_1621);
nor U1656 (N_1656,N_1617,N_1607);
or U1657 (N_1657,N_1614,N_1646);
nand U1658 (N_1658,N_1602,N_1644);
and U1659 (N_1659,N_1642,N_1624);
nor U1660 (N_1660,N_1601,N_1645);
xor U1661 (N_1661,N_1647,N_1637);
nand U1662 (N_1662,N_1608,N_1623);
and U1663 (N_1663,N_1625,N_1627);
and U1664 (N_1664,N_1640,N_1613);
nand U1665 (N_1665,N_1618,N_1634);
and U1666 (N_1666,N_1610,N_1612);
nand U1667 (N_1667,N_1639,N_1630);
or U1668 (N_1668,N_1609,N_1605);
nor U1669 (N_1669,N_1626,N_1619);
or U1670 (N_1670,N_1600,N_1620);
nor U1671 (N_1671,N_1628,N_1622);
nor U1672 (N_1672,N_1632,N_1611);
nor U1673 (N_1673,N_1606,N_1631);
and U1674 (N_1674,N_1603,N_1635);
and U1675 (N_1675,N_1621,N_1639);
nor U1676 (N_1676,N_1638,N_1623);
nor U1677 (N_1677,N_1623,N_1626);
nor U1678 (N_1678,N_1632,N_1608);
or U1679 (N_1679,N_1646,N_1628);
and U1680 (N_1680,N_1627,N_1629);
nor U1681 (N_1681,N_1636,N_1615);
nor U1682 (N_1682,N_1624,N_1600);
nand U1683 (N_1683,N_1612,N_1611);
and U1684 (N_1684,N_1649,N_1604);
or U1685 (N_1685,N_1635,N_1637);
or U1686 (N_1686,N_1647,N_1622);
nand U1687 (N_1687,N_1619,N_1638);
or U1688 (N_1688,N_1648,N_1605);
nor U1689 (N_1689,N_1634,N_1613);
nand U1690 (N_1690,N_1648,N_1639);
nor U1691 (N_1691,N_1604,N_1617);
and U1692 (N_1692,N_1621,N_1635);
or U1693 (N_1693,N_1634,N_1642);
and U1694 (N_1694,N_1641,N_1608);
and U1695 (N_1695,N_1646,N_1648);
xnor U1696 (N_1696,N_1610,N_1633);
nor U1697 (N_1697,N_1618,N_1619);
nor U1698 (N_1698,N_1623,N_1624);
nor U1699 (N_1699,N_1606,N_1617);
or U1700 (N_1700,N_1653,N_1675);
nand U1701 (N_1701,N_1660,N_1654);
nand U1702 (N_1702,N_1682,N_1689);
nor U1703 (N_1703,N_1696,N_1657);
and U1704 (N_1704,N_1699,N_1673);
and U1705 (N_1705,N_1670,N_1693);
or U1706 (N_1706,N_1679,N_1656);
or U1707 (N_1707,N_1659,N_1694);
nand U1708 (N_1708,N_1672,N_1652);
and U1709 (N_1709,N_1684,N_1695);
or U1710 (N_1710,N_1683,N_1666);
nor U1711 (N_1711,N_1669,N_1698);
nor U1712 (N_1712,N_1692,N_1678);
nand U1713 (N_1713,N_1688,N_1665);
or U1714 (N_1714,N_1680,N_1671);
or U1715 (N_1715,N_1677,N_1651);
and U1716 (N_1716,N_1691,N_1681);
nor U1717 (N_1717,N_1662,N_1674);
and U1718 (N_1718,N_1690,N_1650);
and U1719 (N_1719,N_1687,N_1697);
nor U1720 (N_1720,N_1676,N_1661);
nor U1721 (N_1721,N_1668,N_1664);
nand U1722 (N_1722,N_1685,N_1663);
and U1723 (N_1723,N_1667,N_1655);
nor U1724 (N_1724,N_1658,N_1686);
nand U1725 (N_1725,N_1676,N_1685);
nor U1726 (N_1726,N_1675,N_1661);
nor U1727 (N_1727,N_1661,N_1682);
nand U1728 (N_1728,N_1696,N_1697);
or U1729 (N_1729,N_1685,N_1690);
nand U1730 (N_1730,N_1671,N_1666);
and U1731 (N_1731,N_1659,N_1652);
or U1732 (N_1732,N_1660,N_1651);
or U1733 (N_1733,N_1674,N_1657);
nor U1734 (N_1734,N_1697,N_1677);
nor U1735 (N_1735,N_1673,N_1657);
nor U1736 (N_1736,N_1667,N_1698);
nor U1737 (N_1737,N_1680,N_1696);
and U1738 (N_1738,N_1667,N_1664);
or U1739 (N_1739,N_1676,N_1678);
nand U1740 (N_1740,N_1674,N_1688);
nor U1741 (N_1741,N_1657,N_1660);
nand U1742 (N_1742,N_1668,N_1663);
xnor U1743 (N_1743,N_1692,N_1679);
or U1744 (N_1744,N_1657,N_1668);
or U1745 (N_1745,N_1679,N_1653);
nand U1746 (N_1746,N_1666,N_1693);
and U1747 (N_1747,N_1676,N_1696);
or U1748 (N_1748,N_1684,N_1679);
or U1749 (N_1749,N_1695,N_1654);
or U1750 (N_1750,N_1740,N_1726);
nor U1751 (N_1751,N_1705,N_1716);
nand U1752 (N_1752,N_1713,N_1701);
nand U1753 (N_1753,N_1719,N_1742);
or U1754 (N_1754,N_1729,N_1711);
nand U1755 (N_1755,N_1741,N_1732);
nand U1756 (N_1756,N_1706,N_1738);
and U1757 (N_1757,N_1700,N_1745);
nand U1758 (N_1758,N_1704,N_1724);
or U1759 (N_1759,N_1743,N_1747);
nand U1760 (N_1760,N_1735,N_1723);
nand U1761 (N_1761,N_1708,N_1712);
or U1762 (N_1762,N_1739,N_1718);
nand U1763 (N_1763,N_1736,N_1749);
xor U1764 (N_1764,N_1710,N_1707);
and U1765 (N_1765,N_1720,N_1727);
xnor U1766 (N_1766,N_1733,N_1715);
nor U1767 (N_1767,N_1734,N_1725);
nand U1768 (N_1768,N_1714,N_1709);
nor U1769 (N_1769,N_1746,N_1731);
or U1770 (N_1770,N_1722,N_1702);
nor U1771 (N_1771,N_1717,N_1737);
or U1772 (N_1772,N_1748,N_1744);
or U1773 (N_1773,N_1730,N_1728);
or U1774 (N_1774,N_1703,N_1721);
and U1775 (N_1775,N_1732,N_1724);
nand U1776 (N_1776,N_1702,N_1704);
nand U1777 (N_1777,N_1716,N_1701);
nor U1778 (N_1778,N_1701,N_1703);
or U1779 (N_1779,N_1748,N_1710);
nand U1780 (N_1780,N_1739,N_1720);
or U1781 (N_1781,N_1739,N_1713);
nand U1782 (N_1782,N_1720,N_1706);
nor U1783 (N_1783,N_1716,N_1724);
nand U1784 (N_1784,N_1741,N_1731);
nor U1785 (N_1785,N_1700,N_1735);
nor U1786 (N_1786,N_1718,N_1715);
or U1787 (N_1787,N_1708,N_1715);
and U1788 (N_1788,N_1722,N_1729);
nand U1789 (N_1789,N_1708,N_1705);
nand U1790 (N_1790,N_1718,N_1740);
nand U1791 (N_1791,N_1712,N_1748);
nand U1792 (N_1792,N_1746,N_1724);
or U1793 (N_1793,N_1737,N_1749);
nor U1794 (N_1794,N_1708,N_1727);
nor U1795 (N_1795,N_1709,N_1716);
or U1796 (N_1796,N_1745,N_1704);
and U1797 (N_1797,N_1740,N_1730);
or U1798 (N_1798,N_1714,N_1728);
and U1799 (N_1799,N_1711,N_1746);
and U1800 (N_1800,N_1789,N_1776);
or U1801 (N_1801,N_1758,N_1759);
and U1802 (N_1802,N_1753,N_1788);
and U1803 (N_1803,N_1792,N_1790);
and U1804 (N_1804,N_1779,N_1775);
nor U1805 (N_1805,N_1754,N_1791);
nor U1806 (N_1806,N_1798,N_1766);
and U1807 (N_1807,N_1787,N_1780);
nor U1808 (N_1808,N_1767,N_1794);
xnor U1809 (N_1809,N_1769,N_1771);
nand U1810 (N_1810,N_1762,N_1799);
or U1811 (N_1811,N_1781,N_1763);
or U1812 (N_1812,N_1797,N_1782);
or U1813 (N_1813,N_1783,N_1761);
nor U1814 (N_1814,N_1774,N_1778);
and U1815 (N_1815,N_1770,N_1768);
or U1816 (N_1816,N_1755,N_1760);
nor U1817 (N_1817,N_1777,N_1786);
nor U1818 (N_1818,N_1757,N_1750);
xnor U1819 (N_1819,N_1772,N_1756);
nor U1820 (N_1820,N_1784,N_1765);
nand U1821 (N_1821,N_1796,N_1764);
and U1822 (N_1822,N_1785,N_1793);
nand U1823 (N_1823,N_1752,N_1773);
and U1824 (N_1824,N_1795,N_1751);
or U1825 (N_1825,N_1752,N_1788);
nand U1826 (N_1826,N_1786,N_1751);
or U1827 (N_1827,N_1794,N_1797);
nor U1828 (N_1828,N_1764,N_1784);
nor U1829 (N_1829,N_1764,N_1797);
and U1830 (N_1830,N_1774,N_1784);
or U1831 (N_1831,N_1797,N_1754);
or U1832 (N_1832,N_1751,N_1780);
nand U1833 (N_1833,N_1769,N_1757);
nor U1834 (N_1834,N_1785,N_1757);
nand U1835 (N_1835,N_1756,N_1757);
or U1836 (N_1836,N_1751,N_1794);
or U1837 (N_1837,N_1791,N_1774);
nor U1838 (N_1838,N_1765,N_1799);
nand U1839 (N_1839,N_1787,N_1776);
or U1840 (N_1840,N_1765,N_1773);
nor U1841 (N_1841,N_1754,N_1794);
or U1842 (N_1842,N_1769,N_1758);
nand U1843 (N_1843,N_1752,N_1766);
and U1844 (N_1844,N_1779,N_1794);
nor U1845 (N_1845,N_1762,N_1754);
and U1846 (N_1846,N_1787,N_1758);
nand U1847 (N_1847,N_1790,N_1762);
or U1848 (N_1848,N_1790,N_1751);
or U1849 (N_1849,N_1769,N_1767);
nand U1850 (N_1850,N_1812,N_1810);
or U1851 (N_1851,N_1820,N_1841);
nor U1852 (N_1852,N_1803,N_1842);
or U1853 (N_1853,N_1832,N_1809);
nor U1854 (N_1854,N_1844,N_1801);
or U1855 (N_1855,N_1846,N_1823);
and U1856 (N_1856,N_1825,N_1814);
nand U1857 (N_1857,N_1802,N_1834);
nand U1858 (N_1858,N_1843,N_1811);
nor U1859 (N_1859,N_1817,N_1847);
xnor U1860 (N_1860,N_1815,N_1827);
nand U1861 (N_1861,N_1833,N_1849);
nor U1862 (N_1862,N_1807,N_1806);
and U1863 (N_1863,N_1845,N_1804);
nor U1864 (N_1864,N_1805,N_1829);
nor U1865 (N_1865,N_1837,N_1836);
nand U1866 (N_1866,N_1824,N_1813);
and U1867 (N_1867,N_1840,N_1821);
nand U1868 (N_1868,N_1831,N_1800);
or U1869 (N_1869,N_1822,N_1818);
nor U1870 (N_1870,N_1839,N_1830);
xnor U1871 (N_1871,N_1838,N_1835);
nor U1872 (N_1872,N_1819,N_1848);
xnor U1873 (N_1873,N_1828,N_1826);
nor U1874 (N_1874,N_1816,N_1808);
and U1875 (N_1875,N_1810,N_1807);
and U1876 (N_1876,N_1808,N_1804);
nand U1877 (N_1877,N_1838,N_1833);
and U1878 (N_1878,N_1819,N_1833);
and U1879 (N_1879,N_1824,N_1814);
nand U1880 (N_1880,N_1811,N_1814);
xor U1881 (N_1881,N_1845,N_1837);
or U1882 (N_1882,N_1832,N_1819);
nor U1883 (N_1883,N_1805,N_1831);
and U1884 (N_1884,N_1849,N_1811);
and U1885 (N_1885,N_1835,N_1802);
nand U1886 (N_1886,N_1820,N_1828);
nand U1887 (N_1887,N_1809,N_1846);
nand U1888 (N_1888,N_1841,N_1801);
and U1889 (N_1889,N_1815,N_1814);
nand U1890 (N_1890,N_1831,N_1819);
nand U1891 (N_1891,N_1828,N_1804);
and U1892 (N_1892,N_1823,N_1848);
and U1893 (N_1893,N_1810,N_1827);
or U1894 (N_1894,N_1845,N_1807);
or U1895 (N_1895,N_1802,N_1801);
or U1896 (N_1896,N_1840,N_1804);
and U1897 (N_1897,N_1843,N_1828);
nor U1898 (N_1898,N_1809,N_1801);
nor U1899 (N_1899,N_1820,N_1840);
nor U1900 (N_1900,N_1859,N_1858);
nand U1901 (N_1901,N_1882,N_1868);
and U1902 (N_1902,N_1897,N_1872);
or U1903 (N_1903,N_1891,N_1857);
and U1904 (N_1904,N_1880,N_1869);
and U1905 (N_1905,N_1894,N_1896);
or U1906 (N_1906,N_1884,N_1899);
nor U1907 (N_1907,N_1850,N_1863);
or U1908 (N_1908,N_1893,N_1898);
and U1909 (N_1909,N_1879,N_1881);
nor U1910 (N_1910,N_1889,N_1854);
and U1911 (N_1911,N_1886,N_1873);
or U1912 (N_1912,N_1865,N_1852);
nor U1913 (N_1913,N_1877,N_1856);
or U1914 (N_1914,N_1892,N_1860);
and U1915 (N_1915,N_1895,N_1861);
nand U1916 (N_1916,N_1862,N_1851);
and U1917 (N_1917,N_1878,N_1867);
nor U1918 (N_1918,N_1864,N_1887);
nand U1919 (N_1919,N_1874,N_1875);
or U1920 (N_1920,N_1855,N_1888);
nand U1921 (N_1921,N_1883,N_1853);
nor U1922 (N_1922,N_1870,N_1890);
and U1923 (N_1923,N_1885,N_1871);
or U1924 (N_1924,N_1866,N_1876);
or U1925 (N_1925,N_1876,N_1882);
nand U1926 (N_1926,N_1862,N_1870);
or U1927 (N_1927,N_1850,N_1884);
nor U1928 (N_1928,N_1858,N_1856);
nor U1929 (N_1929,N_1873,N_1864);
or U1930 (N_1930,N_1889,N_1876);
and U1931 (N_1931,N_1893,N_1867);
or U1932 (N_1932,N_1859,N_1872);
and U1933 (N_1933,N_1877,N_1887);
nand U1934 (N_1934,N_1856,N_1861);
and U1935 (N_1935,N_1885,N_1881);
and U1936 (N_1936,N_1863,N_1860);
or U1937 (N_1937,N_1863,N_1859);
and U1938 (N_1938,N_1868,N_1871);
or U1939 (N_1939,N_1861,N_1874);
nand U1940 (N_1940,N_1898,N_1867);
nor U1941 (N_1941,N_1870,N_1860);
nor U1942 (N_1942,N_1853,N_1876);
and U1943 (N_1943,N_1879,N_1865);
and U1944 (N_1944,N_1895,N_1857);
or U1945 (N_1945,N_1882,N_1871);
nor U1946 (N_1946,N_1885,N_1890);
nand U1947 (N_1947,N_1862,N_1876);
nor U1948 (N_1948,N_1860,N_1887);
or U1949 (N_1949,N_1850,N_1886);
and U1950 (N_1950,N_1928,N_1910);
nor U1951 (N_1951,N_1922,N_1906);
nor U1952 (N_1952,N_1902,N_1916);
nand U1953 (N_1953,N_1942,N_1925);
nand U1954 (N_1954,N_1903,N_1921);
nor U1955 (N_1955,N_1900,N_1914);
nor U1956 (N_1956,N_1941,N_1927);
nor U1957 (N_1957,N_1944,N_1913);
nor U1958 (N_1958,N_1934,N_1949);
nor U1959 (N_1959,N_1948,N_1947);
nand U1960 (N_1960,N_1918,N_1932);
nor U1961 (N_1961,N_1936,N_1915);
nand U1962 (N_1962,N_1905,N_1939);
nand U1963 (N_1963,N_1937,N_1907);
or U1964 (N_1964,N_1909,N_1908);
or U1965 (N_1965,N_1911,N_1912);
nor U1966 (N_1966,N_1933,N_1930);
xor U1967 (N_1967,N_1920,N_1940);
nand U1968 (N_1968,N_1935,N_1901);
and U1969 (N_1969,N_1943,N_1938);
and U1970 (N_1970,N_1919,N_1931);
nand U1971 (N_1971,N_1926,N_1924);
nand U1972 (N_1972,N_1945,N_1946);
and U1973 (N_1973,N_1904,N_1917);
and U1974 (N_1974,N_1929,N_1923);
nand U1975 (N_1975,N_1930,N_1942);
nor U1976 (N_1976,N_1911,N_1930);
or U1977 (N_1977,N_1949,N_1942);
nor U1978 (N_1978,N_1935,N_1934);
nand U1979 (N_1979,N_1922,N_1915);
nand U1980 (N_1980,N_1946,N_1924);
and U1981 (N_1981,N_1914,N_1910);
or U1982 (N_1982,N_1909,N_1934);
nand U1983 (N_1983,N_1924,N_1927);
or U1984 (N_1984,N_1927,N_1913);
nor U1985 (N_1985,N_1934,N_1916);
xor U1986 (N_1986,N_1943,N_1909);
nor U1987 (N_1987,N_1928,N_1943);
nor U1988 (N_1988,N_1942,N_1923);
and U1989 (N_1989,N_1912,N_1943);
or U1990 (N_1990,N_1922,N_1917);
nor U1991 (N_1991,N_1947,N_1911);
nor U1992 (N_1992,N_1910,N_1936);
or U1993 (N_1993,N_1915,N_1931);
nor U1994 (N_1994,N_1941,N_1939);
nor U1995 (N_1995,N_1914,N_1923);
nor U1996 (N_1996,N_1907,N_1913);
or U1997 (N_1997,N_1924,N_1903);
or U1998 (N_1998,N_1924,N_1943);
and U1999 (N_1999,N_1910,N_1940);
nor U2000 (N_2000,N_1979,N_1993);
and U2001 (N_2001,N_1962,N_1995);
and U2002 (N_2002,N_1994,N_1951);
or U2003 (N_2003,N_1973,N_1977);
or U2004 (N_2004,N_1985,N_1961);
nor U2005 (N_2005,N_1983,N_1958);
or U2006 (N_2006,N_1967,N_1960);
and U2007 (N_2007,N_1998,N_1971);
or U2008 (N_2008,N_1956,N_1999);
and U2009 (N_2009,N_1978,N_1975);
or U2010 (N_2010,N_1984,N_1991);
and U2011 (N_2011,N_1981,N_1954);
nand U2012 (N_2012,N_1996,N_1986);
nor U2013 (N_2013,N_1966,N_1990);
xnor U2014 (N_2014,N_1988,N_1980);
nor U2015 (N_2015,N_1989,N_1987);
or U2016 (N_2016,N_1997,N_1992);
nor U2017 (N_2017,N_1970,N_1953);
nor U2018 (N_2018,N_1952,N_1974);
or U2019 (N_2019,N_1964,N_1976);
nor U2020 (N_2020,N_1982,N_1950);
or U2021 (N_2021,N_1957,N_1972);
or U2022 (N_2022,N_1969,N_1959);
and U2023 (N_2023,N_1965,N_1955);
and U2024 (N_2024,N_1968,N_1963);
and U2025 (N_2025,N_1969,N_1951);
nor U2026 (N_2026,N_1982,N_1958);
or U2027 (N_2027,N_1974,N_1982);
nand U2028 (N_2028,N_1963,N_1967);
or U2029 (N_2029,N_1985,N_1975);
nor U2030 (N_2030,N_1989,N_1982);
or U2031 (N_2031,N_1968,N_1964);
and U2032 (N_2032,N_1977,N_1992);
nand U2033 (N_2033,N_1975,N_1972);
nand U2034 (N_2034,N_1996,N_1995);
nand U2035 (N_2035,N_1991,N_1970);
nand U2036 (N_2036,N_1974,N_1955);
nand U2037 (N_2037,N_1960,N_1961);
or U2038 (N_2038,N_1976,N_1967);
or U2039 (N_2039,N_1956,N_1992);
nor U2040 (N_2040,N_1998,N_1950);
and U2041 (N_2041,N_1988,N_1996);
nor U2042 (N_2042,N_1987,N_1972);
and U2043 (N_2043,N_1989,N_1988);
nor U2044 (N_2044,N_1985,N_1991);
and U2045 (N_2045,N_1952,N_1999);
nand U2046 (N_2046,N_1961,N_1996);
nor U2047 (N_2047,N_1991,N_1963);
nand U2048 (N_2048,N_1977,N_1970);
and U2049 (N_2049,N_1981,N_1957);
and U2050 (N_2050,N_2023,N_2027);
and U2051 (N_2051,N_2006,N_2031);
or U2052 (N_2052,N_2022,N_2025);
or U2053 (N_2053,N_2024,N_2020);
nor U2054 (N_2054,N_2000,N_2029);
nand U2055 (N_2055,N_2017,N_2011);
and U2056 (N_2056,N_2002,N_2041);
nor U2057 (N_2057,N_2015,N_2033);
nand U2058 (N_2058,N_2018,N_2039);
nor U2059 (N_2059,N_2046,N_2036);
nand U2060 (N_2060,N_2005,N_2004);
and U2061 (N_2061,N_2007,N_2047);
nor U2062 (N_2062,N_2010,N_2012);
or U2063 (N_2063,N_2001,N_2016);
or U2064 (N_2064,N_2035,N_2037);
nor U2065 (N_2065,N_2030,N_2049);
xor U2066 (N_2066,N_2008,N_2014);
or U2067 (N_2067,N_2026,N_2040);
nand U2068 (N_2068,N_2043,N_2009);
nor U2069 (N_2069,N_2034,N_2042);
nand U2070 (N_2070,N_2003,N_2038);
nor U2071 (N_2071,N_2028,N_2019);
nor U2072 (N_2072,N_2044,N_2048);
nand U2073 (N_2073,N_2045,N_2013);
nor U2074 (N_2074,N_2021,N_2032);
and U2075 (N_2075,N_2049,N_2021);
nand U2076 (N_2076,N_2047,N_2017);
nand U2077 (N_2077,N_2029,N_2006);
and U2078 (N_2078,N_2046,N_2003);
and U2079 (N_2079,N_2046,N_2011);
and U2080 (N_2080,N_2000,N_2011);
nor U2081 (N_2081,N_2042,N_2025);
and U2082 (N_2082,N_2005,N_2026);
or U2083 (N_2083,N_2044,N_2022);
nor U2084 (N_2084,N_2017,N_2019);
nor U2085 (N_2085,N_2025,N_2040);
nor U2086 (N_2086,N_2045,N_2039);
nand U2087 (N_2087,N_2047,N_2018);
nor U2088 (N_2088,N_2033,N_2034);
and U2089 (N_2089,N_2040,N_2020);
nand U2090 (N_2090,N_2016,N_2024);
xor U2091 (N_2091,N_2009,N_2035);
nand U2092 (N_2092,N_2041,N_2022);
nand U2093 (N_2093,N_2010,N_2023);
nand U2094 (N_2094,N_2015,N_2039);
nor U2095 (N_2095,N_2003,N_2039);
nand U2096 (N_2096,N_2048,N_2020);
and U2097 (N_2097,N_2027,N_2031);
or U2098 (N_2098,N_2023,N_2030);
or U2099 (N_2099,N_2004,N_2013);
nand U2100 (N_2100,N_2082,N_2060);
and U2101 (N_2101,N_2086,N_2097);
or U2102 (N_2102,N_2084,N_2091);
nor U2103 (N_2103,N_2070,N_2052);
nor U2104 (N_2104,N_2088,N_2096);
and U2105 (N_2105,N_2063,N_2056);
nor U2106 (N_2106,N_2094,N_2077);
or U2107 (N_2107,N_2081,N_2064);
xnor U2108 (N_2108,N_2074,N_2062);
nor U2109 (N_2109,N_2069,N_2098);
nor U2110 (N_2110,N_2080,N_2078);
nand U2111 (N_2111,N_2076,N_2054);
or U2112 (N_2112,N_2090,N_2089);
nor U2113 (N_2113,N_2057,N_2087);
nand U2114 (N_2114,N_2061,N_2051);
nand U2115 (N_2115,N_2053,N_2083);
nand U2116 (N_2116,N_2055,N_2067);
and U2117 (N_2117,N_2092,N_2073);
and U2118 (N_2118,N_2093,N_2085);
nand U2119 (N_2119,N_2059,N_2058);
nand U2120 (N_2120,N_2066,N_2072);
nor U2121 (N_2121,N_2099,N_2068);
nand U2122 (N_2122,N_2050,N_2075);
nand U2123 (N_2123,N_2095,N_2079);
and U2124 (N_2124,N_2065,N_2071);
nor U2125 (N_2125,N_2068,N_2051);
nor U2126 (N_2126,N_2052,N_2064);
and U2127 (N_2127,N_2053,N_2051);
or U2128 (N_2128,N_2098,N_2077);
and U2129 (N_2129,N_2081,N_2080);
xnor U2130 (N_2130,N_2072,N_2085);
nor U2131 (N_2131,N_2076,N_2096);
nand U2132 (N_2132,N_2080,N_2057);
nor U2133 (N_2133,N_2050,N_2070);
nand U2134 (N_2134,N_2057,N_2093);
and U2135 (N_2135,N_2060,N_2073);
and U2136 (N_2136,N_2081,N_2050);
nor U2137 (N_2137,N_2091,N_2058);
and U2138 (N_2138,N_2073,N_2058);
or U2139 (N_2139,N_2095,N_2073);
nor U2140 (N_2140,N_2063,N_2087);
xnor U2141 (N_2141,N_2077,N_2087);
nor U2142 (N_2142,N_2063,N_2057);
nand U2143 (N_2143,N_2054,N_2063);
nor U2144 (N_2144,N_2052,N_2090);
nor U2145 (N_2145,N_2083,N_2067);
nor U2146 (N_2146,N_2076,N_2087);
nand U2147 (N_2147,N_2067,N_2077);
nor U2148 (N_2148,N_2088,N_2069);
nor U2149 (N_2149,N_2087,N_2079);
and U2150 (N_2150,N_2105,N_2112);
nor U2151 (N_2151,N_2142,N_2130);
nand U2152 (N_2152,N_2111,N_2121);
nor U2153 (N_2153,N_2116,N_2141);
or U2154 (N_2154,N_2110,N_2124);
and U2155 (N_2155,N_2138,N_2127);
nand U2156 (N_2156,N_2148,N_2134);
or U2157 (N_2157,N_2132,N_2108);
and U2158 (N_2158,N_2146,N_2139);
nand U2159 (N_2159,N_2109,N_2115);
and U2160 (N_2160,N_2104,N_2145);
nor U2161 (N_2161,N_2140,N_2144);
and U2162 (N_2162,N_2113,N_2137);
or U2163 (N_2163,N_2103,N_2136);
and U2164 (N_2164,N_2102,N_2107);
nand U2165 (N_2165,N_2119,N_2147);
or U2166 (N_2166,N_2149,N_2120);
or U2167 (N_2167,N_2123,N_2131);
and U2168 (N_2168,N_2143,N_2118);
or U2169 (N_2169,N_2129,N_2128);
nand U2170 (N_2170,N_2135,N_2114);
nand U2171 (N_2171,N_2117,N_2122);
xnor U2172 (N_2172,N_2126,N_2100);
nand U2173 (N_2173,N_2133,N_2101);
nand U2174 (N_2174,N_2125,N_2106);
or U2175 (N_2175,N_2132,N_2129);
nand U2176 (N_2176,N_2143,N_2105);
nor U2177 (N_2177,N_2146,N_2104);
and U2178 (N_2178,N_2118,N_2122);
or U2179 (N_2179,N_2111,N_2108);
or U2180 (N_2180,N_2142,N_2118);
nor U2181 (N_2181,N_2113,N_2145);
nor U2182 (N_2182,N_2134,N_2144);
xor U2183 (N_2183,N_2119,N_2141);
and U2184 (N_2184,N_2147,N_2103);
and U2185 (N_2185,N_2144,N_2115);
nand U2186 (N_2186,N_2148,N_2124);
or U2187 (N_2187,N_2133,N_2119);
nand U2188 (N_2188,N_2148,N_2100);
nor U2189 (N_2189,N_2108,N_2138);
nand U2190 (N_2190,N_2112,N_2111);
nor U2191 (N_2191,N_2149,N_2130);
or U2192 (N_2192,N_2105,N_2145);
nand U2193 (N_2193,N_2103,N_2107);
nor U2194 (N_2194,N_2118,N_2147);
and U2195 (N_2195,N_2130,N_2145);
and U2196 (N_2196,N_2117,N_2138);
or U2197 (N_2197,N_2106,N_2123);
nor U2198 (N_2198,N_2106,N_2133);
or U2199 (N_2199,N_2128,N_2124);
nor U2200 (N_2200,N_2183,N_2166);
nor U2201 (N_2201,N_2185,N_2186);
and U2202 (N_2202,N_2150,N_2176);
and U2203 (N_2203,N_2198,N_2153);
or U2204 (N_2204,N_2194,N_2163);
nand U2205 (N_2205,N_2193,N_2167);
nor U2206 (N_2206,N_2172,N_2179);
and U2207 (N_2207,N_2152,N_2154);
nand U2208 (N_2208,N_2171,N_2191);
or U2209 (N_2209,N_2168,N_2187);
and U2210 (N_2210,N_2192,N_2164);
or U2211 (N_2211,N_2190,N_2151);
and U2212 (N_2212,N_2157,N_2197);
or U2213 (N_2213,N_2159,N_2165);
nor U2214 (N_2214,N_2196,N_2174);
or U2215 (N_2215,N_2177,N_2158);
or U2216 (N_2216,N_2170,N_2195);
nand U2217 (N_2217,N_2181,N_2189);
nor U2218 (N_2218,N_2173,N_2160);
nor U2219 (N_2219,N_2188,N_2155);
nor U2220 (N_2220,N_2162,N_2199);
nor U2221 (N_2221,N_2169,N_2161);
and U2222 (N_2222,N_2184,N_2175);
nand U2223 (N_2223,N_2178,N_2182);
or U2224 (N_2224,N_2180,N_2156);
nor U2225 (N_2225,N_2189,N_2164);
nand U2226 (N_2226,N_2173,N_2155);
nand U2227 (N_2227,N_2166,N_2153);
nor U2228 (N_2228,N_2184,N_2160);
nor U2229 (N_2229,N_2192,N_2195);
or U2230 (N_2230,N_2189,N_2187);
and U2231 (N_2231,N_2160,N_2182);
nor U2232 (N_2232,N_2182,N_2157);
or U2233 (N_2233,N_2195,N_2162);
and U2234 (N_2234,N_2194,N_2174);
and U2235 (N_2235,N_2182,N_2170);
nor U2236 (N_2236,N_2156,N_2191);
nand U2237 (N_2237,N_2150,N_2185);
or U2238 (N_2238,N_2169,N_2196);
nand U2239 (N_2239,N_2156,N_2194);
xor U2240 (N_2240,N_2189,N_2155);
nor U2241 (N_2241,N_2179,N_2153);
or U2242 (N_2242,N_2174,N_2166);
xor U2243 (N_2243,N_2196,N_2175);
and U2244 (N_2244,N_2161,N_2181);
nand U2245 (N_2245,N_2173,N_2194);
or U2246 (N_2246,N_2154,N_2189);
nand U2247 (N_2247,N_2151,N_2186);
or U2248 (N_2248,N_2190,N_2157);
nor U2249 (N_2249,N_2182,N_2198);
or U2250 (N_2250,N_2245,N_2220);
or U2251 (N_2251,N_2225,N_2215);
and U2252 (N_2252,N_2223,N_2201);
nor U2253 (N_2253,N_2229,N_2210);
or U2254 (N_2254,N_2238,N_2216);
and U2255 (N_2255,N_2202,N_2228);
or U2256 (N_2256,N_2241,N_2240);
and U2257 (N_2257,N_2247,N_2218);
or U2258 (N_2258,N_2248,N_2224);
nand U2259 (N_2259,N_2222,N_2243);
and U2260 (N_2260,N_2207,N_2213);
nand U2261 (N_2261,N_2242,N_2200);
nand U2262 (N_2262,N_2214,N_2211);
or U2263 (N_2263,N_2219,N_2217);
nand U2264 (N_2264,N_2235,N_2203);
nor U2265 (N_2265,N_2239,N_2221);
xnor U2266 (N_2266,N_2246,N_2244);
nand U2267 (N_2267,N_2249,N_2230);
or U2268 (N_2268,N_2212,N_2205);
nor U2269 (N_2269,N_2226,N_2231);
or U2270 (N_2270,N_2227,N_2236);
and U2271 (N_2271,N_2233,N_2208);
and U2272 (N_2272,N_2237,N_2209);
or U2273 (N_2273,N_2204,N_2232);
and U2274 (N_2274,N_2234,N_2206);
or U2275 (N_2275,N_2246,N_2214);
or U2276 (N_2276,N_2230,N_2226);
or U2277 (N_2277,N_2206,N_2239);
or U2278 (N_2278,N_2239,N_2246);
or U2279 (N_2279,N_2202,N_2238);
or U2280 (N_2280,N_2246,N_2202);
and U2281 (N_2281,N_2210,N_2228);
nand U2282 (N_2282,N_2228,N_2222);
and U2283 (N_2283,N_2241,N_2200);
nor U2284 (N_2284,N_2244,N_2207);
and U2285 (N_2285,N_2245,N_2204);
and U2286 (N_2286,N_2238,N_2242);
and U2287 (N_2287,N_2240,N_2229);
or U2288 (N_2288,N_2225,N_2245);
nor U2289 (N_2289,N_2216,N_2235);
nand U2290 (N_2290,N_2224,N_2227);
nand U2291 (N_2291,N_2242,N_2203);
or U2292 (N_2292,N_2207,N_2246);
nand U2293 (N_2293,N_2249,N_2245);
nand U2294 (N_2294,N_2216,N_2228);
nor U2295 (N_2295,N_2218,N_2205);
and U2296 (N_2296,N_2202,N_2233);
nor U2297 (N_2297,N_2224,N_2238);
nand U2298 (N_2298,N_2244,N_2221);
nor U2299 (N_2299,N_2226,N_2232);
nor U2300 (N_2300,N_2292,N_2294);
and U2301 (N_2301,N_2271,N_2293);
and U2302 (N_2302,N_2266,N_2262);
and U2303 (N_2303,N_2283,N_2291);
and U2304 (N_2304,N_2250,N_2259);
nor U2305 (N_2305,N_2268,N_2277);
and U2306 (N_2306,N_2255,N_2265);
and U2307 (N_2307,N_2269,N_2288);
and U2308 (N_2308,N_2257,N_2263);
or U2309 (N_2309,N_2289,N_2290);
nor U2310 (N_2310,N_2273,N_2285);
and U2311 (N_2311,N_2296,N_2260);
nand U2312 (N_2312,N_2272,N_2267);
or U2313 (N_2313,N_2274,N_2284);
nor U2314 (N_2314,N_2281,N_2278);
nor U2315 (N_2315,N_2264,N_2270);
or U2316 (N_2316,N_2252,N_2275);
nor U2317 (N_2317,N_2251,N_2298);
or U2318 (N_2318,N_2299,N_2254);
and U2319 (N_2319,N_2295,N_2253);
and U2320 (N_2320,N_2258,N_2276);
nor U2321 (N_2321,N_2297,N_2286);
nor U2322 (N_2322,N_2287,N_2279);
nor U2323 (N_2323,N_2256,N_2282);
nand U2324 (N_2324,N_2280,N_2261);
nor U2325 (N_2325,N_2289,N_2288);
nand U2326 (N_2326,N_2275,N_2265);
nand U2327 (N_2327,N_2269,N_2275);
nor U2328 (N_2328,N_2280,N_2291);
and U2329 (N_2329,N_2282,N_2279);
nor U2330 (N_2330,N_2277,N_2280);
and U2331 (N_2331,N_2266,N_2259);
nand U2332 (N_2332,N_2298,N_2267);
nand U2333 (N_2333,N_2282,N_2276);
nand U2334 (N_2334,N_2256,N_2270);
nand U2335 (N_2335,N_2278,N_2250);
or U2336 (N_2336,N_2282,N_2278);
nand U2337 (N_2337,N_2256,N_2290);
nor U2338 (N_2338,N_2294,N_2276);
and U2339 (N_2339,N_2255,N_2266);
and U2340 (N_2340,N_2261,N_2260);
or U2341 (N_2341,N_2250,N_2280);
nand U2342 (N_2342,N_2261,N_2270);
nand U2343 (N_2343,N_2285,N_2274);
nor U2344 (N_2344,N_2256,N_2291);
nor U2345 (N_2345,N_2263,N_2296);
nor U2346 (N_2346,N_2259,N_2265);
nor U2347 (N_2347,N_2257,N_2264);
or U2348 (N_2348,N_2285,N_2295);
or U2349 (N_2349,N_2283,N_2265);
or U2350 (N_2350,N_2316,N_2342);
nor U2351 (N_2351,N_2338,N_2326);
nor U2352 (N_2352,N_2334,N_2308);
or U2353 (N_2353,N_2325,N_2301);
and U2354 (N_2354,N_2322,N_2335);
nor U2355 (N_2355,N_2315,N_2328);
and U2356 (N_2356,N_2339,N_2349);
or U2357 (N_2357,N_2337,N_2303);
and U2358 (N_2358,N_2317,N_2311);
nand U2359 (N_2359,N_2304,N_2302);
and U2360 (N_2360,N_2320,N_2347);
and U2361 (N_2361,N_2323,N_2324);
or U2362 (N_2362,N_2345,N_2331);
or U2363 (N_2363,N_2321,N_2300);
nand U2364 (N_2364,N_2343,N_2313);
or U2365 (N_2365,N_2329,N_2341);
and U2366 (N_2366,N_2314,N_2318);
and U2367 (N_2367,N_2309,N_2327);
xor U2368 (N_2368,N_2332,N_2340);
and U2369 (N_2369,N_2333,N_2306);
or U2370 (N_2370,N_2305,N_2310);
or U2371 (N_2371,N_2346,N_2344);
nor U2372 (N_2372,N_2330,N_2312);
nor U2373 (N_2373,N_2336,N_2307);
and U2374 (N_2374,N_2348,N_2319);
and U2375 (N_2375,N_2332,N_2349);
and U2376 (N_2376,N_2331,N_2336);
nor U2377 (N_2377,N_2325,N_2341);
nor U2378 (N_2378,N_2343,N_2305);
or U2379 (N_2379,N_2300,N_2326);
nor U2380 (N_2380,N_2336,N_2330);
and U2381 (N_2381,N_2336,N_2338);
nand U2382 (N_2382,N_2335,N_2309);
or U2383 (N_2383,N_2320,N_2300);
nand U2384 (N_2384,N_2301,N_2332);
nor U2385 (N_2385,N_2323,N_2345);
or U2386 (N_2386,N_2333,N_2343);
and U2387 (N_2387,N_2340,N_2336);
nand U2388 (N_2388,N_2345,N_2343);
nand U2389 (N_2389,N_2338,N_2329);
or U2390 (N_2390,N_2344,N_2308);
nand U2391 (N_2391,N_2320,N_2305);
or U2392 (N_2392,N_2306,N_2345);
xor U2393 (N_2393,N_2328,N_2347);
nand U2394 (N_2394,N_2313,N_2318);
nor U2395 (N_2395,N_2315,N_2311);
nor U2396 (N_2396,N_2321,N_2335);
nor U2397 (N_2397,N_2348,N_2332);
and U2398 (N_2398,N_2317,N_2316);
or U2399 (N_2399,N_2342,N_2301);
and U2400 (N_2400,N_2391,N_2385);
or U2401 (N_2401,N_2350,N_2370);
and U2402 (N_2402,N_2359,N_2354);
and U2403 (N_2403,N_2363,N_2360);
or U2404 (N_2404,N_2390,N_2361);
nor U2405 (N_2405,N_2395,N_2386);
and U2406 (N_2406,N_2366,N_2353);
and U2407 (N_2407,N_2355,N_2392);
or U2408 (N_2408,N_2373,N_2371);
or U2409 (N_2409,N_2357,N_2399);
or U2410 (N_2410,N_2376,N_2394);
or U2411 (N_2411,N_2398,N_2362);
nand U2412 (N_2412,N_2356,N_2382);
and U2413 (N_2413,N_2389,N_2374);
and U2414 (N_2414,N_2358,N_2397);
and U2415 (N_2415,N_2372,N_2377);
nor U2416 (N_2416,N_2383,N_2368);
nand U2417 (N_2417,N_2378,N_2367);
or U2418 (N_2418,N_2384,N_2369);
or U2419 (N_2419,N_2352,N_2387);
nor U2420 (N_2420,N_2379,N_2364);
and U2421 (N_2421,N_2351,N_2375);
and U2422 (N_2422,N_2380,N_2393);
nor U2423 (N_2423,N_2365,N_2388);
nor U2424 (N_2424,N_2381,N_2396);
nand U2425 (N_2425,N_2371,N_2350);
and U2426 (N_2426,N_2354,N_2367);
and U2427 (N_2427,N_2366,N_2383);
nand U2428 (N_2428,N_2396,N_2362);
and U2429 (N_2429,N_2369,N_2390);
or U2430 (N_2430,N_2376,N_2399);
and U2431 (N_2431,N_2357,N_2392);
nand U2432 (N_2432,N_2372,N_2351);
or U2433 (N_2433,N_2394,N_2396);
nand U2434 (N_2434,N_2354,N_2387);
nand U2435 (N_2435,N_2360,N_2359);
xnor U2436 (N_2436,N_2379,N_2381);
or U2437 (N_2437,N_2366,N_2364);
or U2438 (N_2438,N_2350,N_2390);
nand U2439 (N_2439,N_2382,N_2376);
and U2440 (N_2440,N_2366,N_2382);
nor U2441 (N_2441,N_2387,N_2394);
and U2442 (N_2442,N_2380,N_2370);
or U2443 (N_2443,N_2398,N_2357);
nor U2444 (N_2444,N_2360,N_2357);
and U2445 (N_2445,N_2350,N_2382);
nand U2446 (N_2446,N_2350,N_2377);
or U2447 (N_2447,N_2397,N_2394);
nor U2448 (N_2448,N_2395,N_2382);
nand U2449 (N_2449,N_2351,N_2367);
and U2450 (N_2450,N_2438,N_2436);
nor U2451 (N_2451,N_2406,N_2403);
xnor U2452 (N_2452,N_2411,N_2442);
nor U2453 (N_2453,N_2448,N_2429);
and U2454 (N_2454,N_2419,N_2412);
or U2455 (N_2455,N_2430,N_2423);
nand U2456 (N_2456,N_2418,N_2422);
or U2457 (N_2457,N_2428,N_2431);
nand U2458 (N_2458,N_2420,N_2408);
and U2459 (N_2459,N_2425,N_2437);
nor U2460 (N_2460,N_2427,N_2435);
nand U2461 (N_2461,N_2416,N_2413);
nand U2462 (N_2462,N_2444,N_2401);
nand U2463 (N_2463,N_2414,N_2421);
and U2464 (N_2464,N_2434,N_2415);
or U2465 (N_2465,N_2417,N_2432);
and U2466 (N_2466,N_2400,N_2405);
and U2467 (N_2467,N_2407,N_2426);
and U2468 (N_2468,N_2443,N_2424);
or U2469 (N_2469,N_2402,N_2404);
nand U2470 (N_2470,N_2445,N_2446);
and U2471 (N_2471,N_2433,N_2440);
nor U2472 (N_2472,N_2410,N_2441);
nand U2473 (N_2473,N_2449,N_2439);
nand U2474 (N_2474,N_2447,N_2409);
xnor U2475 (N_2475,N_2415,N_2401);
nand U2476 (N_2476,N_2417,N_2410);
or U2477 (N_2477,N_2407,N_2436);
nand U2478 (N_2478,N_2422,N_2437);
nor U2479 (N_2479,N_2446,N_2416);
nor U2480 (N_2480,N_2408,N_2406);
nor U2481 (N_2481,N_2441,N_2401);
nand U2482 (N_2482,N_2407,N_2401);
nor U2483 (N_2483,N_2412,N_2406);
nor U2484 (N_2484,N_2422,N_2412);
or U2485 (N_2485,N_2449,N_2411);
nand U2486 (N_2486,N_2410,N_2404);
nor U2487 (N_2487,N_2448,N_2423);
nand U2488 (N_2488,N_2431,N_2440);
nand U2489 (N_2489,N_2409,N_2421);
and U2490 (N_2490,N_2432,N_2439);
nor U2491 (N_2491,N_2410,N_2408);
and U2492 (N_2492,N_2426,N_2403);
or U2493 (N_2493,N_2400,N_2433);
nand U2494 (N_2494,N_2437,N_2448);
or U2495 (N_2495,N_2438,N_2415);
nand U2496 (N_2496,N_2408,N_2440);
nand U2497 (N_2497,N_2419,N_2409);
or U2498 (N_2498,N_2411,N_2402);
or U2499 (N_2499,N_2449,N_2408);
or U2500 (N_2500,N_2498,N_2454);
nor U2501 (N_2501,N_2486,N_2451);
nand U2502 (N_2502,N_2487,N_2465);
nand U2503 (N_2503,N_2461,N_2478);
nand U2504 (N_2504,N_2481,N_2488);
nand U2505 (N_2505,N_2452,N_2453);
and U2506 (N_2506,N_2476,N_2468);
or U2507 (N_2507,N_2460,N_2496);
nand U2508 (N_2508,N_2471,N_2491);
nor U2509 (N_2509,N_2492,N_2469);
and U2510 (N_2510,N_2499,N_2467);
nor U2511 (N_2511,N_2472,N_2495);
and U2512 (N_2512,N_2485,N_2466);
nor U2513 (N_2513,N_2489,N_2456);
nand U2514 (N_2514,N_2493,N_2483);
xor U2515 (N_2515,N_2470,N_2477);
nand U2516 (N_2516,N_2455,N_2490);
nor U2517 (N_2517,N_2480,N_2494);
and U2518 (N_2518,N_2484,N_2458);
and U2519 (N_2519,N_2479,N_2457);
or U2520 (N_2520,N_2463,N_2497);
or U2521 (N_2521,N_2450,N_2482);
nor U2522 (N_2522,N_2459,N_2474);
nand U2523 (N_2523,N_2475,N_2464);
nand U2524 (N_2524,N_2462,N_2473);
nand U2525 (N_2525,N_2464,N_2480);
xor U2526 (N_2526,N_2452,N_2461);
nand U2527 (N_2527,N_2497,N_2479);
nand U2528 (N_2528,N_2486,N_2463);
or U2529 (N_2529,N_2496,N_2498);
and U2530 (N_2530,N_2496,N_2478);
nand U2531 (N_2531,N_2492,N_2471);
nand U2532 (N_2532,N_2457,N_2490);
or U2533 (N_2533,N_2461,N_2463);
and U2534 (N_2534,N_2451,N_2484);
nand U2535 (N_2535,N_2462,N_2464);
and U2536 (N_2536,N_2471,N_2497);
or U2537 (N_2537,N_2464,N_2472);
and U2538 (N_2538,N_2477,N_2495);
nand U2539 (N_2539,N_2474,N_2465);
and U2540 (N_2540,N_2489,N_2458);
and U2541 (N_2541,N_2489,N_2460);
or U2542 (N_2542,N_2464,N_2497);
nand U2543 (N_2543,N_2491,N_2494);
and U2544 (N_2544,N_2454,N_2465);
nand U2545 (N_2545,N_2488,N_2459);
nand U2546 (N_2546,N_2472,N_2468);
xnor U2547 (N_2547,N_2489,N_2494);
nand U2548 (N_2548,N_2468,N_2453);
nor U2549 (N_2549,N_2476,N_2454);
xnor U2550 (N_2550,N_2501,N_2526);
xnor U2551 (N_2551,N_2517,N_2544);
nand U2552 (N_2552,N_2529,N_2527);
nor U2553 (N_2553,N_2537,N_2541);
nand U2554 (N_2554,N_2539,N_2508);
nand U2555 (N_2555,N_2548,N_2521);
and U2556 (N_2556,N_2519,N_2514);
and U2557 (N_2557,N_2533,N_2549);
nand U2558 (N_2558,N_2522,N_2518);
or U2559 (N_2559,N_2540,N_2504);
and U2560 (N_2560,N_2511,N_2506);
and U2561 (N_2561,N_2500,N_2532);
nand U2562 (N_2562,N_2520,N_2538);
nor U2563 (N_2563,N_2509,N_2546);
and U2564 (N_2564,N_2542,N_2512);
and U2565 (N_2565,N_2547,N_2513);
nand U2566 (N_2566,N_2536,N_2534);
or U2567 (N_2567,N_2505,N_2543);
or U2568 (N_2568,N_2545,N_2530);
and U2569 (N_2569,N_2528,N_2531);
nand U2570 (N_2570,N_2516,N_2503);
or U2571 (N_2571,N_2515,N_2507);
or U2572 (N_2572,N_2510,N_2502);
nand U2573 (N_2573,N_2524,N_2525);
nor U2574 (N_2574,N_2535,N_2523);
and U2575 (N_2575,N_2543,N_2518);
nor U2576 (N_2576,N_2500,N_2510);
and U2577 (N_2577,N_2509,N_2538);
xnor U2578 (N_2578,N_2517,N_2511);
or U2579 (N_2579,N_2532,N_2545);
nand U2580 (N_2580,N_2546,N_2528);
and U2581 (N_2581,N_2510,N_2548);
nand U2582 (N_2582,N_2526,N_2533);
and U2583 (N_2583,N_2519,N_2521);
nand U2584 (N_2584,N_2525,N_2538);
or U2585 (N_2585,N_2541,N_2536);
nand U2586 (N_2586,N_2515,N_2539);
and U2587 (N_2587,N_2513,N_2509);
or U2588 (N_2588,N_2516,N_2528);
and U2589 (N_2589,N_2503,N_2526);
nand U2590 (N_2590,N_2537,N_2534);
xnor U2591 (N_2591,N_2532,N_2542);
or U2592 (N_2592,N_2526,N_2540);
nor U2593 (N_2593,N_2517,N_2501);
and U2594 (N_2594,N_2506,N_2523);
nand U2595 (N_2595,N_2548,N_2539);
and U2596 (N_2596,N_2513,N_2522);
nor U2597 (N_2597,N_2521,N_2501);
and U2598 (N_2598,N_2510,N_2522);
and U2599 (N_2599,N_2532,N_2546);
and U2600 (N_2600,N_2595,N_2574);
or U2601 (N_2601,N_2573,N_2581);
nand U2602 (N_2602,N_2562,N_2557);
nand U2603 (N_2603,N_2551,N_2568);
nand U2604 (N_2604,N_2559,N_2579);
nand U2605 (N_2605,N_2560,N_2594);
and U2606 (N_2606,N_2550,N_2566);
nor U2607 (N_2607,N_2590,N_2575);
or U2608 (N_2608,N_2591,N_2565);
or U2609 (N_2609,N_2597,N_2584);
nor U2610 (N_2610,N_2558,N_2578);
nor U2611 (N_2611,N_2582,N_2585);
or U2612 (N_2612,N_2556,N_2599);
nand U2613 (N_2613,N_2586,N_2583);
or U2614 (N_2614,N_2571,N_2592);
nand U2615 (N_2615,N_2553,N_2563);
or U2616 (N_2616,N_2555,N_2598);
or U2617 (N_2617,N_2561,N_2572);
and U2618 (N_2618,N_2589,N_2577);
nor U2619 (N_2619,N_2587,N_2576);
and U2620 (N_2620,N_2564,N_2580);
nor U2621 (N_2621,N_2554,N_2588);
or U2622 (N_2622,N_2570,N_2596);
and U2623 (N_2623,N_2567,N_2552);
nor U2624 (N_2624,N_2593,N_2569);
nand U2625 (N_2625,N_2599,N_2583);
and U2626 (N_2626,N_2553,N_2566);
nand U2627 (N_2627,N_2557,N_2585);
and U2628 (N_2628,N_2583,N_2594);
or U2629 (N_2629,N_2579,N_2569);
nand U2630 (N_2630,N_2559,N_2564);
nand U2631 (N_2631,N_2592,N_2574);
and U2632 (N_2632,N_2586,N_2599);
and U2633 (N_2633,N_2559,N_2556);
or U2634 (N_2634,N_2575,N_2567);
or U2635 (N_2635,N_2588,N_2590);
nand U2636 (N_2636,N_2559,N_2558);
nor U2637 (N_2637,N_2591,N_2586);
nor U2638 (N_2638,N_2559,N_2577);
nand U2639 (N_2639,N_2593,N_2562);
or U2640 (N_2640,N_2587,N_2573);
nor U2641 (N_2641,N_2583,N_2577);
and U2642 (N_2642,N_2595,N_2571);
and U2643 (N_2643,N_2565,N_2588);
nor U2644 (N_2644,N_2551,N_2556);
and U2645 (N_2645,N_2551,N_2581);
or U2646 (N_2646,N_2555,N_2576);
and U2647 (N_2647,N_2596,N_2562);
and U2648 (N_2648,N_2590,N_2560);
xor U2649 (N_2649,N_2569,N_2578);
nor U2650 (N_2650,N_2634,N_2622);
nand U2651 (N_2651,N_2614,N_2649);
or U2652 (N_2652,N_2601,N_2619);
or U2653 (N_2653,N_2644,N_2610);
nor U2654 (N_2654,N_2621,N_2616);
and U2655 (N_2655,N_2602,N_2611);
nand U2656 (N_2656,N_2606,N_2636);
nand U2657 (N_2657,N_2626,N_2618);
or U2658 (N_2658,N_2642,N_2632);
and U2659 (N_2659,N_2639,N_2600);
nor U2660 (N_2660,N_2605,N_2608);
or U2661 (N_2661,N_2623,N_2607);
nand U2662 (N_2662,N_2641,N_2645);
nor U2663 (N_2663,N_2647,N_2630);
nor U2664 (N_2664,N_2624,N_2603);
nor U2665 (N_2665,N_2643,N_2612);
nor U2666 (N_2666,N_2638,N_2615);
nor U2667 (N_2667,N_2625,N_2648);
nor U2668 (N_2668,N_2640,N_2637);
nor U2669 (N_2669,N_2617,N_2604);
and U2670 (N_2670,N_2627,N_2629);
and U2671 (N_2671,N_2635,N_2609);
or U2672 (N_2672,N_2628,N_2613);
nand U2673 (N_2673,N_2631,N_2620);
nand U2674 (N_2674,N_2633,N_2646);
nor U2675 (N_2675,N_2640,N_2636);
or U2676 (N_2676,N_2623,N_2635);
nand U2677 (N_2677,N_2603,N_2617);
or U2678 (N_2678,N_2602,N_2619);
nand U2679 (N_2679,N_2600,N_2636);
nor U2680 (N_2680,N_2630,N_2644);
or U2681 (N_2681,N_2610,N_2617);
nor U2682 (N_2682,N_2612,N_2630);
nand U2683 (N_2683,N_2641,N_2642);
nand U2684 (N_2684,N_2636,N_2647);
nor U2685 (N_2685,N_2614,N_2622);
or U2686 (N_2686,N_2606,N_2604);
and U2687 (N_2687,N_2620,N_2635);
nor U2688 (N_2688,N_2612,N_2637);
nand U2689 (N_2689,N_2626,N_2632);
and U2690 (N_2690,N_2640,N_2644);
and U2691 (N_2691,N_2603,N_2640);
or U2692 (N_2692,N_2624,N_2632);
nor U2693 (N_2693,N_2619,N_2641);
or U2694 (N_2694,N_2644,N_2616);
or U2695 (N_2695,N_2610,N_2618);
nand U2696 (N_2696,N_2615,N_2611);
nor U2697 (N_2697,N_2603,N_2641);
nand U2698 (N_2698,N_2606,N_2643);
or U2699 (N_2699,N_2629,N_2600);
or U2700 (N_2700,N_2685,N_2652);
and U2701 (N_2701,N_2650,N_2691);
nand U2702 (N_2702,N_2662,N_2696);
nor U2703 (N_2703,N_2697,N_2677);
nor U2704 (N_2704,N_2689,N_2660);
or U2705 (N_2705,N_2658,N_2693);
nor U2706 (N_2706,N_2665,N_2666);
nor U2707 (N_2707,N_2684,N_2663);
and U2708 (N_2708,N_2656,N_2699);
or U2709 (N_2709,N_2688,N_2698);
nand U2710 (N_2710,N_2664,N_2686);
and U2711 (N_2711,N_2687,N_2671);
or U2712 (N_2712,N_2673,N_2659);
and U2713 (N_2713,N_2680,N_2654);
and U2714 (N_2714,N_2694,N_2676);
and U2715 (N_2715,N_2692,N_2674);
and U2716 (N_2716,N_2653,N_2655);
or U2717 (N_2717,N_2679,N_2682);
nand U2718 (N_2718,N_2670,N_2661);
nor U2719 (N_2719,N_2668,N_2651);
nor U2720 (N_2720,N_2695,N_2678);
or U2721 (N_2721,N_2667,N_2683);
or U2722 (N_2722,N_2690,N_2675);
nand U2723 (N_2723,N_2681,N_2669);
or U2724 (N_2724,N_2657,N_2672);
or U2725 (N_2725,N_2681,N_2682);
or U2726 (N_2726,N_2690,N_2668);
and U2727 (N_2727,N_2657,N_2680);
or U2728 (N_2728,N_2650,N_2679);
and U2729 (N_2729,N_2689,N_2673);
nand U2730 (N_2730,N_2672,N_2683);
and U2731 (N_2731,N_2692,N_2684);
or U2732 (N_2732,N_2687,N_2653);
nand U2733 (N_2733,N_2676,N_2665);
nand U2734 (N_2734,N_2654,N_2675);
nor U2735 (N_2735,N_2691,N_2681);
and U2736 (N_2736,N_2690,N_2689);
nand U2737 (N_2737,N_2652,N_2669);
nor U2738 (N_2738,N_2675,N_2665);
or U2739 (N_2739,N_2661,N_2690);
nor U2740 (N_2740,N_2685,N_2680);
nor U2741 (N_2741,N_2698,N_2671);
or U2742 (N_2742,N_2692,N_2689);
xnor U2743 (N_2743,N_2660,N_2673);
and U2744 (N_2744,N_2679,N_2653);
nor U2745 (N_2745,N_2675,N_2685);
or U2746 (N_2746,N_2656,N_2662);
xor U2747 (N_2747,N_2674,N_2696);
and U2748 (N_2748,N_2682,N_2685);
and U2749 (N_2749,N_2654,N_2653);
or U2750 (N_2750,N_2733,N_2735);
nand U2751 (N_2751,N_2730,N_2705);
nor U2752 (N_2752,N_2711,N_2729);
nor U2753 (N_2753,N_2739,N_2747);
nor U2754 (N_2754,N_2722,N_2701);
and U2755 (N_2755,N_2734,N_2702);
nor U2756 (N_2756,N_2745,N_2717);
and U2757 (N_2757,N_2703,N_2736);
nor U2758 (N_2758,N_2746,N_2708);
nor U2759 (N_2759,N_2720,N_2741);
or U2760 (N_2760,N_2712,N_2738);
or U2761 (N_2761,N_2704,N_2727);
nor U2762 (N_2762,N_2725,N_2724);
or U2763 (N_2763,N_2706,N_2721);
and U2764 (N_2764,N_2715,N_2719);
nor U2765 (N_2765,N_2732,N_2713);
nand U2766 (N_2766,N_2731,N_2744);
and U2767 (N_2767,N_2737,N_2743);
nor U2768 (N_2768,N_2726,N_2740);
and U2769 (N_2769,N_2707,N_2716);
nor U2770 (N_2770,N_2748,N_2728);
nor U2771 (N_2771,N_2742,N_2700);
nor U2772 (N_2772,N_2718,N_2749);
nand U2773 (N_2773,N_2723,N_2709);
nand U2774 (N_2774,N_2710,N_2714);
nor U2775 (N_2775,N_2726,N_2725);
nand U2776 (N_2776,N_2706,N_2726);
or U2777 (N_2777,N_2724,N_2742);
nand U2778 (N_2778,N_2735,N_2712);
nor U2779 (N_2779,N_2723,N_2744);
or U2780 (N_2780,N_2721,N_2720);
nand U2781 (N_2781,N_2710,N_2726);
nand U2782 (N_2782,N_2718,N_2726);
and U2783 (N_2783,N_2749,N_2740);
and U2784 (N_2784,N_2713,N_2747);
nand U2785 (N_2785,N_2743,N_2714);
or U2786 (N_2786,N_2740,N_2724);
or U2787 (N_2787,N_2701,N_2749);
nand U2788 (N_2788,N_2729,N_2714);
and U2789 (N_2789,N_2744,N_2720);
or U2790 (N_2790,N_2725,N_2747);
and U2791 (N_2791,N_2719,N_2708);
nand U2792 (N_2792,N_2744,N_2719);
and U2793 (N_2793,N_2740,N_2703);
or U2794 (N_2794,N_2715,N_2717);
and U2795 (N_2795,N_2735,N_2747);
or U2796 (N_2796,N_2737,N_2746);
or U2797 (N_2797,N_2711,N_2720);
nor U2798 (N_2798,N_2744,N_2732);
or U2799 (N_2799,N_2708,N_2745);
or U2800 (N_2800,N_2785,N_2755);
nand U2801 (N_2801,N_2784,N_2780);
xor U2802 (N_2802,N_2753,N_2790);
nand U2803 (N_2803,N_2788,N_2795);
nand U2804 (N_2804,N_2765,N_2760);
or U2805 (N_2805,N_2787,N_2772);
nor U2806 (N_2806,N_2782,N_2789);
or U2807 (N_2807,N_2775,N_2773);
nor U2808 (N_2808,N_2777,N_2776);
or U2809 (N_2809,N_2783,N_2757);
nor U2810 (N_2810,N_2768,N_2762);
nor U2811 (N_2811,N_2766,N_2786);
or U2812 (N_2812,N_2796,N_2764);
or U2813 (N_2813,N_2752,N_2798);
or U2814 (N_2814,N_2763,N_2767);
xor U2815 (N_2815,N_2756,N_2799);
nand U2816 (N_2816,N_2791,N_2761);
nand U2817 (N_2817,N_2771,N_2794);
or U2818 (N_2818,N_2793,N_2797);
or U2819 (N_2819,N_2758,N_2770);
nand U2820 (N_2820,N_2778,N_2779);
nor U2821 (N_2821,N_2781,N_2754);
xor U2822 (N_2822,N_2750,N_2751);
nor U2823 (N_2823,N_2792,N_2759);
nor U2824 (N_2824,N_2774,N_2769);
and U2825 (N_2825,N_2765,N_2773);
or U2826 (N_2826,N_2751,N_2767);
and U2827 (N_2827,N_2776,N_2753);
or U2828 (N_2828,N_2765,N_2798);
xnor U2829 (N_2829,N_2758,N_2763);
nand U2830 (N_2830,N_2765,N_2781);
nor U2831 (N_2831,N_2798,N_2761);
or U2832 (N_2832,N_2763,N_2789);
nor U2833 (N_2833,N_2781,N_2767);
or U2834 (N_2834,N_2756,N_2797);
xnor U2835 (N_2835,N_2772,N_2770);
or U2836 (N_2836,N_2767,N_2789);
or U2837 (N_2837,N_2765,N_2768);
nand U2838 (N_2838,N_2764,N_2777);
nand U2839 (N_2839,N_2792,N_2780);
nor U2840 (N_2840,N_2752,N_2769);
or U2841 (N_2841,N_2752,N_2771);
nand U2842 (N_2842,N_2752,N_2750);
or U2843 (N_2843,N_2771,N_2792);
xnor U2844 (N_2844,N_2796,N_2776);
and U2845 (N_2845,N_2792,N_2785);
and U2846 (N_2846,N_2767,N_2750);
nor U2847 (N_2847,N_2763,N_2793);
nand U2848 (N_2848,N_2779,N_2774);
and U2849 (N_2849,N_2793,N_2786);
nor U2850 (N_2850,N_2802,N_2837);
or U2851 (N_2851,N_2815,N_2818);
or U2852 (N_2852,N_2836,N_2812);
nor U2853 (N_2853,N_2801,N_2828);
or U2854 (N_2854,N_2829,N_2806);
or U2855 (N_2855,N_2816,N_2838);
and U2856 (N_2856,N_2813,N_2833);
nor U2857 (N_2857,N_2830,N_2804);
nor U2858 (N_2858,N_2846,N_2824);
nor U2859 (N_2859,N_2807,N_2821);
and U2860 (N_2860,N_2844,N_2820);
nor U2861 (N_2861,N_2803,N_2832);
nand U2862 (N_2862,N_2835,N_2805);
or U2863 (N_2863,N_2839,N_2840);
nor U2864 (N_2864,N_2834,N_2848);
nor U2865 (N_2865,N_2814,N_2809);
nand U2866 (N_2866,N_2843,N_2823);
nand U2867 (N_2867,N_2845,N_2819);
or U2868 (N_2868,N_2800,N_2847);
nand U2869 (N_2869,N_2822,N_2849);
nand U2870 (N_2870,N_2825,N_2842);
nor U2871 (N_2871,N_2808,N_2811);
or U2872 (N_2872,N_2810,N_2817);
and U2873 (N_2873,N_2841,N_2831);
or U2874 (N_2874,N_2826,N_2827);
nand U2875 (N_2875,N_2815,N_2813);
nand U2876 (N_2876,N_2848,N_2817);
nor U2877 (N_2877,N_2846,N_2808);
or U2878 (N_2878,N_2810,N_2813);
or U2879 (N_2879,N_2847,N_2839);
nor U2880 (N_2880,N_2829,N_2841);
or U2881 (N_2881,N_2834,N_2825);
or U2882 (N_2882,N_2817,N_2813);
nor U2883 (N_2883,N_2827,N_2833);
xnor U2884 (N_2884,N_2842,N_2805);
nand U2885 (N_2885,N_2848,N_2827);
and U2886 (N_2886,N_2801,N_2803);
nor U2887 (N_2887,N_2833,N_2837);
and U2888 (N_2888,N_2845,N_2835);
or U2889 (N_2889,N_2831,N_2824);
nor U2890 (N_2890,N_2800,N_2815);
or U2891 (N_2891,N_2827,N_2837);
nand U2892 (N_2892,N_2822,N_2828);
and U2893 (N_2893,N_2834,N_2846);
nand U2894 (N_2894,N_2834,N_2843);
nor U2895 (N_2895,N_2804,N_2828);
xnor U2896 (N_2896,N_2832,N_2828);
nand U2897 (N_2897,N_2835,N_2849);
and U2898 (N_2898,N_2823,N_2835);
or U2899 (N_2899,N_2817,N_2808);
nand U2900 (N_2900,N_2878,N_2898);
nand U2901 (N_2901,N_2867,N_2881);
or U2902 (N_2902,N_2897,N_2857);
nor U2903 (N_2903,N_2854,N_2870);
or U2904 (N_2904,N_2863,N_2895);
or U2905 (N_2905,N_2861,N_2896);
or U2906 (N_2906,N_2873,N_2875);
nand U2907 (N_2907,N_2865,N_2877);
nor U2908 (N_2908,N_2850,N_2890);
and U2909 (N_2909,N_2891,N_2882);
xnor U2910 (N_2910,N_2866,N_2893);
nor U2911 (N_2911,N_2894,N_2856);
nor U2912 (N_2912,N_2855,N_2889);
nor U2913 (N_2913,N_2885,N_2851);
or U2914 (N_2914,N_2879,N_2872);
nor U2915 (N_2915,N_2864,N_2888);
or U2916 (N_2916,N_2859,N_2884);
or U2917 (N_2917,N_2874,N_2876);
xnor U2918 (N_2918,N_2880,N_2886);
or U2919 (N_2919,N_2869,N_2868);
nor U2920 (N_2920,N_2853,N_2887);
nor U2921 (N_2921,N_2871,N_2899);
or U2922 (N_2922,N_2862,N_2892);
nor U2923 (N_2923,N_2858,N_2852);
or U2924 (N_2924,N_2883,N_2860);
nor U2925 (N_2925,N_2852,N_2880);
nor U2926 (N_2926,N_2869,N_2895);
nand U2927 (N_2927,N_2899,N_2865);
or U2928 (N_2928,N_2871,N_2857);
and U2929 (N_2929,N_2893,N_2854);
nand U2930 (N_2930,N_2854,N_2897);
nor U2931 (N_2931,N_2886,N_2854);
and U2932 (N_2932,N_2861,N_2865);
or U2933 (N_2933,N_2891,N_2895);
and U2934 (N_2934,N_2879,N_2890);
and U2935 (N_2935,N_2855,N_2852);
and U2936 (N_2936,N_2893,N_2882);
nand U2937 (N_2937,N_2864,N_2863);
nor U2938 (N_2938,N_2890,N_2856);
or U2939 (N_2939,N_2852,N_2894);
and U2940 (N_2940,N_2877,N_2872);
nor U2941 (N_2941,N_2891,N_2880);
or U2942 (N_2942,N_2857,N_2889);
nor U2943 (N_2943,N_2889,N_2859);
and U2944 (N_2944,N_2867,N_2861);
nand U2945 (N_2945,N_2877,N_2852);
or U2946 (N_2946,N_2855,N_2880);
or U2947 (N_2947,N_2889,N_2881);
nand U2948 (N_2948,N_2883,N_2885);
nand U2949 (N_2949,N_2867,N_2856);
and U2950 (N_2950,N_2949,N_2915);
or U2951 (N_2951,N_2908,N_2940);
and U2952 (N_2952,N_2932,N_2905);
nand U2953 (N_2953,N_2931,N_2902);
nor U2954 (N_2954,N_2924,N_2937);
nor U2955 (N_2955,N_2909,N_2918);
or U2956 (N_2956,N_2938,N_2930);
nand U2957 (N_2957,N_2947,N_2903);
and U2958 (N_2958,N_2941,N_2943);
nand U2959 (N_2959,N_2935,N_2928);
or U2960 (N_2960,N_2934,N_2900);
and U2961 (N_2961,N_2922,N_2911);
nor U2962 (N_2962,N_2901,N_2917);
or U2963 (N_2963,N_2948,N_2912);
or U2964 (N_2964,N_2914,N_2904);
or U2965 (N_2965,N_2929,N_2945);
nand U2966 (N_2966,N_2916,N_2927);
nor U2967 (N_2967,N_2913,N_2942);
nand U2968 (N_2968,N_2906,N_2944);
and U2969 (N_2969,N_2919,N_2946);
nor U2970 (N_2970,N_2910,N_2923);
nand U2971 (N_2971,N_2939,N_2933);
nor U2972 (N_2972,N_2920,N_2907);
nand U2973 (N_2973,N_2926,N_2921);
or U2974 (N_2974,N_2936,N_2925);
nand U2975 (N_2975,N_2938,N_2935);
nand U2976 (N_2976,N_2921,N_2903);
or U2977 (N_2977,N_2914,N_2942);
xnor U2978 (N_2978,N_2913,N_2938);
and U2979 (N_2979,N_2948,N_2943);
nand U2980 (N_2980,N_2900,N_2909);
nor U2981 (N_2981,N_2927,N_2929);
nand U2982 (N_2982,N_2926,N_2932);
nand U2983 (N_2983,N_2912,N_2941);
nand U2984 (N_2984,N_2917,N_2946);
nor U2985 (N_2985,N_2925,N_2915);
or U2986 (N_2986,N_2907,N_2902);
nand U2987 (N_2987,N_2902,N_2937);
or U2988 (N_2988,N_2936,N_2942);
xor U2989 (N_2989,N_2903,N_2942);
nor U2990 (N_2990,N_2900,N_2924);
or U2991 (N_2991,N_2934,N_2918);
nand U2992 (N_2992,N_2920,N_2930);
xor U2993 (N_2993,N_2928,N_2949);
nand U2994 (N_2994,N_2941,N_2902);
nand U2995 (N_2995,N_2903,N_2914);
or U2996 (N_2996,N_2914,N_2947);
nand U2997 (N_2997,N_2948,N_2928);
and U2998 (N_2998,N_2902,N_2943);
xor U2999 (N_2999,N_2940,N_2901);
nor UO_0 (O_0,N_2966,N_2971);
and UO_1 (O_1,N_2992,N_2958);
nand UO_2 (O_2,N_2974,N_2993);
or UO_3 (O_3,N_2994,N_2990);
nor UO_4 (O_4,N_2962,N_2998);
and UO_5 (O_5,N_2996,N_2987);
or UO_6 (O_6,N_2964,N_2973);
nand UO_7 (O_7,N_2988,N_2978);
nand UO_8 (O_8,N_2975,N_2955);
and UO_9 (O_9,N_2953,N_2968);
nand UO_10 (O_10,N_2980,N_2969);
or UO_11 (O_11,N_2982,N_2952);
and UO_12 (O_12,N_2967,N_2960);
and UO_13 (O_13,N_2959,N_2950);
nand UO_14 (O_14,N_2956,N_2963);
or UO_15 (O_15,N_2972,N_2986);
nor UO_16 (O_16,N_2970,N_2984);
and UO_17 (O_17,N_2983,N_2989);
and UO_18 (O_18,N_2981,N_2979);
or UO_19 (O_19,N_2991,N_2997);
and UO_20 (O_20,N_2995,N_2957);
xor UO_21 (O_21,N_2961,N_2999);
nor UO_22 (O_22,N_2985,N_2954);
or UO_23 (O_23,N_2976,N_2951);
nor UO_24 (O_24,N_2977,N_2965);
xor UO_25 (O_25,N_2990,N_2989);
nor UO_26 (O_26,N_2962,N_2986);
nor UO_27 (O_27,N_2952,N_2954);
nand UO_28 (O_28,N_2952,N_2953);
or UO_29 (O_29,N_2963,N_2958);
or UO_30 (O_30,N_2982,N_2966);
nor UO_31 (O_31,N_2980,N_2997);
xor UO_32 (O_32,N_2994,N_2996);
or UO_33 (O_33,N_2987,N_2952);
nor UO_34 (O_34,N_2974,N_2967);
and UO_35 (O_35,N_2972,N_2971);
nand UO_36 (O_36,N_2953,N_2989);
and UO_37 (O_37,N_2992,N_2993);
or UO_38 (O_38,N_2993,N_2991);
or UO_39 (O_39,N_2997,N_2994);
nor UO_40 (O_40,N_2955,N_2987);
or UO_41 (O_41,N_2990,N_2981);
nand UO_42 (O_42,N_2955,N_2978);
and UO_43 (O_43,N_2997,N_2993);
and UO_44 (O_44,N_2988,N_2998);
nand UO_45 (O_45,N_2973,N_2977);
nor UO_46 (O_46,N_2962,N_2954);
or UO_47 (O_47,N_2954,N_2994);
nor UO_48 (O_48,N_2985,N_2986);
and UO_49 (O_49,N_2953,N_2985);
or UO_50 (O_50,N_2988,N_2951);
and UO_51 (O_51,N_2963,N_2969);
nor UO_52 (O_52,N_2960,N_2997);
nor UO_53 (O_53,N_2986,N_2996);
and UO_54 (O_54,N_2976,N_2963);
or UO_55 (O_55,N_2960,N_2990);
or UO_56 (O_56,N_2981,N_2997);
nor UO_57 (O_57,N_2965,N_2979);
and UO_58 (O_58,N_2959,N_2992);
or UO_59 (O_59,N_2992,N_2996);
and UO_60 (O_60,N_2995,N_2969);
nand UO_61 (O_61,N_2981,N_2983);
or UO_62 (O_62,N_2953,N_2999);
or UO_63 (O_63,N_2962,N_2991);
nand UO_64 (O_64,N_2980,N_2972);
nand UO_65 (O_65,N_2973,N_2972);
or UO_66 (O_66,N_2958,N_2955);
and UO_67 (O_67,N_2962,N_2969);
or UO_68 (O_68,N_2999,N_2981);
and UO_69 (O_69,N_2976,N_2975);
nand UO_70 (O_70,N_2967,N_2976);
nor UO_71 (O_71,N_2998,N_2980);
nor UO_72 (O_72,N_2986,N_2958);
nor UO_73 (O_73,N_2988,N_2974);
and UO_74 (O_74,N_2969,N_2956);
or UO_75 (O_75,N_2995,N_2996);
nor UO_76 (O_76,N_2973,N_2954);
or UO_77 (O_77,N_2965,N_2987);
nor UO_78 (O_78,N_2996,N_2969);
nand UO_79 (O_79,N_2968,N_2962);
nor UO_80 (O_80,N_2950,N_2974);
nand UO_81 (O_81,N_2981,N_2996);
nor UO_82 (O_82,N_2997,N_2999);
and UO_83 (O_83,N_2957,N_2968);
or UO_84 (O_84,N_2953,N_2977);
nand UO_85 (O_85,N_2985,N_2951);
and UO_86 (O_86,N_2959,N_2974);
nor UO_87 (O_87,N_2964,N_2959);
or UO_88 (O_88,N_2996,N_2993);
nand UO_89 (O_89,N_2982,N_2998);
xor UO_90 (O_90,N_2959,N_2976);
nand UO_91 (O_91,N_2961,N_2975);
nor UO_92 (O_92,N_2964,N_2953);
nor UO_93 (O_93,N_2973,N_2951);
or UO_94 (O_94,N_2958,N_2984);
or UO_95 (O_95,N_2961,N_2990);
and UO_96 (O_96,N_2993,N_2978);
and UO_97 (O_97,N_2974,N_2991);
nand UO_98 (O_98,N_2967,N_2994);
or UO_99 (O_99,N_2969,N_2988);
and UO_100 (O_100,N_2992,N_2988);
nand UO_101 (O_101,N_2977,N_2956);
xnor UO_102 (O_102,N_2961,N_2996);
nand UO_103 (O_103,N_2952,N_2951);
and UO_104 (O_104,N_2963,N_2979);
or UO_105 (O_105,N_2960,N_2963);
nand UO_106 (O_106,N_2956,N_2971);
nor UO_107 (O_107,N_2989,N_2982);
or UO_108 (O_108,N_2960,N_2978);
or UO_109 (O_109,N_2959,N_2957);
or UO_110 (O_110,N_2997,N_2989);
and UO_111 (O_111,N_2991,N_2961);
nand UO_112 (O_112,N_2957,N_2985);
nor UO_113 (O_113,N_2984,N_2972);
or UO_114 (O_114,N_2957,N_2975);
nand UO_115 (O_115,N_2969,N_2952);
and UO_116 (O_116,N_2973,N_2961);
nor UO_117 (O_117,N_2959,N_2982);
nor UO_118 (O_118,N_2992,N_2971);
or UO_119 (O_119,N_2963,N_2957);
nand UO_120 (O_120,N_2996,N_2975);
or UO_121 (O_121,N_2997,N_2976);
or UO_122 (O_122,N_2977,N_2994);
nand UO_123 (O_123,N_2971,N_2983);
nor UO_124 (O_124,N_2970,N_2965);
nor UO_125 (O_125,N_2972,N_2963);
nand UO_126 (O_126,N_2979,N_2952);
or UO_127 (O_127,N_2980,N_2964);
or UO_128 (O_128,N_2985,N_2988);
and UO_129 (O_129,N_2975,N_2952);
and UO_130 (O_130,N_2962,N_2950);
nand UO_131 (O_131,N_2967,N_2961);
nand UO_132 (O_132,N_2995,N_2984);
and UO_133 (O_133,N_2968,N_2966);
nor UO_134 (O_134,N_2977,N_2978);
nor UO_135 (O_135,N_2999,N_2954);
nand UO_136 (O_136,N_2950,N_2951);
nor UO_137 (O_137,N_2980,N_2982);
and UO_138 (O_138,N_2967,N_2987);
or UO_139 (O_139,N_2995,N_2986);
or UO_140 (O_140,N_2952,N_2988);
nor UO_141 (O_141,N_2992,N_2978);
or UO_142 (O_142,N_2993,N_2959);
nor UO_143 (O_143,N_2951,N_2974);
and UO_144 (O_144,N_2995,N_2970);
and UO_145 (O_145,N_2999,N_2952);
nor UO_146 (O_146,N_2960,N_2981);
or UO_147 (O_147,N_2962,N_2997);
and UO_148 (O_148,N_2987,N_2992);
nand UO_149 (O_149,N_2964,N_2988);
nand UO_150 (O_150,N_2984,N_2964);
or UO_151 (O_151,N_2998,N_2974);
nor UO_152 (O_152,N_2965,N_2968);
or UO_153 (O_153,N_2973,N_2952);
and UO_154 (O_154,N_2994,N_2991);
or UO_155 (O_155,N_2983,N_2996);
or UO_156 (O_156,N_2974,N_2973);
and UO_157 (O_157,N_2967,N_2996);
nand UO_158 (O_158,N_2987,N_2995);
and UO_159 (O_159,N_2954,N_2961);
or UO_160 (O_160,N_2990,N_2979);
or UO_161 (O_161,N_2950,N_2984);
nand UO_162 (O_162,N_2980,N_2975);
nor UO_163 (O_163,N_2980,N_2989);
nand UO_164 (O_164,N_2997,N_2963);
and UO_165 (O_165,N_2953,N_2991);
nand UO_166 (O_166,N_2981,N_2970);
or UO_167 (O_167,N_2951,N_2977);
and UO_168 (O_168,N_2967,N_2965);
nor UO_169 (O_169,N_2958,N_2991);
and UO_170 (O_170,N_2988,N_2970);
or UO_171 (O_171,N_2998,N_2971);
or UO_172 (O_172,N_2978,N_2976);
nand UO_173 (O_173,N_2968,N_2981);
nand UO_174 (O_174,N_2956,N_2950);
nand UO_175 (O_175,N_2987,N_2956);
and UO_176 (O_176,N_2950,N_2952);
or UO_177 (O_177,N_2996,N_2974);
and UO_178 (O_178,N_2967,N_2998);
and UO_179 (O_179,N_2979,N_2985);
xor UO_180 (O_180,N_2969,N_2999);
and UO_181 (O_181,N_2958,N_2966);
or UO_182 (O_182,N_2960,N_2984);
nor UO_183 (O_183,N_2953,N_2995);
or UO_184 (O_184,N_2991,N_2957);
nor UO_185 (O_185,N_2985,N_2967);
nor UO_186 (O_186,N_2962,N_2989);
nand UO_187 (O_187,N_2980,N_2996);
or UO_188 (O_188,N_2968,N_2988);
nand UO_189 (O_189,N_2955,N_2985);
or UO_190 (O_190,N_2961,N_2965);
nor UO_191 (O_191,N_2963,N_2962);
nand UO_192 (O_192,N_2953,N_2972);
nor UO_193 (O_193,N_2957,N_2988);
and UO_194 (O_194,N_2973,N_2962);
nor UO_195 (O_195,N_2956,N_2980);
nand UO_196 (O_196,N_2992,N_2965);
and UO_197 (O_197,N_2981,N_2975);
and UO_198 (O_198,N_2971,N_2976);
nor UO_199 (O_199,N_2956,N_2976);
xor UO_200 (O_200,N_2971,N_2953);
nand UO_201 (O_201,N_2986,N_2997);
nor UO_202 (O_202,N_2981,N_2951);
or UO_203 (O_203,N_2960,N_2956);
nor UO_204 (O_204,N_2987,N_2968);
or UO_205 (O_205,N_2979,N_2983);
nor UO_206 (O_206,N_2974,N_2968);
and UO_207 (O_207,N_2978,N_2990);
and UO_208 (O_208,N_2958,N_2994);
and UO_209 (O_209,N_2993,N_2969);
nor UO_210 (O_210,N_2972,N_2966);
nor UO_211 (O_211,N_2968,N_2970);
nand UO_212 (O_212,N_2963,N_2983);
or UO_213 (O_213,N_2976,N_2996);
nand UO_214 (O_214,N_2985,N_2956);
and UO_215 (O_215,N_2990,N_2957);
nand UO_216 (O_216,N_2988,N_2966);
nor UO_217 (O_217,N_2993,N_2981);
nand UO_218 (O_218,N_2980,N_2973);
and UO_219 (O_219,N_2995,N_2971);
or UO_220 (O_220,N_2961,N_2955);
or UO_221 (O_221,N_2977,N_2979);
and UO_222 (O_222,N_2979,N_2951);
nand UO_223 (O_223,N_2977,N_2967);
and UO_224 (O_224,N_2994,N_2968);
nand UO_225 (O_225,N_2960,N_2971);
or UO_226 (O_226,N_2969,N_2965);
or UO_227 (O_227,N_2975,N_2987);
nand UO_228 (O_228,N_2981,N_2961);
or UO_229 (O_229,N_2977,N_2983);
nand UO_230 (O_230,N_2964,N_2995);
nand UO_231 (O_231,N_2972,N_2969);
nand UO_232 (O_232,N_2988,N_2954);
and UO_233 (O_233,N_2965,N_2971);
or UO_234 (O_234,N_2957,N_2970);
nor UO_235 (O_235,N_2984,N_2957);
and UO_236 (O_236,N_2997,N_2972);
or UO_237 (O_237,N_2992,N_2981);
nor UO_238 (O_238,N_2961,N_2982);
nand UO_239 (O_239,N_2970,N_2976);
or UO_240 (O_240,N_2977,N_2991);
nand UO_241 (O_241,N_2955,N_2999);
nor UO_242 (O_242,N_2980,N_2988);
nor UO_243 (O_243,N_2969,N_2961);
or UO_244 (O_244,N_2994,N_2992);
or UO_245 (O_245,N_2963,N_2989);
and UO_246 (O_246,N_2954,N_2986);
nand UO_247 (O_247,N_2993,N_2983);
or UO_248 (O_248,N_2960,N_2968);
or UO_249 (O_249,N_2973,N_2982);
nor UO_250 (O_250,N_2998,N_2984);
nor UO_251 (O_251,N_2970,N_2950);
nand UO_252 (O_252,N_2986,N_2950);
nand UO_253 (O_253,N_2994,N_2956);
or UO_254 (O_254,N_2963,N_2970);
and UO_255 (O_255,N_2977,N_2968);
and UO_256 (O_256,N_2987,N_2993);
and UO_257 (O_257,N_2965,N_2954);
nand UO_258 (O_258,N_2997,N_2966);
and UO_259 (O_259,N_2963,N_2955);
or UO_260 (O_260,N_2955,N_2972);
and UO_261 (O_261,N_2985,N_2975);
or UO_262 (O_262,N_2985,N_2961);
nand UO_263 (O_263,N_2997,N_2987);
and UO_264 (O_264,N_2973,N_2998);
nor UO_265 (O_265,N_2978,N_2956);
or UO_266 (O_266,N_2991,N_2975);
and UO_267 (O_267,N_2981,N_2966);
or UO_268 (O_268,N_2990,N_2971);
or UO_269 (O_269,N_2951,N_2970);
nor UO_270 (O_270,N_2984,N_2979);
nor UO_271 (O_271,N_2984,N_2991);
nor UO_272 (O_272,N_2998,N_2952);
nor UO_273 (O_273,N_2979,N_2956);
and UO_274 (O_274,N_2959,N_2954);
or UO_275 (O_275,N_2961,N_2997);
or UO_276 (O_276,N_2965,N_2975);
nand UO_277 (O_277,N_2955,N_2960);
nor UO_278 (O_278,N_2994,N_2966);
or UO_279 (O_279,N_2995,N_2982);
nand UO_280 (O_280,N_2959,N_2971);
nand UO_281 (O_281,N_2985,N_2980);
or UO_282 (O_282,N_2960,N_2988);
nand UO_283 (O_283,N_2958,N_2954);
nand UO_284 (O_284,N_2992,N_2984);
nor UO_285 (O_285,N_2955,N_2951);
nand UO_286 (O_286,N_2992,N_2950);
nor UO_287 (O_287,N_2965,N_2960);
nor UO_288 (O_288,N_2996,N_2999);
and UO_289 (O_289,N_2988,N_2981);
or UO_290 (O_290,N_2973,N_2957);
and UO_291 (O_291,N_2965,N_2950);
and UO_292 (O_292,N_2989,N_2965);
nand UO_293 (O_293,N_2996,N_2962);
nand UO_294 (O_294,N_2969,N_2954);
and UO_295 (O_295,N_2951,N_2963);
nor UO_296 (O_296,N_2964,N_2950);
or UO_297 (O_297,N_2999,N_2958);
and UO_298 (O_298,N_2975,N_2982);
nand UO_299 (O_299,N_2958,N_2957);
or UO_300 (O_300,N_2955,N_2968);
nand UO_301 (O_301,N_2960,N_2973);
or UO_302 (O_302,N_2956,N_2975);
nand UO_303 (O_303,N_2963,N_2982);
or UO_304 (O_304,N_2957,N_2972);
and UO_305 (O_305,N_2978,N_2967);
nor UO_306 (O_306,N_2966,N_2955);
nor UO_307 (O_307,N_2972,N_2987);
nor UO_308 (O_308,N_2997,N_2955);
and UO_309 (O_309,N_2993,N_2967);
nor UO_310 (O_310,N_2958,N_2960);
and UO_311 (O_311,N_2987,N_2988);
nand UO_312 (O_312,N_2952,N_2984);
nor UO_313 (O_313,N_2976,N_2990);
nor UO_314 (O_314,N_2999,N_2998);
nor UO_315 (O_315,N_2965,N_2988);
nor UO_316 (O_316,N_2991,N_2966);
xor UO_317 (O_317,N_2959,N_2952);
or UO_318 (O_318,N_2985,N_2966);
and UO_319 (O_319,N_2962,N_2952);
and UO_320 (O_320,N_2964,N_2992);
nand UO_321 (O_321,N_2965,N_2995);
nor UO_322 (O_322,N_2971,N_2952);
and UO_323 (O_323,N_2974,N_2999);
and UO_324 (O_324,N_2964,N_2969);
nand UO_325 (O_325,N_2999,N_2994);
or UO_326 (O_326,N_2990,N_2958);
or UO_327 (O_327,N_2953,N_2951);
nor UO_328 (O_328,N_2953,N_2958);
and UO_329 (O_329,N_2997,N_2985);
or UO_330 (O_330,N_2955,N_2983);
and UO_331 (O_331,N_2955,N_2989);
or UO_332 (O_332,N_2996,N_2956);
nor UO_333 (O_333,N_2977,N_2987);
or UO_334 (O_334,N_2990,N_2982);
nor UO_335 (O_335,N_2967,N_2952);
or UO_336 (O_336,N_2958,N_2975);
and UO_337 (O_337,N_2963,N_2978);
nor UO_338 (O_338,N_2953,N_2994);
nor UO_339 (O_339,N_2999,N_2989);
and UO_340 (O_340,N_2956,N_2999);
or UO_341 (O_341,N_2983,N_2988);
nand UO_342 (O_342,N_2976,N_2965);
nand UO_343 (O_343,N_2975,N_2983);
or UO_344 (O_344,N_2987,N_2964);
nor UO_345 (O_345,N_2988,N_2973);
nor UO_346 (O_346,N_2966,N_2983);
xor UO_347 (O_347,N_2999,N_2991);
and UO_348 (O_348,N_2953,N_2979);
or UO_349 (O_349,N_2999,N_2962);
xnor UO_350 (O_350,N_2974,N_2997);
nor UO_351 (O_351,N_2969,N_2955);
or UO_352 (O_352,N_2989,N_2996);
nor UO_353 (O_353,N_2998,N_2986);
or UO_354 (O_354,N_2955,N_2965);
nand UO_355 (O_355,N_2983,N_2990);
or UO_356 (O_356,N_2998,N_2950);
nor UO_357 (O_357,N_2977,N_2990);
or UO_358 (O_358,N_2962,N_2978);
or UO_359 (O_359,N_2977,N_2988);
and UO_360 (O_360,N_2959,N_2956);
and UO_361 (O_361,N_2971,N_2985);
nand UO_362 (O_362,N_2967,N_2981);
or UO_363 (O_363,N_2974,N_2984);
and UO_364 (O_364,N_2986,N_2988);
nand UO_365 (O_365,N_2952,N_2977);
nor UO_366 (O_366,N_2953,N_2973);
and UO_367 (O_367,N_2952,N_2978);
and UO_368 (O_368,N_2977,N_2999);
nor UO_369 (O_369,N_2977,N_2997);
or UO_370 (O_370,N_2960,N_2969);
nor UO_371 (O_371,N_2982,N_2950);
nand UO_372 (O_372,N_2973,N_2976);
nand UO_373 (O_373,N_2970,N_2962);
and UO_374 (O_374,N_2992,N_2968);
nand UO_375 (O_375,N_2964,N_2993);
nand UO_376 (O_376,N_2988,N_2975);
or UO_377 (O_377,N_2957,N_2994);
or UO_378 (O_378,N_2984,N_2978);
nand UO_379 (O_379,N_2955,N_2984);
or UO_380 (O_380,N_2981,N_2985);
and UO_381 (O_381,N_2985,N_2987);
nor UO_382 (O_382,N_2995,N_2960);
or UO_383 (O_383,N_2972,N_2965);
and UO_384 (O_384,N_2977,N_2966);
or UO_385 (O_385,N_2957,N_2950);
or UO_386 (O_386,N_2978,N_2966);
and UO_387 (O_387,N_2992,N_2982);
nand UO_388 (O_388,N_2953,N_2990);
nor UO_389 (O_389,N_2988,N_2994);
nand UO_390 (O_390,N_2977,N_2955);
or UO_391 (O_391,N_2990,N_2967);
or UO_392 (O_392,N_2955,N_2971);
and UO_393 (O_393,N_2972,N_2951);
nand UO_394 (O_394,N_2958,N_2962);
nand UO_395 (O_395,N_2982,N_2964);
or UO_396 (O_396,N_2958,N_2964);
or UO_397 (O_397,N_2995,N_2994);
and UO_398 (O_398,N_2996,N_2979);
or UO_399 (O_399,N_2970,N_2961);
or UO_400 (O_400,N_2985,N_2963);
nand UO_401 (O_401,N_2978,N_2950);
nand UO_402 (O_402,N_2999,N_2951);
xnor UO_403 (O_403,N_2987,N_2982);
and UO_404 (O_404,N_2983,N_2953);
and UO_405 (O_405,N_2976,N_2969);
xor UO_406 (O_406,N_2981,N_2954);
or UO_407 (O_407,N_2993,N_2976);
or UO_408 (O_408,N_2950,N_2991);
nor UO_409 (O_409,N_2986,N_2992);
and UO_410 (O_410,N_2953,N_2956);
nor UO_411 (O_411,N_2999,N_2985);
and UO_412 (O_412,N_2980,N_2965);
or UO_413 (O_413,N_2961,N_2962);
and UO_414 (O_414,N_2985,N_2998);
or UO_415 (O_415,N_2988,N_2995);
or UO_416 (O_416,N_2982,N_2981);
nand UO_417 (O_417,N_2964,N_2963);
nor UO_418 (O_418,N_2958,N_2993);
and UO_419 (O_419,N_2960,N_2964);
nor UO_420 (O_420,N_2966,N_2986);
nor UO_421 (O_421,N_2997,N_2992);
nor UO_422 (O_422,N_2986,N_2963);
or UO_423 (O_423,N_2954,N_2972);
or UO_424 (O_424,N_2970,N_2990);
nor UO_425 (O_425,N_2962,N_2983);
xnor UO_426 (O_426,N_2995,N_2954);
and UO_427 (O_427,N_2991,N_2986);
and UO_428 (O_428,N_2973,N_2981);
nor UO_429 (O_429,N_2983,N_2984);
and UO_430 (O_430,N_2979,N_2968);
nor UO_431 (O_431,N_2972,N_2961);
nand UO_432 (O_432,N_2952,N_2995);
nor UO_433 (O_433,N_2953,N_2957);
or UO_434 (O_434,N_2980,N_2951);
and UO_435 (O_435,N_2977,N_2960);
and UO_436 (O_436,N_2970,N_2967);
nor UO_437 (O_437,N_2999,N_2972);
nor UO_438 (O_438,N_2965,N_2999);
and UO_439 (O_439,N_2953,N_2954);
and UO_440 (O_440,N_2971,N_2968);
nor UO_441 (O_441,N_2955,N_2959);
or UO_442 (O_442,N_2972,N_2981);
or UO_443 (O_443,N_2964,N_2956);
nand UO_444 (O_444,N_2972,N_2983);
nor UO_445 (O_445,N_2953,N_2966);
or UO_446 (O_446,N_2984,N_2988);
nor UO_447 (O_447,N_2958,N_2988);
nor UO_448 (O_448,N_2950,N_2961);
or UO_449 (O_449,N_2974,N_2958);
and UO_450 (O_450,N_2981,N_2987);
nand UO_451 (O_451,N_2952,N_2972);
nor UO_452 (O_452,N_2997,N_2958);
and UO_453 (O_453,N_2993,N_2982);
nand UO_454 (O_454,N_2983,N_2965);
nand UO_455 (O_455,N_2989,N_2951);
nand UO_456 (O_456,N_2966,N_2984);
and UO_457 (O_457,N_2998,N_2964);
or UO_458 (O_458,N_2956,N_2970);
and UO_459 (O_459,N_2997,N_2998);
and UO_460 (O_460,N_2965,N_2993);
and UO_461 (O_461,N_2978,N_2995);
nor UO_462 (O_462,N_2953,N_2986);
nand UO_463 (O_463,N_2954,N_2964);
or UO_464 (O_464,N_2986,N_2956);
nor UO_465 (O_465,N_2979,N_2988);
or UO_466 (O_466,N_2995,N_2975);
xor UO_467 (O_467,N_2986,N_2980);
nand UO_468 (O_468,N_2977,N_2992);
and UO_469 (O_469,N_2978,N_2961);
and UO_470 (O_470,N_2974,N_2979);
nor UO_471 (O_471,N_2991,N_2996);
and UO_472 (O_472,N_2971,N_2977);
nor UO_473 (O_473,N_2965,N_2966);
nand UO_474 (O_474,N_2956,N_2984);
xnor UO_475 (O_475,N_2954,N_2987);
xor UO_476 (O_476,N_2960,N_2980);
nand UO_477 (O_477,N_2989,N_2966);
or UO_478 (O_478,N_2979,N_2997);
and UO_479 (O_479,N_2967,N_2950);
nor UO_480 (O_480,N_2967,N_2995);
and UO_481 (O_481,N_2984,N_2968);
or UO_482 (O_482,N_2973,N_2969);
nor UO_483 (O_483,N_2984,N_2973);
or UO_484 (O_484,N_2961,N_2994);
or UO_485 (O_485,N_2956,N_2982);
and UO_486 (O_486,N_2994,N_2998);
or UO_487 (O_487,N_2973,N_2970);
nand UO_488 (O_488,N_2965,N_2986);
nor UO_489 (O_489,N_2969,N_2959);
or UO_490 (O_490,N_2960,N_2974);
or UO_491 (O_491,N_2979,N_2971);
or UO_492 (O_492,N_2974,N_2982);
and UO_493 (O_493,N_2991,N_2972);
and UO_494 (O_494,N_2959,N_2998);
or UO_495 (O_495,N_2955,N_2970);
nor UO_496 (O_496,N_2976,N_2991);
nand UO_497 (O_497,N_2966,N_2950);
or UO_498 (O_498,N_2968,N_2989);
nand UO_499 (O_499,N_2960,N_2972);
endmodule