module basic_750_5000_1000_25_levels_2xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
nor U0 (N_0,In_262,In_120);
and U1 (N_1,In_107,In_260);
nor U2 (N_2,In_466,In_241);
or U3 (N_3,In_292,In_287);
nor U4 (N_4,In_457,In_207);
and U5 (N_5,In_444,In_326);
or U6 (N_6,In_228,In_151);
nand U7 (N_7,In_180,In_42);
nor U8 (N_8,In_740,In_514);
or U9 (N_9,In_523,In_675);
and U10 (N_10,In_177,In_539);
xor U11 (N_11,In_565,In_604);
or U12 (N_12,In_90,In_4);
or U13 (N_13,In_254,In_76);
and U14 (N_14,In_233,In_208);
nor U15 (N_15,In_469,In_306);
and U16 (N_16,In_415,In_141);
nor U17 (N_17,In_737,In_619);
nand U18 (N_18,In_150,In_229);
nor U19 (N_19,In_316,In_723);
and U20 (N_20,In_164,In_673);
and U21 (N_21,In_9,In_621);
or U22 (N_22,In_452,In_303);
and U23 (N_23,In_243,In_531);
nor U24 (N_24,In_548,In_356);
or U25 (N_25,In_77,In_47);
nand U26 (N_26,In_111,In_304);
xor U27 (N_27,In_537,In_580);
or U28 (N_28,In_89,In_209);
or U29 (N_29,In_15,In_330);
nor U30 (N_30,In_124,In_496);
and U31 (N_31,In_202,In_329);
nand U32 (N_32,In_176,In_680);
or U33 (N_33,In_583,In_308);
nor U34 (N_34,In_428,In_590);
or U35 (N_35,In_342,In_648);
nand U36 (N_36,In_335,In_87);
and U37 (N_37,In_392,In_456);
nor U38 (N_38,In_574,In_60);
nand U39 (N_39,In_437,In_106);
or U40 (N_40,In_424,In_67);
or U41 (N_41,In_189,In_88);
or U42 (N_42,In_192,In_512);
nand U43 (N_43,In_480,In_259);
and U44 (N_44,In_190,In_232);
or U45 (N_45,In_423,In_692);
nor U46 (N_46,In_498,In_285);
and U47 (N_47,In_408,In_485);
nand U48 (N_48,In_310,In_614);
or U49 (N_49,In_473,In_462);
nor U50 (N_50,In_579,In_311);
or U51 (N_51,In_645,In_251);
nor U52 (N_52,In_382,In_109);
nor U53 (N_53,In_439,In_519);
and U54 (N_54,In_581,In_373);
and U55 (N_55,In_70,In_244);
or U56 (N_56,In_635,In_299);
nand U57 (N_57,In_79,In_203);
and U58 (N_58,In_718,In_598);
or U59 (N_59,In_295,In_706);
and U60 (N_60,In_484,In_436);
and U61 (N_61,In_429,In_185);
and U62 (N_62,In_724,In_98);
nor U63 (N_63,In_159,In_472);
or U64 (N_64,In_41,In_385);
or U65 (N_65,In_257,In_296);
nor U66 (N_66,In_56,In_334);
nor U67 (N_67,In_602,In_697);
and U68 (N_68,In_488,In_39);
nor U69 (N_69,In_122,In_414);
nor U70 (N_70,In_525,In_301);
and U71 (N_71,In_664,In_395);
xor U72 (N_72,In_250,In_361);
nor U73 (N_73,In_249,In_701);
and U74 (N_74,In_104,In_46);
nand U75 (N_75,In_80,In_520);
nand U76 (N_76,In_119,In_163);
or U77 (N_77,In_671,In_500);
or U78 (N_78,In_704,In_570);
or U79 (N_79,In_169,In_245);
nor U80 (N_80,In_355,In_127);
nand U81 (N_81,In_137,In_234);
nor U82 (N_82,In_551,In_143);
nor U83 (N_83,In_369,In_629);
or U84 (N_84,In_144,In_594);
nor U85 (N_85,In_641,In_650);
nand U86 (N_86,In_401,In_603);
nor U87 (N_87,In_347,In_434);
and U88 (N_88,In_68,In_430);
or U89 (N_89,In_86,In_659);
nor U90 (N_90,In_707,In_665);
or U91 (N_91,In_595,In_688);
nor U92 (N_92,In_588,In_607);
and U93 (N_93,In_610,In_142);
nor U94 (N_94,In_147,In_735);
and U95 (N_95,In_33,In_78);
nor U96 (N_96,In_246,In_64);
or U97 (N_97,In_48,In_231);
or U98 (N_98,In_378,In_383);
nor U99 (N_99,In_562,In_721);
nand U100 (N_100,In_442,In_25);
nor U101 (N_101,In_210,In_327);
nor U102 (N_102,In_678,In_309);
and U103 (N_103,In_427,In_677);
nand U104 (N_104,In_217,In_242);
and U105 (N_105,In_402,In_560);
nor U106 (N_106,In_267,In_503);
or U107 (N_107,In_399,In_256);
and U108 (N_108,In_608,In_59);
and U109 (N_109,In_128,In_420);
nor U110 (N_110,In_546,In_352);
nand U111 (N_111,In_32,In_12);
or U112 (N_112,In_194,In_405);
nand U113 (N_113,In_613,In_129);
nor U114 (N_114,In_685,In_719);
nor U115 (N_115,In_471,In_170);
or U116 (N_116,In_625,In_646);
nor U117 (N_117,In_200,In_341);
or U118 (N_118,In_417,In_84);
or U119 (N_119,In_75,In_85);
or U120 (N_120,In_575,In_74);
or U121 (N_121,In_362,In_467);
and U122 (N_122,In_201,In_175);
nor U123 (N_123,In_722,In_596);
or U124 (N_124,In_669,In_631);
or U125 (N_125,In_172,In_513);
and U126 (N_126,In_130,In_363);
nand U127 (N_127,In_351,In_691);
or U128 (N_128,In_184,In_213);
or U129 (N_129,In_495,In_44);
or U130 (N_130,In_446,In_283);
nand U131 (N_131,In_475,In_632);
nand U132 (N_132,In_505,In_366);
nand U133 (N_133,In_318,In_374);
nor U134 (N_134,In_421,In_291);
or U135 (N_135,In_672,In_284);
nor U136 (N_136,In_689,In_138);
and U137 (N_137,In_367,In_220);
nand U138 (N_138,In_305,In_453);
nand U139 (N_139,In_563,In_100);
nor U140 (N_140,In_344,In_38);
nand U141 (N_141,In_5,In_370);
nand U142 (N_142,In_511,In_276);
nand U143 (N_143,In_624,In_431);
nor U144 (N_144,In_554,In_204);
nand U145 (N_145,In_381,In_620);
nand U146 (N_146,In_440,In_131);
or U147 (N_147,In_435,In_394);
nor U148 (N_148,In_699,In_263);
or U149 (N_149,In_686,In_167);
or U150 (N_150,In_441,In_670);
and U151 (N_151,In_725,In_270);
or U152 (N_152,In_464,In_388);
or U153 (N_153,In_188,In_507);
nor U154 (N_154,In_23,In_69);
nand U155 (N_155,In_123,In_384);
nand U156 (N_156,In_657,In_393);
and U157 (N_157,In_448,In_555);
nand U158 (N_158,In_487,In_668);
and U159 (N_159,In_8,In_57);
or U160 (N_160,In_535,In_418);
or U161 (N_161,In_372,In_509);
nand U162 (N_162,In_696,In_628);
nor U163 (N_163,In_7,In_741);
nor U164 (N_164,In_736,In_586);
xnor U165 (N_165,In_211,In_125);
nand U166 (N_166,In_101,In_536);
or U167 (N_167,In_58,In_656);
nand U168 (N_168,In_593,In_708);
or U169 (N_169,In_528,In_547);
or U170 (N_170,In_340,In_21);
or U171 (N_171,In_447,In_438);
and U172 (N_172,In_389,In_585);
nor U173 (N_173,In_157,In_568);
nand U174 (N_174,In_313,In_684);
nor U175 (N_175,In_542,In_102);
nand U176 (N_176,In_386,In_687);
nor U177 (N_177,In_416,In_526);
and U178 (N_178,In_314,In_333);
or U179 (N_179,In_481,In_567);
nand U180 (N_180,In_636,In_53);
or U181 (N_181,In_223,In_298);
nor U182 (N_182,In_561,In_550);
nand U183 (N_183,In_73,In_622);
nor U184 (N_184,In_40,In_300);
and U185 (N_185,In_746,In_508);
or U186 (N_186,In_281,In_379);
and U187 (N_187,In_571,In_713);
and U188 (N_188,In_156,In_716);
nand U189 (N_189,In_108,In_179);
nand U190 (N_190,In_272,In_403);
or U191 (N_191,In_286,In_694);
nor U192 (N_192,In_654,In_275);
nand U193 (N_193,In_35,In_215);
and U194 (N_194,In_152,In_693);
or U195 (N_195,In_569,In_55);
or U196 (N_196,In_350,In_271);
and U197 (N_197,In_591,In_212);
nor U198 (N_198,In_516,In_703);
nor U199 (N_199,In_196,In_332);
or U200 (N_200,N_5,N_158);
or U201 (N_201,In_726,In_178);
nor U202 (N_202,In_371,In_168);
or U203 (N_203,N_194,In_95);
nand U204 (N_204,In_37,In_651);
or U205 (N_205,In_118,In_126);
nor U206 (N_206,In_490,In_617);
and U207 (N_207,In_627,In_34);
or U208 (N_208,N_69,In_255);
and U209 (N_209,In_155,In_600);
nand U210 (N_210,In_476,In_18);
nor U211 (N_211,In_376,N_109);
and U212 (N_212,In_640,N_101);
or U213 (N_213,In_349,N_18);
nand U214 (N_214,N_187,In_404);
and U215 (N_215,In_99,N_149);
nand U216 (N_216,In_248,In_317);
nand U217 (N_217,In_407,In_454);
or U218 (N_218,In_734,In_307);
nor U219 (N_219,In_2,N_179);
xor U220 (N_220,In_727,In_559);
nand U221 (N_221,N_95,In_748);
and U222 (N_222,In_337,N_104);
or U223 (N_223,In_540,N_52);
nand U224 (N_224,In_52,N_62);
nand U225 (N_225,N_82,In_458);
or U226 (N_226,In_698,In_3);
nand U227 (N_227,In_449,In_410);
and U228 (N_228,N_47,N_71);
or U229 (N_229,In_146,In_577);
and U230 (N_230,In_566,In_552);
or U231 (N_231,N_105,In_470);
nor U232 (N_232,N_181,In_277);
nand U233 (N_233,In_544,N_49);
and U234 (N_234,N_193,In_312);
nand U235 (N_235,N_88,N_146);
nor U236 (N_236,In_162,N_30);
and U237 (N_237,N_173,In_236);
nand U238 (N_238,In_348,In_279);
nor U239 (N_239,In_160,In_463);
and U240 (N_240,In_510,In_486);
nand U241 (N_241,N_112,In_91);
nor U242 (N_242,In_413,N_119);
and U243 (N_243,N_29,N_120);
or U244 (N_244,In_63,In_238);
or U245 (N_245,In_132,N_137);
nand U246 (N_246,In_529,N_170);
or U247 (N_247,In_338,N_57);
nand U248 (N_248,N_19,In_601);
nor U249 (N_249,In_247,In_216);
and U250 (N_250,In_611,In_532);
xnor U251 (N_251,N_167,N_97);
nor U252 (N_252,In_663,N_40);
nor U253 (N_253,In_166,N_99);
nor U254 (N_254,In_50,In_564);
and U255 (N_255,In_158,In_666);
and U256 (N_256,N_183,In_320);
or U257 (N_257,In_92,N_38);
and U258 (N_258,N_157,In_135);
nand U259 (N_259,In_538,In_682);
or U260 (N_260,N_3,In_116);
and U261 (N_261,In_97,N_154);
nor U262 (N_262,In_578,In_661);
nor U263 (N_263,In_465,In_460);
and U264 (N_264,In_710,N_46);
nand U265 (N_265,In_700,In_433);
nand U266 (N_266,In_148,In_743);
and U267 (N_267,In_115,In_261);
and U268 (N_268,In_482,N_190);
nand U269 (N_269,N_60,In_183);
nand U270 (N_270,In_679,N_16);
or U271 (N_271,In_199,In_584);
nor U272 (N_272,N_180,N_26);
nor U273 (N_273,In_319,In_409);
and U274 (N_274,N_153,In_589);
nand U275 (N_275,N_93,N_68);
nand U276 (N_276,In_702,In_280);
nor U277 (N_277,N_116,In_556);
or U278 (N_278,In_27,In_732);
nor U279 (N_279,In_149,In_705);
nor U280 (N_280,In_31,N_117);
or U281 (N_281,In_278,In_489);
nor U282 (N_282,N_192,In_461);
or U283 (N_283,In_674,N_44);
nand U284 (N_284,N_17,In_174);
or U285 (N_285,N_185,In_226);
nor U286 (N_286,N_2,In_182);
and U287 (N_287,N_25,N_21);
nand U288 (N_288,N_169,N_10);
nor U289 (N_289,In_154,In_747);
nor U290 (N_290,In_96,In_749);
nand U291 (N_291,In_218,In_478);
nand U292 (N_292,In_266,In_10);
xnor U293 (N_293,N_125,In_504);
or U294 (N_294,In_524,In_61);
nand U295 (N_295,In_597,In_642);
nor U296 (N_296,N_160,In_558);
or U297 (N_297,N_86,N_0);
nor U298 (N_298,N_20,In_695);
nor U299 (N_299,In_325,In_221);
nor U300 (N_300,In_43,N_118);
nor U301 (N_301,In_345,In_274);
nand U302 (N_302,In_419,In_499);
or U303 (N_303,In_653,In_136);
nor U304 (N_304,In_28,N_84);
and U305 (N_305,In_26,N_163);
nand U306 (N_306,In_81,In_745);
and U307 (N_307,N_196,In_521);
nand U308 (N_308,In_29,In_171);
nand U309 (N_309,N_165,In_549);
nor U310 (N_310,In_609,In_422);
nor U311 (N_311,N_7,N_91);
nor U312 (N_312,N_184,In_667);
nor U313 (N_313,In_406,N_134);
nor U314 (N_314,N_136,In_13);
and U315 (N_315,In_375,In_599);
and U316 (N_316,N_177,In_515);
or U317 (N_317,In_451,In_545);
nand U318 (N_318,N_58,N_115);
nor U319 (N_319,N_130,In_359);
nand U320 (N_320,In_66,N_36);
or U321 (N_321,N_43,N_11);
nor U322 (N_322,N_141,In_728);
or U323 (N_323,In_239,In_396);
and U324 (N_324,N_51,In_357);
xnor U325 (N_325,In_506,In_206);
or U326 (N_326,In_527,In_94);
and U327 (N_327,N_63,In_36);
or U328 (N_328,N_128,In_293);
nor U329 (N_329,N_89,N_50);
or U330 (N_330,N_140,In_214);
nand U331 (N_331,N_188,N_144);
or U332 (N_332,In_541,In_638);
nand U333 (N_333,In_518,In_83);
nand U334 (N_334,In_302,In_230);
and U335 (N_335,In_22,In_6);
nand U336 (N_336,In_288,In_623);
or U337 (N_337,In_139,In_324);
or U338 (N_338,N_122,N_162);
or U339 (N_339,In_105,N_23);
nand U340 (N_340,N_151,In_165);
or U341 (N_341,In_187,In_644);
or U342 (N_342,N_176,N_110);
or U343 (N_343,N_55,In_533);
or U344 (N_344,In_153,In_445);
and U345 (N_345,N_67,N_108);
nor U346 (N_346,N_175,In_522);
and U347 (N_347,N_113,In_543);
nand U348 (N_348,N_77,In_606);
and U349 (N_349,N_90,N_54);
or U350 (N_350,In_346,In_494);
and U351 (N_351,N_102,N_59);
nand U352 (N_352,In_553,In_683);
and U353 (N_353,In_117,N_189);
nor U354 (N_354,N_131,N_135);
and U355 (N_355,In_240,In_634);
or U356 (N_356,In_432,In_572);
or U357 (N_357,N_138,In_258);
or U358 (N_358,In_711,In_502);
or U359 (N_359,In_328,In_615);
nand U360 (N_360,In_681,In_455);
or U361 (N_361,In_398,N_197);
nand U362 (N_362,In_733,N_64);
and U363 (N_363,In_17,In_637);
nand U364 (N_364,N_107,In_652);
nand U365 (N_365,In_181,In_198);
or U366 (N_366,In_391,In_323);
nor U367 (N_367,N_74,N_87);
or U368 (N_368,N_80,N_139);
nor U369 (N_369,In_647,In_612);
nor U370 (N_370,In_658,In_690);
and U371 (N_371,N_53,In_65);
nor U372 (N_372,N_37,In_720);
nand U373 (N_373,N_83,In_744);
nand U374 (N_374,N_34,In_24);
or U375 (N_375,In_365,N_4);
nor U376 (N_376,In_517,N_174);
nor U377 (N_377,In_195,N_15);
nor U378 (N_378,In_353,N_72);
nand U379 (N_379,N_195,N_155);
nand U380 (N_380,In_268,N_32);
or U381 (N_381,In_331,In_315);
nand U382 (N_382,In_425,In_224);
and U383 (N_383,In_269,In_265);
nor U384 (N_384,In_161,In_14);
or U385 (N_385,In_739,In_573);
nor U386 (N_386,N_33,In_714);
and U387 (N_387,In_110,In_364);
or U388 (N_388,N_126,In_479);
and U389 (N_389,In_397,In_20);
or U390 (N_390,N_78,In_173);
nand U391 (N_391,In_649,In_11);
and U392 (N_392,In_358,N_79);
nor U393 (N_393,N_100,N_22);
and U394 (N_394,In_121,In_93);
nand U395 (N_395,In_717,In_191);
nand U396 (N_396,In_491,N_75);
and U397 (N_397,N_98,N_27);
and U398 (N_398,N_41,N_31);
or U399 (N_399,In_322,In_459);
nand U400 (N_400,In_377,N_392);
and U401 (N_401,N_326,In_443);
nor U402 (N_402,N_256,N_230);
or U403 (N_403,N_123,N_229);
nand U404 (N_404,In_709,N_209);
nand U405 (N_405,N_311,N_343);
or U406 (N_406,N_270,In_237);
nand U407 (N_407,N_85,In_219);
or U408 (N_408,N_312,N_309);
and U409 (N_409,In_72,N_73);
and U410 (N_410,N_248,In_273);
nor U411 (N_411,N_275,N_293);
nand U412 (N_412,N_226,N_210);
nor U413 (N_413,N_356,N_334);
nor U414 (N_414,N_299,N_222);
nand U415 (N_415,In_294,N_106);
nand U416 (N_416,In_71,N_289);
or U417 (N_417,N_96,N_280);
and U418 (N_418,N_370,In_412);
nor U419 (N_419,N_368,N_365);
nand U420 (N_420,In_738,N_220);
and U421 (N_421,N_267,N_243);
nor U422 (N_422,N_66,N_316);
and U423 (N_423,In_643,N_357);
nand U424 (N_424,N_381,N_327);
and U425 (N_425,In_193,In_51);
and U426 (N_426,N_81,N_379);
nor U427 (N_427,N_344,N_200);
or U428 (N_428,N_352,N_254);
and U429 (N_429,N_202,In_82);
and U430 (N_430,N_234,In_354);
or U431 (N_431,In_477,N_264);
and U432 (N_432,N_318,N_150);
and U433 (N_433,N_164,In_587);
xnor U434 (N_434,N_224,N_304);
or U435 (N_435,N_1,In_343);
nand U436 (N_436,In_715,N_186);
and U437 (N_437,N_147,N_345);
and U438 (N_438,N_212,N_262);
and U439 (N_439,N_127,N_132);
and U440 (N_440,In_390,In_222);
or U441 (N_441,N_272,In_450);
and U442 (N_442,N_76,In_186);
nor U443 (N_443,N_333,N_305);
xnor U444 (N_444,N_394,N_295);
nand U445 (N_445,In_235,N_285);
nand U446 (N_446,In_112,N_143);
nand U447 (N_447,N_263,N_341);
nor U448 (N_448,N_148,N_395);
or U449 (N_449,In_626,N_145);
and U450 (N_450,In_712,In_290);
xor U451 (N_451,In_16,N_258);
or U452 (N_452,In_582,N_213);
nor U453 (N_453,N_353,N_322);
nand U454 (N_454,N_278,N_70);
or U455 (N_455,N_279,N_214);
nand U456 (N_456,N_282,N_315);
or U457 (N_457,In_134,N_133);
or U458 (N_458,N_359,N_240);
or U459 (N_459,N_351,In_19);
nand U460 (N_460,N_39,N_245);
or U461 (N_461,N_288,N_332);
nand U462 (N_462,In_145,N_389);
or U463 (N_463,N_244,N_265);
or U464 (N_464,N_361,N_355);
nor U465 (N_465,In_339,In_205);
nand U466 (N_466,N_374,N_297);
nor U467 (N_467,In_530,N_391);
or U468 (N_468,N_317,N_301);
and U469 (N_469,N_324,In_426);
and U470 (N_470,In_468,N_191);
and U471 (N_471,N_261,N_65);
nor U472 (N_472,In_227,N_178);
and U473 (N_473,N_382,N_387);
nand U474 (N_474,In_113,N_114);
and U475 (N_475,In_45,N_199);
nor U476 (N_476,N_383,In_103);
or U477 (N_477,N_372,N_390);
nor U478 (N_478,N_12,In_630);
and U479 (N_479,N_48,N_371);
or U480 (N_480,N_94,N_266);
nor U481 (N_481,N_377,N_384);
or U482 (N_482,N_269,In_534);
xor U483 (N_483,N_228,N_227);
and U484 (N_484,In_264,N_349);
nor U485 (N_485,N_225,In_576);
nor U486 (N_486,N_292,N_166);
or U487 (N_487,N_239,In_639);
nand U488 (N_488,In_592,N_253);
or U489 (N_489,N_217,N_338);
or U490 (N_490,In_501,N_367);
and U491 (N_491,N_242,N_283);
nor U492 (N_492,N_323,N_376);
and U493 (N_493,In_380,N_393);
or U494 (N_494,N_346,N_201);
and U495 (N_495,In_114,N_249);
or U496 (N_496,In_729,N_364);
nand U497 (N_497,N_250,N_287);
and U498 (N_498,N_260,N_232);
nand U499 (N_499,In_225,N_362);
and U500 (N_500,In_742,In_676);
and U501 (N_501,N_276,In_62);
and U502 (N_502,N_198,N_325);
xnor U503 (N_503,N_373,N_14);
nand U504 (N_504,In_297,N_378);
nor U505 (N_505,In_662,N_255);
and U506 (N_506,N_223,N_121);
or U507 (N_507,N_366,N_340);
nor U508 (N_508,In_633,N_219);
nor U509 (N_509,In_387,N_360);
nor U510 (N_510,In_140,In_321);
nand U511 (N_511,N_161,N_296);
and U512 (N_512,N_237,N_124);
or U513 (N_513,N_271,N_291);
or U514 (N_514,In_360,In_133);
nand U515 (N_515,N_45,In_497);
and U516 (N_516,In_474,N_168);
and U517 (N_517,N_24,N_328);
or U518 (N_518,N_302,N_216);
nor U519 (N_519,N_331,N_218);
nand U520 (N_520,N_208,N_342);
or U521 (N_521,In_368,N_286);
or U522 (N_522,In_616,N_336);
or U523 (N_523,N_313,N_281);
nand U524 (N_524,N_306,N_252);
and U525 (N_525,In_49,N_204);
and U526 (N_526,In_1,In_483);
or U527 (N_527,In_30,In_336);
xor U528 (N_528,In_54,N_369);
nand U529 (N_529,N_129,N_111);
and U530 (N_530,N_35,In_253);
or U531 (N_531,N_156,N_339);
nor U532 (N_532,N_375,N_103);
nor U533 (N_533,N_56,N_348);
nand U534 (N_534,N_236,N_330);
and U535 (N_535,In_655,N_159);
and U536 (N_536,In_492,N_203);
nand U537 (N_537,N_257,N_61);
nor U538 (N_538,N_284,In_730);
and U539 (N_539,N_172,N_300);
nand U540 (N_540,N_206,N_337);
or U541 (N_541,N_215,N_380);
nand U542 (N_542,N_247,N_319);
or U543 (N_543,In_605,In_197);
nand U544 (N_544,N_251,N_335);
nand U545 (N_545,N_221,In_0);
nand U546 (N_546,N_358,N_231);
or U547 (N_547,N_9,In_618);
or U548 (N_548,N_246,In_400);
nor U549 (N_549,In_557,N_350);
and U550 (N_550,N_6,In_282);
nand U551 (N_551,N_308,N_385);
and U552 (N_552,N_303,N_310);
nand U553 (N_553,N_28,N_347);
or U554 (N_554,In_660,N_290);
or U555 (N_555,N_314,N_354);
and U556 (N_556,N_152,In_493);
nor U557 (N_557,N_207,N_388);
or U558 (N_558,N_329,N_321);
nor U559 (N_559,N_398,N_274);
nand U560 (N_560,N_307,N_241);
and U561 (N_561,N_396,N_259);
nand U562 (N_562,N_233,In_252);
and U563 (N_563,N_8,N_399);
nor U564 (N_564,N_273,N_171);
nand U565 (N_565,N_142,In_289);
xnor U566 (N_566,N_294,N_13);
nand U567 (N_567,N_397,N_205);
nor U568 (N_568,N_386,N_92);
or U569 (N_569,N_363,N_182);
nor U570 (N_570,N_238,N_298);
and U571 (N_571,In_411,N_42);
and U572 (N_572,N_277,N_320);
and U573 (N_573,N_211,N_268);
and U574 (N_574,N_235,In_731);
nand U575 (N_575,N_161,In_54);
nand U576 (N_576,N_252,In_530);
or U577 (N_577,N_392,N_307);
and U578 (N_578,In_45,N_235);
nor U579 (N_579,In_140,N_232);
or U580 (N_580,N_147,N_305);
or U581 (N_581,N_250,In_712);
nand U582 (N_582,N_65,N_269);
nand U583 (N_583,In_660,N_148);
nand U584 (N_584,In_639,In_450);
nor U585 (N_585,In_227,N_363);
and U586 (N_586,N_205,N_129);
and U587 (N_587,N_242,N_227);
nand U588 (N_588,N_313,N_303);
or U589 (N_589,N_369,N_247);
nand U590 (N_590,N_191,N_256);
nor U591 (N_591,N_216,N_182);
nand U592 (N_592,N_6,N_85);
or U593 (N_593,In_235,N_133);
and U594 (N_594,N_66,N_237);
nor U595 (N_595,N_243,In_222);
nor U596 (N_596,N_315,N_306);
nand U597 (N_597,In_103,N_45);
or U598 (N_598,N_150,N_208);
nor U599 (N_599,In_477,N_280);
nor U600 (N_600,N_409,N_425);
or U601 (N_601,N_487,N_526);
nor U602 (N_602,N_552,N_470);
and U603 (N_603,N_560,N_597);
nand U604 (N_604,N_571,N_501);
nand U605 (N_605,N_563,N_458);
nand U606 (N_606,N_553,N_440);
nor U607 (N_607,N_536,N_407);
nand U608 (N_608,N_576,N_404);
and U609 (N_609,N_585,N_406);
and U610 (N_610,N_413,N_517);
nand U611 (N_611,N_558,N_494);
or U612 (N_612,N_543,N_463);
or U613 (N_613,N_528,N_562);
nor U614 (N_614,N_586,N_532);
nand U615 (N_615,N_461,N_491);
and U616 (N_616,N_550,N_596);
nor U617 (N_617,N_531,N_431);
or U618 (N_618,N_509,N_414);
or U619 (N_619,N_444,N_497);
or U620 (N_620,N_466,N_492);
and U621 (N_621,N_599,N_498);
and U622 (N_622,N_513,N_419);
nand U623 (N_623,N_515,N_555);
and U624 (N_624,N_478,N_418);
nand U625 (N_625,N_474,N_544);
nand U626 (N_626,N_556,N_589);
and U627 (N_627,N_403,N_401);
nand U628 (N_628,N_575,N_462);
or U629 (N_629,N_546,N_460);
nand U630 (N_630,N_545,N_493);
nor U631 (N_631,N_446,N_527);
nor U632 (N_632,N_496,N_443);
nand U633 (N_633,N_566,N_479);
and U634 (N_634,N_472,N_438);
nor U635 (N_635,N_452,N_583);
nor U636 (N_636,N_450,N_584);
or U637 (N_637,N_572,N_426);
or U638 (N_638,N_529,N_468);
nor U639 (N_639,N_590,N_489);
nor U640 (N_640,N_417,N_416);
and U641 (N_641,N_511,N_453);
nand U642 (N_642,N_408,N_410);
nand U643 (N_643,N_594,N_445);
and U644 (N_644,N_588,N_433);
nor U645 (N_645,N_565,N_402);
or U646 (N_646,N_522,N_551);
nor U647 (N_647,N_534,N_483);
or U648 (N_648,N_424,N_557);
nor U649 (N_649,N_471,N_535);
or U650 (N_650,N_580,N_554);
nand U651 (N_651,N_400,N_537);
nand U652 (N_652,N_533,N_422);
or U653 (N_653,N_423,N_539);
and U654 (N_654,N_598,N_569);
nor U655 (N_655,N_541,N_579);
nor U656 (N_656,N_481,N_508);
nor U657 (N_657,N_574,N_499);
and U658 (N_658,N_495,N_430);
nand U659 (N_659,N_432,N_475);
nand U660 (N_660,N_591,N_427);
nor U661 (N_661,N_577,N_485);
nand U662 (N_662,N_568,N_503);
nand U663 (N_663,N_480,N_454);
or U664 (N_664,N_435,N_473);
nand U665 (N_665,N_459,N_507);
or U666 (N_666,N_587,N_510);
nand U667 (N_667,N_488,N_504);
nand U668 (N_668,N_500,N_415);
or U669 (N_669,N_411,N_519);
nand U670 (N_670,N_484,N_429);
nor U671 (N_671,N_592,N_434);
nor U672 (N_672,N_567,N_582);
nor U673 (N_673,N_412,N_441);
nor U674 (N_674,N_524,N_578);
nand U675 (N_675,N_447,N_548);
and U676 (N_676,N_520,N_467);
and U677 (N_677,N_559,N_437);
and U678 (N_678,N_439,N_549);
and U679 (N_679,N_564,N_523);
nand U680 (N_680,N_540,N_516);
nand U681 (N_681,N_573,N_542);
nand U682 (N_682,N_570,N_538);
or U683 (N_683,N_451,N_464);
and U684 (N_684,N_506,N_561);
and U685 (N_685,N_486,N_436);
and U686 (N_686,N_490,N_469);
nor U687 (N_687,N_512,N_420);
nor U688 (N_688,N_442,N_593);
nor U689 (N_689,N_547,N_581);
or U690 (N_690,N_476,N_518);
xor U691 (N_691,N_421,N_521);
nor U692 (N_692,N_502,N_456);
nor U693 (N_693,N_405,N_514);
or U694 (N_694,N_428,N_457);
xnor U695 (N_695,N_505,N_482);
or U696 (N_696,N_448,N_530);
or U697 (N_697,N_525,N_449);
nor U698 (N_698,N_595,N_477);
nor U699 (N_699,N_465,N_455);
or U700 (N_700,N_576,N_475);
and U701 (N_701,N_564,N_538);
nand U702 (N_702,N_440,N_492);
or U703 (N_703,N_423,N_571);
or U704 (N_704,N_508,N_437);
nand U705 (N_705,N_568,N_523);
or U706 (N_706,N_412,N_575);
or U707 (N_707,N_589,N_554);
or U708 (N_708,N_489,N_595);
nand U709 (N_709,N_533,N_427);
or U710 (N_710,N_585,N_516);
and U711 (N_711,N_459,N_490);
nand U712 (N_712,N_564,N_566);
or U713 (N_713,N_499,N_444);
nor U714 (N_714,N_456,N_552);
and U715 (N_715,N_473,N_568);
and U716 (N_716,N_466,N_427);
nor U717 (N_717,N_487,N_462);
nand U718 (N_718,N_445,N_478);
nor U719 (N_719,N_575,N_556);
nor U720 (N_720,N_503,N_413);
nand U721 (N_721,N_401,N_495);
or U722 (N_722,N_411,N_462);
nor U723 (N_723,N_500,N_481);
nand U724 (N_724,N_432,N_405);
or U725 (N_725,N_596,N_506);
nor U726 (N_726,N_402,N_594);
and U727 (N_727,N_436,N_442);
nand U728 (N_728,N_416,N_463);
nand U729 (N_729,N_408,N_466);
or U730 (N_730,N_563,N_554);
xnor U731 (N_731,N_522,N_464);
nand U732 (N_732,N_550,N_440);
xnor U733 (N_733,N_578,N_433);
nor U734 (N_734,N_510,N_414);
nor U735 (N_735,N_490,N_442);
and U736 (N_736,N_553,N_421);
or U737 (N_737,N_555,N_440);
xnor U738 (N_738,N_511,N_484);
nand U739 (N_739,N_496,N_434);
nand U740 (N_740,N_487,N_488);
nand U741 (N_741,N_452,N_447);
and U742 (N_742,N_592,N_553);
or U743 (N_743,N_402,N_451);
nand U744 (N_744,N_516,N_464);
nand U745 (N_745,N_514,N_431);
nand U746 (N_746,N_452,N_435);
nand U747 (N_747,N_599,N_566);
or U748 (N_748,N_580,N_471);
xor U749 (N_749,N_551,N_582);
and U750 (N_750,N_519,N_586);
and U751 (N_751,N_502,N_594);
and U752 (N_752,N_574,N_506);
or U753 (N_753,N_571,N_459);
and U754 (N_754,N_433,N_574);
nand U755 (N_755,N_471,N_443);
or U756 (N_756,N_479,N_477);
nor U757 (N_757,N_578,N_561);
nor U758 (N_758,N_512,N_573);
or U759 (N_759,N_424,N_586);
nor U760 (N_760,N_483,N_420);
nor U761 (N_761,N_471,N_502);
or U762 (N_762,N_495,N_473);
or U763 (N_763,N_591,N_540);
nand U764 (N_764,N_468,N_514);
or U765 (N_765,N_572,N_457);
or U766 (N_766,N_407,N_420);
nand U767 (N_767,N_434,N_505);
nor U768 (N_768,N_584,N_405);
or U769 (N_769,N_443,N_512);
nor U770 (N_770,N_421,N_585);
nor U771 (N_771,N_598,N_445);
nor U772 (N_772,N_598,N_543);
and U773 (N_773,N_467,N_547);
or U774 (N_774,N_599,N_545);
nor U775 (N_775,N_407,N_571);
and U776 (N_776,N_513,N_422);
nor U777 (N_777,N_414,N_438);
or U778 (N_778,N_498,N_518);
nor U779 (N_779,N_473,N_406);
nor U780 (N_780,N_456,N_477);
and U781 (N_781,N_455,N_432);
nand U782 (N_782,N_556,N_569);
or U783 (N_783,N_409,N_441);
nand U784 (N_784,N_417,N_516);
nand U785 (N_785,N_405,N_449);
and U786 (N_786,N_587,N_488);
and U787 (N_787,N_410,N_570);
and U788 (N_788,N_590,N_417);
nand U789 (N_789,N_461,N_536);
nand U790 (N_790,N_501,N_431);
nor U791 (N_791,N_499,N_570);
and U792 (N_792,N_466,N_414);
nor U793 (N_793,N_511,N_529);
and U794 (N_794,N_439,N_500);
or U795 (N_795,N_406,N_574);
nor U796 (N_796,N_498,N_542);
nand U797 (N_797,N_426,N_500);
and U798 (N_798,N_538,N_519);
xnor U799 (N_799,N_403,N_594);
and U800 (N_800,N_790,N_701);
or U801 (N_801,N_631,N_721);
or U802 (N_802,N_731,N_666);
nor U803 (N_803,N_604,N_773);
nor U804 (N_804,N_644,N_730);
and U805 (N_805,N_671,N_766);
and U806 (N_806,N_752,N_610);
nand U807 (N_807,N_776,N_613);
nor U808 (N_808,N_706,N_694);
nor U809 (N_809,N_625,N_749);
or U810 (N_810,N_677,N_712);
or U811 (N_811,N_637,N_692);
or U812 (N_812,N_630,N_643);
and U813 (N_813,N_709,N_662);
nor U814 (N_814,N_645,N_735);
or U815 (N_815,N_789,N_663);
and U816 (N_816,N_769,N_668);
and U817 (N_817,N_601,N_682);
nor U818 (N_818,N_711,N_628);
and U819 (N_819,N_750,N_695);
nor U820 (N_820,N_762,N_702);
nor U821 (N_821,N_633,N_777);
nand U822 (N_822,N_618,N_765);
or U823 (N_823,N_683,N_659);
and U824 (N_824,N_600,N_640);
nand U825 (N_825,N_715,N_719);
and U826 (N_826,N_723,N_727);
and U827 (N_827,N_665,N_664);
or U828 (N_828,N_737,N_717);
and U829 (N_829,N_639,N_676);
or U830 (N_830,N_713,N_669);
or U831 (N_831,N_748,N_626);
nor U832 (N_832,N_674,N_747);
nand U833 (N_833,N_673,N_722);
nand U834 (N_834,N_739,N_621);
xor U835 (N_835,N_745,N_693);
nand U836 (N_836,N_679,N_704);
nor U837 (N_837,N_767,N_661);
or U838 (N_838,N_609,N_688);
nand U839 (N_839,N_636,N_696);
nand U840 (N_840,N_622,N_726);
nor U841 (N_841,N_611,N_738);
nand U842 (N_842,N_623,N_606);
or U843 (N_843,N_728,N_753);
or U844 (N_844,N_798,N_697);
xnor U845 (N_845,N_655,N_672);
nor U846 (N_846,N_732,N_689);
or U847 (N_847,N_699,N_710);
and U848 (N_848,N_714,N_743);
and U849 (N_849,N_660,N_729);
nor U850 (N_850,N_770,N_651);
and U851 (N_851,N_678,N_687);
and U852 (N_852,N_707,N_755);
nand U853 (N_853,N_741,N_703);
nor U854 (N_854,N_646,N_705);
and U855 (N_855,N_657,N_638);
xor U856 (N_856,N_634,N_768);
nand U857 (N_857,N_751,N_720);
and U858 (N_858,N_733,N_691);
or U859 (N_859,N_736,N_744);
nor U860 (N_860,N_761,N_700);
nand U861 (N_861,N_656,N_781);
and U862 (N_862,N_740,N_650);
nor U863 (N_863,N_795,N_775);
nor U864 (N_864,N_785,N_793);
and U865 (N_865,N_724,N_686);
nand U866 (N_866,N_652,N_763);
nand U867 (N_867,N_734,N_614);
or U868 (N_868,N_782,N_642);
nand U869 (N_869,N_786,N_616);
nand U870 (N_870,N_607,N_635);
nand U871 (N_871,N_780,N_675);
nor U872 (N_872,N_718,N_648);
and U873 (N_873,N_603,N_615);
nor U874 (N_874,N_772,N_757);
or U875 (N_875,N_799,N_779);
or U876 (N_876,N_629,N_708);
and U877 (N_877,N_788,N_760);
and U878 (N_878,N_641,N_754);
nand U879 (N_879,N_619,N_758);
or U880 (N_880,N_620,N_756);
or U881 (N_881,N_647,N_791);
and U882 (N_882,N_667,N_602);
and U883 (N_883,N_684,N_716);
nor U884 (N_884,N_796,N_725);
nor U885 (N_885,N_690,N_759);
or U886 (N_886,N_627,N_612);
or U887 (N_887,N_605,N_624);
or U888 (N_888,N_654,N_658);
nand U889 (N_889,N_792,N_653);
or U890 (N_890,N_787,N_746);
nor U891 (N_891,N_670,N_797);
or U892 (N_892,N_794,N_783);
or U893 (N_893,N_784,N_617);
and U894 (N_894,N_698,N_632);
nor U895 (N_895,N_685,N_608);
or U896 (N_896,N_742,N_764);
nor U897 (N_897,N_774,N_649);
nand U898 (N_898,N_771,N_681);
nor U899 (N_899,N_778,N_680);
nand U900 (N_900,N_784,N_666);
nor U901 (N_901,N_643,N_687);
nand U902 (N_902,N_604,N_741);
nand U903 (N_903,N_741,N_796);
nor U904 (N_904,N_714,N_748);
nand U905 (N_905,N_775,N_664);
or U906 (N_906,N_644,N_688);
xor U907 (N_907,N_676,N_704);
nor U908 (N_908,N_704,N_726);
nand U909 (N_909,N_789,N_738);
nor U910 (N_910,N_609,N_772);
nor U911 (N_911,N_753,N_699);
xor U912 (N_912,N_665,N_742);
nor U913 (N_913,N_647,N_680);
or U914 (N_914,N_743,N_678);
nor U915 (N_915,N_739,N_607);
nand U916 (N_916,N_643,N_609);
and U917 (N_917,N_763,N_752);
and U918 (N_918,N_643,N_738);
nand U919 (N_919,N_794,N_743);
or U920 (N_920,N_789,N_788);
or U921 (N_921,N_771,N_619);
nor U922 (N_922,N_651,N_752);
nand U923 (N_923,N_682,N_799);
and U924 (N_924,N_775,N_673);
and U925 (N_925,N_650,N_709);
and U926 (N_926,N_610,N_688);
and U927 (N_927,N_773,N_694);
or U928 (N_928,N_607,N_772);
or U929 (N_929,N_776,N_717);
nor U930 (N_930,N_785,N_719);
or U931 (N_931,N_721,N_799);
and U932 (N_932,N_730,N_671);
nand U933 (N_933,N_615,N_612);
or U934 (N_934,N_777,N_656);
and U935 (N_935,N_657,N_729);
and U936 (N_936,N_669,N_792);
xnor U937 (N_937,N_648,N_695);
or U938 (N_938,N_682,N_743);
nand U939 (N_939,N_759,N_732);
nor U940 (N_940,N_648,N_745);
nor U941 (N_941,N_737,N_747);
and U942 (N_942,N_799,N_768);
nor U943 (N_943,N_763,N_728);
or U944 (N_944,N_687,N_662);
or U945 (N_945,N_746,N_604);
and U946 (N_946,N_654,N_643);
or U947 (N_947,N_683,N_682);
nand U948 (N_948,N_638,N_602);
or U949 (N_949,N_617,N_743);
nand U950 (N_950,N_721,N_621);
or U951 (N_951,N_685,N_691);
nor U952 (N_952,N_752,N_769);
and U953 (N_953,N_734,N_795);
nor U954 (N_954,N_746,N_717);
or U955 (N_955,N_614,N_672);
or U956 (N_956,N_666,N_619);
or U957 (N_957,N_702,N_655);
nor U958 (N_958,N_709,N_731);
and U959 (N_959,N_760,N_685);
nand U960 (N_960,N_741,N_772);
nor U961 (N_961,N_736,N_689);
nor U962 (N_962,N_658,N_717);
nor U963 (N_963,N_600,N_767);
and U964 (N_964,N_712,N_742);
and U965 (N_965,N_616,N_610);
nor U966 (N_966,N_768,N_661);
and U967 (N_967,N_699,N_654);
nor U968 (N_968,N_628,N_605);
nor U969 (N_969,N_745,N_706);
or U970 (N_970,N_761,N_672);
and U971 (N_971,N_712,N_700);
or U972 (N_972,N_717,N_602);
and U973 (N_973,N_690,N_715);
nor U974 (N_974,N_611,N_799);
and U975 (N_975,N_775,N_698);
or U976 (N_976,N_611,N_691);
or U977 (N_977,N_620,N_657);
nand U978 (N_978,N_696,N_629);
and U979 (N_979,N_729,N_626);
or U980 (N_980,N_707,N_652);
nand U981 (N_981,N_767,N_716);
nand U982 (N_982,N_611,N_613);
or U983 (N_983,N_792,N_708);
or U984 (N_984,N_680,N_756);
or U985 (N_985,N_720,N_622);
nor U986 (N_986,N_654,N_690);
or U987 (N_987,N_730,N_717);
or U988 (N_988,N_663,N_705);
nor U989 (N_989,N_620,N_676);
or U990 (N_990,N_771,N_695);
and U991 (N_991,N_740,N_782);
nor U992 (N_992,N_642,N_797);
nand U993 (N_993,N_651,N_686);
nand U994 (N_994,N_658,N_650);
or U995 (N_995,N_754,N_605);
and U996 (N_996,N_644,N_782);
or U997 (N_997,N_782,N_620);
and U998 (N_998,N_675,N_656);
nand U999 (N_999,N_646,N_687);
nand U1000 (N_1000,N_824,N_845);
nand U1001 (N_1001,N_882,N_800);
nand U1002 (N_1002,N_958,N_982);
nor U1003 (N_1003,N_962,N_840);
and U1004 (N_1004,N_880,N_996);
and U1005 (N_1005,N_825,N_842);
or U1006 (N_1006,N_969,N_852);
or U1007 (N_1007,N_837,N_858);
and U1008 (N_1008,N_972,N_967);
nand U1009 (N_1009,N_817,N_892);
or U1010 (N_1010,N_853,N_873);
nand U1011 (N_1011,N_823,N_989);
nor U1012 (N_1012,N_843,N_801);
or U1013 (N_1013,N_862,N_975);
or U1014 (N_1014,N_928,N_864);
nor U1015 (N_1015,N_894,N_942);
nor U1016 (N_1016,N_919,N_805);
nor U1017 (N_1017,N_953,N_872);
or U1018 (N_1018,N_907,N_991);
or U1019 (N_1019,N_951,N_970);
nor U1020 (N_1020,N_878,N_946);
nor U1021 (N_1021,N_956,N_994);
or U1022 (N_1022,N_890,N_984);
and U1023 (N_1023,N_847,N_997);
or U1024 (N_1024,N_939,N_877);
or U1025 (N_1025,N_810,N_911);
nand U1026 (N_1026,N_941,N_808);
and U1027 (N_1027,N_908,N_979);
nand U1028 (N_1028,N_833,N_871);
and U1029 (N_1029,N_902,N_895);
and U1030 (N_1030,N_978,N_983);
nand U1031 (N_1031,N_802,N_959);
and U1032 (N_1032,N_990,N_883);
nand U1033 (N_1033,N_900,N_812);
nor U1034 (N_1034,N_934,N_950);
nor U1035 (N_1035,N_992,N_857);
nor U1036 (N_1036,N_955,N_917);
and U1037 (N_1037,N_910,N_960);
or U1038 (N_1038,N_881,N_828);
nand U1039 (N_1039,N_988,N_918);
or U1040 (N_1040,N_809,N_807);
or U1041 (N_1041,N_844,N_803);
nand U1042 (N_1042,N_947,N_846);
nor U1043 (N_1043,N_806,N_903);
or U1044 (N_1044,N_921,N_974);
nor U1045 (N_1045,N_826,N_897);
or U1046 (N_1046,N_865,N_986);
or U1047 (N_1047,N_924,N_944);
or U1048 (N_1048,N_977,N_855);
nand U1049 (N_1049,N_898,N_856);
nor U1050 (N_1050,N_961,N_906);
or U1051 (N_1051,N_981,N_887);
and U1052 (N_1052,N_987,N_896);
xnor U1053 (N_1053,N_968,N_860);
or U1054 (N_1054,N_816,N_999);
and U1055 (N_1055,N_804,N_869);
nor U1056 (N_1056,N_914,N_831);
xnor U1057 (N_1057,N_861,N_913);
or U1058 (N_1058,N_850,N_814);
and U1059 (N_1059,N_940,N_935);
xnor U1060 (N_1060,N_849,N_888);
nor U1061 (N_1061,N_879,N_835);
nand U1062 (N_1062,N_899,N_841);
or U1063 (N_1063,N_893,N_832);
nand U1064 (N_1064,N_851,N_966);
or U1065 (N_1065,N_945,N_909);
and U1066 (N_1066,N_822,N_932);
nand U1067 (N_1067,N_963,N_859);
and U1068 (N_1068,N_957,N_848);
nor U1069 (N_1069,N_834,N_854);
nor U1070 (N_1070,N_931,N_875);
and U1071 (N_1071,N_954,N_891);
nor U1072 (N_1072,N_927,N_912);
nor U1073 (N_1073,N_870,N_811);
nor U1074 (N_1074,N_930,N_922);
and U1075 (N_1075,N_838,N_876);
nand U1076 (N_1076,N_813,N_868);
or U1077 (N_1077,N_993,N_916);
nand U1078 (N_1078,N_948,N_923);
or U1079 (N_1079,N_821,N_985);
nand U1080 (N_1080,N_998,N_905);
or U1081 (N_1081,N_863,N_943);
nor U1082 (N_1082,N_829,N_973);
or U1083 (N_1083,N_889,N_885);
nand U1084 (N_1084,N_886,N_866);
and U1085 (N_1085,N_938,N_915);
nor U1086 (N_1086,N_936,N_949);
or U1087 (N_1087,N_976,N_839);
or U1088 (N_1088,N_920,N_926);
nor U1089 (N_1089,N_971,N_980);
and U1090 (N_1090,N_836,N_995);
or U1091 (N_1091,N_884,N_933);
nor U1092 (N_1092,N_827,N_965);
and U1093 (N_1093,N_964,N_952);
or U1094 (N_1094,N_818,N_901);
and U1095 (N_1095,N_830,N_874);
nor U1096 (N_1096,N_925,N_820);
or U1097 (N_1097,N_867,N_815);
and U1098 (N_1098,N_929,N_904);
and U1099 (N_1099,N_819,N_937);
or U1100 (N_1100,N_956,N_947);
xnor U1101 (N_1101,N_922,N_939);
nand U1102 (N_1102,N_897,N_813);
and U1103 (N_1103,N_964,N_853);
and U1104 (N_1104,N_913,N_836);
or U1105 (N_1105,N_851,N_927);
and U1106 (N_1106,N_880,N_889);
or U1107 (N_1107,N_816,N_846);
and U1108 (N_1108,N_822,N_829);
and U1109 (N_1109,N_867,N_944);
nor U1110 (N_1110,N_919,N_862);
and U1111 (N_1111,N_954,N_964);
and U1112 (N_1112,N_867,N_969);
nor U1113 (N_1113,N_956,N_854);
nor U1114 (N_1114,N_895,N_935);
nand U1115 (N_1115,N_928,N_931);
nand U1116 (N_1116,N_957,N_822);
and U1117 (N_1117,N_913,N_822);
and U1118 (N_1118,N_873,N_919);
nand U1119 (N_1119,N_861,N_865);
nor U1120 (N_1120,N_903,N_874);
nand U1121 (N_1121,N_850,N_816);
nor U1122 (N_1122,N_967,N_810);
and U1123 (N_1123,N_873,N_958);
and U1124 (N_1124,N_976,N_953);
and U1125 (N_1125,N_860,N_849);
or U1126 (N_1126,N_895,N_900);
or U1127 (N_1127,N_967,N_844);
or U1128 (N_1128,N_864,N_863);
or U1129 (N_1129,N_915,N_931);
or U1130 (N_1130,N_995,N_849);
nand U1131 (N_1131,N_800,N_818);
nor U1132 (N_1132,N_959,N_943);
nor U1133 (N_1133,N_814,N_998);
or U1134 (N_1134,N_965,N_985);
or U1135 (N_1135,N_909,N_882);
nand U1136 (N_1136,N_823,N_872);
or U1137 (N_1137,N_838,N_901);
xnor U1138 (N_1138,N_812,N_847);
nor U1139 (N_1139,N_937,N_877);
and U1140 (N_1140,N_987,N_873);
and U1141 (N_1141,N_998,N_952);
nand U1142 (N_1142,N_979,N_876);
nor U1143 (N_1143,N_898,N_817);
and U1144 (N_1144,N_980,N_966);
xnor U1145 (N_1145,N_876,N_972);
and U1146 (N_1146,N_999,N_809);
nand U1147 (N_1147,N_812,N_852);
and U1148 (N_1148,N_848,N_887);
or U1149 (N_1149,N_922,N_877);
or U1150 (N_1150,N_833,N_962);
nor U1151 (N_1151,N_940,N_832);
nand U1152 (N_1152,N_842,N_871);
and U1153 (N_1153,N_898,N_918);
or U1154 (N_1154,N_856,N_933);
and U1155 (N_1155,N_937,N_830);
nor U1156 (N_1156,N_838,N_854);
nor U1157 (N_1157,N_943,N_822);
xor U1158 (N_1158,N_864,N_927);
nand U1159 (N_1159,N_836,N_979);
xnor U1160 (N_1160,N_802,N_862);
nor U1161 (N_1161,N_908,N_859);
nor U1162 (N_1162,N_829,N_969);
nand U1163 (N_1163,N_943,N_826);
nand U1164 (N_1164,N_940,N_863);
and U1165 (N_1165,N_878,N_934);
nand U1166 (N_1166,N_871,N_892);
xor U1167 (N_1167,N_963,N_938);
nor U1168 (N_1168,N_837,N_856);
or U1169 (N_1169,N_828,N_839);
nor U1170 (N_1170,N_803,N_906);
nor U1171 (N_1171,N_981,N_971);
or U1172 (N_1172,N_897,N_965);
or U1173 (N_1173,N_994,N_912);
and U1174 (N_1174,N_958,N_952);
nand U1175 (N_1175,N_979,N_838);
nand U1176 (N_1176,N_917,N_839);
xor U1177 (N_1177,N_960,N_840);
nand U1178 (N_1178,N_839,N_924);
nand U1179 (N_1179,N_863,N_961);
nand U1180 (N_1180,N_946,N_933);
nand U1181 (N_1181,N_803,N_990);
xnor U1182 (N_1182,N_943,N_988);
nand U1183 (N_1183,N_955,N_908);
and U1184 (N_1184,N_970,N_870);
nor U1185 (N_1185,N_834,N_981);
nor U1186 (N_1186,N_979,N_955);
or U1187 (N_1187,N_955,N_952);
nand U1188 (N_1188,N_994,N_983);
nor U1189 (N_1189,N_966,N_853);
nand U1190 (N_1190,N_891,N_809);
or U1191 (N_1191,N_963,N_928);
or U1192 (N_1192,N_842,N_807);
nand U1193 (N_1193,N_843,N_995);
and U1194 (N_1194,N_918,N_943);
nand U1195 (N_1195,N_965,N_835);
nand U1196 (N_1196,N_945,N_992);
and U1197 (N_1197,N_922,N_849);
and U1198 (N_1198,N_855,N_952);
or U1199 (N_1199,N_844,N_853);
or U1200 (N_1200,N_1183,N_1185);
nand U1201 (N_1201,N_1144,N_1163);
or U1202 (N_1202,N_1145,N_1141);
or U1203 (N_1203,N_1026,N_1174);
or U1204 (N_1204,N_1077,N_1184);
or U1205 (N_1205,N_1052,N_1090);
and U1206 (N_1206,N_1119,N_1007);
or U1207 (N_1207,N_1188,N_1057);
nor U1208 (N_1208,N_1017,N_1045);
and U1209 (N_1209,N_1053,N_1033);
nand U1210 (N_1210,N_1056,N_1100);
and U1211 (N_1211,N_1051,N_1086);
or U1212 (N_1212,N_1061,N_1170);
nor U1213 (N_1213,N_1175,N_1084);
nor U1214 (N_1214,N_1194,N_1187);
or U1215 (N_1215,N_1089,N_1028);
nand U1216 (N_1216,N_1124,N_1004);
and U1217 (N_1217,N_1066,N_1158);
or U1218 (N_1218,N_1074,N_1073);
nand U1219 (N_1219,N_1039,N_1070);
and U1220 (N_1220,N_1103,N_1147);
or U1221 (N_1221,N_1037,N_1035);
or U1222 (N_1222,N_1142,N_1038);
or U1223 (N_1223,N_1022,N_1101);
or U1224 (N_1224,N_1027,N_1156);
nand U1225 (N_1225,N_1139,N_1064);
or U1226 (N_1226,N_1161,N_1008);
nand U1227 (N_1227,N_1166,N_1012);
or U1228 (N_1228,N_1058,N_1047);
nor U1229 (N_1229,N_1136,N_1195);
nand U1230 (N_1230,N_1099,N_1079);
or U1231 (N_1231,N_1189,N_1190);
nand U1232 (N_1232,N_1126,N_1009);
nor U1233 (N_1233,N_1067,N_1143);
nor U1234 (N_1234,N_1010,N_1002);
or U1235 (N_1235,N_1111,N_1042);
or U1236 (N_1236,N_1078,N_1034);
and U1237 (N_1237,N_1081,N_1133);
nand U1238 (N_1238,N_1129,N_1065);
nand U1239 (N_1239,N_1054,N_1121);
xnor U1240 (N_1240,N_1006,N_1076);
and U1241 (N_1241,N_1000,N_1036);
and U1242 (N_1242,N_1193,N_1055);
and U1243 (N_1243,N_1113,N_1062);
and U1244 (N_1244,N_1085,N_1025);
nor U1245 (N_1245,N_1063,N_1160);
and U1246 (N_1246,N_1082,N_1107);
nor U1247 (N_1247,N_1146,N_1180);
and U1248 (N_1248,N_1024,N_1023);
nor U1249 (N_1249,N_1117,N_1095);
nand U1250 (N_1250,N_1131,N_1182);
and U1251 (N_1251,N_1106,N_1165);
and U1252 (N_1252,N_1071,N_1114);
or U1253 (N_1253,N_1031,N_1198);
nand U1254 (N_1254,N_1177,N_1016);
nand U1255 (N_1255,N_1197,N_1030);
nand U1256 (N_1256,N_1186,N_1029);
and U1257 (N_1257,N_1068,N_1155);
or U1258 (N_1258,N_1151,N_1118);
and U1259 (N_1259,N_1132,N_1092);
xor U1260 (N_1260,N_1072,N_1087);
and U1261 (N_1261,N_1169,N_1013);
nor U1262 (N_1262,N_1032,N_1152);
or U1263 (N_1263,N_1014,N_1130);
and U1264 (N_1264,N_1199,N_1043);
and U1265 (N_1265,N_1097,N_1148);
and U1266 (N_1266,N_1019,N_1179);
or U1267 (N_1267,N_1112,N_1011);
nor U1268 (N_1268,N_1167,N_1127);
or U1269 (N_1269,N_1021,N_1005);
and U1270 (N_1270,N_1088,N_1003);
nand U1271 (N_1271,N_1134,N_1049);
and U1272 (N_1272,N_1162,N_1122);
nand U1273 (N_1273,N_1080,N_1060);
nor U1274 (N_1274,N_1181,N_1140);
nor U1275 (N_1275,N_1115,N_1135);
or U1276 (N_1276,N_1120,N_1123);
or U1277 (N_1277,N_1105,N_1137);
and U1278 (N_1278,N_1116,N_1171);
nor U1279 (N_1279,N_1048,N_1096);
nand U1280 (N_1280,N_1157,N_1075);
and U1281 (N_1281,N_1018,N_1150);
nor U1282 (N_1282,N_1091,N_1154);
nor U1283 (N_1283,N_1098,N_1196);
nor U1284 (N_1284,N_1041,N_1138);
or U1285 (N_1285,N_1176,N_1153);
nand U1286 (N_1286,N_1125,N_1172);
xnor U1287 (N_1287,N_1173,N_1040);
or U1288 (N_1288,N_1159,N_1164);
and U1289 (N_1289,N_1108,N_1102);
or U1290 (N_1290,N_1192,N_1069);
nand U1291 (N_1291,N_1149,N_1059);
nand U1292 (N_1292,N_1093,N_1015);
nand U1293 (N_1293,N_1191,N_1104);
nor U1294 (N_1294,N_1109,N_1128);
and U1295 (N_1295,N_1001,N_1046);
xnor U1296 (N_1296,N_1094,N_1083);
and U1297 (N_1297,N_1168,N_1178);
nand U1298 (N_1298,N_1044,N_1110);
xor U1299 (N_1299,N_1050,N_1020);
xor U1300 (N_1300,N_1109,N_1161);
nand U1301 (N_1301,N_1054,N_1179);
and U1302 (N_1302,N_1142,N_1139);
or U1303 (N_1303,N_1010,N_1035);
and U1304 (N_1304,N_1044,N_1125);
nor U1305 (N_1305,N_1054,N_1188);
and U1306 (N_1306,N_1098,N_1047);
or U1307 (N_1307,N_1157,N_1009);
nor U1308 (N_1308,N_1044,N_1106);
and U1309 (N_1309,N_1166,N_1014);
and U1310 (N_1310,N_1170,N_1185);
nand U1311 (N_1311,N_1179,N_1191);
nor U1312 (N_1312,N_1143,N_1198);
or U1313 (N_1313,N_1051,N_1032);
and U1314 (N_1314,N_1138,N_1064);
or U1315 (N_1315,N_1035,N_1154);
and U1316 (N_1316,N_1096,N_1166);
or U1317 (N_1317,N_1163,N_1116);
nor U1318 (N_1318,N_1183,N_1179);
or U1319 (N_1319,N_1124,N_1111);
and U1320 (N_1320,N_1075,N_1064);
nand U1321 (N_1321,N_1179,N_1164);
and U1322 (N_1322,N_1127,N_1134);
nor U1323 (N_1323,N_1024,N_1015);
or U1324 (N_1324,N_1108,N_1119);
nand U1325 (N_1325,N_1055,N_1049);
or U1326 (N_1326,N_1193,N_1002);
nor U1327 (N_1327,N_1002,N_1016);
nor U1328 (N_1328,N_1003,N_1017);
and U1329 (N_1329,N_1164,N_1121);
nand U1330 (N_1330,N_1099,N_1134);
nor U1331 (N_1331,N_1157,N_1028);
and U1332 (N_1332,N_1046,N_1062);
or U1333 (N_1333,N_1034,N_1062);
or U1334 (N_1334,N_1113,N_1129);
and U1335 (N_1335,N_1005,N_1084);
and U1336 (N_1336,N_1114,N_1100);
or U1337 (N_1337,N_1129,N_1071);
and U1338 (N_1338,N_1146,N_1029);
and U1339 (N_1339,N_1053,N_1045);
and U1340 (N_1340,N_1013,N_1175);
and U1341 (N_1341,N_1091,N_1039);
nand U1342 (N_1342,N_1099,N_1155);
and U1343 (N_1343,N_1186,N_1015);
nor U1344 (N_1344,N_1022,N_1192);
and U1345 (N_1345,N_1057,N_1092);
nor U1346 (N_1346,N_1076,N_1128);
and U1347 (N_1347,N_1045,N_1080);
and U1348 (N_1348,N_1024,N_1124);
or U1349 (N_1349,N_1194,N_1039);
and U1350 (N_1350,N_1077,N_1056);
nor U1351 (N_1351,N_1032,N_1064);
or U1352 (N_1352,N_1013,N_1093);
nand U1353 (N_1353,N_1073,N_1121);
or U1354 (N_1354,N_1162,N_1168);
or U1355 (N_1355,N_1075,N_1178);
and U1356 (N_1356,N_1139,N_1162);
and U1357 (N_1357,N_1058,N_1106);
nand U1358 (N_1358,N_1113,N_1197);
or U1359 (N_1359,N_1143,N_1007);
xor U1360 (N_1360,N_1058,N_1060);
and U1361 (N_1361,N_1137,N_1018);
nor U1362 (N_1362,N_1121,N_1151);
and U1363 (N_1363,N_1163,N_1185);
nand U1364 (N_1364,N_1042,N_1067);
xnor U1365 (N_1365,N_1000,N_1175);
nand U1366 (N_1366,N_1183,N_1012);
nand U1367 (N_1367,N_1134,N_1135);
nand U1368 (N_1368,N_1116,N_1026);
nand U1369 (N_1369,N_1160,N_1143);
nor U1370 (N_1370,N_1062,N_1152);
or U1371 (N_1371,N_1019,N_1075);
and U1372 (N_1372,N_1040,N_1022);
or U1373 (N_1373,N_1043,N_1133);
or U1374 (N_1374,N_1007,N_1079);
nand U1375 (N_1375,N_1081,N_1165);
or U1376 (N_1376,N_1133,N_1188);
nand U1377 (N_1377,N_1121,N_1071);
or U1378 (N_1378,N_1180,N_1102);
xnor U1379 (N_1379,N_1193,N_1178);
nor U1380 (N_1380,N_1006,N_1173);
and U1381 (N_1381,N_1054,N_1013);
nor U1382 (N_1382,N_1001,N_1024);
nand U1383 (N_1383,N_1161,N_1141);
or U1384 (N_1384,N_1008,N_1139);
nand U1385 (N_1385,N_1099,N_1047);
nand U1386 (N_1386,N_1104,N_1100);
and U1387 (N_1387,N_1012,N_1152);
and U1388 (N_1388,N_1123,N_1092);
or U1389 (N_1389,N_1097,N_1028);
or U1390 (N_1390,N_1032,N_1175);
or U1391 (N_1391,N_1010,N_1018);
or U1392 (N_1392,N_1185,N_1023);
or U1393 (N_1393,N_1133,N_1000);
nand U1394 (N_1394,N_1124,N_1157);
nor U1395 (N_1395,N_1085,N_1133);
or U1396 (N_1396,N_1137,N_1111);
and U1397 (N_1397,N_1176,N_1177);
nand U1398 (N_1398,N_1104,N_1019);
and U1399 (N_1399,N_1143,N_1045);
nand U1400 (N_1400,N_1360,N_1316);
nor U1401 (N_1401,N_1386,N_1392);
and U1402 (N_1402,N_1319,N_1367);
nor U1403 (N_1403,N_1331,N_1333);
nand U1404 (N_1404,N_1325,N_1390);
nand U1405 (N_1405,N_1362,N_1312);
nor U1406 (N_1406,N_1346,N_1223);
xnor U1407 (N_1407,N_1222,N_1322);
nand U1408 (N_1408,N_1289,N_1294);
nor U1409 (N_1409,N_1241,N_1343);
nand U1410 (N_1410,N_1368,N_1206);
and U1411 (N_1411,N_1345,N_1204);
or U1412 (N_1412,N_1202,N_1363);
or U1413 (N_1413,N_1259,N_1359);
nor U1414 (N_1414,N_1284,N_1209);
or U1415 (N_1415,N_1290,N_1315);
nor U1416 (N_1416,N_1364,N_1227);
or U1417 (N_1417,N_1366,N_1313);
and U1418 (N_1418,N_1354,N_1207);
and U1419 (N_1419,N_1212,N_1302);
nor U1420 (N_1420,N_1306,N_1340);
nand U1421 (N_1421,N_1213,N_1371);
xnor U1422 (N_1422,N_1307,N_1246);
or U1423 (N_1423,N_1234,N_1327);
and U1424 (N_1424,N_1203,N_1385);
nor U1425 (N_1425,N_1298,N_1239);
nand U1426 (N_1426,N_1244,N_1301);
nand U1427 (N_1427,N_1262,N_1278);
and U1428 (N_1428,N_1361,N_1226);
and U1429 (N_1429,N_1251,N_1281);
nand U1430 (N_1430,N_1231,N_1374);
nand U1431 (N_1431,N_1372,N_1376);
nor U1432 (N_1432,N_1344,N_1309);
nor U1433 (N_1433,N_1394,N_1377);
nor U1434 (N_1434,N_1342,N_1381);
or U1435 (N_1435,N_1242,N_1235);
nand U1436 (N_1436,N_1237,N_1317);
and U1437 (N_1437,N_1349,N_1238);
nand U1438 (N_1438,N_1250,N_1382);
nand U1439 (N_1439,N_1240,N_1264);
nand U1440 (N_1440,N_1348,N_1395);
nor U1441 (N_1441,N_1308,N_1283);
nand U1442 (N_1442,N_1273,N_1351);
nand U1443 (N_1443,N_1224,N_1274);
or U1444 (N_1444,N_1225,N_1334);
nand U1445 (N_1445,N_1350,N_1339);
and U1446 (N_1446,N_1379,N_1230);
or U1447 (N_1447,N_1297,N_1210);
nand U1448 (N_1448,N_1338,N_1214);
and U1449 (N_1449,N_1287,N_1201);
or U1450 (N_1450,N_1275,N_1292);
nor U1451 (N_1451,N_1326,N_1229);
or U1452 (N_1452,N_1286,N_1267);
and U1453 (N_1453,N_1279,N_1356);
or U1454 (N_1454,N_1268,N_1398);
or U1455 (N_1455,N_1248,N_1258);
nand U1456 (N_1456,N_1249,N_1310);
nor U1457 (N_1457,N_1216,N_1266);
nor U1458 (N_1458,N_1300,N_1329);
nand U1459 (N_1459,N_1369,N_1221);
nand U1460 (N_1460,N_1337,N_1296);
or U1461 (N_1461,N_1393,N_1357);
nor U1462 (N_1462,N_1263,N_1341);
nand U1463 (N_1463,N_1358,N_1208);
nand U1464 (N_1464,N_1270,N_1261);
nand U1465 (N_1465,N_1311,N_1236);
nor U1466 (N_1466,N_1255,N_1330);
and U1467 (N_1467,N_1220,N_1388);
and U1468 (N_1468,N_1355,N_1254);
and U1469 (N_1469,N_1397,N_1277);
and U1470 (N_1470,N_1218,N_1257);
and U1471 (N_1471,N_1347,N_1217);
or U1472 (N_1472,N_1352,N_1332);
or U1473 (N_1473,N_1387,N_1378);
and U1474 (N_1474,N_1375,N_1205);
nand U1475 (N_1475,N_1276,N_1291);
nor U1476 (N_1476,N_1314,N_1233);
nor U1477 (N_1477,N_1324,N_1280);
xor U1478 (N_1478,N_1293,N_1336);
or U1479 (N_1479,N_1320,N_1295);
nor U1480 (N_1480,N_1271,N_1399);
and U1481 (N_1481,N_1200,N_1282);
and U1482 (N_1482,N_1365,N_1335);
and U1483 (N_1483,N_1305,N_1391);
nand U1484 (N_1484,N_1256,N_1260);
nor U1485 (N_1485,N_1396,N_1228);
nor U1486 (N_1486,N_1373,N_1253);
nand U1487 (N_1487,N_1243,N_1323);
nand U1488 (N_1488,N_1252,N_1389);
or U1489 (N_1489,N_1318,N_1219);
nand U1490 (N_1490,N_1353,N_1272);
nand U1491 (N_1491,N_1211,N_1304);
or U1492 (N_1492,N_1299,N_1232);
nor U1493 (N_1493,N_1328,N_1380);
nor U1494 (N_1494,N_1303,N_1215);
or U1495 (N_1495,N_1370,N_1288);
and U1496 (N_1496,N_1321,N_1265);
nor U1497 (N_1497,N_1285,N_1269);
and U1498 (N_1498,N_1247,N_1383);
nor U1499 (N_1499,N_1384,N_1245);
or U1500 (N_1500,N_1217,N_1224);
nor U1501 (N_1501,N_1216,N_1374);
and U1502 (N_1502,N_1228,N_1359);
nand U1503 (N_1503,N_1368,N_1346);
or U1504 (N_1504,N_1319,N_1281);
nand U1505 (N_1505,N_1364,N_1279);
and U1506 (N_1506,N_1395,N_1224);
and U1507 (N_1507,N_1230,N_1399);
nor U1508 (N_1508,N_1335,N_1278);
and U1509 (N_1509,N_1253,N_1255);
or U1510 (N_1510,N_1351,N_1241);
or U1511 (N_1511,N_1287,N_1369);
nor U1512 (N_1512,N_1350,N_1248);
or U1513 (N_1513,N_1295,N_1225);
or U1514 (N_1514,N_1367,N_1228);
xor U1515 (N_1515,N_1299,N_1270);
or U1516 (N_1516,N_1335,N_1284);
or U1517 (N_1517,N_1261,N_1316);
and U1518 (N_1518,N_1240,N_1279);
or U1519 (N_1519,N_1284,N_1321);
nand U1520 (N_1520,N_1240,N_1208);
and U1521 (N_1521,N_1276,N_1391);
and U1522 (N_1522,N_1381,N_1247);
nand U1523 (N_1523,N_1300,N_1267);
nor U1524 (N_1524,N_1382,N_1348);
nand U1525 (N_1525,N_1371,N_1271);
nor U1526 (N_1526,N_1273,N_1377);
and U1527 (N_1527,N_1222,N_1380);
nor U1528 (N_1528,N_1298,N_1335);
nor U1529 (N_1529,N_1308,N_1334);
or U1530 (N_1530,N_1392,N_1270);
nand U1531 (N_1531,N_1202,N_1373);
and U1532 (N_1532,N_1260,N_1287);
or U1533 (N_1533,N_1207,N_1383);
nand U1534 (N_1534,N_1379,N_1260);
or U1535 (N_1535,N_1381,N_1323);
xor U1536 (N_1536,N_1288,N_1385);
and U1537 (N_1537,N_1345,N_1286);
nand U1538 (N_1538,N_1201,N_1375);
or U1539 (N_1539,N_1316,N_1242);
or U1540 (N_1540,N_1371,N_1369);
nor U1541 (N_1541,N_1283,N_1311);
and U1542 (N_1542,N_1217,N_1207);
nor U1543 (N_1543,N_1310,N_1313);
or U1544 (N_1544,N_1256,N_1392);
or U1545 (N_1545,N_1229,N_1270);
nand U1546 (N_1546,N_1363,N_1304);
or U1547 (N_1547,N_1214,N_1388);
nand U1548 (N_1548,N_1280,N_1272);
nand U1549 (N_1549,N_1323,N_1340);
nand U1550 (N_1550,N_1379,N_1220);
nand U1551 (N_1551,N_1399,N_1298);
or U1552 (N_1552,N_1310,N_1268);
and U1553 (N_1553,N_1283,N_1224);
and U1554 (N_1554,N_1350,N_1360);
nor U1555 (N_1555,N_1272,N_1322);
nor U1556 (N_1556,N_1226,N_1391);
nor U1557 (N_1557,N_1328,N_1318);
or U1558 (N_1558,N_1328,N_1284);
or U1559 (N_1559,N_1322,N_1294);
or U1560 (N_1560,N_1202,N_1302);
and U1561 (N_1561,N_1257,N_1364);
nor U1562 (N_1562,N_1363,N_1365);
nor U1563 (N_1563,N_1372,N_1391);
xor U1564 (N_1564,N_1315,N_1341);
xor U1565 (N_1565,N_1259,N_1362);
and U1566 (N_1566,N_1326,N_1314);
nor U1567 (N_1567,N_1383,N_1295);
nor U1568 (N_1568,N_1254,N_1371);
nor U1569 (N_1569,N_1304,N_1370);
or U1570 (N_1570,N_1313,N_1299);
or U1571 (N_1571,N_1280,N_1385);
and U1572 (N_1572,N_1366,N_1247);
nand U1573 (N_1573,N_1321,N_1324);
nor U1574 (N_1574,N_1212,N_1219);
or U1575 (N_1575,N_1311,N_1284);
or U1576 (N_1576,N_1322,N_1285);
or U1577 (N_1577,N_1215,N_1321);
or U1578 (N_1578,N_1254,N_1294);
or U1579 (N_1579,N_1315,N_1249);
nor U1580 (N_1580,N_1289,N_1356);
nand U1581 (N_1581,N_1322,N_1271);
nor U1582 (N_1582,N_1341,N_1253);
and U1583 (N_1583,N_1345,N_1336);
and U1584 (N_1584,N_1396,N_1330);
nor U1585 (N_1585,N_1392,N_1280);
or U1586 (N_1586,N_1252,N_1265);
nand U1587 (N_1587,N_1315,N_1378);
nand U1588 (N_1588,N_1269,N_1267);
nand U1589 (N_1589,N_1343,N_1393);
nor U1590 (N_1590,N_1352,N_1274);
nand U1591 (N_1591,N_1348,N_1248);
nor U1592 (N_1592,N_1395,N_1209);
nor U1593 (N_1593,N_1238,N_1311);
and U1594 (N_1594,N_1343,N_1377);
or U1595 (N_1595,N_1320,N_1242);
and U1596 (N_1596,N_1215,N_1371);
nand U1597 (N_1597,N_1282,N_1254);
nor U1598 (N_1598,N_1257,N_1388);
nand U1599 (N_1599,N_1251,N_1259);
and U1600 (N_1600,N_1439,N_1477);
nand U1601 (N_1601,N_1554,N_1447);
or U1602 (N_1602,N_1536,N_1540);
nand U1603 (N_1603,N_1524,N_1589);
nor U1604 (N_1604,N_1487,N_1517);
xor U1605 (N_1605,N_1598,N_1462);
or U1606 (N_1606,N_1522,N_1456);
nand U1607 (N_1607,N_1430,N_1472);
nor U1608 (N_1608,N_1491,N_1459);
nor U1609 (N_1609,N_1575,N_1461);
nand U1610 (N_1610,N_1452,N_1403);
and U1611 (N_1611,N_1486,N_1577);
nor U1612 (N_1612,N_1493,N_1564);
or U1613 (N_1613,N_1431,N_1531);
or U1614 (N_1614,N_1543,N_1547);
or U1615 (N_1615,N_1586,N_1545);
and U1616 (N_1616,N_1433,N_1469);
nand U1617 (N_1617,N_1408,N_1597);
nand U1618 (N_1618,N_1502,N_1466);
nand U1619 (N_1619,N_1425,N_1513);
nand U1620 (N_1620,N_1407,N_1457);
nor U1621 (N_1621,N_1500,N_1595);
nor U1622 (N_1622,N_1567,N_1555);
nor U1623 (N_1623,N_1497,N_1580);
and U1624 (N_1624,N_1578,N_1458);
nor U1625 (N_1625,N_1551,N_1561);
xnor U1626 (N_1626,N_1473,N_1516);
nand U1627 (N_1627,N_1566,N_1599);
and U1628 (N_1628,N_1539,N_1406);
nor U1629 (N_1629,N_1441,N_1581);
nand U1630 (N_1630,N_1585,N_1565);
nor U1631 (N_1631,N_1488,N_1549);
nor U1632 (N_1632,N_1507,N_1440);
nor U1633 (N_1633,N_1509,N_1557);
nand U1634 (N_1634,N_1498,N_1501);
nand U1635 (N_1635,N_1423,N_1404);
or U1636 (N_1636,N_1582,N_1448);
and U1637 (N_1637,N_1527,N_1492);
or U1638 (N_1638,N_1427,N_1428);
and U1639 (N_1639,N_1515,N_1568);
or U1640 (N_1640,N_1400,N_1401);
nand U1641 (N_1641,N_1533,N_1437);
nand U1642 (N_1642,N_1429,N_1525);
nand U1643 (N_1643,N_1519,N_1411);
and U1644 (N_1644,N_1419,N_1454);
and U1645 (N_1645,N_1446,N_1535);
and U1646 (N_1646,N_1420,N_1546);
nand U1647 (N_1647,N_1479,N_1591);
nand U1648 (N_1648,N_1444,N_1475);
and U1649 (N_1649,N_1442,N_1559);
nor U1650 (N_1650,N_1571,N_1542);
nand U1651 (N_1651,N_1592,N_1482);
and U1652 (N_1652,N_1421,N_1504);
or U1653 (N_1653,N_1455,N_1460);
and U1654 (N_1654,N_1449,N_1453);
nor U1655 (N_1655,N_1529,N_1410);
nor U1656 (N_1656,N_1481,N_1450);
or U1657 (N_1657,N_1537,N_1532);
and U1658 (N_1658,N_1424,N_1576);
nand U1659 (N_1659,N_1484,N_1414);
or U1660 (N_1660,N_1534,N_1463);
xnor U1661 (N_1661,N_1478,N_1587);
or U1662 (N_1662,N_1583,N_1518);
and U1663 (N_1663,N_1584,N_1552);
and U1664 (N_1664,N_1499,N_1530);
nor U1665 (N_1665,N_1467,N_1569);
and U1666 (N_1666,N_1574,N_1523);
nand U1667 (N_1667,N_1505,N_1512);
nor U1668 (N_1668,N_1506,N_1415);
and U1669 (N_1669,N_1483,N_1538);
nand U1670 (N_1670,N_1476,N_1528);
nand U1671 (N_1671,N_1511,N_1548);
and U1672 (N_1672,N_1405,N_1544);
nor U1673 (N_1673,N_1560,N_1471);
nor U1674 (N_1674,N_1572,N_1418);
and U1675 (N_1675,N_1485,N_1436);
nor U1676 (N_1676,N_1489,N_1470);
or U1677 (N_1677,N_1556,N_1417);
and U1678 (N_1678,N_1520,N_1496);
nor U1679 (N_1679,N_1490,N_1553);
and U1680 (N_1680,N_1503,N_1445);
nor U1681 (N_1681,N_1521,N_1426);
nand U1682 (N_1682,N_1413,N_1579);
and U1683 (N_1683,N_1468,N_1465);
or U1684 (N_1684,N_1573,N_1435);
nor U1685 (N_1685,N_1588,N_1443);
or U1686 (N_1686,N_1409,N_1495);
nand U1687 (N_1687,N_1422,N_1590);
and U1688 (N_1688,N_1510,N_1563);
or U1689 (N_1689,N_1412,N_1451);
nand U1690 (N_1690,N_1416,N_1494);
nor U1691 (N_1691,N_1526,N_1402);
and U1692 (N_1692,N_1558,N_1593);
and U1693 (N_1693,N_1562,N_1514);
nand U1694 (N_1694,N_1432,N_1541);
nand U1695 (N_1695,N_1594,N_1438);
and U1696 (N_1696,N_1474,N_1596);
or U1697 (N_1697,N_1434,N_1508);
and U1698 (N_1698,N_1464,N_1570);
nand U1699 (N_1699,N_1550,N_1480);
nor U1700 (N_1700,N_1555,N_1443);
nor U1701 (N_1701,N_1410,N_1556);
and U1702 (N_1702,N_1499,N_1452);
and U1703 (N_1703,N_1451,N_1529);
nand U1704 (N_1704,N_1597,N_1561);
xor U1705 (N_1705,N_1555,N_1562);
nor U1706 (N_1706,N_1589,N_1473);
nor U1707 (N_1707,N_1553,N_1561);
or U1708 (N_1708,N_1411,N_1504);
and U1709 (N_1709,N_1410,N_1547);
or U1710 (N_1710,N_1476,N_1409);
xor U1711 (N_1711,N_1445,N_1528);
nor U1712 (N_1712,N_1557,N_1497);
or U1713 (N_1713,N_1577,N_1561);
nor U1714 (N_1714,N_1429,N_1454);
nand U1715 (N_1715,N_1464,N_1467);
or U1716 (N_1716,N_1414,N_1428);
nor U1717 (N_1717,N_1444,N_1472);
and U1718 (N_1718,N_1571,N_1494);
and U1719 (N_1719,N_1491,N_1462);
nand U1720 (N_1720,N_1599,N_1440);
nor U1721 (N_1721,N_1592,N_1411);
nand U1722 (N_1722,N_1525,N_1509);
or U1723 (N_1723,N_1492,N_1458);
or U1724 (N_1724,N_1509,N_1503);
nor U1725 (N_1725,N_1578,N_1450);
or U1726 (N_1726,N_1567,N_1546);
nor U1727 (N_1727,N_1581,N_1521);
and U1728 (N_1728,N_1459,N_1407);
nand U1729 (N_1729,N_1427,N_1441);
nor U1730 (N_1730,N_1575,N_1424);
and U1731 (N_1731,N_1440,N_1418);
and U1732 (N_1732,N_1594,N_1536);
nand U1733 (N_1733,N_1473,N_1436);
and U1734 (N_1734,N_1452,N_1434);
nor U1735 (N_1735,N_1508,N_1401);
and U1736 (N_1736,N_1543,N_1569);
and U1737 (N_1737,N_1400,N_1438);
nand U1738 (N_1738,N_1557,N_1570);
and U1739 (N_1739,N_1559,N_1450);
nand U1740 (N_1740,N_1538,N_1584);
and U1741 (N_1741,N_1472,N_1576);
and U1742 (N_1742,N_1585,N_1480);
nor U1743 (N_1743,N_1591,N_1464);
and U1744 (N_1744,N_1591,N_1506);
or U1745 (N_1745,N_1446,N_1505);
nand U1746 (N_1746,N_1518,N_1447);
or U1747 (N_1747,N_1479,N_1533);
nand U1748 (N_1748,N_1426,N_1474);
and U1749 (N_1749,N_1586,N_1408);
or U1750 (N_1750,N_1409,N_1452);
and U1751 (N_1751,N_1478,N_1504);
and U1752 (N_1752,N_1471,N_1459);
or U1753 (N_1753,N_1578,N_1537);
and U1754 (N_1754,N_1585,N_1578);
and U1755 (N_1755,N_1499,N_1412);
nand U1756 (N_1756,N_1586,N_1594);
nor U1757 (N_1757,N_1552,N_1448);
and U1758 (N_1758,N_1474,N_1574);
nand U1759 (N_1759,N_1507,N_1451);
nor U1760 (N_1760,N_1582,N_1570);
nor U1761 (N_1761,N_1556,N_1503);
or U1762 (N_1762,N_1511,N_1555);
nor U1763 (N_1763,N_1408,N_1580);
or U1764 (N_1764,N_1528,N_1414);
nor U1765 (N_1765,N_1474,N_1484);
or U1766 (N_1766,N_1519,N_1560);
or U1767 (N_1767,N_1469,N_1456);
or U1768 (N_1768,N_1573,N_1599);
or U1769 (N_1769,N_1484,N_1430);
nand U1770 (N_1770,N_1449,N_1548);
nor U1771 (N_1771,N_1595,N_1449);
and U1772 (N_1772,N_1542,N_1519);
nand U1773 (N_1773,N_1425,N_1497);
or U1774 (N_1774,N_1599,N_1477);
or U1775 (N_1775,N_1480,N_1541);
and U1776 (N_1776,N_1517,N_1418);
nand U1777 (N_1777,N_1573,N_1438);
nand U1778 (N_1778,N_1404,N_1474);
and U1779 (N_1779,N_1408,N_1503);
and U1780 (N_1780,N_1580,N_1491);
and U1781 (N_1781,N_1539,N_1450);
nand U1782 (N_1782,N_1581,N_1571);
xor U1783 (N_1783,N_1416,N_1483);
nor U1784 (N_1784,N_1419,N_1472);
or U1785 (N_1785,N_1477,N_1579);
or U1786 (N_1786,N_1458,N_1432);
nor U1787 (N_1787,N_1402,N_1560);
or U1788 (N_1788,N_1405,N_1450);
nand U1789 (N_1789,N_1522,N_1587);
and U1790 (N_1790,N_1442,N_1517);
nand U1791 (N_1791,N_1514,N_1538);
or U1792 (N_1792,N_1402,N_1489);
and U1793 (N_1793,N_1531,N_1430);
and U1794 (N_1794,N_1411,N_1435);
nor U1795 (N_1795,N_1505,N_1527);
nor U1796 (N_1796,N_1544,N_1486);
or U1797 (N_1797,N_1488,N_1575);
or U1798 (N_1798,N_1564,N_1456);
nand U1799 (N_1799,N_1431,N_1532);
nor U1800 (N_1800,N_1724,N_1718);
nor U1801 (N_1801,N_1684,N_1733);
nor U1802 (N_1802,N_1672,N_1632);
or U1803 (N_1803,N_1622,N_1601);
nand U1804 (N_1804,N_1625,N_1780);
nand U1805 (N_1805,N_1777,N_1668);
or U1806 (N_1806,N_1706,N_1669);
or U1807 (N_1807,N_1652,N_1716);
nand U1808 (N_1808,N_1645,N_1756);
nand U1809 (N_1809,N_1656,N_1770);
and U1810 (N_1810,N_1795,N_1758);
nand U1811 (N_1811,N_1776,N_1786);
and U1812 (N_1812,N_1736,N_1710);
and U1813 (N_1813,N_1760,N_1750);
or U1814 (N_1814,N_1778,N_1737);
and U1815 (N_1815,N_1738,N_1744);
nand U1816 (N_1816,N_1748,N_1794);
nand U1817 (N_1817,N_1621,N_1779);
nand U1818 (N_1818,N_1715,N_1717);
nor U1819 (N_1819,N_1730,N_1734);
nand U1820 (N_1820,N_1785,N_1757);
nor U1821 (N_1821,N_1679,N_1709);
and U1822 (N_1822,N_1728,N_1775);
nand U1823 (N_1823,N_1612,N_1708);
or U1824 (N_1824,N_1751,N_1651);
nand U1825 (N_1825,N_1725,N_1713);
nor U1826 (N_1826,N_1610,N_1722);
nand U1827 (N_1827,N_1766,N_1634);
nand U1828 (N_1828,N_1793,N_1694);
and U1829 (N_1829,N_1602,N_1620);
nor U1830 (N_1830,N_1765,N_1752);
xor U1831 (N_1831,N_1721,N_1664);
nand U1832 (N_1832,N_1673,N_1646);
nor U1833 (N_1833,N_1675,N_1735);
or U1834 (N_1834,N_1643,N_1712);
and U1835 (N_1835,N_1799,N_1642);
nor U1836 (N_1836,N_1665,N_1663);
nor U1837 (N_1837,N_1636,N_1635);
or U1838 (N_1838,N_1661,N_1639);
nand U1839 (N_1839,N_1792,N_1696);
nand U1840 (N_1840,N_1617,N_1774);
or U1841 (N_1841,N_1747,N_1729);
or U1842 (N_1842,N_1726,N_1787);
nor U1843 (N_1843,N_1740,N_1743);
nor U1844 (N_1844,N_1703,N_1604);
nor U1845 (N_1845,N_1631,N_1692);
nor U1846 (N_1846,N_1682,N_1781);
or U1847 (N_1847,N_1678,N_1783);
nand U1848 (N_1848,N_1723,N_1633);
nor U1849 (N_1849,N_1666,N_1767);
or U1850 (N_1850,N_1640,N_1641);
and U1851 (N_1851,N_1627,N_1690);
or U1852 (N_1852,N_1687,N_1732);
nor U1853 (N_1853,N_1741,N_1659);
nor U1854 (N_1854,N_1600,N_1603);
and U1855 (N_1855,N_1768,N_1697);
or U1856 (N_1856,N_1688,N_1790);
nor U1857 (N_1857,N_1662,N_1611);
or U1858 (N_1858,N_1615,N_1624);
nor U1859 (N_1859,N_1759,N_1686);
nor U1860 (N_1860,N_1771,N_1745);
nand U1861 (N_1861,N_1711,N_1784);
or U1862 (N_1862,N_1695,N_1755);
nor U1863 (N_1863,N_1658,N_1764);
nand U1864 (N_1864,N_1613,N_1731);
nand U1865 (N_1865,N_1677,N_1763);
and U1866 (N_1866,N_1623,N_1693);
and U1867 (N_1867,N_1796,N_1773);
and U1868 (N_1868,N_1788,N_1618);
nand U1869 (N_1869,N_1655,N_1746);
or U1870 (N_1870,N_1648,N_1791);
or U1871 (N_1871,N_1691,N_1720);
nand U1872 (N_1872,N_1647,N_1742);
nand U1873 (N_1873,N_1689,N_1671);
nor U1874 (N_1874,N_1719,N_1714);
nand U1875 (N_1875,N_1685,N_1700);
and U1876 (N_1876,N_1749,N_1619);
or U1877 (N_1877,N_1630,N_1654);
nor U1878 (N_1878,N_1680,N_1705);
and U1879 (N_1879,N_1609,N_1704);
or U1880 (N_1880,N_1681,N_1606);
or U1881 (N_1881,N_1761,N_1614);
nand U1882 (N_1882,N_1739,N_1650);
or U1883 (N_1883,N_1653,N_1789);
nand U1884 (N_1884,N_1667,N_1616);
nand U1885 (N_1885,N_1699,N_1798);
nand U1886 (N_1886,N_1660,N_1782);
or U1887 (N_1887,N_1674,N_1762);
or U1888 (N_1888,N_1683,N_1637);
nand U1889 (N_1889,N_1707,N_1626);
nor U1890 (N_1890,N_1607,N_1702);
nand U1891 (N_1891,N_1605,N_1769);
or U1892 (N_1892,N_1644,N_1629);
and U1893 (N_1893,N_1676,N_1608);
and U1894 (N_1894,N_1638,N_1657);
and U1895 (N_1895,N_1772,N_1727);
nand U1896 (N_1896,N_1754,N_1797);
or U1897 (N_1897,N_1649,N_1698);
nand U1898 (N_1898,N_1628,N_1753);
nand U1899 (N_1899,N_1701,N_1670);
xnor U1900 (N_1900,N_1655,N_1628);
nor U1901 (N_1901,N_1611,N_1716);
or U1902 (N_1902,N_1604,N_1718);
and U1903 (N_1903,N_1783,N_1645);
or U1904 (N_1904,N_1675,N_1604);
nand U1905 (N_1905,N_1605,N_1638);
nand U1906 (N_1906,N_1641,N_1693);
or U1907 (N_1907,N_1731,N_1615);
nand U1908 (N_1908,N_1607,N_1652);
nor U1909 (N_1909,N_1755,N_1737);
nand U1910 (N_1910,N_1673,N_1698);
and U1911 (N_1911,N_1725,N_1763);
nor U1912 (N_1912,N_1704,N_1786);
nand U1913 (N_1913,N_1624,N_1621);
xnor U1914 (N_1914,N_1757,N_1776);
and U1915 (N_1915,N_1787,N_1679);
and U1916 (N_1916,N_1743,N_1791);
and U1917 (N_1917,N_1652,N_1677);
and U1918 (N_1918,N_1625,N_1684);
nor U1919 (N_1919,N_1668,N_1639);
or U1920 (N_1920,N_1640,N_1688);
or U1921 (N_1921,N_1629,N_1759);
nand U1922 (N_1922,N_1622,N_1740);
nand U1923 (N_1923,N_1746,N_1706);
and U1924 (N_1924,N_1759,N_1683);
or U1925 (N_1925,N_1743,N_1776);
nor U1926 (N_1926,N_1655,N_1767);
and U1927 (N_1927,N_1737,N_1784);
nor U1928 (N_1928,N_1797,N_1666);
and U1929 (N_1929,N_1727,N_1612);
or U1930 (N_1930,N_1753,N_1777);
nor U1931 (N_1931,N_1705,N_1713);
or U1932 (N_1932,N_1708,N_1699);
or U1933 (N_1933,N_1724,N_1788);
and U1934 (N_1934,N_1744,N_1684);
nor U1935 (N_1935,N_1728,N_1656);
nor U1936 (N_1936,N_1701,N_1721);
and U1937 (N_1937,N_1627,N_1651);
nand U1938 (N_1938,N_1782,N_1690);
and U1939 (N_1939,N_1791,N_1766);
nor U1940 (N_1940,N_1686,N_1697);
and U1941 (N_1941,N_1635,N_1725);
nor U1942 (N_1942,N_1665,N_1771);
nand U1943 (N_1943,N_1760,N_1675);
nand U1944 (N_1944,N_1716,N_1706);
or U1945 (N_1945,N_1768,N_1791);
nor U1946 (N_1946,N_1760,N_1681);
and U1947 (N_1947,N_1770,N_1612);
nand U1948 (N_1948,N_1619,N_1781);
nand U1949 (N_1949,N_1646,N_1763);
and U1950 (N_1950,N_1764,N_1679);
and U1951 (N_1951,N_1664,N_1694);
nand U1952 (N_1952,N_1730,N_1614);
nor U1953 (N_1953,N_1610,N_1739);
nand U1954 (N_1954,N_1632,N_1726);
nand U1955 (N_1955,N_1696,N_1636);
and U1956 (N_1956,N_1702,N_1789);
and U1957 (N_1957,N_1631,N_1769);
nor U1958 (N_1958,N_1646,N_1724);
nor U1959 (N_1959,N_1719,N_1695);
nand U1960 (N_1960,N_1707,N_1652);
or U1961 (N_1961,N_1629,N_1645);
and U1962 (N_1962,N_1736,N_1756);
xnor U1963 (N_1963,N_1756,N_1793);
and U1964 (N_1964,N_1759,N_1782);
nor U1965 (N_1965,N_1735,N_1766);
and U1966 (N_1966,N_1633,N_1791);
and U1967 (N_1967,N_1629,N_1718);
nand U1968 (N_1968,N_1799,N_1751);
or U1969 (N_1969,N_1624,N_1627);
and U1970 (N_1970,N_1654,N_1675);
nor U1971 (N_1971,N_1748,N_1674);
and U1972 (N_1972,N_1679,N_1613);
nand U1973 (N_1973,N_1719,N_1792);
and U1974 (N_1974,N_1731,N_1739);
nand U1975 (N_1975,N_1730,N_1765);
nand U1976 (N_1976,N_1777,N_1613);
nor U1977 (N_1977,N_1713,N_1720);
nor U1978 (N_1978,N_1624,N_1654);
or U1979 (N_1979,N_1796,N_1757);
nor U1980 (N_1980,N_1623,N_1774);
nand U1981 (N_1981,N_1637,N_1730);
and U1982 (N_1982,N_1636,N_1629);
or U1983 (N_1983,N_1699,N_1640);
nand U1984 (N_1984,N_1770,N_1703);
and U1985 (N_1985,N_1704,N_1738);
nor U1986 (N_1986,N_1793,N_1664);
nand U1987 (N_1987,N_1604,N_1719);
and U1988 (N_1988,N_1790,N_1605);
nand U1989 (N_1989,N_1758,N_1770);
and U1990 (N_1990,N_1678,N_1772);
and U1991 (N_1991,N_1610,N_1789);
nand U1992 (N_1992,N_1724,N_1684);
xor U1993 (N_1993,N_1687,N_1740);
nand U1994 (N_1994,N_1653,N_1713);
nor U1995 (N_1995,N_1714,N_1723);
nor U1996 (N_1996,N_1739,N_1666);
nor U1997 (N_1997,N_1659,N_1604);
or U1998 (N_1998,N_1740,N_1708);
nand U1999 (N_1999,N_1645,N_1609);
nor U2000 (N_2000,N_1839,N_1891);
or U2001 (N_2001,N_1847,N_1994);
nand U2002 (N_2002,N_1889,N_1898);
nor U2003 (N_2003,N_1935,N_1834);
or U2004 (N_2004,N_1992,N_1915);
and U2005 (N_2005,N_1830,N_1993);
and U2006 (N_2006,N_1905,N_1972);
nand U2007 (N_2007,N_1958,N_1946);
nor U2008 (N_2008,N_1963,N_1996);
or U2009 (N_2009,N_1979,N_1883);
nand U2010 (N_2010,N_1916,N_1820);
and U2011 (N_2011,N_1838,N_1987);
and U2012 (N_2012,N_1878,N_1922);
and U2013 (N_2013,N_1876,N_1846);
or U2014 (N_2014,N_1999,N_1831);
and U2015 (N_2015,N_1814,N_1873);
and U2016 (N_2016,N_1908,N_1854);
nand U2017 (N_2017,N_1969,N_1892);
or U2018 (N_2018,N_1802,N_1800);
xnor U2019 (N_2019,N_1986,N_1909);
and U2020 (N_2020,N_1813,N_1938);
or U2021 (N_2021,N_1991,N_1936);
or U2022 (N_2022,N_1875,N_1869);
and U2023 (N_2023,N_1881,N_1983);
nand U2024 (N_2024,N_1807,N_1977);
nand U2025 (N_2025,N_1812,N_1928);
nand U2026 (N_2026,N_1921,N_1859);
or U2027 (N_2027,N_1947,N_1841);
nand U2028 (N_2028,N_1912,N_1966);
nand U2029 (N_2029,N_1903,N_1997);
nand U2030 (N_2030,N_1879,N_1937);
and U2031 (N_2031,N_1913,N_1801);
or U2032 (N_2032,N_1853,N_1957);
and U2033 (N_2033,N_1920,N_1871);
and U2034 (N_2034,N_1927,N_1811);
or U2035 (N_2035,N_1817,N_1819);
or U2036 (N_2036,N_1872,N_1944);
nor U2037 (N_2037,N_1925,N_1933);
and U2038 (N_2038,N_1941,N_1952);
nor U2039 (N_2039,N_1978,N_1924);
nor U2040 (N_2040,N_1899,N_1914);
and U2041 (N_2041,N_1990,N_1960);
nor U2042 (N_2042,N_1829,N_1852);
or U2043 (N_2043,N_1906,N_1860);
nand U2044 (N_2044,N_1967,N_1981);
nand U2045 (N_2045,N_1956,N_1953);
and U2046 (N_2046,N_1855,N_1858);
or U2047 (N_2047,N_1806,N_1955);
and U2048 (N_2048,N_1837,N_1850);
or U2049 (N_2049,N_1893,N_1917);
nor U2050 (N_2050,N_1880,N_1822);
nand U2051 (N_2051,N_1886,N_1882);
nor U2052 (N_2052,N_1929,N_1862);
nand U2053 (N_2053,N_1976,N_1942);
nor U2054 (N_2054,N_1919,N_1870);
nand U2055 (N_2055,N_1961,N_1931);
nand U2056 (N_2056,N_1836,N_1815);
and U2057 (N_2057,N_1932,N_1900);
nand U2058 (N_2058,N_1888,N_1902);
and U2059 (N_2059,N_1842,N_1845);
nand U2060 (N_2060,N_1864,N_1843);
or U2061 (N_2061,N_1840,N_1973);
xnor U2062 (N_2062,N_1894,N_1989);
nand U2063 (N_2063,N_1844,N_1975);
and U2064 (N_2064,N_1835,N_1911);
and U2065 (N_2065,N_1863,N_1988);
nand U2066 (N_2066,N_1849,N_1974);
nand U2067 (N_2067,N_1861,N_1887);
and U2068 (N_2068,N_1832,N_1965);
nand U2069 (N_2069,N_1985,N_1964);
or U2070 (N_2070,N_1874,N_1848);
nand U2071 (N_2071,N_1959,N_1810);
nand U2072 (N_2072,N_1901,N_1884);
nor U2073 (N_2073,N_1998,N_1950);
xnor U2074 (N_2074,N_1982,N_1904);
nand U2075 (N_2075,N_1803,N_1918);
and U2076 (N_2076,N_1808,N_1926);
and U2077 (N_2077,N_1968,N_1867);
and U2078 (N_2078,N_1823,N_1949);
nand U2079 (N_2079,N_1907,N_1827);
nor U2080 (N_2080,N_1825,N_1954);
and U2081 (N_2081,N_1865,N_1948);
nand U2082 (N_2082,N_1856,N_1962);
nor U2083 (N_2083,N_1877,N_1833);
nand U2084 (N_2084,N_1857,N_1940);
and U2085 (N_2085,N_1818,N_1809);
or U2086 (N_2086,N_1930,N_1945);
nor U2087 (N_2087,N_1910,N_1805);
nand U2088 (N_2088,N_1866,N_1934);
or U2089 (N_2089,N_1851,N_1896);
and U2090 (N_2090,N_1885,N_1826);
nand U2091 (N_2091,N_1895,N_1868);
nand U2092 (N_2092,N_1984,N_1951);
and U2093 (N_2093,N_1970,N_1943);
nor U2094 (N_2094,N_1980,N_1897);
or U2095 (N_2095,N_1804,N_1890);
nand U2096 (N_2096,N_1816,N_1995);
and U2097 (N_2097,N_1923,N_1971);
nor U2098 (N_2098,N_1939,N_1828);
nor U2099 (N_2099,N_1821,N_1824);
and U2100 (N_2100,N_1810,N_1873);
nor U2101 (N_2101,N_1905,N_1934);
nor U2102 (N_2102,N_1927,N_1878);
or U2103 (N_2103,N_1858,N_1857);
nor U2104 (N_2104,N_1884,N_1931);
or U2105 (N_2105,N_1918,N_1814);
and U2106 (N_2106,N_1959,N_1866);
or U2107 (N_2107,N_1927,N_1864);
and U2108 (N_2108,N_1810,N_1831);
nor U2109 (N_2109,N_1965,N_1834);
and U2110 (N_2110,N_1910,N_1810);
nand U2111 (N_2111,N_1934,N_1878);
and U2112 (N_2112,N_1952,N_1970);
or U2113 (N_2113,N_1806,N_1924);
or U2114 (N_2114,N_1902,N_1848);
nand U2115 (N_2115,N_1953,N_1862);
or U2116 (N_2116,N_1842,N_1835);
nand U2117 (N_2117,N_1902,N_1891);
or U2118 (N_2118,N_1801,N_1949);
nand U2119 (N_2119,N_1953,N_1950);
and U2120 (N_2120,N_1922,N_1975);
nor U2121 (N_2121,N_1871,N_1840);
nor U2122 (N_2122,N_1886,N_1893);
nor U2123 (N_2123,N_1907,N_1997);
nor U2124 (N_2124,N_1935,N_1887);
or U2125 (N_2125,N_1963,N_1829);
or U2126 (N_2126,N_1969,N_1809);
nand U2127 (N_2127,N_1960,N_1864);
nand U2128 (N_2128,N_1981,N_1829);
nor U2129 (N_2129,N_1862,N_1985);
nand U2130 (N_2130,N_1833,N_1991);
nor U2131 (N_2131,N_1934,N_1871);
and U2132 (N_2132,N_1829,N_1822);
nor U2133 (N_2133,N_1858,N_1853);
and U2134 (N_2134,N_1951,N_1956);
nor U2135 (N_2135,N_1960,N_1845);
nand U2136 (N_2136,N_1904,N_1952);
or U2137 (N_2137,N_1926,N_1943);
nor U2138 (N_2138,N_1929,N_1955);
nand U2139 (N_2139,N_1902,N_1837);
and U2140 (N_2140,N_1970,N_1947);
nor U2141 (N_2141,N_1893,N_1919);
nor U2142 (N_2142,N_1800,N_1849);
nor U2143 (N_2143,N_1940,N_1946);
and U2144 (N_2144,N_1853,N_1913);
or U2145 (N_2145,N_1892,N_1863);
or U2146 (N_2146,N_1992,N_1876);
nand U2147 (N_2147,N_1836,N_1998);
and U2148 (N_2148,N_1990,N_1999);
nor U2149 (N_2149,N_1834,N_1879);
nor U2150 (N_2150,N_1868,N_1944);
nor U2151 (N_2151,N_1855,N_1937);
nand U2152 (N_2152,N_1967,N_1936);
nor U2153 (N_2153,N_1875,N_1823);
nand U2154 (N_2154,N_1850,N_1939);
and U2155 (N_2155,N_1911,N_1840);
and U2156 (N_2156,N_1991,N_1921);
and U2157 (N_2157,N_1936,N_1973);
nor U2158 (N_2158,N_1888,N_1952);
and U2159 (N_2159,N_1938,N_1948);
nor U2160 (N_2160,N_1986,N_1879);
or U2161 (N_2161,N_1890,N_1994);
nand U2162 (N_2162,N_1992,N_1849);
and U2163 (N_2163,N_1940,N_1870);
nand U2164 (N_2164,N_1982,N_1956);
or U2165 (N_2165,N_1988,N_1959);
nor U2166 (N_2166,N_1851,N_1806);
nor U2167 (N_2167,N_1896,N_1821);
and U2168 (N_2168,N_1999,N_1929);
nand U2169 (N_2169,N_1963,N_1864);
nand U2170 (N_2170,N_1997,N_1865);
and U2171 (N_2171,N_1861,N_1841);
nand U2172 (N_2172,N_1999,N_1924);
and U2173 (N_2173,N_1982,N_1860);
or U2174 (N_2174,N_1907,N_1931);
or U2175 (N_2175,N_1922,N_1813);
nand U2176 (N_2176,N_1858,N_1808);
nor U2177 (N_2177,N_1914,N_1851);
nand U2178 (N_2178,N_1945,N_1964);
nor U2179 (N_2179,N_1957,N_1841);
or U2180 (N_2180,N_1833,N_1883);
and U2181 (N_2181,N_1800,N_1985);
nor U2182 (N_2182,N_1808,N_1853);
nand U2183 (N_2183,N_1824,N_1948);
or U2184 (N_2184,N_1863,N_1855);
nor U2185 (N_2185,N_1990,N_1923);
and U2186 (N_2186,N_1973,N_1953);
nand U2187 (N_2187,N_1914,N_1940);
or U2188 (N_2188,N_1994,N_1897);
or U2189 (N_2189,N_1965,N_1879);
nor U2190 (N_2190,N_1921,N_1848);
nor U2191 (N_2191,N_1808,N_1800);
nor U2192 (N_2192,N_1951,N_1824);
nand U2193 (N_2193,N_1808,N_1939);
or U2194 (N_2194,N_1962,N_1914);
nand U2195 (N_2195,N_1947,N_1920);
or U2196 (N_2196,N_1905,N_1807);
and U2197 (N_2197,N_1851,N_1869);
or U2198 (N_2198,N_1993,N_1955);
or U2199 (N_2199,N_1953,N_1876);
nand U2200 (N_2200,N_2154,N_2070);
nor U2201 (N_2201,N_2043,N_2026);
nor U2202 (N_2202,N_2149,N_2041);
or U2203 (N_2203,N_2045,N_2105);
nand U2204 (N_2204,N_2151,N_2012);
and U2205 (N_2205,N_2058,N_2034);
or U2206 (N_2206,N_2093,N_2004);
nor U2207 (N_2207,N_2096,N_2089);
nor U2208 (N_2208,N_2003,N_2082);
nand U2209 (N_2209,N_2115,N_2141);
nand U2210 (N_2210,N_2170,N_2106);
nor U2211 (N_2211,N_2165,N_2114);
or U2212 (N_2212,N_2128,N_2021);
nand U2213 (N_2213,N_2052,N_2168);
or U2214 (N_2214,N_2131,N_2077);
and U2215 (N_2215,N_2173,N_2116);
and U2216 (N_2216,N_2076,N_2123);
nand U2217 (N_2217,N_2179,N_2010);
nor U2218 (N_2218,N_2140,N_2056);
nor U2219 (N_2219,N_2002,N_2008);
or U2220 (N_2220,N_2142,N_2192);
nor U2221 (N_2221,N_2175,N_2118);
nand U2222 (N_2222,N_2135,N_2157);
nor U2223 (N_2223,N_2074,N_2100);
nand U2224 (N_2224,N_2150,N_2036);
or U2225 (N_2225,N_2022,N_2065);
and U2226 (N_2226,N_2174,N_2028);
nand U2227 (N_2227,N_2144,N_2018);
and U2228 (N_2228,N_2049,N_2068);
nor U2229 (N_2229,N_2094,N_2067);
nor U2230 (N_2230,N_2199,N_2009);
nor U2231 (N_2231,N_2129,N_2148);
nand U2232 (N_2232,N_2006,N_2062);
xnor U2233 (N_2233,N_2011,N_2042);
nand U2234 (N_2234,N_2095,N_2098);
and U2235 (N_2235,N_2088,N_2153);
xor U2236 (N_2236,N_2120,N_2103);
and U2237 (N_2237,N_2104,N_2017);
nor U2238 (N_2238,N_2015,N_2160);
nand U2239 (N_2239,N_2184,N_2187);
nor U2240 (N_2240,N_2000,N_2081);
nor U2241 (N_2241,N_2112,N_2057);
xnor U2242 (N_2242,N_2127,N_2145);
xor U2243 (N_2243,N_2078,N_2169);
or U2244 (N_2244,N_2124,N_2064);
nor U2245 (N_2245,N_2066,N_2090);
nor U2246 (N_2246,N_2134,N_2029);
and U2247 (N_2247,N_2055,N_2047);
nand U2248 (N_2248,N_2063,N_2189);
or U2249 (N_2249,N_2044,N_2117);
nand U2250 (N_2250,N_2176,N_2019);
and U2251 (N_2251,N_2059,N_2024);
nand U2252 (N_2252,N_2001,N_2137);
or U2253 (N_2253,N_2087,N_2183);
nand U2254 (N_2254,N_2158,N_2014);
nand U2255 (N_2255,N_2113,N_2069);
nor U2256 (N_2256,N_2193,N_2188);
nand U2257 (N_2257,N_2198,N_2121);
nor U2258 (N_2258,N_2166,N_2091);
or U2259 (N_2259,N_2023,N_2185);
nand U2260 (N_2260,N_2111,N_2092);
nor U2261 (N_2261,N_2037,N_2025);
nor U2262 (N_2262,N_2030,N_2099);
nand U2263 (N_2263,N_2152,N_2051);
nor U2264 (N_2264,N_2050,N_2107);
and U2265 (N_2265,N_2110,N_2083);
and U2266 (N_2266,N_2180,N_2155);
or U2267 (N_2267,N_2054,N_2138);
or U2268 (N_2268,N_2143,N_2162);
or U2269 (N_2269,N_2147,N_2194);
nand U2270 (N_2270,N_2119,N_2164);
or U2271 (N_2271,N_2102,N_2146);
and U2272 (N_2272,N_2005,N_2039);
or U2273 (N_2273,N_2080,N_2053);
nor U2274 (N_2274,N_2177,N_2060);
nand U2275 (N_2275,N_2033,N_2172);
or U2276 (N_2276,N_2126,N_2084);
and U2277 (N_2277,N_2061,N_2073);
or U2278 (N_2278,N_2032,N_2156);
nor U2279 (N_2279,N_2132,N_2136);
or U2280 (N_2280,N_2020,N_2159);
xor U2281 (N_2281,N_2040,N_2182);
or U2282 (N_2282,N_2196,N_2130);
or U2283 (N_2283,N_2161,N_2197);
and U2284 (N_2284,N_2072,N_2101);
nand U2285 (N_2285,N_2038,N_2027);
nand U2286 (N_2286,N_2016,N_2186);
nand U2287 (N_2287,N_2122,N_2190);
and U2288 (N_2288,N_2048,N_2046);
nor U2289 (N_2289,N_2108,N_2031);
nor U2290 (N_2290,N_2163,N_2035);
or U2291 (N_2291,N_2075,N_2133);
nand U2292 (N_2292,N_2125,N_2178);
or U2293 (N_2293,N_2007,N_2109);
nand U2294 (N_2294,N_2071,N_2171);
nand U2295 (N_2295,N_2079,N_2086);
and U2296 (N_2296,N_2191,N_2181);
nand U2297 (N_2297,N_2167,N_2097);
and U2298 (N_2298,N_2085,N_2139);
or U2299 (N_2299,N_2013,N_2195);
and U2300 (N_2300,N_2105,N_2019);
nand U2301 (N_2301,N_2021,N_2196);
or U2302 (N_2302,N_2106,N_2145);
nor U2303 (N_2303,N_2082,N_2005);
nor U2304 (N_2304,N_2023,N_2137);
nand U2305 (N_2305,N_2074,N_2166);
or U2306 (N_2306,N_2025,N_2001);
nand U2307 (N_2307,N_2131,N_2151);
and U2308 (N_2308,N_2034,N_2169);
nand U2309 (N_2309,N_2012,N_2184);
nor U2310 (N_2310,N_2034,N_2009);
or U2311 (N_2311,N_2198,N_2133);
or U2312 (N_2312,N_2173,N_2059);
or U2313 (N_2313,N_2182,N_2075);
or U2314 (N_2314,N_2104,N_2047);
and U2315 (N_2315,N_2023,N_2168);
nand U2316 (N_2316,N_2166,N_2048);
nand U2317 (N_2317,N_2199,N_2133);
nor U2318 (N_2318,N_2012,N_2018);
nor U2319 (N_2319,N_2179,N_2037);
or U2320 (N_2320,N_2149,N_2030);
nand U2321 (N_2321,N_2005,N_2037);
and U2322 (N_2322,N_2150,N_2019);
nor U2323 (N_2323,N_2007,N_2132);
or U2324 (N_2324,N_2094,N_2080);
nand U2325 (N_2325,N_2134,N_2157);
nor U2326 (N_2326,N_2125,N_2037);
or U2327 (N_2327,N_2117,N_2166);
or U2328 (N_2328,N_2084,N_2059);
or U2329 (N_2329,N_2159,N_2096);
and U2330 (N_2330,N_2144,N_2083);
or U2331 (N_2331,N_2071,N_2100);
or U2332 (N_2332,N_2162,N_2001);
nor U2333 (N_2333,N_2045,N_2059);
and U2334 (N_2334,N_2061,N_2110);
and U2335 (N_2335,N_2046,N_2065);
nor U2336 (N_2336,N_2073,N_2105);
nand U2337 (N_2337,N_2077,N_2196);
nor U2338 (N_2338,N_2086,N_2161);
or U2339 (N_2339,N_2059,N_2021);
xor U2340 (N_2340,N_2096,N_2015);
nor U2341 (N_2341,N_2071,N_2128);
and U2342 (N_2342,N_2174,N_2103);
nor U2343 (N_2343,N_2141,N_2096);
and U2344 (N_2344,N_2066,N_2177);
nor U2345 (N_2345,N_2166,N_2101);
nand U2346 (N_2346,N_2041,N_2083);
and U2347 (N_2347,N_2072,N_2074);
nand U2348 (N_2348,N_2182,N_2124);
or U2349 (N_2349,N_2045,N_2176);
nor U2350 (N_2350,N_2008,N_2050);
nand U2351 (N_2351,N_2088,N_2082);
nand U2352 (N_2352,N_2167,N_2159);
and U2353 (N_2353,N_2001,N_2079);
or U2354 (N_2354,N_2029,N_2062);
or U2355 (N_2355,N_2122,N_2185);
or U2356 (N_2356,N_2133,N_2048);
and U2357 (N_2357,N_2107,N_2112);
nor U2358 (N_2358,N_2196,N_2054);
nor U2359 (N_2359,N_2090,N_2157);
nand U2360 (N_2360,N_2121,N_2181);
and U2361 (N_2361,N_2121,N_2117);
and U2362 (N_2362,N_2117,N_2081);
nand U2363 (N_2363,N_2098,N_2086);
or U2364 (N_2364,N_2136,N_2055);
nand U2365 (N_2365,N_2072,N_2097);
nand U2366 (N_2366,N_2121,N_2038);
xnor U2367 (N_2367,N_2051,N_2075);
and U2368 (N_2368,N_2108,N_2198);
or U2369 (N_2369,N_2041,N_2158);
or U2370 (N_2370,N_2009,N_2100);
nand U2371 (N_2371,N_2132,N_2104);
and U2372 (N_2372,N_2141,N_2087);
or U2373 (N_2373,N_2124,N_2021);
nand U2374 (N_2374,N_2093,N_2118);
nor U2375 (N_2375,N_2195,N_2014);
nor U2376 (N_2376,N_2109,N_2133);
or U2377 (N_2377,N_2013,N_2182);
nand U2378 (N_2378,N_2067,N_2119);
nor U2379 (N_2379,N_2057,N_2086);
nand U2380 (N_2380,N_2089,N_2033);
or U2381 (N_2381,N_2087,N_2093);
and U2382 (N_2382,N_2127,N_2000);
nor U2383 (N_2383,N_2026,N_2075);
or U2384 (N_2384,N_2092,N_2048);
xor U2385 (N_2385,N_2005,N_2129);
and U2386 (N_2386,N_2085,N_2144);
nand U2387 (N_2387,N_2173,N_2041);
or U2388 (N_2388,N_2086,N_2142);
and U2389 (N_2389,N_2041,N_2127);
or U2390 (N_2390,N_2000,N_2099);
nand U2391 (N_2391,N_2164,N_2081);
nand U2392 (N_2392,N_2094,N_2114);
nand U2393 (N_2393,N_2062,N_2076);
nand U2394 (N_2394,N_2053,N_2006);
nor U2395 (N_2395,N_2107,N_2174);
or U2396 (N_2396,N_2060,N_2063);
xnor U2397 (N_2397,N_2006,N_2085);
nand U2398 (N_2398,N_2028,N_2173);
or U2399 (N_2399,N_2018,N_2110);
or U2400 (N_2400,N_2263,N_2324);
or U2401 (N_2401,N_2309,N_2251);
or U2402 (N_2402,N_2257,N_2276);
nand U2403 (N_2403,N_2303,N_2348);
nor U2404 (N_2404,N_2218,N_2374);
nand U2405 (N_2405,N_2329,N_2349);
nand U2406 (N_2406,N_2397,N_2335);
nor U2407 (N_2407,N_2331,N_2394);
and U2408 (N_2408,N_2298,N_2295);
nand U2409 (N_2409,N_2302,N_2314);
nand U2410 (N_2410,N_2236,N_2287);
nor U2411 (N_2411,N_2339,N_2215);
nand U2412 (N_2412,N_2344,N_2270);
nand U2413 (N_2413,N_2212,N_2360);
and U2414 (N_2414,N_2227,N_2375);
and U2415 (N_2415,N_2203,N_2352);
xnor U2416 (N_2416,N_2201,N_2376);
nand U2417 (N_2417,N_2363,N_2357);
nor U2418 (N_2418,N_2272,N_2209);
nor U2419 (N_2419,N_2225,N_2387);
and U2420 (N_2420,N_2299,N_2249);
nand U2421 (N_2421,N_2328,N_2350);
and U2422 (N_2422,N_2278,N_2305);
and U2423 (N_2423,N_2318,N_2234);
and U2424 (N_2424,N_2356,N_2213);
nor U2425 (N_2425,N_2208,N_2355);
nand U2426 (N_2426,N_2260,N_2346);
and U2427 (N_2427,N_2381,N_2285);
nor U2428 (N_2428,N_2241,N_2300);
nor U2429 (N_2429,N_2223,N_2222);
and U2430 (N_2430,N_2367,N_2268);
or U2431 (N_2431,N_2281,N_2231);
nand U2432 (N_2432,N_2221,N_2229);
or U2433 (N_2433,N_2271,N_2320);
and U2434 (N_2434,N_2366,N_2254);
or U2435 (N_2435,N_2313,N_2341);
and U2436 (N_2436,N_2390,N_2330);
and U2437 (N_2437,N_2351,N_2343);
nor U2438 (N_2438,N_2258,N_2286);
nor U2439 (N_2439,N_2277,N_2382);
or U2440 (N_2440,N_2217,N_2373);
and U2441 (N_2441,N_2396,N_2392);
or U2442 (N_2442,N_2284,N_2274);
or U2443 (N_2443,N_2290,N_2383);
and U2444 (N_2444,N_2380,N_2315);
nand U2445 (N_2445,N_2202,N_2399);
nor U2446 (N_2446,N_2235,N_2368);
or U2447 (N_2447,N_2369,N_2243);
and U2448 (N_2448,N_2311,N_2325);
or U2449 (N_2449,N_2259,N_2322);
nand U2450 (N_2450,N_2389,N_2306);
nor U2451 (N_2451,N_2266,N_2354);
or U2452 (N_2452,N_2280,N_2279);
nand U2453 (N_2453,N_2245,N_2326);
and U2454 (N_2454,N_2395,N_2207);
nor U2455 (N_2455,N_2321,N_2388);
and U2456 (N_2456,N_2247,N_2301);
nor U2457 (N_2457,N_2293,N_2333);
nor U2458 (N_2458,N_2214,N_2262);
and U2459 (N_2459,N_2398,N_2359);
nor U2460 (N_2460,N_2307,N_2246);
nand U2461 (N_2461,N_2228,N_2233);
nor U2462 (N_2462,N_2255,N_2216);
and U2463 (N_2463,N_2283,N_2219);
and U2464 (N_2464,N_2248,N_2204);
and U2465 (N_2465,N_2224,N_2345);
and U2466 (N_2466,N_2261,N_2265);
nand U2467 (N_2467,N_2338,N_2361);
and U2468 (N_2468,N_2364,N_2379);
nor U2469 (N_2469,N_2317,N_2294);
and U2470 (N_2470,N_2362,N_2353);
and U2471 (N_2471,N_2372,N_2312);
nor U2472 (N_2472,N_2342,N_2253);
xnor U2473 (N_2473,N_2291,N_2347);
nand U2474 (N_2474,N_2240,N_2340);
xnor U2475 (N_2475,N_2337,N_2316);
nor U2476 (N_2476,N_2365,N_2358);
nor U2477 (N_2477,N_2211,N_2242);
nand U2478 (N_2478,N_2206,N_2250);
xor U2479 (N_2479,N_2289,N_2297);
xor U2480 (N_2480,N_2282,N_2273);
xnor U2481 (N_2481,N_2336,N_2378);
xor U2482 (N_2482,N_2220,N_2238);
nand U2483 (N_2483,N_2230,N_2232);
nand U2484 (N_2484,N_2205,N_2327);
or U2485 (N_2485,N_2385,N_2296);
nand U2486 (N_2486,N_2264,N_2391);
nor U2487 (N_2487,N_2332,N_2239);
nand U2488 (N_2488,N_2226,N_2384);
or U2489 (N_2489,N_2323,N_2393);
or U2490 (N_2490,N_2334,N_2377);
and U2491 (N_2491,N_2256,N_2244);
or U2492 (N_2492,N_2308,N_2319);
or U2493 (N_2493,N_2371,N_2292);
nor U2494 (N_2494,N_2269,N_2267);
nand U2495 (N_2495,N_2275,N_2200);
nor U2496 (N_2496,N_2210,N_2386);
nor U2497 (N_2497,N_2370,N_2304);
nor U2498 (N_2498,N_2252,N_2288);
nand U2499 (N_2499,N_2237,N_2310);
nand U2500 (N_2500,N_2350,N_2310);
xor U2501 (N_2501,N_2338,N_2318);
and U2502 (N_2502,N_2284,N_2251);
xor U2503 (N_2503,N_2202,N_2335);
and U2504 (N_2504,N_2369,N_2261);
nor U2505 (N_2505,N_2305,N_2287);
nand U2506 (N_2506,N_2263,N_2373);
and U2507 (N_2507,N_2249,N_2396);
nor U2508 (N_2508,N_2224,N_2310);
nand U2509 (N_2509,N_2336,N_2358);
and U2510 (N_2510,N_2249,N_2284);
nand U2511 (N_2511,N_2210,N_2326);
and U2512 (N_2512,N_2245,N_2225);
nor U2513 (N_2513,N_2320,N_2313);
nand U2514 (N_2514,N_2277,N_2361);
or U2515 (N_2515,N_2372,N_2385);
or U2516 (N_2516,N_2218,N_2397);
nand U2517 (N_2517,N_2222,N_2394);
or U2518 (N_2518,N_2328,N_2356);
nand U2519 (N_2519,N_2332,N_2382);
and U2520 (N_2520,N_2202,N_2384);
and U2521 (N_2521,N_2279,N_2298);
nor U2522 (N_2522,N_2280,N_2313);
nor U2523 (N_2523,N_2358,N_2327);
nor U2524 (N_2524,N_2373,N_2330);
and U2525 (N_2525,N_2325,N_2259);
nor U2526 (N_2526,N_2298,N_2339);
and U2527 (N_2527,N_2345,N_2257);
or U2528 (N_2528,N_2206,N_2387);
or U2529 (N_2529,N_2366,N_2243);
and U2530 (N_2530,N_2343,N_2315);
and U2531 (N_2531,N_2311,N_2277);
or U2532 (N_2532,N_2362,N_2283);
nand U2533 (N_2533,N_2278,N_2376);
nand U2534 (N_2534,N_2216,N_2317);
nand U2535 (N_2535,N_2322,N_2302);
nand U2536 (N_2536,N_2398,N_2380);
and U2537 (N_2537,N_2237,N_2324);
nand U2538 (N_2538,N_2339,N_2237);
and U2539 (N_2539,N_2327,N_2379);
and U2540 (N_2540,N_2213,N_2226);
or U2541 (N_2541,N_2312,N_2394);
nand U2542 (N_2542,N_2205,N_2325);
or U2543 (N_2543,N_2374,N_2207);
nor U2544 (N_2544,N_2356,N_2327);
nand U2545 (N_2545,N_2355,N_2261);
nor U2546 (N_2546,N_2215,N_2245);
xor U2547 (N_2547,N_2390,N_2380);
nor U2548 (N_2548,N_2259,N_2215);
xnor U2549 (N_2549,N_2217,N_2396);
and U2550 (N_2550,N_2309,N_2234);
nor U2551 (N_2551,N_2226,N_2221);
and U2552 (N_2552,N_2360,N_2279);
or U2553 (N_2553,N_2231,N_2391);
and U2554 (N_2554,N_2268,N_2249);
and U2555 (N_2555,N_2247,N_2210);
nor U2556 (N_2556,N_2358,N_2299);
or U2557 (N_2557,N_2388,N_2242);
nor U2558 (N_2558,N_2326,N_2337);
nor U2559 (N_2559,N_2347,N_2251);
nand U2560 (N_2560,N_2273,N_2391);
nand U2561 (N_2561,N_2304,N_2384);
nor U2562 (N_2562,N_2280,N_2217);
nor U2563 (N_2563,N_2204,N_2236);
or U2564 (N_2564,N_2248,N_2337);
xnor U2565 (N_2565,N_2330,N_2227);
nand U2566 (N_2566,N_2344,N_2368);
nand U2567 (N_2567,N_2311,N_2262);
nand U2568 (N_2568,N_2279,N_2214);
nand U2569 (N_2569,N_2394,N_2256);
or U2570 (N_2570,N_2234,N_2235);
and U2571 (N_2571,N_2352,N_2379);
or U2572 (N_2572,N_2273,N_2336);
nand U2573 (N_2573,N_2314,N_2254);
or U2574 (N_2574,N_2234,N_2272);
nand U2575 (N_2575,N_2333,N_2339);
nand U2576 (N_2576,N_2202,N_2242);
nand U2577 (N_2577,N_2333,N_2251);
or U2578 (N_2578,N_2365,N_2282);
or U2579 (N_2579,N_2280,N_2329);
and U2580 (N_2580,N_2359,N_2262);
nand U2581 (N_2581,N_2291,N_2343);
nor U2582 (N_2582,N_2257,N_2250);
and U2583 (N_2583,N_2361,N_2208);
and U2584 (N_2584,N_2396,N_2272);
nor U2585 (N_2585,N_2369,N_2327);
nor U2586 (N_2586,N_2257,N_2287);
or U2587 (N_2587,N_2341,N_2254);
or U2588 (N_2588,N_2240,N_2276);
xor U2589 (N_2589,N_2361,N_2239);
or U2590 (N_2590,N_2214,N_2309);
nor U2591 (N_2591,N_2378,N_2363);
and U2592 (N_2592,N_2211,N_2269);
nand U2593 (N_2593,N_2340,N_2396);
nor U2594 (N_2594,N_2323,N_2360);
or U2595 (N_2595,N_2291,N_2398);
or U2596 (N_2596,N_2272,N_2319);
nor U2597 (N_2597,N_2375,N_2200);
or U2598 (N_2598,N_2206,N_2265);
nand U2599 (N_2599,N_2248,N_2354);
or U2600 (N_2600,N_2520,N_2524);
and U2601 (N_2601,N_2424,N_2510);
or U2602 (N_2602,N_2415,N_2571);
nand U2603 (N_2603,N_2581,N_2432);
or U2604 (N_2604,N_2474,N_2428);
nor U2605 (N_2605,N_2501,N_2537);
nor U2606 (N_2606,N_2549,N_2542);
nand U2607 (N_2607,N_2497,N_2412);
nor U2608 (N_2608,N_2489,N_2484);
and U2609 (N_2609,N_2465,N_2503);
nand U2610 (N_2610,N_2512,N_2461);
and U2611 (N_2611,N_2414,N_2429);
and U2612 (N_2612,N_2403,N_2554);
or U2613 (N_2613,N_2586,N_2491);
nand U2614 (N_2614,N_2444,N_2529);
nand U2615 (N_2615,N_2580,N_2570);
or U2616 (N_2616,N_2443,N_2599);
nor U2617 (N_2617,N_2453,N_2557);
or U2618 (N_2618,N_2454,N_2540);
or U2619 (N_2619,N_2583,N_2508);
and U2620 (N_2620,N_2456,N_2413);
nor U2621 (N_2621,N_2574,N_2544);
or U2622 (N_2622,N_2595,N_2452);
nand U2623 (N_2623,N_2506,N_2566);
nor U2624 (N_2624,N_2502,N_2430);
and U2625 (N_2625,N_2499,N_2558);
and U2626 (N_2626,N_2597,N_2483);
nor U2627 (N_2627,N_2553,N_2400);
nor U2628 (N_2628,N_2539,N_2417);
or U2629 (N_2629,N_2561,N_2578);
nand U2630 (N_2630,N_2492,N_2434);
nand U2631 (N_2631,N_2589,N_2500);
or U2632 (N_2632,N_2446,N_2593);
and U2633 (N_2633,N_2402,N_2547);
or U2634 (N_2634,N_2528,N_2556);
or U2635 (N_2635,N_2555,N_2479);
nand U2636 (N_2636,N_2573,N_2419);
or U2637 (N_2637,N_2533,N_2538);
xor U2638 (N_2638,N_2598,N_2447);
nand U2639 (N_2639,N_2587,N_2523);
or U2640 (N_2640,N_2433,N_2439);
nor U2641 (N_2641,N_2449,N_2463);
or U2642 (N_2642,N_2468,N_2577);
and U2643 (N_2643,N_2584,N_2420);
and U2644 (N_2644,N_2585,N_2478);
and U2645 (N_2645,N_2576,N_2519);
nor U2646 (N_2646,N_2511,N_2427);
nand U2647 (N_2647,N_2460,N_2592);
and U2648 (N_2648,N_2441,N_2477);
and U2649 (N_2649,N_2480,N_2548);
and U2650 (N_2650,N_2564,N_2550);
and U2651 (N_2651,N_2559,N_2409);
or U2652 (N_2652,N_2466,N_2481);
and U2653 (N_2653,N_2493,N_2525);
nand U2654 (N_2654,N_2515,N_2521);
nor U2655 (N_2655,N_2445,N_2567);
or U2656 (N_2656,N_2488,N_2536);
nand U2657 (N_2657,N_2563,N_2437);
and U2658 (N_2658,N_2575,N_2591);
nor U2659 (N_2659,N_2572,N_2535);
or U2660 (N_2660,N_2459,N_2408);
nor U2661 (N_2661,N_2457,N_2467);
nor U2662 (N_2662,N_2440,N_2534);
and U2663 (N_2663,N_2464,N_2405);
or U2664 (N_2664,N_2531,N_2494);
and U2665 (N_2665,N_2543,N_2516);
nor U2666 (N_2666,N_2490,N_2487);
and U2667 (N_2667,N_2579,N_2410);
and U2668 (N_2668,N_2552,N_2513);
nor U2669 (N_2669,N_2406,N_2518);
or U2670 (N_2670,N_2482,N_2426);
and U2671 (N_2671,N_2562,N_2435);
or U2672 (N_2672,N_2423,N_2507);
xnor U2673 (N_2673,N_2401,N_2569);
nor U2674 (N_2674,N_2458,N_2404);
or U2675 (N_2675,N_2568,N_2451);
xor U2676 (N_2676,N_2588,N_2407);
nand U2677 (N_2677,N_2517,N_2473);
and U2678 (N_2678,N_2530,N_2496);
and U2679 (N_2679,N_2545,N_2495);
or U2680 (N_2680,N_2475,N_2436);
nor U2681 (N_2681,N_2425,N_2442);
and U2682 (N_2682,N_2527,N_2470);
nor U2683 (N_2683,N_2438,N_2431);
nor U2684 (N_2684,N_2514,N_2469);
and U2685 (N_2685,N_2596,N_2504);
nand U2686 (N_2686,N_2421,N_2416);
nor U2687 (N_2687,N_2486,N_2594);
and U2688 (N_2688,N_2565,N_2560);
nand U2689 (N_2689,N_2472,N_2462);
nor U2690 (N_2690,N_2418,N_2532);
and U2691 (N_2691,N_2541,N_2582);
or U2692 (N_2692,N_2509,N_2450);
or U2693 (N_2693,N_2448,N_2422);
or U2694 (N_2694,N_2546,N_2590);
nor U2695 (N_2695,N_2476,N_2455);
nand U2696 (N_2696,N_2551,N_2498);
or U2697 (N_2697,N_2411,N_2485);
nor U2698 (N_2698,N_2526,N_2471);
xor U2699 (N_2699,N_2505,N_2522);
and U2700 (N_2700,N_2454,N_2574);
nand U2701 (N_2701,N_2532,N_2470);
nand U2702 (N_2702,N_2546,N_2522);
nand U2703 (N_2703,N_2418,N_2588);
nand U2704 (N_2704,N_2535,N_2560);
nor U2705 (N_2705,N_2560,N_2495);
or U2706 (N_2706,N_2414,N_2464);
and U2707 (N_2707,N_2529,N_2499);
or U2708 (N_2708,N_2542,N_2598);
xnor U2709 (N_2709,N_2461,N_2535);
or U2710 (N_2710,N_2438,N_2481);
or U2711 (N_2711,N_2450,N_2495);
nor U2712 (N_2712,N_2558,N_2440);
or U2713 (N_2713,N_2574,N_2565);
or U2714 (N_2714,N_2586,N_2455);
nand U2715 (N_2715,N_2551,N_2582);
nand U2716 (N_2716,N_2568,N_2498);
or U2717 (N_2717,N_2560,N_2555);
xnor U2718 (N_2718,N_2535,N_2446);
and U2719 (N_2719,N_2475,N_2400);
nor U2720 (N_2720,N_2452,N_2589);
or U2721 (N_2721,N_2443,N_2530);
nand U2722 (N_2722,N_2545,N_2423);
nor U2723 (N_2723,N_2511,N_2459);
nand U2724 (N_2724,N_2447,N_2554);
nand U2725 (N_2725,N_2568,N_2424);
nand U2726 (N_2726,N_2565,N_2463);
or U2727 (N_2727,N_2472,N_2554);
nand U2728 (N_2728,N_2547,N_2558);
nand U2729 (N_2729,N_2478,N_2417);
nor U2730 (N_2730,N_2453,N_2496);
or U2731 (N_2731,N_2580,N_2490);
nor U2732 (N_2732,N_2460,N_2421);
nand U2733 (N_2733,N_2505,N_2405);
or U2734 (N_2734,N_2528,N_2420);
and U2735 (N_2735,N_2436,N_2529);
nor U2736 (N_2736,N_2424,N_2579);
nand U2737 (N_2737,N_2493,N_2579);
or U2738 (N_2738,N_2472,N_2533);
or U2739 (N_2739,N_2417,N_2497);
or U2740 (N_2740,N_2424,N_2468);
nor U2741 (N_2741,N_2568,N_2519);
or U2742 (N_2742,N_2506,N_2593);
nor U2743 (N_2743,N_2474,N_2519);
or U2744 (N_2744,N_2476,N_2543);
and U2745 (N_2745,N_2569,N_2435);
and U2746 (N_2746,N_2573,N_2534);
nor U2747 (N_2747,N_2414,N_2501);
xnor U2748 (N_2748,N_2491,N_2559);
nand U2749 (N_2749,N_2434,N_2401);
and U2750 (N_2750,N_2584,N_2434);
nand U2751 (N_2751,N_2592,N_2479);
nor U2752 (N_2752,N_2570,N_2542);
or U2753 (N_2753,N_2466,N_2580);
nand U2754 (N_2754,N_2552,N_2515);
nand U2755 (N_2755,N_2593,N_2476);
and U2756 (N_2756,N_2565,N_2501);
nor U2757 (N_2757,N_2461,N_2582);
nand U2758 (N_2758,N_2560,N_2578);
and U2759 (N_2759,N_2486,N_2576);
and U2760 (N_2760,N_2472,N_2471);
and U2761 (N_2761,N_2485,N_2572);
nor U2762 (N_2762,N_2509,N_2552);
and U2763 (N_2763,N_2439,N_2528);
and U2764 (N_2764,N_2450,N_2543);
or U2765 (N_2765,N_2446,N_2464);
and U2766 (N_2766,N_2425,N_2524);
nand U2767 (N_2767,N_2561,N_2488);
nand U2768 (N_2768,N_2470,N_2463);
and U2769 (N_2769,N_2407,N_2507);
nor U2770 (N_2770,N_2555,N_2494);
or U2771 (N_2771,N_2448,N_2452);
nor U2772 (N_2772,N_2420,N_2482);
or U2773 (N_2773,N_2560,N_2519);
or U2774 (N_2774,N_2401,N_2594);
nand U2775 (N_2775,N_2589,N_2488);
xor U2776 (N_2776,N_2469,N_2564);
or U2777 (N_2777,N_2485,N_2507);
xnor U2778 (N_2778,N_2595,N_2588);
or U2779 (N_2779,N_2503,N_2421);
nand U2780 (N_2780,N_2554,N_2455);
or U2781 (N_2781,N_2595,N_2567);
and U2782 (N_2782,N_2537,N_2546);
or U2783 (N_2783,N_2581,N_2594);
or U2784 (N_2784,N_2513,N_2531);
or U2785 (N_2785,N_2552,N_2571);
nand U2786 (N_2786,N_2479,N_2559);
nand U2787 (N_2787,N_2528,N_2591);
nand U2788 (N_2788,N_2428,N_2408);
or U2789 (N_2789,N_2528,N_2577);
nand U2790 (N_2790,N_2492,N_2533);
nor U2791 (N_2791,N_2593,N_2584);
and U2792 (N_2792,N_2483,N_2465);
and U2793 (N_2793,N_2426,N_2454);
or U2794 (N_2794,N_2575,N_2572);
and U2795 (N_2795,N_2481,N_2439);
nand U2796 (N_2796,N_2485,N_2528);
nor U2797 (N_2797,N_2505,N_2403);
nand U2798 (N_2798,N_2527,N_2544);
and U2799 (N_2799,N_2488,N_2453);
nand U2800 (N_2800,N_2798,N_2636);
nor U2801 (N_2801,N_2727,N_2643);
nor U2802 (N_2802,N_2781,N_2786);
nand U2803 (N_2803,N_2728,N_2637);
or U2804 (N_2804,N_2709,N_2664);
nand U2805 (N_2805,N_2777,N_2617);
nand U2806 (N_2806,N_2660,N_2742);
or U2807 (N_2807,N_2644,N_2656);
or U2808 (N_2808,N_2695,N_2683);
or U2809 (N_2809,N_2747,N_2611);
nor U2810 (N_2810,N_2640,N_2629);
or U2811 (N_2811,N_2659,N_2748);
or U2812 (N_2812,N_2774,N_2779);
nor U2813 (N_2813,N_2638,N_2794);
and U2814 (N_2814,N_2657,N_2651);
nor U2815 (N_2815,N_2761,N_2745);
nand U2816 (N_2816,N_2628,N_2738);
and U2817 (N_2817,N_2652,N_2620);
or U2818 (N_2818,N_2688,N_2627);
and U2819 (N_2819,N_2699,N_2749);
and U2820 (N_2820,N_2790,N_2678);
nor U2821 (N_2821,N_2765,N_2658);
nand U2822 (N_2822,N_2604,N_2713);
and U2823 (N_2823,N_2718,N_2703);
and U2824 (N_2824,N_2601,N_2714);
nand U2825 (N_2825,N_2619,N_2625);
or U2826 (N_2826,N_2600,N_2792);
nand U2827 (N_2827,N_2755,N_2720);
or U2828 (N_2828,N_2692,N_2743);
nor U2829 (N_2829,N_2759,N_2693);
nor U2830 (N_2830,N_2752,N_2634);
and U2831 (N_2831,N_2783,N_2618);
nor U2832 (N_2832,N_2641,N_2780);
nand U2833 (N_2833,N_2679,N_2613);
nand U2834 (N_2834,N_2632,N_2698);
and U2835 (N_2835,N_2711,N_2724);
nor U2836 (N_2836,N_2772,N_2754);
nand U2837 (N_2837,N_2622,N_2766);
nor U2838 (N_2838,N_2753,N_2681);
and U2839 (N_2839,N_2690,N_2722);
or U2840 (N_2840,N_2689,N_2776);
nor U2841 (N_2841,N_2633,N_2669);
nand U2842 (N_2842,N_2671,N_2707);
or U2843 (N_2843,N_2715,N_2680);
nor U2844 (N_2844,N_2677,N_2685);
and U2845 (N_2845,N_2675,N_2799);
and U2846 (N_2846,N_2701,N_2673);
nand U2847 (N_2847,N_2649,N_2672);
or U2848 (N_2848,N_2646,N_2788);
nor U2849 (N_2849,N_2764,N_2687);
or U2850 (N_2850,N_2726,N_2645);
nor U2851 (N_2851,N_2741,N_2609);
nand U2852 (N_2852,N_2712,N_2782);
nor U2853 (N_2853,N_2686,N_2697);
nor U2854 (N_2854,N_2735,N_2696);
or U2855 (N_2855,N_2740,N_2674);
and U2856 (N_2856,N_2631,N_2758);
and U2857 (N_2857,N_2736,N_2706);
nand U2858 (N_2858,N_2654,N_2616);
and U2859 (N_2859,N_2667,N_2682);
nor U2860 (N_2860,N_2731,N_2716);
or U2861 (N_2861,N_2784,N_2665);
and U2862 (N_2862,N_2642,N_2608);
or U2863 (N_2863,N_2639,N_2648);
or U2864 (N_2864,N_2615,N_2670);
or U2865 (N_2865,N_2773,N_2621);
or U2866 (N_2866,N_2663,N_2647);
or U2867 (N_2867,N_2791,N_2756);
nor U2868 (N_2868,N_2721,N_2610);
and U2869 (N_2869,N_2676,N_2750);
and U2870 (N_2870,N_2769,N_2694);
and U2871 (N_2871,N_2606,N_2723);
nor U2872 (N_2872,N_2796,N_2603);
and U2873 (N_2873,N_2797,N_2746);
nand U2874 (N_2874,N_2719,N_2612);
or U2875 (N_2875,N_2624,N_2705);
and U2876 (N_2876,N_2733,N_2734);
nand U2877 (N_2877,N_2684,N_2666);
or U2878 (N_2878,N_2655,N_2661);
or U2879 (N_2879,N_2668,N_2739);
nor U2880 (N_2880,N_2717,N_2737);
and U2881 (N_2881,N_2757,N_2789);
or U2882 (N_2882,N_2732,N_2662);
xor U2883 (N_2883,N_2793,N_2630);
nor U2884 (N_2884,N_2626,N_2710);
nor U2885 (N_2885,N_2607,N_2730);
and U2886 (N_2886,N_2760,N_2602);
or U2887 (N_2887,N_2729,N_2700);
or U2888 (N_2888,N_2770,N_2650);
nand U2889 (N_2889,N_2744,N_2635);
or U2890 (N_2890,N_2691,N_2763);
nand U2891 (N_2891,N_2785,N_2767);
or U2892 (N_2892,N_2768,N_2771);
or U2893 (N_2893,N_2614,N_2623);
nor U2894 (N_2894,N_2775,N_2653);
nand U2895 (N_2895,N_2751,N_2778);
or U2896 (N_2896,N_2702,N_2725);
or U2897 (N_2897,N_2708,N_2605);
or U2898 (N_2898,N_2787,N_2795);
nand U2899 (N_2899,N_2704,N_2762);
and U2900 (N_2900,N_2675,N_2790);
and U2901 (N_2901,N_2753,N_2603);
or U2902 (N_2902,N_2727,N_2662);
or U2903 (N_2903,N_2634,N_2670);
and U2904 (N_2904,N_2619,N_2784);
nor U2905 (N_2905,N_2649,N_2620);
nand U2906 (N_2906,N_2632,N_2790);
nor U2907 (N_2907,N_2665,N_2775);
or U2908 (N_2908,N_2758,N_2635);
nor U2909 (N_2909,N_2766,N_2695);
nand U2910 (N_2910,N_2612,N_2746);
nor U2911 (N_2911,N_2652,N_2729);
nor U2912 (N_2912,N_2771,N_2725);
and U2913 (N_2913,N_2653,N_2743);
and U2914 (N_2914,N_2619,N_2627);
nor U2915 (N_2915,N_2690,N_2739);
nor U2916 (N_2916,N_2734,N_2751);
or U2917 (N_2917,N_2621,N_2799);
and U2918 (N_2918,N_2620,N_2723);
or U2919 (N_2919,N_2661,N_2615);
nand U2920 (N_2920,N_2645,N_2600);
and U2921 (N_2921,N_2752,N_2604);
nor U2922 (N_2922,N_2665,N_2737);
xnor U2923 (N_2923,N_2739,N_2781);
nor U2924 (N_2924,N_2773,N_2686);
and U2925 (N_2925,N_2682,N_2658);
nand U2926 (N_2926,N_2727,N_2794);
nand U2927 (N_2927,N_2650,N_2709);
nand U2928 (N_2928,N_2711,N_2652);
nand U2929 (N_2929,N_2606,N_2797);
or U2930 (N_2930,N_2665,N_2653);
and U2931 (N_2931,N_2772,N_2792);
nand U2932 (N_2932,N_2622,N_2616);
nor U2933 (N_2933,N_2655,N_2664);
or U2934 (N_2934,N_2623,N_2694);
nor U2935 (N_2935,N_2639,N_2642);
or U2936 (N_2936,N_2696,N_2716);
nor U2937 (N_2937,N_2698,N_2744);
or U2938 (N_2938,N_2787,N_2734);
nand U2939 (N_2939,N_2650,N_2776);
and U2940 (N_2940,N_2677,N_2749);
nand U2941 (N_2941,N_2661,N_2761);
nor U2942 (N_2942,N_2727,N_2613);
nand U2943 (N_2943,N_2672,N_2755);
nor U2944 (N_2944,N_2607,N_2622);
or U2945 (N_2945,N_2762,N_2697);
xnor U2946 (N_2946,N_2716,N_2640);
and U2947 (N_2947,N_2760,N_2788);
or U2948 (N_2948,N_2728,N_2606);
and U2949 (N_2949,N_2647,N_2624);
nand U2950 (N_2950,N_2721,N_2656);
or U2951 (N_2951,N_2755,N_2618);
or U2952 (N_2952,N_2693,N_2645);
or U2953 (N_2953,N_2664,N_2741);
nand U2954 (N_2954,N_2620,N_2717);
and U2955 (N_2955,N_2647,N_2693);
nor U2956 (N_2956,N_2721,N_2623);
nand U2957 (N_2957,N_2763,N_2660);
or U2958 (N_2958,N_2663,N_2603);
and U2959 (N_2959,N_2688,N_2677);
and U2960 (N_2960,N_2658,N_2724);
and U2961 (N_2961,N_2779,N_2667);
xor U2962 (N_2962,N_2726,N_2669);
nor U2963 (N_2963,N_2791,N_2613);
nand U2964 (N_2964,N_2723,N_2641);
nand U2965 (N_2965,N_2645,N_2774);
and U2966 (N_2966,N_2722,N_2637);
or U2967 (N_2967,N_2622,N_2737);
or U2968 (N_2968,N_2706,N_2772);
or U2969 (N_2969,N_2719,N_2600);
or U2970 (N_2970,N_2771,N_2793);
nor U2971 (N_2971,N_2626,N_2618);
or U2972 (N_2972,N_2733,N_2739);
nand U2973 (N_2973,N_2763,N_2712);
nand U2974 (N_2974,N_2627,N_2625);
or U2975 (N_2975,N_2726,N_2637);
nand U2976 (N_2976,N_2676,N_2738);
nor U2977 (N_2977,N_2759,N_2611);
or U2978 (N_2978,N_2655,N_2634);
or U2979 (N_2979,N_2752,N_2779);
nor U2980 (N_2980,N_2697,N_2784);
or U2981 (N_2981,N_2730,N_2623);
nor U2982 (N_2982,N_2746,N_2752);
and U2983 (N_2983,N_2708,N_2721);
nor U2984 (N_2984,N_2703,N_2724);
nand U2985 (N_2985,N_2759,N_2772);
nand U2986 (N_2986,N_2749,N_2664);
nand U2987 (N_2987,N_2613,N_2781);
and U2988 (N_2988,N_2606,N_2706);
nor U2989 (N_2989,N_2634,N_2631);
nand U2990 (N_2990,N_2795,N_2737);
nor U2991 (N_2991,N_2784,N_2786);
and U2992 (N_2992,N_2663,N_2688);
nor U2993 (N_2993,N_2605,N_2728);
nor U2994 (N_2994,N_2616,N_2727);
or U2995 (N_2995,N_2746,N_2712);
nand U2996 (N_2996,N_2656,N_2660);
or U2997 (N_2997,N_2765,N_2629);
or U2998 (N_2998,N_2620,N_2763);
nor U2999 (N_2999,N_2614,N_2774);
and U3000 (N_3000,N_2897,N_2850);
nand U3001 (N_3001,N_2979,N_2879);
nand U3002 (N_3002,N_2944,N_2825);
nor U3003 (N_3003,N_2805,N_2876);
nand U3004 (N_3004,N_2994,N_2836);
and U3005 (N_3005,N_2887,N_2875);
nor U3006 (N_3006,N_2931,N_2856);
nor U3007 (N_3007,N_2802,N_2917);
and U3008 (N_3008,N_2828,N_2950);
nor U3009 (N_3009,N_2821,N_2945);
or U3010 (N_3010,N_2936,N_2848);
nor U3011 (N_3011,N_2860,N_2996);
nand U3012 (N_3012,N_2803,N_2977);
nand U3013 (N_3013,N_2822,N_2906);
nor U3014 (N_3014,N_2873,N_2854);
or U3015 (N_3015,N_2993,N_2868);
nor U3016 (N_3016,N_2989,N_2910);
and U3017 (N_3017,N_2867,N_2998);
or U3018 (N_3018,N_2874,N_2813);
nor U3019 (N_3019,N_2956,N_2893);
and U3020 (N_3020,N_2954,N_2997);
nand U3021 (N_3021,N_2863,N_2991);
nor U3022 (N_3022,N_2973,N_2878);
nor U3023 (N_3023,N_2970,N_2861);
and U3024 (N_3024,N_2833,N_2943);
and U3025 (N_3025,N_2890,N_2814);
and U3026 (N_3026,N_2962,N_2896);
nor U3027 (N_3027,N_2984,N_2978);
and U3028 (N_3028,N_2811,N_2930);
nor U3029 (N_3029,N_2992,N_2969);
nor U3030 (N_3030,N_2940,N_2899);
and U3031 (N_3031,N_2830,N_2918);
nand U3032 (N_3032,N_2841,N_2902);
nand U3033 (N_3033,N_2972,N_2832);
nand U3034 (N_3034,N_2818,N_2851);
and U3035 (N_3035,N_2842,N_2949);
nor U3036 (N_3036,N_2847,N_2871);
nand U3037 (N_3037,N_2809,N_2831);
and U3038 (N_3038,N_2933,N_2963);
nand U3039 (N_3039,N_2865,N_2932);
nand U3040 (N_3040,N_2838,N_2824);
nand U3041 (N_3041,N_2965,N_2892);
nor U3042 (N_3042,N_2988,N_2835);
or U3043 (N_3043,N_2881,N_2806);
nand U3044 (N_3044,N_2987,N_2929);
nand U3045 (N_3045,N_2857,N_2957);
nor U3046 (N_3046,N_2883,N_2900);
nor U3047 (N_3047,N_2928,N_2958);
or U3048 (N_3048,N_2974,N_2801);
or U3049 (N_3049,N_2921,N_2916);
or U3050 (N_3050,N_2815,N_2869);
or U3051 (N_3051,N_2826,N_2985);
nor U3052 (N_3052,N_2862,N_2823);
or U3053 (N_3053,N_2808,N_2853);
nand U3054 (N_3054,N_2880,N_2912);
or U3055 (N_3055,N_2990,N_2870);
nand U3056 (N_3056,N_2827,N_2971);
or U3057 (N_3057,N_2807,N_2904);
or U3058 (N_3058,N_2852,N_2829);
nor U3059 (N_3059,N_2849,N_2866);
nor U3060 (N_3060,N_2911,N_2925);
or U3061 (N_3061,N_2905,N_2903);
nand U3062 (N_3062,N_2981,N_2859);
nand U3063 (N_3063,N_2983,N_2946);
and U3064 (N_3064,N_2820,N_2999);
nor U3065 (N_3065,N_2924,N_2800);
or U3066 (N_3066,N_2920,N_2845);
nor U3067 (N_3067,N_2952,N_2941);
nor U3068 (N_3068,N_2942,N_2927);
nand U3069 (N_3069,N_2953,N_2947);
nor U3070 (N_3070,N_2982,N_2967);
and U3071 (N_3071,N_2948,N_2884);
nand U3072 (N_3072,N_2810,N_2938);
and U3073 (N_3073,N_2907,N_2895);
nand U3074 (N_3074,N_2864,N_2817);
nand U3075 (N_3075,N_2844,N_2889);
nand U3076 (N_3076,N_2964,N_2888);
nor U3077 (N_3077,N_2846,N_2812);
nor U3078 (N_3078,N_2885,N_2995);
nor U3079 (N_3079,N_2914,N_2901);
and U3080 (N_3080,N_2951,N_2840);
and U3081 (N_3081,N_2908,N_2959);
nand U3082 (N_3082,N_2960,N_2839);
and U3083 (N_3083,N_2976,N_2894);
nand U3084 (N_3084,N_2922,N_2955);
nor U3085 (N_3085,N_2923,N_2898);
or U3086 (N_3086,N_2926,N_2919);
or U3087 (N_3087,N_2939,N_2882);
nor U3088 (N_3088,N_2886,N_2843);
nor U3089 (N_3089,N_2891,N_2834);
or U3090 (N_3090,N_2837,N_2961);
nand U3091 (N_3091,N_2877,N_2966);
nand U3092 (N_3092,N_2872,N_2980);
nand U3093 (N_3093,N_2915,N_2819);
nand U3094 (N_3094,N_2935,N_2968);
or U3095 (N_3095,N_2937,N_2913);
or U3096 (N_3096,N_2858,N_2986);
or U3097 (N_3097,N_2816,N_2855);
nor U3098 (N_3098,N_2804,N_2909);
nand U3099 (N_3099,N_2975,N_2934);
or U3100 (N_3100,N_2809,N_2966);
nand U3101 (N_3101,N_2806,N_2915);
nand U3102 (N_3102,N_2939,N_2952);
or U3103 (N_3103,N_2841,N_2840);
and U3104 (N_3104,N_2920,N_2900);
nor U3105 (N_3105,N_2865,N_2828);
nor U3106 (N_3106,N_2900,N_2846);
nand U3107 (N_3107,N_2877,N_2993);
and U3108 (N_3108,N_2881,N_2962);
nor U3109 (N_3109,N_2970,N_2924);
nand U3110 (N_3110,N_2869,N_2879);
nand U3111 (N_3111,N_2966,N_2990);
nor U3112 (N_3112,N_2815,N_2966);
nor U3113 (N_3113,N_2877,N_2863);
nand U3114 (N_3114,N_2854,N_2966);
or U3115 (N_3115,N_2888,N_2913);
or U3116 (N_3116,N_2963,N_2979);
or U3117 (N_3117,N_2820,N_2977);
or U3118 (N_3118,N_2883,N_2939);
nand U3119 (N_3119,N_2897,N_2965);
and U3120 (N_3120,N_2828,N_2891);
and U3121 (N_3121,N_2942,N_2996);
or U3122 (N_3122,N_2859,N_2822);
nor U3123 (N_3123,N_2826,N_2996);
nor U3124 (N_3124,N_2846,N_2924);
and U3125 (N_3125,N_2823,N_2956);
and U3126 (N_3126,N_2824,N_2953);
nor U3127 (N_3127,N_2899,N_2894);
nand U3128 (N_3128,N_2905,N_2894);
nand U3129 (N_3129,N_2991,N_2955);
nand U3130 (N_3130,N_2981,N_2901);
or U3131 (N_3131,N_2915,N_2893);
nor U3132 (N_3132,N_2967,N_2920);
nand U3133 (N_3133,N_2964,N_2861);
xnor U3134 (N_3134,N_2836,N_2823);
and U3135 (N_3135,N_2973,N_2997);
or U3136 (N_3136,N_2816,N_2907);
or U3137 (N_3137,N_2954,N_2827);
and U3138 (N_3138,N_2923,N_2902);
nor U3139 (N_3139,N_2833,N_2920);
nand U3140 (N_3140,N_2898,N_2967);
or U3141 (N_3141,N_2836,N_2896);
or U3142 (N_3142,N_2848,N_2883);
and U3143 (N_3143,N_2850,N_2928);
and U3144 (N_3144,N_2884,N_2813);
nand U3145 (N_3145,N_2886,N_2941);
and U3146 (N_3146,N_2883,N_2895);
and U3147 (N_3147,N_2989,N_2985);
nand U3148 (N_3148,N_2804,N_2913);
and U3149 (N_3149,N_2804,N_2917);
or U3150 (N_3150,N_2911,N_2828);
nand U3151 (N_3151,N_2850,N_2835);
and U3152 (N_3152,N_2818,N_2916);
and U3153 (N_3153,N_2951,N_2969);
or U3154 (N_3154,N_2876,N_2900);
and U3155 (N_3155,N_2972,N_2831);
and U3156 (N_3156,N_2935,N_2834);
xor U3157 (N_3157,N_2956,N_2987);
and U3158 (N_3158,N_2829,N_2880);
and U3159 (N_3159,N_2876,N_2840);
nor U3160 (N_3160,N_2810,N_2866);
and U3161 (N_3161,N_2939,N_2819);
nor U3162 (N_3162,N_2963,N_2850);
or U3163 (N_3163,N_2916,N_2938);
xor U3164 (N_3164,N_2810,N_2826);
or U3165 (N_3165,N_2990,N_2911);
nor U3166 (N_3166,N_2912,N_2991);
nor U3167 (N_3167,N_2811,N_2815);
or U3168 (N_3168,N_2999,N_2876);
or U3169 (N_3169,N_2954,N_2961);
nand U3170 (N_3170,N_2807,N_2987);
nor U3171 (N_3171,N_2869,N_2893);
and U3172 (N_3172,N_2816,N_2859);
nand U3173 (N_3173,N_2994,N_2887);
nand U3174 (N_3174,N_2822,N_2875);
or U3175 (N_3175,N_2820,N_2996);
and U3176 (N_3176,N_2996,N_2998);
nand U3177 (N_3177,N_2900,N_2824);
nor U3178 (N_3178,N_2934,N_2937);
and U3179 (N_3179,N_2873,N_2942);
nand U3180 (N_3180,N_2947,N_2940);
or U3181 (N_3181,N_2995,N_2878);
or U3182 (N_3182,N_2856,N_2957);
or U3183 (N_3183,N_2986,N_2833);
nand U3184 (N_3184,N_2897,N_2839);
nand U3185 (N_3185,N_2881,N_2976);
nand U3186 (N_3186,N_2992,N_2998);
and U3187 (N_3187,N_2960,N_2967);
nand U3188 (N_3188,N_2948,N_2831);
and U3189 (N_3189,N_2860,N_2846);
nor U3190 (N_3190,N_2963,N_2939);
nor U3191 (N_3191,N_2812,N_2857);
and U3192 (N_3192,N_2929,N_2863);
nor U3193 (N_3193,N_2816,N_2891);
nand U3194 (N_3194,N_2815,N_2863);
nand U3195 (N_3195,N_2935,N_2966);
nand U3196 (N_3196,N_2868,N_2839);
nand U3197 (N_3197,N_2875,N_2878);
or U3198 (N_3198,N_2800,N_2833);
nor U3199 (N_3199,N_2976,N_2981);
nand U3200 (N_3200,N_3152,N_3175);
or U3201 (N_3201,N_3052,N_3173);
and U3202 (N_3202,N_3078,N_3132);
or U3203 (N_3203,N_3119,N_3155);
nand U3204 (N_3204,N_3099,N_3053);
and U3205 (N_3205,N_3063,N_3080);
nand U3206 (N_3206,N_3019,N_3151);
nor U3207 (N_3207,N_3006,N_3084);
nor U3208 (N_3208,N_3020,N_3074);
nor U3209 (N_3209,N_3178,N_3017);
and U3210 (N_3210,N_3001,N_3032);
and U3211 (N_3211,N_3035,N_3086);
and U3212 (N_3212,N_3114,N_3136);
or U3213 (N_3213,N_3058,N_3158);
nor U3214 (N_3214,N_3166,N_3168);
and U3215 (N_3215,N_3143,N_3077);
and U3216 (N_3216,N_3033,N_3054);
nor U3217 (N_3217,N_3096,N_3009);
or U3218 (N_3218,N_3180,N_3056);
nor U3219 (N_3219,N_3062,N_3179);
xor U3220 (N_3220,N_3100,N_3103);
or U3221 (N_3221,N_3163,N_3002);
or U3222 (N_3222,N_3190,N_3102);
nand U3223 (N_3223,N_3192,N_3048);
nand U3224 (N_3224,N_3036,N_3115);
nand U3225 (N_3225,N_3150,N_3174);
nand U3226 (N_3226,N_3011,N_3161);
and U3227 (N_3227,N_3188,N_3037);
nand U3228 (N_3228,N_3061,N_3075);
or U3229 (N_3229,N_3170,N_3144);
nand U3230 (N_3230,N_3027,N_3087);
nor U3231 (N_3231,N_3128,N_3124);
or U3232 (N_3232,N_3177,N_3184);
and U3233 (N_3233,N_3113,N_3133);
and U3234 (N_3234,N_3145,N_3157);
nor U3235 (N_3235,N_3051,N_3094);
and U3236 (N_3236,N_3055,N_3183);
or U3237 (N_3237,N_3066,N_3187);
or U3238 (N_3238,N_3014,N_3024);
and U3239 (N_3239,N_3159,N_3122);
xnor U3240 (N_3240,N_3003,N_3149);
and U3241 (N_3241,N_3081,N_3076);
nand U3242 (N_3242,N_3041,N_3073);
and U3243 (N_3243,N_3182,N_3046);
or U3244 (N_3244,N_3164,N_3044);
and U3245 (N_3245,N_3069,N_3111);
or U3246 (N_3246,N_3194,N_3082);
or U3247 (N_3247,N_3071,N_3015);
or U3248 (N_3248,N_3116,N_3092);
or U3249 (N_3249,N_3167,N_3064);
and U3250 (N_3250,N_3049,N_3018);
nand U3251 (N_3251,N_3043,N_3107);
nand U3252 (N_3252,N_3176,N_3068);
nand U3253 (N_3253,N_3146,N_3195);
and U3254 (N_3254,N_3067,N_3045);
nand U3255 (N_3255,N_3105,N_3160);
or U3256 (N_3256,N_3186,N_3034);
nor U3257 (N_3257,N_3140,N_3199);
and U3258 (N_3258,N_3172,N_3093);
nor U3259 (N_3259,N_3108,N_3121);
nor U3260 (N_3260,N_3169,N_3125);
nand U3261 (N_3261,N_3142,N_3141);
and U3262 (N_3262,N_3090,N_3057);
nand U3263 (N_3263,N_3112,N_3127);
or U3264 (N_3264,N_3029,N_3156);
or U3265 (N_3265,N_3123,N_3109);
or U3266 (N_3266,N_3031,N_3040);
nand U3267 (N_3267,N_3138,N_3021);
and U3268 (N_3268,N_3007,N_3005);
and U3269 (N_3269,N_3097,N_3131);
and U3270 (N_3270,N_3028,N_3013);
nand U3271 (N_3271,N_3026,N_3091);
nor U3272 (N_3272,N_3197,N_3104);
and U3273 (N_3273,N_3171,N_3198);
nor U3274 (N_3274,N_3196,N_3000);
and U3275 (N_3275,N_3079,N_3126);
and U3276 (N_3276,N_3130,N_3010);
nor U3277 (N_3277,N_3085,N_3110);
nor U3278 (N_3278,N_3022,N_3193);
nand U3279 (N_3279,N_3148,N_3038);
nor U3280 (N_3280,N_3118,N_3050);
and U3281 (N_3281,N_3004,N_3016);
and U3282 (N_3282,N_3098,N_3162);
and U3283 (N_3283,N_3030,N_3135);
and U3284 (N_3284,N_3147,N_3072);
nor U3285 (N_3285,N_3137,N_3070);
nand U3286 (N_3286,N_3088,N_3025);
nand U3287 (N_3287,N_3117,N_3089);
and U3288 (N_3288,N_3154,N_3060);
and U3289 (N_3289,N_3181,N_3106);
or U3290 (N_3290,N_3095,N_3023);
or U3291 (N_3291,N_3191,N_3065);
or U3292 (N_3292,N_3012,N_3059);
and U3293 (N_3293,N_3042,N_3039);
and U3294 (N_3294,N_3129,N_3120);
or U3295 (N_3295,N_3185,N_3083);
nor U3296 (N_3296,N_3139,N_3134);
nand U3297 (N_3297,N_3047,N_3101);
nor U3298 (N_3298,N_3165,N_3189);
nand U3299 (N_3299,N_3153,N_3008);
or U3300 (N_3300,N_3165,N_3101);
and U3301 (N_3301,N_3113,N_3140);
nand U3302 (N_3302,N_3152,N_3046);
and U3303 (N_3303,N_3062,N_3078);
nand U3304 (N_3304,N_3007,N_3018);
and U3305 (N_3305,N_3178,N_3031);
and U3306 (N_3306,N_3019,N_3073);
nand U3307 (N_3307,N_3083,N_3110);
nand U3308 (N_3308,N_3077,N_3166);
or U3309 (N_3309,N_3158,N_3089);
nand U3310 (N_3310,N_3115,N_3096);
or U3311 (N_3311,N_3012,N_3192);
nand U3312 (N_3312,N_3088,N_3064);
and U3313 (N_3313,N_3179,N_3064);
nand U3314 (N_3314,N_3156,N_3137);
and U3315 (N_3315,N_3032,N_3016);
nand U3316 (N_3316,N_3120,N_3090);
nor U3317 (N_3317,N_3022,N_3031);
nand U3318 (N_3318,N_3122,N_3028);
xnor U3319 (N_3319,N_3158,N_3051);
nand U3320 (N_3320,N_3076,N_3054);
and U3321 (N_3321,N_3143,N_3186);
nand U3322 (N_3322,N_3126,N_3092);
nand U3323 (N_3323,N_3009,N_3153);
and U3324 (N_3324,N_3129,N_3117);
nand U3325 (N_3325,N_3012,N_3170);
or U3326 (N_3326,N_3085,N_3034);
or U3327 (N_3327,N_3084,N_3041);
nor U3328 (N_3328,N_3161,N_3172);
nand U3329 (N_3329,N_3165,N_3033);
and U3330 (N_3330,N_3120,N_3008);
nand U3331 (N_3331,N_3103,N_3067);
nor U3332 (N_3332,N_3026,N_3083);
nand U3333 (N_3333,N_3157,N_3096);
nor U3334 (N_3334,N_3017,N_3053);
nand U3335 (N_3335,N_3189,N_3168);
and U3336 (N_3336,N_3089,N_3136);
and U3337 (N_3337,N_3069,N_3014);
nand U3338 (N_3338,N_3153,N_3137);
nand U3339 (N_3339,N_3184,N_3166);
nor U3340 (N_3340,N_3186,N_3100);
and U3341 (N_3341,N_3062,N_3136);
and U3342 (N_3342,N_3102,N_3135);
nor U3343 (N_3343,N_3174,N_3152);
and U3344 (N_3344,N_3152,N_3114);
or U3345 (N_3345,N_3043,N_3102);
nand U3346 (N_3346,N_3114,N_3194);
xor U3347 (N_3347,N_3016,N_3036);
and U3348 (N_3348,N_3043,N_3049);
nand U3349 (N_3349,N_3180,N_3054);
or U3350 (N_3350,N_3021,N_3198);
and U3351 (N_3351,N_3131,N_3089);
nor U3352 (N_3352,N_3182,N_3192);
and U3353 (N_3353,N_3197,N_3037);
and U3354 (N_3354,N_3040,N_3174);
nand U3355 (N_3355,N_3145,N_3051);
and U3356 (N_3356,N_3152,N_3016);
or U3357 (N_3357,N_3131,N_3123);
or U3358 (N_3358,N_3029,N_3088);
and U3359 (N_3359,N_3071,N_3116);
nand U3360 (N_3360,N_3103,N_3069);
nor U3361 (N_3361,N_3074,N_3057);
nand U3362 (N_3362,N_3081,N_3018);
and U3363 (N_3363,N_3132,N_3043);
nand U3364 (N_3364,N_3070,N_3133);
or U3365 (N_3365,N_3038,N_3083);
or U3366 (N_3366,N_3100,N_3121);
nand U3367 (N_3367,N_3022,N_3099);
nor U3368 (N_3368,N_3019,N_3164);
or U3369 (N_3369,N_3134,N_3037);
nor U3370 (N_3370,N_3070,N_3140);
nor U3371 (N_3371,N_3078,N_3074);
and U3372 (N_3372,N_3145,N_3185);
or U3373 (N_3373,N_3182,N_3078);
and U3374 (N_3374,N_3075,N_3097);
and U3375 (N_3375,N_3013,N_3085);
and U3376 (N_3376,N_3004,N_3072);
or U3377 (N_3377,N_3187,N_3079);
and U3378 (N_3378,N_3131,N_3088);
and U3379 (N_3379,N_3015,N_3049);
xnor U3380 (N_3380,N_3000,N_3095);
and U3381 (N_3381,N_3007,N_3136);
and U3382 (N_3382,N_3133,N_3068);
and U3383 (N_3383,N_3138,N_3075);
nor U3384 (N_3384,N_3188,N_3101);
nor U3385 (N_3385,N_3007,N_3092);
nor U3386 (N_3386,N_3019,N_3118);
or U3387 (N_3387,N_3028,N_3082);
or U3388 (N_3388,N_3150,N_3099);
nor U3389 (N_3389,N_3157,N_3009);
nand U3390 (N_3390,N_3174,N_3024);
nor U3391 (N_3391,N_3124,N_3150);
and U3392 (N_3392,N_3097,N_3135);
nor U3393 (N_3393,N_3016,N_3013);
nand U3394 (N_3394,N_3063,N_3138);
and U3395 (N_3395,N_3180,N_3006);
and U3396 (N_3396,N_3063,N_3013);
or U3397 (N_3397,N_3011,N_3115);
nor U3398 (N_3398,N_3199,N_3057);
and U3399 (N_3399,N_3040,N_3036);
nor U3400 (N_3400,N_3249,N_3224);
nand U3401 (N_3401,N_3309,N_3225);
nand U3402 (N_3402,N_3219,N_3335);
nand U3403 (N_3403,N_3380,N_3367);
nand U3404 (N_3404,N_3291,N_3236);
or U3405 (N_3405,N_3237,N_3305);
nand U3406 (N_3406,N_3233,N_3362);
nand U3407 (N_3407,N_3358,N_3332);
and U3408 (N_3408,N_3329,N_3286);
nand U3409 (N_3409,N_3384,N_3349);
nand U3410 (N_3410,N_3378,N_3360);
nand U3411 (N_3411,N_3299,N_3379);
or U3412 (N_3412,N_3206,N_3375);
or U3413 (N_3413,N_3242,N_3326);
or U3414 (N_3414,N_3231,N_3355);
nor U3415 (N_3415,N_3210,N_3234);
or U3416 (N_3416,N_3325,N_3247);
and U3417 (N_3417,N_3287,N_3339);
or U3418 (N_3418,N_3398,N_3382);
and U3419 (N_3419,N_3356,N_3273);
and U3420 (N_3420,N_3353,N_3227);
nand U3421 (N_3421,N_3293,N_3301);
and U3422 (N_3422,N_3303,N_3274);
nor U3423 (N_3423,N_3359,N_3290);
nand U3424 (N_3424,N_3207,N_3283);
nor U3425 (N_3425,N_3387,N_3289);
and U3426 (N_3426,N_3240,N_3363);
and U3427 (N_3427,N_3328,N_3279);
nor U3428 (N_3428,N_3221,N_3282);
nor U3429 (N_3429,N_3269,N_3220);
nand U3430 (N_3430,N_3372,N_3288);
or U3431 (N_3431,N_3370,N_3205);
nor U3432 (N_3432,N_3228,N_3369);
nand U3433 (N_3433,N_3331,N_3250);
and U3434 (N_3434,N_3376,N_3350);
and U3435 (N_3435,N_3397,N_3256);
nor U3436 (N_3436,N_3336,N_3213);
and U3437 (N_3437,N_3211,N_3351);
nor U3438 (N_3438,N_3347,N_3212);
nand U3439 (N_3439,N_3229,N_3364);
xor U3440 (N_3440,N_3238,N_3343);
or U3441 (N_3441,N_3203,N_3396);
and U3442 (N_3442,N_3338,N_3346);
and U3443 (N_3443,N_3204,N_3352);
nor U3444 (N_3444,N_3313,N_3395);
nand U3445 (N_3445,N_3318,N_3366);
nor U3446 (N_3446,N_3312,N_3292);
nor U3447 (N_3447,N_3334,N_3389);
or U3448 (N_3448,N_3278,N_3266);
nor U3449 (N_3449,N_3337,N_3295);
nor U3450 (N_3450,N_3252,N_3248);
nor U3451 (N_3451,N_3268,N_3342);
or U3452 (N_3452,N_3230,N_3253);
and U3453 (N_3453,N_3263,N_3232);
and U3454 (N_3454,N_3304,N_3264);
or U3455 (N_3455,N_3386,N_3285);
nand U3456 (N_3456,N_3244,N_3259);
nand U3457 (N_3457,N_3281,N_3323);
or U3458 (N_3458,N_3317,N_3381);
nand U3459 (N_3459,N_3391,N_3255);
nand U3460 (N_3460,N_3223,N_3275);
nor U3461 (N_3461,N_3315,N_3383);
or U3462 (N_3462,N_3316,N_3393);
and U3463 (N_3463,N_3209,N_3201);
nor U3464 (N_3464,N_3214,N_3307);
nand U3465 (N_3465,N_3399,N_3365);
and U3466 (N_3466,N_3348,N_3235);
or U3467 (N_3467,N_3361,N_3302);
or U3468 (N_3468,N_3344,N_3377);
nand U3469 (N_3469,N_3330,N_3319);
and U3470 (N_3470,N_3371,N_3340);
and U3471 (N_3471,N_3310,N_3320);
nor U3472 (N_3472,N_3333,N_3239);
nand U3473 (N_3473,N_3322,N_3202);
or U3474 (N_3474,N_3300,N_3388);
and U3475 (N_3475,N_3200,N_3222);
nor U3476 (N_3476,N_3321,N_3265);
nand U3477 (N_3477,N_3298,N_3280);
or U3478 (N_3478,N_3284,N_3374);
nand U3479 (N_3479,N_3385,N_3373);
xor U3480 (N_3480,N_3216,N_3261);
or U3481 (N_3481,N_3271,N_3226);
nor U3482 (N_3482,N_3394,N_3270);
and U3483 (N_3483,N_3260,N_3392);
and U3484 (N_3484,N_3245,N_3311);
nor U3485 (N_3485,N_3296,N_3251);
nand U3486 (N_3486,N_3243,N_3314);
or U3487 (N_3487,N_3345,N_3354);
and U3488 (N_3488,N_3258,N_3277);
and U3489 (N_3489,N_3241,N_3368);
nand U3490 (N_3490,N_3217,N_3297);
and U3491 (N_3491,N_3357,N_3306);
and U3492 (N_3492,N_3276,N_3208);
nand U3493 (N_3493,N_3267,N_3246);
nand U3494 (N_3494,N_3254,N_3257);
nand U3495 (N_3495,N_3215,N_3390);
nand U3496 (N_3496,N_3272,N_3218);
or U3497 (N_3497,N_3294,N_3327);
nor U3498 (N_3498,N_3308,N_3262);
and U3499 (N_3499,N_3324,N_3341);
nor U3500 (N_3500,N_3343,N_3313);
or U3501 (N_3501,N_3359,N_3322);
nor U3502 (N_3502,N_3220,N_3251);
and U3503 (N_3503,N_3293,N_3322);
nand U3504 (N_3504,N_3239,N_3201);
or U3505 (N_3505,N_3232,N_3223);
and U3506 (N_3506,N_3305,N_3216);
or U3507 (N_3507,N_3282,N_3379);
and U3508 (N_3508,N_3293,N_3228);
nand U3509 (N_3509,N_3290,N_3319);
nand U3510 (N_3510,N_3209,N_3381);
and U3511 (N_3511,N_3374,N_3278);
nand U3512 (N_3512,N_3290,N_3243);
nand U3513 (N_3513,N_3397,N_3368);
or U3514 (N_3514,N_3236,N_3368);
nor U3515 (N_3515,N_3360,N_3214);
nand U3516 (N_3516,N_3385,N_3216);
nand U3517 (N_3517,N_3319,N_3298);
nand U3518 (N_3518,N_3228,N_3259);
or U3519 (N_3519,N_3270,N_3298);
nand U3520 (N_3520,N_3371,N_3234);
nor U3521 (N_3521,N_3335,N_3391);
nor U3522 (N_3522,N_3368,N_3240);
and U3523 (N_3523,N_3222,N_3271);
and U3524 (N_3524,N_3214,N_3242);
nand U3525 (N_3525,N_3203,N_3370);
nor U3526 (N_3526,N_3321,N_3327);
nor U3527 (N_3527,N_3397,N_3247);
and U3528 (N_3528,N_3261,N_3376);
nand U3529 (N_3529,N_3338,N_3314);
or U3530 (N_3530,N_3202,N_3306);
and U3531 (N_3531,N_3267,N_3392);
and U3532 (N_3532,N_3258,N_3244);
and U3533 (N_3533,N_3270,N_3205);
and U3534 (N_3534,N_3351,N_3285);
xor U3535 (N_3535,N_3300,N_3319);
nor U3536 (N_3536,N_3227,N_3380);
or U3537 (N_3537,N_3276,N_3377);
nand U3538 (N_3538,N_3378,N_3331);
nand U3539 (N_3539,N_3365,N_3273);
and U3540 (N_3540,N_3349,N_3250);
nor U3541 (N_3541,N_3220,N_3333);
or U3542 (N_3542,N_3225,N_3288);
or U3543 (N_3543,N_3399,N_3369);
and U3544 (N_3544,N_3301,N_3252);
nor U3545 (N_3545,N_3260,N_3243);
and U3546 (N_3546,N_3320,N_3319);
nand U3547 (N_3547,N_3377,N_3240);
nor U3548 (N_3548,N_3284,N_3390);
and U3549 (N_3549,N_3269,N_3324);
nand U3550 (N_3550,N_3231,N_3259);
xor U3551 (N_3551,N_3311,N_3361);
or U3552 (N_3552,N_3235,N_3224);
nand U3553 (N_3553,N_3395,N_3311);
or U3554 (N_3554,N_3294,N_3355);
nor U3555 (N_3555,N_3282,N_3366);
and U3556 (N_3556,N_3381,N_3241);
nor U3557 (N_3557,N_3216,N_3325);
nand U3558 (N_3558,N_3237,N_3211);
and U3559 (N_3559,N_3270,N_3214);
nand U3560 (N_3560,N_3313,N_3242);
or U3561 (N_3561,N_3266,N_3324);
nand U3562 (N_3562,N_3380,N_3332);
and U3563 (N_3563,N_3354,N_3303);
or U3564 (N_3564,N_3238,N_3326);
and U3565 (N_3565,N_3299,N_3262);
nor U3566 (N_3566,N_3307,N_3237);
and U3567 (N_3567,N_3389,N_3210);
and U3568 (N_3568,N_3267,N_3257);
nand U3569 (N_3569,N_3354,N_3323);
or U3570 (N_3570,N_3284,N_3244);
nor U3571 (N_3571,N_3322,N_3364);
or U3572 (N_3572,N_3379,N_3286);
and U3573 (N_3573,N_3270,N_3311);
nor U3574 (N_3574,N_3353,N_3254);
or U3575 (N_3575,N_3203,N_3392);
nor U3576 (N_3576,N_3261,N_3365);
nand U3577 (N_3577,N_3203,N_3306);
nand U3578 (N_3578,N_3260,N_3267);
nor U3579 (N_3579,N_3311,N_3370);
or U3580 (N_3580,N_3397,N_3227);
or U3581 (N_3581,N_3257,N_3282);
or U3582 (N_3582,N_3358,N_3330);
nand U3583 (N_3583,N_3205,N_3312);
and U3584 (N_3584,N_3208,N_3247);
or U3585 (N_3585,N_3358,N_3215);
nand U3586 (N_3586,N_3296,N_3244);
or U3587 (N_3587,N_3286,N_3320);
nand U3588 (N_3588,N_3225,N_3298);
nand U3589 (N_3589,N_3242,N_3383);
or U3590 (N_3590,N_3254,N_3207);
and U3591 (N_3591,N_3203,N_3384);
nor U3592 (N_3592,N_3211,N_3229);
nand U3593 (N_3593,N_3221,N_3350);
nor U3594 (N_3594,N_3278,N_3384);
nand U3595 (N_3595,N_3276,N_3319);
nand U3596 (N_3596,N_3369,N_3307);
nor U3597 (N_3597,N_3345,N_3286);
and U3598 (N_3598,N_3380,N_3271);
nor U3599 (N_3599,N_3208,N_3342);
nand U3600 (N_3600,N_3522,N_3456);
nor U3601 (N_3601,N_3521,N_3585);
or U3602 (N_3602,N_3534,N_3535);
or U3603 (N_3603,N_3455,N_3536);
or U3604 (N_3604,N_3510,N_3516);
or U3605 (N_3605,N_3409,N_3464);
and U3606 (N_3606,N_3441,N_3462);
and U3607 (N_3607,N_3403,N_3400);
and U3608 (N_3608,N_3527,N_3555);
nand U3609 (N_3609,N_3405,N_3471);
nand U3610 (N_3610,N_3570,N_3429);
or U3611 (N_3611,N_3439,N_3571);
or U3612 (N_3612,N_3416,N_3572);
nor U3613 (N_3613,N_3406,N_3562);
and U3614 (N_3614,N_3577,N_3497);
and U3615 (N_3615,N_3436,N_3424);
or U3616 (N_3616,N_3586,N_3569);
nor U3617 (N_3617,N_3457,N_3538);
and U3618 (N_3618,N_3465,N_3531);
and U3619 (N_3619,N_3501,N_3448);
nand U3620 (N_3620,N_3559,N_3575);
nor U3621 (N_3621,N_3410,N_3589);
or U3622 (N_3622,N_3469,N_3496);
or U3623 (N_3623,N_3453,N_3446);
and U3624 (N_3624,N_3461,N_3508);
and U3625 (N_3625,N_3599,N_3594);
nor U3626 (N_3626,N_3408,N_3458);
and U3627 (N_3627,N_3505,N_3493);
nand U3628 (N_3628,N_3475,N_3427);
or U3629 (N_3629,N_3428,N_3590);
nand U3630 (N_3630,N_3499,N_3454);
or U3631 (N_3631,N_3419,N_3504);
nand U3632 (N_3632,N_3494,N_3533);
nor U3633 (N_3633,N_3554,N_3430);
or U3634 (N_3634,N_3511,N_3546);
nand U3635 (N_3635,N_3483,N_3420);
nor U3636 (N_3636,N_3418,N_3451);
and U3637 (N_3637,N_3593,N_3574);
and U3638 (N_3638,N_3438,N_3490);
and U3639 (N_3639,N_3423,N_3415);
xor U3640 (N_3640,N_3547,N_3582);
and U3641 (N_3641,N_3411,N_3549);
and U3642 (N_3642,N_3530,N_3445);
and U3643 (N_3643,N_3517,N_3459);
nand U3644 (N_3644,N_3491,N_3584);
or U3645 (N_3645,N_3532,N_3467);
xnor U3646 (N_3646,N_3502,N_3515);
nor U3647 (N_3647,N_3477,N_3579);
or U3648 (N_3648,N_3402,N_3413);
and U3649 (N_3649,N_3443,N_3523);
or U3650 (N_3650,N_3537,N_3544);
nor U3651 (N_3651,N_3592,N_3404);
nor U3652 (N_3652,N_3492,N_3513);
and U3653 (N_3653,N_3525,N_3503);
or U3654 (N_3654,N_3449,N_3528);
or U3655 (N_3655,N_3548,N_3550);
and U3656 (N_3656,N_3563,N_3595);
nand U3657 (N_3657,N_3426,N_3509);
nor U3658 (N_3658,N_3553,N_3540);
nand U3659 (N_3659,N_3431,N_3434);
and U3660 (N_3660,N_3485,N_3519);
and U3661 (N_3661,N_3468,N_3591);
nor U3662 (N_3662,N_3564,N_3543);
nor U3663 (N_3663,N_3588,N_3460);
or U3664 (N_3664,N_3597,N_3520);
nand U3665 (N_3665,N_3583,N_3541);
and U3666 (N_3666,N_3421,N_3567);
and U3667 (N_3667,N_3425,N_3542);
and U3668 (N_3668,N_3442,N_3482);
or U3669 (N_3669,N_3512,N_3440);
nor U3670 (N_3670,N_3598,N_3578);
and U3671 (N_3671,N_3487,N_3506);
or U3672 (N_3672,N_3407,N_3529);
and U3673 (N_3673,N_3488,N_3433);
or U3674 (N_3674,N_3526,N_3566);
or U3675 (N_3675,N_3507,N_3484);
and U3676 (N_3676,N_3481,N_3524);
nand U3677 (N_3677,N_3514,N_3556);
nor U3678 (N_3678,N_3444,N_3561);
or U3679 (N_3679,N_3552,N_3466);
and U3680 (N_3680,N_3573,N_3476);
nor U3681 (N_3681,N_3498,N_3500);
nor U3682 (N_3682,N_3470,N_3412);
nand U3683 (N_3683,N_3435,N_3414);
nor U3684 (N_3684,N_3565,N_3474);
nor U3685 (N_3685,N_3568,N_3545);
and U3686 (N_3686,N_3518,N_3452);
nor U3687 (N_3687,N_3450,N_3486);
nor U3688 (N_3688,N_3447,N_3539);
and U3689 (N_3689,N_3463,N_3480);
nand U3690 (N_3690,N_3587,N_3473);
or U3691 (N_3691,N_3489,N_3479);
or U3692 (N_3692,N_3557,N_3472);
and U3693 (N_3693,N_3581,N_3495);
and U3694 (N_3694,N_3596,N_3576);
and U3695 (N_3695,N_3551,N_3478);
and U3696 (N_3696,N_3580,N_3417);
nor U3697 (N_3697,N_3437,N_3432);
nor U3698 (N_3698,N_3422,N_3558);
or U3699 (N_3699,N_3401,N_3560);
nand U3700 (N_3700,N_3494,N_3522);
nand U3701 (N_3701,N_3425,N_3497);
and U3702 (N_3702,N_3414,N_3492);
nor U3703 (N_3703,N_3538,N_3417);
nor U3704 (N_3704,N_3402,N_3543);
nand U3705 (N_3705,N_3593,N_3459);
nand U3706 (N_3706,N_3512,N_3498);
nor U3707 (N_3707,N_3573,N_3452);
or U3708 (N_3708,N_3515,N_3440);
nor U3709 (N_3709,N_3414,N_3514);
and U3710 (N_3710,N_3466,N_3577);
or U3711 (N_3711,N_3515,N_3471);
nor U3712 (N_3712,N_3540,N_3515);
and U3713 (N_3713,N_3543,N_3510);
nand U3714 (N_3714,N_3462,N_3549);
and U3715 (N_3715,N_3405,N_3579);
or U3716 (N_3716,N_3558,N_3480);
nor U3717 (N_3717,N_3455,N_3559);
nor U3718 (N_3718,N_3514,N_3562);
nor U3719 (N_3719,N_3489,N_3552);
or U3720 (N_3720,N_3519,N_3575);
or U3721 (N_3721,N_3498,N_3533);
nand U3722 (N_3722,N_3492,N_3496);
nand U3723 (N_3723,N_3595,N_3461);
or U3724 (N_3724,N_3472,N_3539);
nand U3725 (N_3725,N_3497,N_3520);
nor U3726 (N_3726,N_3473,N_3430);
nor U3727 (N_3727,N_3522,N_3569);
and U3728 (N_3728,N_3464,N_3558);
nand U3729 (N_3729,N_3454,N_3445);
or U3730 (N_3730,N_3420,N_3423);
nand U3731 (N_3731,N_3497,N_3557);
nand U3732 (N_3732,N_3553,N_3491);
or U3733 (N_3733,N_3525,N_3596);
or U3734 (N_3734,N_3414,N_3486);
and U3735 (N_3735,N_3475,N_3488);
nand U3736 (N_3736,N_3474,N_3422);
nand U3737 (N_3737,N_3532,N_3408);
and U3738 (N_3738,N_3504,N_3486);
nor U3739 (N_3739,N_3549,N_3455);
nand U3740 (N_3740,N_3579,N_3465);
nand U3741 (N_3741,N_3450,N_3518);
or U3742 (N_3742,N_3535,N_3547);
nand U3743 (N_3743,N_3434,N_3596);
nand U3744 (N_3744,N_3596,N_3598);
nor U3745 (N_3745,N_3579,N_3568);
nor U3746 (N_3746,N_3576,N_3483);
xnor U3747 (N_3747,N_3530,N_3481);
and U3748 (N_3748,N_3512,N_3479);
or U3749 (N_3749,N_3592,N_3437);
nor U3750 (N_3750,N_3428,N_3493);
or U3751 (N_3751,N_3482,N_3422);
or U3752 (N_3752,N_3523,N_3562);
or U3753 (N_3753,N_3500,N_3573);
and U3754 (N_3754,N_3582,N_3565);
nand U3755 (N_3755,N_3484,N_3488);
nor U3756 (N_3756,N_3492,N_3533);
nand U3757 (N_3757,N_3548,N_3422);
or U3758 (N_3758,N_3490,N_3444);
nand U3759 (N_3759,N_3495,N_3491);
and U3760 (N_3760,N_3489,N_3437);
and U3761 (N_3761,N_3483,N_3538);
or U3762 (N_3762,N_3553,N_3450);
nand U3763 (N_3763,N_3506,N_3583);
or U3764 (N_3764,N_3582,N_3509);
nand U3765 (N_3765,N_3550,N_3415);
or U3766 (N_3766,N_3543,N_3438);
nand U3767 (N_3767,N_3439,N_3487);
nand U3768 (N_3768,N_3426,N_3433);
nor U3769 (N_3769,N_3469,N_3501);
nor U3770 (N_3770,N_3455,N_3576);
nor U3771 (N_3771,N_3534,N_3420);
and U3772 (N_3772,N_3479,N_3551);
or U3773 (N_3773,N_3410,N_3592);
nor U3774 (N_3774,N_3428,N_3423);
nand U3775 (N_3775,N_3407,N_3462);
nor U3776 (N_3776,N_3436,N_3429);
or U3777 (N_3777,N_3489,N_3522);
and U3778 (N_3778,N_3401,N_3511);
nor U3779 (N_3779,N_3514,N_3597);
or U3780 (N_3780,N_3432,N_3538);
nand U3781 (N_3781,N_3585,N_3468);
and U3782 (N_3782,N_3478,N_3503);
nand U3783 (N_3783,N_3412,N_3587);
and U3784 (N_3784,N_3405,N_3595);
nor U3785 (N_3785,N_3540,N_3528);
xor U3786 (N_3786,N_3404,N_3490);
nor U3787 (N_3787,N_3588,N_3538);
or U3788 (N_3788,N_3485,N_3521);
nand U3789 (N_3789,N_3446,N_3517);
and U3790 (N_3790,N_3519,N_3596);
and U3791 (N_3791,N_3466,N_3487);
nor U3792 (N_3792,N_3431,N_3507);
and U3793 (N_3793,N_3442,N_3573);
and U3794 (N_3794,N_3484,N_3574);
and U3795 (N_3795,N_3492,N_3523);
nor U3796 (N_3796,N_3433,N_3410);
xnor U3797 (N_3797,N_3404,N_3548);
or U3798 (N_3798,N_3528,N_3573);
and U3799 (N_3799,N_3459,N_3492);
nand U3800 (N_3800,N_3626,N_3779);
nand U3801 (N_3801,N_3646,N_3785);
nand U3802 (N_3802,N_3717,N_3694);
or U3803 (N_3803,N_3676,N_3647);
nand U3804 (N_3804,N_3727,N_3730);
and U3805 (N_3805,N_3629,N_3794);
nor U3806 (N_3806,N_3619,N_3639);
nor U3807 (N_3807,N_3738,N_3614);
and U3808 (N_3808,N_3799,N_3702);
or U3809 (N_3809,N_3624,N_3737);
and U3810 (N_3810,N_3697,N_3611);
and U3811 (N_3811,N_3643,N_3612);
nand U3812 (N_3812,N_3608,N_3719);
or U3813 (N_3813,N_3743,N_3712);
and U3814 (N_3814,N_3628,N_3782);
and U3815 (N_3815,N_3795,N_3663);
nand U3816 (N_3816,N_3631,N_3723);
nand U3817 (N_3817,N_3791,N_3780);
nor U3818 (N_3818,N_3600,N_3681);
or U3819 (N_3819,N_3653,N_3733);
or U3820 (N_3820,N_3759,N_3739);
or U3821 (N_3821,N_3678,N_3732);
and U3822 (N_3822,N_3709,N_3749);
nand U3823 (N_3823,N_3720,N_3746);
or U3824 (N_3824,N_3696,N_3679);
nor U3825 (N_3825,N_3661,N_3683);
or U3826 (N_3826,N_3635,N_3790);
nand U3827 (N_3827,N_3770,N_3705);
nor U3828 (N_3828,N_3672,N_3698);
or U3829 (N_3829,N_3704,N_3662);
or U3830 (N_3830,N_3740,N_3616);
nand U3831 (N_3831,N_3687,N_3685);
nand U3832 (N_3832,N_3788,N_3715);
nand U3833 (N_3833,N_3638,N_3615);
nand U3834 (N_3834,N_3689,N_3718);
nand U3835 (N_3835,N_3659,N_3701);
or U3836 (N_3836,N_3714,N_3750);
or U3837 (N_3837,N_3633,N_3748);
nand U3838 (N_3838,N_3691,N_3729);
or U3839 (N_3839,N_3753,N_3747);
or U3840 (N_3840,N_3642,N_3652);
or U3841 (N_3841,N_3786,N_3664);
nand U3842 (N_3842,N_3617,N_3630);
nand U3843 (N_3843,N_3657,N_3756);
nand U3844 (N_3844,N_3618,N_3649);
or U3845 (N_3845,N_3675,N_3695);
and U3846 (N_3846,N_3609,N_3601);
and U3847 (N_3847,N_3722,N_3768);
nand U3848 (N_3848,N_3674,N_3673);
or U3849 (N_3849,N_3767,N_3724);
nor U3850 (N_3850,N_3744,N_3706);
and U3851 (N_3851,N_3669,N_3764);
and U3852 (N_3852,N_3620,N_3796);
or U3853 (N_3853,N_3680,N_3650);
nor U3854 (N_3854,N_3745,N_3632);
or U3855 (N_3855,N_3686,N_3752);
nor U3856 (N_3856,N_3707,N_3700);
and U3857 (N_3857,N_3625,N_3684);
nand U3858 (N_3858,N_3742,N_3658);
nand U3859 (N_3859,N_3713,N_3622);
and U3860 (N_3860,N_3668,N_3604);
nor U3861 (N_3861,N_3793,N_3797);
nor U3862 (N_3862,N_3734,N_3711);
nand U3863 (N_3863,N_3654,N_3644);
and U3864 (N_3864,N_3725,N_3634);
nor U3865 (N_3865,N_3602,N_3751);
nand U3866 (N_3866,N_3773,N_3741);
or U3867 (N_3867,N_3671,N_3757);
and U3868 (N_3868,N_3623,N_3606);
or U3869 (N_3869,N_3670,N_3641);
and U3870 (N_3870,N_3798,N_3610);
and U3871 (N_3871,N_3726,N_3693);
xor U3872 (N_3872,N_3636,N_3665);
xnor U3873 (N_3873,N_3735,N_3775);
nor U3874 (N_3874,N_3692,N_3667);
nand U3875 (N_3875,N_3666,N_3637);
or U3876 (N_3876,N_3789,N_3771);
and U3877 (N_3877,N_3762,N_3716);
or U3878 (N_3878,N_3651,N_3607);
and U3879 (N_3879,N_3656,N_3660);
xnor U3880 (N_3880,N_3721,N_3690);
and U3881 (N_3881,N_3777,N_3688);
nand U3882 (N_3882,N_3655,N_3778);
nand U3883 (N_3883,N_3792,N_3703);
nor U3884 (N_3884,N_3731,N_3682);
or U3885 (N_3885,N_3772,N_3603);
or U3886 (N_3886,N_3784,N_3766);
nor U3887 (N_3887,N_3677,N_3774);
nand U3888 (N_3888,N_3710,N_3761);
and U3889 (N_3889,N_3728,N_3613);
nand U3890 (N_3890,N_3758,N_3763);
or U3891 (N_3891,N_3776,N_3754);
and U3892 (N_3892,N_3760,N_3783);
and U3893 (N_3893,N_3736,N_3605);
and U3894 (N_3894,N_3708,N_3640);
or U3895 (N_3895,N_3648,N_3699);
and U3896 (N_3896,N_3769,N_3627);
nand U3897 (N_3897,N_3755,N_3621);
or U3898 (N_3898,N_3781,N_3765);
nand U3899 (N_3899,N_3645,N_3787);
nand U3900 (N_3900,N_3772,N_3780);
nor U3901 (N_3901,N_3605,N_3661);
and U3902 (N_3902,N_3622,N_3602);
and U3903 (N_3903,N_3796,N_3793);
nor U3904 (N_3904,N_3710,N_3777);
nand U3905 (N_3905,N_3677,N_3725);
or U3906 (N_3906,N_3651,N_3740);
and U3907 (N_3907,N_3790,N_3612);
nor U3908 (N_3908,N_3730,N_3640);
and U3909 (N_3909,N_3736,N_3659);
nor U3910 (N_3910,N_3604,N_3705);
or U3911 (N_3911,N_3623,N_3793);
nor U3912 (N_3912,N_3663,N_3772);
or U3913 (N_3913,N_3694,N_3799);
or U3914 (N_3914,N_3694,N_3660);
nor U3915 (N_3915,N_3764,N_3712);
xor U3916 (N_3916,N_3678,N_3660);
or U3917 (N_3917,N_3681,N_3606);
or U3918 (N_3918,N_3670,N_3692);
nand U3919 (N_3919,N_3682,N_3669);
and U3920 (N_3920,N_3793,N_3672);
and U3921 (N_3921,N_3753,N_3702);
nor U3922 (N_3922,N_3616,N_3750);
nor U3923 (N_3923,N_3628,N_3612);
and U3924 (N_3924,N_3721,N_3792);
or U3925 (N_3925,N_3747,N_3622);
xor U3926 (N_3926,N_3609,N_3716);
nor U3927 (N_3927,N_3732,N_3755);
and U3928 (N_3928,N_3616,N_3715);
or U3929 (N_3929,N_3688,N_3684);
nor U3930 (N_3930,N_3616,N_3719);
nor U3931 (N_3931,N_3702,N_3641);
and U3932 (N_3932,N_3625,N_3738);
nor U3933 (N_3933,N_3702,N_3788);
nor U3934 (N_3934,N_3642,N_3600);
nand U3935 (N_3935,N_3621,N_3690);
or U3936 (N_3936,N_3637,N_3644);
nor U3937 (N_3937,N_3790,N_3705);
or U3938 (N_3938,N_3792,N_3757);
nand U3939 (N_3939,N_3633,N_3614);
or U3940 (N_3940,N_3687,N_3731);
nor U3941 (N_3941,N_3608,N_3628);
or U3942 (N_3942,N_3711,N_3736);
nand U3943 (N_3943,N_3605,N_3791);
and U3944 (N_3944,N_3686,N_3673);
nor U3945 (N_3945,N_3776,N_3758);
nor U3946 (N_3946,N_3658,N_3727);
nor U3947 (N_3947,N_3693,N_3760);
or U3948 (N_3948,N_3770,N_3609);
or U3949 (N_3949,N_3787,N_3639);
or U3950 (N_3950,N_3781,N_3729);
and U3951 (N_3951,N_3728,N_3765);
nand U3952 (N_3952,N_3703,N_3783);
and U3953 (N_3953,N_3653,N_3629);
nor U3954 (N_3954,N_3759,N_3645);
or U3955 (N_3955,N_3698,N_3786);
and U3956 (N_3956,N_3655,N_3681);
or U3957 (N_3957,N_3690,N_3698);
or U3958 (N_3958,N_3745,N_3624);
and U3959 (N_3959,N_3697,N_3789);
nand U3960 (N_3960,N_3671,N_3691);
or U3961 (N_3961,N_3780,N_3724);
nand U3962 (N_3962,N_3786,N_3666);
or U3963 (N_3963,N_3668,N_3602);
or U3964 (N_3964,N_3763,N_3619);
nor U3965 (N_3965,N_3651,N_3695);
nor U3966 (N_3966,N_3789,N_3648);
nor U3967 (N_3967,N_3700,N_3673);
and U3968 (N_3968,N_3679,N_3629);
and U3969 (N_3969,N_3659,N_3757);
and U3970 (N_3970,N_3794,N_3724);
nor U3971 (N_3971,N_3702,N_3793);
nand U3972 (N_3972,N_3714,N_3767);
and U3973 (N_3973,N_3664,N_3649);
or U3974 (N_3974,N_3760,N_3764);
and U3975 (N_3975,N_3726,N_3770);
or U3976 (N_3976,N_3715,N_3704);
and U3977 (N_3977,N_3799,N_3603);
nand U3978 (N_3978,N_3713,N_3742);
and U3979 (N_3979,N_3690,N_3731);
or U3980 (N_3980,N_3678,N_3666);
and U3981 (N_3981,N_3736,N_3644);
or U3982 (N_3982,N_3788,N_3795);
and U3983 (N_3983,N_3699,N_3760);
nand U3984 (N_3984,N_3734,N_3730);
and U3985 (N_3985,N_3629,N_3638);
nand U3986 (N_3986,N_3790,N_3711);
xor U3987 (N_3987,N_3602,N_3699);
xor U3988 (N_3988,N_3692,N_3621);
and U3989 (N_3989,N_3672,N_3786);
nand U3990 (N_3990,N_3627,N_3749);
or U3991 (N_3991,N_3717,N_3692);
nand U3992 (N_3992,N_3786,N_3622);
or U3993 (N_3993,N_3680,N_3658);
or U3994 (N_3994,N_3626,N_3607);
or U3995 (N_3995,N_3601,N_3700);
nor U3996 (N_3996,N_3736,N_3741);
nor U3997 (N_3997,N_3646,N_3654);
or U3998 (N_3998,N_3686,N_3610);
nor U3999 (N_3999,N_3623,N_3614);
or U4000 (N_4000,N_3898,N_3923);
nor U4001 (N_4001,N_3930,N_3817);
or U4002 (N_4002,N_3880,N_3889);
nand U4003 (N_4003,N_3944,N_3849);
nor U4004 (N_4004,N_3801,N_3978);
or U4005 (N_4005,N_3818,N_3934);
or U4006 (N_4006,N_3883,N_3848);
nand U4007 (N_4007,N_3825,N_3999);
nor U4008 (N_4008,N_3949,N_3840);
and U4009 (N_4009,N_3933,N_3813);
and U4010 (N_4010,N_3920,N_3969);
and U4011 (N_4011,N_3902,N_3987);
and U4012 (N_4012,N_3986,N_3876);
nand U4013 (N_4013,N_3894,N_3867);
nor U4014 (N_4014,N_3841,N_3870);
nor U4015 (N_4015,N_3937,N_3907);
nand U4016 (N_4016,N_3882,N_3895);
nor U4017 (N_4017,N_3928,N_3808);
nand U4018 (N_4018,N_3957,N_3862);
or U4019 (N_4019,N_3822,N_3942);
nand U4020 (N_4020,N_3991,N_3909);
or U4021 (N_4021,N_3858,N_3886);
nor U4022 (N_4022,N_3828,N_3956);
nor U4023 (N_4023,N_3989,N_3900);
nor U4024 (N_4024,N_3976,N_3963);
nor U4025 (N_4025,N_3852,N_3936);
or U4026 (N_4026,N_3981,N_3885);
or U4027 (N_4027,N_3940,N_3854);
nand U4028 (N_4028,N_3827,N_3853);
or U4029 (N_4029,N_3977,N_3831);
or U4030 (N_4030,N_3918,N_3872);
and U4031 (N_4031,N_3863,N_3924);
nand U4032 (N_4032,N_3819,N_3985);
and U4033 (N_4033,N_3922,N_3892);
and U4034 (N_4034,N_3806,N_3905);
or U4035 (N_4035,N_3802,N_3800);
nor U4036 (N_4036,N_3998,N_3954);
and U4037 (N_4037,N_3973,N_3943);
and U4038 (N_4038,N_3856,N_3916);
or U4039 (N_4039,N_3997,N_3869);
and U4040 (N_4040,N_3829,N_3821);
or U4041 (N_4041,N_3903,N_3958);
or U4042 (N_4042,N_3845,N_3955);
nor U4043 (N_4043,N_3877,N_3935);
nor U4044 (N_4044,N_3993,N_3893);
or U4045 (N_4045,N_3995,N_3988);
nor U4046 (N_4046,N_3833,N_3910);
nand U4047 (N_4047,N_3938,N_3899);
and U4048 (N_4048,N_3911,N_3824);
and U4049 (N_4049,N_3932,N_3915);
or U4050 (N_4050,N_3951,N_3803);
and U4051 (N_4051,N_3809,N_3891);
nand U4052 (N_4052,N_3908,N_3971);
nor U4053 (N_4053,N_3979,N_3921);
or U4054 (N_4054,N_3835,N_3887);
nand U4055 (N_4055,N_3834,N_3855);
or U4056 (N_4056,N_3975,N_3990);
or U4057 (N_4057,N_3996,N_3890);
and U4058 (N_4058,N_3967,N_3980);
nand U4059 (N_4059,N_3873,N_3945);
and U4060 (N_4060,N_3866,N_3917);
or U4061 (N_4061,N_3811,N_3972);
and U4062 (N_4062,N_3865,N_3875);
nand U4063 (N_4063,N_3914,N_3896);
nor U4064 (N_4064,N_3857,N_3844);
nor U4065 (N_4065,N_3837,N_3970);
or U4066 (N_4066,N_3859,N_3839);
or U4067 (N_4067,N_3964,N_3847);
and U4068 (N_4068,N_3906,N_3947);
and U4069 (N_4069,N_3929,N_3982);
or U4070 (N_4070,N_3953,N_3874);
or U4071 (N_4071,N_3807,N_3836);
and U4072 (N_4072,N_3812,N_3919);
nand U4073 (N_4073,N_3832,N_3966);
xnor U4074 (N_4074,N_3960,N_3884);
and U4075 (N_4075,N_3961,N_3974);
or U4076 (N_4076,N_3950,N_3994);
nand U4077 (N_4077,N_3897,N_3959);
or U4078 (N_4078,N_3925,N_3814);
nor U4079 (N_4079,N_3968,N_3842);
or U4080 (N_4080,N_3983,N_3913);
nand U4081 (N_4081,N_3815,N_3965);
nand U4082 (N_4082,N_3962,N_3846);
nor U4083 (N_4083,N_3843,N_3912);
xnor U4084 (N_4084,N_3850,N_3931);
or U4085 (N_4085,N_3823,N_3868);
and U4086 (N_4086,N_3826,N_3864);
and U4087 (N_4087,N_3838,N_3984);
nor U4088 (N_4088,N_3888,N_3804);
xnor U4089 (N_4089,N_3926,N_3820);
nor U4090 (N_4090,N_3901,N_3927);
xor U4091 (N_4091,N_3881,N_3851);
nor U4092 (N_4092,N_3992,N_3871);
nand U4093 (N_4093,N_3948,N_3810);
or U4094 (N_4094,N_3816,N_3946);
and U4095 (N_4095,N_3952,N_3805);
nand U4096 (N_4096,N_3904,N_3879);
nor U4097 (N_4097,N_3941,N_3878);
xnor U4098 (N_4098,N_3830,N_3861);
or U4099 (N_4099,N_3860,N_3939);
nand U4100 (N_4100,N_3862,N_3971);
or U4101 (N_4101,N_3940,N_3924);
or U4102 (N_4102,N_3920,N_3863);
nand U4103 (N_4103,N_3836,N_3937);
and U4104 (N_4104,N_3834,N_3804);
nor U4105 (N_4105,N_3841,N_3837);
or U4106 (N_4106,N_3866,N_3835);
nor U4107 (N_4107,N_3983,N_3869);
nor U4108 (N_4108,N_3853,N_3897);
nor U4109 (N_4109,N_3807,N_3893);
and U4110 (N_4110,N_3985,N_3854);
nor U4111 (N_4111,N_3908,N_3893);
or U4112 (N_4112,N_3831,N_3815);
and U4113 (N_4113,N_3968,N_3997);
and U4114 (N_4114,N_3811,N_3849);
nor U4115 (N_4115,N_3866,N_3845);
nand U4116 (N_4116,N_3941,N_3914);
and U4117 (N_4117,N_3806,N_3949);
nor U4118 (N_4118,N_3939,N_3879);
or U4119 (N_4119,N_3839,N_3964);
and U4120 (N_4120,N_3865,N_3858);
nor U4121 (N_4121,N_3854,N_3947);
nand U4122 (N_4122,N_3973,N_3921);
xor U4123 (N_4123,N_3984,N_3936);
or U4124 (N_4124,N_3821,N_3878);
or U4125 (N_4125,N_3964,N_3811);
or U4126 (N_4126,N_3957,N_3931);
nor U4127 (N_4127,N_3827,N_3982);
nor U4128 (N_4128,N_3812,N_3918);
or U4129 (N_4129,N_3833,N_3965);
nand U4130 (N_4130,N_3808,N_3972);
and U4131 (N_4131,N_3964,N_3976);
xnor U4132 (N_4132,N_3994,N_3836);
and U4133 (N_4133,N_3889,N_3985);
or U4134 (N_4134,N_3977,N_3921);
or U4135 (N_4135,N_3813,N_3977);
nor U4136 (N_4136,N_3858,N_3950);
and U4137 (N_4137,N_3828,N_3993);
nand U4138 (N_4138,N_3876,N_3893);
nand U4139 (N_4139,N_3841,N_3873);
or U4140 (N_4140,N_3897,N_3879);
or U4141 (N_4141,N_3802,N_3883);
nand U4142 (N_4142,N_3889,N_3933);
and U4143 (N_4143,N_3805,N_3806);
nor U4144 (N_4144,N_3822,N_3873);
nor U4145 (N_4145,N_3832,N_3834);
nand U4146 (N_4146,N_3934,N_3954);
nand U4147 (N_4147,N_3975,N_3985);
or U4148 (N_4148,N_3845,N_3863);
or U4149 (N_4149,N_3966,N_3918);
xnor U4150 (N_4150,N_3922,N_3976);
nand U4151 (N_4151,N_3830,N_3923);
or U4152 (N_4152,N_3817,N_3868);
nand U4153 (N_4153,N_3805,N_3988);
nand U4154 (N_4154,N_3960,N_3802);
nor U4155 (N_4155,N_3865,N_3883);
nand U4156 (N_4156,N_3954,N_3955);
and U4157 (N_4157,N_3829,N_3816);
nand U4158 (N_4158,N_3860,N_3920);
or U4159 (N_4159,N_3857,N_3893);
nand U4160 (N_4160,N_3989,N_3830);
nand U4161 (N_4161,N_3861,N_3828);
and U4162 (N_4162,N_3995,N_3854);
or U4163 (N_4163,N_3870,N_3859);
nor U4164 (N_4164,N_3939,N_3922);
nor U4165 (N_4165,N_3856,N_3950);
nand U4166 (N_4166,N_3985,N_3853);
nand U4167 (N_4167,N_3970,N_3816);
or U4168 (N_4168,N_3993,N_3974);
and U4169 (N_4169,N_3914,N_3999);
nand U4170 (N_4170,N_3974,N_3801);
xor U4171 (N_4171,N_3862,N_3901);
or U4172 (N_4172,N_3814,N_3918);
nor U4173 (N_4173,N_3839,N_3814);
or U4174 (N_4174,N_3931,N_3871);
and U4175 (N_4175,N_3962,N_3918);
or U4176 (N_4176,N_3948,N_3917);
nor U4177 (N_4177,N_3807,N_3949);
nor U4178 (N_4178,N_3993,N_3908);
nor U4179 (N_4179,N_3998,N_3923);
nor U4180 (N_4180,N_3848,N_3937);
or U4181 (N_4181,N_3941,N_3929);
or U4182 (N_4182,N_3861,N_3911);
or U4183 (N_4183,N_3929,N_3894);
nand U4184 (N_4184,N_3836,N_3879);
or U4185 (N_4185,N_3881,N_3853);
nor U4186 (N_4186,N_3868,N_3847);
nand U4187 (N_4187,N_3838,N_3813);
and U4188 (N_4188,N_3911,N_3837);
nand U4189 (N_4189,N_3832,N_3902);
and U4190 (N_4190,N_3912,N_3826);
or U4191 (N_4191,N_3890,N_3801);
or U4192 (N_4192,N_3870,N_3930);
nor U4193 (N_4193,N_3972,N_3979);
nand U4194 (N_4194,N_3951,N_3800);
nand U4195 (N_4195,N_3947,N_3926);
and U4196 (N_4196,N_3852,N_3861);
nand U4197 (N_4197,N_3865,N_3829);
and U4198 (N_4198,N_3924,N_3983);
or U4199 (N_4199,N_3945,N_3823);
nand U4200 (N_4200,N_4033,N_4104);
nand U4201 (N_4201,N_4002,N_4196);
and U4202 (N_4202,N_4011,N_4082);
nand U4203 (N_4203,N_4112,N_4094);
nor U4204 (N_4204,N_4019,N_4168);
or U4205 (N_4205,N_4118,N_4126);
nand U4206 (N_4206,N_4023,N_4108);
and U4207 (N_4207,N_4180,N_4163);
nor U4208 (N_4208,N_4065,N_4184);
nor U4209 (N_4209,N_4187,N_4006);
nand U4210 (N_4210,N_4154,N_4115);
and U4211 (N_4211,N_4151,N_4063);
nor U4212 (N_4212,N_4067,N_4077);
or U4213 (N_4213,N_4164,N_4027);
nor U4214 (N_4214,N_4092,N_4128);
and U4215 (N_4215,N_4093,N_4156);
nand U4216 (N_4216,N_4125,N_4143);
nand U4217 (N_4217,N_4012,N_4040);
or U4218 (N_4218,N_4064,N_4142);
or U4219 (N_4219,N_4121,N_4129);
nand U4220 (N_4220,N_4001,N_4017);
nor U4221 (N_4221,N_4042,N_4056);
or U4222 (N_4222,N_4100,N_4049);
nand U4223 (N_4223,N_4198,N_4197);
nor U4224 (N_4224,N_4024,N_4188);
nand U4225 (N_4225,N_4003,N_4034);
nand U4226 (N_4226,N_4075,N_4171);
or U4227 (N_4227,N_4014,N_4052);
or U4228 (N_4228,N_4130,N_4181);
or U4229 (N_4229,N_4140,N_4069);
nand U4230 (N_4230,N_4183,N_4105);
or U4231 (N_4231,N_4098,N_4095);
nor U4232 (N_4232,N_4070,N_4160);
nand U4233 (N_4233,N_4195,N_4020);
nand U4234 (N_4234,N_4127,N_4159);
and U4235 (N_4235,N_4177,N_4178);
nor U4236 (N_4236,N_4037,N_4057);
nor U4237 (N_4237,N_4016,N_4035);
and U4238 (N_4238,N_4007,N_4120);
or U4239 (N_4239,N_4138,N_4041);
nand U4240 (N_4240,N_4144,N_4149);
and U4241 (N_4241,N_4074,N_4122);
or U4242 (N_4242,N_4146,N_4038);
and U4243 (N_4243,N_4123,N_4060);
nand U4244 (N_4244,N_4000,N_4134);
or U4245 (N_4245,N_4175,N_4044);
nand U4246 (N_4246,N_4072,N_4114);
or U4247 (N_4247,N_4097,N_4008);
nor U4248 (N_4248,N_4119,N_4021);
nand U4249 (N_4249,N_4109,N_4106);
or U4250 (N_4250,N_4145,N_4152);
and U4251 (N_4251,N_4148,N_4046);
nor U4252 (N_4252,N_4107,N_4111);
nand U4253 (N_4253,N_4135,N_4172);
and U4254 (N_4254,N_4158,N_4132);
and U4255 (N_4255,N_4078,N_4084);
nand U4256 (N_4256,N_4031,N_4058);
or U4257 (N_4257,N_4102,N_4173);
nand U4258 (N_4258,N_4045,N_4174);
or U4259 (N_4259,N_4055,N_4062);
and U4260 (N_4260,N_4085,N_4194);
or U4261 (N_4261,N_4089,N_4015);
or U4262 (N_4262,N_4090,N_4088);
or U4263 (N_4263,N_4170,N_4185);
nand U4264 (N_4264,N_4166,N_4147);
or U4265 (N_4265,N_4080,N_4054);
and U4266 (N_4266,N_4068,N_4022);
nand U4267 (N_4267,N_4073,N_4169);
nand U4268 (N_4268,N_4009,N_4199);
and U4269 (N_4269,N_4076,N_4179);
nor U4270 (N_4270,N_4039,N_4059);
or U4271 (N_4271,N_4167,N_4189);
nand U4272 (N_4272,N_4028,N_4137);
nand U4273 (N_4273,N_4004,N_4186);
or U4274 (N_4274,N_4013,N_4182);
nor U4275 (N_4275,N_4005,N_4066);
nand U4276 (N_4276,N_4133,N_4025);
nand U4277 (N_4277,N_4139,N_4116);
nor U4278 (N_4278,N_4165,N_4155);
xor U4279 (N_4279,N_4081,N_4029);
nand U4280 (N_4280,N_4176,N_4190);
or U4281 (N_4281,N_4048,N_4061);
nor U4282 (N_4282,N_4141,N_4053);
and U4283 (N_4283,N_4083,N_4051);
or U4284 (N_4284,N_4157,N_4103);
or U4285 (N_4285,N_4030,N_4026);
nand U4286 (N_4286,N_4086,N_4071);
nor U4287 (N_4287,N_4050,N_4192);
nor U4288 (N_4288,N_4047,N_4161);
nand U4289 (N_4289,N_4191,N_4110);
nor U4290 (N_4290,N_4136,N_4124);
nor U4291 (N_4291,N_4162,N_4036);
and U4292 (N_4292,N_4193,N_4091);
nor U4293 (N_4293,N_4099,N_4113);
and U4294 (N_4294,N_4096,N_4131);
nand U4295 (N_4295,N_4117,N_4010);
nand U4296 (N_4296,N_4079,N_4150);
and U4297 (N_4297,N_4087,N_4032);
or U4298 (N_4298,N_4101,N_4043);
nor U4299 (N_4299,N_4153,N_4018);
nor U4300 (N_4300,N_4072,N_4187);
nor U4301 (N_4301,N_4019,N_4059);
nor U4302 (N_4302,N_4079,N_4107);
nand U4303 (N_4303,N_4067,N_4120);
and U4304 (N_4304,N_4007,N_4148);
nand U4305 (N_4305,N_4104,N_4145);
nand U4306 (N_4306,N_4178,N_4149);
and U4307 (N_4307,N_4101,N_4158);
nand U4308 (N_4308,N_4193,N_4135);
and U4309 (N_4309,N_4151,N_4047);
nand U4310 (N_4310,N_4153,N_4022);
and U4311 (N_4311,N_4030,N_4196);
or U4312 (N_4312,N_4166,N_4195);
or U4313 (N_4313,N_4164,N_4141);
or U4314 (N_4314,N_4158,N_4170);
xnor U4315 (N_4315,N_4030,N_4050);
or U4316 (N_4316,N_4097,N_4013);
nand U4317 (N_4317,N_4177,N_4152);
and U4318 (N_4318,N_4170,N_4070);
and U4319 (N_4319,N_4062,N_4164);
nor U4320 (N_4320,N_4186,N_4064);
nor U4321 (N_4321,N_4027,N_4058);
nor U4322 (N_4322,N_4074,N_4011);
or U4323 (N_4323,N_4091,N_4038);
and U4324 (N_4324,N_4186,N_4078);
nor U4325 (N_4325,N_4057,N_4114);
nor U4326 (N_4326,N_4144,N_4071);
nor U4327 (N_4327,N_4075,N_4027);
and U4328 (N_4328,N_4034,N_4117);
nor U4329 (N_4329,N_4002,N_4061);
nor U4330 (N_4330,N_4034,N_4016);
nor U4331 (N_4331,N_4165,N_4146);
nand U4332 (N_4332,N_4028,N_4084);
and U4333 (N_4333,N_4005,N_4177);
nand U4334 (N_4334,N_4023,N_4111);
or U4335 (N_4335,N_4092,N_4088);
nor U4336 (N_4336,N_4154,N_4016);
nor U4337 (N_4337,N_4095,N_4178);
nand U4338 (N_4338,N_4134,N_4002);
or U4339 (N_4339,N_4040,N_4097);
nor U4340 (N_4340,N_4025,N_4080);
nand U4341 (N_4341,N_4177,N_4190);
xor U4342 (N_4342,N_4019,N_4009);
nor U4343 (N_4343,N_4120,N_4056);
and U4344 (N_4344,N_4166,N_4018);
and U4345 (N_4345,N_4097,N_4171);
or U4346 (N_4346,N_4177,N_4103);
and U4347 (N_4347,N_4144,N_4197);
and U4348 (N_4348,N_4174,N_4005);
nor U4349 (N_4349,N_4087,N_4081);
nand U4350 (N_4350,N_4153,N_4038);
xor U4351 (N_4351,N_4150,N_4047);
nand U4352 (N_4352,N_4110,N_4049);
xor U4353 (N_4353,N_4059,N_4011);
nand U4354 (N_4354,N_4172,N_4177);
nand U4355 (N_4355,N_4170,N_4056);
or U4356 (N_4356,N_4092,N_4070);
nand U4357 (N_4357,N_4162,N_4138);
or U4358 (N_4358,N_4180,N_4130);
nor U4359 (N_4359,N_4088,N_4060);
or U4360 (N_4360,N_4195,N_4060);
nor U4361 (N_4361,N_4041,N_4071);
or U4362 (N_4362,N_4045,N_4052);
or U4363 (N_4363,N_4091,N_4103);
nand U4364 (N_4364,N_4148,N_4056);
nand U4365 (N_4365,N_4033,N_4141);
nand U4366 (N_4366,N_4130,N_4023);
nor U4367 (N_4367,N_4162,N_4116);
or U4368 (N_4368,N_4002,N_4087);
and U4369 (N_4369,N_4118,N_4119);
and U4370 (N_4370,N_4180,N_4145);
or U4371 (N_4371,N_4001,N_4119);
nand U4372 (N_4372,N_4082,N_4091);
nor U4373 (N_4373,N_4117,N_4079);
or U4374 (N_4374,N_4026,N_4080);
nor U4375 (N_4375,N_4092,N_4032);
nor U4376 (N_4376,N_4058,N_4190);
or U4377 (N_4377,N_4107,N_4018);
nor U4378 (N_4378,N_4160,N_4185);
nor U4379 (N_4379,N_4069,N_4102);
or U4380 (N_4380,N_4198,N_4065);
and U4381 (N_4381,N_4036,N_4199);
nor U4382 (N_4382,N_4122,N_4002);
nor U4383 (N_4383,N_4167,N_4098);
xor U4384 (N_4384,N_4059,N_4016);
and U4385 (N_4385,N_4140,N_4058);
nor U4386 (N_4386,N_4150,N_4195);
xor U4387 (N_4387,N_4106,N_4051);
nand U4388 (N_4388,N_4081,N_4152);
and U4389 (N_4389,N_4148,N_4031);
or U4390 (N_4390,N_4002,N_4034);
nor U4391 (N_4391,N_4147,N_4021);
nor U4392 (N_4392,N_4112,N_4176);
or U4393 (N_4393,N_4119,N_4117);
and U4394 (N_4394,N_4023,N_4000);
or U4395 (N_4395,N_4110,N_4015);
and U4396 (N_4396,N_4103,N_4036);
nor U4397 (N_4397,N_4116,N_4058);
nor U4398 (N_4398,N_4007,N_4096);
and U4399 (N_4399,N_4109,N_4120);
nand U4400 (N_4400,N_4270,N_4349);
nand U4401 (N_4401,N_4380,N_4222);
nor U4402 (N_4402,N_4309,N_4343);
and U4403 (N_4403,N_4387,N_4345);
nand U4404 (N_4404,N_4214,N_4333);
nand U4405 (N_4405,N_4238,N_4303);
nor U4406 (N_4406,N_4285,N_4229);
nor U4407 (N_4407,N_4227,N_4286);
nor U4408 (N_4408,N_4255,N_4302);
nor U4409 (N_4409,N_4208,N_4379);
and U4410 (N_4410,N_4396,N_4213);
nand U4411 (N_4411,N_4278,N_4252);
and U4412 (N_4412,N_4246,N_4293);
nor U4413 (N_4413,N_4305,N_4217);
and U4414 (N_4414,N_4319,N_4267);
and U4415 (N_4415,N_4381,N_4326);
and U4416 (N_4416,N_4323,N_4236);
nor U4417 (N_4417,N_4220,N_4315);
nand U4418 (N_4418,N_4391,N_4261);
nand U4419 (N_4419,N_4389,N_4276);
nand U4420 (N_4420,N_4228,N_4274);
nand U4421 (N_4421,N_4316,N_4353);
and U4422 (N_4422,N_4271,N_4307);
nor U4423 (N_4423,N_4280,N_4386);
nand U4424 (N_4424,N_4321,N_4288);
and U4425 (N_4425,N_4248,N_4364);
and U4426 (N_4426,N_4292,N_4335);
or U4427 (N_4427,N_4283,N_4240);
or U4428 (N_4428,N_4210,N_4395);
or U4429 (N_4429,N_4269,N_4397);
nand U4430 (N_4430,N_4212,N_4332);
nand U4431 (N_4431,N_4231,N_4350);
or U4432 (N_4432,N_4223,N_4264);
nand U4433 (N_4433,N_4233,N_4275);
or U4434 (N_4434,N_4203,N_4361);
nor U4435 (N_4435,N_4291,N_4357);
and U4436 (N_4436,N_4363,N_4378);
nand U4437 (N_4437,N_4304,N_4394);
nor U4438 (N_4438,N_4254,N_4341);
or U4439 (N_4439,N_4358,N_4221);
or U4440 (N_4440,N_4297,N_4294);
and U4441 (N_4441,N_4237,N_4310);
nor U4442 (N_4442,N_4211,N_4336);
and U4443 (N_4443,N_4247,N_4268);
or U4444 (N_4444,N_4334,N_4360);
nor U4445 (N_4445,N_4317,N_4262);
xor U4446 (N_4446,N_4322,N_4253);
nand U4447 (N_4447,N_4354,N_4249);
nand U4448 (N_4448,N_4299,N_4351);
nor U4449 (N_4449,N_4306,N_4205);
nor U4450 (N_4450,N_4340,N_4352);
and U4451 (N_4451,N_4202,N_4375);
and U4452 (N_4452,N_4235,N_4344);
nor U4453 (N_4453,N_4216,N_4372);
nor U4454 (N_4454,N_4384,N_4392);
and U4455 (N_4455,N_4298,N_4281);
and U4456 (N_4456,N_4284,N_4279);
nor U4457 (N_4457,N_4245,N_4242);
nor U4458 (N_4458,N_4265,N_4257);
nor U4459 (N_4459,N_4277,N_4215);
nor U4460 (N_4460,N_4328,N_4390);
nor U4461 (N_4461,N_4383,N_4218);
nand U4462 (N_4462,N_4243,N_4226);
or U4463 (N_4463,N_4347,N_4201);
or U4464 (N_4464,N_4377,N_4331);
or U4465 (N_4465,N_4374,N_4393);
nor U4466 (N_4466,N_4368,N_4399);
and U4467 (N_4467,N_4366,N_4365);
xor U4468 (N_4468,N_4337,N_4263);
xnor U4469 (N_4469,N_4206,N_4325);
and U4470 (N_4470,N_4287,N_4209);
nor U4471 (N_4471,N_4200,N_4327);
or U4472 (N_4472,N_4272,N_4355);
and U4473 (N_4473,N_4258,N_4388);
nor U4474 (N_4474,N_4311,N_4266);
nor U4475 (N_4475,N_4232,N_4382);
and U4476 (N_4476,N_4373,N_4385);
nor U4477 (N_4477,N_4225,N_4290);
nand U4478 (N_4478,N_4359,N_4224);
or U4479 (N_4479,N_4313,N_4348);
nor U4480 (N_4480,N_4250,N_4234);
nand U4481 (N_4481,N_4207,N_4239);
nor U4482 (N_4482,N_4362,N_4273);
nand U4483 (N_4483,N_4219,N_4376);
and U4484 (N_4484,N_4295,N_4371);
nor U4485 (N_4485,N_4301,N_4339);
xnor U4486 (N_4486,N_4260,N_4312);
nand U4487 (N_4487,N_4330,N_4346);
nand U4488 (N_4488,N_4369,N_4244);
or U4489 (N_4489,N_4296,N_4398);
and U4490 (N_4490,N_4367,N_4300);
or U4491 (N_4491,N_4256,N_4308);
and U4492 (N_4492,N_4282,N_4342);
and U4493 (N_4493,N_4324,N_4314);
nand U4494 (N_4494,N_4318,N_4230);
and U4495 (N_4495,N_4320,N_4370);
and U4496 (N_4496,N_4251,N_4289);
or U4497 (N_4497,N_4329,N_4241);
nor U4498 (N_4498,N_4338,N_4259);
or U4499 (N_4499,N_4356,N_4204);
nand U4500 (N_4500,N_4263,N_4257);
and U4501 (N_4501,N_4329,N_4343);
nand U4502 (N_4502,N_4213,N_4264);
nand U4503 (N_4503,N_4318,N_4379);
or U4504 (N_4504,N_4310,N_4366);
or U4505 (N_4505,N_4319,N_4357);
or U4506 (N_4506,N_4309,N_4291);
and U4507 (N_4507,N_4315,N_4328);
or U4508 (N_4508,N_4373,N_4340);
nor U4509 (N_4509,N_4397,N_4204);
nor U4510 (N_4510,N_4261,N_4390);
and U4511 (N_4511,N_4386,N_4246);
or U4512 (N_4512,N_4328,N_4323);
or U4513 (N_4513,N_4220,N_4242);
and U4514 (N_4514,N_4233,N_4266);
nand U4515 (N_4515,N_4299,N_4234);
nor U4516 (N_4516,N_4230,N_4325);
and U4517 (N_4517,N_4220,N_4225);
nand U4518 (N_4518,N_4392,N_4368);
nor U4519 (N_4519,N_4229,N_4231);
or U4520 (N_4520,N_4320,N_4215);
or U4521 (N_4521,N_4279,N_4312);
nand U4522 (N_4522,N_4345,N_4389);
nand U4523 (N_4523,N_4368,N_4209);
nand U4524 (N_4524,N_4277,N_4219);
or U4525 (N_4525,N_4290,N_4222);
or U4526 (N_4526,N_4300,N_4290);
or U4527 (N_4527,N_4332,N_4250);
nand U4528 (N_4528,N_4225,N_4204);
nor U4529 (N_4529,N_4258,N_4356);
nor U4530 (N_4530,N_4245,N_4352);
nor U4531 (N_4531,N_4249,N_4226);
and U4532 (N_4532,N_4281,N_4367);
nand U4533 (N_4533,N_4384,N_4382);
or U4534 (N_4534,N_4202,N_4348);
nor U4535 (N_4535,N_4266,N_4284);
or U4536 (N_4536,N_4308,N_4241);
or U4537 (N_4537,N_4229,N_4307);
or U4538 (N_4538,N_4397,N_4373);
nand U4539 (N_4539,N_4251,N_4353);
and U4540 (N_4540,N_4343,N_4277);
and U4541 (N_4541,N_4284,N_4325);
and U4542 (N_4542,N_4239,N_4224);
and U4543 (N_4543,N_4389,N_4323);
or U4544 (N_4544,N_4285,N_4378);
or U4545 (N_4545,N_4361,N_4228);
nand U4546 (N_4546,N_4335,N_4260);
or U4547 (N_4547,N_4343,N_4397);
and U4548 (N_4548,N_4322,N_4316);
or U4549 (N_4549,N_4394,N_4207);
and U4550 (N_4550,N_4254,N_4201);
and U4551 (N_4551,N_4265,N_4218);
and U4552 (N_4552,N_4345,N_4347);
nor U4553 (N_4553,N_4238,N_4273);
or U4554 (N_4554,N_4320,N_4360);
or U4555 (N_4555,N_4326,N_4225);
nand U4556 (N_4556,N_4231,N_4230);
nand U4557 (N_4557,N_4232,N_4312);
or U4558 (N_4558,N_4359,N_4395);
or U4559 (N_4559,N_4342,N_4293);
nand U4560 (N_4560,N_4356,N_4274);
nand U4561 (N_4561,N_4287,N_4300);
nor U4562 (N_4562,N_4329,N_4392);
nor U4563 (N_4563,N_4316,N_4341);
xor U4564 (N_4564,N_4233,N_4287);
and U4565 (N_4565,N_4227,N_4387);
nor U4566 (N_4566,N_4235,N_4226);
and U4567 (N_4567,N_4311,N_4393);
and U4568 (N_4568,N_4304,N_4237);
nor U4569 (N_4569,N_4377,N_4277);
nand U4570 (N_4570,N_4386,N_4277);
nand U4571 (N_4571,N_4312,N_4340);
and U4572 (N_4572,N_4294,N_4370);
nor U4573 (N_4573,N_4244,N_4344);
and U4574 (N_4574,N_4354,N_4327);
nor U4575 (N_4575,N_4287,N_4397);
nand U4576 (N_4576,N_4278,N_4251);
nor U4577 (N_4577,N_4372,N_4277);
nand U4578 (N_4578,N_4362,N_4357);
nor U4579 (N_4579,N_4307,N_4249);
nor U4580 (N_4580,N_4392,N_4243);
nor U4581 (N_4581,N_4318,N_4275);
nand U4582 (N_4582,N_4365,N_4334);
and U4583 (N_4583,N_4303,N_4361);
or U4584 (N_4584,N_4313,N_4264);
or U4585 (N_4585,N_4229,N_4360);
nor U4586 (N_4586,N_4339,N_4272);
nor U4587 (N_4587,N_4298,N_4367);
nor U4588 (N_4588,N_4233,N_4232);
nor U4589 (N_4589,N_4373,N_4378);
or U4590 (N_4590,N_4399,N_4207);
nor U4591 (N_4591,N_4296,N_4250);
and U4592 (N_4592,N_4303,N_4227);
or U4593 (N_4593,N_4399,N_4262);
nor U4594 (N_4594,N_4253,N_4224);
and U4595 (N_4595,N_4326,N_4293);
or U4596 (N_4596,N_4243,N_4343);
nor U4597 (N_4597,N_4212,N_4389);
nor U4598 (N_4598,N_4201,N_4385);
or U4599 (N_4599,N_4217,N_4313);
or U4600 (N_4600,N_4546,N_4528);
or U4601 (N_4601,N_4593,N_4450);
nand U4602 (N_4602,N_4422,N_4427);
nor U4603 (N_4603,N_4409,N_4440);
xor U4604 (N_4604,N_4584,N_4442);
nand U4605 (N_4605,N_4502,N_4437);
or U4606 (N_4606,N_4478,N_4581);
nor U4607 (N_4607,N_4536,N_4544);
and U4608 (N_4608,N_4460,N_4432);
nor U4609 (N_4609,N_4557,N_4413);
and U4610 (N_4610,N_4482,N_4529);
xnor U4611 (N_4611,N_4596,N_4564);
and U4612 (N_4612,N_4516,N_4507);
nor U4613 (N_4613,N_4588,N_4512);
nor U4614 (N_4614,N_4477,N_4594);
nor U4615 (N_4615,N_4453,N_4591);
nand U4616 (N_4616,N_4447,N_4423);
nand U4617 (N_4617,N_4540,N_4424);
or U4618 (N_4618,N_4467,N_4506);
nor U4619 (N_4619,N_4524,N_4587);
and U4620 (N_4620,N_4403,N_4439);
and U4621 (N_4621,N_4518,N_4459);
and U4622 (N_4622,N_4497,N_4574);
nor U4623 (N_4623,N_4575,N_4498);
nand U4624 (N_4624,N_4465,N_4515);
nor U4625 (N_4625,N_4547,N_4463);
and U4626 (N_4626,N_4405,N_4471);
nand U4627 (N_4627,N_4457,N_4435);
or U4628 (N_4628,N_4476,N_4579);
or U4629 (N_4629,N_4425,N_4549);
xor U4630 (N_4630,N_4599,N_4472);
nand U4631 (N_4631,N_4452,N_4551);
or U4632 (N_4632,N_4531,N_4486);
and U4633 (N_4633,N_4415,N_4508);
nor U4634 (N_4634,N_4525,N_4475);
nor U4635 (N_4635,N_4573,N_4541);
nor U4636 (N_4636,N_4441,N_4590);
and U4637 (N_4637,N_4481,N_4500);
or U4638 (N_4638,N_4499,N_4426);
or U4639 (N_4639,N_4402,N_4454);
nor U4640 (N_4640,N_4410,N_4533);
nor U4641 (N_4641,N_4535,N_4434);
or U4642 (N_4642,N_4532,N_4495);
nand U4643 (N_4643,N_4578,N_4561);
nor U4644 (N_4644,N_4462,N_4530);
nor U4645 (N_4645,N_4568,N_4404);
nand U4646 (N_4646,N_4414,N_4451);
nor U4647 (N_4647,N_4534,N_4586);
nor U4648 (N_4648,N_4443,N_4567);
nand U4649 (N_4649,N_4565,N_4513);
or U4650 (N_4650,N_4455,N_4537);
and U4651 (N_4651,N_4558,N_4519);
nor U4652 (N_4652,N_4461,N_4577);
nand U4653 (N_4653,N_4542,N_4485);
and U4654 (N_4654,N_4416,N_4521);
or U4655 (N_4655,N_4583,N_4469);
nand U4656 (N_4656,N_4444,N_4527);
nor U4657 (N_4657,N_4582,N_4449);
nand U4658 (N_4658,N_4493,N_4563);
or U4659 (N_4659,N_4548,N_4552);
or U4660 (N_4660,N_4448,N_4474);
nor U4661 (N_4661,N_4496,N_4401);
or U4662 (N_4662,N_4554,N_4420);
nor U4663 (N_4663,N_4458,N_4419);
nand U4664 (N_4664,N_4456,N_4411);
nand U4665 (N_4665,N_4494,N_4501);
or U4666 (N_4666,N_4572,N_4514);
and U4667 (N_4667,N_4464,N_4580);
xnor U4668 (N_4668,N_4592,N_4569);
or U4669 (N_4669,N_4429,N_4509);
nor U4670 (N_4670,N_4491,N_4492);
nor U4671 (N_4671,N_4445,N_4560);
nor U4672 (N_4672,N_4484,N_4517);
and U4673 (N_4673,N_4553,N_4487);
nor U4674 (N_4674,N_4408,N_4522);
and U4675 (N_4675,N_4488,N_4559);
nor U4676 (N_4676,N_4407,N_4412);
nor U4677 (N_4677,N_4421,N_4585);
nand U4678 (N_4678,N_4566,N_4545);
nor U4679 (N_4679,N_4430,N_4490);
nor U4680 (N_4680,N_4428,N_4595);
and U4681 (N_4681,N_4479,N_4483);
and U4682 (N_4682,N_4418,N_4597);
nand U4683 (N_4683,N_4436,N_4550);
nor U4684 (N_4684,N_4526,N_4468);
nand U4685 (N_4685,N_4510,N_4598);
or U4686 (N_4686,N_4406,N_4504);
nor U4687 (N_4687,N_4470,N_4589);
nor U4688 (N_4688,N_4523,N_4539);
or U4689 (N_4689,N_4511,N_4400);
or U4690 (N_4690,N_4571,N_4489);
nor U4691 (N_4691,N_4520,N_4503);
or U4692 (N_4692,N_4417,N_4562);
nand U4693 (N_4693,N_4576,N_4473);
or U4694 (N_4694,N_4480,N_4466);
nor U4695 (N_4695,N_4555,N_4570);
and U4696 (N_4696,N_4431,N_4538);
nor U4697 (N_4697,N_4505,N_4446);
nor U4698 (N_4698,N_4433,N_4543);
and U4699 (N_4699,N_4556,N_4438);
nand U4700 (N_4700,N_4545,N_4483);
or U4701 (N_4701,N_4434,N_4517);
or U4702 (N_4702,N_4495,N_4529);
nor U4703 (N_4703,N_4418,N_4596);
and U4704 (N_4704,N_4435,N_4466);
or U4705 (N_4705,N_4567,N_4580);
and U4706 (N_4706,N_4521,N_4514);
nor U4707 (N_4707,N_4429,N_4524);
or U4708 (N_4708,N_4498,N_4447);
or U4709 (N_4709,N_4408,N_4579);
nand U4710 (N_4710,N_4503,N_4463);
nand U4711 (N_4711,N_4563,N_4568);
nand U4712 (N_4712,N_4457,N_4594);
nor U4713 (N_4713,N_4591,N_4510);
nor U4714 (N_4714,N_4485,N_4467);
nand U4715 (N_4715,N_4458,N_4585);
xnor U4716 (N_4716,N_4445,N_4499);
or U4717 (N_4717,N_4447,N_4541);
and U4718 (N_4718,N_4474,N_4511);
or U4719 (N_4719,N_4598,N_4561);
nor U4720 (N_4720,N_4444,N_4521);
nor U4721 (N_4721,N_4400,N_4498);
and U4722 (N_4722,N_4451,N_4529);
nand U4723 (N_4723,N_4403,N_4538);
or U4724 (N_4724,N_4530,N_4580);
and U4725 (N_4725,N_4475,N_4567);
or U4726 (N_4726,N_4551,N_4483);
nand U4727 (N_4727,N_4421,N_4523);
nor U4728 (N_4728,N_4415,N_4489);
or U4729 (N_4729,N_4500,N_4560);
or U4730 (N_4730,N_4501,N_4453);
nor U4731 (N_4731,N_4512,N_4533);
nand U4732 (N_4732,N_4471,N_4412);
or U4733 (N_4733,N_4485,N_4525);
and U4734 (N_4734,N_4470,N_4555);
or U4735 (N_4735,N_4414,N_4597);
and U4736 (N_4736,N_4461,N_4490);
nand U4737 (N_4737,N_4539,N_4527);
or U4738 (N_4738,N_4510,N_4535);
xor U4739 (N_4739,N_4553,N_4522);
nand U4740 (N_4740,N_4456,N_4596);
or U4741 (N_4741,N_4460,N_4420);
nor U4742 (N_4742,N_4506,N_4444);
and U4743 (N_4743,N_4518,N_4427);
or U4744 (N_4744,N_4566,N_4471);
nand U4745 (N_4745,N_4493,N_4491);
and U4746 (N_4746,N_4565,N_4463);
or U4747 (N_4747,N_4537,N_4536);
nor U4748 (N_4748,N_4407,N_4441);
nor U4749 (N_4749,N_4545,N_4448);
and U4750 (N_4750,N_4576,N_4589);
and U4751 (N_4751,N_4491,N_4428);
nand U4752 (N_4752,N_4529,N_4472);
and U4753 (N_4753,N_4430,N_4535);
or U4754 (N_4754,N_4455,N_4539);
and U4755 (N_4755,N_4468,N_4551);
nand U4756 (N_4756,N_4443,N_4429);
and U4757 (N_4757,N_4453,N_4556);
and U4758 (N_4758,N_4423,N_4427);
nor U4759 (N_4759,N_4465,N_4477);
and U4760 (N_4760,N_4581,N_4468);
nand U4761 (N_4761,N_4531,N_4483);
nor U4762 (N_4762,N_4584,N_4519);
nor U4763 (N_4763,N_4556,N_4420);
nand U4764 (N_4764,N_4591,N_4416);
nand U4765 (N_4765,N_4565,N_4566);
and U4766 (N_4766,N_4464,N_4458);
or U4767 (N_4767,N_4542,N_4594);
nor U4768 (N_4768,N_4576,N_4447);
nand U4769 (N_4769,N_4414,N_4401);
or U4770 (N_4770,N_4537,N_4550);
nand U4771 (N_4771,N_4462,N_4549);
nor U4772 (N_4772,N_4596,N_4451);
or U4773 (N_4773,N_4582,N_4503);
nor U4774 (N_4774,N_4427,N_4503);
and U4775 (N_4775,N_4432,N_4500);
and U4776 (N_4776,N_4420,N_4551);
nor U4777 (N_4777,N_4519,N_4467);
or U4778 (N_4778,N_4490,N_4587);
nand U4779 (N_4779,N_4524,N_4480);
or U4780 (N_4780,N_4448,N_4432);
and U4781 (N_4781,N_4574,N_4573);
or U4782 (N_4782,N_4460,N_4466);
nand U4783 (N_4783,N_4566,N_4540);
or U4784 (N_4784,N_4434,N_4411);
nor U4785 (N_4785,N_4465,N_4522);
nor U4786 (N_4786,N_4522,N_4505);
and U4787 (N_4787,N_4514,N_4543);
and U4788 (N_4788,N_4508,N_4550);
and U4789 (N_4789,N_4510,N_4435);
or U4790 (N_4790,N_4542,N_4499);
nor U4791 (N_4791,N_4476,N_4416);
or U4792 (N_4792,N_4563,N_4576);
or U4793 (N_4793,N_4420,N_4599);
nor U4794 (N_4794,N_4595,N_4403);
and U4795 (N_4795,N_4542,N_4538);
nand U4796 (N_4796,N_4428,N_4570);
or U4797 (N_4797,N_4536,N_4528);
or U4798 (N_4798,N_4525,N_4425);
and U4799 (N_4799,N_4554,N_4573);
nand U4800 (N_4800,N_4696,N_4789);
nand U4801 (N_4801,N_4766,N_4711);
or U4802 (N_4802,N_4604,N_4701);
nand U4803 (N_4803,N_4762,N_4690);
or U4804 (N_4804,N_4695,N_4652);
nor U4805 (N_4805,N_4760,N_4645);
nand U4806 (N_4806,N_4644,N_4691);
or U4807 (N_4807,N_4758,N_4640);
or U4808 (N_4808,N_4735,N_4602);
or U4809 (N_4809,N_4631,N_4608);
or U4810 (N_4810,N_4717,N_4779);
nor U4811 (N_4811,N_4739,N_4646);
and U4812 (N_4812,N_4719,N_4728);
nand U4813 (N_4813,N_4630,N_4681);
and U4814 (N_4814,N_4693,N_4712);
and U4815 (N_4815,N_4751,N_4622);
and U4816 (N_4816,N_4685,N_4707);
nand U4817 (N_4817,N_4659,N_4749);
or U4818 (N_4818,N_4674,N_4725);
and U4819 (N_4819,N_4692,N_4768);
nand U4820 (N_4820,N_4651,N_4661);
or U4821 (N_4821,N_4752,N_4729);
nand U4822 (N_4822,N_4638,N_4670);
or U4823 (N_4823,N_4654,N_4764);
and U4824 (N_4824,N_4618,N_4731);
and U4825 (N_4825,N_4778,N_4665);
or U4826 (N_4826,N_4628,N_4675);
or U4827 (N_4827,N_4641,N_4797);
nor U4828 (N_4828,N_4703,N_4677);
nor U4829 (N_4829,N_4656,N_4611);
nor U4830 (N_4830,N_4600,N_4747);
nor U4831 (N_4831,N_4720,N_4738);
nor U4832 (N_4832,N_4698,N_4775);
nand U4833 (N_4833,N_4607,N_4671);
nand U4834 (N_4834,N_4759,N_4649);
and U4835 (N_4835,N_4705,N_4774);
nor U4836 (N_4836,N_4754,N_4723);
or U4837 (N_4837,N_4669,N_4730);
and U4838 (N_4838,N_4613,N_4635);
nand U4839 (N_4839,N_4697,N_4684);
or U4840 (N_4840,N_4624,N_4744);
nor U4841 (N_4841,N_4704,N_4794);
and U4842 (N_4842,N_4773,N_4786);
nor U4843 (N_4843,N_4666,N_4658);
nand U4844 (N_4844,N_4603,N_4627);
nand U4845 (N_4845,N_4615,N_4715);
and U4846 (N_4846,N_4662,N_4629);
nor U4847 (N_4847,N_4643,N_4795);
or U4848 (N_4848,N_4626,N_4612);
or U4849 (N_4849,N_4702,N_4726);
nor U4850 (N_4850,N_4799,N_4741);
and U4851 (N_4851,N_4625,N_4755);
nor U4852 (N_4852,N_4706,N_4672);
and U4853 (N_4853,N_4714,N_4791);
nand U4854 (N_4854,N_4761,N_4756);
nor U4855 (N_4855,N_4718,N_4614);
nand U4856 (N_4856,N_4694,N_4660);
and U4857 (N_4857,N_4753,N_4687);
and U4858 (N_4858,N_4683,N_4619);
and U4859 (N_4859,N_4617,N_4686);
or U4860 (N_4860,N_4732,N_4777);
nor U4861 (N_4861,N_4734,N_4650);
nor U4862 (N_4862,N_4606,N_4637);
nand U4863 (N_4863,N_4689,N_4616);
nand U4864 (N_4864,N_4748,N_4710);
nand U4865 (N_4865,N_4776,N_4743);
nand U4866 (N_4866,N_4796,N_4745);
nand U4867 (N_4867,N_4639,N_4634);
or U4868 (N_4868,N_4699,N_4657);
nor U4869 (N_4869,N_4721,N_4772);
or U4870 (N_4870,N_4724,N_4655);
nor U4871 (N_4871,N_4667,N_4716);
or U4872 (N_4872,N_4788,N_4623);
nor U4873 (N_4873,N_4700,N_4785);
and U4874 (N_4874,N_4784,N_4722);
nor U4875 (N_4875,N_4601,N_4632);
nor U4876 (N_4876,N_4680,N_4708);
nor U4877 (N_4877,N_4678,N_4781);
and U4878 (N_4878,N_4757,N_4767);
and U4879 (N_4879,N_4787,N_4620);
or U4880 (N_4880,N_4780,N_4769);
nor U4881 (N_4881,N_4647,N_4798);
nand U4882 (N_4882,N_4770,N_4653);
nor U4883 (N_4883,N_4790,N_4782);
nand U4884 (N_4884,N_4742,N_4642);
or U4885 (N_4885,N_4727,N_4750);
nor U4886 (N_4886,N_4621,N_4733);
nor U4887 (N_4887,N_4610,N_4771);
nand U4888 (N_4888,N_4792,N_4740);
nand U4889 (N_4889,N_4688,N_4609);
and U4890 (N_4890,N_4783,N_4663);
nand U4891 (N_4891,N_4736,N_4633);
or U4892 (N_4892,N_4648,N_4793);
nor U4893 (N_4893,N_4737,N_4673);
nor U4894 (N_4894,N_4679,N_4664);
or U4895 (N_4895,N_4709,N_4713);
nand U4896 (N_4896,N_4746,N_4765);
and U4897 (N_4897,N_4668,N_4763);
or U4898 (N_4898,N_4676,N_4682);
nor U4899 (N_4899,N_4636,N_4605);
nand U4900 (N_4900,N_4777,N_4760);
or U4901 (N_4901,N_4605,N_4689);
and U4902 (N_4902,N_4751,N_4726);
or U4903 (N_4903,N_4724,N_4729);
nor U4904 (N_4904,N_4667,N_4796);
or U4905 (N_4905,N_4630,N_4621);
and U4906 (N_4906,N_4688,N_4799);
or U4907 (N_4907,N_4742,N_4639);
or U4908 (N_4908,N_4772,N_4773);
or U4909 (N_4909,N_4769,N_4622);
nor U4910 (N_4910,N_4777,N_4639);
nor U4911 (N_4911,N_4673,N_4662);
and U4912 (N_4912,N_4602,N_4648);
or U4913 (N_4913,N_4665,N_4666);
nor U4914 (N_4914,N_4614,N_4644);
nand U4915 (N_4915,N_4764,N_4623);
and U4916 (N_4916,N_4629,N_4626);
or U4917 (N_4917,N_4656,N_4691);
and U4918 (N_4918,N_4645,N_4624);
nor U4919 (N_4919,N_4681,N_4774);
or U4920 (N_4920,N_4646,N_4797);
nand U4921 (N_4921,N_4609,N_4607);
nor U4922 (N_4922,N_4704,N_4601);
and U4923 (N_4923,N_4790,N_4653);
and U4924 (N_4924,N_4698,N_4617);
nor U4925 (N_4925,N_4610,N_4684);
nor U4926 (N_4926,N_4633,N_4705);
nand U4927 (N_4927,N_4746,N_4645);
and U4928 (N_4928,N_4654,N_4666);
and U4929 (N_4929,N_4787,N_4746);
nand U4930 (N_4930,N_4791,N_4659);
nand U4931 (N_4931,N_4765,N_4718);
nand U4932 (N_4932,N_4660,N_4676);
nand U4933 (N_4933,N_4662,N_4746);
and U4934 (N_4934,N_4656,N_4790);
or U4935 (N_4935,N_4761,N_4680);
and U4936 (N_4936,N_4773,N_4611);
and U4937 (N_4937,N_4720,N_4618);
or U4938 (N_4938,N_4723,N_4624);
nor U4939 (N_4939,N_4633,N_4794);
or U4940 (N_4940,N_4696,N_4705);
and U4941 (N_4941,N_4653,N_4610);
nor U4942 (N_4942,N_4761,N_4708);
and U4943 (N_4943,N_4753,N_4633);
nor U4944 (N_4944,N_4704,N_4764);
and U4945 (N_4945,N_4719,N_4757);
nand U4946 (N_4946,N_4628,N_4605);
nand U4947 (N_4947,N_4750,N_4772);
or U4948 (N_4948,N_4696,N_4719);
and U4949 (N_4949,N_4671,N_4676);
nor U4950 (N_4950,N_4799,N_4638);
and U4951 (N_4951,N_4752,N_4634);
nor U4952 (N_4952,N_4634,N_4748);
nor U4953 (N_4953,N_4786,N_4715);
nand U4954 (N_4954,N_4773,N_4654);
nand U4955 (N_4955,N_4778,N_4746);
or U4956 (N_4956,N_4681,N_4763);
nor U4957 (N_4957,N_4765,N_4655);
and U4958 (N_4958,N_4658,N_4753);
nand U4959 (N_4959,N_4769,N_4715);
and U4960 (N_4960,N_4709,N_4652);
and U4961 (N_4961,N_4768,N_4675);
and U4962 (N_4962,N_4715,N_4797);
and U4963 (N_4963,N_4669,N_4697);
nand U4964 (N_4964,N_4699,N_4770);
or U4965 (N_4965,N_4765,N_4616);
or U4966 (N_4966,N_4702,N_4765);
and U4967 (N_4967,N_4646,N_4667);
or U4968 (N_4968,N_4735,N_4691);
or U4969 (N_4969,N_4647,N_4616);
xor U4970 (N_4970,N_4639,N_4709);
or U4971 (N_4971,N_4605,N_4637);
and U4972 (N_4972,N_4753,N_4677);
or U4973 (N_4973,N_4637,N_4664);
or U4974 (N_4974,N_4779,N_4711);
nor U4975 (N_4975,N_4605,N_4615);
and U4976 (N_4976,N_4663,N_4668);
and U4977 (N_4977,N_4713,N_4708);
nand U4978 (N_4978,N_4746,N_4782);
nand U4979 (N_4979,N_4602,N_4694);
nand U4980 (N_4980,N_4603,N_4744);
nor U4981 (N_4981,N_4662,N_4618);
nor U4982 (N_4982,N_4613,N_4739);
and U4983 (N_4983,N_4752,N_4793);
or U4984 (N_4984,N_4679,N_4722);
nand U4985 (N_4985,N_4698,N_4767);
nor U4986 (N_4986,N_4790,N_4639);
nor U4987 (N_4987,N_4764,N_4631);
nand U4988 (N_4988,N_4754,N_4706);
and U4989 (N_4989,N_4718,N_4650);
and U4990 (N_4990,N_4646,N_4623);
or U4991 (N_4991,N_4699,N_4645);
nand U4992 (N_4992,N_4664,N_4687);
nand U4993 (N_4993,N_4695,N_4616);
nand U4994 (N_4994,N_4684,N_4672);
nor U4995 (N_4995,N_4629,N_4616);
nor U4996 (N_4996,N_4720,N_4654);
nor U4997 (N_4997,N_4675,N_4649);
nand U4998 (N_4998,N_4742,N_4647);
or U4999 (N_4999,N_4743,N_4796);
or UO_0 (O_0,N_4922,N_4921);
nand UO_1 (O_1,N_4833,N_4826);
xnor UO_2 (O_2,N_4946,N_4959);
nor UO_3 (O_3,N_4877,N_4857);
nand UO_4 (O_4,N_4881,N_4823);
nor UO_5 (O_5,N_4926,N_4927);
nor UO_6 (O_6,N_4804,N_4942);
or UO_7 (O_7,N_4909,N_4917);
nand UO_8 (O_8,N_4848,N_4847);
or UO_9 (O_9,N_4990,N_4969);
and UO_10 (O_10,N_4984,N_4965);
nand UO_11 (O_11,N_4979,N_4805);
and UO_12 (O_12,N_4824,N_4830);
nor UO_13 (O_13,N_4947,N_4944);
nor UO_14 (O_14,N_4836,N_4885);
and UO_15 (O_15,N_4800,N_4861);
nor UO_16 (O_16,N_4981,N_4970);
xor UO_17 (O_17,N_4991,N_4975);
or UO_18 (O_18,N_4980,N_4878);
or UO_19 (O_19,N_4825,N_4801);
nor UO_20 (O_20,N_4988,N_4894);
nor UO_21 (O_21,N_4892,N_4879);
nand UO_22 (O_22,N_4820,N_4956);
nor UO_23 (O_23,N_4943,N_4911);
nor UO_24 (O_24,N_4815,N_4950);
and UO_25 (O_25,N_4953,N_4871);
nand UO_26 (O_26,N_4949,N_4916);
nor UO_27 (O_27,N_4827,N_4872);
nand UO_28 (O_28,N_4995,N_4869);
and UO_29 (O_29,N_4841,N_4906);
or UO_30 (O_30,N_4868,N_4890);
nand UO_31 (O_31,N_4832,N_4889);
and UO_32 (O_32,N_4813,N_4985);
nand UO_33 (O_33,N_4802,N_4851);
or UO_34 (O_34,N_4971,N_4930);
or UO_35 (O_35,N_4849,N_4814);
and UO_36 (O_36,N_4838,N_4846);
and UO_37 (O_37,N_4888,N_4897);
and UO_38 (O_38,N_4997,N_4902);
and UO_39 (O_39,N_4937,N_4907);
nor UO_40 (O_40,N_4835,N_4931);
nor UO_41 (O_41,N_4912,N_4963);
and UO_42 (O_42,N_4929,N_4875);
nand UO_43 (O_43,N_4905,N_4915);
nor UO_44 (O_44,N_4962,N_4925);
nand UO_45 (O_45,N_4908,N_4874);
or UO_46 (O_46,N_4865,N_4939);
and UO_47 (O_47,N_4859,N_4831);
nand UO_48 (O_48,N_4863,N_4934);
nor UO_49 (O_49,N_4966,N_4961);
nand UO_50 (O_50,N_4935,N_4843);
and UO_51 (O_51,N_4895,N_4828);
or UO_52 (O_52,N_4996,N_4940);
or UO_53 (O_53,N_4948,N_4850);
nor UO_54 (O_54,N_4982,N_4900);
nor UO_55 (O_55,N_4919,N_4803);
nand UO_56 (O_56,N_4818,N_4977);
xor UO_57 (O_57,N_4834,N_4974);
nand UO_58 (O_58,N_4867,N_4913);
nand UO_59 (O_59,N_4910,N_4973);
nor UO_60 (O_60,N_4964,N_4840);
nor UO_61 (O_61,N_4992,N_4976);
and UO_62 (O_62,N_4967,N_4887);
nor UO_63 (O_63,N_4855,N_4936);
or UO_64 (O_64,N_4924,N_4958);
nand UO_65 (O_65,N_4938,N_4886);
nand UO_66 (O_66,N_4978,N_4852);
nor UO_67 (O_67,N_4812,N_4819);
or UO_68 (O_68,N_4941,N_4955);
nor UO_69 (O_69,N_4993,N_4808);
and UO_70 (O_70,N_4968,N_4870);
or UO_71 (O_71,N_4951,N_4989);
and UO_72 (O_72,N_4960,N_4904);
and UO_73 (O_73,N_4862,N_4896);
nand UO_74 (O_74,N_4839,N_4994);
nand UO_75 (O_75,N_4893,N_4883);
nor UO_76 (O_76,N_4918,N_4864);
nand UO_77 (O_77,N_4891,N_4933);
nand UO_78 (O_78,N_4829,N_4853);
and UO_79 (O_79,N_4957,N_4817);
and UO_80 (O_80,N_4858,N_4923);
or UO_81 (O_81,N_4809,N_4952);
or UO_82 (O_82,N_4860,N_4810);
nor UO_83 (O_83,N_4987,N_4903);
nor UO_84 (O_84,N_4856,N_4873);
nor UO_85 (O_85,N_4876,N_4914);
nor UO_86 (O_86,N_4882,N_4928);
nor UO_87 (O_87,N_4845,N_4920);
or UO_88 (O_88,N_4854,N_4972);
or UO_89 (O_89,N_4998,N_4837);
or UO_90 (O_90,N_4822,N_4811);
nor UO_91 (O_91,N_4983,N_4844);
and UO_92 (O_92,N_4986,N_4806);
or UO_93 (O_93,N_4816,N_4880);
or UO_94 (O_94,N_4898,N_4932);
or UO_95 (O_95,N_4866,N_4899);
and UO_96 (O_96,N_4842,N_4821);
or UO_97 (O_97,N_4901,N_4807);
nor UO_98 (O_98,N_4954,N_4999);
and UO_99 (O_99,N_4945,N_4884);
and UO_100 (O_100,N_4963,N_4860);
or UO_101 (O_101,N_4803,N_4904);
nand UO_102 (O_102,N_4801,N_4842);
and UO_103 (O_103,N_4985,N_4834);
or UO_104 (O_104,N_4874,N_4907);
nor UO_105 (O_105,N_4851,N_4894);
xor UO_106 (O_106,N_4911,N_4992);
and UO_107 (O_107,N_4903,N_4881);
nand UO_108 (O_108,N_4900,N_4846);
nor UO_109 (O_109,N_4936,N_4945);
and UO_110 (O_110,N_4935,N_4891);
or UO_111 (O_111,N_4812,N_4879);
and UO_112 (O_112,N_4984,N_4831);
nand UO_113 (O_113,N_4985,N_4998);
nand UO_114 (O_114,N_4823,N_4994);
nand UO_115 (O_115,N_4828,N_4901);
nand UO_116 (O_116,N_4821,N_4983);
nor UO_117 (O_117,N_4831,N_4900);
or UO_118 (O_118,N_4807,N_4830);
or UO_119 (O_119,N_4938,N_4976);
or UO_120 (O_120,N_4819,N_4944);
and UO_121 (O_121,N_4857,N_4958);
nand UO_122 (O_122,N_4926,N_4823);
and UO_123 (O_123,N_4947,N_4925);
and UO_124 (O_124,N_4826,N_4806);
nand UO_125 (O_125,N_4862,N_4995);
or UO_126 (O_126,N_4957,N_4910);
or UO_127 (O_127,N_4803,N_4913);
or UO_128 (O_128,N_4823,N_4861);
nand UO_129 (O_129,N_4824,N_4930);
nand UO_130 (O_130,N_4968,N_4806);
nor UO_131 (O_131,N_4880,N_4926);
or UO_132 (O_132,N_4840,N_4955);
nand UO_133 (O_133,N_4800,N_4968);
nor UO_134 (O_134,N_4998,N_4817);
nor UO_135 (O_135,N_4921,N_4973);
nor UO_136 (O_136,N_4866,N_4987);
nand UO_137 (O_137,N_4911,N_4808);
or UO_138 (O_138,N_4918,N_4810);
or UO_139 (O_139,N_4860,N_4965);
nor UO_140 (O_140,N_4873,N_4925);
or UO_141 (O_141,N_4828,N_4998);
nor UO_142 (O_142,N_4900,N_4830);
or UO_143 (O_143,N_4930,N_4842);
nand UO_144 (O_144,N_4894,N_4822);
nand UO_145 (O_145,N_4843,N_4998);
nand UO_146 (O_146,N_4870,N_4877);
or UO_147 (O_147,N_4901,N_4908);
and UO_148 (O_148,N_4949,N_4841);
and UO_149 (O_149,N_4891,N_4860);
or UO_150 (O_150,N_4833,N_4841);
nand UO_151 (O_151,N_4801,N_4919);
nor UO_152 (O_152,N_4840,N_4858);
nand UO_153 (O_153,N_4856,N_4945);
nor UO_154 (O_154,N_4852,N_4845);
nor UO_155 (O_155,N_4992,N_4805);
nand UO_156 (O_156,N_4816,N_4978);
and UO_157 (O_157,N_4822,N_4865);
nand UO_158 (O_158,N_4902,N_4970);
and UO_159 (O_159,N_4887,N_4867);
nand UO_160 (O_160,N_4877,N_4976);
nor UO_161 (O_161,N_4978,N_4926);
or UO_162 (O_162,N_4996,N_4992);
nor UO_163 (O_163,N_4877,N_4874);
and UO_164 (O_164,N_4905,N_4840);
nand UO_165 (O_165,N_4973,N_4985);
and UO_166 (O_166,N_4982,N_4953);
nand UO_167 (O_167,N_4989,N_4929);
and UO_168 (O_168,N_4884,N_4951);
nand UO_169 (O_169,N_4871,N_4952);
nor UO_170 (O_170,N_4938,N_4966);
and UO_171 (O_171,N_4881,N_4872);
and UO_172 (O_172,N_4989,N_4997);
and UO_173 (O_173,N_4835,N_4882);
nand UO_174 (O_174,N_4926,N_4928);
nand UO_175 (O_175,N_4870,N_4883);
or UO_176 (O_176,N_4969,N_4872);
nor UO_177 (O_177,N_4845,N_4860);
nand UO_178 (O_178,N_4865,N_4853);
and UO_179 (O_179,N_4891,N_4835);
or UO_180 (O_180,N_4980,N_4829);
nand UO_181 (O_181,N_4852,N_4862);
nand UO_182 (O_182,N_4878,N_4996);
nor UO_183 (O_183,N_4958,N_4910);
nor UO_184 (O_184,N_4884,N_4898);
or UO_185 (O_185,N_4941,N_4971);
and UO_186 (O_186,N_4954,N_4822);
or UO_187 (O_187,N_4940,N_4976);
nand UO_188 (O_188,N_4813,N_4866);
nor UO_189 (O_189,N_4935,N_4901);
or UO_190 (O_190,N_4812,N_4826);
or UO_191 (O_191,N_4958,N_4882);
or UO_192 (O_192,N_4826,N_4968);
nor UO_193 (O_193,N_4941,N_4965);
nor UO_194 (O_194,N_4894,N_4952);
or UO_195 (O_195,N_4956,N_4936);
xnor UO_196 (O_196,N_4968,N_4808);
or UO_197 (O_197,N_4932,N_4816);
or UO_198 (O_198,N_4956,N_4863);
or UO_199 (O_199,N_4858,N_4894);
or UO_200 (O_200,N_4889,N_4921);
and UO_201 (O_201,N_4869,N_4889);
nor UO_202 (O_202,N_4966,N_4994);
nor UO_203 (O_203,N_4843,N_4913);
nor UO_204 (O_204,N_4817,N_4858);
nand UO_205 (O_205,N_4961,N_4955);
nor UO_206 (O_206,N_4815,N_4980);
and UO_207 (O_207,N_4804,N_4892);
nand UO_208 (O_208,N_4950,N_4849);
nand UO_209 (O_209,N_4802,N_4818);
nor UO_210 (O_210,N_4913,N_4980);
nor UO_211 (O_211,N_4809,N_4908);
and UO_212 (O_212,N_4857,N_4828);
xor UO_213 (O_213,N_4877,N_4945);
nand UO_214 (O_214,N_4915,N_4857);
nand UO_215 (O_215,N_4841,N_4867);
or UO_216 (O_216,N_4960,N_4842);
or UO_217 (O_217,N_4823,N_4937);
xor UO_218 (O_218,N_4817,N_4906);
nand UO_219 (O_219,N_4860,N_4930);
or UO_220 (O_220,N_4883,N_4803);
or UO_221 (O_221,N_4934,N_4848);
or UO_222 (O_222,N_4993,N_4946);
and UO_223 (O_223,N_4801,N_4866);
and UO_224 (O_224,N_4856,N_4835);
and UO_225 (O_225,N_4811,N_4982);
and UO_226 (O_226,N_4966,N_4882);
nor UO_227 (O_227,N_4972,N_4839);
nand UO_228 (O_228,N_4826,N_4835);
and UO_229 (O_229,N_4942,N_4909);
and UO_230 (O_230,N_4979,N_4801);
nand UO_231 (O_231,N_4921,N_4865);
or UO_232 (O_232,N_4863,N_4938);
or UO_233 (O_233,N_4994,N_4848);
or UO_234 (O_234,N_4867,N_4920);
nor UO_235 (O_235,N_4843,N_4887);
or UO_236 (O_236,N_4803,N_4902);
or UO_237 (O_237,N_4840,N_4908);
nand UO_238 (O_238,N_4864,N_4993);
or UO_239 (O_239,N_4842,N_4866);
nand UO_240 (O_240,N_4813,N_4812);
and UO_241 (O_241,N_4913,N_4860);
and UO_242 (O_242,N_4914,N_4853);
or UO_243 (O_243,N_4863,N_4802);
nand UO_244 (O_244,N_4995,N_4998);
xor UO_245 (O_245,N_4826,N_4843);
or UO_246 (O_246,N_4851,N_4857);
nor UO_247 (O_247,N_4927,N_4887);
and UO_248 (O_248,N_4969,N_4925);
or UO_249 (O_249,N_4870,N_4855);
nor UO_250 (O_250,N_4945,N_4974);
nor UO_251 (O_251,N_4837,N_4997);
nand UO_252 (O_252,N_4815,N_4909);
and UO_253 (O_253,N_4887,N_4947);
or UO_254 (O_254,N_4926,N_4992);
nor UO_255 (O_255,N_4836,N_4978);
and UO_256 (O_256,N_4811,N_4838);
nand UO_257 (O_257,N_4867,N_4906);
nor UO_258 (O_258,N_4932,N_4808);
nor UO_259 (O_259,N_4983,N_4889);
nand UO_260 (O_260,N_4822,N_4806);
and UO_261 (O_261,N_4916,N_4991);
or UO_262 (O_262,N_4801,N_4812);
nand UO_263 (O_263,N_4839,N_4953);
or UO_264 (O_264,N_4997,N_4803);
nand UO_265 (O_265,N_4839,N_4903);
nor UO_266 (O_266,N_4858,N_4937);
xnor UO_267 (O_267,N_4977,N_4879);
nor UO_268 (O_268,N_4941,N_4815);
and UO_269 (O_269,N_4915,N_4975);
nor UO_270 (O_270,N_4805,N_4883);
or UO_271 (O_271,N_4963,N_4876);
nor UO_272 (O_272,N_4958,N_4907);
nor UO_273 (O_273,N_4963,N_4826);
or UO_274 (O_274,N_4938,N_4968);
nor UO_275 (O_275,N_4876,N_4919);
nand UO_276 (O_276,N_4872,N_4948);
or UO_277 (O_277,N_4898,N_4905);
or UO_278 (O_278,N_4814,N_4990);
nor UO_279 (O_279,N_4954,N_4902);
nor UO_280 (O_280,N_4973,N_4898);
nor UO_281 (O_281,N_4976,N_4838);
nand UO_282 (O_282,N_4810,N_4914);
nand UO_283 (O_283,N_4832,N_4892);
or UO_284 (O_284,N_4984,N_4943);
nand UO_285 (O_285,N_4864,N_4979);
nand UO_286 (O_286,N_4947,N_4978);
nor UO_287 (O_287,N_4817,N_4900);
nor UO_288 (O_288,N_4961,N_4811);
or UO_289 (O_289,N_4883,N_4980);
and UO_290 (O_290,N_4980,N_4916);
or UO_291 (O_291,N_4990,N_4882);
or UO_292 (O_292,N_4955,N_4949);
and UO_293 (O_293,N_4847,N_4896);
or UO_294 (O_294,N_4981,N_4858);
nand UO_295 (O_295,N_4932,N_4802);
nor UO_296 (O_296,N_4810,N_4826);
nand UO_297 (O_297,N_4884,N_4858);
and UO_298 (O_298,N_4812,N_4811);
nor UO_299 (O_299,N_4806,N_4889);
nand UO_300 (O_300,N_4917,N_4922);
or UO_301 (O_301,N_4830,N_4986);
nand UO_302 (O_302,N_4985,N_4978);
or UO_303 (O_303,N_4940,N_4861);
nor UO_304 (O_304,N_4887,N_4808);
or UO_305 (O_305,N_4898,N_4862);
nand UO_306 (O_306,N_4995,N_4812);
nor UO_307 (O_307,N_4954,N_4916);
and UO_308 (O_308,N_4832,N_4831);
or UO_309 (O_309,N_4931,N_4937);
nand UO_310 (O_310,N_4962,N_4995);
or UO_311 (O_311,N_4801,N_4938);
nand UO_312 (O_312,N_4965,N_4980);
nand UO_313 (O_313,N_4915,N_4957);
nor UO_314 (O_314,N_4979,N_4955);
and UO_315 (O_315,N_4926,N_4987);
nor UO_316 (O_316,N_4850,N_4817);
nand UO_317 (O_317,N_4862,N_4861);
or UO_318 (O_318,N_4841,N_4808);
nor UO_319 (O_319,N_4923,N_4979);
or UO_320 (O_320,N_4845,N_4877);
and UO_321 (O_321,N_4866,N_4820);
or UO_322 (O_322,N_4947,N_4907);
nand UO_323 (O_323,N_4915,N_4886);
nand UO_324 (O_324,N_4932,N_4857);
nand UO_325 (O_325,N_4928,N_4920);
nor UO_326 (O_326,N_4848,N_4932);
or UO_327 (O_327,N_4876,N_4921);
and UO_328 (O_328,N_4856,N_4959);
nand UO_329 (O_329,N_4915,N_4953);
and UO_330 (O_330,N_4825,N_4945);
and UO_331 (O_331,N_4924,N_4935);
nand UO_332 (O_332,N_4878,N_4897);
xnor UO_333 (O_333,N_4921,N_4919);
and UO_334 (O_334,N_4970,N_4915);
and UO_335 (O_335,N_4924,N_4845);
and UO_336 (O_336,N_4971,N_4812);
nand UO_337 (O_337,N_4942,N_4997);
nor UO_338 (O_338,N_4977,N_4987);
or UO_339 (O_339,N_4812,N_4952);
or UO_340 (O_340,N_4811,N_4895);
and UO_341 (O_341,N_4881,N_4969);
nor UO_342 (O_342,N_4858,N_4912);
or UO_343 (O_343,N_4843,N_4946);
nand UO_344 (O_344,N_4937,N_4898);
nor UO_345 (O_345,N_4971,N_4996);
and UO_346 (O_346,N_4835,N_4972);
or UO_347 (O_347,N_4931,N_4896);
nand UO_348 (O_348,N_4853,N_4952);
nand UO_349 (O_349,N_4912,N_4937);
or UO_350 (O_350,N_4955,N_4945);
nor UO_351 (O_351,N_4828,N_4999);
nor UO_352 (O_352,N_4841,N_4893);
or UO_353 (O_353,N_4930,N_4889);
nand UO_354 (O_354,N_4935,N_4914);
nand UO_355 (O_355,N_4949,N_4883);
or UO_356 (O_356,N_4877,N_4912);
nand UO_357 (O_357,N_4807,N_4871);
nor UO_358 (O_358,N_4987,N_4917);
or UO_359 (O_359,N_4888,N_4927);
or UO_360 (O_360,N_4960,N_4888);
nand UO_361 (O_361,N_4970,N_4872);
or UO_362 (O_362,N_4833,N_4905);
and UO_363 (O_363,N_4984,N_4812);
nand UO_364 (O_364,N_4824,N_4935);
and UO_365 (O_365,N_4970,N_4822);
or UO_366 (O_366,N_4913,N_4908);
and UO_367 (O_367,N_4818,N_4994);
nor UO_368 (O_368,N_4917,N_4954);
or UO_369 (O_369,N_4800,N_4910);
or UO_370 (O_370,N_4844,N_4918);
nor UO_371 (O_371,N_4805,N_4968);
and UO_372 (O_372,N_4876,N_4997);
nor UO_373 (O_373,N_4921,N_4923);
nor UO_374 (O_374,N_4990,N_4877);
nor UO_375 (O_375,N_4805,N_4907);
nand UO_376 (O_376,N_4864,N_4897);
or UO_377 (O_377,N_4880,N_4938);
nand UO_378 (O_378,N_4882,N_4840);
nand UO_379 (O_379,N_4961,N_4938);
nand UO_380 (O_380,N_4860,N_4970);
nor UO_381 (O_381,N_4987,N_4931);
nor UO_382 (O_382,N_4910,N_4815);
nand UO_383 (O_383,N_4827,N_4961);
nor UO_384 (O_384,N_4869,N_4830);
and UO_385 (O_385,N_4988,N_4919);
nor UO_386 (O_386,N_4872,N_4880);
or UO_387 (O_387,N_4868,N_4880);
and UO_388 (O_388,N_4933,N_4909);
nor UO_389 (O_389,N_4996,N_4880);
nand UO_390 (O_390,N_4900,N_4838);
and UO_391 (O_391,N_4900,N_4801);
and UO_392 (O_392,N_4908,N_4839);
nand UO_393 (O_393,N_4822,N_4852);
nor UO_394 (O_394,N_4944,N_4835);
nor UO_395 (O_395,N_4914,N_4998);
and UO_396 (O_396,N_4881,N_4854);
nor UO_397 (O_397,N_4899,N_4909);
and UO_398 (O_398,N_4947,N_4982);
nor UO_399 (O_399,N_4946,N_4954);
and UO_400 (O_400,N_4992,N_4822);
and UO_401 (O_401,N_4828,N_4994);
or UO_402 (O_402,N_4976,N_4970);
nor UO_403 (O_403,N_4943,N_4981);
and UO_404 (O_404,N_4814,N_4994);
nor UO_405 (O_405,N_4874,N_4925);
and UO_406 (O_406,N_4870,N_4918);
nand UO_407 (O_407,N_4931,N_4860);
and UO_408 (O_408,N_4986,N_4815);
nand UO_409 (O_409,N_4932,N_4878);
and UO_410 (O_410,N_4990,N_4857);
and UO_411 (O_411,N_4885,N_4955);
nor UO_412 (O_412,N_4908,N_4886);
or UO_413 (O_413,N_4905,N_4882);
nor UO_414 (O_414,N_4804,N_4843);
nor UO_415 (O_415,N_4988,N_4935);
or UO_416 (O_416,N_4854,N_4908);
nand UO_417 (O_417,N_4977,N_4855);
nand UO_418 (O_418,N_4828,N_4876);
nand UO_419 (O_419,N_4947,N_4933);
nor UO_420 (O_420,N_4970,N_4836);
and UO_421 (O_421,N_4905,N_4831);
nor UO_422 (O_422,N_4916,N_4979);
and UO_423 (O_423,N_4901,N_4848);
nand UO_424 (O_424,N_4871,N_4982);
nand UO_425 (O_425,N_4872,N_4997);
nand UO_426 (O_426,N_4904,N_4912);
or UO_427 (O_427,N_4829,N_4804);
and UO_428 (O_428,N_4813,N_4829);
nand UO_429 (O_429,N_4958,N_4898);
and UO_430 (O_430,N_4807,N_4847);
and UO_431 (O_431,N_4915,N_4849);
nand UO_432 (O_432,N_4828,N_4838);
and UO_433 (O_433,N_4888,N_4801);
nor UO_434 (O_434,N_4955,N_4974);
and UO_435 (O_435,N_4980,N_4902);
and UO_436 (O_436,N_4929,N_4838);
and UO_437 (O_437,N_4839,N_4886);
or UO_438 (O_438,N_4862,N_4882);
or UO_439 (O_439,N_4804,N_4931);
xor UO_440 (O_440,N_4848,N_4963);
nand UO_441 (O_441,N_4924,N_4811);
nor UO_442 (O_442,N_4800,N_4977);
nor UO_443 (O_443,N_4985,N_4820);
or UO_444 (O_444,N_4941,N_4991);
and UO_445 (O_445,N_4804,N_4911);
nor UO_446 (O_446,N_4889,N_4845);
or UO_447 (O_447,N_4894,N_4923);
xnor UO_448 (O_448,N_4900,N_4808);
nor UO_449 (O_449,N_4843,N_4870);
and UO_450 (O_450,N_4917,N_4970);
nand UO_451 (O_451,N_4842,N_4989);
nor UO_452 (O_452,N_4974,N_4941);
nand UO_453 (O_453,N_4841,N_4851);
and UO_454 (O_454,N_4982,N_4821);
or UO_455 (O_455,N_4823,N_4871);
nand UO_456 (O_456,N_4969,N_4888);
xor UO_457 (O_457,N_4945,N_4803);
or UO_458 (O_458,N_4963,N_4990);
or UO_459 (O_459,N_4874,N_4842);
nor UO_460 (O_460,N_4853,N_4951);
nand UO_461 (O_461,N_4962,N_4911);
nand UO_462 (O_462,N_4896,N_4920);
nand UO_463 (O_463,N_4953,N_4861);
or UO_464 (O_464,N_4871,N_4996);
nor UO_465 (O_465,N_4901,N_4926);
nor UO_466 (O_466,N_4944,N_4930);
nor UO_467 (O_467,N_4833,N_4856);
nand UO_468 (O_468,N_4852,N_4929);
or UO_469 (O_469,N_4912,N_4980);
or UO_470 (O_470,N_4999,N_4854);
xnor UO_471 (O_471,N_4904,N_4918);
or UO_472 (O_472,N_4829,N_4869);
nor UO_473 (O_473,N_4803,N_4955);
nand UO_474 (O_474,N_4942,N_4881);
and UO_475 (O_475,N_4832,N_4980);
nand UO_476 (O_476,N_4962,N_4978);
or UO_477 (O_477,N_4984,N_4905);
nand UO_478 (O_478,N_4809,N_4829);
nand UO_479 (O_479,N_4944,N_4946);
nand UO_480 (O_480,N_4919,N_4870);
and UO_481 (O_481,N_4853,N_4945);
nand UO_482 (O_482,N_4801,N_4881);
nand UO_483 (O_483,N_4855,N_4839);
and UO_484 (O_484,N_4886,N_4900);
and UO_485 (O_485,N_4980,N_4816);
nand UO_486 (O_486,N_4870,N_4873);
nor UO_487 (O_487,N_4905,N_4814);
nor UO_488 (O_488,N_4898,N_4969);
and UO_489 (O_489,N_4947,N_4910);
nand UO_490 (O_490,N_4994,N_4996);
and UO_491 (O_491,N_4948,N_4890);
nand UO_492 (O_492,N_4944,N_4984);
or UO_493 (O_493,N_4865,N_4967);
nor UO_494 (O_494,N_4840,N_4892);
nand UO_495 (O_495,N_4904,N_4843);
nand UO_496 (O_496,N_4863,N_4927);
and UO_497 (O_497,N_4810,N_4838);
nor UO_498 (O_498,N_4861,N_4931);
and UO_499 (O_499,N_4893,N_4928);
nand UO_500 (O_500,N_4849,N_4933);
and UO_501 (O_501,N_4865,N_4819);
nand UO_502 (O_502,N_4898,N_4842);
or UO_503 (O_503,N_4958,N_4827);
and UO_504 (O_504,N_4837,N_4968);
nor UO_505 (O_505,N_4828,N_4808);
or UO_506 (O_506,N_4872,N_4908);
or UO_507 (O_507,N_4822,N_4860);
and UO_508 (O_508,N_4935,N_4962);
nor UO_509 (O_509,N_4987,N_4817);
and UO_510 (O_510,N_4988,N_4953);
or UO_511 (O_511,N_4906,N_4891);
nand UO_512 (O_512,N_4856,N_4804);
or UO_513 (O_513,N_4967,N_4904);
nand UO_514 (O_514,N_4968,N_4883);
nor UO_515 (O_515,N_4950,N_4952);
or UO_516 (O_516,N_4879,N_4865);
nand UO_517 (O_517,N_4859,N_4849);
and UO_518 (O_518,N_4918,N_4832);
nand UO_519 (O_519,N_4885,N_4906);
and UO_520 (O_520,N_4932,N_4855);
xor UO_521 (O_521,N_4802,N_4966);
nand UO_522 (O_522,N_4949,N_4893);
and UO_523 (O_523,N_4814,N_4939);
nor UO_524 (O_524,N_4993,N_4983);
nand UO_525 (O_525,N_4926,N_4832);
and UO_526 (O_526,N_4856,N_4863);
or UO_527 (O_527,N_4901,N_4802);
nand UO_528 (O_528,N_4878,N_4950);
and UO_529 (O_529,N_4914,N_4970);
nor UO_530 (O_530,N_4969,N_4960);
nor UO_531 (O_531,N_4923,N_4896);
nand UO_532 (O_532,N_4905,N_4977);
or UO_533 (O_533,N_4988,N_4965);
nand UO_534 (O_534,N_4806,N_4884);
nand UO_535 (O_535,N_4913,N_4815);
nand UO_536 (O_536,N_4808,N_4850);
and UO_537 (O_537,N_4972,N_4866);
and UO_538 (O_538,N_4863,N_4960);
nor UO_539 (O_539,N_4925,N_4957);
nand UO_540 (O_540,N_4865,N_4988);
nor UO_541 (O_541,N_4984,N_4958);
or UO_542 (O_542,N_4909,N_4929);
nor UO_543 (O_543,N_4925,N_4982);
or UO_544 (O_544,N_4832,N_4820);
nor UO_545 (O_545,N_4894,N_4872);
nor UO_546 (O_546,N_4827,N_4813);
or UO_547 (O_547,N_4941,N_4914);
or UO_548 (O_548,N_4868,N_4987);
nand UO_549 (O_549,N_4980,N_4820);
and UO_550 (O_550,N_4850,N_4941);
or UO_551 (O_551,N_4873,N_4975);
nor UO_552 (O_552,N_4966,N_4903);
or UO_553 (O_553,N_4850,N_4873);
nor UO_554 (O_554,N_4857,N_4874);
nor UO_555 (O_555,N_4995,N_4985);
nand UO_556 (O_556,N_4970,N_4841);
xor UO_557 (O_557,N_4959,N_4951);
nor UO_558 (O_558,N_4816,N_4938);
and UO_559 (O_559,N_4996,N_4957);
or UO_560 (O_560,N_4969,N_4993);
nand UO_561 (O_561,N_4969,N_4923);
or UO_562 (O_562,N_4968,N_4958);
nand UO_563 (O_563,N_4851,N_4888);
nand UO_564 (O_564,N_4971,N_4907);
and UO_565 (O_565,N_4892,N_4900);
nor UO_566 (O_566,N_4966,N_4878);
and UO_567 (O_567,N_4811,N_4867);
and UO_568 (O_568,N_4811,N_4861);
or UO_569 (O_569,N_4978,N_4912);
and UO_570 (O_570,N_4910,N_4937);
nand UO_571 (O_571,N_4999,N_4861);
nor UO_572 (O_572,N_4835,N_4884);
and UO_573 (O_573,N_4817,N_4988);
and UO_574 (O_574,N_4853,N_4974);
nor UO_575 (O_575,N_4950,N_4922);
nor UO_576 (O_576,N_4988,N_4917);
or UO_577 (O_577,N_4983,N_4892);
and UO_578 (O_578,N_4960,N_4921);
nand UO_579 (O_579,N_4939,N_4855);
nand UO_580 (O_580,N_4966,N_4831);
or UO_581 (O_581,N_4902,N_4950);
nand UO_582 (O_582,N_4951,N_4920);
nand UO_583 (O_583,N_4932,N_4977);
xnor UO_584 (O_584,N_4854,N_4814);
and UO_585 (O_585,N_4867,N_4956);
and UO_586 (O_586,N_4900,N_4963);
nor UO_587 (O_587,N_4906,N_4851);
or UO_588 (O_588,N_4816,N_4841);
and UO_589 (O_589,N_4989,N_4970);
nand UO_590 (O_590,N_4914,N_4895);
or UO_591 (O_591,N_4904,N_4982);
and UO_592 (O_592,N_4985,N_4805);
nor UO_593 (O_593,N_4844,N_4896);
or UO_594 (O_594,N_4986,N_4847);
nand UO_595 (O_595,N_4965,N_4829);
nand UO_596 (O_596,N_4970,N_4852);
nor UO_597 (O_597,N_4910,N_4812);
nor UO_598 (O_598,N_4941,N_4841);
or UO_599 (O_599,N_4811,N_4885);
and UO_600 (O_600,N_4818,N_4989);
nor UO_601 (O_601,N_4926,N_4982);
or UO_602 (O_602,N_4985,N_4860);
nand UO_603 (O_603,N_4961,N_4991);
nor UO_604 (O_604,N_4978,N_4965);
nor UO_605 (O_605,N_4988,N_4806);
nor UO_606 (O_606,N_4938,N_4932);
and UO_607 (O_607,N_4929,N_4905);
or UO_608 (O_608,N_4820,N_4948);
or UO_609 (O_609,N_4954,N_4876);
or UO_610 (O_610,N_4813,N_4876);
or UO_611 (O_611,N_4996,N_4934);
or UO_612 (O_612,N_4920,N_4811);
and UO_613 (O_613,N_4934,N_4877);
and UO_614 (O_614,N_4896,N_4911);
and UO_615 (O_615,N_4871,N_4969);
xnor UO_616 (O_616,N_4906,N_4983);
nand UO_617 (O_617,N_4878,N_4999);
xor UO_618 (O_618,N_4962,N_4827);
nor UO_619 (O_619,N_4947,N_4995);
nand UO_620 (O_620,N_4912,N_4845);
and UO_621 (O_621,N_4977,N_4952);
or UO_622 (O_622,N_4962,N_4940);
or UO_623 (O_623,N_4877,N_4816);
nor UO_624 (O_624,N_4995,N_4963);
or UO_625 (O_625,N_4805,N_4801);
nor UO_626 (O_626,N_4891,N_4837);
nand UO_627 (O_627,N_4836,N_4877);
or UO_628 (O_628,N_4857,N_4998);
and UO_629 (O_629,N_4879,N_4917);
and UO_630 (O_630,N_4819,N_4985);
nand UO_631 (O_631,N_4909,N_4950);
or UO_632 (O_632,N_4801,N_4869);
and UO_633 (O_633,N_4814,N_4862);
nor UO_634 (O_634,N_4880,N_4806);
nor UO_635 (O_635,N_4986,N_4878);
and UO_636 (O_636,N_4929,N_4934);
nand UO_637 (O_637,N_4887,N_4869);
and UO_638 (O_638,N_4960,N_4898);
nand UO_639 (O_639,N_4900,N_4802);
or UO_640 (O_640,N_4989,N_4958);
nand UO_641 (O_641,N_4802,N_4975);
nand UO_642 (O_642,N_4990,N_4910);
and UO_643 (O_643,N_4922,N_4836);
nand UO_644 (O_644,N_4813,N_4888);
nor UO_645 (O_645,N_4830,N_4895);
or UO_646 (O_646,N_4967,N_4929);
or UO_647 (O_647,N_4896,N_4888);
xnor UO_648 (O_648,N_4904,N_4935);
or UO_649 (O_649,N_4930,N_4865);
and UO_650 (O_650,N_4945,N_4841);
and UO_651 (O_651,N_4904,N_4964);
nand UO_652 (O_652,N_4861,N_4949);
nand UO_653 (O_653,N_4817,N_4914);
nand UO_654 (O_654,N_4860,N_4817);
and UO_655 (O_655,N_4829,N_4864);
or UO_656 (O_656,N_4972,N_4896);
and UO_657 (O_657,N_4989,N_4946);
or UO_658 (O_658,N_4984,N_4945);
nor UO_659 (O_659,N_4806,N_4922);
and UO_660 (O_660,N_4868,N_4927);
nor UO_661 (O_661,N_4946,N_4894);
or UO_662 (O_662,N_4959,N_4837);
nor UO_663 (O_663,N_4933,N_4864);
or UO_664 (O_664,N_4914,N_4939);
nor UO_665 (O_665,N_4950,N_4900);
or UO_666 (O_666,N_4898,N_4852);
and UO_667 (O_667,N_4949,N_4885);
nand UO_668 (O_668,N_4841,N_4865);
or UO_669 (O_669,N_4846,N_4864);
nand UO_670 (O_670,N_4832,N_4894);
and UO_671 (O_671,N_4920,N_4812);
nand UO_672 (O_672,N_4948,N_4871);
or UO_673 (O_673,N_4960,N_4899);
nor UO_674 (O_674,N_4823,N_4897);
nor UO_675 (O_675,N_4836,N_4837);
nand UO_676 (O_676,N_4897,N_4934);
and UO_677 (O_677,N_4957,N_4810);
nor UO_678 (O_678,N_4863,N_4941);
xor UO_679 (O_679,N_4837,N_4817);
or UO_680 (O_680,N_4839,N_4898);
and UO_681 (O_681,N_4933,N_4898);
and UO_682 (O_682,N_4849,N_4843);
xor UO_683 (O_683,N_4873,N_4942);
nand UO_684 (O_684,N_4955,N_4918);
nand UO_685 (O_685,N_4826,N_4958);
or UO_686 (O_686,N_4880,N_4981);
nor UO_687 (O_687,N_4993,N_4881);
and UO_688 (O_688,N_4821,N_4856);
nand UO_689 (O_689,N_4884,N_4923);
or UO_690 (O_690,N_4925,N_4967);
nand UO_691 (O_691,N_4921,N_4855);
nand UO_692 (O_692,N_4880,N_4931);
or UO_693 (O_693,N_4991,N_4871);
nor UO_694 (O_694,N_4933,N_4893);
or UO_695 (O_695,N_4838,N_4920);
or UO_696 (O_696,N_4973,N_4975);
xor UO_697 (O_697,N_4910,N_4887);
nor UO_698 (O_698,N_4980,N_4818);
nor UO_699 (O_699,N_4861,N_4919);
nor UO_700 (O_700,N_4855,N_4867);
nand UO_701 (O_701,N_4850,N_4940);
nand UO_702 (O_702,N_4883,N_4898);
nand UO_703 (O_703,N_4885,N_4993);
or UO_704 (O_704,N_4936,N_4857);
nor UO_705 (O_705,N_4965,N_4851);
nand UO_706 (O_706,N_4946,N_4974);
or UO_707 (O_707,N_4936,N_4897);
nor UO_708 (O_708,N_4930,N_4955);
and UO_709 (O_709,N_4963,N_4971);
nor UO_710 (O_710,N_4990,N_4916);
nand UO_711 (O_711,N_4853,N_4969);
nor UO_712 (O_712,N_4863,N_4872);
or UO_713 (O_713,N_4904,N_4850);
or UO_714 (O_714,N_4887,N_4825);
and UO_715 (O_715,N_4868,N_4993);
and UO_716 (O_716,N_4958,N_4873);
or UO_717 (O_717,N_4812,N_4973);
nor UO_718 (O_718,N_4933,N_4837);
nor UO_719 (O_719,N_4885,N_4806);
and UO_720 (O_720,N_4927,N_4925);
nand UO_721 (O_721,N_4959,N_4940);
nand UO_722 (O_722,N_4999,N_4912);
or UO_723 (O_723,N_4962,N_4889);
nand UO_724 (O_724,N_4973,N_4949);
xnor UO_725 (O_725,N_4854,N_4969);
and UO_726 (O_726,N_4831,N_4919);
or UO_727 (O_727,N_4938,N_4964);
nand UO_728 (O_728,N_4921,N_4853);
and UO_729 (O_729,N_4964,N_4810);
and UO_730 (O_730,N_4873,N_4821);
and UO_731 (O_731,N_4824,N_4941);
nand UO_732 (O_732,N_4969,N_4918);
nor UO_733 (O_733,N_4968,N_4928);
or UO_734 (O_734,N_4910,N_4941);
nand UO_735 (O_735,N_4855,N_4997);
and UO_736 (O_736,N_4876,N_4870);
and UO_737 (O_737,N_4815,N_4862);
or UO_738 (O_738,N_4977,N_4981);
or UO_739 (O_739,N_4900,N_4974);
or UO_740 (O_740,N_4992,N_4868);
and UO_741 (O_741,N_4938,N_4995);
and UO_742 (O_742,N_4960,N_4827);
nand UO_743 (O_743,N_4867,N_4854);
and UO_744 (O_744,N_4897,N_4845);
xor UO_745 (O_745,N_4927,N_4801);
and UO_746 (O_746,N_4946,N_4986);
nor UO_747 (O_747,N_4902,N_4925);
nand UO_748 (O_748,N_4812,N_4838);
or UO_749 (O_749,N_4948,N_4994);
and UO_750 (O_750,N_4814,N_4954);
nand UO_751 (O_751,N_4808,N_4879);
and UO_752 (O_752,N_4994,N_4819);
or UO_753 (O_753,N_4939,N_4866);
or UO_754 (O_754,N_4865,N_4875);
nor UO_755 (O_755,N_4942,N_4831);
nand UO_756 (O_756,N_4883,N_4916);
xor UO_757 (O_757,N_4855,N_4987);
nand UO_758 (O_758,N_4821,N_4823);
nor UO_759 (O_759,N_4862,N_4800);
nand UO_760 (O_760,N_4889,N_4837);
nand UO_761 (O_761,N_4973,N_4877);
nor UO_762 (O_762,N_4820,N_4977);
or UO_763 (O_763,N_4845,N_4815);
nand UO_764 (O_764,N_4959,N_4886);
xnor UO_765 (O_765,N_4833,N_4881);
and UO_766 (O_766,N_4839,N_4997);
or UO_767 (O_767,N_4957,N_4818);
or UO_768 (O_768,N_4991,N_4923);
or UO_769 (O_769,N_4886,N_4978);
nor UO_770 (O_770,N_4891,N_4809);
nand UO_771 (O_771,N_4879,N_4810);
and UO_772 (O_772,N_4978,N_4934);
and UO_773 (O_773,N_4967,N_4935);
nor UO_774 (O_774,N_4883,N_4850);
and UO_775 (O_775,N_4909,N_4972);
or UO_776 (O_776,N_4810,N_4999);
and UO_777 (O_777,N_4866,N_4902);
nor UO_778 (O_778,N_4850,N_4807);
and UO_779 (O_779,N_4921,N_4884);
nor UO_780 (O_780,N_4945,N_4852);
nand UO_781 (O_781,N_4813,N_4803);
nor UO_782 (O_782,N_4896,N_4884);
and UO_783 (O_783,N_4825,N_4817);
nand UO_784 (O_784,N_4924,N_4921);
and UO_785 (O_785,N_4826,N_4927);
nand UO_786 (O_786,N_4909,N_4831);
nor UO_787 (O_787,N_4875,N_4882);
nor UO_788 (O_788,N_4935,N_4805);
nand UO_789 (O_789,N_4834,N_4953);
nand UO_790 (O_790,N_4903,N_4820);
and UO_791 (O_791,N_4808,N_4888);
nor UO_792 (O_792,N_4937,N_4964);
or UO_793 (O_793,N_4968,N_4842);
nand UO_794 (O_794,N_4869,N_4860);
or UO_795 (O_795,N_4835,N_4911);
and UO_796 (O_796,N_4921,N_4979);
or UO_797 (O_797,N_4986,N_4960);
and UO_798 (O_798,N_4935,N_4898);
or UO_799 (O_799,N_4996,N_4870);
or UO_800 (O_800,N_4903,N_4929);
or UO_801 (O_801,N_4925,N_4849);
and UO_802 (O_802,N_4864,N_4831);
or UO_803 (O_803,N_4818,N_4930);
nor UO_804 (O_804,N_4900,N_4990);
nor UO_805 (O_805,N_4904,N_4839);
and UO_806 (O_806,N_4876,N_4832);
nand UO_807 (O_807,N_4918,N_4806);
nor UO_808 (O_808,N_4953,N_4814);
nor UO_809 (O_809,N_4827,N_4916);
nand UO_810 (O_810,N_4818,N_4928);
and UO_811 (O_811,N_4955,N_4800);
nor UO_812 (O_812,N_4944,N_4989);
nand UO_813 (O_813,N_4808,N_4917);
nand UO_814 (O_814,N_4875,N_4994);
and UO_815 (O_815,N_4873,N_4982);
and UO_816 (O_816,N_4806,N_4850);
and UO_817 (O_817,N_4866,N_4864);
nor UO_818 (O_818,N_4894,N_4968);
nor UO_819 (O_819,N_4971,N_4852);
and UO_820 (O_820,N_4862,N_4974);
nand UO_821 (O_821,N_4854,N_4831);
or UO_822 (O_822,N_4897,N_4928);
and UO_823 (O_823,N_4944,N_4822);
nor UO_824 (O_824,N_4943,N_4810);
nor UO_825 (O_825,N_4923,N_4815);
nand UO_826 (O_826,N_4942,N_4815);
nand UO_827 (O_827,N_4908,N_4969);
or UO_828 (O_828,N_4954,N_4842);
and UO_829 (O_829,N_4972,N_4938);
nand UO_830 (O_830,N_4989,N_4816);
or UO_831 (O_831,N_4934,N_4922);
and UO_832 (O_832,N_4913,N_4851);
nand UO_833 (O_833,N_4807,N_4957);
nand UO_834 (O_834,N_4841,N_4955);
nand UO_835 (O_835,N_4990,N_4936);
and UO_836 (O_836,N_4872,N_4975);
and UO_837 (O_837,N_4983,N_4972);
nand UO_838 (O_838,N_4984,N_4805);
nor UO_839 (O_839,N_4980,N_4896);
and UO_840 (O_840,N_4854,N_4971);
nor UO_841 (O_841,N_4801,N_4903);
or UO_842 (O_842,N_4982,N_4843);
nand UO_843 (O_843,N_4872,N_4861);
or UO_844 (O_844,N_4887,N_4983);
and UO_845 (O_845,N_4819,N_4975);
and UO_846 (O_846,N_4953,N_4828);
xor UO_847 (O_847,N_4949,N_4938);
or UO_848 (O_848,N_4937,N_4866);
nor UO_849 (O_849,N_4993,N_4836);
nor UO_850 (O_850,N_4955,N_4834);
and UO_851 (O_851,N_4967,N_4907);
and UO_852 (O_852,N_4941,N_4950);
nand UO_853 (O_853,N_4984,N_4859);
or UO_854 (O_854,N_4933,N_4886);
nand UO_855 (O_855,N_4880,N_4974);
and UO_856 (O_856,N_4866,N_4867);
or UO_857 (O_857,N_4976,N_4889);
and UO_858 (O_858,N_4820,N_4847);
and UO_859 (O_859,N_4998,N_4804);
and UO_860 (O_860,N_4988,N_4915);
and UO_861 (O_861,N_4926,N_4967);
or UO_862 (O_862,N_4925,N_4977);
and UO_863 (O_863,N_4921,N_4838);
and UO_864 (O_864,N_4970,N_4979);
nand UO_865 (O_865,N_4816,N_4918);
or UO_866 (O_866,N_4863,N_4985);
or UO_867 (O_867,N_4812,N_4901);
and UO_868 (O_868,N_4829,N_4934);
and UO_869 (O_869,N_4967,N_4946);
nand UO_870 (O_870,N_4981,N_4815);
nand UO_871 (O_871,N_4873,N_4990);
and UO_872 (O_872,N_4967,N_4961);
or UO_873 (O_873,N_4938,N_4984);
nand UO_874 (O_874,N_4965,N_4920);
nand UO_875 (O_875,N_4979,N_4951);
xnor UO_876 (O_876,N_4827,N_4957);
or UO_877 (O_877,N_4841,N_4852);
nand UO_878 (O_878,N_4889,N_4981);
nor UO_879 (O_879,N_4870,N_4910);
nand UO_880 (O_880,N_4983,N_4985);
and UO_881 (O_881,N_4888,N_4819);
or UO_882 (O_882,N_4852,N_4827);
or UO_883 (O_883,N_4852,N_4869);
nor UO_884 (O_884,N_4876,N_4972);
and UO_885 (O_885,N_4896,N_4857);
and UO_886 (O_886,N_4982,N_4848);
nor UO_887 (O_887,N_4928,N_4886);
nand UO_888 (O_888,N_4968,N_4817);
and UO_889 (O_889,N_4919,N_4964);
nor UO_890 (O_890,N_4840,N_4829);
nand UO_891 (O_891,N_4802,N_4880);
and UO_892 (O_892,N_4831,N_4958);
nor UO_893 (O_893,N_4821,N_4859);
nand UO_894 (O_894,N_4852,N_4983);
and UO_895 (O_895,N_4834,N_4918);
nand UO_896 (O_896,N_4953,N_4929);
or UO_897 (O_897,N_4803,N_4872);
nor UO_898 (O_898,N_4925,N_4815);
xor UO_899 (O_899,N_4958,N_4949);
or UO_900 (O_900,N_4880,N_4874);
nor UO_901 (O_901,N_4898,N_4872);
and UO_902 (O_902,N_4900,N_4924);
nand UO_903 (O_903,N_4801,N_4901);
nor UO_904 (O_904,N_4983,N_4865);
and UO_905 (O_905,N_4887,N_4975);
xnor UO_906 (O_906,N_4843,N_4920);
nand UO_907 (O_907,N_4913,N_4936);
nand UO_908 (O_908,N_4886,N_4977);
and UO_909 (O_909,N_4861,N_4877);
xor UO_910 (O_910,N_4836,N_4985);
and UO_911 (O_911,N_4988,N_4994);
xor UO_912 (O_912,N_4891,N_4869);
nor UO_913 (O_913,N_4998,N_4847);
or UO_914 (O_914,N_4856,N_4928);
nor UO_915 (O_915,N_4968,N_4839);
nor UO_916 (O_916,N_4808,N_4959);
or UO_917 (O_917,N_4911,N_4865);
nor UO_918 (O_918,N_4915,N_4960);
and UO_919 (O_919,N_4812,N_4857);
nor UO_920 (O_920,N_4823,N_4847);
or UO_921 (O_921,N_4986,N_4934);
nor UO_922 (O_922,N_4897,N_4921);
or UO_923 (O_923,N_4842,N_4864);
and UO_924 (O_924,N_4911,N_4944);
and UO_925 (O_925,N_4831,N_4802);
and UO_926 (O_926,N_4979,N_4914);
or UO_927 (O_927,N_4980,N_4851);
and UO_928 (O_928,N_4888,N_4828);
or UO_929 (O_929,N_4900,N_4857);
and UO_930 (O_930,N_4994,N_4916);
and UO_931 (O_931,N_4995,N_4892);
and UO_932 (O_932,N_4832,N_4898);
nor UO_933 (O_933,N_4815,N_4973);
or UO_934 (O_934,N_4996,N_4863);
or UO_935 (O_935,N_4947,N_4828);
nor UO_936 (O_936,N_4999,N_4941);
xor UO_937 (O_937,N_4821,N_4967);
nor UO_938 (O_938,N_4851,N_4981);
and UO_939 (O_939,N_4876,N_4875);
and UO_940 (O_940,N_4968,N_4980);
nor UO_941 (O_941,N_4936,N_4843);
and UO_942 (O_942,N_4801,N_4854);
and UO_943 (O_943,N_4917,N_4951);
and UO_944 (O_944,N_4844,N_4985);
nand UO_945 (O_945,N_4989,N_4982);
nand UO_946 (O_946,N_4977,N_4960);
or UO_947 (O_947,N_4914,N_4833);
or UO_948 (O_948,N_4874,N_4946);
nand UO_949 (O_949,N_4875,N_4866);
nand UO_950 (O_950,N_4813,N_4843);
nand UO_951 (O_951,N_4814,N_4821);
nand UO_952 (O_952,N_4967,N_4808);
or UO_953 (O_953,N_4964,N_4838);
nor UO_954 (O_954,N_4934,N_4828);
or UO_955 (O_955,N_4947,N_4906);
xnor UO_956 (O_956,N_4829,N_4810);
xnor UO_957 (O_957,N_4929,N_4861);
xor UO_958 (O_958,N_4877,N_4956);
xnor UO_959 (O_959,N_4932,N_4900);
nand UO_960 (O_960,N_4861,N_4913);
nand UO_961 (O_961,N_4897,N_4962);
or UO_962 (O_962,N_4871,N_4980);
nor UO_963 (O_963,N_4966,N_4996);
or UO_964 (O_964,N_4918,N_4869);
or UO_965 (O_965,N_4990,N_4961);
nor UO_966 (O_966,N_4823,N_4854);
and UO_967 (O_967,N_4827,N_4997);
nor UO_968 (O_968,N_4938,N_4872);
nor UO_969 (O_969,N_4833,N_4845);
or UO_970 (O_970,N_4978,N_4918);
nand UO_971 (O_971,N_4843,N_4884);
nor UO_972 (O_972,N_4931,N_4956);
nor UO_973 (O_973,N_4972,N_4904);
xor UO_974 (O_974,N_4906,N_4970);
or UO_975 (O_975,N_4951,N_4837);
or UO_976 (O_976,N_4955,N_4914);
and UO_977 (O_977,N_4920,N_4930);
and UO_978 (O_978,N_4975,N_4841);
xnor UO_979 (O_979,N_4917,N_4995);
nand UO_980 (O_980,N_4934,N_4927);
nand UO_981 (O_981,N_4928,N_4829);
and UO_982 (O_982,N_4964,N_4849);
or UO_983 (O_983,N_4919,N_4999);
nor UO_984 (O_984,N_4983,N_4815);
nor UO_985 (O_985,N_4930,N_4848);
xor UO_986 (O_986,N_4928,N_4956);
or UO_987 (O_987,N_4882,N_4852);
nor UO_988 (O_988,N_4842,N_4840);
nor UO_989 (O_989,N_4982,N_4938);
nor UO_990 (O_990,N_4914,N_4860);
nor UO_991 (O_991,N_4817,N_4867);
and UO_992 (O_992,N_4912,N_4939);
nand UO_993 (O_993,N_4832,N_4861);
nor UO_994 (O_994,N_4858,N_4971);
nor UO_995 (O_995,N_4819,N_4955);
nor UO_996 (O_996,N_4937,N_4821);
or UO_997 (O_997,N_4818,N_4969);
or UO_998 (O_998,N_4845,N_4871);
or UO_999 (O_999,N_4912,N_4838);
endmodule