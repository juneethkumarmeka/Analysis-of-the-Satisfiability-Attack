module basic_2000_20000_2500_5_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
or U0 (N_0,In_1802,In_218);
nor U1 (N_1,In_183,In_671);
xnor U2 (N_2,In_543,In_1376);
or U3 (N_3,In_1873,In_231);
xnor U4 (N_4,In_497,In_1514);
and U5 (N_5,In_392,In_48);
and U6 (N_6,In_1721,In_357);
and U7 (N_7,In_840,In_1250);
or U8 (N_8,In_522,In_1320);
xnor U9 (N_9,In_1226,In_35);
and U10 (N_10,In_1961,In_534);
or U11 (N_11,In_7,In_1241);
nor U12 (N_12,In_918,In_526);
xnor U13 (N_13,In_1187,In_774);
xor U14 (N_14,In_1259,In_894);
or U15 (N_15,In_483,In_1644);
nand U16 (N_16,In_1550,In_1010);
nor U17 (N_17,In_253,In_1963);
nor U18 (N_18,In_920,In_1493);
or U19 (N_19,In_1256,In_427);
xor U20 (N_20,In_551,In_226);
nand U21 (N_21,In_595,In_1);
and U22 (N_22,In_244,In_393);
xor U23 (N_23,In_1385,In_1069);
xnor U24 (N_24,In_1617,In_454);
nand U25 (N_25,In_1946,In_475);
nor U26 (N_26,In_558,In_1281);
xor U27 (N_27,In_1660,In_795);
nand U28 (N_28,In_1889,In_866);
and U29 (N_29,In_438,In_1654);
xnor U30 (N_30,In_836,In_1835);
and U31 (N_31,In_981,In_1176);
nor U32 (N_32,In_892,In_1999);
nand U33 (N_33,In_1569,In_684);
xor U34 (N_34,In_1439,In_1536);
nand U35 (N_35,In_584,In_1397);
nor U36 (N_36,In_1322,In_954);
nor U37 (N_37,In_246,In_1708);
and U38 (N_38,In_749,In_1403);
nand U39 (N_39,In_1503,In_1723);
xnor U40 (N_40,In_1347,In_1152);
xor U41 (N_41,In_1809,In_1150);
or U42 (N_42,In_1497,In_1715);
nand U43 (N_43,In_528,In_1477);
or U44 (N_44,In_1876,In_1843);
nand U45 (N_45,In_776,In_1167);
xor U46 (N_46,In_1217,In_536);
nor U47 (N_47,In_345,In_816);
nand U48 (N_48,In_582,In_623);
nand U49 (N_49,In_1437,In_1292);
xnor U50 (N_50,In_1460,In_1599);
nand U51 (N_51,In_1053,In_425);
nor U52 (N_52,In_624,In_770);
and U53 (N_53,In_407,In_1340);
nor U54 (N_54,In_539,In_1712);
nor U55 (N_55,In_247,In_885);
and U56 (N_56,In_1329,In_1034);
and U57 (N_57,In_440,In_1185);
and U58 (N_58,In_727,In_107);
or U59 (N_59,In_472,In_1379);
nand U60 (N_60,In_945,In_384);
nand U61 (N_61,In_609,In_1778);
nor U62 (N_62,In_1291,In_887);
or U63 (N_63,In_1529,In_1666);
nor U64 (N_64,In_1746,In_4);
and U65 (N_65,In_1832,In_293);
xor U66 (N_66,In_1979,In_1282);
and U67 (N_67,In_697,In_903);
xnor U68 (N_68,In_1002,In_900);
or U69 (N_69,In_1810,In_78);
xnor U70 (N_70,In_1841,In_1021);
xor U71 (N_71,In_882,In_1283);
xor U72 (N_72,In_1290,In_287);
nand U73 (N_73,In_768,In_1014);
and U74 (N_74,In_318,In_1751);
and U75 (N_75,In_1001,In_1211);
nand U76 (N_76,In_1044,In_1970);
nand U77 (N_77,In_1787,In_1694);
and U78 (N_78,In_1052,In_660);
nand U79 (N_79,In_1412,In_1507);
nand U80 (N_80,In_1155,In_908);
xor U81 (N_81,In_1370,In_890);
nor U82 (N_82,In_1271,In_680);
nand U83 (N_83,In_1727,In_154);
xor U84 (N_84,In_370,In_1177);
xnor U85 (N_85,In_1381,In_1188);
nand U86 (N_86,In_1878,In_23);
or U87 (N_87,In_1011,In_49);
and U88 (N_88,In_321,In_1824);
and U89 (N_89,In_1844,In_650);
and U90 (N_90,In_983,In_135);
nand U91 (N_91,In_262,In_1196);
and U92 (N_92,In_388,In_978);
nand U93 (N_93,In_1730,In_1990);
xnor U94 (N_94,In_1888,In_1095);
nor U95 (N_95,In_99,In_1936);
nand U96 (N_96,In_1697,In_269);
nand U97 (N_97,In_674,In_1985);
nand U98 (N_98,In_1111,In_9);
nand U99 (N_99,In_656,In_872);
xnor U100 (N_100,In_1974,In_106);
or U101 (N_101,In_670,In_310);
nor U102 (N_102,In_640,In_1962);
or U103 (N_103,In_811,In_1781);
nor U104 (N_104,In_1992,In_187);
or U105 (N_105,In_306,In_819);
or U106 (N_106,In_40,In_859);
or U107 (N_107,In_1890,In_631);
and U108 (N_108,In_1797,In_1079);
nor U109 (N_109,In_494,In_1452);
xor U110 (N_110,In_1704,In_1958);
nand U111 (N_111,In_397,In_1473);
and U112 (N_112,In_951,In_672);
or U113 (N_113,In_1931,In_997);
nor U114 (N_114,In_330,In_821);
or U115 (N_115,In_1816,In_202);
or U116 (N_116,In_1659,In_1035);
xor U117 (N_117,In_337,In_898);
nand U118 (N_118,In_1462,In_1692);
nand U119 (N_119,In_1297,In_1233);
nor U120 (N_120,In_1264,In_1565);
xor U121 (N_121,In_1975,In_747);
nor U122 (N_122,In_1072,In_1578);
or U123 (N_123,In_915,In_433);
nand U124 (N_124,In_1251,In_1582);
xor U125 (N_125,In_220,In_174);
and U126 (N_126,In_1857,In_1771);
nand U127 (N_127,In_1212,In_1877);
nor U128 (N_128,In_962,In_815);
nand U129 (N_129,In_1823,In_46);
xor U130 (N_130,In_1016,In_1828);
and U131 (N_131,In_316,In_530);
xor U132 (N_132,In_1634,In_132);
nor U133 (N_133,In_517,In_1764);
or U134 (N_134,In_1899,In_143);
and U135 (N_135,In_1068,In_1935);
and U136 (N_136,In_1033,In_1592);
nand U137 (N_137,In_878,In_781);
and U138 (N_138,In_468,In_1589);
and U139 (N_139,In_987,In_1918);
nand U140 (N_140,In_649,In_1351);
and U141 (N_141,In_426,In_1517);
nand U142 (N_142,In_444,In_1467);
nand U143 (N_143,In_1213,In_998);
and U144 (N_144,In_385,In_185);
nand U145 (N_145,In_557,In_1800);
or U146 (N_146,In_709,In_1720);
or U147 (N_147,In_1729,In_1137);
and U148 (N_148,In_1235,In_1651);
nand U149 (N_149,In_214,In_1556);
or U150 (N_150,In_1768,In_615);
nor U151 (N_151,In_1490,In_1971);
nor U152 (N_152,In_495,In_1997);
nand U153 (N_153,In_1732,In_1986);
xor U154 (N_154,In_1570,In_549);
or U155 (N_155,In_1656,In_1829);
nand U156 (N_156,In_939,In_493);
nand U157 (N_157,In_323,In_1948);
and U158 (N_158,In_1885,In_1554);
xor U159 (N_159,In_950,In_44);
nand U160 (N_160,In_668,In_326);
nor U161 (N_161,In_798,In_1615);
or U162 (N_162,In_34,In_996);
nor U163 (N_163,In_216,In_1312);
or U164 (N_164,In_91,In_1195);
and U165 (N_165,In_1458,In_1363);
or U166 (N_166,In_1197,In_568);
xor U167 (N_167,In_1788,In_1350);
and U168 (N_168,In_1025,In_1309);
and U169 (N_169,In_1173,In_698);
nor U170 (N_170,In_554,In_773);
and U171 (N_171,In_1400,In_1042);
or U172 (N_172,In_1293,In_1475);
and U173 (N_173,In_1194,In_739);
nor U174 (N_174,In_1145,In_955);
or U175 (N_175,In_735,In_1080);
and U176 (N_176,In_1396,In_1041);
and U177 (N_177,In_1066,In_1261);
and U178 (N_178,In_1134,In_36);
nor U179 (N_179,In_579,In_1834);
nand U180 (N_180,In_450,In_729);
nor U181 (N_181,In_1995,In_161);
xnor U182 (N_182,In_946,In_1806);
or U183 (N_183,In_1776,In_1031);
and U184 (N_184,In_547,In_502);
nand U185 (N_185,In_402,In_1605);
nand U186 (N_186,In_1366,In_827);
nand U187 (N_187,In_1013,In_934);
and U188 (N_188,In_678,In_380);
nand U189 (N_189,In_1190,In_245);
nor U190 (N_190,In_1484,In_249);
or U191 (N_191,In_1557,In_1853);
or U192 (N_192,In_1608,In_1837);
or U193 (N_193,In_1562,In_1210);
nor U194 (N_194,In_291,In_1638);
nand U195 (N_195,In_1100,In_446);
or U196 (N_196,In_375,In_1920);
or U197 (N_197,In_870,In_1623);
nor U198 (N_198,In_1548,In_1149);
nand U199 (N_199,In_307,In_234);
or U200 (N_200,In_1722,In_914);
or U201 (N_201,In_369,In_1005);
nand U202 (N_202,In_700,In_474);
or U203 (N_203,In_1595,In_356);
and U204 (N_204,In_1774,In_263);
and U205 (N_205,In_1371,In_1154);
and U206 (N_206,In_1133,In_47);
nor U207 (N_207,In_1945,In_991);
or U208 (N_208,In_1189,In_599);
nand U209 (N_209,In_209,In_689);
xor U210 (N_210,In_157,In_527);
or U211 (N_211,In_1022,In_794);
or U212 (N_212,In_875,In_1941);
and U213 (N_213,In_1372,In_276);
xnor U214 (N_214,In_42,In_90);
and U215 (N_215,In_655,In_1140);
nand U216 (N_216,In_1906,In_626);
xnor U217 (N_217,In_1308,In_1461);
and U218 (N_218,In_274,In_862);
nand U219 (N_219,In_273,In_1951);
and U220 (N_220,In_1472,In_1319);
nand U221 (N_221,In_1652,In_664);
nor U222 (N_222,In_1489,In_1984);
or U223 (N_223,In_1126,In_886);
and U224 (N_224,In_208,In_740);
xnor U225 (N_225,In_1242,In_240);
xor U226 (N_226,In_1561,In_491);
nor U227 (N_227,In_1328,In_513);
or U228 (N_228,In_65,In_685);
or U229 (N_229,In_583,In_1808);
nor U230 (N_230,In_464,In_966);
or U231 (N_231,In_1485,In_930);
and U232 (N_232,In_1246,In_1169);
nand U233 (N_233,In_1639,In_531);
nor U234 (N_234,In_101,In_591);
or U235 (N_235,In_1425,In_1738);
nand U236 (N_236,In_511,In_328);
nor U237 (N_237,In_1944,In_1040);
or U238 (N_238,In_1682,In_1258);
xor U239 (N_239,In_172,In_498);
and U240 (N_240,In_1048,In_1421);
nand U241 (N_241,In_1663,In_471);
nand U242 (N_242,In_149,In_1676);
or U243 (N_243,In_1273,In_302);
nand U244 (N_244,In_1735,In_1620);
or U245 (N_245,In_1520,In_559);
or U246 (N_246,In_1224,In_145);
and U247 (N_247,In_566,In_96);
and U248 (N_248,In_1600,In_1408);
and U249 (N_249,In_902,In_264);
xnor U250 (N_250,In_1168,In_546);
nand U251 (N_251,In_753,In_818);
or U252 (N_252,In_1938,In_1129);
or U253 (N_253,In_417,In_1051);
nand U254 (N_254,In_1494,In_45);
nand U255 (N_255,In_56,In_720);
xor U256 (N_256,In_1348,In_21);
and U257 (N_257,In_1586,In_1094);
and U258 (N_258,In_270,In_2);
xor U259 (N_259,In_723,In_959);
and U260 (N_260,In_125,In_1665);
or U261 (N_261,In_627,In_288);
nand U262 (N_262,In_1967,In_1953);
and U263 (N_263,In_435,In_1216);
or U264 (N_264,In_294,In_386);
and U265 (N_265,In_704,In_1192);
xnor U266 (N_266,In_1792,In_1921);
nor U267 (N_267,In_1934,In_424);
nor U268 (N_268,In_97,In_779);
nor U269 (N_269,In_404,In_578);
and U270 (N_270,In_1588,In_57);
and U271 (N_271,In_1672,In_507);
and U272 (N_272,In_1894,In_594);
xnor U273 (N_273,In_204,In_1277);
nor U274 (N_274,In_104,In_1763);
nor U275 (N_275,In_289,In_113);
xnor U276 (N_276,In_1220,In_876);
and U277 (N_277,In_140,In_1922);
nand U278 (N_278,In_77,In_422);
nor U279 (N_279,In_254,In_279);
xnor U280 (N_280,In_341,In_159);
nor U281 (N_281,In_1471,In_917);
and U282 (N_282,In_1706,In_1686);
nand U283 (N_283,In_1247,In_391);
and U284 (N_284,In_995,In_967);
nand U285 (N_285,In_1534,In_1649);
and U286 (N_286,In_1757,In_1081);
nor U287 (N_287,In_1927,In_1773);
xor U288 (N_288,In_1869,In_1530);
nor U289 (N_289,In_848,In_1897);
nor U290 (N_290,In_86,In_1904);
nor U291 (N_291,In_1333,In_1510);
nor U292 (N_292,In_1142,In_1765);
nor U293 (N_293,In_1380,In_1766);
xor U294 (N_294,In_1455,In_1017);
nand U295 (N_295,In_1318,In_437);
or U296 (N_296,In_1463,In_223);
and U297 (N_297,In_673,In_1270);
or U298 (N_298,In_856,In_1544);
or U299 (N_299,In_1110,In_1614);
or U300 (N_300,In_1257,In_351);
nand U301 (N_301,In_1560,In_659);
nand U302 (N_302,In_1861,In_1337);
nand U303 (N_303,In_575,In_1761);
and U304 (N_304,In_1917,In_545);
or U305 (N_305,In_1862,In_969);
nand U306 (N_306,In_478,In_889);
or U307 (N_307,In_782,In_1770);
xor U308 (N_308,In_1083,In_1830);
nand U309 (N_309,In_1276,In_1976);
or U310 (N_310,In_362,In_1880);
or U311 (N_311,In_948,In_1891);
nand U312 (N_312,In_508,In_1524);
nand U313 (N_313,In_1601,In_347);
and U314 (N_314,In_1981,In_1346);
and U315 (N_315,In_1505,In_195);
nand U316 (N_316,In_473,In_1249);
xnor U317 (N_317,In_1143,In_620);
nand U318 (N_318,In_1977,In_8);
nor U319 (N_319,In_428,In_320);
nand U320 (N_320,In_1334,In_926);
nand U321 (N_321,In_1581,In_58);
and U322 (N_322,In_610,In_1252);
nor U323 (N_323,In_1914,In_1688);
or U324 (N_324,In_1236,In_592);
nand U325 (N_325,In_1690,In_1858);
nand U326 (N_326,In_761,In_284);
nor U327 (N_327,In_30,In_941);
nor U328 (N_328,In_1637,In_1508);
or U329 (N_329,In_1699,In_845);
or U330 (N_330,In_1789,In_120);
and U331 (N_331,In_577,In_1313);
or U332 (N_332,In_802,In_873);
and U333 (N_333,In_1426,In_1643);
xnor U334 (N_334,In_363,In_1952);
xor U335 (N_335,In_420,In_841);
xor U336 (N_336,In_1267,In_83);
nor U337 (N_337,In_448,In_1105);
nand U338 (N_338,In_1470,In_963);
and U339 (N_339,In_238,In_309);
nand U340 (N_340,In_124,In_1390);
xnor U341 (N_341,In_1838,In_1209);
xor U342 (N_342,In_193,In_1059);
xnor U343 (N_343,In_1499,In_1479);
or U344 (N_344,In_186,In_797);
xor U345 (N_345,In_1310,In_1947);
xnor U346 (N_346,In_888,In_1302);
nand U347 (N_347,In_1063,In_1102);
nand U348 (N_348,In_100,In_325);
xnor U349 (N_349,In_462,In_1228);
nor U350 (N_350,In_1815,In_1084);
or U351 (N_351,In_1612,In_89);
nand U352 (N_352,In_1428,In_1448);
or U353 (N_353,In_194,In_1512);
xor U354 (N_354,In_1162,In_1405);
and U355 (N_355,In_1046,In_1610);
and U356 (N_356,In_1410,In_1404);
or U357 (N_357,In_116,In_24);
and U358 (N_358,In_211,In_1275);
or U359 (N_359,In_374,In_399);
nand U360 (N_360,In_1354,In_1998);
nand U361 (N_361,In_98,In_400);
or U362 (N_362,In_658,In_317);
or U363 (N_363,In_617,In_642);
and U364 (N_364,In_1551,In_550);
nor U365 (N_365,In_931,In_1866);
xnor U366 (N_366,In_1924,In_1796);
nor U367 (N_367,In_803,In_339);
and U368 (N_368,In_1675,In_405);
nand U369 (N_369,In_992,In_523);
nand U370 (N_370,In_1653,In_994);
xor U371 (N_371,In_979,In_224);
and U372 (N_372,In_1465,In_947);
or U373 (N_373,In_314,In_1423);
or U374 (N_374,In_1369,In_1625);
or U375 (N_375,In_335,In_153);
and U376 (N_376,In_748,In_1633);
nand U377 (N_377,In_28,In_929);
nor U378 (N_378,In_943,In_461);
or U379 (N_379,In_1159,In_780);
nand U380 (N_380,In_414,In_198);
nor U381 (N_381,In_1123,In_769);
nor U382 (N_382,In_38,In_1875);
nor U383 (N_383,In_968,In_665);
or U384 (N_384,In_1476,In_66);
nor U385 (N_385,In_850,In_662);
and U386 (N_386,In_679,In_171);
or U387 (N_387,In_1628,In_1928);
xnor U388 (N_388,In_1887,In_492);
nand U389 (N_389,In_879,In_922);
nand U390 (N_390,In_1669,In_590);
xnor U391 (N_391,In_1604,In_1910);
nor U392 (N_392,In_1820,In_778);
xor U393 (N_393,In_1067,In_694);
and U394 (N_394,In_1905,In_509);
or U395 (N_395,In_1255,In_864);
nand U396 (N_396,In_713,In_160);
nor U397 (N_397,In_205,In_828);
xnor U398 (N_398,In_1685,In_155);
and U399 (N_399,In_1045,In_1039);
nor U400 (N_400,In_327,In_607);
xor U401 (N_401,In_1419,In_1916);
and U402 (N_402,In_719,In_261);
nor U403 (N_403,In_506,In_1157);
nor U404 (N_404,In_25,In_629);
and U405 (N_405,In_788,In_1799);
nor U406 (N_406,In_651,In_1739);
nand U407 (N_407,In_1631,In_1138);
and U408 (N_408,In_1836,In_1330);
or U409 (N_409,In_382,In_1882);
nor U410 (N_410,In_280,In_257);
and U411 (N_411,In_666,In_168);
or U412 (N_412,In_88,In_1868);
nand U413 (N_413,In_957,In_1092);
nand U414 (N_414,In_1214,In_250);
xnor U415 (N_415,In_225,In_366);
nor U416 (N_416,In_1532,In_1695);
nand U417 (N_417,In_1336,In_1469);
or U418 (N_418,In_1433,In_1574);
or U419 (N_419,In_1344,In_1972);
xnor U420 (N_420,In_927,In_1012);
nand U421 (N_421,In_1427,In_1074);
and U422 (N_422,In_529,In_308);
xor U423 (N_423,In_708,In_221);
nand U424 (N_424,In_182,In_1020);
xor U425 (N_425,In_561,In_822);
nand U426 (N_426,In_1487,In_151);
or U427 (N_427,In_1087,In_162);
xnor U428 (N_428,In_1019,In_608);
xor U429 (N_429,In_1043,In_1125);
nand U430 (N_430,In_1430,In_228);
xnor U431 (N_431,In_169,In_1496);
or U432 (N_432,In_1568,In_1714);
xnor U433 (N_433,In_580,In_129);
xnor U434 (N_434,In_1980,In_215);
or U435 (N_435,In_871,In_519);
and U436 (N_436,In_923,In_458);
or U437 (N_437,In_1447,In_938);
nor U438 (N_438,In_1449,In_861);
or U439 (N_439,In_1057,In_1222);
and U440 (N_440,In_1872,In_164);
and U441 (N_441,In_1422,In_1870);
nor U442 (N_442,In_1709,In_297);
xnor U443 (N_443,In_597,In_63);
nor U444 (N_444,In_1368,In_1388);
nand U445 (N_445,In_1741,In_177);
and U446 (N_446,In_1245,In_1538);
and U447 (N_447,In_232,In_156);
xnor U448 (N_448,In_488,In_336);
nand U449 (N_449,In_1395,In_826);
and U450 (N_450,In_701,In_1122);
xor U451 (N_451,In_1029,In_1109);
nor U452 (N_452,In_1420,In_1362);
or U453 (N_453,In_1795,In_1908);
and U454 (N_454,In_1003,In_1645);
nand U455 (N_455,In_0,In_1901);
and U456 (N_456,In_1779,In_1128);
or U457 (N_457,In_1287,In_625);
and U458 (N_458,In_1148,In_1749);
nand U459 (N_459,In_1191,In_1968);
or U460 (N_460,In_1907,In_1794);
nor U461 (N_461,In_1166,In_754);
xor U462 (N_462,In_20,In_296);
xor U463 (N_463,In_842,In_682);
nand U464 (N_464,In_1117,In_210);
or U465 (N_465,In_50,In_176);
xor U466 (N_466,In_857,In_1677);
and U467 (N_467,In_503,In_70);
xnor U468 (N_468,In_1156,In_411);
and U469 (N_469,In_1969,In_1204);
or U470 (N_470,In_771,In_85);
nand U471 (N_471,In_467,In_1221);
and U472 (N_472,In_80,In_235);
and U473 (N_473,In_290,In_1198);
nand U474 (N_474,In_1902,In_355);
and U475 (N_475,In_1725,In_1698);
xor U476 (N_476,In_524,In_1993);
or U477 (N_477,In_1624,In_138);
nand U478 (N_478,In_1925,In_1547);
xor U479 (N_479,In_764,In_1519);
or U480 (N_480,In_1254,In_1552);
xor U481 (N_481,In_1865,In_1942);
xnor U482 (N_482,In_1662,In_786);
and U483 (N_483,In_117,In_863);
and U484 (N_484,In_820,In_611);
or U485 (N_485,In_1856,In_1762);
nor U486 (N_486,In_1088,In_716);
or U487 (N_487,In_789,In_332);
xnor U488 (N_488,In_904,In_1491);
xor U489 (N_489,In_311,In_847);
or U490 (N_490,In_756,In_15);
or U491 (N_491,In_26,In_1782);
or U492 (N_492,In_533,In_1630);
and U493 (N_493,In_1587,In_1501);
nor U494 (N_494,In_1987,In_358);
or U495 (N_495,In_501,In_1736);
or U496 (N_496,In_1681,In_1000);
nor U497 (N_497,In_352,In_993);
xor U498 (N_498,In_102,In_481);
or U499 (N_499,In_486,In_1988);
nand U500 (N_500,In_346,In_190);
xor U501 (N_501,In_602,In_1316);
nand U502 (N_502,In_1667,In_552);
and U503 (N_503,In_251,In_200);
or U504 (N_504,In_1518,In_616);
nor U505 (N_505,In_1387,In_984);
and U506 (N_506,In_1006,In_219);
xnor U507 (N_507,In_1718,In_1324);
nand U508 (N_508,In_22,In_470);
or U509 (N_509,In_271,In_1365);
and U510 (N_510,In_587,In_906);
nor U511 (N_511,In_377,In_1513);
nand U512 (N_512,In_977,In_242);
nor U513 (N_513,In_852,In_278);
xor U514 (N_514,In_544,In_765);
or U515 (N_515,In_436,In_647);
or U516 (N_516,In_141,In_256);
or U517 (N_517,In_933,In_1136);
nand U518 (N_518,In_32,In_884);
and U519 (N_519,In_548,In_880);
nand U520 (N_520,In_79,In_1358);
nor U521 (N_521,In_410,In_1234);
nor U522 (N_522,In_111,In_500);
nor U523 (N_523,In_1441,In_342);
and U524 (N_524,In_1703,In_1431);
xnor U525 (N_525,In_68,In_830);
nor U526 (N_526,In_833,In_338);
nand U527 (N_527,In_808,In_1146);
or U528 (N_528,In_1626,In_1065);
xor U529 (N_529,In_1456,In_1598);
xnor U530 (N_530,In_1804,In_989);
xnor U531 (N_531,In_1818,In_1121);
and U532 (N_532,In_1451,In_1064);
nor U533 (N_533,In_696,In_686);
nor U534 (N_534,In_1027,In_1713);
nand U535 (N_535,In_1883,In_173);
or U536 (N_536,In_542,In_1378);
nor U537 (N_537,In_965,In_1266);
nand U538 (N_538,In_233,In_150);
nand U539 (N_539,In_1096,In_1244);
nand U540 (N_540,In_834,In_1576);
or U541 (N_541,In_365,In_1759);
or U542 (N_542,In_343,In_695);
and U543 (N_543,In_1575,In_144);
nor U544 (N_544,In_601,In_212);
nor U545 (N_545,In_1867,In_301);
nand U546 (N_546,In_940,In_1893);
xnor U547 (N_547,In_831,In_1060);
xor U548 (N_548,In_1413,In_1535);
and U549 (N_549,In_1284,In_199);
and U550 (N_550,In_1114,In_1445);
nor U551 (N_551,In_1647,In_333);
nand U552 (N_552,In_1260,In_1680);
or U553 (N_553,In_895,In_521);
xnor U554 (N_554,In_305,In_295);
nand U555 (N_555,In_430,In_1132);
nor U556 (N_556,In_1817,In_401);
or U557 (N_557,In_746,In_1478);
and U558 (N_558,In_1265,In_851);
and U559 (N_559,In_1107,In_490);
nand U560 (N_560,In_722,In_331);
xor U561 (N_561,In_1296,In_567);
nor U562 (N_562,In_1186,In_1393);
or U563 (N_563,In_1183,In_81);
xor U564 (N_564,In_1417,In_1840);
or U565 (N_565,In_637,In_1450);
xor U566 (N_566,In_1937,In_1089);
xnor U567 (N_567,In_39,In_64);
xnor U568 (N_568,In_1982,In_441);
xor U569 (N_569,In_1566,In_1786);
nor U570 (N_570,In_793,In_460);
xnor U571 (N_571,In_1812,In_1165);
or U572 (N_572,In_1201,In_869);
xnor U573 (N_573,In_217,In_312);
xnor U574 (N_574,In_1061,In_1616);
nor U575 (N_575,In_733,In_361);
nor U576 (N_576,In_1689,In_324);
nor U577 (N_577,In_734,In_105);
nor U578 (N_578,In_1139,In_359);
or U579 (N_579,In_59,In_976);
nor U580 (N_580,In_442,In_1374);
nand U581 (N_581,In_646,In_1673);
nand U582 (N_582,In_1627,In_667);
nand U583 (N_583,In_1153,In_1268);
nand U584 (N_584,In_1416,In_1317);
nand U585 (N_585,In_16,In_1343);
nor U586 (N_586,In_883,In_657);
xnor U587 (N_587,In_114,In_823);
xor U588 (N_588,In_1203,In_800);
nor U589 (N_589,In_570,In_956);
or U590 (N_590,In_1594,In_329);
nand U591 (N_591,In_1648,In_555);
nand U592 (N_592,In_1700,In_1112);
nor U593 (N_593,In_538,In_1299);
or U594 (N_594,In_368,In_853);
xnor U595 (N_595,In_844,In_367);
and U596 (N_596,In_1364,In_1609);
xnor U597 (N_597,In_1750,In_18);
and U598 (N_598,In_1705,In_1018);
and U599 (N_599,In_499,In_37);
xnor U600 (N_600,In_1965,In_1522);
nand U601 (N_601,In_1504,In_801);
nor U602 (N_602,In_1632,In_1325);
or U603 (N_603,In_10,In_1315);
nand U604 (N_604,In_849,In_1955);
or U605 (N_605,In_1007,In_728);
or U606 (N_606,In_614,In_612);
and U607 (N_607,In_964,In_372);
and U608 (N_608,In_687,In_1178);
xnor U609 (N_609,In_1075,In_179);
xnor U610 (N_610,In_1959,In_1394);
nor U611 (N_611,In_41,In_525);
or U612 (N_612,In_553,In_1391);
or U613 (N_613,In_1684,In_618);
xnor U614 (N_614,In_421,In_303);
nor U615 (N_615,In_449,In_737);
and U616 (N_616,In_1772,In_1545);
nand U617 (N_617,In_19,In_1208);
nor U618 (N_618,In_724,In_1119);
or U619 (N_619,In_910,In_1541);
xnor U620 (N_620,In_1436,In_1913);
and U621 (N_621,In_480,In_148);
and U622 (N_622,In_285,In_1670);
nor U623 (N_623,In_1055,In_1269);
xnor U624 (N_624,In_1826,In_630);
nor U625 (N_625,In_1406,In_1141);
and U626 (N_626,In_197,In_1555);
nor U627 (N_627,In_838,In_896);
nand U628 (N_628,In_258,In_796);
and U629 (N_629,In_663,In_1338);
or U630 (N_630,In_1193,In_574);
xnor U631 (N_631,In_974,In_711);
nand U632 (N_632,In_868,In_1819);
or U633 (N_633,In_804,In_504);
and U634 (N_634,In_1657,In_732);
nor U635 (N_635,In_596,In_1650);
and U636 (N_636,In_121,In_505);
xnor U637 (N_637,In_1332,In_564);
or U638 (N_638,In_415,In_1884);
nor U639 (N_639,In_1842,In_275);
and U640 (N_640,In_1492,In_1949);
xor U641 (N_641,In_1622,In_1671);
and U642 (N_642,In_932,In_1147);
and U643 (N_643,In_103,In_621);
nand U644 (N_644,In_72,In_792);
nor U645 (N_645,In_790,In_489);
xor U646 (N_646,In_1206,In_537);
nand U647 (N_647,In_1717,In_447);
xor U648 (N_648,In_1215,In_1641);
nor U649 (N_649,In_87,In_1898);
nand U650 (N_650,In_1923,In_901);
or U651 (N_651,In_829,In_1077);
xor U652 (N_652,In_158,In_1326);
or U653 (N_653,In_958,In_451);
nor U654 (N_654,In_1373,In_785);
nor U655 (N_655,In_1116,In_1078);
or U656 (N_656,In_1640,In_999);
nand U657 (N_657,In_1097,In_560);
nand U658 (N_658,In_1327,In_61);
nand U659 (N_659,In_1199,In_184);
nand U660 (N_660,In_1780,In_1546);
nand U661 (N_661,In_1502,In_371);
nand U662 (N_662,In_459,In_360);
nand U663 (N_663,In_936,In_791);
or U664 (N_664,In_1964,In_860);
or U665 (N_665,In_572,In_180);
xor U666 (N_666,In_652,In_181);
nor U667 (N_667,In_1498,In_286);
nand U668 (N_668,In_907,In_373);
and U669 (N_669,In_924,In_1182);
nor U670 (N_670,In_1375,In_1531);
nand U671 (N_671,In_1983,In_344);
or U672 (N_672,In_43,In_1085);
nand U673 (N_673,In_1767,In_515);
nand U674 (N_674,In_1683,In_1805);
or U675 (N_675,In_1811,In_975);
or U676 (N_676,In_1131,In_1754);
and U677 (N_677,In_139,In_738);
xnor U678 (N_678,In_354,In_835);
nand U679 (N_679,In_51,In_762);
nor U680 (N_680,In_1345,In_429);
nand U681 (N_681,In_1537,In_1822);
nand U682 (N_682,In_322,In_518);
nand U683 (N_683,In_1050,In_1572);
nand U684 (N_684,In_1164,In_690);
nand U685 (N_685,In_745,In_1108);
nor U686 (N_686,In_705,In_600);
and U687 (N_687,In_299,In_982);
and U688 (N_688,In_921,In_1446);
or U689 (N_689,In_319,In_905);
and U690 (N_690,In_163,In_986);
nand U691 (N_691,In_1728,In_453);
nand U692 (N_692,In_1389,In_17);
nand U693 (N_693,In_751,In_252);
or U694 (N_694,In_11,In_1454);
xnor U695 (N_695,In_1457,In_632);
nand U696 (N_696,In_1747,In_1943);
or U697 (N_697,In_653,In_403);
and U698 (N_698,In_1170,In_1860);
or U699 (N_699,In_1239,In_340);
or U700 (N_700,In_972,In_1526);
xnor U701 (N_701,In_817,In_1752);
xor U702 (N_702,In_980,In_477);
or U703 (N_703,In_432,In_313);
nor U704 (N_704,In_165,In_1966);
nor U705 (N_705,In_1298,In_752);
nand U706 (N_706,In_1272,In_142);
nor U707 (N_707,In_1733,In_1912);
nand U708 (N_708,In_364,In_1418);
and U709 (N_709,In_230,In_1542);
nor U710 (N_710,In_1783,In_1731);
nand U711 (N_711,In_29,In_112);
xnor U712 (N_712,In_1120,In_1793);
xnor U713 (N_713,In_589,In_603);
nand U714 (N_714,In_573,In_1026);
xor U715 (N_715,In_476,In_760);
or U716 (N_716,In_1758,In_717);
xor U717 (N_717,In_1070,In_1303);
and U718 (N_718,In_431,In_512);
nand U719 (N_719,In_1726,In_832);
and U720 (N_720,In_1527,In_1847);
nor U721 (N_721,In_1056,In_1424);
nand U722 (N_722,In_1008,In_1593);
or U723 (N_723,In_1495,In_1090);
nor U724 (N_724,In_1991,In_1331);
or U725 (N_725,In_418,In_1696);
nor U726 (N_726,In_1174,In_130);
nand U727 (N_727,In_990,In_973);
and U728 (N_728,In_1207,In_1263);
xor U729 (N_729,In_1978,In_1321);
and U730 (N_730,In_236,In_1278);
and U731 (N_731,In_758,In_1933);
or U732 (N_732,In_283,In_766);
xnor U733 (N_733,In_1939,In_119);
nor U734 (N_734,In_1335,In_268);
or U735 (N_735,In_565,In_1693);
nor U736 (N_736,In_1248,In_260);
xor U737 (N_737,In_389,In_1506);
or U738 (N_738,In_731,In_1459);
or U739 (N_739,In_1024,In_925);
nand U740 (N_740,In_1383,In_1262);
or U741 (N_741,In_912,In_1442);
or U742 (N_742,In_1367,In_604);
nor U743 (N_743,In_911,In_891);
nor U744 (N_744,In_1590,In_681);
xor U745 (N_745,In_1909,In_334);
xor U746 (N_746,In_207,In_1280);
and U747 (N_747,In_767,In_95);
and U748 (N_748,In_784,In_1036);
and U749 (N_749,In_541,In_1716);
nor U750 (N_750,In_1237,In_1435);
and U751 (N_751,In_569,In_1401);
or U752 (N_752,In_1629,In_1274);
nor U753 (N_753,In_485,In_6);
xnor U754 (N_754,In_777,In_267);
nor U755 (N_755,In_1597,In_1619);
and U756 (N_756,In_759,In_1540);
nand U757 (N_757,In_613,In_1086);
xor U758 (N_758,In_469,In_1850);
nand U759 (N_759,In_636,In_408);
and U760 (N_760,In_1253,In_413);
xor U761 (N_761,In_843,In_1171);
nor U762 (N_762,In_1352,In_1585);
nand U763 (N_763,In_27,In_648);
or U764 (N_764,In_807,In_1444);
nor U765 (N_765,In_586,In_1859);
xnor U766 (N_766,In_1956,In_645);
xnor U767 (N_767,In_443,In_191);
and U768 (N_768,In_1879,In_1553);
and U769 (N_769,In_799,In_874);
nor U770 (N_770,In_1748,In_1611);
xor U771 (N_771,In_1443,In_1438);
xnor U772 (N_772,In_1037,In_1511);
nand U773 (N_773,In_277,In_1356);
nor U774 (N_774,In_839,In_1886);
nor U775 (N_775,In_1099,In_855);
nand U776 (N_776,In_1161,In_1742);
or U777 (N_777,In_1740,In_1777);
nand U778 (N_778,In_1306,In_1073);
nand U779 (N_779,In_1603,In_439);
nand U780 (N_780,In_82,In_1871);
nand U781 (N_781,In_1175,In_1785);
nand U782 (N_782,In_1602,In_292);
nor U783 (N_783,In_304,In_605);
xnor U784 (N_784,In_1833,In_1098);
or U785 (N_785,In_1734,In_692);
or U786 (N_786,In_899,In_206);
xor U787 (N_787,In_949,In_1062);
xor U788 (N_788,In_1851,In_406);
nand U789 (N_789,In_1784,In_1646);
or U790 (N_790,In_837,In_742);
xnor U791 (N_791,In_1311,In_1353);
or U792 (N_792,In_644,In_1549);
and U793 (N_793,In_1791,In_622);
nor U794 (N_794,In_1813,In_62);
xor U795 (N_795,In_1954,In_1661);
nand U796 (N_796,In_1486,In_1521);
xor U797 (N_797,In_31,In_1558);
or U798 (N_798,In_919,In_1895);
and U799 (N_799,In_1803,In_757);
xnor U800 (N_800,In_726,In_1678);
and U801 (N_801,In_1202,In_387);
and U802 (N_802,In_635,In_1855);
or U803 (N_803,In_315,In_1571);
xor U804 (N_804,In_1106,In_1184);
xnor U805 (N_805,In_496,In_482);
or U806 (N_806,In_1205,In_1231);
nor U807 (N_807,In_1200,In_1474);
xor U808 (N_808,In_1009,In_1973);
or U809 (N_809,In_985,In_693);
xnor U810 (N_810,In_1591,In_1118);
and U811 (N_811,In_350,In_487);
nand U812 (N_812,In_1225,In_1091);
nor U813 (N_813,In_281,In_571);
and U814 (N_814,In_714,In_730);
xnor U815 (N_815,In_76,In_1480);
or U816 (N_816,In_937,In_699);
xor U817 (N_817,In_628,In_1848);
xor U818 (N_818,In_581,In_69);
xor U819 (N_819,In_935,In_1144);
or U820 (N_820,In_702,In_1596);
or U821 (N_821,In_3,In_510);
nand U822 (N_822,In_381,In_133);
xor U823 (N_823,In_669,In_812);
nor U824 (N_824,In_349,In_806);
nand U825 (N_825,In_881,In_641);
or U826 (N_826,In_1807,In_1642);
and U827 (N_827,In_53,In_1960);
or U828 (N_828,In_192,In_916);
or U829 (N_829,In_1054,In_718);
nor U830 (N_830,In_854,In_12);
or U831 (N_831,In_813,In_1892);
nand U832 (N_832,In_465,In_824);
xor U833 (N_833,In_1584,In_858);
and U834 (N_834,In_1737,In_1516);
or U835 (N_835,In_1415,In_1104);
nor U836 (N_836,In_1790,In_123);
xnor U837 (N_837,In_1915,In_1468);
nor U838 (N_838,In_1032,In_1305);
nor U839 (N_839,In_237,In_970);
nand U840 (N_840,In_94,In_1314);
nand U841 (N_841,In_1158,In_452);
nand U842 (N_842,In_638,In_588);
nor U843 (N_843,In_189,In_741);
or U844 (N_844,In_1223,In_1607);
or U845 (N_845,In_222,In_1567);
or U846 (N_846,In_1533,In_706);
nor U847 (N_847,In_633,In_455);
or U848 (N_848,In_1525,In_516);
nor U849 (N_849,In_952,In_825);
or U850 (N_850,In_744,In_556);
nand U851 (N_851,In_1115,In_115);
or U852 (N_852,In_703,In_707);
and U853 (N_853,In_1846,In_1355);
nand U854 (N_854,In_1687,In_1932);
xor U855 (N_855,In_298,In_1180);
or U856 (N_856,In_118,In_152);
or U857 (N_857,In_1047,In_928);
or U858 (N_858,In_535,In_961);
nand U859 (N_859,In_971,In_1058);
nand U860 (N_860,In_1523,In_188);
xnor U861 (N_861,In_1753,In_1071);
nand U862 (N_862,In_282,In_1093);
nand U863 (N_863,In_167,In_1294);
xnor U864 (N_864,In_1429,In_398);
nor U865 (N_865,In_772,In_1163);
nand U866 (N_866,In_1515,In_1635);
and U867 (N_867,In_1361,In_1724);
or U868 (N_868,In_1398,In_126);
nor U869 (N_869,In_1295,In_147);
and U870 (N_870,In_108,In_1409);
nand U871 (N_871,In_865,In_1719);
nor U872 (N_872,In_1798,In_348);
nor U873 (N_873,In_201,In_423);
nand U874 (N_874,In_1432,In_585);
and U875 (N_875,In_127,In_634);
nor U876 (N_876,In_1227,In_1342);
xor U877 (N_877,In_1151,In_1341);
or U878 (N_878,In_1076,In_239);
nand U879 (N_879,In_60,In_1240);
nand U880 (N_880,In_1488,In_178);
xnor U881 (N_881,In_942,In_606);
xnor U882 (N_882,In_1814,In_175);
nor U883 (N_883,In_1613,In_33);
and U884 (N_884,In_988,In_259);
nand U885 (N_885,In_378,In_1082);
and U886 (N_886,In_1130,In_1386);
or U887 (N_887,In_1172,In_1852);
nand U888 (N_888,In_1543,In_379);
nor U889 (N_889,In_1744,In_710);
nor U890 (N_890,In_563,In_514);
nand U891 (N_891,In_14,In_71);
and U892 (N_892,In_1481,In_73);
nand U893 (N_893,In_1482,In_1825);
xnor U894 (N_894,In_1359,In_170);
and U895 (N_895,In_55,In_736);
or U896 (N_896,In_1004,In_1881);
or U897 (N_897,In_1940,In_1658);
nand U898 (N_898,In_1500,In_479);
xor U899 (N_899,In_1564,In_122);
xor U900 (N_900,In_661,In_1580);
nand U901 (N_901,In_688,In_1989);
nand U902 (N_902,In_1181,In_1453);
or U903 (N_903,In_809,In_1219);
xor U904 (N_904,In_1483,In_272);
or U905 (N_905,In_396,In_1357);
or U906 (N_906,In_1528,In_540);
nor U907 (N_907,In_1950,In_1845);
nand U908 (N_908,In_110,In_1903);
nand U909 (N_909,In_1926,In_1957);
or U910 (N_910,In_1664,In_562);
xor U911 (N_911,In_1618,In_394);
and U912 (N_912,In_1218,In_1113);
and U913 (N_913,In_1711,In_576);
and U914 (N_914,In_814,In_755);
xnor U915 (N_915,In_1655,In_1127);
xnor U916 (N_916,In_13,In_1414);
nor U917 (N_917,In_867,In_897);
or U918 (N_918,In_805,In_1103);
and U919 (N_919,In_265,In_146);
nor U920 (N_920,In_52,In_639);
nand U921 (N_921,In_227,In_1304);
nor U922 (N_922,In_1573,In_677);
nor U923 (N_923,In_654,In_1539);
or U924 (N_924,In_893,In_593);
and U925 (N_925,In_1232,In_1691);
and U926 (N_926,In_1015,In_54);
or U927 (N_927,In_1755,In_1407);
nor U928 (N_928,In_1030,In_619);
or U929 (N_929,In_166,In_1300);
nor U930 (N_930,In_1279,In_1023);
nor U931 (N_931,In_1702,In_416);
nor U932 (N_932,In_846,In_1900);
and U933 (N_933,In_128,In_74);
nand U934 (N_934,In_783,In_691);
nor U935 (N_935,In_84,In_1038);
nand U936 (N_936,In_67,In_953);
and U937 (N_937,In_1230,In_1863);
and U938 (N_938,In_1679,In_248);
or U939 (N_939,In_675,In_743);
xor U940 (N_940,In_1559,In_1929);
or U941 (N_941,In_1124,In_750);
nand U942 (N_942,In_1411,In_456);
nand U943 (N_943,In_243,In_1821);
nor U944 (N_944,In_1579,In_1179);
xnor U945 (N_945,In_676,In_1701);
xnor U946 (N_946,In_1831,In_466);
nor U947 (N_947,In_419,In_598);
and U948 (N_948,In_960,In_136);
nor U949 (N_949,In_1399,In_412);
nor U950 (N_950,In_683,In_787);
or U951 (N_951,In_1621,In_1440);
nand U952 (N_952,In_1577,In_1849);
nand U953 (N_953,In_213,In_1911);
or U954 (N_954,In_944,In_1243);
or U955 (N_955,In_5,In_1864);
nor U956 (N_956,In_131,In_376);
and U957 (N_957,In_229,In_1745);
nor U958 (N_958,In_445,In_353);
or U959 (N_959,In_1101,In_810);
nand U960 (N_960,In_1563,In_241);
nand U961 (N_961,In_913,In_1238);
xnor U962 (N_962,In_457,In_1392);
nor U963 (N_963,In_532,In_1769);
nor U964 (N_964,In_1994,In_1930);
nor U965 (N_965,In_1919,In_1377);
or U966 (N_966,In_1301,In_1668);
xnor U967 (N_967,In_712,In_434);
xnor U968 (N_968,In_1896,In_1839);
nor U969 (N_969,In_203,In_721);
nor U970 (N_970,In_1384,In_725);
nor U971 (N_971,In_1349,In_1775);
nand U972 (N_972,In_1743,In_1049);
or U973 (N_973,In_877,In_390);
or U974 (N_974,In_1801,In_1307);
nand U975 (N_975,In_1760,In_775);
and U976 (N_976,In_1756,In_1323);
and U977 (N_977,In_1464,In_92);
nor U978 (N_978,In_1288,In_1382);
xnor U979 (N_979,In_763,In_484);
nand U980 (N_980,In_383,In_1583);
and U981 (N_981,In_137,In_1509);
nor U982 (N_982,In_715,In_196);
nand U983 (N_983,In_1229,In_1636);
nand U984 (N_984,In_1707,In_75);
or U985 (N_985,In_1028,In_1339);
xor U986 (N_986,In_395,In_1160);
or U987 (N_987,In_1606,In_1466);
xor U988 (N_988,In_1434,In_1854);
nor U989 (N_989,In_1827,In_520);
or U990 (N_990,In_1135,In_643);
xor U991 (N_991,In_109,In_909);
nand U992 (N_992,In_134,In_1710);
or U993 (N_993,In_1286,In_1874);
and U994 (N_994,In_463,In_1674);
nor U995 (N_995,In_409,In_1360);
nor U996 (N_996,In_255,In_1289);
nor U997 (N_997,In_1996,In_1285);
nand U998 (N_998,In_266,In_93);
xnor U999 (N_999,In_300,In_1402);
xor U1000 (N_1000,In_596,In_1363);
and U1001 (N_1001,In_904,In_1338);
xor U1002 (N_1002,In_555,In_56);
nand U1003 (N_1003,In_1124,In_964);
nor U1004 (N_1004,In_903,In_486);
nor U1005 (N_1005,In_1169,In_439);
nand U1006 (N_1006,In_1444,In_74);
nand U1007 (N_1007,In_743,In_1342);
nand U1008 (N_1008,In_669,In_1103);
nor U1009 (N_1009,In_623,In_564);
nor U1010 (N_1010,In_855,In_416);
or U1011 (N_1011,In_448,In_1427);
nand U1012 (N_1012,In_1774,In_724);
and U1013 (N_1013,In_344,In_1469);
nor U1014 (N_1014,In_23,In_1996);
and U1015 (N_1015,In_702,In_1027);
nand U1016 (N_1016,In_1526,In_1521);
xnor U1017 (N_1017,In_1662,In_215);
or U1018 (N_1018,In_421,In_1163);
nand U1019 (N_1019,In_1642,In_1448);
nor U1020 (N_1020,In_869,In_432);
and U1021 (N_1021,In_1487,In_830);
or U1022 (N_1022,In_1902,In_836);
nor U1023 (N_1023,In_481,In_1836);
or U1024 (N_1024,In_276,In_1019);
nand U1025 (N_1025,In_71,In_365);
nor U1026 (N_1026,In_1424,In_866);
nor U1027 (N_1027,In_1169,In_1);
xnor U1028 (N_1028,In_1937,In_100);
and U1029 (N_1029,In_810,In_414);
nor U1030 (N_1030,In_385,In_413);
and U1031 (N_1031,In_404,In_325);
xor U1032 (N_1032,In_1327,In_528);
xnor U1033 (N_1033,In_412,In_587);
xnor U1034 (N_1034,In_337,In_346);
nand U1035 (N_1035,In_531,In_38);
nor U1036 (N_1036,In_1006,In_1762);
xnor U1037 (N_1037,In_1128,In_500);
xnor U1038 (N_1038,In_1444,In_805);
and U1039 (N_1039,In_320,In_1350);
xor U1040 (N_1040,In_520,In_293);
xnor U1041 (N_1041,In_1446,In_1792);
and U1042 (N_1042,In_1082,In_1833);
nand U1043 (N_1043,In_95,In_1743);
nor U1044 (N_1044,In_442,In_1450);
or U1045 (N_1045,In_1006,In_831);
xnor U1046 (N_1046,In_1204,In_1426);
nand U1047 (N_1047,In_1754,In_258);
and U1048 (N_1048,In_621,In_1454);
nand U1049 (N_1049,In_111,In_1007);
or U1050 (N_1050,In_938,In_852);
nand U1051 (N_1051,In_444,In_1719);
xor U1052 (N_1052,In_354,In_1444);
nor U1053 (N_1053,In_1928,In_199);
nand U1054 (N_1054,In_1720,In_1597);
or U1055 (N_1055,In_771,In_880);
nor U1056 (N_1056,In_778,In_998);
nor U1057 (N_1057,In_1017,In_84);
nor U1058 (N_1058,In_1341,In_1141);
xor U1059 (N_1059,In_1958,In_1591);
xor U1060 (N_1060,In_1482,In_212);
and U1061 (N_1061,In_1193,In_1796);
and U1062 (N_1062,In_651,In_468);
or U1063 (N_1063,In_1573,In_374);
or U1064 (N_1064,In_563,In_1016);
xnor U1065 (N_1065,In_1592,In_24);
and U1066 (N_1066,In_511,In_545);
or U1067 (N_1067,In_749,In_260);
nand U1068 (N_1068,In_316,In_1746);
xor U1069 (N_1069,In_378,In_119);
nand U1070 (N_1070,In_898,In_1235);
or U1071 (N_1071,In_1306,In_240);
or U1072 (N_1072,In_557,In_267);
nand U1073 (N_1073,In_640,In_1659);
and U1074 (N_1074,In_497,In_1799);
or U1075 (N_1075,In_1448,In_161);
and U1076 (N_1076,In_1814,In_433);
and U1077 (N_1077,In_957,In_1661);
nor U1078 (N_1078,In_1693,In_1775);
nand U1079 (N_1079,In_712,In_629);
and U1080 (N_1080,In_1270,In_1803);
nor U1081 (N_1081,In_1867,In_944);
and U1082 (N_1082,In_1399,In_1165);
and U1083 (N_1083,In_1301,In_1827);
nand U1084 (N_1084,In_277,In_1286);
nand U1085 (N_1085,In_1294,In_1812);
xnor U1086 (N_1086,In_1336,In_1879);
and U1087 (N_1087,In_96,In_1180);
nor U1088 (N_1088,In_1151,In_150);
or U1089 (N_1089,In_892,In_1846);
nand U1090 (N_1090,In_434,In_439);
and U1091 (N_1091,In_899,In_26);
and U1092 (N_1092,In_1771,In_1232);
nand U1093 (N_1093,In_1619,In_716);
nor U1094 (N_1094,In_1767,In_292);
or U1095 (N_1095,In_1190,In_337);
or U1096 (N_1096,In_1365,In_1360);
nand U1097 (N_1097,In_1723,In_415);
nand U1098 (N_1098,In_301,In_1427);
and U1099 (N_1099,In_949,In_279);
xnor U1100 (N_1100,In_1298,In_1386);
nor U1101 (N_1101,In_917,In_1660);
and U1102 (N_1102,In_667,In_1688);
or U1103 (N_1103,In_1380,In_915);
xor U1104 (N_1104,In_1999,In_1195);
nand U1105 (N_1105,In_1368,In_1326);
xnor U1106 (N_1106,In_1862,In_1381);
nor U1107 (N_1107,In_1815,In_646);
xor U1108 (N_1108,In_184,In_1218);
or U1109 (N_1109,In_453,In_1405);
or U1110 (N_1110,In_467,In_1655);
xnor U1111 (N_1111,In_191,In_815);
nand U1112 (N_1112,In_321,In_174);
xnor U1113 (N_1113,In_1843,In_1482);
nor U1114 (N_1114,In_202,In_1660);
and U1115 (N_1115,In_1431,In_824);
xnor U1116 (N_1116,In_1115,In_1301);
nor U1117 (N_1117,In_598,In_1718);
nand U1118 (N_1118,In_711,In_265);
or U1119 (N_1119,In_583,In_11);
nand U1120 (N_1120,In_1201,In_1311);
nand U1121 (N_1121,In_1242,In_634);
and U1122 (N_1122,In_727,In_1623);
nand U1123 (N_1123,In_1662,In_534);
xnor U1124 (N_1124,In_613,In_560);
or U1125 (N_1125,In_1432,In_1399);
nor U1126 (N_1126,In_475,In_707);
and U1127 (N_1127,In_780,In_879);
nor U1128 (N_1128,In_1646,In_537);
nor U1129 (N_1129,In_1822,In_835);
and U1130 (N_1130,In_1136,In_1636);
nor U1131 (N_1131,In_1127,In_1487);
nor U1132 (N_1132,In_23,In_465);
nor U1133 (N_1133,In_567,In_701);
or U1134 (N_1134,In_971,In_1696);
xnor U1135 (N_1135,In_1477,In_390);
and U1136 (N_1136,In_1273,In_631);
and U1137 (N_1137,In_1458,In_907);
nand U1138 (N_1138,In_1063,In_1184);
or U1139 (N_1139,In_620,In_1574);
xor U1140 (N_1140,In_1237,In_1537);
nor U1141 (N_1141,In_641,In_380);
xor U1142 (N_1142,In_776,In_95);
xnor U1143 (N_1143,In_703,In_309);
and U1144 (N_1144,In_739,In_1024);
nor U1145 (N_1145,In_1145,In_1692);
nor U1146 (N_1146,In_758,In_1831);
or U1147 (N_1147,In_889,In_1241);
xnor U1148 (N_1148,In_1418,In_320);
nor U1149 (N_1149,In_1923,In_1110);
nor U1150 (N_1150,In_826,In_168);
nor U1151 (N_1151,In_1666,In_168);
and U1152 (N_1152,In_668,In_1861);
nor U1153 (N_1153,In_1535,In_1308);
nand U1154 (N_1154,In_410,In_740);
or U1155 (N_1155,In_878,In_820);
and U1156 (N_1156,In_1752,In_659);
nand U1157 (N_1157,In_207,In_843);
xor U1158 (N_1158,In_1116,In_1904);
xnor U1159 (N_1159,In_1275,In_932);
xor U1160 (N_1160,In_460,In_719);
nor U1161 (N_1161,In_273,In_459);
nor U1162 (N_1162,In_1822,In_1759);
or U1163 (N_1163,In_67,In_694);
and U1164 (N_1164,In_286,In_426);
nand U1165 (N_1165,In_1524,In_1420);
xor U1166 (N_1166,In_49,In_1475);
or U1167 (N_1167,In_717,In_1677);
or U1168 (N_1168,In_1414,In_908);
and U1169 (N_1169,In_1167,In_169);
xor U1170 (N_1170,In_1182,In_6);
nand U1171 (N_1171,In_700,In_444);
or U1172 (N_1172,In_1263,In_1905);
nand U1173 (N_1173,In_1011,In_679);
nor U1174 (N_1174,In_944,In_1617);
or U1175 (N_1175,In_711,In_1784);
or U1176 (N_1176,In_1426,In_1029);
and U1177 (N_1177,In_1911,In_1488);
nor U1178 (N_1178,In_1408,In_1466);
nand U1179 (N_1179,In_961,In_1955);
nor U1180 (N_1180,In_758,In_615);
nor U1181 (N_1181,In_1246,In_580);
or U1182 (N_1182,In_1431,In_1199);
nand U1183 (N_1183,In_906,In_848);
and U1184 (N_1184,In_1922,In_1572);
or U1185 (N_1185,In_1075,In_1535);
and U1186 (N_1186,In_1724,In_751);
nand U1187 (N_1187,In_1149,In_647);
nor U1188 (N_1188,In_1135,In_436);
nor U1189 (N_1189,In_642,In_261);
and U1190 (N_1190,In_12,In_1633);
nor U1191 (N_1191,In_815,In_396);
and U1192 (N_1192,In_1244,In_415);
and U1193 (N_1193,In_1335,In_1178);
nand U1194 (N_1194,In_253,In_591);
and U1195 (N_1195,In_863,In_1278);
and U1196 (N_1196,In_1457,In_1602);
nor U1197 (N_1197,In_1915,In_773);
and U1198 (N_1198,In_1379,In_1344);
or U1199 (N_1199,In_473,In_458);
nor U1200 (N_1200,In_1101,In_1719);
nor U1201 (N_1201,In_1460,In_1960);
nand U1202 (N_1202,In_1711,In_1769);
or U1203 (N_1203,In_16,In_384);
or U1204 (N_1204,In_1499,In_609);
nand U1205 (N_1205,In_479,In_1314);
nor U1206 (N_1206,In_1466,In_1123);
xnor U1207 (N_1207,In_142,In_1232);
nor U1208 (N_1208,In_922,In_709);
xor U1209 (N_1209,In_954,In_721);
nor U1210 (N_1210,In_1437,In_1490);
nand U1211 (N_1211,In_277,In_1101);
and U1212 (N_1212,In_1628,In_269);
and U1213 (N_1213,In_761,In_402);
or U1214 (N_1214,In_1232,In_1150);
xor U1215 (N_1215,In_253,In_1628);
nand U1216 (N_1216,In_297,In_991);
or U1217 (N_1217,In_928,In_476);
and U1218 (N_1218,In_388,In_195);
or U1219 (N_1219,In_178,In_812);
nor U1220 (N_1220,In_798,In_1287);
xnor U1221 (N_1221,In_1768,In_838);
nand U1222 (N_1222,In_1758,In_1186);
xnor U1223 (N_1223,In_1044,In_347);
nor U1224 (N_1224,In_218,In_1713);
nor U1225 (N_1225,In_802,In_1846);
nand U1226 (N_1226,In_580,In_1058);
and U1227 (N_1227,In_512,In_441);
or U1228 (N_1228,In_1392,In_1555);
nand U1229 (N_1229,In_259,In_1350);
and U1230 (N_1230,In_1241,In_1244);
xor U1231 (N_1231,In_412,In_1112);
nor U1232 (N_1232,In_543,In_1357);
and U1233 (N_1233,In_994,In_1179);
nor U1234 (N_1234,In_1586,In_5);
nor U1235 (N_1235,In_1571,In_1448);
or U1236 (N_1236,In_138,In_1687);
or U1237 (N_1237,In_9,In_1288);
xnor U1238 (N_1238,In_1769,In_882);
nor U1239 (N_1239,In_445,In_286);
nor U1240 (N_1240,In_1761,In_94);
and U1241 (N_1241,In_820,In_1353);
nand U1242 (N_1242,In_1440,In_1511);
nor U1243 (N_1243,In_668,In_1052);
nand U1244 (N_1244,In_612,In_1274);
or U1245 (N_1245,In_368,In_777);
or U1246 (N_1246,In_35,In_1297);
nor U1247 (N_1247,In_324,In_1125);
xnor U1248 (N_1248,In_1611,In_826);
and U1249 (N_1249,In_129,In_1204);
and U1250 (N_1250,In_1269,In_923);
nand U1251 (N_1251,In_407,In_1238);
nand U1252 (N_1252,In_1521,In_1246);
nand U1253 (N_1253,In_1884,In_399);
nor U1254 (N_1254,In_87,In_525);
xor U1255 (N_1255,In_1139,In_896);
or U1256 (N_1256,In_1218,In_1970);
or U1257 (N_1257,In_132,In_1202);
and U1258 (N_1258,In_311,In_1373);
nor U1259 (N_1259,In_97,In_1419);
nand U1260 (N_1260,In_1908,In_1474);
and U1261 (N_1261,In_75,In_1589);
or U1262 (N_1262,In_642,In_355);
xor U1263 (N_1263,In_514,In_329);
or U1264 (N_1264,In_256,In_995);
xnor U1265 (N_1265,In_677,In_1930);
nand U1266 (N_1266,In_1072,In_806);
nor U1267 (N_1267,In_64,In_749);
or U1268 (N_1268,In_898,In_1942);
nand U1269 (N_1269,In_1188,In_1379);
and U1270 (N_1270,In_329,In_157);
xnor U1271 (N_1271,In_1362,In_1724);
or U1272 (N_1272,In_467,In_803);
nand U1273 (N_1273,In_1718,In_1470);
nor U1274 (N_1274,In_22,In_318);
xnor U1275 (N_1275,In_7,In_1607);
or U1276 (N_1276,In_700,In_735);
nor U1277 (N_1277,In_1913,In_802);
nand U1278 (N_1278,In_1351,In_98);
nand U1279 (N_1279,In_1085,In_144);
or U1280 (N_1280,In_1518,In_1371);
or U1281 (N_1281,In_505,In_1946);
xor U1282 (N_1282,In_1605,In_244);
nor U1283 (N_1283,In_340,In_404);
and U1284 (N_1284,In_1021,In_714);
or U1285 (N_1285,In_1306,In_1212);
nand U1286 (N_1286,In_102,In_234);
or U1287 (N_1287,In_1893,In_572);
nor U1288 (N_1288,In_446,In_1197);
nor U1289 (N_1289,In_977,In_509);
nor U1290 (N_1290,In_804,In_1508);
or U1291 (N_1291,In_647,In_1781);
nor U1292 (N_1292,In_1877,In_203);
and U1293 (N_1293,In_257,In_267);
xor U1294 (N_1294,In_117,In_172);
or U1295 (N_1295,In_1553,In_1238);
xnor U1296 (N_1296,In_1129,In_1312);
nand U1297 (N_1297,In_376,In_1556);
nand U1298 (N_1298,In_1221,In_786);
or U1299 (N_1299,In_1089,In_796);
xor U1300 (N_1300,In_1680,In_273);
nor U1301 (N_1301,In_301,In_906);
or U1302 (N_1302,In_1505,In_1913);
xnor U1303 (N_1303,In_307,In_1748);
nor U1304 (N_1304,In_1608,In_222);
or U1305 (N_1305,In_914,In_1787);
nand U1306 (N_1306,In_1801,In_1558);
xnor U1307 (N_1307,In_288,In_1149);
xnor U1308 (N_1308,In_1283,In_427);
xor U1309 (N_1309,In_1296,In_126);
nor U1310 (N_1310,In_148,In_952);
nor U1311 (N_1311,In_300,In_1765);
xor U1312 (N_1312,In_576,In_524);
or U1313 (N_1313,In_1490,In_1821);
nor U1314 (N_1314,In_1546,In_1019);
nor U1315 (N_1315,In_435,In_1570);
or U1316 (N_1316,In_1306,In_1497);
xor U1317 (N_1317,In_1762,In_1443);
nor U1318 (N_1318,In_985,In_1793);
nor U1319 (N_1319,In_430,In_1481);
and U1320 (N_1320,In_704,In_889);
and U1321 (N_1321,In_1654,In_596);
nand U1322 (N_1322,In_1425,In_1043);
xor U1323 (N_1323,In_127,In_1659);
and U1324 (N_1324,In_399,In_1264);
nor U1325 (N_1325,In_1506,In_1007);
nor U1326 (N_1326,In_1339,In_62);
and U1327 (N_1327,In_62,In_574);
and U1328 (N_1328,In_1957,In_449);
nor U1329 (N_1329,In_1179,In_1691);
nand U1330 (N_1330,In_17,In_515);
or U1331 (N_1331,In_527,In_979);
and U1332 (N_1332,In_1691,In_794);
xor U1333 (N_1333,In_1093,In_946);
nor U1334 (N_1334,In_1824,In_239);
and U1335 (N_1335,In_21,In_71);
and U1336 (N_1336,In_1320,In_1470);
or U1337 (N_1337,In_956,In_1971);
xnor U1338 (N_1338,In_661,In_1192);
nor U1339 (N_1339,In_629,In_128);
xnor U1340 (N_1340,In_1338,In_1748);
or U1341 (N_1341,In_969,In_885);
xor U1342 (N_1342,In_1381,In_1063);
xnor U1343 (N_1343,In_1034,In_346);
nand U1344 (N_1344,In_1446,In_1955);
nand U1345 (N_1345,In_741,In_1452);
nor U1346 (N_1346,In_617,In_1377);
nand U1347 (N_1347,In_749,In_185);
nor U1348 (N_1348,In_1658,In_1305);
xor U1349 (N_1349,In_1557,In_729);
or U1350 (N_1350,In_422,In_1365);
nand U1351 (N_1351,In_1681,In_497);
nand U1352 (N_1352,In_1150,In_1718);
nor U1353 (N_1353,In_1162,In_597);
or U1354 (N_1354,In_1780,In_439);
or U1355 (N_1355,In_1563,In_1921);
nor U1356 (N_1356,In_1356,In_1690);
nor U1357 (N_1357,In_509,In_274);
nor U1358 (N_1358,In_145,In_241);
xnor U1359 (N_1359,In_868,In_443);
and U1360 (N_1360,In_1166,In_1574);
nor U1361 (N_1361,In_1152,In_180);
xor U1362 (N_1362,In_627,In_645);
nor U1363 (N_1363,In_1200,In_1020);
xor U1364 (N_1364,In_1433,In_30);
and U1365 (N_1365,In_1404,In_21);
and U1366 (N_1366,In_1393,In_758);
xnor U1367 (N_1367,In_167,In_294);
nand U1368 (N_1368,In_1757,In_1811);
nand U1369 (N_1369,In_864,In_443);
or U1370 (N_1370,In_1023,In_1054);
nand U1371 (N_1371,In_946,In_824);
and U1372 (N_1372,In_1186,In_754);
nand U1373 (N_1373,In_652,In_946);
nor U1374 (N_1374,In_239,In_1185);
and U1375 (N_1375,In_1794,In_1063);
nand U1376 (N_1376,In_1107,In_31);
xor U1377 (N_1377,In_1938,In_1540);
xor U1378 (N_1378,In_905,In_398);
nor U1379 (N_1379,In_1189,In_1971);
nor U1380 (N_1380,In_522,In_169);
or U1381 (N_1381,In_488,In_124);
nand U1382 (N_1382,In_1560,In_706);
nand U1383 (N_1383,In_13,In_1888);
nand U1384 (N_1384,In_1901,In_1912);
xnor U1385 (N_1385,In_141,In_569);
xnor U1386 (N_1386,In_1705,In_1448);
nor U1387 (N_1387,In_1865,In_968);
nor U1388 (N_1388,In_92,In_1530);
nand U1389 (N_1389,In_255,In_31);
nor U1390 (N_1390,In_338,In_1461);
and U1391 (N_1391,In_199,In_1069);
and U1392 (N_1392,In_1355,In_125);
nor U1393 (N_1393,In_241,In_1848);
and U1394 (N_1394,In_1630,In_256);
and U1395 (N_1395,In_387,In_182);
and U1396 (N_1396,In_408,In_1640);
or U1397 (N_1397,In_1067,In_1747);
or U1398 (N_1398,In_368,In_1827);
nand U1399 (N_1399,In_544,In_1252);
nand U1400 (N_1400,In_1812,In_240);
nand U1401 (N_1401,In_762,In_1128);
nor U1402 (N_1402,In_1549,In_916);
and U1403 (N_1403,In_255,In_40);
nand U1404 (N_1404,In_130,In_496);
xor U1405 (N_1405,In_176,In_1576);
nor U1406 (N_1406,In_531,In_571);
nor U1407 (N_1407,In_548,In_237);
nor U1408 (N_1408,In_1313,In_544);
nor U1409 (N_1409,In_1403,In_1179);
nand U1410 (N_1410,In_1513,In_1307);
nand U1411 (N_1411,In_1974,In_1575);
and U1412 (N_1412,In_680,In_1990);
nand U1413 (N_1413,In_1338,In_954);
nor U1414 (N_1414,In_1318,In_1772);
or U1415 (N_1415,In_1575,In_962);
nand U1416 (N_1416,In_1905,In_1740);
xor U1417 (N_1417,In_857,In_1948);
and U1418 (N_1418,In_325,In_427);
nor U1419 (N_1419,In_762,In_1240);
and U1420 (N_1420,In_783,In_915);
xor U1421 (N_1421,In_1084,In_1499);
nor U1422 (N_1422,In_1361,In_844);
nor U1423 (N_1423,In_23,In_1209);
nand U1424 (N_1424,In_1609,In_1303);
nand U1425 (N_1425,In_1476,In_728);
and U1426 (N_1426,In_592,In_798);
or U1427 (N_1427,In_1956,In_1389);
and U1428 (N_1428,In_72,In_187);
xor U1429 (N_1429,In_701,In_977);
xnor U1430 (N_1430,In_641,In_705);
and U1431 (N_1431,In_473,In_390);
nor U1432 (N_1432,In_420,In_766);
nor U1433 (N_1433,In_783,In_1584);
or U1434 (N_1434,In_680,In_325);
and U1435 (N_1435,In_582,In_1249);
nand U1436 (N_1436,In_105,In_613);
and U1437 (N_1437,In_1599,In_173);
nand U1438 (N_1438,In_507,In_154);
or U1439 (N_1439,In_213,In_1750);
and U1440 (N_1440,In_230,In_26);
and U1441 (N_1441,In_812,In_802);
and U1442 (N_1442,In_609,In_638);
nand U1443 (N_1443,In_907,In_885);
nand U1444 (N_1444,In_1538,In_211);
nor U1445 (N_1445,In_1780,In_1650);
and U1446 (N_1446,In_1065,In_66);
nand U1447 (N_1447,In_1439,In_800);
nand U1448 (N_1448,In_1571,In_865);
or U1449 (N_1449,In_382,In_1294);
nor U1450 (N_1450,In_1101,In_1409);
or U1451 (N_1451,In_1815,In_649);
xor U1452 (N_1452,In_1847,In_522);
xor U1453 (N_1453,In_245,In_479);
or U1454 (N_1454,In_169,In_4);
nor U1455 (N_1455,In_776,In_827);
nor U1456 (N_1456,In_1600,In_981);
xor U1457 (N_1457,In_298,In_1056);
and U1458 (N_1458,In_1431,In_1374);
nand U1459 (N_1459,In_1467,In_1299);
nor U1460 (N_1460,In_1511,In_17);
xor U1461 (N_1461,In_853,In_1097);
nand U1462 (N_1462,In_1900,In_1497);
and U1463 (N_1463,In_72,In_122);
nand U1464 (N_1464,In_1376,In_1029);
xor U1465 (N_1465,In_60,In_1361);
nand U1466 (N_1466,In_1575,In_1695);
and U1467 (N_1467,In_792,In_665);
and U1468 (N_1468,In_1630,In_412);
and U1469 (N_1469,In_1730,In_614);
xor U1470 (N_1470,In_20,In_1553);
and U1471 (N_1471,In_32,In_871);
xor U1472 (N_1472,In_771,In_633);
or U1473 (N_1473,In_1711,In_745);
and U1474 (N_1474,In_7,In_918);
nor U1475 (N_1475,In_1017,In_565);
and U1476 (N_1476,In_1294,In_1689);
nand U1477 (N_1477,In_386,In_730);
nor U1478 (N_1478,In_372,In_1065);
or U1479 (N_1479,In_299,In_145);
and U1480 (N_1480,In_67,In_1989);
xnor U1481 (N_1481,In_170,In_1617);
nand U1482 (N_1482,In_1699,In_525);
nand U1483 (N_1483,In_1531,In_1636);
nor U1484 (N_1484,In_287,In_397);
nor U1485 (N_1485,In_1284,In_1448);
or U1486 (N_1486,In_781,In_193);
xnor U1487 (N_1487,In_334,In_1530);
and U1488 (N_1488,In_1143,In_1896);
nand U1489 (N_1489,In_410,In_115);
xnor U1490 (N_1490,In_274,In_984);
or U1491 (N_1491,In_1879,In_608);
or U1492 (N_1492,In_1250,In_120);
xor U1493 (N_1493,In_710,In_674);
or U1494 (N_1494,In_1279,In_782);
nand U1495 (N_1495,In_1511,In_118);
nor U1496 (N_1496,In_154,In_188);
nor U1497 (N_1497,In_1728,In_1902);
and U1498 (N_1498,In_1067,In_1874);
nor U1499 (N_1499,In_991,In_1227);
or U1500 (N_1500,In_708,In_349);
and U1501 (N_1501,In_682,In_1543);
nand U1502 (N_1502,In_27,In_1376);
xor U1503 (N_1503,In_1617,In_1006);
nor U1504 (N_1504,In_749,In_1613);
nand U1505 (N_1505,In_1778,In_1790);
and U1506 (N_1506,In_14,In_1063);
nand U1507 (N_1507,In_406,In_1529);
xor U1508 (N_1508,In_1643,In_197);
and U1509 (N_1509,In_282,In_87);
or U1510 (N_1510,In_1662,In_290);
xor U1511 (N_1511,In_819,In_274);
nor U1512 (N_1512,In_1812,In_1524);
and U1513 (N_1513,In_1069,In_175);
nor U1514 (N_1514,In_750,In_962);
or U1515 (N_1515,In_269,In_706);
xnor U1516 (N_1516,In_945,In_881);
nand U1517 (N_1517,In_124,In_692);
or U1518 (N_1518,In_622,In_1960);
nand U1519 (N_1519,In_1936,In_1092);
xor U1520 (N_1520,In_1370,In_1418);
nand U1521 (N_1521,In_766,In_55);
or U1522 (N_1522,In_1112,In_1242);
or U1523 (N_1523,In_260,In_1105);
and U1524 (N_1524,In_1703,In_1253);
or U1525 (N_1525,In_1188,In_1392);
xnor U1526 (N_1526,In_5,In_1081);
nor U1527 (N_1527,In_67,In_1348);
and U1528 (N_1528,In_822,In_1472);
xor U1529 (N_1529,In_95,In_59);
and U1530 (N_1530,In_589,In_1042);
or U1531 (N_1531,In_1045,In_1201);
nand U1532 (N_1532,In_729,In_841);
nand U1533 (N_1533,In_1421,In_1782);
xor U1534 (N_1534,In_148,In_161);
nor U1535 (N_1535,In_1068,In_1358);
nand U1536 (N_1536,In_486,In_1276);
or U1537 (N_1537,In_324,In_907);
nor U1538 (N_1538,In_1115,In_1873);
or U1539 (N_1539,In_1396,In_609);
or U1540 (N_1540,In_1477,In_411);
or U1541 (N_1541,In_1721,In_981);
nand U1542 (N_1542,In_464,In_1167);
xor U1543 (N_1543,In_1796,In_1442);
nor U1544 (N_1544,In_678,In_1428);
nand U1545 (N_1545,In_1937,In_1559);
xnor U1546 (N_1546,In_1951,In_452);
xor U1547 (N_1547,In_343,In_1820);
xor U1548 (N_1548,In_470,In_272);
nor U1549 (N_1549,In_1384,In_1307);
or U1550 (N_1550,In_625,In_1502);
nand U1551 (N_1551,In_257,In_1333);
or U1552 (N_1552,In_991,In_369);
and U1553 (N_1553,In_87,In_965);
nor U1554 (N_1554,In_548,In_1618);
and U1555 (N_1555,In_1753,In_565);
nor U1556 (N_1556,In_280,In_1006);
xnor U1557 (N_1557,In_426,In_3);
or U1558 (N_1558,In_185,In_1917);
or U1559 (N_1559,In_802,In_1288);
nand U1560 (N_1560,In_130,In_1216);
xor U1561 (N_1561,In_1371,In_1607);
or U1562 (N_1562,In_236,In_672);
nor U1563 (N_1563,In_711,In_1193);
nand U1564 (N_1564,In_1966,In_85);
xor U1565 (N_1565,In_1658,In_686);
or U1566 (N_1566,In_623,In_1296);
xnor U1567 (N_1567,In_1733,In_210);
and U1568 (N_1568,In_526,In_1109);
and U1569 (N_1569,In_338,In_688);
nand U1570 (N_1570,In_790,In_1107);
nand U1571 (N_1571,In_40,In_270);
xor U1572 (N_1572,In_1772,In_1110);
or U1573 (N_1573,In_1146,In_1144);
nand U1574 (N_1574,In_918,In_485);
xnor U1575 (N_1575,In_346,In_827);
and U1576 (N_1576,In_1020,In_1189);
xnor U1577 (N_1577,In_239,In_741);
nor U1578 (N_1578,In_1766,In_587);
xor U1579 (N_1579,In_64,In_815);
nor U1580 (N_1580,In_361,In_1873);
xnor U1581 (N_1581,In_946,In_1170);
and U1582 (N_1582,In_1998,In_570);
or U1583 (N_1583,In_1747,In_1087);
and U1584 (N_1584,In_223,In_1991);
nand U1585 (N_1585,In_1693,In_559);
or U1586 (N_1586,In_417,In_893);
and U1587 (N_1587,In_935,In_1724);
nand U1588 (N_1588,In_1547,In_1653);
xor U1589 (N_1589,In_821,In_925);
or U1590 (N_1590,In_1140,In_833);
nand U1591 (N_1591,In_274,In_1599);
nor U1592 (N_1592,In_655,In_470);
nand U1593 (N_1593,In_239,In_1607);
nor U1594 (N_1594,In_1361,In_1478);
and U1595 (N_1595,In_167,In_863);
and U1596 (N_1596,In_1216,In_995);
nor U1597 (N_1597,In_1900,In_69);
nand U1598 (N_1598,In_1344,In_245);
nand U1599 (N_1599,In_677,In_834);
and U1600 (N_1600,In_1340,In_116);
or U1601 (N_1601,In_335,In_710);
nor U1602 (N_1602,In_746,In_510);
nand U1603 (N_1603,In_1317,In_787);
and U1604 (N_1604,In_1607,In_408);
xor U1605 (N_1605,In_213,In_283);
nand U1606 (N_1606,In_780,In_1888);
or U1607 (N_1607,In_38,In_1665);
and U1608 (N_1608,In_294,In_893);
nor U1609 (N_1609,In_1858,In_1394);
or U1610 (N_1610,In_691,In_200);
and U1611 (N_1611,In_1327,In_1358);
nor U1612 (N_1612,In_741,In_577);
xor U1613 (N_1613,In_1074,In_1833);
xnor U1614 (N_1614,In_1524,In_1941);
nand U1615 (N_1615,In_1946,In_17);
nand U1616 (N_1616,In_1008,In_1349);
nor U1617 (N_1617,In_1239,In_1214);
xor U1618 (N_1618,In_958,In_655);
or U1619 (N_1619,In_406,In_1402);
nand U1620 (N_1620,In_1379,In_679);
and U1621 (N_1621,In_482,In_810);
xor U1622 (N_1622,In_459,In_69);
xnor U1623 (N_1623,In_74,In_1617);
nor U1624 (N_1624,In_947,In_1194);
nand U1625 (N_1625,In_1224,In_1162);
nand U1626 (N_1626,In_533,In_1849);
nor U1627 (N_1627,In_998,In_414);
xor U1628 (N_1628,In_846,In_1769);
or U1629 (N_1629,In_713,In_1228);
nor U1630 (N_1630,In_565,In_1472);
xnor U1631 (N_1631,In_606,In_963);
or U1632 (N_1632,In_837,In_1230);
xor U1633 (N_1633,In_1252,In_929);
xnor U1634 (N_1634,In_295,In_1551);
and U1635 (N_1635,In_713,In_275);
xnor U1636 (N_1636,In_1961,In_801);
nor U1637 (N_1637,In_388,In_266);
nand U1638 (N_1638,In_1780,In_802);
nand U1639 (N_1639,In_1980,In_765);
xor U1640 (N_1640,In_264,In_1628);
or U1641 (N_1641,In_1060,In_1063);
nor U1642 (N_1642,In_472,In_1973);
nand U1643 (N_1643,In_52,In_1172);
nand U1644 (N_1644,In_920,In_1208);
or U1645 (N_1645,In_805,In_68);
and U1646 (N_1646,In_1584,In_1203);
xor U1647 (N_1647,In_1030,In_275);
nand U1648 (N_1648,In_133,In_1417);
nor U1649 (N_1649,In_1554,In_1781);
xor U1650 (N_1650,In_625,In_593);
nand U1651 (N_1651,In_195,In_70);
nand U1652 (N_1652,In_945,In_916);
nand U1653 (N_1653,In_744,In_501);
nor U1654 (N_1654,In_726,In_699);
or U1655 (N_1655,In_450,In_1818);
or U1656 (N_1656,In_332,In_1289);
nor U1657 (N_1657,In_1254,In_404);
nor U1658 (N_1658,In_424,In_1619);
xnor U1659 (N_1659,In_437,In_39);
or U1660 (N_1660,In_1952,In_769);
nand U1661 (N_1661,In_1845,In_585);
nor U1662 (N_1662,In_585,In_1869);
xor U1663 (N_1663,In_1077,In_1838);
and U1664 (N_1664,In_474,In_1694);
and U1665 (N_1665,In_954,In_1901);
nand U1666 (N_1666,In_1858,In_1165);
xnor U1667 (N_1667,In_602,In_1473);
and U1668 (N_1668,In_357,In_1423);
nor U1669 (N_1669,In_1771,In_966);
nand U1670 (N_1670,In_1359,In_358);
or U1671 (N_1671,In_343,In_737);
nor U1672 (N_1672,In_1779,In_1553);
nor U1673 (N_1673,In_707,In_1241);
or U1674 (N_1674,In_1809,In_1374);
xnor U1675 (N_1675,In_1976,In_714);
or U1676 (N_1676,In_448,In_1507);
nor U1677 (N_1677,In_500,In_325);
or U1678 (N_1678,In_776,In_987);
nand U1679 (N_1679,In_21,In_376);
or U1680 (N_1680,In_375,In_112);
or U1681 (N_1681,In_798,In_419);
nand U1682 (N_1682,In_472,In_1099);
or U1683 (N_1683,In_1566,In_1396);
nor U1684 (N_1684,In_348,In_1785);
nand U1685 (N_1685,In_100,In_914);
nor U1686 (N_1686,In_425,In_226);
and U1687 (N_1687,In_1226,In_49);
nor U1688 (N_1688,In_519,In_1917);
or U1689 (N_1689,In_1883,In_1855);
and U1690 (N_1690,In_1743,In_1644);
xnor U1691 (N_1691,In_806,In_561);
and U1692 (N_1692,In_1159,In_362);
and U1693 (N_1693,In_551,In_933);
nand U1694 (N_1694,In_1572,In_541);
and U1695 (N_1695,In_341,In_1090);
nor U1696 (N_1696,In_117,In_1530);
and U1697 (N_1697,In_1596,In_1126);
xnor U1698 (N_1698,In_1013,In_1249);
or U1699 (N_1699,In_1984,In_211);
nand U1700 (N_1700,In_1294,In_517);
nor U1701 (N_1701,In_1461,In_122);
nand U1702 (N_1702,In_1983,In_1598);
and U1703 (N_1703,In_1015,In_118);
nand U1704 (N_1704,In_1620,In_242);
or U1705 (N_1705,In_1298,In_1752);
or U1706 (N_1706,In_1936,In_1350);
and U1707 (N_1707,In_33,In_160);
nor U1708 (N_1708,In_1792,In_1775);
xor U1709 (N_1709,In_1514,In_1619);
nor U1710 (N_1710,In_618,In_965);
nand U1711 (N_1711,In_1156,In_1866);
nor U1712 (N_1712,In_1156,In_1759);
xor U1713 (N_1713,In_374,In_1722);
and U1714 (N_1714,In_912,In_1054);
and U1715 (N_1715,In_532,In_427);
nor U1716 (N_1716,In_140,In_1684);
nor U1717 (N_1717,In_85,In_1546);
xnor U1718 (N_1718,In_1747,In_440);
and U1719 (N_1719,In_469,In_1151);
nor U1720 (N_1720,In_1151,In_1966);
nand U1721 (N_1721,In_132,In_1351);
nor U1722 (N_1722,In_389,In_623);
nor U1723 (N_1723,In_167,In_671);
and U1724 (N_1724,In_907,In_280);
and U1725 (N_1725,In_287,In_1365);
and U1726 (N_1726,In_1816,In_122);
nor U1727 (N_1727,In_763,In_979);
or U1728 (N_1728,In_631,In_938);
and U1729 (N_1729,In_587,In_1203);
nor U1730 (N_1730,In_815,In_990);
nor U1731 (N_1731,In_980,In_385);
xnor U1732 (N_1732,In_1139,In_1684);
nor U1733 (N_1733,In_1830,In_630);
or U1734 (N_1734,In_827,In_1218);
xor U1735 (N_1735,In_1087,In_262);
and U1736 (N_1736,In_948,In_1718);
nor U1737 (N_1737,In_1124,In_746);
or U1738 (N_1738,In_1828,In_16);
and U1739 (N_1739,In_1925,In_993);
or U1740 (N_1740,In_106,In_1052);
nand U1741 (N_1741,In_200,In_190);
nor U1742 (N_1742,In_577,In_1562);
nor U1743 (N_1743,In_469,In_1347);
xnor U1744 (N_1744,In_302,In_483);
nor U1745 (N_1745,In_1629,In_1127);
xnor U1746 (N_1746,In_1526,In_1851);
and U1747 (N_1747,In_106,In_286);
nor U1748 (N_1748,In_739,In_744);
xor U1749 (N_1749,In_1665,In_1919);
or U1750 (N_1750,In_1887,In_885);
nor U1751 (N_1751,In_1674,In_196);
nand U1752 (N_1752,In_814,In_1482);
nand U1753 (N_1753,In_1719,In_1512);
or U1754 (N_1754,In_299,In_609);
nand U1755 (N_1755,In_1553,In_532);
and U1756 (N_1756,In_1522,In_1725);
xor U1757 (N_1757,In_1727,In_1538);
nand U1758 (N_1758,In_583,In_454);
nor U1759 (N_1759,In_1555,In_1153);
and U1760 (N_1760,In_38,In_1917);
xor U1761 (N_1761,In_785,In_918);
or U1762 (N_1762,In_1365,In_698);
and U1763 (N_1763,In_1106,In_1754);
nor U1764 (N_1764,In_1665,In_1047);
nand U1765 (N_1765,In_1438,In_1990);
nor U1766 (N_1766,In_1522,In_45);
nor U1767 (N_1767,In_1372,In_226);
nand U1768 (N_1768,In_1866,In_1678);
or U1769 (N_1769,In_257,In_199);
nor U1770 (N_1770,In_1200,In_72);
or U1771 (N_1771,In_920,In_1546);
or U1772 (N_1772,In_942,In_1189);
nor U1773 (N_1773,In_479,In_1186);
or U1774 (N_1774,In_1599,In_843);
nand U1775 (N_1775,In_847,In_1727);
nand U1776 (N_1776,In_1443,In_897);
and U1777 (N_1777,In_1740,In_843);
or U1778 (N_1778,In_252,In_1636);
or U1779 (N_1779,In_1120,In_1517);
nor U1780 (N_1780,In_1209,In_1833);
nand U1781 (N_1781,In_1024,In_1247);
or U1782 (N_1782,In_1613,In_105);
and U1783 (N_1783,In_366,In_1265);
xnor U1784 (N_1784,In_1781,In_1194);
and U1785 (N_1785,In_666,In_45);
or U1786 (N_1786,In_80,In_148);
xnor U1787 (N_1787,In_356,In_934);
xor U1788 (N_1788,In_473,In_1185);
xnor U1789 (N_1789,In_1267,In_1968);
nand U1790 (N_1790,In_1965,In_1758);
and U1791 (N_1791,In_1516,In_1859);
nand U1792 (N_1792,In_844,In_9);
and U1793 (N_1793,In_1191,In_951);
xnor U1794 (N_1794,In_1813,In_1455);
and U1795 (N_1795,In_1360,In_308);
and U1796 (N_1796,In_81,In_1850);
and U1797 (N_1797,In_809,In_440);
or U1798 (N_1798,In_559,In_1449);
nand U1799 (N_1799,In_211,In_1369);
nand U1800 (N_1800,In_1751,In_132);
and U1801 (N_1801,In_283,In_1588);
nor U1802 (N_1802,In_150,In_1193);
nor U1803 (N_1803,In_785,In_791);
or U1804 (N_1804,In_62,In_1961);
and U1805 (N_1805,In_503,In_1047);
or U1806 (N_1806,In_1784,In_1117);
and U1807 (N_1807,In_1548,In_1174);
nand U1808 (N_1808,In_134,In_322);
xor U1809 (N_1809,In_120,In_542);
xnor U1810 (N_1810,In_984,In_697);
and U1811 (N_1811,In_523,In_1311);
xor U1812 (N_1812,In_1747,In_1788);
and U1813 (N_1813,In_1558,In_123);
nor U1814 (N_1814,In_1416,In_1668);
and U1815 (N_1815,In_1421,In_89);
and U1816 (N_1816,In_771,In_265);
xor U1817 (N_1817,In_480,In_143);
nor U1818 (N_1818,In_1609,In_1976);
or U1819 (N_1819,In_31,In_1765);
or U1820 (N_1820,In_129,In_797);
or U1821 (N_1821,In_28,In_1010);
nor U1822 (N_1822,In_1178,In_1641);
nand U1823 (N_1823,In_881,In_1668);
or U1824 (N_1824,In_1136,In_1011);
xor U1825 (N_1825,In_1903,In_485);
and U1826 (N_1826,In_1870,In_1484);
and U1827 (N_1827,In_522,In_1675);
nand U1828 (N_1828,In_627,In_228);
nor U1829 (N_1829,In_1746,In_200);
and U1830 (N_1830,In_1197,In_1916);
xnor U1831 (N_1831,In_1090,In_485);
nor U1832 (N_1832,In_1468,In_909);
nand U1833 (N_1833,In_591,In_641);
and U1834 (N_1834,In_1017,In_506);
nand U1835 (N_1835,In_736,In_1119);
and U1836 (N_1836,In_1766,In_1610);
nand U1837 (N_1837,In_1006,In_67);
nand U1838 (N_1838,In_3,In_1023);
xnor U1839 (N_1839,In_1454,In_818);
nand U1840 (N_1840,In_904,In_653);
nor U1841 (N_1841,In_1362,In_820);
or U1842 (N_1842,In_1560,In_1060);
or U1843 (N_1843,In_1011,In_391);
nand U1844 (N_1844,In_367,In_530);
nand U1845 (N_1845,In_428,In_774);
nor U1846 (N_1846,In_1695,In_1245);
and U1847 (N_1847,In_1445,In_1180);
nand U1848 (N_1848,In_903,In_871);
nor U1849 (N_1849,In_427,In_1426);
nand U1850 (N_1850,In_1286,In_1520);
nand U1851 (N_1851,In_1850,In_1181);
nand U1852 (N_1852,In_20,In_340);
xnor U1853 (N_1853,In_1766,In_1294);
nor U1854 (N_1854,In_1011,In_1608);
nand U1855 (N_1855,In_504,In_15);
xnor U1856 (N_1856,In_905,In_275);
nand U1857 (N_1857,In_566,In_1014);
nand U1858 (N_1858,In_548,In_543);
nand U1859 (N_1859,In_548,In_929);
xnor U1860 (N_1860,In_1004,In_72);
or U1861 (N_1861,In_1271,In_1710);
nor U1862 (N_1862,In_571,In_1268);
and U1863 (N_1863,In_1481,In_1489);
xor U1864 (N_1864,In_1792,In_423);
xor U1865 (N_1865,In_1207,In_551);
nor U1866 (N_1866,In_503,In_1452);
and U1867 (N_1867,In_718,In_713);
and U1868 (N_1868,In_665,In_1347);
and U1869 (N_1869,In_1485,In_243);
and U1870 (N_1870,In_619,In_1795);
xnor U1871 (N_1871,In_1953,In_749);
nor U1872 (N_1872,In_925,In_467);
xnor U1873 (N_1873,In_1595,In_547);
and U1874 (N_1874,In_1150,In_97);
nand U1875 (N_1875,In_796,In_1356);
nor U1876 (N_1876,In_1879,In_1170);
or U1877 (N_1877,In_1843,In_1743);
and U1878 (N_1878,In_1811,In_1891);
nand U1879 (N_1879,In_1752,In_1537);
nand U1880 (N_1880,In_513,In_1894);
or U1881 (N_1881,In_1293,In_29);
and U1882 (N_1882,In_808,In_1661);
nand U1883 (N_1883,In_454,In_1101);
nor U1884 (N_1884,In_841,In_8);
nand U1885 (N_1885,In_1708,In_1969);
nor U1886 (N_1886,In_1595,In_638);
xor U1887 (N_1887,In_1740,In_1037);
nor U1888 (N_1888,In_1402,In_684);
nand U1889 (N_1889,In_1416,In_1986);
nor U1890 (N_1890,In_274,In_880);
and U1891 (N_1891,In_1187,In_125);
xor U1892 (N_1892,In_1593,In_836);
nand U1893 (N_1893,In_710,In_191);
xor U1894 (N_1894,In_1343,In_1996);
or U1895 (N_1895,In_855,In_298);
nand U1896 (N_1896,In_1940,In_187);
or U1897 (N_1897,In_1197,In_1954);
nor U1898 (N_1898,In_1916,In_1928);
xor U1899 (N_1899,In_1745,In_161);
nor U1900 (N_1900,In_1883,In_431);
nor U1901 (N_1901,In_567,In_33);
xnor U1902 (N_1902,In_1946,In_158);
nand U1903 (N_1903,In_346,In_1284);
xnor U1904 (N_1904,In_665,In_1530);
xor U1905 (N_1905,In_1339,In_1590);
or U1906 (N_1906,In_1152,In_1918);
and U1907 (N_1907,In_277,In_1553);
and U1908 (N_1908,In_821,In_1322);
xnor U1909 (N_1909,In_909,In_1704);
or U1910 (N_1910,In_1021,In_629);
and U1911 (N_1911,In_310,In_516);
nand U1912 (N_1912,In_390,In_185);
nand U1913 (N_1913,In_1632,In_1033);
or U1914 (N_1914,In_853,In_667);
nor U1915 (N_1915,In_1830,In_251);
or U1916 (N_1916,In_664,In_1373);
and U1917 (N_1917,In_795,In_1774);
and U1918 (N_1918,In_453,In_1055);
and U1919 (N_1919,In_1782,In_108);
or U1920 (N_1920,In_1311,In_419);
nand U1921 (N_1921,In_1808,In_87);
and U1922 (N_1922,In_1437,In_1253);
xor U1923 (N_1923,In_1692,In_1821);
xor U1924 (N_1924,In_492,In_86);
or U1925 (N_1925,In_424,In_532);
and U1926 (N_1926,In_1096,In_1561);
and U1927 (N_1927,In_1384,In_994);
and U1928 (N_1928,In_946,In_358);
nor U1929 (N_1929,In_1139,In_1262);
nand U1930 (N_1930,In_612,In_673);
and U1931 (N_1931,In_1517,In_1174);
xnor U1932 (N_1932,In_306,In_1985);
nor U1933 (N_1933,In_1478,In_1448);
xnor U1934 (N_1934,In_942,In_21);
nand U1935 (N_1935,In_265,In_955);
nor U1936 (N_1936,In_1326,In_1001);
nand U1937 (N_1937,In_1409,In_1498);
nand U1938 (N_1938,In_196,In_774);
nor U1939 (N_1939,In_803,In_1345);
and U1940 (N_1940,In_175,In_440);
nor U1941 (N_1941,In_973,In_1891);
or U1942 (N_1942,In_278,In_851);
or U1943 (N_1943,In_1404,In_460);
nand U1944 (N_1944,In_975,In_693);
nor U1945 (N_1945,In_655,In_574);
nand U1946 (N_1946,In_1511,In_1659);
or U1947 (N_1947,In_1166,In_1219);
nand U1948 (N_1948,In_626,In_1557);
or U1949 (N_1949,In_722,In_1578);
nor U1950 (N_1950,In_401,In_473);
nor U1951 (N_1951,In_1738,In_592);
nor U1952 (N_1952,In_1509,In_756);
nor U1953 (N_1953,In_524,In_1762);
and U1954 (N_1954,In_950,In_117);
or U1955 (N_1955,In_1208,In_1343);
and U1956 (N_1956,In_559,In_1197);
nand U1957 (N_1957,In_1645,In_1057);
xnor U1958 (N_1958,In_192,In_1120);
nor U1959 (N_1959,In_1598,In_582);
and U1960 (N_1960,In_1206,In_1529);
nand U1961 (N_1961,In_430,In_1011);
or U1962 (N_1962,In_830,In_1445);
nand U1963 (N_1963,In_704,In_1732);
xnor U1964 (N_1964,In_1125,In_281);
xnor U1965 (N_1965,In_109,In_401);
xnor U1966 (N_1966,In_159,In_1039);
or U1967 (N_1967,In_1461,In_456);
xor U1968 (N_1968,In_1555,In_1984);
or U1969 (N_1969,In_1932,In_85);
or U1970 (N_1970,In_1349,In_1375);
nand U1971 (N_1971,In_1556,In_810);
nor U1972 (N_1972,In_177,In_624);
and U1973 (N_1973,In_847,In_949);
or U1974 (N_1974,In_99,In_447);
nor U1975 (N_1975,In_1430,In_248);
xor U1976 (N_1976,In_1115,In_1215);
or U1977 (N_1977,In_841,In_162);
nand U1978 (N_1978,In_1909,In_1899);
and U1979 (N_1979,In_220,In_1017);
or U1980 (N_1980,In_1439,In_1706);
nor U1981 (N_1981,In_1173,In_1077);
nor U1982 (N_1982,In_213,In_189);
or U1983 (N_1983,In_1331,In_241);
and U1984 (N_1984,In_304,In_176);
nor U1985 (N_1985,In_1853,In_1472);
and U1986 (N_1986,In_880,In_658);
nor U1987 (N_1987,In_644,In_1711);
and U1988 (N_1988,In_613,In_666);
or U1989 (N_1989,In_553,In_215);
xor U1990 (N_1990,In_1418,In_649);
nor U1991 (N_1991,In_1803,In_382);
and U1992 (N_1992,In_767,In_1380);
and U1993 (N_1993,In_113,In_881);
nand U1994 (N_1994,In_321,In_885);
xnor U1995 (N_1995,In_1883,In_1919);
xor U1996 (N_1996,In_1024,In_1572);
nand U1997 (N_1997,In_457,In_74);
xnor U1998 (N_1998,In_434,In_1452);
nor U1999 (N_1999,In_1939,In_951);
nor U2000 (N_2000,In_347,In_1401);
or U2001 (N_2001,In_968,In_1443);
nor U2002 (N_2002,In_990,In_1406);
or U2003 (N_2003,In_420,In_727);
nand U2004 (N_2004,In_113,In_296);
or U2005 (N_2005,In_1847,In_708);
and U2006 (N_2006,In_1458,In_1156);
or U2007 (N_2007,In_733,In_416);
nor U2008 (N_2008,In_1821,In_1783);
xor U2009 (N_2009,In_1377,In_833);
nor U2010 (N_2010,In_103,In_779);
nand U2011 (N_2011,In_690,In_1291);
nand U2012 (N_2012,In_443,In_1403);
nor U2013 (N_2013,In_1036,In_867);
and U2014 (N_2014,In_1085,In_243);
xnor U2015 (N_2015,In_1300,In_1391);
nand U2016 (N_2016,In_672,In_49);
or U2017 (N_2017,In_1806,In_371);
xnor U2018 (N_2018,In_563,In_1381);
and U2019 (N_2019,In_125,In_1777);
nor U2020 (N_2020,In_1899,In_820);
or U2021 (N_2021,In_137,In_1969);
and U2022 (N_2022,In_1224,In_331);
and U2023 (N_2023,In_294,In_33);
nor U2024 (N_2024,In_208,In_830);
xor U2025 (N_2025,In_1766,In_840);
nand U2026 (N_2026,In_217,In_1668);
xnor U2027 (N_2027,In_57,In_193);
or U2028 (N_2028,In_292,In_531);
nor U2029 (N_2029,In_1365,In_1852);
and U2030 (N_2030,In_290,In_1509);
xnor U2031 (N_2031,In_681,In_1351);
nand U2032 (N_2032,In_1298,In_1866);
and U2033 (N_2033,In_1237,In_505);
nor U2034 (N_2034,In_1079,In_716);
nand U2035 (N_2035,In_1858,In_663);
and U2036 (N_2036,In_1110,In_887);
nand U2037 (N_2037,In_888,In_1712);
or U2038 (N_2038,In_599,In_528);
nand U2039 (N_2039,In_1460,In_879);
nor U2040 (N_2040,In_800,In_1989);
or U2041 (N_2041,In_641,In_596);
nor U2042 (N_2042,In_1407,In_927);
xnor U2043 (N_2043,In_707,In_1603);
or U2044 (N_2044,In_1653,In_251);
or U2045 (N_2045,In_1705,In_1900);
or U2046 (N_2046,In_243,In_1673);
or U2047 (N_2047,In_409,In_1684);
or U2048 (N_2048,In_1051,In_1763);
and U2049 (N_2049,In_136,In_732);
xnor U2050 (N_2050,In_820,In_1179);
or U2051 (N_2051,In_956,In_1707);
nand U2052 (N_2052,In_1911,In_389);
xor U2053 (N_2053,In_1457,In_814);
and U2054 (N_2054,In_1852,In_456);
nor U2055 (N_2055,In_1189,In_808);
nor U2056 (N_2056,In_1362,In_1025);
nor U2057 (N_2057,In_1193,In_813);
or U2058 (N_2058,In_262,In_729);
and U2059 (N_2059,In_122,In_1052);
nand U2060 (N_2060,In_187,In_1266);
nand U2061 (N_2061,In_550,In_1242);
xnor U2062 (N_2062,In_982,In_489);
and U2063 (N_2063,In_225,In_1325);
xnor U2064 (N_2064,In_878,In_1161);
nand U2065 (N_2065,In_813,In_1709);
nand U2066 (N_2066,In_377,In_844);
or U2067 (N_2067,In_1720,In_1850);
and U2068 (N_2068,In_350,In_732);
and U2069 (N_2069,In_1652,In_1765);
nand U2070 (N_2070,In_1790,In_1640);
or U2071 (N_2071,In_1355,In_508);
or U2072 (N_2072,In_1580,In_1668);
and U2073 (N_2073,In_619,In_1181);
nand U2074 (N_2074,In_677,In_1767);
nor U2075 (N_2075,In_1873,In_997);
and U2076 (N_2076,In_117,In_1680);
nor U2077 (N_2077,In_1285,In_557);
nand U2078 (N_2078,In_774,In_1367);
nand U2079 (N_2079,In_253,In_1781);
nor U2080 (N_2080,In_1901,In_679);
nor U2081 (N_2081,In_26,In_1993);
nor U2082 (N_2082,In_1922,In_1421);
nand U2083 (N_2083,In_1978,In_1445);
xor U2084 (N_2084,In_1301,In_1893);
and U2085 (N_2085,In_1411,In_52);
nor U2086 (N_2086,In_439,In_1196);
nor U2087 (N_2087,In_1108,In_100);
nand U2088 (N_2088,In_1982,In_225);
xor U2089 (N_2089,In_1523,In_1715);
xor U2090 (N_2090,In_698,In_1290);
and U2091 (N_2091,In_251,In_204);
nor U2092 (N_2092,In_317,In_403);
xnor U2093 (N_2093,In_1587,In_339);
nor U2094 (N_2094,In_1101,In_1836);
nor U2095 (N_2095,In_1078,In_927);
or U2096 (N_2096,In_602,In_1817);
xnor U2097 (N_2097,In_1101,In_1449);
nor U2098 (N_2098,In_1119,In_1599);
xor U2099 (N_2099,In_1779,In_665);
nor U2100 (N_2100,In_1894,In_1395);
xor U2101 (N_2101,In_519,In_939);
xor U2102 (N_2102,In_242,In_179);
and U2103 (N_2103,In_35,In_945);
and U2104 (N_2104,In_977,In_1227);
and U2105 (N_2105,In_1619,In_1401);
and U2106 (N_2106,In_1438,In_368);
or U2107 (N_2107,In_1573,In_97);
nor U2108 (N_2108,In_265,In_1021);
or U2109 (N_2109,In_1116,In_359);
nor U2110 (N_2110,In_203,In_1166);
nor U2111 (N_2111,In_1257,In_1192);
nor U2112 (N_2112,In_634,In_1883);
and U2113 (N_2113,In_1525,In_1973);
nand U2114 (N_2114,In_1111,In_174);
xnor U2115 (N_2115,In_1439,In_446);
and U2116 (N_2116,In_372,In_267);
or U2117 (N_2117,In_688,In_1106);
and U2118 (N_2118,In_1184,In_556);
nor U2119 (N_2119,In_1528,In_801);
xnor U2120 (N_2120,In_1186,In_1467);
nand U2121 (N_2121,In_477,In_1754);
nor U2122 (N_2122,In_1085,In_16);
nor U2123 (N_2123,In_825,In_1646);
or U2124 (N_2124,In_1516,In_1259);
nor U2125 (N_2125,In_1981,In_661);
nand U2126 (N_2126,In_307,In_1561);
and U2127 (N_2127,In_1216,In_385);
or U2128 (N_2128,In_1773,In_1836);
and U2129 (N_2129,In_1655,In_460);
or U2130 (N_2130,In_38,In_258);
xor U2131 (N_2131,In_672,In_724);
nand U2132 (N_2132,In_1509,In_467);
nand U2133 (N_2133,In_293,In_1500);
xor U2134 (N_2134,In_950,In_1887);
nand U2135 (N_2135,In_990,In_1245);
nor U2136 (N_2136,In_227,In_900);
nor U2137 (N_2137,In_1706,In_410);
xnor U2138 (N_2138,In_1950,In_967);
or U2139 (N_2139,In_613,In_939);
nand U2140 (N_2140,In_1110,In_1695);
or U2141 (N_2141,In_1377,In_1588);
or U2142 (N_2142,In_1267,In_50);
or U2143 (N_2143,In_322,In_297);
xnor U2144 (N_2144,In_227,In_1632);
and U2145 (N_2145,In_1745,In_1320);
nand U2146 (N_2146,In_1639,In_909);
xor U2147 (N_2147,In_126,In_33);
or U2148 (N_2148,In_324,In_572);
nand U2149 (N_2149,In_1834,In_925);
xor U2150 (N_2150,In_1371,In_452);
or U2151 (N_2151,In_1601,In_128);
or U2152 (N_2152,In_954,In_534);
and U2153 (N_2153,In_1254,In_68);
nor U2154 (N_2154,In_1251,In_413);
xnor U2155 (N_2155,In_1175,In_539);
or U2156 (N_2156,In_125,In_1551);
nor U2157 (N_2157,In_1447,In_647);
or U2158 (N_2158,In_329,In_290);
nand U2159 (N_2159,In_1649,In_387);
xnor U2160 (N_2160,In_919,In_1757);
nor U2161 (N_2161,In_1534,In_31);
nand U2162 (N_2162,In_688,In_151);
and U2163 (N_2163,In_1343,In_821);
and U2164 (N_2164,In_784,In_825);
and U2165 (N_2165,In_116,In_1065);
nor U2166 (N_2166,In_1014,In_35);
nand U2167 (N_2167,In_724,In_1825);
and U2168 (N_2168,In_1352,In_1390);
nor U2169 (N_2169,In_1468,In_417);
and U2170 (N_2170,In_1407,In_205);
nor U2171 (N_2171,In_208,In_1727);
nand U2172 (N_2172,In_676,In_385);
or U2173 (N_2173,In_1421,In_384);
nand U2174 (N_2174,In_541,In_1385);
and U2175 (N_2175,In_1,In_1934);
xnor U2176 (N_2176,In_1861,In_1029);
and U2177 (N_2177,In_624,In_1597);
nor U2178 (N_2178,In_548,In_678);
nand U2179 (N_2179,In_460,In_959);
and U2180 (N_2180,In_824,In_967);
nor U2181 (N_2181,In_1633,In_475);
xnor U2182 (N_2182,In_194,In_752);
or U2183 (N_2183,In_246,In_1824);
or U2184 (N_2184,In_21,In_1401);
or U2185 (N_2185,In_45,In_1580);
or U2186 (N_2186,In_1580,In_1669);
and U2187 (N_2187,In_935,In_1022);
or U2188 (N_2188,In_358,In_1736);
and U2189 (N_2189,In_211,In_1584);
or U2190 (N_2190,In_126,In_120);
nor U2191 (N_2191,In_1826,In_1781);
or U2192 (N_2192,In_409,In_1649);
xor U2193 (N_2193,In_465,In_1978);
nand U2194 (N_2194,In_803,In_616);
nand U2195 (N_2195,In_821,In_1259);
and U2196 (N_2196,In_31,In_790);
nor U2197 (N_2197,In_1759,In_201);
nor U2198 (N_2198,In_1094,In_1974);
xor U2199 (N_2199,In_1994,In_1626);
xnor U2200 (N_2200,In_1459,In_216);
and U2201 (N_2201,In_1329,In_935);
nor U2202 (N_2202,In_1713,In_1228);
nand U2203 (N_2203,In_1670,In_250);
or U2204 (N_2204,In_1794,In_11);
xor U2205 (N_2205,In_1567,In_304);
xnor U2206 (N_2206,In_517,In_2);
and U2207 (N_2207,In_1086,In_215);
nor U2208 (N_2208,In_1210,In_1030);
nor U2209 (N_2209,In_725,In_1936);
and U2210 (N_2210,In_1205,In_323);
or U2211 (N_2211,In_1930,In_584);
xnor U2212 (N_2212,In_1730,In_793);
and U2213 (N_2213,In_1349,In_1755);
nand U2214 (N_2214,In_295,In_769);
nor U2215 (N_2215,In_1362,In_1051);
nor U2216 (N_2216,In_745,In_491);
or U2217 (N_2217,In_508,In_269);
nand U2218 (N_2218,In_569,In_590);
or U2219 (N_2219,In_1950,In_786);
or U2220 (N_2220,In_1032,In_14);
nand U2221 (N_2221,In_1945,In_775);
nor U2222 (N_2222,In_48,In_1956);
nor U2223 (N_2223,In_1473,In_1038);
nand U2224 (N_2224,In_1264,In_702);
xor U2225 (N_2225,In_830,In_1968);
and U2226 (N_2226,In_1706,In_1030);
nand U2227 (N_2227,In_410,In_884);
or U2228 (N_2228,In_763,In_197);
nor U2229 (N_2229,In_1855,In_343);
xor U2230 (N_2230,In_1195,In_678);
and U2231 (N_2231,In_499,In_1884);
xnor U2232 (N_2232,In_1496,In_4);
nor U2233 (N_2233,In_1742,In_799);
nand U2234 (N_2234,In_1454,In_577);
xnor U2235 (N_2235,In_577,In_66);
and U2236 (N_2236,In_549,In_784);
or U2237 (N_2237,In_1827,In_1719);
nor U2238 (N_2238,In_145,In_549);
or U2239 (N_2239,In_341,In_1795);
nor U2240 (N_2240,In_258,In_377);
or U2241 (N_2241,In_1205,In_1953);
and U2242 (N_2242,In_423,In_276);
or U2243 (N_2243,In_126,In_1665);
or U2244 (N_2244,In_62,In_862);
or U2245 (N_2245,In_1458,In_191);
xnor U2246 (N_2246,In_1096,In_608);
xnor U2247 (N_2247,In_899,In_1515);
xnor U2248 (N_2248,In_1920,In_293);
and U2249 (N_2249,In_1216,In_1174);
nand U2250 (N_2250,In_1002,In_77);
xnor U2251 (N_2251,In_668,In_1803);
nand U2252 (N_2252,In_473,In_1231);
nor U2253 (N_2253,In_1292,In_993);
nor U2254 (N_2254,In_250,In_1934);
and U2255 (N_2255,In_525,In_164);
nand U2256 (N_2256,In_479,In_371);
and U2257 (N_2257,In_1509,In_1761);
xor U2258 (N_2258,In_1624,In_333);
or U2259 (N_2259,In_143,In_1383);
nor U2260 (N_2260,In_661,In_1649);
nor U2261 (N_2261,In_1673,In_589);
xnor U2262 (N_2262,In_322,In_854);
nor U2263 (N_2263,In_1975,In_443);
xor U2264 (N_2264,In_478,In_1068);
xor U2265 (N_2265,In_160,In_1948);
xnor U2266 (N_2266,In_535,In_1837);
or U2267 (N_2267,In_1378,In_633);
and U2268 (N_2268,In_646,In_1600);
nand U2269 (N_2269,In_826,In_1265);
or U2270 (N_2270,In_1295,In_162);
nor U2271 (N_2271,In_603,In_1563);
xnor U2272 (N_2272,In_420,In_1632);
or U2273 (N_2273,In_846,In_1369);
nor U2274 (N_2274,In_781,In_635);
and U2275 (N_2275,In_1585,In_42);
nor U2276 (N_2276,In_1594,In_1383);
nor U2277 (N_2277,In_89,In_1038);
or U2278 (N_2278,In_527,In_1141);
nand U2279 (N_2279,In_57,In_1705);
xor U2280 (N_2280,In_963,In_1518);
nand U2281 (N_2281,In_1396,In_1571);
xor U2282 (N_2282,In_681,In_1330);
nor U2283 (N_2283,In_1330,In_413);
or U2284 (N_2284,In_55,In_386);
xnor U2285 (N_2285,In_284,In_1037);
nor U2286 (N_2286,In_1271,In_1377);
or U2287 (N_2287,In_413,In_849);
xnor U2288 (N_2288,In_1691,In_1924);
nand U2289 (N_2289,In_454,In_457);
or U2290 (N_2290,In_1964,In_1956);
and U2291 (N_2291,In_516,In_1598);
or U2292 (N_2292,In_194,In_545);
or U2293 (N_2293,In_1970,In_1175);
nand U2294 (N_2294,In_1583,In_796);
and U2295 (N_2295,In_48,In_1105);
xor U2296 (N_2296,In_1056,In_1965);
xor U2297 (N_2297,In_391,In_332);
and U2298 (N_2298,In_1329,In_523);
and U2299 (N_2299,In_549,In_294);
nor U2300 (N_2300,In_1776,In_1942);
nor U2301 (N_2301,In_101,In_1541);
nand U2302 (N_2302,In_917,In_1614);
xor U2303 (N_2303,In_1349,In_491);
and U2304 (N_2304,In_1685,In_1654);
and U2305 (N_2305,In_49,In_536);
and U2306 (N_2306,In_1131,In_568);
and U2307 (N_2307,In_1197,In_1061);
nor U2308 (N_2308,In_1008,In_859);
or U2309 (N_2309,In_991,In_1219);
xnor U2310 (N_2310,In_1289,In_1531);
nor U2311 (N_2311,In_812,In_1163);
and U2312 (N_2312,In_935,In_1114);
or U2313 (N_2313,In_9,In_1067);
or U2314 (N_2314,In_1510,In_1716);
or U2315 (N_2315,In_707,In_153);
nand U2316 (N_2316,In_701,In_302);
and U2317 (N_2317,In_1593,In_369);
nand U2318 (N_2318,In_1122,In_1671);
or U2319 (N_2319,In_1329,In_1357);
nor U2320 (N_2320,In_1929,In_1487);
nor U2321 (N_2321,In_801,In_1267);
nor U2322 (N_2322,In_717,In_1247);
nand U2323 (N_2323,In_655,In_692);
nor U2324 (N_2324,In_512,In_1016);
nor U2325 (N_2325,In_181,In_454);
or U2326 (N_2326,In_978,In_990);
nand U2327 (N_2327,In_1743,In_501);
xnor U2328 (N_2328,In_909,In_1517);
xnor U2329 (N_2329,In_969,In_1315);
or U2330 (N_2330,In_1551,In_735);
nor U2331 (N_2331,In_1458,In_1348);
and U2332 (N_2332,In_1681,In_425);
and U2333 (N_2333,In_1405,In_1043);
nand U2334 (N_2334,In_240,In_1846);
and U2335 (N_2335,In_112,In_293);
xnor U2336 (N_2336,In_1208,In_379);
and U2337 (N_2337,In_1241,In_47);
nor U2338 (N_2338,In_546,In_1764);
nor U2339 (N_2339,In_969,In_1816);
or U2340 (N_2340,In_1054,In_1548);
nor U2341 (N_2341,In_1795,In_432);
nor U2342 (N_2342,In_1043,In_12);
or U2343 (N_2343,In_1655,In_1640);
nand U2344 (N_2344,In_1266,In_1333);
and U2345 (N_2345,In_1050,In_1758);
xnor U2346 (N_2346,In_994,In_1257);
nor U2347 (N_2347,In_325,In_1710);
nand U2348 (N_2348,In_741,In_198);
or U2349 (N_2349,In_1554,In_693);
and U2350 (N_2350,In_1712,In_592);
or U2351 (N_2351,In_833,In_1305);
xnor U2352 (N_2352,In_1926,In_24);
nor U2353 (N_2353,In_1012,In_1827);
and U2354 (N_2354,In_497,In_1880);
or U2355 (N_2355,In_624,In_909);
or U2356 (N_2356,In_1950,In_738);
nand U2357 (N_2357,In_948,In_234);
xnor U2358 (N_2358,In_808,In_478);
nand U2359 (N_2359,In_1191,In_403);
xnor U2360 (N_2360,In_423,In_989);
or U2361 (N_2361,In_1455,In_748);
nor U2362 (N_2362,In_1342,In_1539);
nand U2363 (N_2363,In_926,In_1639);
and U2364 (N_2364,In_1260,In_333);
xor U2365 (N_2365,In_1084,In_1691);
and U2366 (N_2366,In_1615,In_830);
nand U2367 (N_2367,In_671,In_1716);
xor U2368 (N_2368,In_341,In_892);
and U2369 (N_2369,In_1621,In_1081);
nand U2370 (N_2370,In_1347,In_1377);
and U2371 (N_2371,In_980,In_1893);
xor U2372 (N_2372,In_1031,In_82);
and U2373 (N_2373,In_1905,In_1463);
and U2374 (N_2374,In_1793,In_1101);
xor U2375 (N_2375,In_738,In_178);
xor U2376 (N_2376,In_1439,In_1324);
or U2377 (N_2377,In_303,In_989);
and U2378 (N_2378,In_673,In_1438);
and U2379 (N_2379,In_1406,In_314);
xnor U2380 (N_2380,In_1756,In_885);
xnor U2381 (N_2381,In_1004,In_1885);
or U2382 (N_2382,In_1664,In_1083);
and U2383 (N_2383,In_974,In_386);
nand U2384 (N_2384,In_25,In_530);
xnor U2385 (N_2385,In_274,In_1113);
and U2386 (N_2386,In_1528,In_991);
nor U2387 (N_2387,In_920,In_256);
nand U2388 (N_2388,In_70,In_147);
nand U2389 (N_2389,In_813,In_339);
or U2390 (N_2390,In_1546,In_674);
xnor U2391 (N_2391,In_3,In_168);
nor U2392 (N_2392,In_604,In_1382);
nand U2393 (N_2393,In_1794,In_945);
or U2394 (N_2394,In_455,In_1646);
or U2395 (N_2395,In_1916,In_1688);
nand U2396 (N_2396,In_1490,In_1747);
nand U2397 (N_2397,In_118,In_899);
or U2398 (N_2398,In_1618,In_1247);
xnor U2399 (N_2399,In_822,In_114);
and U2400 (N_2400,In_931,In_586);
nor U2401 (N_2401,In_951,In_953);
and U2402 (N_2402,In_1042,In_1314);
and U2403 (N_2403,In_660,In_566);
nor U2404 (N_2404,In_873,In_981);
xor U2405 (N_2405,In_344,In_821);
xnor U2406 (N_2406,In_605,In_719);
nand U2407 (N_2407,In_71,In_827);
nor U2408 (N_2408,In_1732,In_1113);
or U2409 (N_2409,In_729,In_1440);
xnor U2410 (N_2410,In_236,In_758);
nand U2411 (N_2411,In_778,In_1350);
and U2412 (N_2412,In_1665,In_1772);
nand U2413 (N_2413,In_1662,In_895);
xnor U2414 (N_2414,In_1223,In_1744);
and U2415 (N_2415,In_1672,In_589);
or U2416 (N_2416,In_1060,In_1859);
xnor U2417 (N_2417,In_348,In_1472);
nor U2418 (N_2418,In_1187,In_838);
nor U2419 (N_2419,In_314,In_213);
nand U2420 (N_2420,In_1229,In_1580);
nand U2421 (N_2421,In_1053,In_203);
nand U2422 (N_2422,In_964,In_207);
xor U2423 (N_2423,In_1076,In_1137);
and U2424 (N_2424,In_447,In_592);
and U2425 (N_2425,In_1700,In_99);
nor U2426 (N_2426,In_1938,In_736);
or U2427 (N_2427,In_1683,In_471);
nor U2428 (N_2428,In_1247,In_1088);
xor U2429 (N_2429,In_727,In_1276);
or U2430 (N_2430,In_1567,In_1662);
or U2431 (N_2431,In_489,In_1373);
nand U2432 (N_2432,In_1963,In_1782);
xor U2433 (N_2433,In_590,In_1589);
xnor U2434 (N_2434,In_1127,In_575);
xor U2435 (N_2435,In_955,In_1516);
nand U2436 (N_2436,In_1415,In_1736);
or U2437 (N_2437,In_1512,In_1849);
or U2438 (N_2438,In_1321,In_723);
xnor U2439 (N_2439,In_427,In_1185);
and U2440 (N_2440,In_1603,In_203);
and U2441 (N_2441,In_512,In_1191);
xor U2442 (N_2442,In_1394,In_1788);
nand U2443 (N_2443,In_1413,In_1184);
and U2444 (N_2444,In_1677,In_753);
and U2445 (N_2445,In_1404,In_393);
nand U2446 (N_2446,In_564,In_757);
xnor U2447 (N_2447,In_371,In_85);
nor U2448 (N_2448,In_400,In_1975);
and U2449 (N_2449,In_914,In_60);
nor U2450 (N_2450,In_234,In_596);
nor U2451 (N_2451,In_788,In_571);
xnor U2452 (N_2452,In_484,In_487);
nor U2453 (N_2453,In_1111,In_1012);
or U2454 (N_2454,In_278,In_1089);
nand U2455 (N_2455,In_1785,In_927);
and U2456 (N_2456,In_1973,In_471);
or U2457 (N_2457,In_1409,In_1376);
and U2458 (N_2458,In_905,In_860);
and U2459 (N_2459,In_529,In_1920);
or U2460 (N_2460,In_853,In_1279);
and U2461 (N_2461,In_544,In_1223);
or U2462 (N_2462,In_313,In_1169);
or U2463 (N_2463,In_1714,In_1689);
or U2464 (N_2464,In_1357,In_1762);
nand U2465 (N_2465,In_742,In_1276);
nor U2466 (N_2466,In_63,In_1939);
nand U2467 (N_2467,In_1998,In_1975);
and U2468 (N_2468,In_42,In_1637);
nor U2469 (N_2469,In_169,In_341);
nor U2470 (N_2470,In_1525,In_1455);
nand U2471 (N_2471,In_1901,In_1798);
nand U2472 (N_2472,In_1573,In_606);
and U2473 (N_2473,In_1328,In_979);
xor U2474 (N_2474,In_1819,In_839);
and U2475 (N_2475,In_299,In_1137);
xor U2476 (N_2476,In_227,In_855);
and U2477 (N_2477,In_591,In_1663);
and U2478 (N_2478,In_1330,In_1296);
nand U2479 (N_2479,In_1703,In_800);
nand U2480 (N_2480,In_1286,In_1249);
nor U2481 (N_2481,In_1269,In_1586);
and U2482 (N_2482,In_564,In_1378);
nand U2483 (N_2483,In_1318,In_1254);
or U2484 (N_2484,In_1494,In_1044);
and U2485 (N_2485,In_177,In_535);
and U2486 (N_2486,In_1492,In_1220);
nor U2487 (N_2487,In_1522,In_1375);
xnor U2488 (N_2488,In_166,In_410);
or U2489 (N_2489,In_187,In_1637);
nand U2490 (N_2490,In_219,In_631);
or U2491 (N_2491,In_1197,In_353);
and U2492 (N_2492,In_1568,In_1622);
xor U2493 (N_2493,In_1389,In_57);
or U2494 (N_2494,In_821,In_291);
and U2495 (N_2495,In_593,In_163);
or U2496 (N_2496,In_1107,In_874);
xnor U2497 (N_2497,In_1719,In_1757);
and U2498 (N_2498,In_521,In_788);
or U2499 (N_2499,In_1236,In_632);
xor U2500 (N_2500,In_396,In_1725);
nand U2501 (N_2501,In_555,In_769);
and U2502 (N_2502,In_814,In_1007);
nand U2503 (N_2503,In_977,In_515);
xnor U2504 (N_2504,In_495,In_1024);
nand U2505 (N_2505,In_518,In_1140);
xnor U2506 (N_2506,In_822,In_854);
nand U2507 (N_2507,In_1761,In_1459);
or U2508 (N_2508,In_1281,In_1051);
or U2509 (N_2509,In_226,In_48);
and U2510 (N_2510,In_117,In_699);
or U2511 (N_2511,In_378,In_469);
and U2512 (N_2512,In_1520,In_1483);
nand U2513 (N_2513,In_1819,In_72);
nor U2514 (N_2514,In_566,In_562);
and U2515 (N_2515,In_1249,In_489);
and U2516 (N_2516,In_164,In_1914);
nand U2517 (N_2517,In_1215,In_780);
nand U2518 (N_2518,In_861,In_714);
and U2519 (N_2519,In_813,In_1426);
nand U2520 (N_2520,In_98,In_918);
nand U2521 (N_2521,In_1745,In_1030);
nand U2522 (N_2522,In_638,In_1774);
and U2523 (N_2523,In_145,In_705);
nor U2524 (N_2524,In_1668,In_1465);
or U2525 (N_2525,In_668,In_1182);
and U2526 (N_2526,In_1257,In_1953);
nand U2527 (N_2527,In_603,In_1987);
or U2528 (N_2528,In_1284,In_204);
xor U2529 (N_2529,In_1024,In_215);
xor U2530 (N_2530,In_1509,In_1974);
or U2531 (N_2531,In_101,In_134);
nand U2532 (N_2532,In_282,In_1267);
xnor U2533 (N_2533,In_1343,In_1887);
or U2534 (N_2534,In_1877,In_370);
nand U2535 (N_2535,In_1342,In_1951);
and U2536 (N_2536,In_618,In_1845);
nor U2537 (N_2537,In_1868,In_321);
nor U2538 (N_2538,In_1343,In_573);
nor U2539 (N_2539,In_1187,In_210);
xnor U2540 (N_2540,In_988,In_1578);
nand U2541 (N_2541,In_456,In_679);
nand U2542 (N_2542,In_1194,In_1112);
nor U2543 (N_2543,In_412,In_363);
or U2544 (N_2544,In_224,In_1548);
or U2545 (N_2545,In_1738,In_1704);
nand U2546 (N_2546,In_1590,In_324);
nor U2547 (N_2547,In_1692,In_461);
nor U2548 (N_2548,In_1724,In_1647);
and U2549 (N_2549,In_1469,In_140);
and U2550 (N_2550,In_711,In_433);
nor U2551 (N_2551,In_1224,In_1972);
xor U2552 (N_2552,In_150,In_796);
nor U2553 (N_2553,In_464,In_1401);
or U2554 (N_2554,In_166,In_1145);
and U2555 (N_2555,In_778,In_1140);
nor U2556 (N_2556,In_1107,In_1900);
nor U2557 (N_2557,In_61,In_45);
and U2558 (N_2558,In_1513,In_771);
xnor U2559 (N_2559,In_349,In_126);
nor U2560 (N_2560,In_446,In_1865);
or U2561 (N_2561,In_941,In_72);
nand U2562 (N_2562,In_1788,In_679);
nand U2563 (N_2563,In_1104,In_43);
nor U2564 (N_2564,In_481,In_889);
or U2565 (N_2565,In_1480,In_1363);
and U2566 (N_2566,In_999,In_47);
xnor U2567 (N_2567,In_1981,In_1438);
xnor U2568 (N_2568,In_1275,In_1526);
nand U2569 (N_2569,In_1571,In_1788);
xnor U2570 (N_2570,In_594,In_1644);
xnor U2571 (N_2571,In_1668,In_1188);
and U2572 (N_2572,In_204,In_85);
or U2573 (N_2573,In_1740,In_1721);
nor U2574 (N_2574,In_1861,In_842);
nor U2575 (N_2575,In_820,In_1099);
or U2576 (N_2576,In_1834,In_1534);
nand U2577 (N_2577,In_507,In_330);
xor U2578 (N_2578,In_177,In_290);
nor U2579 (N_2579,In_1874,In_1040);
and U2580 (N_2580,In_196,In_1766);
nor U2581 (N_2581,In_112,In_1412);
and U2582 (N_2582,In_228,In_1416);
or U2583 (N_2583,In_1359,In_274);
or U2584 (N_2584,In_1058,In_54);
nor U2585 (N_2585,In_1842,In_596);
and U2586 (N_2586,In_369,In_1435);
nor U2587 (N_2587,In_29,In_1694);
or U2588 (N_2588,In_828,In_714);
and U2589 (N_2589,In_1717,In_1364);
nand U2590 (N_2590,In_1659,In_1209);
or U2591 (N_2591,In_677,In_181);
nor U2592 (N_2592,In_1637,In_1655);
nor U2593 (N_2593,In_1871,In_565);
nor U2594 (N_2594,In_1784,In_331);
xor U2595 (N_2595,In_90,In_663);
nor U2596 (N_2596,In_1403,In_1005);
or U2597 (N_2597,In_718,In_826);
or U2598 (N_2598,In_1806,In_813);
nor U2599 (N_2599,In_1989,In_1168);
or U2600 (N_2600,In_940,In_350);
and U2601 (N_2601,In_1586,In_525);
or U2602 (N_2602,In_774,In_1421);
or U2603 (N_2603,In_1144,In_1602);
or U2604 (N_2604,In_753,In_26);
nand U2605 (N_2605,In_1657,In_1807);
and U2606 (N_2606,In_1909,In_1847);
nor U2607 (N_2607,In_246,In_1234);
and U2608 (N_2608,In_110,In_1642);
nor U2609 (N_2609,In_1468,In_1980);
nand U2610 (N_2610,In_14,In_1296);
nor U2611 (N_2611,In_932,In_460);
nand U2612 (N_2612,In_1962,In_943);
nand U2613 (N_2613,In_1968,In_628);
nor U2614 (N_2614,In_1053,In_1275);
nor U2615 (N_2615,In_1459,In_795);
or U2616 (N_2616,In_1930,In_321);
or U2617 (N_2617,In_1210,In_1609);
and U2618 (N_2618,In_1097,In_34);
xor U2619 (N_2619,In_1330,In_85);
nor U2620 (N_2620,In_1594,In_1160);
or U2621 (N_2621,In_1022,In_372);
nand U2622 (N_2622,In_1514,In_1450);
and U2623 (N_2623,In_1518,In_308);
nand U2624 (N_2624,In_1323,In_1182);
nand U2625 (N_2625,In_298,In_1751);
nor U2626 (N_2626,In_1942,In_804);
nor U2627 (N_2627,In_335,In_1268);
xnor U2628 (N_2628,In_990,In_1619);
or U2629 (N_2629,In_1631,In_1859);
xor U2630 (N_2630,In_1608,In_562);
nor U2631 (N_2631,In_1494,In_559);
or U2632 (N_2632,In_733,In_700);
nor U2633 (N_2633,In_63,In_1020);
nand U2634 (N_2634,In_85,In_1463);
nand U2635 (N_2635,In_106,In_1172);
nor U2636 (N_2636,In_1856,In_514);
nand U2637 (N_2637,In_1558,In_6);
nand U2638 (N_2638,In_1123,In_1094);
or U2639 (N_2639,In_559,In_1175);
and U2640 (N_2640,In_166,In_1990);
or U2641 (N_2641,In_1982,In_1751);
xnor U2642 (N_2642,In_1665,In_198);
nand U2643 (N_2643,In_1565,In_1018);
nand U2644 (N_2644,In_1449,In_692);
nor U2645 (N_2645,In_290,In_420);
nor U2646 (N_2646,In_555,In_186);
xor U2647 (N_2647,In_334,In_940);
xor U2648 (N_2648,In_1457,In_1135);
xor U2649 (N_2649,In_416,In_1865);
nor U2650 (N_2650,In_142,In_1333);
and U2651 (N_2651,In_1281,In_726);
xor U2652 (N_2652,In_1395,In_233);
nor U2653 (N_2653,In_955,In_160);
nand U2654 (N_2654,In_1557,In_1058);
nand U2655 (N_2655,In_336,In_1575);
or U2656 (N_2656,In_1967,In_1187);
nor U2657 (N_2657,In_1588,In_1663);
xor U2658 (N_2658,In_1275,In_1097);
or U2659 (N_2659,In_1148,In_1942);
or U2660 (N_2660,In_1942,In_703);
xnor U2661 (N_2661,In_1953,In_1654);
xnor U2662 (N_2662,In_1297,In_1415);
nor U2663 (N_2663,In_1566,In_1717);
and U2664 (N_2664,In_1661,In_807);
and U2665 (N_2665,In_31,In_1834);
or U2666 (N_2666,In_536,In_1801);
and U2667 (N_2667,In_1707,In_382);
and U2668 (N_2668,In_1980,In_1593);
or U2669 (N_2669,In_225,In_1343);
and U2670 (N_2670,In_1977,In_803);
nand U2671 (N_2671,In_281,In_1005);
or U2672 (N_2672,In_704,In_142);
or U2673 (N_2673,In_1039,In_1274);
and U2674 (N_2674,In_1754,In_1433);
nand U2675 (N_2675,In_83,In_1911);
or U2676 (N_2676,In_554,In_38);
or U2677 (N_2677,In_246,In_293);
and U2678 (N_2678,In_1586,In_261);
nand U2679 (N_2679,In_1717,In_941);
and U2680 (N_2680,In_1834,In_1702);
nor U2681 (N_2681,In_1498,In_1249);
nand U2682 (N_2682,In_580,In_912);
or U2683 (N_2683,In_731,In_1045);
or U2684 (N_2684,In_822,In_1802);
and U2685 (N_2685,In_1364,In_1225);
nand U2686 (N_2686,In_14,In_652);
xnor U2687 (N_2687,In_1573,In_1374);
xor U2688 (N_2688,In_405,In_1732);
nand U2689 (N_2689,In_1345,In_1675);
and U2690 (N_2690,In_319,In_1552);
and U2691 (N_2691,In_801,In_1723);
xnor U2692 (N_2692,In_1825,In_240);
xor U2693 (N_2693,In_516,In_436);
and U2694 (N_2694,In_153,In_173);
and U2695 (N_2695,In_1464,In_1971);
and U2696 (N_2696,In_1033,In_1264);
or U2697 (N_2697,In_167,In_695);
xnor U2698 (N_2698,In_1926,In_1445);
and U2699 (N_2699,In_713,In_446);
nand U2700 (N_2700,In_1039,In_1377);
or U2701 (N_2701,In_105,In_572);
xnor U2702 (N_2702,In_16,In_1709);
nor U2703 (N_2703,In_495,In_1148);
and U2704 (N_2704,In_659,In_1055);
or U2705 (N_2705,In_1308,In_1419);
nor U2706 (N_2706,In_1536,In_1999);
nor U2707 (N_2707,In_1475,In_784);
nor U2708 (N_2708,In_456,In_431);
nand U2709 (N_2709,In_1994,In_556);
nor U2710 (N_2710,In_202,In_1826);
nand U2711 (N_2711,In_507,In_891);
and U2712 (N_2712,In_186,In_839);
nand U2713 (N_2713,In_1018,In_655);
nor U2714 (N_2714,In_1629,In_1974);
or U2715 (N_2715,In_312,In_1527);
nand U2716 (N_2716,In_1708,In_1358);
xor U2717 (N_2717,In_977,In_1710);
nand U2718 (N_2718,In_493,In_999);
nor U2719 (N_2719,In_602,In_616);
or U2720 (N_2720,In_823,In_1816);
or U2721 (N_2721,In_813,In_552);
and U2722 (N_2722,In_299,In_1217);
xnor U2723 (N_2723,In_65,In_1175);
nor U2724 (N_2724,In_1313,In_14);
or U2725 (N_2725,In_1943,In_1326);
nand U2726 (N_2726,In_1489,In_1106);
and U2727 (N_2727,In_139,In_779);
or U2728 (N_2728,In_713,In_971);
and U2729 (N_2729,In_1538,In_885);
or U2730 (N_2730,In_1894,In_1241);
or U2731 (N_2731,In_209,In_79);
nor U2732 (N_2732,In_39,In_1263);
nor U2733 (N_2733,In_1198,In_114);
xnor U2734 (N_2734,In_1313,In_1502);
nand U2735 (N_2735,In_1467,In_717);
nor U2736 (N_2736,In_15,In_838);
xor U2737 (N_2737,In_764,In_1439);
nand U2738 (N_2738,In_890,In_1482);
nand U2739 (N_2739,In_1444,In_560);
nor U2740 (N_2740,In_1656,In_1006);
nor U2741 (N_2741,In_491,In_286);
or U2742 (N_2742,In_848,In_434);
xor U2743 (N_2743,In_1674,In_1356);
and U2744 (N_2744,In_1572,In_1820);
xor U2745 (N_2745,In_1591,In_301);
xnor U2746 (N_2746,In_742,In_1627);
xnor U2747 (N_2747,In_640,In_562);
and U2748 (N_2748,In_1462,In_221);
nand U2749 (N_2749,In_911,In_1007);
nor U2750 (N_2750,In_1664,In_416);
or U2751 (N_2751,In_1486,In_226);
and U2752 (N_2752,In_1484,In_1568);
and U2753 (N_2753,In_500,In_1005);
and U2754 (N_2754,In_837,In_313);
or U2755 (N_2755,In_1029,In_760);
and U2756 (N_2756,In_1668,In_1878);
and U2757 (N_2757,In_1728,In_758);
nor U2758 (N_2758,In_844,In_1305);
nor U2759 (N_2759,In_735,In_1954);
xor U2760 (N_2760,In_62,In_1201);
or U2761 (N_2761,In_1044,In_536);
or U2762 (N_2762,In_1107,In_523);
and U2763 (N_2763,In_1239,In_1842);
nand U2764 (N_2764,In_225,In_314);
or U2765 (N_2765,In_143,In_615);
nand U2766 (N_2766,In_1633,In_1018);
nand U2767 (N_2767,In_776,In_1175);
nor U2768 (N_2768,In_671,In_940);
nand U2769 (N_2769,In_1215,In_1297);
nor U2770 (N_2770,In_1402,In_1405);
nand U2771 (N_2771,In_275,In_1773);
nor U2772 (N_2772,In_1939,In_628);
or U2773 (N_2773,In_536,In_393);
nand U2774 (N_2774,In_929,In_1826);
nor U2775 (N_2775,In_582,In_1295);
nand U2776 (N_2776,In_440,In_991);
or U2777 (N_2777,In_1020,In_185);
nand U2778 (N_2778,In_1320,In_829);
xnor U2779 (N_2779,In_1127,In_1186);
nor U2780 (N_2780,In_1509,In_316);
and U2781 (N_2781,In_1828,In_1358);
xor U2782 (N_2782,In_1260,In_1652);
or U2783 (N_2783,In_885,In_491);
and U2784 (N_2784,In_834,In_577);
or U2785 (N_2785,In_325,In_213);
xor U2786 (N_2786,In_771,In_1567);
nor U2787 (N_2787,In_1649,In_959);
nand U2788 (N_2788,In_934,In_1184);
xnor U2789 (N_2789,In_222,In_1751);
nor U2790 (N_2790,In_1858,In_178);
nor U2791 (N_2791,In_1581,In_497);
and U2792 (N_2792,In_317,In_310);
nor U2793 (N_2793,In_304,In_58);
or U2794 (N_2794,In_1456,In_1943);
nor U2795 (N_2795,In_1181,In_1083);
and U2796 (N_2796,In_1828,In_1468);
or U2797 (N_2797,In_1925,In_307);
xnor U2798 (N_2798,In_716,In_1944);
nor U2799 (N_2799,In_1395,In_1108);
or U2800 (N_2800,In_1900,In_1591);
nor U2801 (N_2801,In_1365,In_1517);
and U2802 (N_2802,In_365,In_1591);
nor U2803 (N_2803,In_1714,In_29);
or U2804 (N_2804,In_810,In_309);
nand U2805 (N_2805,In_1926,In_69);
xnor U2806 (N_2806,In_966,In_113);
nand U2807 (N_2807,In_884,In_22);
and U2808 (N_2808,In_1463,In_1162);
and U2809 (N_2809,In_1264,In_1098);
or U2810 (N_2810,In_1846,In_521);
and U2811 (N_2811,In_315,In_695);
xor U2812 (N_2812,In_1028,In_261);
and U2813 (N_2813,In_783,In_324);
xor U2814 (N_2814,In_1824,In_1139);
xnor U2815 (N_2815,In_1813,In_369);
xor U2816 (N_2816,In_526,In_1300);
and U2817 (N_2817,In_1875,In_1509);
nand U2818 (N_2818,In_780,In_493);
xor U2819 (N_2819,In_1124,In_1600);
and U2820 (N_2820,In_1798,In_1090);
and U2821 (N_2821,In_713,In_1483);
and U2822 (N_2822,In_1907,In_1594);
and U2823 (N_2823,In_1395,In_1353);
and U2824 (N_2824,In_721,In_672);
and U2825 (N_2825,In_58,In_1414);
or U2826 (N_2826,In_681,In_134);
nand U2827 (N_2827,In_566,In_827);
xor U2828 (N_2828,In_588,In_1921);
and U2829 (N_2829,In_619,In_1529);
xnor U2830 (N_2830,In_1286,In_254);
or U2831 (N_2831,In_1104,In_1192);
and U2832 (N_2832,In_349,In_1159);
or U2833 (N_2833,In_146,In_692);
nand U2834 (N_2834,In_861,In_1379);
nor U2835 (N_2835,In_1414,In_1393);
and U2836 (N_2836,In_69,In_18);
nand U2837 (N_2837,In_1982,In_82);
or U2838 (N_2838,In_1811,In_34);
nand U2839 (N_2839,In_428,In_1842);
and U2840 (N_2840,In_423,In_296);
nand U2841 (N_2841,In_1793,In_682);
xor U2842 (N_2842,In_1130,In_1401);
xor U2843 (N_2843,In_350,In_30);
xor U2844 (N_2844,In_941,In_1858);
nor U2845 (N_2845,In_430,In_1594);
or U2846 (N_2846,In_125,In_1991);
nor U2847 (N_2847,In_1969,In_1003);
nor U2848 (N_2848,In_973,In_1730);
and U2849 (N_2849,In_252,In_769);
or U2850 (N_2850,In_799,In_1908);
nand U2851 (N_2851,In_1166,In_304);
or U2852 (N_2852,In_299,In_1058);
nand U2853 (N_2853,In_1520,In_1058);
nand U2854 (N_2854,In_1932,In_877);
or U2855 (N_2855,In_170,In_921);
nand U2856 (N_2856,In_1111,In_117);
and U2857 (N_2857,In_1209,In_1363);
or U2858 (N_2858,In_898,In_1119);
nor U2859 (N_2859,In_2,In_77);
or U2860 (N_2860,In_1152,In_601);
nor U2861 (N_2861,In_1370,In_429);
or U2862 (N_2862,In_1478,In_453);
or U2863 (N_2863,In_1425,In_1212);
or U2864 (N_2864,In_792,In_435);
nor U2865 (N_2865,In_1569,In_908);
nand U2866 (N_2866,In_1048,In_1114);
nand U2867 (N_2867,In_544,In_1599);
and U2868 (N_2868,In_1093,In_136);
or U2869 (N_2869,In_1,In_278);
nand U2870 (N_2870,In_1431,In_771);
and U2871 (N_2871,In_963,In_664);
xor U2872 (N_2872,In_627,In_437);
xnor U2873 (N_2873,In_1667,In_454);
xnor U2874 (N_2874,In_130,In_1772);
xnor U2875 (N_2875,In_924,In_1782);
xnor U2876 (N_2876,In_1939,In_274);
or U2877 (N_2877,In_247,In_950);
or U2878 (N_2878,In_477,In_1435);
xor U2879 (N_2879,In_1865,In_1762);
xor U2880 (N_2880,In_1198,In_212);
and U2881 (N_2881,In_79,In_1702);
nand U2882 (N_2882,In_1483,In_1090);
nor U2883 (N_2883,In_110,In_1318);
xor U2884 (N_2884,In_115,In_949);
nand U2885 (N_2885,In_1367,In_1845);
or U2886 (N_2886,In_573,In_1249);
nor U2887 (N_2887,In_425,In_279);
and U2888 (N_2888,In_247,In_762);
or U2889 (N_2889,In_1759,In_99);
xor U2890 (N_2890,In_1022,In_747);
or U2891 (N_2891,In_1169,In_902);
and U2892 (N_2892,In_1007,In_925);
nor U2893 (N_2893,In_1037,In_1818);
nor U2894 (N_2894,In_1112,In_1776);
xor U2895 (N_2895,In_1354,In_1092);
or U2896 (N_2896,In_218,In_343);
and U2897 (N_2897,In_1618,In_1468);
xnor U2898 (N_2898,In_29,In_176);
nor U2899 (N_2899,In_552,In_418);
nor U2900 (N_2900,In_222,In_882);
nor U2901 (N_2901,In_315,In_1980);
or U2902 (N_2902,In_591,In_798);
nor U2903 (N_2903,In_1109,In_1060);
or U2904 (N_2904,In_351,In_377);
nor U2905 (N_2905,In_324,In_440);
and U2906 (N_2906,In_1129,In_979);
and U2907 (N_2907,In_289,In_450);
xor U2908 (N_2908,In_888,In_1433);
xor U2909 (N_2909,In_656,In_210);
xnor U2910 (N_2910,In_494,In_1461);
xnor U2911 (N_2911,In_1783,In_415);
and U2912 (N_2912,In_1263,In_644);
or U2913 (N_2913,In_1868,In_1007);
or U2914 (N_2914,In_516,In_1208);
xnor U2915 (N_2915,In_396,In_1993);
xnor U2916 (N_2916,In_875,In_1120);
nand U2917 (N_2917,In_460,In_1675);
or U2918 (N_2918,In_1501,In_201);
or U2919 (N_2919,In_1516,In_1024);
or U2920 (N_2920,In_1790,In_1872);
and U2921 (N_2921,In_71,In_1261);
nor U2922 (N_2922,In_214,In_503);
or U2923 (N_2923,In_1019,In_1933);
or U2924 (N_2924,In_743,In_1114);
nor U2925 (N_2925,In_1313,In_1487);
xnor U2926 (N_2926,In_196,In_1465);
and U2927 (N_2927,In_1777,In_112);
nor U2928 (N_2928,In_492,In_251);
nor U2929 (N_2929,In_1147,In_1569);
and U2930 (N_2930,In_1000,In_971);
nor U2931 (N_2931,In_1967,In_1477);
xor U2932 (N_2932,In_1434,In_54);
and U2933 (N_2933,In_1672,In_1758);
nand U2934 (N_2934,In_810,In_1804);
nand U2935 (N_2935,In_340,In_1045);
and U2936 (N_2936,In_308,In_1956);
nor U2937 (N_2937,In_455,In_118);
or U2938 (N_2938,In_426,In_1437);
nand U2939 (N_2939,In_553,In_1934);
nand U2940 (N_2940,In_370,In_245);
or U2941 (N_2941,In_1078,In_761);
and U2942 (N_2942,In_1597,In_702);
nor U2943 (N_2943,In_1106,In_607);
xnor U2944 (N_2944,In_988,In_643);
nand U2945 (N_2945,In_70,In_291);
xnor U2946 (N_2946,In_1556,In_695);
xnor U2947 (N_2947,In_1304,In_768);
or U2948 (N_2948,In_799,In_1014);
or U2949 (N_2949,In_1480,In_1724);
xnor U2950 (N_2950,In_1635,In_1897);
and U2951 (N_2951,In_1161,In_1025);
nor U2952 (N_2952,In_232,In_1558);
nand U2953 (N_2953,In_1065,In_193);
xor U2954 (N_2954,In_554,In_264);
or U2955 (N_2955,In_1093,In_826);
or U2956 (N_2956,In_1326,In_1638);
and U2957 (N_2957,In_1676,In_1687);
nor U2958 (N_2958,In_1415,In_1429);
nor U2959 (N_2959,In_1979,In_1537);
nor U2960 (N_2960,In_142,In_1289);
xor U2961 (N_2961,In_1570,In_821);
nor U2962 (N_2962,In_1317,In_933);
and U2963 (N_2963,In_401,In_779);
or U2964 (N_2964,In_1348,In_155);
and U2965 (N_2965,In_993,In_288);
nand U2966 (N_2966,In_1529,In_547);
or U2967 (N_2967,In_1791,In_349);
nand U2968 (N_2968,In_1035,In_1033);
and U2969 (N_2969,In_164,In_1361);
nor U2970 (N_2970,In_552,In_1590);
and U2971 (N_2971,In_458,In_1325);
and U2972 (N_2972,In_1255,In_932);
and U2973 (N_2973,In_1890,In_803);
and U2974 (N_2974,In_137,In_1578);
nand U2975 (N_2975,In_1756,In_75);
or U2976 (N_2976,In_1354,In_173);
xnor U2977 (N_2977,In_888,In_1983);
nor U2978 (N_2978,In_791,In_1910);
or U2979 (N_2979,In_1808,In_1446);
and U2980 (N_2980,In_931,In_964);
xnor U2981 (N_2981,In_292,In_437);
xnor U2982 (N_2982,In_1843,In_1919);
or U2983 (N_2983,In_1109,In_833);
nand U2984 (N_2984,In_1127,In_1581);
nand U2985 (N_2985,In_258,In_1);
and U2986 (N_2986,In_1289,In_471);
xnor U2987 (N_2987,In_169,In_260);
nor U2988 (N_2988,In_1645,In_1838);
and U2989 (N_2989,In_456,In_648);
nor U2990 (N_2990,In_1593,In_2);
and U2991 (N_2991,In_459,In_1899);
xnor U2992 (N_2992,In_1592,In_1935);
xnor U2993 (N_2993,In_1244,In_512);
or U2994 (N_2994,In_473,In_1923);
xor U2995 (N_2995,In_660,In_719);
xor U2996 (N_2996,In_1855,In_811);
nor U2997 (N_2997,In_226,In_1681);
and U2998 (N_2998,In_173,In_648);
and U2999 (N_2999,In_1802,In_1381);
and U3000 (N_3000,In_1475,In_844);
xnor U3001 (N_3001,In_967,In_1242);
nor U3002 (N_3002,In_420,In_125);
xor U3003 (N_3003,In_1112,In_1609);
xnor U3004 (N_3004,In_335,In_1248);
and U3005 (N_3005,In_385,In_138);
or U3006 (N_3006,In_1188,In_815);
nand U3007 (N_3007,In_853,In_809);
nand U3008 (N_3008,In_1671,In_1068);
or U3009 (N_3009,In_772,In_9);
nand U3010 (N_3010,In_886,In_1850);
nor U3011 (N_3011,In_1489,In_425);
nor U3012 (N_3012,In_1763,In_1011);
and U3013 (N_3013,In_1669,In_331);
nor U3014 (N_3014,In_1161,In_153);
nor U3015 (N_3015,In_699,In_273);
xor U3016 (N_3016,In_1287,In_375);
nor U3017 (N_3017,In_564,In_1387);
or U3018 (N_3018,In_1259,In_1306);
xor U3019 (N_3019,In_831,In_1184);
xnor U3020 (N_3020,In_653,In_96);
nor U3021 (N_3021,In_1052,In_971);
nand U3022 (N_3022,In_1664,In_1670);
and U3023 (N_3023,In_235,In_115);
or U3024 (N_3024,In_393,In_277);
nand U3025 (N_3025,In_1315,In_541);
or U3026 (N_3026,In_563,In_483);
or U3027 (N_3027,In_1008,In_1408);
and U3028 (N_3028,In_969,In_138);
nor U3029 (N_3029,In_108,In_1392);
xor U3030 (N_3030,In_861,In_752);
nand U3031 (N_3031,In_1226,In_1885);
nand U3032 (N_3032,In_1727,In_981);
nand U3033 (N_3033,In_1306,In_1346);
xor U3034 (N_3034,In_651,In_1784);
and U3035 (N_3035,In_926,In_623);
nand U3036 (N_3036,In_1747,In_734);
nor U3037 (N_3037,In_419,In_1439);
nand U3038 (N_3038,In_558,In_705);
xor U3039 (N_3039,In_184,In_1306);
nand U3040 (N_3040,In_842,In_1119);
nand U3041 (N_3041,In_604,In_169);
or U3042 (N_3042,In_481,In_1671);
and U3043 (N_3043,In_404,In_1849);
and U3044 (N_3044,In_503,In_1180);
nand U3045 (N_3045,In_240,In_1476);
and U3046 (N_3046,In_584,In_1705);
or U3047 (N_3047,In_1960,In_1936);
and U3048 (N_3048,In_1762,In_167);
xnor U3049 (N_3049,In_988,In_1430);
nor U3050 (N_3050,In_1748,In_149);
xor U3051 (N_3051,In_1551,In_307);
and U3052 (N_3052,In_1808,In_650);
nand U3053 (N_3053,In_1920,In_1226);
or U3054 (N_3054,In_492,In_35);
xor U3055 (N_3055,In_1232,In_1854);
and U3056 (N_3056,In_1652,In_371);
and U3057 (N_3057,In_603,In_130);
nor U3058 (N_3058,In_86,In_489);
and U3059 (N_3059,In_640,In_1616);
and U3060 (N_3060,In_240,In_855);
and U3061 (N_3061,In_613,In_871);
and U3062 (N_3062,In_1503,In_35);
xor U3063 (N_3063,In_863,In_431);
and U3064 (N_3064,In_1885,In_1564);
and U3065 (N_3065,In_1917,In_483);
xor U3066 (N_3066,In_12,In_1262);
or U3067 (N_3067,In_1324,In_880);
and U3068 (N_3068,In_747,In_194);
nand U3069 (N_3069,In_1714,In_980);
nand U3070 (N_3070,In_1717,In_288);
nand U3071 (N_3071,In_93,In_637);
xnor U3072 (N_3072,In_1072,In_1315);
or U3073 (N_3073,In_1616,In_1129);
and U3074 (N_3074,In_160,In_1658);
xnor U3075 (N_3075,In_323,In_378);
nand U3076 (N_3076,In_55,In_1131);
xnor U3077 (N_3077,In_942,In_1489);
nor U3078 (N_3078,In_1801,In_971);
nor U3079 (N_3079,In_1754,In_530);
or U3080 (N_3080,In_599,In_122);
nand U3081 (N_3081,In_1990,In_1155);
xnor U3082 (N_3082,In_1700,In_1087);
nand U3083 (N_3083,In_1326,In_1075);
or U3084 (N_3084,In_1482,In_23);
xor U3085 (N_3085,In_1654,In_342);
xor U3086 (N_3086,In_954,In_1022);
or U3087 (N_3087,In_211,In_733);
xnor U3088 (N_3088,In_293,In_67);
nand U3089 (N_3089,In_1401,In_493);
and U3090 (N_3090,In_396,In_1033);
or U3091 (N_3091,In_739,In_514);
and U3092 (N_3092,In_59,In_354);
and U3093 (N_3093,In_1094,In_1957);
nor U3094 (N_3094,In_1209,In_141);
xnor U3095 (N_3095,In_180,In_479);
or U3096 (N_3096,In_1535,In_458);
xor U3097 (N_3097,In_1940,In_1007);
xnor U3098 (N_3098,In_527,In_638);
nor U3099 (N_3099,In_767,In_1687);
xnor U3100 (N_3100,In_285,In_1493);
or U3101 (N_3101,In_879,In_1555);
or U3102 (N_3102,In_1448,In_843);
nor U3103 (N_3103,In_1250,In_971);
xnor U3104 (N_3104,In_446,In_1510);
and U3105 (N_3105,In_522,In_99);
nor U3106 (N_3106,In_1258,In_639);
and U3107 (N_3107,In_225,In_1192);
nor U3108 (N_3108,In_1253,In_116);
xor U3109 (N_3109,In_924,In_1897);
or U3110 (N_3110,In_322,In_561);
xor U3111 (N_3111,In_1706,In_71);
nand U3112 (N_3112,In_548,In_1201);
and U3113 (N_3113,In_1324,In_1873);
nor U3114 (N_3114,In_91,In_266);
xor U3115 (N_3115,In_659,In_325);
nand U3116 (N_3116,In_893,In_934);
nand U3117 (N_3117,In_1979,In_728);
and U3118 (N_3118,In_1600,In_677);
or U3119 (N_3119,In_590,In_1828);
or U3120 (N_3120,In_1698,In_1825);
nand U3121 (N_3121,In_1357,In_965);
xor U3122 (N_3122,In_952,In_995);
nor U3123 (N_3123,In_359,In_514);
nand U3124 (N_3124,In_1574,In_1920);
nor U3125 (N_3125,In_783,In_1868);
xnor U3126 (N_3126,In_1357,In_804);
xnor U3127 (N_3127,In_1625,In_1352);
nand U3128 (N_3128,In_457,In_204);
or U3129 (N_3129,In_1557,In_394);
nor U3130 (N_3130,In_1233,In_1970);
nor U3131 (N_3131,In_1458,In_890);
and U3132 (N_3132,In_1416,In_1854);
or U3133 (N_3133,In_1205,In_1194);
nor U3134 (N_3134,In_1805,In_835);
and U3135 (N_3135,In_1137,In_1213);
and U3136 (N_3136,In_1157,In_1623);
nand U3137 (N_3137,In_286,In_1069);
and U3138 (N_3138,In_960,In_339);
nand U3139 (N_3139,In_184,In_1821);
and U3140 (N_3140,In_1323,In_557);
xnor U3141 (N_3141,In_393,In_1930);
or U3142 (N_3142,In_1638,In_777);
nand U3143 (N_3143,In_280,In_200);
nand U3144 (N_3144,In_245,In_1094);
or U3145 (N_3145,In_1666,In_542);
and U3146 (N_3146,In_1555,In_1702);
xor U3147 (N_3147,In_211,In_1267);
nor U3148 (N_3148,In_935,In_664);
nand U3149 (N_3149,In_1401,In_946);
nand U3150 (N_3150,In_376,In_1845);
nand U3151 (N_3151,In_1061,In_97);
or U3152 (N_3152,In_50,In_56);
nor U3153 (N_3153,In_1449,In_145);
or U3154 (N_3154,In_927,In_706);
or U3155 (N_3155,In_602,In_141);
nor U3156 (N_3156,In_438,In_1121);
nand U3157 (N_3157,In_1016,In_1175);
nand U3158 (N_3158,In_1870,In_837);
nor U3159 (N_3159,In_1000,In_1327);
or U3160 (N_3160,In_616,In_659);
nand U3161 (N_3161,In_567,In_796);
and U3162 (N_3162,In_1076,In_350);
and U3163 (N_3163,In_1083,In_945);
nor U3164 (N_3164,In_1528,In_1244);
or U3165 (N_3165,In_241,In_1533);
and U3166 (N_3166,In_231,In_640);
nor U3167 (N_3167,In_417,In_1108);
nor U3168 (N_3168,In_1828,In_1764);
or U3169 (N_3169,In_1906,In_1003);
or U3170 (N_3170,In_323,In_1983);
nor U3171 (N_3171,In_23,In_1702);
nand U3172 (N_3172,In_469,In_322);
xnor U3173 (N_3173,In_321,In_1984);
xor U3174 (N_3174,In_922,In_791);
xor U3175 (N_3175,In_570,In_1030);
and U3176 (N_3176,In_1865,In_873);
or U3177 (N_3177,In_1019,In_1271);
or U3178 (N_3178,In_92,In_413);
xnor U3179 (N_3179,In_1664,In_699);
nor U3180 (N_3180,In_1276,In_544);
nand U3181 (N_3181,In_1230,In_412);
xnor U3182 (N_3182,In_53,In_961);
or U3183 (N_3183,In_340,In_1714);
and U3184 (N_3184,In_598,In_695);
xor U3185 (N_3185,In_1245,In_1981);
or U3186 (N_3186,In_1708,In_88);
or U3187 (N_3187,In_456,In_1284);
nand U3188 (N_3188,In_267,In_1533);
nand U3189 (N_3189,In_1247,In_145);
nor U3190 (N_3190,In_1801,In_1421);
nor U3191 (N_3191,In_1222,In_1781);
nand U3192 (N_3192,In_1704,In_1993);
and U3193 (N_3193,In_1001,In_1728);
or U3194 (N_3194,In_713,In_949);
xor U3195 (N_3195,In_1964,In_839);
xor U3196 (N_3196,In_457,In_1250);
xor U3197 (N_3197,In_1785,In_637);
nand U3198 (N_3198,In_1598,In_765);
xor U3199 (N_3199,In_1484,In_1848);
or U3200 (N_3200,In_1985,In_1887);
or U3201 (N_3201,In_1503,In_46);
and U3202 (N_3202,In_140,In_1739);
or U3203 (N_3203,In_42,In_1413);
or U3204 (N_3204,In_265,In_1666);
or U3205 (N_3205,In_166,In_169);
nor U3206 (N_3206,In_1718,In_366);
nand U3207 (N_3207,In_59,In_1338);
or U3208 (N_3208,In_998,In_758);
and U3209 (N_3209,In_1912,In_825);
or U3210 (N_3210,In_1093,In_281);
and U3211 (N_3211,In_1699,In_1942);
nand U3212 (N_3212,In_877,In_1678);
nand U3213 (N_3213,In_137,In_66);
xor U3214 (N_3214,In_984,In_1717);
or U3215 (N_3215,In_539,In_1430);
xnor U3216 (N_3216,In_1256,In_1280);
xnor U3217 (N_3217,In_473,In_670);
nand U3218 (N_3218,In_797,In_1671);
nor U3219 (N_3219,In_1881,In_1493);
and U3220 (N_3220,In_1711,In_1170);
nor U3221 (N_3221,In_402,In_1924);
xnor U3222 (N_3222,In_1619,In_1578);
xor U3223 (N_3223,In_1259,In_822);
xor U3224 (N_3224,In_403,In_1117);
nor U3225 (N_3225,In_1005,In_1811);
xnor U3226 (N_3226,In_1954,In_1380);
nand U3227 (N_3227,In_639,In_1067);
xor U3228 (N_3228,In_1102,In_1156);
nor U3229 (N_3229,In_913,In_127);
nand U3230 (N_3230,In_1277,In_1544);
nor U3231 (N_3231,In_994,In_1132);
or U3232 (N_3232,In_18,In_736);
and U3233 (N_3233,In_1732,In_1742);
nand U3234 (N_3234,In_89,In_1439);
nand U3235 (N_3235,In_975,In_461);
and U3236 (N_3236,In_1518,In_1683);
nand U3237 (N_3237,In_1977,In_114);
and U3238 (N_3238,In_1908,In_121);
nor U3239 (N_3239,In_1838,In_394);
and U3240 (N_3240,In_1005,In_635);
xor U3241 (N_3241,In_1229,In_1769);
and U3242 (N_3242,In_1459,In_1938);
nand U3243 (N_3243,In_1561,In_312);
or U3244 (N_3244,In_1475,In_2);
nand U3245 (N_3245,In_189,In_1159);
xor U3246 (N_3246,In_1202,In_297);
xor U3247 (N_3247,In_1188,In_406);
or U3248 (N_3248,In_1276,In_236);
and U3249 (N_3249,In_1315,In_1716);
nand U3250 (N_3250,In_1429,In_1619);
nand U3251 (N_3251,In_633,In_81);
or U3252 (N_3252,In_265,In_1714);
or U3253 (N_3253,In_303,In_1649);
xor U3254 (N_3254,In_1311,In_697);
xor U3255 (N_3255,In_150,In_304);
nand U3256 (N_3256,In_1992,In_1091);
xor U3257 (N_3257,In_1833,In_363);
xor U3258 (N_3258,In_246,In_1027);
nor U3259 (N_3259,In_97,In_1601);
nand U3260 (N_3260,In_915,In_529);
or U3261 (N_3261,In_1686,In_255);
nor U3262 (N_3262,In_610,In_1067);
and U3263 (N_3263,In_877,In_695);
xor U3264 (N_3264,In_48,In_1566);
and U3265 (N_3265,In_125,In_1788);
xor U3266 (N_3266,In_1167,In_932);
or U3267 (N_3267,In_327,In_8);
and U3268 (N_3268,In_1622,In_1935);
nand U3269 (N_3269,In_222,In_347);
nand U3270 (N_3270,In_1582,In_13);
nand U3271 (N_3271,In_962,In_519);
or U3272 (N_3272,In_814,In_1648);
and U3273 (N_3273,In_77,In_1843);
xnor U3274 (N_3274,In_963,In_439);
xor U3275 (N_3275,In_283,In_1455);
nor U3276 (N_3276,In_1891,In_1399);
nand U3277 (N_3277,In_902,In_1165);
xor U3278 (N_3278,In_1987,In_292);
xor U3279 (N_3279,In_1838,In_1984);
nand U3280 (N_3280,In_561,In_1993);
xor U3281 (N_3281,In_1972,In_698);
xnor U3282 (N_3282,In_1718,In_1244);
nand U3283 (N_3283,In_610,In_186);
or U3284 (N_3284,In_1463,In_1965);
and U3285 (N_3285,In_1351,In_1061);
or U3286 (N_3286,In_753,In_808);
xnor U3287 (N_3287,In_791,In_1593);
nor U3288 (N_3288,In_1431,In_850);
nor U3289 (N_3289,In_1126,In_1350);
or U3290 (N_3290,In_690,In_401);
and U3291 (N_3291,In_1913,In_624);
nand U3292 (N_3292,In_1016,In_1110);
xor U3293 (N_3293,In_1367,In_1800);
or U3294 (N_3294,In_1985,In_571);
or U3295 (N_3295,In_1703,In_769);
nor U3296 (N_3296,In_1450,In_1902);
and U3297 (N_3297,In_747,In_1524);
and U3298 (N_3298,In_1746,In_929);
nand U3299 (N_3299,In_1206,In_1356);
nor U3300 (N_3300,In_610,In_1);
and U3301 (N_3301,In_1690,In_33);
nand U3302 (N_3302,In_888,In_1584);
nor U3303 (N_3303,In_1461,In_1665);
nor U3304 (N_3304,In_553,In_962);
xor U3305 (N_3305,In_1434,In_1846);
nand U3306 (N_3306,In_709,In_1595);
nand U3307 (N_3307,In_717,In_1352);
nor U3308 (N_3308,In_879,In_1715);
and U3309 (N_3309,In_1503,In_119);
nand U3310 (N_3310,In_295,In_641);
nand U3311 (N_3311,In_94,In_545);
nand U3312 (N_3312,In_1509,In_171);
nor U3313 (N_3313,In_1236,In_1962);
and U3314 (N_3314,In_310,In_1736);
nor U3315 (N_3315,In_393,In_926);
xor U3316 (N_3316,In_1198,In_966);
nor U3317 (N_3317,In_1974,In_818);
xor U3318 (N_3318,In_152,In_196);
or U3319 (N_3319,In_300,In_194);
xor U3320 (N_3320,In_242,In_1498);
nor U3321 (N_3321,In_1664,In_388);
nand U3322 (N_3322,In_1625,In_1351);
nor U3323 (N_3323,In_629,In_506);
nand U3324 (N_3324,In_844,In_1322);
xor U3325 (N_3325,In_1932,In_685);
xnor U3326 (N_3326,In_1437,In_1524);
and U3327 (N_3327,In_1065,In_204);
nand U3328 (N_3328,In_1363,In_142);
or U3329 (N_3329,In_449,In_1241);
or U3330 (N_3330,In_1880,In_1921);
or U3331 (N_3331,In_1821,In_295);
xor U3332 (N_3332,In_1337,In_1788);
and U3333 (N_3333,In_716,In_1477);
nand U3334 (N_3334,In_1220,In_1335);
xor U3335 (N_3335,In_1833,In_1308);
and U3336 (N_3336,In_992,In_798);
xor U3337 (N_3337,In_72,In_1072);
xnor U3338 (N_3338,In_1523,In_1976);
or U3339 (N_3339,In_1144,In_255);
and U3340 (N_3340,In_1952,In_1550);
or U3341 (N_3341,In_1521,In_877);
nand U3342 (N_3342,In_224,In_1063);
nand U3343 (N_3343,In_307,In_196);
nand U3344 (N_3344,In_1795,In_291);
nand U3345 (N_3345,In_1361,In_317);
nor U3346 (N_3346,In_1557,In_846);
xnor U3347 (N_3347,In_1543,In_756);
and U3348 (N_3348,In_996,In_282);
xor U3349 (N_3349,In_1648,In_504);
nand U3350 (N_3350,In_1878,In_541);
nor U3351 (N_3351,In_477,In_97);
xor U3352 (N_3352,In_564,In_552);
or U3353 (N_3353,In_107,In_874);
nor U3354 (N_3354,In_1760,In_235);
and U3355 (N_3355,In_1212,In_1405);
nand U3356 (N_3356,In_1330,In_534);
nand U3357 (N_3357,In_965,In_852);
nor U3358 (N_3358,In_1115,In_1514);
xor U3359 (N_3359,In_1947,In_1080);
or U3360 (N_3360,In_394,In_351);
or U3361 (N_3361,In_1976,In_831);
nor U3362 (N_3362,In_684,In_880);
nand U3363 (N_3363,In_1272,In_133);
nand U3364 (N_3364,In_205,In_91);
nand U3365 (N_3365,In_1257,In_701);
nor U3366 (N_3366,In_986,In_620);
xnor U3367 (N_3367,In_31,In_224);
or U3368 (N_3368,In_468,In_789);
xor U3369 (N_3369,In_196,In_68);
and U3370 (N_3370,In_1046,In_1788);
nor U3371 (N_3371,In_1795,In_30);
xnor U3372 (N_3372,In_1646,In_551);
xor U3373 (N_3373,In_1419,In_488);
xnor U3374 (N_3374,In_1723,In_1665);
and U3375 (N_3375,In_1152,In_962);
and U3376 (N_3376,In_1927,In_1333);
nor U3377 (N_3377,In_441,In_1557);
and U3378 (N_3378,In_1767,In_197);
and U3379 (N_3379,In_584,In_1786);
xnor U3380 (N_3380,In_589,In_1190);
and U3381 (N_3381,In_1370,In_331);
nand U3382 (N_3382,In_1271,In_452);
and U3383 (N_3383,In_337,In_1148);
xor U3384 (N_3384,In_660,In_827);
xor U3385 (N_3385,In_838,In_1333);
or U3386 (N_3386,In_490,In_907);
and U3387 (N_3387,In_292,In_1729);
or U3388 (N_3388,In_1262,In_352);
and U3389 (N_3389,In_1680,In_1707);
xor U3390 (N_3390,In_505,In_1737);
xnor U3391 (N_3391,In_89,In_1413);
and U3392 (N_3392,In_1484,In_1618);
nor U3393 (N_3393,In_994,In_892);
or U3394 (N_3394,In_1132,In_1019);
nand U3395 (N_3395,In_992,In_439);
nor U3396 (N_3396,In_749,In_711);
xor U3397 (N_3397,In_1853,In_1143);
or U3398 (N_3398,In_1177,In_1403);
nand U3399 (N_3399,In_1586,In_1918);
nor U3400 (N_3400,In_240,In_809);
nand U3401 (N_3401,In_1796,In_1275);
and U3402 (N_3402,In_309,In_807);
or U3403 (N_3403,In_26,In_1744);
xor U3404 (N_3404,In_1007,In_927);
nand U3405 (N_3405,In_1775,In_1109);
and U3406 (N_3406,In_497,In_1212);
nand U3407 (N_3407,In_1540,In_990);
or U3408 (N_3408,In_737,In_901);
nor U3409 (N_3409,In_1083,In_931);
or U3410 (N_3410,In_1126,In_175);
and U3411 (N_3411,In_363,In_1777);
or U3412 (N_3412,In_1909,In_1482);
nand U3413 (N_3413,In_400,In_270);
or U3414 (N_3414,In_1316,In_1352);
or U3415 (N_3415,In_489,In_1469);
xnor U3416 (N_3416,In_239,In_1789);
or U3417 (N_3417,In_308,In_1678);
or U3418 (N_3418,In_1442,In_614);
nor U3419 (N_3419,In_1348,In_1182);
nand U3420 (N_3420,In_1347,In_1234);
or U3421 (N_3421,In_1361,In_181);
nand U3422 (N_3422,In_683,In_5);
and U3423 (N_3423,In_1596,In_1676);
and U3424 (N_3424,In_394,In_27);
nor U3425 (N_3425,In_935,In_1227);
xnor U3426 (N_3426,In_595,In_1293);
or U3427 (N_3427,In_1514,In_805);
and U3428 (N_3428,In_1378,In_896);
xor U3429 (N_3429,In_560,In_441);
and U3430 (N_3430,In_891,In_578);
nand U3431 (N_3431,In_1508,In_1238);
and U3432 (N_3432,In_133,In_1438);
and U3433 (N_3433,In_205,In_1746);
nor U3434 (N_3434,In_1321,In_585);
nor U3435 (N_3435,In_519,In_1142);
and U3436 (N_3436,In_609,In_166);
xnor U3437 (N_3437,In_406,In_1130);
nand U3438 (N_3438,In_1434,In_512);
nor U3439 (N_3439,In_537,In_454);
nand U3440 (N_3440,In_1907,In_1936);
or U3441 (N_3441,In_1764,In_376);
nor U3442 (N_3442,In_1584,In_1780);
nand U3443 (N_3443,In_688,In_228);
nand U3444 (N_3444,In_345,In_1833);
nand U3445 (N_3445,In_169,In_1658);
or U3446 (N_3446,In_1406,In_709);
or U3447 (N_3447,In_1057,In_1549);
or U3448 (N_3448,In_660,In_1317);
nand U3449 (N_3449,In_649,In_301);
and U3450 (N_3450,In_671,In_326);
xor U3451 (N_3451,In_247,In_377);
and U3452 (N_3452,In_1455,In_584);
and U3453 (N_3453,In_843,In_485);
nand U3454 (N_3454,In_920,In_536);
xnor U3455 (N_3455,In_642,In_600);
and U3456 (N_3456,In_1716,In_249);
xnor U3457 (N_3457,In_1563,In_1604);
xnor U3458 (N_3458,In_598,In_211);
and U3459 (N_3459,In_1718,In_1274);
nor U3460 (N_3460,In_757,In_1875);
or U3461 (N_3461,In_945,In_110);
and U3462 (N_3462,In_1485,In_347);
nor U3463 (N_3463,In_1024,In_676);
xnor U3464 (N_3464,In_524,In_1939);
xnor U3465 (N_3465,In_1095,In_1419);
xor U3466 (N_3466,In_1031,In_1046);
xor U3467 (N_3467,In_1644,In_265);
nand U3468 (N_3468,In_1642,In_1193);
and U3469 (N_3469,In_1049,In_1965);
nand U3470 (N_3470,In_200,In_1333);
nor U3471 (N_3471,In_1700,In_1556);
or U3472 (N_3472,In_1446,In_1471);
or U3473 (N_3473,In_723,In_1641);
or U3474 (N_3474,In_309,In_1069);
nand U3475 (N_3475,In_108,In_243);
and U3476 (N_3476,In_509,In_1747);
nor U3477 (N_3477,In_410,In_1945);
and U3478 (N_3478,In_1935,In_307);
nor U3479 (N_3479,In_1150,In_664);
and U3480 (N_3480,In_377,In_1601);
and U3481 (N_3481,In_755,In_189);
or U3482 (N_3482,In_315,In_1359);
or U3483 (N_3483,In_1769,In_54);
or U3484 (N_3484,In_1383,In_104);
and U3485 (N_3485,In_662,In_266);
xnor U3486 (N_3486,In_57,In_1678);
nor U3487 (N_3487,In_778,In_363);
nand U3488 (N_3488,In_1506,In_927);
and U3489 (N_3489,In_1893,In_414);
nor U3490 (N_3490,In_1740,In_1717);
nor U3491 (N_3491,In_1859,In_1112);
nor U3492 (N_3492,In_1837,In_1546);
or U3493 (N_3493,In_917,In_250);
xor U3494 (N_3494,In_1651,In_1661);
or U3495 (N_3495,In_858,In_1558);
or U3496 (N_3496,In_143,In_1949);
or U3497 (N_3497,In_340,In_783);
nand U3498 (N_3498,In_1190,In_1364);
nand U3499 (N_3499,In_1534,In_1208);
or U3500 (N_3500,In_306,In_170);
nor U3501 (N_3501,In_661,In_929);
nor U3502 (N_3502,In_37,In_1473);
xor U3503 (N_3503,In_1070,In_981);
nor U3504 (N_3504,In_1119,In_1201);
or U3505 (N_3505,In_126,In_580);
xnor U3506 (N_3506,In_182,In_1416);
and U3507 (N_3507,In_1726,In_1222);
or U3508 (N_3508,In_249,In_793);
and U3509 (N_3509,In_129,In_325);
nor U3510 (N_3510,In_1184,In_1029);
and U3511 (N_3511,In_765,In_380);
nand U3512 (N_3512,In_71,In_484);
nor U3513 (N_3513,In_997,In_303);
xnor U3514 (N_3514,In_1615,In_531);
xor U3515 (N_3515,In_992,In_384);
nor U3516 (N_3516,In_487,In_1161);
and U3517 (N_3517,In_842,In_1481);
and U3518 (N_3518,In_226,In_1397);
nand U3519 (N_3519,In_824,In_1012);
xor U3520 (N_3520,In_1983,In_1859);
nor U3521 (N_3521,In_76,In_1555);
xor U3522 (N_3522,In_463,In_692);
xor U3523 (N_3523,In_125,In_1152);
and U3524 (N_3524,In_898,In_733);
and U3525 (N_3525,In_126,In_1837);
and U3526 (N_3526,In_1068,In_1944);
xor U3527 (N_3527,In_1774,In_1921);
and U3528 (N_3528,In_1527,In_334);
or U3529 (N_3529,In_412,In_1200);
or U3530 (N_3530,In_365,In_181);
xor U3531 (N_3531,In_867,In_966);
nand U3532 (N_3532,In_1132,In_804);
nor U3533 (N_3533,In_737,In_998);
and U3534 (N_3534,In_528,In_1072);
and U3535 (N_3535,In_1859,In_1367);
xor U3536 (N_3536,In_1403,In_796);
and U3537 (N_3537,In_95,In_359);
nand U3538 (N_3538,In_74,In_299);
xor U3539 (N_3539,In_1019,In_1340);
xnor U3540 (N_3540,In_1853,In_707);
xnor U3541 (N_3541,In_1706,In_1936);
or U3542 (N_3542,In_1509,In_994);
or U3543 (N_3543,In_1793,In_343);
nor U3544 (N_3544,In_83,In_1240);
xnor U3545 (N_3545,In_1540,In_133);
nand U3546 (N_3546,In_242,In_867);
nor U3547 (N_3547,In_1287,In_345);
nand U3548 (N_3548,In_52,In_487);
nor U3549 (N_3549,In_1041,In_1864);
nand U3550 (N_3550,In_1922,In_1147);
and U3551 (N_3551,In_1961,In_163);
nand U3552 (N_3552,In_1743,In_1934);
nor U3553 (N_3553,In_177,In_1651);
xor U3554 (N_3554,In_264,In_634);
nor U3555 (N_3555,In_632,In_606);
and U3556 (N_3556,In_800,In_705);
xor U3557 (N_3557,In_87,In_1850);
nor U3558 (N_3558,In_1575,In_211);
and U3559 (N_3559,In_205,In_1787);
or U3560 (N_3560,In_578,In_917);
nor U3561 (N_3561,In_1616,In_272);
and U3562 (N_3562,In_1536,In_489);
nand U3563 (N_3563,In_788,In_1326);
xnor U3564 (N_3564,In_1927,In_516);
and U3565 (N_3565,In_946,In_407);
nand U3566 (N_3566,In_1618,In_559);
nor U3567 (N_3567,In_843,In_411);
or U3568 (N_3568,In_345,In_875);
xor U3569 (N_3569,In_311,In_1245);
or U3570 (N_3570,In_1862,In_160);
xor U3571 (N_3571,In_527,In_436);
xor U3572 (N_3572,In_582,In_1643);
xnor U3573 (N_3573,In_1111,In_419);
xor U3574 (N_3574,In_1038,In_971);
nor U3575 (N_3575,In_657,In_1965);
or U3576 (N_3576,In_1664,In_390);
nand U3577 (N_3577,In_1018,In_1304);
and U3578 (N_3578,In_636,In_992);
nand U3579 (N_3579,In_1708,In_324);
and U3580 (N_3580,In_1734,In_641);
nand U3581 (N_3581,In_426,In_649);
and U3582 (N_3582,In_483,In_1131);
xnor U3583 (N_3583,In_1517,In_1233);
nand U3584 (N_3584,In_1965,In_903);
nor U3585 (N_3585,In_572,In_1026);
nor U3586 (N_3586,In_30,In_497);
nand U3587 (N_3587,In_1615,In_761);
xor U3588 (N_3588,In_1711,In_413);
and U3589 (N_3589,In_1556,In_1232);
or U3590 (N_3590,In_1949,In_833);
nand U3591 (N_3591,In_1329,In_1521);
xnor U3592 (N_3592,In_1199,In_1634);
nand U3593 (N_3593,In_1069,In_1168);
nor U3594 (N_3594,In_1149,In_1037);
or U3595 (N_3595,In_1114,In_1410);
or U3596 (N_3596,In_1525,In_154);
nor U3597 (N_3597,In_424,In_1697);
nand U3598 (N_3598,In_1777,In_360);
xnor U3599 (N_3599,In_1836,In_1593);
or U3600 (N_3600,In_87,In_904);
nor U3601 (N_3601,In_835,In_77);
nand U3602 (N_3602,In_986,In_54);
or U3603 (N_3603,In_719,In_1084);
xnor U3604 (N_3604,In_915,In_148);
xnor U3605 (N_3605,In_941,In_641);
nor U3606 (N_3606,In_938,In_1146);
nor U3607 (N_3607,In_385,In_1255);
and U3608 (N_3608,In_82,In_94);
nor U3609 (N_3609,In_836,In_897);
or U3610 (N_3610,In_309,In_906);
or U3611 (N_3611,In_1988,In_228);
xnor U3612 (N_3612,In_1813,In_95);
xor U3613 (N_3613,In_1465,In_1866);
and U3614 (N_3614,In_1018,In_851);
and U3615 (N_3615,In_279,In_1561);
xnor U3616 (N_3616,In_970,In_1160);
nand U3617 (N_3617,In_1347,In_981);
or U3618 (N_3618,In_1363,In_1379);
xor U3619 (N_3619,In_1345,In_1774);
and U3620 (N_3620,In_1752,In_1516);
and U3621 (N_3621,In_975,In_697);
or U3622 (N_3622,In_431,In_1225);
or U3623 (N_3623,In_311,In_590);
and U3624 (N_3624,In_772,In_1834);
xnor U3625 (N_3625,In_455,In_707);
nor U3626 (N_3626,In_901,In_1905);
or U3627 (N_3627,In_1565,In_161);
nor U3628 (N_3628,In_221,In_1224);
xnor U3629 (N_3629,In_1179,In_1406);
nand U3630 (N_3630,In_92,In_352);
or U3631 (N_3631,In_1665,In_591);
nand U3632 (N_3632,In_589,In_1050);
and U3633 (N_3633,In_334,In_1283);
xor U3634 (N_3634,In_1981,In_710);
nor U3635 (N_3635,In_791,In_1082);
xor U3636 (N_3636,In_1425,In_1611);
nor U3637 (N_3637,In_1531,In_1444);
nand U3638 (N_3638,In_143,In_1979);
nor U3639 (N_3639,In_1442,In_1419);
and U3640 (N_3640,In_1758,In_1415);
xor U3641 (N_3641,In_1055,In_1118);
and U3642 (N_3642,In_685,In_53);
nor U3643 (N_3643,In_122,In_1105);
and U3644 (N_3644,In_940,In_1949);
and U3645 (N_3645,In_1902,In_770);
xnor U3646 (N_3646,In_51,In_1612);
and U3647 (N_3647,In_890,In_1958);
and U3648 (N_3648,In_1294,In_424);
xnor U3649 (N_3649,In_1091,In_1922);
or U3650 (N_3650,In_1729,In_1323);
or U3651 (N_3651,In_1870,In_945);
xnor U3652 (N_3652,In_1854,In_93);
xnor U3653 (N_3653,In_1954,In_166);
nand U3654 (N_3654,In_279,In_1695);
or U3655 (N_3655,In_765,In_191);
and U3656 (N_3656,In_599,In_126);
nand U3657 (N_3657,In_221,In_832);
xor U3658 (N_3658,In_737,In_550);
nor U3659 (N_3659,In_670,In_1355);
and U3660 (N_3660,In_726,In_312);
and U3661 (N_3661,In_849,In_1573);
nand U3662 (N_3662,In_1925,In_609);
or U3663 (N_3663,In_587,In_1506);
nand U3664 (N_3664,In_1949,In_988);
nor U3665 (N_3665,In_89,In_166);
nor U3666 (N_3666,In_1153,In_1681);
and U3667 (N_3667,In_171,In_66);
nand U3668 (N_3668,In_551,In_876);
nor U3669 (N_3669,In_1574,In_709);
xor U3670 (N_3670,In_1415,In_903);
xor U3671 (N_3671,In_1042,In_613);
or U3672 (N_3672,In_1254,In_1606);
nor U3673 (N_3673,In_958,In_1345);
xor U3674 (N_3674,In_840,In_1785);
or U3675 (N_3675,In_683,In_1990);
and U3676 (N_3676,In_112,In_1109);
xnor U3677 (N_3677,In_1016,In_1958);
nand U3678 (N_3678,In_1493,In_1193);
xor U3679 (N_3679,In_66,In_1071);
nand U3680 (N_3680,In_1573,In_1923);
or U3681 (N_3681,In_59,In_256);
xnor U3682 (N_3682,In_1381,In_263);
nand U3683 (N_3683,In_541,In_1159);
nand U3684 (N_3684,In_1195,In_1205);
nand U3685 (N_3685,In_362,In_883);
nor U3686 (N_3686,In_485,In_1892);
xnor U3687 (N_3687,In_1574,In_60);
or U3688 (N_3688,In_760,In_231);
or U3689 (N_3689,In_259,In_1035);
nor U3690 (N_3690,In_1744,In_1313);
nand U3691 (N_3691,In_1799,In_1038);
nand U3692 (N_3692,In_164,In_1074);
nor U3693 (N_3693,In_15,In_393);
or U3694 (N_3694,In_134,In_63);
nand U3695 (N_3695,In_1452,In_541);
nor U3696 (N_3696,In_172,In_267);
or U3697 (N_3697,In_395,In_974);
or U3698 (N_3698,In_1952,In_498);
xnor U3699 (N_3699,In_322,In_1699);
or U3700 (N_3700,In_1005,In_442);
nand U3701 (N_3701,In_930,In_592);
xor U3702 (N_3702,In_1617,In_1034);
and U3703 (N_3703,In_818,In_634);
or U3704 (N_3704,In_1886,In_909);
and U3705 (N_3705,In_839,In_41);
xor U3706 (N_3706,In_316,In_873);
nand U3707 (N_3707,In_1792,In_633);
nor U3708 (N_3708,In_1052,In_885);
xor U3709 (N_3709,In_675,In_1471);
nand U3710 (N_3710,In_406,In_1848);
and U3711 (N_3711,In_697,In_1787);
nand U3712 (N_3712,In_769,In_629);
or U3713 (N_3713,In_236,In_498);
xnor U3714 (N_3714,In_1869,In_1032);
xnor U3715 (N_3715,In_464,In_410);
and U3716 (N_3716,In_790,In_120);
xnor U3717 (N_3717,In_1743,In_1157);
and U3718 (N_3718,In_798,In_1112);
nor U3719 (N_3719,In_1646,In_980);
xnor U3720 (N_3720,In_1403,In_38);
nand U3721 (N_3721,In_1083,In_1815);
or U3722 (N_3722,In_1448,In_128);
nor U3723 (N_3723,In_716,In_828);
or U3724 (N_3724,In_1120,In_253);
xor U3725 (N_3725,In_452,In_1152);
nand U3726 (N_3726,In_1722,In_1880);
nand U3727 (N_3727,In_718,In_1802);
nand U3728 (N_3728,In_71,In_568);
and U3729 (N_3729,In_1714,In_1407);
nor U3730 (N_3730,In_600,In_713);
nand U3731 (N_3731,In_1684,In_634);
or U3732 (N_3732,In_171,In_1322);
xor U3733 (N_3733,In_1706,In_1722);
nand U3734 (N_3734,In_1682,In_1908);
and U3735 (N_3735,In_699,In_737);
nand U3736 (N_3736,In_505,In_1221);
nand U3737 (N_3737,In_523,In_1241);
or U3738 (N_3738,In_579,In_898);
nor U3739 (N_3739,In_1524,In_1473);
and U3740 (N_3740,In_466,In_398);
nor U3741 (N_3741,In_1944,In_844);
or U3742 (N_3742,In_3,In_1480);
or U3743 (N_3743,In_854,In_272);
nand U3744 (N_3744,In_49,In_630);
nor U3745 (N_3745,In_1220,In_1396);
or U3746 (N_3746,In_244,In_410);
or U3747 (N_3747,In_777,In_520);
or U3748 (N_3748,In_1148,In_563);
and U3749 (N_3749,In_1023,In_357);
nand U3750 (N_3750,In_1561,In_1158);
xnor U3751 (N_3751,In_1547,In_0);
xnor U3752 (N_3752,In_1453,In_1731);
xnor U3753 (N_3753,In_1244,In_1356);
or U3754 (N_3754,In_661,In_453);
or U3755 (N_3755,In_497,In_509);
nand U3756 (N_3756,In_1258,In_305);
xnor U3757 (N_3757,In_609,In_1490);
nand U3758 (N_3758,In_1020,In_1458);
nor U3759 (N_3759,In_1746,In_1142);
and U3760 (N_3760,In_489,In_949);
xor U3761 (N_3761,In_1285,In_577);
nor U3762 (N_3762,In_779,In_949);
and U3763 (N_3763,In_1168,In_1153);
nand U3764 (N_3764,In_527,In_1226);
or U3765 (N_3765,In_180,In_1791);
nor U3766 (N_3766,In_1689,In_151);
xor U3767 (N_3767,In_851,In_1711);
or U3768 (N_3768,In_1,In_764);
or U3769 (N_3769,In_139,In_328);
nor U3770 (N_3770,In_625,In_1452);
or U3771 (N_3771,In_1152,In_1796);
or U3772 (N_3772,In_686,In_1559);
nand U3773 (N_3773,In_280,In_986);
and U3774 (N_3774,In_1362,In_760);
nand U3775 (N_3775,In_1164,In_1621);
or U3776 (N_3776,In_745,In_1898);
and U3777 (N_3777,In_1189,In_1798);
nand U3778 (N_3778,In_1232,In_1293);
or U3779 (N_3779,In_1405,In_1923);
xnor U3780 (N_3780,In_210,In_1657);
nor U3781 (N_3781,In_1937,In_49);
xor U3782 (N_3782,In_1001,In_557);
or U3783 (N_3783,In_770,In_679);
nand U3784 (N_3784,In_1762,In_1958);
nor U3785 (N_3785,In_136,In_947);
or U3786 (N_3786,In_1778,In_114);
nand U3787 (N_3787,In_246,In_47);
and U3788 (N_3788,In_1871,In_1406);
xor U3789 (N_3789,In_1291,In_731);
xnor U3790 (N_3790,In_824,In_1890);
xnor U3791 (N_3791,In_919,In_854);
xor U3792 (N_3792,In_1404,In_978);
and U3793 (N_3793,In_712,In_147);
nor U3794 (N_3794,In_1534,In_1089);
nor U3795 (N_3795,In_1031,In_115);
and U3796 (N_3796,In_1075,In_82);
nor U3797 (N_3797,In_1689,In_671);
nand U3798 (N_3798,In_1636,In_718);
or U3799 (N_3799,In_924,In_115);
and U3800 (N_3800,In_1503,In_832);
xnor U3801 (N_3801,In_975,In_496);
xnor U3802 (N_3802,In_208,In_504);
nand U3803 (N_3803,In_1387,In_12);
nand U3804 (N_3804,In_717,In_240);
nand U3805 (N_3805,In_1267,In_1113);
xnor U3806 (N_3806,In_1725,In_1565);
nand U3807 (N_3807,In_1759,In_229);
nand U3808 (N_3808,In_763,In_1443);
nor U3809 (N_3809,In_501,In_988);
nand U3810 (N_3810,In_646,In_1612);
and U3811 (N_3811,In_79,In_1491);
nor U3812 (N_3812,In_1717,In_119);
nor U3813 (N_3813,In_886,In_1497);
or U3814 (N_3814,In_107,In_172);
or U3815 (N_3815,In_1265,In_942);
and U3816 (N_3816,In_1062,In_1369);
xnor U3817 (N_3817,In_975,In_395);
nand U3818 (N_3818,In_608,In_1364);
or U3819 (N_3819,In_587,In_1776);
or U3820 (N_3820,In_9,In_1844);
nor U3821 (N_3821,In_1068,In_355);
or U3822 (N_3822,In_1625,In_1611);
nor U3823 (N_3823,In_421,In_990);
or U3824 (N_3824,In_781,In_337);
and U3825 (N_3825,In_1430,In_1558);
and U3826 (N_3826,In_1831,In_1858);
nand U3827 (N_3827,In_1072,In_1346);
and U3828 (N_3828,In_1229,In_595);
or U3829 (N_3829,In_693,In_897);
and U3830 (N_3830,In_616,In_296);
or U3831 (N_3831,In_1159,In_600);
xor U3832 (N_3832,In_348,In_1926);
and U3833 (N_3833,In_1646,In_1242);
xor U3834 (N_3834,In_466,In_889);
nand U3835 (N_3835,In_304,In_1778);
nor U3836 (N_3836,In_1269,In_1928);
and U3837 (N_3837,In_523,In_538);
or U3838 (N_3838,In_837,In_1350);
and U3839 (N_3839,In_518,In_948);
and U3840 (N_3840,In_222,In_1680);
nand U3841 (N_3841,In_376,In_1288);
nand U3842 (N_3842,In_1015,In_1994);
and U3843 (N_3843,In_589,In_49);
nor U3844 (N_3844,In_1344,In_1154);
nand U3845 (N_3845,In_1222,In_328);
nand U3846 (N_3846,In_341,In_901);
and U3847 (N_3847,In_1633,In_1319);
and U3848 (N_3848,In_621,In_1261);
nor U3849 (N_3849,In_1647,In_1409);
or U3850 (N_3850,In_743,In_1537);
nor U3851 (N_3851,In_49,In_559);
and U3852 (N_3852,In_331,In_1504);
and U3853 (N_3853,In_784,In_1239);
nor U3854 (N_3854,In_237,In_1974);
nor U3855 (N_3855,In_1317,In_282);
nand U3856 (N_3856,In_1752,In_725);
or U3857 (N_3857,In_1614,In_78);
nand U3858 (N_3858,In_208,In_1513);
and U3859 (N_3859,In_1125,In_983);
or U3860 (N_3860,In_1791,In_247);
and U3861 (N_3861,In_739,In_158);
nor U3862 (N_3862,In_263,In_907);
and U3863 (N_3863,In_1121,In_908);
or U3864 (N_3864,In_741,In_1617);
nor U3865 (N_3865,In_1389,In_1559);
or U3866 (N_3866,In_1160,In_762);
xor U3867 (N_3867,In_206,In_1539);
and U3868 (N_3868,In_1918,In_566);
and U3869 (N_3869,In_1217,In_1430);
and U3870 (N_3870,In_645,In_889);
xnor U3871 (N_3871,In_728,In_622);
xnor U3872 (N_3872,In_1724,In_757);
nand U3873 (N_3873,In_694,In_569);
nand U3874 (N_3874,In_66,In_361);
xnor U3875 (N_3875,In_668,In_510);
or U3876 (N_3876,In_1379,In_478);
nand U3877 (N_3877,In_1553,In_1647);
nor U3878 (N_3878,In_155,In_19);
nand U3879 (N_3879,In_948,In_1694);
and U3880 (N_3880,In_20,In_1391);
nand U3881 (N_3881,In_1882,In_1216);
or U3882 (N_3882,In_541,In_437);
xor U3883 (N_3883,In_617,In_1934);
nor U3884 (N_3884,In_1857,In_1541);
nor U3885 (N_3885,In_529,In_580);
nor U3886 (N_3886,In_428,In_1790);
nor U3887 (N_3887,In_793,In_1438);
and U3888 (N_3888,In_508,In_1235);
or U3889 (N_3889,In_702,In_1278);
xor U3890 (N_3890,In_1393,In_1416);
and U3891 (N_3891,In_1837,In_554);
xnor U3892 (N_3892,In_1559,In_1894);
nor U3893 (N_3893,In_1385,In_1053);
nor U3894 (N_3894,In_328,In_1671);
or U3895 (N_3895,In_1483,In_568);
xnor U3896 (N_3896,In_413,In_1883);
xor U3897 (N_3897,In_590,In_609);
or U3898 (N_3898,In_1233,In_1739);
and U3899 (N_3899,In_447,In_561);
and U3900 (N_3900,In_1532,In_404);
xnor U3901 (N_3901,In_1302,In_396);
nand U3902 (N_3902,In_1540,In_1566);
and U3903 (N_3903,In_464,In_1126);
nand U3904 (N_3904,In_1433,In_1648);
or U3905 (N_3905,In_257,In_1191);
or U3906 (N_3906,In_832,In_762);
and U3907 (N_3907,In_1268,In_1387);
nand U3908 (N_3908,In_76,In_438);
or U3909 (N_3909,In_97,In_1104);
and U3910 (N_3910,In_1588,In_684);
or U3911 (N_3911,In_1552,In_241);
nor U3912 (N_3912,In_1265,In_1747);
nand U3913 (N_3913,In_324,In_707);
and U3914 (N_3914,In_670,In_667);
and U3915 (N_3915,In_633,In_1195);
nand U3916 (N_3916,In_1641,In_1284);
nor U3917 (N_3917,In_711,In_193);
xor U3918 (N_3918,In_983,In_376);
or U3919 (N_3919,In_58,In_1252);
and U3920 (N_3920,In_1470,In_1003);
and U3921 (N_3921,In_172,In_402);
nor U3922 (N_3922,In_1577,In_55);
and U3923 (N_3923,In_782,In_633);
and U3924 (N_3924,In_458,In_1268);
nor U3925 (N_3925,In_1217,In_1913);
xor U3926 (N_3926,In_1676,In_1279);
xor U3927 (N_3927,In_1351,In_1850);
nor U3928 (N_3928,In_996,In_1213);
and U3929 (N_3929,In_774,In_861);
and U3930 (N_3930,In_1974,In_114);
and U3931 (N_3931,In_741,In_265);
or U3932 (N_3932,In_905,In_1331);
nand U3933 (N_3933,In_1958,In_230);
or U3934 (N_3934,In_990,In_912);
nand U3935 (N_3935,In_1884,In_1777);
nor U3936 (N_3936,In_115,In_145);
nor U3937 (N_3937,In_1739,In_442);
nand U3938 (N_3938,In_1605,In_1733);
nor U3939 (N_3939,In_1993,In_1159);
nor U3940 (N_3940,In_1486,In_305);
nand U3941 (N_3941,In_1339,In_532);
nor U3942 (N_3942,In_1706,In_1805);
nor U3943 (N_3943,In_1254,In_161);
nor U3944 (N_3944,In_398,In_1272);
nand U3945 (N_3945,In_325,In_792);
nand U3946 (N_3946,In_269,In_1465);
or U3947 (N_3947,In_1921,In_368);
or U3948 (N_3948,In_1929,In_994);
or U3949 (N_3949,In_1298,In_1665);
xor U3950 (N_3950,In_743,In_208);
or U3951 (N_3951,In_594,In_1445);
or U3952 (N_3952,In_1960,In_581);
nand U3953 (N_3953,In_559,In_1709);
or U3954 (N_3954,In_909,In_1381);
and U3955 (N_3955,In_1054,In_625);
xnor U3956 (N_3956,In_333,In_1273);
nor U3957 (N_3957,In_1453,In_1011);
xnor U3958 (N_3958,In_527,In_17);
nand U3959 (N_3959,In_556,In_550);
nand U3960 (N_3960,In_1076,In_1816);
nand U3961 (N_3961,In_1751,In_1617);
and U3962 (N_3962,In_1881,In_573);
or U3963 (N_3963,In_129,In_1670);
nand U3964 (N_3964,In_1711,In_1633);
nand U3965 (N_3965,In_1984,In_566);
and U3966 (N_3966,In_1301,In_1819);
nor U3967 (N_3967,In_1176,In_1185);
xor U3968 (N_3968,In_883,In_939);
or U3969 (N_3969,In_1491,In_1068);
nor U3970 (N_3970,In_203,In_697);
nor U3971 (N_3971,In_536,In_1197);
nor U3972 (N_3972,In_1704,In_189);
xnor U3973 (N_3973,In_52,In_430);
xor U3974 (N_3974,In_1617,In_187);
and U3975 (N_3975,In_1425,In_972);
nor U3976 (N_3976,In_1038,In_1029);
and U3977 (N_3977,In_1906,In_148);
and U3978 (N_3978,In_1762,In_1899);
xor U3979 (N_3979,In_1687,In_833);
or U3980 (N_3980,In_1315,In_63);
and U3981 (N_3981,In_1876,In_1943);
nor U3982 (N_3982,In_794,In_1825);
xnor U3983 (N_3983,In_457,In_1632);
or U3984 (N_3984,In_1363,In_462);
or U3985 (N_3985,In_1352,In_891);
and U3986 (N_3986,In_1235,In_1339);
nor U3987 (N_3987,In_1698,In_1086);
nor U3988 (N_3988,In_570,In_388);
and U3989 (N_3989,In_1717,In_396);
and U3990 (N_3990,In_1779,In_1361);
xor U3991 (N_3991,In_1373,In_288);
nand U3992 (N_3992,In_1656,In_1284);
and U3993 (N_3993,In_681,In_1427);
nand U3994 (N_3994,In_281,In_758);
or U3995 (N_3995,In_122,In_1037);
or U3996 (N_3996,In_1503,In_385);
nor U3997 (N_3997,In_62,In_1824);
nand U3998 (N_3998,In_1346,In_1999);
and U3999 (N_3999,In_1740,In_1362);
nand U4000 (N_4000,N_3860,N_2182);
nor U4001 (N_4001,N_286,N_1408);
nor U4002 (N_4002,N_2070,N_3762);
or U4003 (N_4003,N_737,N_856);
or U4004 (N_4004,N_1571,N_995);
nand U4005 (N_4005,N_2066,N_1863);
or U4006 (N_4006,N_1412,N_2840);
xnor U4007 (N_4007,N_2845,N_340);
nand U4008 (N_4008,N_827,N_626);
nand U4009 (N_4009,N_1372,N_71);
or U4010 (N_4010,N_2420,N_3061);
xor U4011 (N_4011,N_1790,N_3342);
and U4012 (N_4012,N_3435,N_1186);
and U4013 (N_4013,N_3464,N_3695);
or U4014 (N_4014,N_2065,N_3183);
xnor U4015 (N_4015,N_2057,N_3345);
xnor U4016 (N_4016,N_572,N_1676);
nor U4017 (N_4017,N_1485,N_2698);
nor U4018 (N_4018,N_1061,N_599);
or U4019 (N_4019,N_1470,N_210);
or U4020 (N_4020,N_968,N_1252);
and U4021 (N_4021,N_2823,N_2521);
and U4022 (N_4022,N_3262,N_534);
or U4023 (N_4023,N_613,N_1717);
nand U4024 (N_4024,N_1505,N_557);
and U4025 (N_4025,N_891,N_770);
xnor U4026 (N_4026,N_809,N_387);
and U4027 (N_4027,N_1360,N_3515);
nand U4028 (N_4028,N_3281,N_3601);
and U4029 (N_4029,N_2857,N_2341);
nor U4030 (N_4030,N_2925,N_1887);
nor U4031 (N_4031,N_2826,N_2247);
nor U4032 (N_4032,N_3182,N_2596);
or U4033 (N_4033,N_589,N_1620);
nor U4034 (N_4034,N_3484,N_2536);
nor U4035 (N_4035,N_3699,N_2712);
xnor U4036 (N_4036,N_3880,N_3198);
xor U4037 (N_4037,N_1276,N_2072);
nor U4038 (N_4038,N_2410,N_144);
or U4039 (N_4039,N_704,N_1366);
xnor U4040 (N_4040,N_135,N_2701);
nand U4041 (N_4041,N_406,N_762);
xnor U4042 (N_4042,N_1854,N_3736);
and U4043 (N_4043,N_235,N_2902);
or U4044 (N_4044,N_1472,N_1826);
or U4045 (N_4045,N_1204,N_3790);
nor U4046 (N_4046,N_265,N_3213);
or U4047 (N_4047,N_543,N_571);
and U4048 (N_4048,N_461,N_1179);
xor U4049 (N_4049,N_3275,N_2696);
nand U4050 (N_4050,N_2031,N_1441);
or U4051 (N_4051,N_3993,N_1088);
or U4052 (N_4052,N_2073,N_1110);
and U4053 (N_4053,N_1947,N_3769);
nor U4054 (N_4054,N_2822,N_330);
nand U4055 (N_4055,N_3392,N_1246);
nand U4056 (N_4056,N_3130,N_3765);
and U4057 (N_4057,N_3547,N_2255);
nor U4058 (N_4058,N_917,N_266);
and U4059 (N_4059,N_1296,N_3509);
nor U4060 (N_4060,N_3441,N_1396);
or U4061 (N_4061,N_3384,N_2952);
xor U4062 (N_4062,N_1748,N_3440);
nor U4063 (N_4063,N_444,N_2135);
nor U4064 (N_4064,N_2454,N_3059);
nor U4065 (N_4065,N_1847,N_498);
nand U4066 (N_4066,N_1253,N_3598);
nor U4067 (N_4067,N_2127,N_10);
or U4068 (N_4068,N_3062,N_1593);
xnor U4069 (N_4069,N_434,N_3690);
nand U4070 (N_4070,N_1096,N_2608);
and U4071 (N_4071,N_979,N_1758);
nor U4072 (N_4072,N_1168,N_2002);
xor U4073 (N_4073,N_108,N_1310);
nand U4074 (N_4074,N_1487,N_2688);
xnor U4075 (N_4075,N_919,N_637);
xor U4076 (N_4076,N_148,N_2911);
nand U4077 (N_4077,N_3636,N_3840);
nor U4078 (N_4078,N_769,N_416);
xor U4079 (N_4079,N_2354,N_399);
nor U4080 (N_4080,N_1953,N_1963);
nor U4081 (N_4081,N_173,N_2415);
nor U4082 (N_4082,N_33,N_2981);
and U4083 (N_4083,N_15,N_1226);
nand U4084 (N_4084,N_3206,N_2099);
nand U4085 (N_4085,N_511,N_586);
or U4086 (N_4086,N_2196,N_1386);
or U4087 (N_4087,N_3556,N_3312);
or U4088 (N_4088,N_3569,N_2783);
nand U4089 (N_4089,N_3128,N_3862);
or U4090 (N_4090,N_1741,N_2277);
nor U4091 (N_4091,N_1494,N_2498);
nor U4092 (N_4092,N_2233,N_427);
and U4093 (N_4093,N_1585,N_713);
and U4094 (N_4094,N_2257,N_2625);
or U4095 (N_4095,N_2191,N_2814);
and U4096 (N_4096,N_3521,N_166);
nor U4097 (N_4097,N_963,N_3463);
and U4098 (N_4098,N_3118,N_3063);
and U4099 (N_4099,N_729,N_4);
nand U4100 (N_4100,N_250,N_1903);
xnor U4101 (N_4101,N_3095,N_2437);
nor U4102 (N_4102,N_2392,N_966);
nand U4103 (N_4103,N_2612,N_2560);
and U4104 (N_4104,N_1488,N_3012);
or U4105 (N_4105,N_3592,N_3416);
nor U4106 (N_4106,N_1218,N_2004);
or U4107 (N_4107,N_3496,N_3401);
xor U4108 (N_4108,N_753,N_40);
xnor U4109 (N_4109,N_2744,N_243);
nor U4110 (N_4110,N_843,N_1591);
nor U4111 (N_4111,N_227,N_2000);
or U4112 (N_4112,N_1673,N_3196);
or U4113 (N_4113,N_2644,N_2329);
and U4114 (N_4114,N_1803,N_3498);
nand U4115 (N_4115,N_579,N_186);
nor U4116 (N_4116,N_897,N_3579);
xnor U4117 (N_4117,N_1261,N_411);
nor U4118 (N_4118,N_2846,N_2145);
or U4119 (N_4119,N_1525,N_1848);
nand U4120 (N_4120,N_1931,N_196);
nor U4121 (N_4121,N_1517,N_3574);
nor U4122 (N_4122,N_2890,N_3113);
or U4123 (N_4123,N_3814,N_938);
or U4124 (N_4124,N_1772,N_366);
or U4125 (N_4125,N_3507,N_2317);
xnor U4126 (N_4126,N_1780,N_652);
or U4127 (N_4127,N_3259,N_92);
nor U4128 (N_4128,N_2047,N_2243);
and U4129 (N_4129,N_3677,N_3589);
nor U4130 (N_4130,N_275,N_3044);
nand U4131 (N_4131,N_1180,N_1402);
or U4132 (N_4132,N_2754,N_2969);
and U4133 (N_4133,N_1207,N_3261);
xor U4134 (N_4134,N_2155,N_395);
nor U4135 (N_4135,N_2286,N_2339);
and U4136 (N_4136,N_3249,N_1012);
or U4137 (N_4137,N_3678,N_288);
xor U4138 (N_4138,N_2284,N_794);
xor U4139 (N_4139,N_3223,N_3353);
or U4140 (N_4140,N_192,N_3133);
xnor U4141 (N_4141,N_583,N_1922);
nand U4142 (N_4142,N_428,N_2610);
nand U4143 (N_4143,N_1380,N_338);
xor U4144 (N_4144,N_2595,N_117);
nand U4145 (N_4145,N_1556,N_3268);
xor U4146 (N_4146,N_2861,N_388);
nor U4147 (N_4147,N_3869,N_2051);
xor U4148 (N_4148,N_742,N_2796);
nand U4149 (N_4149,N_170,N_2882);
and U4150 (N_4150,N_1646,N_3181);
and U4151 (N_4151,N_1552,N_956);
or U4152 (N_4152,N_2888,N_2935);
nor U4153 (N_4153,N_3240,N_1073);
and U4154 (N_4154,N_3823,N_2507);
and U4155 (N_4155,N_3174,N_2787);
or U4156 (N_4156,N_535,N_3753);
and U4157 (N_4157,N_2393,N_1794);
and U4158 (N_4158,N_3145,N_3821);
nor U4159 (N_4159,N_3089,N_1555);
nand U4160 (N_4160,N_2776,N_3369);
nand U4161 (N_4161,N_2795,N_582);
nor U4162 (N_4162,N_3479,N_2199);
and U4163 (N_4163,N_736,N_258);
nor U4164 (N_4164,N_1781,N_2742);
nor U4165 (N_4165,N_1216,N_1833);
and U4166 (N_4166,N_1969,N_3287);
xor U4167 (N_4167,N_2734,N_2957);
nand U4168 (N_4168,N_2267,N_2953);
or U4169 (N_4169,N_2631,N_1559);
nand U4170 (N_4170,N_3791,N_1562);
or U4171 (N_4171,N_601,N_3512);
xor U4172 (N_4172,N_510,N_1866);
and U4173 (N_4173,N_3947,N_2933);
xnor U4174 (N_4174,N_871,N_1263);
and U4175 (N_4175,N_2574,N_329);
nand U4176 (N_4176,N_1404,N_1578);
and U4177 (N_4177,N_270,N_2236);
nor U4178 (N_4178,N_2308,N_3140);
and U4179 (N_4179,N_189,N_2697);
or U4180 (N_4180,N_1724,N_442);
and U4181 (N_4181,N_129,N_3684);
and U4182 (N_4182,N_3934,N_1846);
xor U4183 (N_4183,N_3752,N_38);
nand U4184 (N_4184,N_726,N_3717);
and U4185 (N_4185,N_2997,N_905);
nor U4186 (N_4186,N_101,N_2088);
or U4187 (N_4187,N_765,N_3469);
xor U4188 (N_4188,N_3746,N_495);
nor U4189 (N_4189,N_1280,N_1375);
or U4190 (N_4190,N_1669,N_894);
xor U4191 (N_4191,N_487,N_2086);
and U4192 (N_4192,N_3266,N_2683);
nand U4193 (N_4193,N_701,N_230);
or U4194 (N_4194,N_2081,N_294);
or U4195 (N_4195,N_1125,N_2640);
nor U4196 (N_4196,N_3500,N_2011);
or U4197 (N_4197,N_1522,N_2431);
xor U4198 (N_4198,N_1684,N_996);
nand U4199 (N_4199,N_3393,N_2680);
xnor U4200 (N_4200,N_3260,N_1784);
xor U4201 (N_4201,N_3945,N_2654);
or U4202 (N_4202,N_1329,N_3197);
and U4203 (N_4203,N_925,N_3400);
nand U4204 (N_4204,N_2629,N_1840);
nand U4205 (N_4205,N_2567,N_3573);
or U4206 (N_4206,N_54,N_2483);
xor U4207 (N_4207,N_3923,N_763);
nor U4208 (N_4208,N_668,N_1681);
and U4209 (N_4209,N_1190,N_2710);
or U4210 (N_4210,N_3002,N_111);
xor U4211 (N_4211,N_1901,N_1893);
nor U4212 (N_4212,N_1356,N_3562);
or U4213 (N_4213,N_3138,N_1009);
nor U4214 (N_4214,N_1611,N_641);
xor U4215 (N_4215,N_1519,N_1010);
nand U4216 (N_4216,N_2656,N_1182);
and U4217 (N_4217,N_3623,N_2883);
or U4218 (N_4218,N_2623,N_285);
nand U4219 (N_4219,N_1456,N_2666);
or U4220 (N_4220,N_342,N_946);
nand U4221 (N_4221,N_2956,N_426);
xnor U4222 (N_4222,N_1411,N_316);
or U4223 (N_4223,N_2597,N_1136);
and U4224 (N_4224,N_847,N_305);
nor U4225 (N_4225,N_3625,N_527);
nor U4226 (N_4226,N_671,N_2164);
nand U4227 (N_4227,N_1761,N_2537);
or U4228 (N_4228,N_3561,N_324);
nand U4229 (N_4229,N_3426,N_121);
xor U4230 (N_4230,N_3293,N_282);
and U4231 (N_4231,N_1899,N_1816);
xor U4232 (N_4232,N_3570,N_2063);
nand U4233 (N_4233,N_2165,N_3168);
xnor U4234 (N_4234,N_296,N_2841);
and U4235 (N_4235,N_3593,N_2604);
and U4236 (N_4236,N_2098,N_3320);
and U4237 (N_4237,N_562,N_1465);
nor U4238 (N_4238,N_2034,N_3642);
nand U4239 (N_4239,N_2657,N_1231);
or U4240 (N_4240,N_70,N_2865);
nand U4241 (N_4241,N_2777,N_2932);
and U4242 (N_4242,N_2470,N_34);
xor U4243 (N_4243,N_3207,N_3214);
nor U4244 (N_4244,N_1041,N_177);
nand U4245 (N_4245,N_32,N_1510);
nor U4246 (N_4246,N_1564,N_2248);
and U4247 (N_4247,N_1531,N_1900);
xor U4248 (N_4248,N_109,N_3641);
nor U4249 (N_4249,N_2064,N_692);
nor U4250 (N_4250,N_1227,N_3058);
or U4251 (N_4251,N_187,N_717);
and U4252 (N_4252,N_3634,N_740);
and U4253 (N_4253,N_2130,N_3740);
and U4254 (N_4254,N_419,N_2588);
and U4255 (N_4255,N_2318,N_2559);
or U4256 (N_4256,N_3487,N_2213);
nor U4257 (N_4257,N_2557,N_2749);
nand U4258 (N_4258,N_1542,N_799);
or U4259 (N_4259,N_3918,N_538);
or U4260 (N_4260,N_2143,N_1322);
nor U4261 (N_4261,N_2036,N_2812);
nand U4262 (N_4262,N_790,N_3972);
and U4263 (N_4263,N_3730,N_1986);
xor U4264 (N_4264,N_251,N_3616);
or U4265 (N_4265,N_3452,N_2077);
nand U4266 (N_4266,N_1152,N_1979);
xor U4267 (N_4267,N_3368,N_67);
nor U4268 (N_4268,N_876,N_2024);
nor U4269 (N_4269,N_1964,N_2692);
nand U4270 (N_4270,N_569,N_1929);
xor U4271 (N_4271,N_2979,N_3597);
nor U4272 (N_4272,N_1738,N_3729);
or U4273 (N_4273,N_3865,N_3131);
xor U4274 (N_4274,N_1130,N_1289);
or U4275 (N_4275,N_1513,N_677);
or U4276 (N_4276,N_1912,N_3074);
xor U4277 (N_4277,N_1539,N_2529);
nand U4278 (N_4278,N_180,N_3221);
nand U4279 (N_4279,N_1362,N_3780);
or U4280 (N_4280,N_1813,N_2531);
nand U4281 (N_4281,N_1657,N_3427);
nor U4282 (N_4282,N_2091,N_2565);
xor U4283 (N_4283,N_2043,N_2076);
nor U4284 (N_4284,N_1077,N_999);
nor U4285 (N_4285,N_57,N_1504);
xor U4286 (N_4286,N_676,N_1581);
or U4287 (N_4287,N_3888,N_3748);
or U4288 (N_4288,N_568,N_2068);
and U4289 (N_4289,N_530,N_3785);
xor U4290 (N_4290,N_2111,N_649);
nor U4291 (N_4291,N_2179,N_3352);
and U4292 (N_4292,N_3167,N_3478);
and U4293 (N_4293,N_1131,N_371);
nand U4294 (N_4294,N_1115,N_3600);
nand U4295 (N_4295,N_1043,N_3473);
and U4296 (N_4296,N_708,N_2951);
nor U4297 (N_4297,N_2961,N_2092);
nor U4298 (N_4298,N_2627,N_3170);
or U4299 (N_4299,N_942,N_683);
and U4300 (N_4300,N_2722,N_2891);
or U4301 (N_4301,N_307,N_1870);
nor U4302 (N_4302,N_3318,N_1944);
nor U4303 (N_4303,N_2794,N_2601);
xor U4304 (N_4304,N_1316,N_2839);
and U4305 (N_4305,N_2922,N_273);
xnor U4306 (N_4306,N_2575,N_72);
nand U4307 (N_4307,N_935,N_659);
nand U4308 (N_4308,N_1236,N_875);
nor U4309 (N_4309,N_2832,N_3157);
nand U4310 (N_4310,N_801,N_3703);
or U4311 (N_4311,N_1254,N_2869);
or U4312 (N_4312,N_2101,N_2995);
nand U4313 (N_4313,N_1883,N_3870);
or U4314 (N_4314,N_3192,N_1199);
xor U4315 (N_4315,N_1016,N_1732);
nand U4316 (N_4316,N_597,N_2514);
and U4317 (N_4317,N_3661,N_1175);
and U4318 (N_4318,N_3687,N_2798);
and U4319 (N_4319,N_3408,N_616);
or U4320 (N_4320,N_3347,N_1647);
nor U4321 (N_4321,N_482,N_224);
xor U4322 (N_4322,N_1425,N_2301);
xnor U4323 (N_4323,N_2705,N_3257);
and U4324 (N_4324,N_2039,N_2947);
and U4325 (N_4325,N_3,N_1683);
and U4326 (N_4326,N_1224,N_118);
or U4327 (N_4327,N_3913,N_2180);
nand U4328 (N_4328,N_700,N_2365);
nor U4329 (N_4329,N_3404,N_1797);
xor U4330 (N_4330,N_1595,N_382);
or U4331 (N_4331,N_420,N_2381);
nand U4332 (N_4332,N_1331,N_1643);
nand U4333 (N_4333,N_673,N_3092);
xor U4334 (N_4334,N_1975,N_3632);
and U4335 (N_4335,N_413,N_289);
or U4336 (N_4336,N_185,N_1145);
nand U4337 (N_4337,N_3071,N_469);
nand U4338 (N_4338,N_1650,N_59);
or U4339 (N_4339,N_3649,N_2867);
and U4340 (N_4340,N_473,N_2659);
nand U4341 (N_4341,N_3390,N_445);
xnor U4342 (N_4342,N_110,N_3842);
and U4343 (N_4343,N_3151,N_304);
and U4344 (N_4344,N_2040,N_2764);
or U4345 (N_4345,N_3091,N_1134);
or U4346 (N_4346,N_2746,N_1008);
and U4347 (N_4347,N_807,N_3014);
nand U4348 (N_4348,N_1197,N_2745);
and U4349 (N_4349,N_2707,N_2999);
nand U4350 (N_4350,N_3396,N_236);
or U4351 (N_4351,N_1515,N_63);
nand U4352 (N_4352,N_1798,N_605);
or U4353 (N_4353,N_682,N_3009);
nand U4354 (N_4354,N_3005,N_74);
or U4355 (N_4355,N_1704,N_2169);
or U4356 (N_4356,N_238,N_491);
nor U4357 (N_4357,N_648,N_3490);
nand U4358 (N_4358,N_3952,N_2910);
or U4359 (N_4359,N_1292,N_2332);
and U4360 (N_4360,N_1549,N_1279);
and U4361 (N_4361,N_1890,N_3160);
or U4362 (N_4362,N_2584,N_2538);
nand U4363 (N_4363,N_3444,N_1159);
or U4364 (N_4364,N_1727,N_2509);
xor U4365 (N_4365,N_820,N_3545);
nor U4366 (N_4366,N_3800,N_764);
or U4367 (N_4367,N_43,N_379);
xnor U4368 (N_4368,N_585,N_2750);
xor U4369 (N_4369,N_2835,N_3428);
xnor U4370 (N_4370,N_2747,N_323);
xor U4371 (N_4371,N_232,N_1444);
and U4372 (N_4372,N_1089,N_488);
and U4373 (N_4373,N_1660,N_793);
and U4374 (N_4374,N_912,N_2210);
or U4375 (N_4375,N_3462,N_2690);
or U4376 (N_4376,N_2889,N_1264);
nand U4377 (N_4377,N_2782,N_532);
or U4378 (N_4378,N_3658,N_313);
nand U4379 (N_4379,N_1889,N_3238);
nand U4380 (N_4380,N_3638,N_2384);
or U4381 (N_4381,N_940,N_11);
nor U4382 (N_4382,N_1002,N_3606);
or U4383 (N_4383,N_822,N_2512);
xor U4384 (N_4384,N_176,N_774);
xor U4385 (N_4385,N_3410,N_2285);
xnor U4386 (N_4386,N_3297,N_2026);
nand U4387 (N_4387,N_1471,N_1405);
and U4388 (N_4388,N_2194,N_3964);
xor U4389 (N_4389,N_2141,N_934);
xor U4390 (N_4390,N_2972,N_694);
nor U4391 (N_4391,N_1759,N_1084);
xor U4392 (N_4392,N_651,N_2310);
and U4393 (N_4393,N_1267,N_1654);
nand U4394 (N_4394,N_2725,N_2250);
and U4395 (N_4395,N_1733,N_563);
or U4396 (N_4396,N_2927,N_777);
and U4397 (N_4397,N_2637,N_3018);
xor U4398 (N_4398,N_360,N_100);
and U4399 (N_4399,N_1508,N_2809);
and U4400 (N_4400,N_2472,N_6);
nor U4401 (N_4401,N_3115,N_1692);
or U4402 (N_4402,N_457,N_3474);
xor U4403 (N_4403,N_3938,N_122);
xnor U4404 (N_4404,N_888,N_1370);
nor U4405 (N_4405,N_480,N_1358);
and U4406 (N_4406,N_1477,N_2154);
or U4407 (N_4407,N_146,N_3097);
or U4408 (N_4408,N_3055,N_123);
or U4409 (N_4409,N_3256,N_1274);
nand U4410 (N_4410,N_1686,N_143);
nor U4411 (N_4411,N_2815,N_991);
nand U4412 (N_4412,N_2461,N_1055);
xnor U4413 (N_4413,N_2499,N_2589);
and U4414 (N_4414,N_41,N_65);
nand U4415 (N_4415,N_1468,N_3609);
nand U4416 (N_4416,N_981,N_2163);
xnor U4417 (N_4417,N_219,N_522);
xnor U4418 (N_4418,N_529,N_1703);
or U4419 (N_4419,N_937,N_559);
nand U4420 (N_4420,N_560,N_670);
nand U4421 (N_4421,N_643,N_1957);
xnor U4422 (N_4422,N_2937,N_2858);
xor U4423 (N_4423,N_3431,N_2919);
xor U4424 (N_4424,N_314,N_3807);
nand U4425 (N_4425,N_1118,N_1400);
xnor U4426 (N_4426,N_3194,N_2504);
and U4427 (N_4427,N_1906,N_1298);
nor U4428 (N_4428,N_958,N_3417);
and U4429 (N_4429,N_3686,N_267);
or U4430 (N_4430,N_1120,N_2582);
nor U4431 (N_4431,N_1856,N_2990);
or U4432 (N_4432,N_2488,N_497);
nand U4433 (N_4433,N_3219,N_1491);
xor U4434 (N_4434,N_131,N_1339);
xnor U4435 (N_4435,N_2292,N_1171);
or U4436 (N_4436,N_3273,N_253);
nor U4437 (N_4437,N_1910,N_404);
nand U4438 (N_4438,N_3788,N_3761);
nor U4439 (N_4439,N_3681,N_1050);
and U4440 (N_4440,N_3572,N_291);
nand U4441 (N_4441,N_667,N_1235);
nand U4442 (N_4442,N_2594,N_356);
nand U4443 (N_4443,N_103,N_158);
or U4444 (N_4444,N_3323,N_481);
xor U4445 (N_4445,N_3144,N_3715);
nor U4446 (N_4446,N_3920,N_1038);
xor U4447 (N_4447,N_3697,N_872);
xor U4448 (N_4448,N_2544,N_1342);
nor U4449 (N_4449,N_2306,N_3344);
xor U4450 (N_4450,N_3946,N_3873);
nand U4451 (N_4451,N_3422,N_3822);
nor U4452 (N_4452,N_1852,N_2758);
xor U4453 (N_4453,N_3348,N_867);
nand U4454 (N_4454,N_3656,N_2495);
xnor U4455 (N_4455,N_1679,N_309);
and U4456 (N_4456,N_3518,N_1627);
and U4457 (N_4457,N_464,N_1841);
or U4458 (N_4458,N_1034,N_2009);
xor U4459 (N_4459,N_1716,N_284);
and U4460 (N_4460,N_1000,N_1333);
nand U4461 (N_4461,N_982,N_2348);
xor U4462 (N_4462,N_1814,N_2403);
nor U4463 (N_4463,N_3330,N_863);
and U4464 (N_4464,N_2208,N_860);
nor U4465 (N_4465,N_37,N_1385);
nor U4466 (N_4466,N_1312,N_3890);
or U4467 (N_4467,N_1062,N_2192);
or U4468 (N_4468,N_2452,N_3725);
xor U4469 (N_4469,N_2399,N_1458);
nand U4470 (N_4470,N_3666,N_1882);
xor U4471 (N_4471,N_209,N_2870);
nor U4472 (N_4472,N_3726,N_446);
or U4473 (N_4473,N_3853,N_3026);
or U4474 (N_4474,N_3960,N_3508);
and U4475 (N_4475,N_3202,N_1623);
xnor U4476 (N_4476,N_3530,N_1985);
nand U4477 (N_4477,N_161,N_241);
or U4478 (N_4478,N_2252,N_2450);
or U4479 (N_4479,N_2466,N_13);
nor U4480 (N_4480,N_2082,N_1048);
and U4481 (N_4481,N_2107,N_2409);
nand U4482 (N_4482,N_1911,N_720);
nor U4483 (N_4483,N_2030,N_477);
nor U4484 (N_4484,N_3283,N_503);
and U4485 (N_4485,N_1334,N_3010);
nor U4486 (N_4486,N_82,N_1745);
or U4487 (N_4487,N_102,N_622);
or U4488 (N_4488,N_614,N_744);
nand U4489 (N_4489,N_2804,N_3847);
or U4490 (N_4490,N_695,N_1449);
nor U4491 (N_4491,N_1361,N_2885);
and U4492 (N_4492,N_1473,N_1635);
and U4493 (N_4493,N_435,N_1720);
or U4494 (N_4494,N_936,N_3893);
or U4495 (N_4495,N_1169,N_489);
nand U4496 (N_4496,N_2344,N_759);
nor U4497 (N_4497,N_3146,N_369);
nand U4498 (N_4498,N_2364,N_2128);
nand U4499 (N_4499,N_3439,N_1467);
xnor U4500 (N_4500,N_206,N_1994);
nor U4501 (N_4501,N_3653,N_750);
and U4502 (N_4502,N_1415,N_228);
or U4503 (N_4503,N_172,N_3916);
xor U4504 (N_4504,N_1133,N_2383);
and U4505 (N_4505,N_1886,N_3778);
xor U4506 (N_4506,N_2978,N_3090);
xnor U4507 (N_4507,N_3955,N_3109);
nand U4508 (N_4508,N_2877,N_3701);
and U4509 (N_4509,N_3698,N_1445);
or U4510 (N_4510,N_223,N_1222);
nand U4511 (N_4511,N_1005,N_3749);
or U4512 (N_4512,N_1345,N_448);
xnor U4513 (N_4513,N_3728,N_1407);
or U4514 (N_4514,N_1081,N_2387);
and U4515 (N_4515,N_2926,N_932);
and U4516 (N_4516,N_1109,N_3094);
nand U4517 (N_4517,N_1209,N_525);
nor U4518 (N_4518,N_2426,N_2844);
or U4519 (N_4519,N_2501,N_3298);
xor U4520 (N_4520,N_2078,N_2314);
nand U4521 (N_4521,N_524,N_3624);
xnor U4522 (N_4522,N_1767,N_3875);
nand U4523 (N_4523,N_3659,N_2484);
nand U4524 (N_4524,N_2763,N_2541);
xor U4525 (N_4525,N_2693,N_194);
nor U4526 (N_4526,N_2336,N_1988);
xor U4527 (N_4527,N_2510,N_151);
xnor U4528 (N_4528,N_138,N_99);
and U4529 (N_4529,N_3718,N_23);
nand U4530 (N_4530,N_3834,N_2148);
nor U4531 (N_4531,N_1582,N_663);
and U4532 (N_4532,N_2774,N_3053);
nand U4533 (N_4533,N_2649,N_2261);
nand U4534 (N_4534,N_714,N_3626);
nand U4535 (N_4535,N_293,N_689);
xnor U4536 (N_4536,N_812,N_3343);
nor U4537 (N_4537,N_1850,N_3333);
nor U4538 (N_4538,N_1694,N_3466);
and U4539 (N_4539,N_2881,N_2540);
or U4540 (N_4540,N_3774,N_2120);
nand U4541 (N_4541,N_68,N_2170);
or U4542 (N_4542,N_644,N_2166);
nand U4543 (N_4543,N_2188,N_246);
and U4544 (N_4544,N_2711,N_1229);
and U4545 (N_4545,N_2769,N_1156);
nand U4546 (N_4546,N_1424,N_977);
or U4547 (N_4547,N_2337,N_132);
nor U4548 (N_4548,N_2728,N_145);
nor U4549 (N_4549,N_1313,N_3433);
nor U4550 (N_4550,N_549,N_3898);
and U4551 (N_4551,N_500,N_2316);
xnor U4552 (N_4552,N_1563,N_1888);
and U4553 (N_4553,N_1384,N_3905);
nand U4554 (N_4554,N_3252,N_903);
xor U4555 (N_4555,N_456,N_1085);
xor U4556 (N_4556,N_2458,N_1435);
or U4557 (N_4557,N_2123,N_3337);
nand U4558 (N_4558,N_1666,N_988);
nor U4559 (N_4559,N_3326,N_2975);
xor U4560 (N_4560,N_2174,N_1194);
and U4561 (N_4561,N_3526,N_3375);
xnor U4562 (N_4562,N_2859,N_2035);
or U4563 (N_4563,N_1605,N_1897);
nor U4564 (N_4564,N_1020,N_218);
nand U4565 (N_4565,N_1540,N_838);
xor U4566 (N_4566,N_3771,N_782);
nand U4567 (N_4567,N_75,N_2214);
or U4568 (N_4568,N_3077,N_2621);
or U4569 (N_4569,N_2738,N_3171);
and U4570 (N_4570,N_1123,N_1359);
nor U4571 (N_4571,N_1710,N_1212);
nand U4572 (N_4572,N_337,N_2311);
nor U4573 (N_4573,N_3069,N_2448);
or U4574 (N_4574,N_841,N_1439);
xnor U4575 (N_4575,N_3000,N_3969);
nor U4576 (N_4576,N_2185,N_3046);
xnor U4577 (N_4577,N_548,N_3019);
xor U4578 (N_4578,N_2650,N_364);
nor U4579 (N_4579,N_2679,N_3577);
xor U4580 (N_4580,N_3835,N_1336);
nand U4581 (N_4581,N_3406,N_1629);
nand U4582 (N_4582,N_544,N_3123);
or U4583 (N_4583,N_1523,N_1277);
nand U4584 (N_4584,N_2302,N_1328);
and U4585 (N_4585,N_2801,N_2273);
or U4586 (N_4586,N_1398,N_2439);
nand U4587 (N_4587,N_2539,N_2864);
nand U4588 (N_4588,N_792,N_2346);
xnor U4589 (N_4589,N_2949,N_650);
xor U4590 (N_4590,N_1671,N_1828);
xnor U4591 (N_4591,N_1535,N_271);
xnor U4592 (N_4592,N_3644,N_3472);
nor U4593 (N_4593,N_2159,N_1930);
nand U4594 (N_4594,N_3759,N_2807);
or U4595 (N_4595,N_299,N_3650);
xnor U4596 (N_4596,N_3087,N_3806);
nand U4597 (N_4597,N_2331,N_816);
or U4598 (N_4598,N_2241,N_896);
nor U4599 (N_4599,N_3243,N_160);
or U4600 (N_4600,N_3763,N_788);
or U4601 (N_4601,N_2887,N_879);
xnor U4602 (N_4602,N_2225,N_433);
xnor U4603 (N_4603,N_638,N_2830);
or U4604 (N_4604,N_1700,N_2367);
nand U4605 (N_4605,N_247,N_2146);
nand U4606 (N_4606,N_183,N_1350);
nor U4607 (N_4607,N_3395,N_142);
or U4608 (N_4608,N_2058,N_2464);
nand U4609 (N_4609,N_3949,N_3854);
nor U4610 (N_4610,N_2880,N_2767);
and U4611 (N_4611,N_2404,N_2142);
or U4612 (N_4612,N_2398,N_3732);
nor U4613 (N_4613,N_3279,N_1939);
nand U4614 (N_4614,N_373,N_188);
xnor U4615 (N_4615,N_3667,N_939);
nor U4616 (N_4616,N_3637,N_198);
or U4617 (N_4617,N_2222,N_3251);
and U4618 (N_4618,N_609,N_3370);
or U4619 (N_4619,N_1597,N_3445);
nor U4620 (N_4620,N_635,N_930);
or U4621 (N_4621,N_910,N_2868);
nand U4622 (N_4622,N_1651,N_346);
xnor U4623 (N_4623,N_274,N_2183);
nor U4624 (N_4624,N_2987,N_3615);
xor U4625 (N_4625,N_3557,N_191);
nand U4626 (N_4626,N_3544,N_2229);
nor U4627 (N_4627,N_588,N_2232);
or U4628 (N_4628,N_1663,N_1778);
xor U4629 (N_4629,N_2479,N_3008);
nand U4630 (N_4630,N_2761,N_1615);
nor U4631 (N_4631,N_2161,N_590);
xnor U4632 (N_4632,N_3887,N_2239);
and U4633 (N_4633,N_31,N_2634);
or U4634 (N_4634,N_139,N_3450);
nand U4635 (N_4635,N_3709,N_984);
nand U4636 (N_4636,N_1730,N_1205);
nor U4637 (N_4637,N_3576,N_3951);
or U4638 (N_4638,N_3210,N_1189);
nor U4639 (N_4639,N_1383,N_870);
nor U4640 (N_4640,N_414,N_1302);
and U4641 (N_4641,N_1122,N_1343);
xnor U4642 (N_4642,N_789,N_882);
xor U4643 (N_4643,N_3179,N_2114);
and U4644 (N_4644,N_212,N_453);
nor U4645 (N_4645,N_1958,N_1869);
nand U4646 (N_4646,N_214,N_35);
and U4647 (N_4647,N_848,N_1161);
nor U4648 (N_4648,N_2930,N_3801);
and U4649 (N_4649,N_521,N_2517);
xnor U4650 (N_4650,N_1952,N_2295);
or U4651 (N_4651,N_1634,N_615);
nor U4652 (N_4652,N_1655,N_1951);
or U4653 (N_4653,N_1707,N_885);
nand U4654 (N_4654,N_3742,N_2569);
or U4655 (N_4655,N_3465,N_3232);
and U4656 (N_4656,N_1577,N_1721);
xor U4657 (N_4657,N_1891,N_2977);
and U4658 (N_4658,N_3033,N_974);
nand U4659 (N_4659,N_1711,N_3511);
nand U4660 (N_4660,N_768,N_3876);
nor U4661 (N_4661,N_2943,N_2298);
or U4662 (N_4662,N_849,N_2059);
nor U4663 (N_4663,N_1066,N_1588);
xor U4664 (N_4664,N_386,N_2389);
nor U4665 (N_4665,N_2173,N_2819);
xnor U4666 (N_4666,N_239,N_2296);
xnor U4667 (N_4667,N_1622,N_2668);
and U4668 (N_4668,N_1699,N_2918);
and U4669 (N_4669,N_89,N_1075);
and U4670 (N_4670,N_1807,N_1688);
nand U4671 (N_4671,N_5,N_1054);
and U4672 (N_4672,N_3389,N_2689);
and U4673 (N_4673,N_2655,N_127);
xnor U4674 (N_4674,N_800,N_2493);
or U4675 (N_4675,N_2532,N_878);
xor U4676 (N_4676,N_852,N_392);
xnor U4677 (N_4677,N_3602,N_3195);
nand U4678 (N_4678,N_1029,N_391);
and U4679 (N_4679,N_1499,N_175);
xor U4680 (N_4680,N_2394,N_3001);
nand U4681 (N_4681,N_2895,N_29);
xor U4682 (N_4682,N_1753,N_743);
nand U4683 (N_4683,N_1632,N_2427);
nand U4684 (N_4684,N_3350,N_3329);
and U4685 (N_4685,N_331,N_1774);
nor U4686 (N_4686,N_1137,N_216);
or U4687 (N_4687,N_519,N_3039);
and U4688 (N_4688,N_120,N_2743);
and U4689 (N_4689,N_2793,N_703);
or U4690 (N_4690,N_2015,N_1364);
or U4691 (N_4691,N_1022,N_3863);
and U4692 (N_4692,N_2205,N_2276);
xnor U4693 (N_4693,N_1973,N_2849);
xnor U4694 (N_4694,N_1273,N_1291);
and U4695 (N_4695,N_3549,N_1495);
nand U4696 (N_4696,N_2643,N_2137);
nor U4697 (N_4697,N_3582,N_3909);
or U4698 (N_4698,N_2684,N_1414);
and U4699 (N_4699,N_1461,N_2357);
nor U4700 (N_4700,N_541,N_3430);
xor U4701 (N_4701,N_1785,N_3036);
nand U4702 (N_4702,N_1885,N_2576);
and U4703 (N_4703,N_3028,N_3203);
nand U4704 (N_4704,N_2265,N_2737);
xor U4705 (N_4705,N_2682,N_836);
xor U4706 (N_4706,N_2879,N_1589);
nor U4707 (N_4707,N_3075,N_2244);
nand U4708 (N_4708,N_2395,N_2699);
and U4709 (N_4709,N_2027,N_3588);
and U4710 (N_4710,N_1948,N_1512);
nand U4711 (N_4711,N_2486,N_1044);
xnor U4712 (N_4712,N_2465,N_76);
and U4713 (N_4713,N_3527,N_3536);
or U4714 (N_4714,N_325,N_3215);
nand U4715 (N_4715,N_2720,N_2695);
nor U4716 (N_4716,N_748,N_862);
and U4717 (N_4717,N_390,N_3199);
and U4718 (N_4718,N_254,N_1902);
or U4719 (N_4719,N_245,N_1381);
nand U4720 (N_4720,N_3611,N_722);
or U4721 (N_4721,N_971,N_1490);
nand U4722 (N_4722,N_2884,N_1642);
xor U4723 (N_4723,N_1737,N_1422);
or U4724 (N_4724,N_1154,N_3657);
nor U4725 (N_4725,N_3937,N_2817);
xnor U4726 (N_4726,N_1183,N_1693);
nor U4727 (N_4727,N_2903,N_2139);
nor U4728 (N_4728,N_19,N_2347);
nand U4729 (N_4729,N_1132,N_28);
or U4730 (N_4730,N_2843,N_215);
or U4731 (N_4731,N_3942,N_2382);
xor U4732 (N_4732,N_1714,N_2012);
or U4733 (N_4733,N_2813,N_3132);
nor U4734 (N_4734,N_3468,N_3619);
or U4735 (N_4735,N_3317,N_3394);
nand U4736 (N_4736,N_2586,N_1516);
and U4737 (N_4737,N_3321,N_1324);
or U4738 (N_4738,N_1162,N_3832);
nand U4739 (N_4739,N_2379,N_1970);
and U4740 (N_4740,N_3633,N_3603);
and U4741 (N_4741,N_3663,N_1575);
and U4742 (N_4742,N_803,N_2475);
nand U4743 (N_4743,N_1849,N_3669);
nand U4744 (N_4744,N_3407,N_2511);
nand U4745 (N_4745,N_1861,N_2638);
nand U4746 (N_4746,N_2653,N_3981);
nand U4747 (N_4747,N_2253,N_2266);
nor U4748 (N_4748,N_1497,N_3977);
nor U4749 (N_4749,N_3662,N_1104);
nand U4750 (N_4750,N_3193,N_3073);
and U4751 (N_4751,N_2773,N_451);
xor U4752 (N_4752,N_1511,N_499);
and U4753 (N_4753,N_2983,N_2543);
nand U4754 (N_4754,N_1496,N_3953);
xor U4755 (N_4755,N_2001,N_1868);
and U4756 (N_4756,N_260,N_603);
nand U4757 (N_4757,N_3322,N_1286);
and U4758 (N_4758,N_2941,N_252);
or U4759 (N_4759,N_2626,N_3456);
nand U4760 (N_4760,N_1127,N_747);
or U4761 (N_4761,N_3516,N_2056);
xnor U4762 (N_4762,N_2333,N_1113);
or U4763 (N_4763,N_661,N_1801);
nand U4764 (N_4764,N_978,N_3924);
and U4765 (N_4765,N_3340,N_3382);
nand U4766 (N_4766,N_732,N_352);
nand U4767 (N_4767,N_1744,N_2901);
and U4768 (N_4768,N_3757,N_165);
nand U4769 (N_4769,N_1153,N_2768);
xor U4770 (N_4770,N_989,N_1208);
nand U4771 (N_4771,N_3861,N_225);
xnor U4772 (N_4772,N_1188,N_3803);
xnor U4773 (N_4773,N_1550,N_221);
nand U4774 (N_4774,N_3978,N_1129);
nor U4775 (N_4775,N_771,N_2751);
and U4776 (N_4776,N_2374,N_2048);
xnor U4777 (N_4777,N_3672,N_1028);
nand U4778 (N_4778,N_3524,N_2200);
or U4779 (N_4779,N_2046,N_3436);
or U4780 (N_4780,N_1262,N_2263);
nand U4781 (N_4781,N_1463,N_417);
nor U4782 (N_4782,N_3443,N_332);
nor U4783 (N_4783,N_2017,N_1057);
and U4784 (N_4784,N_2850,N_965);
nor U4785 (N_4785,N_2406,N_2436);
nand U4786 (N_4786,N_1762,N_1546);
nand U4787 (N_4787,N_3758,N_3362);
xor U4788 (N_4788,N_3691,N_3029);
nand U4789 (N_4789,N_349,N_1082);
and U4790 (N_4790,N_1892,N_2726);
or U4791 (N_4791,N_685,N_2549);
or U4792 (N_4792,N_1221,N_3901);
and U4793 (N_4793,N_1943,N_3162);
and U4794 (N_4794,N_2408,N_785);
or U4795 (N_4795,N_370,N_1035);
nor U4796 (N_4796,N_3038,N_728);
nor U4797 (N_4797,N_1033,N_351);
nand U4798 (N_4798,N_1311,N_3336);
nand U4799 (N_4799,N_1844,N_1352);
nor U4800 (N_4800,N_1583,N_45);
nor U4801 (N_4801,N_913,N_205);
or U4802 (N_4802,N_62,N_2661);
and U4803 (N_4803,N_2789,N_2456);
or U4804 (N_4804,N_1317,N_51);
or U4805 (N_4805,N_3403,N_1068);
nand U4806 (N_4806,N_2108,N_1723);
nor U4807 (N_4807,N_3139,N_1176);
or U4808 (N_4808,N_845,N_2121);
nand U4809 (N_4809,N_2605,N_2898);
nand U4810 (N_4810,N_2370,N_3083);
or U4811 (N_4811,N_2973,N_2600);
nand U4812 (N_4812,N_1177,N_249);
or U4813 (N_4813,N_203,N_1232);
or U4814 (N_4814,N_3871,N_1288);
xnor U4815 (N_4815,N_167,N_25);
xor U4816 (N_4816,N_1713,N_1545);
nor U4817 (N_4817,N_2503,N_1503);
and U4818 (N_4818,N_1111,N_3676);
and U4819 (N_4819,N_2050,N_2270);
or U4820 (N_4820,N_2825,N_3480);
and U4821 (N_4821,N_3711,N_2240);
nor U4822 (N_4822,N_834,N_240);
nand U4823 (N_4823,N_3912,N_1480);
xnor U4824 (N_4824,N_2694,N_2313);
xor U4825 (N_4825,N_3296,N_79);
nor U4826 (N_4826,N_2212,N_1344);
nand U4827 (N_4827,N_2443,N_691);
nand U4828 (N_4828,N_2432,N_1392);
nor U4829 (N_4829,N_1604,N_1749);
and U4830 (N_4830,N_1047,N_3086);
and U4831 (N_4831,N_1106,N_3745);
or U4832 (N_4832,N_844,N_3510);
or U4833 (N_4833,N_3963,N_2014);
and U4834 (N_4834,N_766,N_3552);
or U4835 (N_4835,N_2592,N_3302);
and U4836 (N_4836,N_3307,N_292);
xnor U4837 (N_4837,N_947,N_1151);
nor U4838 (N_4838,N_567,N_702);
or U4839 (N_4839,N_3041,N_1078);
or U4840 (N_4840,N_909,N_3921);
or U4841 (N_4841,N_3383,N_3907);
or U4842 (N_4842,N_1898,N_2833);
xnor U4843 (N_4843,N_1025,N_546);
and U4844 (N_4844,N_1417,N_1011);
or U4845 (N_4845,N_857,N_2664);
nand U4846 (N_4846,N_1256,N_2866);
and U4847 (N_4847,N_471,N_2727);
nor U4848 (N_4848,N_2279,N_2368);
nor U4849 (N_4849,N_3043,N_1501);
or U4850 (N_4850,N_1644,N_2172);
nor U4851 (N_4851,N_3288,N_1837);
nor U4852 (N_4852,N_1695,N_3295);
xnor U4853 (N_4853,N_2724,N_528);
and U4854 (N_4854,N_1271,N_3359);
or U4855 (N_4855,N_3277,N_3532);
nand U4856 (N_4856,N_565,N_333);
or U4857 (N_4857,N_547,N_2067);
nand U4858 (N_4858,N_892,N_3274);
and U4859 (N_4859,N_3919,N_3451);
or U4860 (N_4860,N_3995,N_3120);
nor U4861 (N_4861,N_3586,N_853);
nand U4862 (N_4862,N_2784,N_3166);
nor U4863 (N_4863,N_1165,N_16);
xnor U4864 (N_4864,N_1543,N_3531);
nor U4865 (N_4865,N_468,N_114);
nor U4866 (N_4866,N_2157,N_2006);
xor U4867 (N_4867,N_3931,N_855);
nor U4868 (N_4868,N_580,N_2520);
and U4869 (N_4869,N_1116,N_3244);
and U4870 (N_4870,N_681,N_3365);
xor U4871 (N_4871,N_3838,N_3415);
and U4872 (N_4872,N_1284,N_884);
nand U4873 (N_4873,N_3023,N_2607);
nand U4874 (N_4874,N_2102,N_2477);
xor U4875 (N_4875,N_2478,N_893);
xor U4876 (N_4876,N_923,N_2467);
or U4877 (N_4877,N_2896,N_1946);
and U4878 (N_4878,N_1982,N_22);
xor U4879 (N_4879,N_3566,N_2294);
and U4880 (N_4880,N_2583,N_1126);
or U4881 (N_4881,N_3239,N_2032);
and U4882 (N_4882,N_561,N_1032);
and U4883 (N_4883,N_2587,N_1907);
xnor U4884 (N_4884,N_2335,N_2652);
xor U4885 (N_4885,N_2429,N_1083);
xor U4886 (N_4886,N_3032,N_3013);
nand U4887 (N_4887,N_2177,N_318);
nor U4888 (N_4888,N_2829,N_2219);
xnor U4889 (N_4889,N_1587,N_140);
or U4890 (N_4890,N_2388,N_1409);
and U4891 (N_4891,N_1594,N_449);
nor U4892 (N_4892,N_2842,N_1860);
and U4893 (N_4893,N_828,N_80);
nand U4894 (N_4894,N_2714,N_1051);
nor U4895 (N_4895,N_1945,N_1815);
nand U4896 (N_4896,N_1315,N_3188);
nor U4897 (N_4897,N_1842,N_1674);
and U4898 (N_4898,N_1925,N_3727);
xnor U4899 (N_4899,N_2441,N_3319);
and U4900 (N_4900,N_1926,N_1751);
and U4901 (N_4901,N_2221,N_3792);
and U4902 (N_4902,N_1648,N_124);
nand U4903 (N_4903,N_3968,N_125);
xnor U4904 (N_4904,N_2455,N_3722);
xor U4905 (N_4905,N_1238,N_914);
nor U4906 (N_4906,N_3129,N_3802);
and U4907 (N_4907,N_705,N_2994);
nor U4908 (N_4908,N_2095,N_2184);
nor U4909 (N_4909,N_1014,N_36);
xnor U4910 (N_4910,N_3973,N_476);
nor U4911 (N_4911,N_1851,N_2019);
or U4912 (N_4912,N_2152,N_795);
and U4913 (N_4913,N_619,N_773);
xor U4914 (N_4914,N_1128,N_751);
and U4915 (N_4915,N_3292,N_1938);
and U4916 (N_4916,N_3982,N_3983);
nand U4917 (N_4917,N_1100,N_2685);
and U4918 (N_4918,N_3693,N_1337);
nor U4919 (N_4919,N_494,N_576);
and U4920 (N_4920,N_3906,N_533);
or U4921 (N_4921,N_881,N_3453);
xor U4922 (N_4922,N_2491,N_1933);
nand U4923 (N_4923,N_2251,N_2489);
or U4924 (N_4924,N_2948,N_3936);
and U4925 (N_4925,N_3327,N_2770);
or U4926 (N_4926,N_3236,N_14);
or U4927 (N_4927,N_2755,N_2433);
or U4928 (N_4928,N_3173,N_1421);
xor U4929 (N_4929,N_3989,N_1102);
nand U4930 (N_4930,N_1139,N_2481);
and U4931 (N_4931,N_1374,N_1696);
or U4932 (N_4932,N_3652,N_3230);
nand U4933 (N_4933,N_3471,N_1661);
or U4934 (N_4934,N_3299,N_2217);
nand U4935 (N_4935,N_1335,N_1341);
and U4936 (N_4936,N_91,N_1529);
xnor U4937 (N_4937,N_2648,N_815);
or U4938 (N_4938,N_2894,N_2852);
xor U4939 (N_4939,N_3776,N_690);
nor U4940 (N_4940,N_2752,N_2138);
or U4941 (N_4941,N_1072,N_24);
nand U4942 (N_4942,N_3607,N_1164);
and U4943 (N_4943,N_1708,N_1995);
or U4944 (N_4944,N_1469,N_359);
and U4945 (N_4945,N_2899,N_900);
or U4946 (N_4946,N_256,N_1895);
nand U4947 (N_4947,N_3374,N_1017);
or U4948 (N_4948,N_3378,N_3939);
or U4949 (N_4949,N_405,N_2061);
xnor U4950 (N_4950,N_2297,N_2938);
and U4951 (N_4951,N_2326,N_1403);
nand U4952 (N_4952,N_107,N_513);
and U4953 (N_4953,N_3683,N_1726);
or U4954 (N_4954,N_2674,N_2305);
or U4955 (N_4955,N_1838,N_3639);
and U4956 (N_4956,N_1756,N_2736);
nor U4957 (N_4957,N_1631,N_2886);
and U4958 (N_4958,N_1006,N_1514);
nor U4959 (N_4959,N_2838,N_1821);
nand U4960 (N_4960,N_3910,N_2580);
xor U4961 (N_4961,N_3209,N_1036);
xnor U4962 (N_4962,N_1616,N_56);
and U4963 (N_4963,N_1018,N_1318);
xnor U4964 (N_4964,N_3714,N_298);
or U4965 (N_4965,N_3843,N_1007);
xnor U4966 (N_4966,N_231,N_1367);
nor U4967 (N_4967,N_3985,N_811);
nor U4968 (N_4968,N_3539,N_1927);
nand U4969 (N_4969,N_2362,N_3553);
or U4970 (N_4970,N_3980,N_628);
or U4971 (N_4971,N_783,N_311);
xnor U4972 (N_4972,N_2291,N_2748);
and U4973 (N_4973,N_3325,N_3878);
nor U4974 (N_4974,N_150,N_467);
xor U4975 (N_4975,N_517,N_3741);
nor U4976 (N_4976,N_278,N_3712);
nor U4977 (N_4977,N_787,N_1247);
nor U4978 (N_4978,N_2550,N_2639);
nand U4979 (N_4979,N_3849,N_2553);
and U4980 (N_4980,N_3640,N_1272);
nor U4981 (N_4981,N_174,N_1193);
or U4982 (N_4982,N_3216,N_1327);
xor U4983 (N_4983,N_983,N_2775);
and U4984 (N_4984,N_640,N_1791);
and U4985 (N_4985,N_361,N_1776);
and U4986 (N_4986,N_3651,N_3413);
xor U4987 (N_4987,N_2469,N_1031);
and U4988 (N_4988,N_3585,N_1282);
nor U4989 (N_4989,N_199,N_1475);
nor U4990 (N_4990,N_2418,N_2677);
xnor U4991 (N_4991,N_3367,N_2319);
nor U4992 (N_4992,N_2363,N_1278);
nand U4993 (N_4993,N_578,N_3764);
and U4994 (N_4994,N_3419,N_3704);
and U4995 (N_4995,N_3328,N_3491);
nor U4996 (N_4996,N_1308,N_2307);
xor U4997 (N_4997,N_1662,N_2496);
and U4998 (N_4998,N_3270,N_3734);
nand U4999 (N_4999,N_948,N_3357);
or U5000 (N_5000,N_2524,N_1824);
nand U5001 (N_5001,N_904,N_3200);
nor U5002 (N_5002,N_2788,N_3399);
or U5003 (N_5003,N_478,N_1287);
nand U5004 (N_5004,N_1181,N_2802);
or U5005 (N_5005,N_678,N_334);
xor U5006 (N_5006,N_317,N_493);
nand U5007 (N_5007,N_1638,N_2780);
xor U5008 (N_5008,N_3258,N_3694);
nor U5009 (N_5009,N_178,N_1800);
nand U5010 (N_5010,N_2878,N_106);
nand U5011 (N_5011,N_1687,N_2606);
nor U5012 (N_5012,N_1357,N_3956);
nor U5013 (N_5013,N_3519,N_207);
xnor U5014 (N_5014,N_2530,N_3313);
nor U5015 (N_5015,N_184,N_2269);
nor U5016 (N_5016,N_3111,N_2008);
nand U5017 (N_5017,N_1112,N_761);
nor U5018 (N_5018,N_1541,N_831);
or U5019 (N_5019,N_2513,N_504);
or U5020 (N_5020,N_3020,N_2871);
and U5021 (N_5021,N_1532,N_3027);
and U5022 (N_5022,N_53,N_2338);
nor U5023 (N_5023,N_1410,N_1266);
xor U5024 (N_5024,N_3186,N_669);
or U5025 (N_5025,N_3398,N_1981);
nand U5026 (N_5026,N_61,N_3580);
nor U5027 (N_5027,N_2062,N_2907);
nand U5028 (N_5028,N_393,N_3017);
nand U5029 (N_5029,N_1793,N_975);
or U5030 (N_5030,N_552,N_666);
nor U5031 (N_5031,N_2921,N_269);
xor U5032 (N_5032,N_1768,N_746);
nor U5033 (N_5033,N_3988,N_632);
xor U5034 (N_5034,N_3246,N_899);
or U5035 (N_5035,N_3795,N_3844);
nand U5036 (N_5036,N_1709,N_42);
nand U5037 (N_5037,N_3954,N_3756);
or U5038 (N_5038,N_2579,N_2206);
nand U5039 (N_5039,N_115,N_3108);
or U5040 (N_5040,N_3706,N_3054);
xnor U5041 (N_5041,N_3812,N_767);
nand U5042 (N_5042,N_3645,N_3253);
nor U5043 (N_5043,N_1147,N_425);
xor U5044 (N_5044,N_3255,N_3915);
and U5045 (N_5045,N_1369,N_772);
xnor U5046 (N_5046,N_1934,N_1326);
nand U5047 (N_5047,N_1998,N_1346);
nand U5048 (N_5048,N_1777,N_709);
and U5049 (N_5049,N_1299,N_1862);
nor U5050 (N_5050,N_506,N_851);
nand U5051 (N_5051,N_155,N_1457);
xnor U5052 (N_5052,N_3499,N_2361);
nand U5053 (N_5053,N_779,N_2970);
nand U5054 (N_5054,N_2345,N_3829);
nand U5055 (N_5055,N_2662,N_3805);
nand U5056 (N_5056,N_1533,N_2349);
nand U5057 (N_5057,N_2546,N_3356);
or U5058 (N_5058,N_484,N_233);
xor U5059 (N_5059,N_2581,N_1086);
nand U5060 (N_5060,N_3620,N_2041);
xor U5061 (N_5061,N_372,N_1971);
and U5062 (N_5062,N_3719,N_1429);
nor U5063 (N_5063,N_1689,N_970);
or U5064 (N_5064,N_1091,N_507);
or U5065 (N_5065,N_94,N_3057);
or U5066 (N_5066,N_3621,N_1223);
or U5067 (N_5067,N_3908,N_1200);
nor U5068 (N_5068,N_1040,N_1466);
and U5069 (N_5069,N_290,N_1195);
nand U5070 (N_5070,N_3941,N_3459);
xnor U5071 (N_5071,N_3674,N_200);
nand U5072 (N_5072,N_3127,N_3925);
xor U5073 (N_5073,N_2405,N_1799);
and U5074 (N_5074,N_1989,N_3148);
nand U5075 (N_5075,N_2434,N_3064);
nand U5076 (N_5076,N_1734,N_3438);
or U5077 (N_5077,N_3364,N_3904);
xor U5078 (N_5078,N_2356,N_3076);
xnor U5079 (N_5079,N_898,N_3301);
and U5080 (N_5080,N_343,N_1294);
xnor U5081 (N_5081,N_556,N_1395);
nand U5082 (N_5082,N_163,N_1095);
xor U5083 (N_5083,N_439,N_3779);
or U5084 (N_5084,N_620,N_3208);
or U5085 (N_5085,N_1300,N_3781);
and U5086 (N_5086,N_2847,N_2555);
xor U5087 (N_5087,N_821,N_778);
or U5088 (N_5088,N_2112,N_3264);
xnor U5089 (N_5089,N_858,N_2052);
and U5090 (N_5090,N_3735,N_3421);
nand U5091 (N_5091,N_512,N_3733);
and U5092 (N_5092,N_2069,N_3354);
nor U5093 (N_5093,N_3004,N_303);
nor U5094 (N_5094,N_696,N_2974);
nor U5095 (N_5095,N_2615,N_3713);
nand U5096 (N_5096,N_3306,N_1244);
nand U5097 (N_5097,N_3191,N_3868);
nand U5098 (N_5098,N_3229,N_915);
nand U5099 (N_5099,N_721,N_2193);
or U5100 (N_5100,N_2673,N_423);
or U5101 (N_5101,N_1260,N_2260);
nor U5102 (N_5102,N_3930,N_2254);
or U5103 (N_5103,N_3220,N_1773);
nand U5104 (N_5104,N_376,N_3314);
and U5105 (N_5105,N_2732,N_3042);
nor U5106 (N_5106,N_2079,N_2482);
nor U5107 (N_5107,N_169,N_217);
nand U5108 (N_5108,N_3700,N_1297);
nor U5109 (N_5109,N_263,N_3373);
xnor U5110 (N_5110,N_2598,N_2617);
and U5111 (N_5111,N_1618,N_3289);
nand U5112 (N_5112,N_2785,N_1452);
or U5113 (N_5113,N_1735,N_3482);
nor U5114 (N_5114,N_2417,N_551);
or U5115 (N_5115,N_780,N_1626);
or U5116 (N_5116,N_734,N_1936);
nand U5117 (N_5117,N_2189,N_154);
nand U5118 (N_5118,N_1561,N_8);
nand U5119 (N_5119,N_2023,N_2924);
or U5120 (N_5120,N_1301,N_3855);
xnor U5121 (N_5121,N_2564,N_301);
nand U5122 (N_5122,N_624,N_2940);
or U5123 (N_5123,N_1349,N_3928);
or U5124 (N_5124,N_986,N_2915);
xor U5125 (N_5125,N_686,N_1770);
nand U5126 (N_5126,N_2740,N_3493);
or U5127 (N_5127,N_1325,N_2669);
and U5128 (N_5128,N_2960,N_60);
xor U5129 (N_5129,N_1431,N_955);
nand U5130 (N_5130,N_1121,N_1918);
or U5131 (N_5131,N_2928,N_1220);
and U5132 (N_5132,N_3992,N_2303);
nand U5133 (N_5133,N_1460,N_2686);
nand U5134 (N_5134,N_1937,N_1609);
or U5135 (N_5135,N_3226,N_96);
and U5136 (N_5136,N_2739,N_2474);
and U5137 (N_5137,N_911,N_2149);
and U5138 (N_5138,N_842,N_2578);
xnor U5139 (N_5139,N_3775,N_2321);
xnor U5140 (N_5140,N_2097,N_964);
and U5141 (N_5141,N_3754,N_656);
or U5142 (N_5142,N_1520,N_1250);
or U5143 (N_5143,N_1572,N_2526);
nand U5144 (N_5144,N_752,N_465);
xnor U5145 (N_5145,N_2323,N_3494);
nor U5146 (N_5146,N_2109,N_3688);
xor U5147 (N_5147,N_617,N_3845);
nor U5148 (N_5148,N_3804,N_833);
nand U5149 (N_5149,N_3670,N_2435);
nor U5150 (N_5150,N_920,N_2315);
or U5151 (N_5151,N_3797,N_864);
nand U5152 (N_5152,N_3836,N_2106);
and U5153 (N_5153,N_3025,N_3476);
or U5154 (N_5154,N_234,N_407);
xnor U5155 (N_5155,N_3172,N_3839);
xnor U5156 (N_5156,N_3975,N_1795);
nor U5157 (N_5157,N_3710,N_3007);
or U5158 (N_5158,N_3523,N_415);
or U5159 (N_5159,N_3587,N_2920);
xnor U5160 (N_5160,N_389,N_1914);
nand U5161 (N_5161,N_1697,N_280);
nand U5162 (N_5162,N_339,N_660);
or U5163 (N_5163,N_3567,N_459);
or U5164 (N_5164,N_2700,N_3550);
nand U5165 (N_5165,N_944,N_3502);
and U5166 (N_5166,N_3442,N_805);
xor U5167 (N_5167,N_3124,N_3248);
or U5168 (N_5168,N_2293,N_429);
or U5169 (N_5169,N_3892,N_584);
nand U5170 (N_5170,N_3555,N_3414);
nand U5171 (N_5171,N_1438,N_3957);
nand U5172 (N_5172,N_2534,N_3994);
xor U5173 (N_5173,N_1557,N_3458);
nand U5174 (N_5174,N_2156,N_3563);
xnor U5175 (N_5175,N_1619,N_1509);
nor U5176 (N_5176,N_587,N_1476);
and U5177 (N_5177,N_2372,N_1804);
or U5178 (N_5178,N_634,N_3630);
or U5179 (N_5179,N_358,N_2862);
xor U5180 (N_5180,N_2860,N_724);
nor U5181 (N_5181,N_2235,N_3770);
nor U5182 (N_5182,N_3884,N_2492);
or U5183 (N_5183,N_3543,N_321);
and U5184 (N_5184,N_3093,N_1879);
or U5185 (N_5185,N_725,N_3629);
nor U5186 (N_5186,N_3254,N_2256);
nor U5187 (N_5187,N_2982,N_2721);
or U5188 (N_5188,N_1553,N_1268);
and U5189 (N_5189,N_97,N_2585);
nand U5190 (N_5190,N_1489,N_202);
nor U5191 (N_5191,N_208,N_1275);
nand U5192 (N_5192,N_2863,N_3962);
nor U5193 (N_5193,N_866,N_952);
nor U5194 (N_5194,N_3738,N_2971);
and U5195 (N_5195,N_1691,N_455);
xor U5196 (N_5196,N_665,N_606);
or U5197 (N_5197,N_1991,N_1419);
and U5198 (N_5198,N_116,N_3827);
or U5199 (N_5199,N_1178,N_368);
and U5200 (N_5200,N_2986,N_3568);
and U5201 (N_5201,N_113,N_1932);
xnor U5202 (N_5202,N_1389,N_2110);
and U5203 (N_5203,N_3604,N_490);
nand U5204 (N_5204,N_3412,N_383);
xnor U5205 (N_5205,N_3241,N_3554);
nor U5206 (N_5206,N_21,N_1255);
or U5207 (N_5207,N_680,N_3596);
nor U5208 (N_5208,N_2518,N_1873);
nand U5209 (N_5209,N_3409,N_1746);
or U5210 (N_5210,N_2730,N_2856);
or U5211 (N_5211,N_3169,N_1428);
and U5212 (N_5212,N_3813,N_3135);
and U5213 (N_5213,N_1305,N_539);
and U5214 (N_5214,N_2136,N_1853);
nor U5215 (N_5215,N_2075,N_1782);
and U5216 (N_5216,N_3338,N_2045);
nand U5217 (N_5217,N_2084,N_1966);
nor U5218 (N_5218,N_3675,N_1464);
and U5219 (N_5219,N_3628,N_1027);
xor U5220 (N_5220,N_1775,N_2220);
nand U5221 (N_5221,N_1916,N_906);
or U5222 (N_5222,N_3432,N_2281);
xnor U5223 (N_5223,N_1004,N_3121);
nand U5224 (N_5224,N_3379,N_326);
nand U5225 (N_5225,N_1967,N_1672);
xor U5226 (N_5226,N_2153,N_2646);
nand U5227 (N_5227,N_1049,N_718);
or U5228 (N_5228,N_2228,N_437);
nand U5229 (N_5229,N_1340,N_1015);
xor U5230 (N_5230,N_1574,N_531);
and U5231 (N_5231,N_3818,N_1820);
nor U5232 (N_5232,N_2445,N_2487);
nor U5233 (N_5233,N_2759,N_2691);
nor U5234 (N_5234,N_1754,N_2523);
nand U5235 (N_5235,N_3152,N_3037);
nor U5236 (N_5236,N_1353,N_1314);
xnor U5237 (N_5237,N_735,N_1060);
and U5238 (N_5238,N_257,N_1955);
nand U5239 (N_5239,N_69,N_2946);
and U5240 (N_5240,N_2203,N_1070);
and U5241 (N_5241,N_450,N_3040);
nand U5242 (N_5242,N_1962,N_1234);
nor U5243 (N_5243,N_3161,N_636);
xor U5244 (N_5244,N_1368,N_2416);
and U5245 (N_5245,N_1167,N_642);
nand U5246 (N_5246,N_3896,N_308);
nor U5247 (N_5247,N_1864,N_901);
nand U5248 (N_5248,N_1281,N_738);
or U5249 (N_5249,N_943,N_441);
or U5250 (N_5250,N_2355,N_2944);
nand U5251 (N_5251,N_1203,N_2330);
nor U5252 (N_5252,N_1528,N_600);
xor U5253 (N_5253,N_3049,N_73);
and U5254 (N_5254,N_3503,N_3104);
or U5255 (N_5255,N_2618,N_403);
xnor U5256 (N_5256,N_2044,N_1114);
xnor U5257 (N_5257,N_1760,N_1243);
or U5258 (N_5258,N_3300,N_1739);
or U5259 (N_5259,N_595,N_3966);
nor U5260 (N_5260,N_2603,N_2670);
xnor U5261 (N_5261,N_3534,N_454);
or U5262 (N_5262,N_657,N_758);
xnor U5263 (N_5263,N_1092,N_2176);
or U5264 (N_5264,N_2535,N_2089);
xnor U5265 (N_5265,N_1192,N_1196);
xnor U5266 (N_5266,N_466,N_1706);
xor U5267 (N_5267,N_1664,N_2628);
or U5268 (N_5268,N_1810,N_3537);
and U5269 (N_5269,N_3696,N_868);
nand U5270 (N_5270,N_1135,N_3271);
and U5271 (N_5271,N_2380,N_1796);
nor U5272 (N_5272,N_3045,N_3355);
and U5273 (N_5273,N_2566,N_1283);
xnor U5274 (N_5274,N_2985,N_2893);
and U5275 (N_5275,N_3467,N_2181);
nor U5276 (N_5276,N_2397,N_3231);
xor U5277 (N_5277,N_2645,N_3750);
nand U5278 (N_5278,N_604,N_3311);
xor U5279 (N_5279,N_3341,N_3212);
nand U5280 (N_5280,N_2334,N_341);
or U5281 (N_5281,N_1825,N_1974);
nor U5282 (N_5282,N_385,N_545);
nand U5283 (N_5283,N_1747,N_629);
nor U5284 (N_5284,N_889,N_922);
and U5285 (N_5285,N_1625,N_526);
or U5286 (N_5286,N_432,N_3360);
xor U5287 (N_5287,N_1479,N_1573);
xnor U5288 (N_5288,N_664,N_78);
and U5289 (N_5289,N_1603,N_2556);
or U5290 (N_5290,N_83,N_2);
nor U5291 (N_5291,N_1668,N_3048);
xor U5292 (N_5292,N_3852,N_7);
nand U5293 (N_5293,N_1915,N_2998);
and U5294 (N_5294,N_3489,N_3885);
xor U5295 (N_5295,N_2289,N_731);
or U5296 (N_5296,N_2473,N_1763);
and U5297 (N_5297,N_2735,N_2274);
or U5298 (N_5298,N_3768,N_2060);
nand U5299 (N_5299,N_1617,N_2402);
nand U5300 (N_5300,N_3967,N_2421);
xor U5301 (N_5301,N_1446,N_2989);
and U5302 (N_5302,N_1872,N_1026);
xnor U5303 (N_5303,N_1413,N_1309);
xor U5304 (N_5304,N_374,N_1119);
xor U5305 (N_5305,N_1242,N_3724);
nand U5306 (N_5306,N_951,N_3739);
or U5307 (N_5307,N_3247,N_1613);
xnor U5308 (N_5308,N_1101,N_3533);
nand U5309 (N_5309,N_447,N_1909);
nor U5310 (N_5310,N_1580,N_1107);
and U5311 (N_5311,N_1493,N_2290);
nand U5312 (N_5312,N_1527,N_3581);
nor U5313 (N_5313,N_2563,N_2954);
and U5314 (N_5314,N_1752,N_182);
and U5315 (N_5315,N_2401,N_2547);
and U5316 (N_5316,N_472,N_1202);
xor U5317 (N_5317,N_2224,N_1858);
and U5318 (N_5318,N_1157,N_3263);
and U5319 (N_5319,N_3610,N_3051);
nor U5320 (N_5320,N_3664,N_961);
or U5321 (N_5321,N_1965,N_566);
nor U5322 (N_5322,N_1094,N_540);
xor U5323 (N_5323,N_2831,N_2676);
nor U5324 (N_5324,N_2340,N_3371);
xor U5325 (N_5325,N_2528,N_1507);
nor U5326 (N_5326,N_3234,N_1319);
nand U5327 (N_5327,N_112,N_2900);
nand U5328 (N_5328,N_2622,N_1430);
nor U5329 (N_5329,N_3857,N_711);
nand U5330 (N_5330,N_81,N_1596);
nor U5331 (N_5331,N_826,N_631);
nor U5332 (N_5332,N_2620,N_1064);
xor U5333 (N_5333,N_3187,N_222);
nor U5334 (N_5334,N_2821,N_1788);
nand U5335 (N_5335,N_3874,N_2449);
and U5336 (N_5336,N_3137,N_3612);
and U5337 (N_5337,N_2234,N_3595);
and U5338 (N_5338,N_2080,N_3125);
and U5339 (N_5339,N_283,N_3159);
nor U5340 (N_5340,N_2460,N_1959);
nor U5341 (N_5341,N_378,N_1950);
nand U5342 (N_5342,N_3851,N_2494);
or U5343 (N_5343,N_1867,N_3648);
or U5344 (N_5344,N_2094,N_1170);
nand U5345 (N_5345,N_602,N_3492);
and U5346 (N_5346,N_1972,N_594);
and U5347 (N_5347,N_1599,N_1987);
nand U5348 (N_5348,N_3457,N_3575);
or U5349 (N_5349,N_164,N_3594);
nand U5350 (N_5350,N_3540,N_2029);
and U5351 (N_5351,N_2671,N_2020);
xnor U5352 (N_5352,N_1537,N_2570);
nand U5353 (N_5353,N_1524,N_2160);
xnor U5354 (N_5354,N_741,N_162);
nor U5355 (N_5355,N_2425,N_2053);
and U5356 (N_5356,N_52,N_1715);
or U5357 (N_5357,N_993,N_1877);
or U5358 (N_5358,N_1865,N_2390);
nor U5359 (N_5359,N_2471,N_1079);
xor U5360 (N_5360,N_2931,N_3034);
nand U5361 (N_5361,N_2320,N_2021);
xor U5362 (N_5362,N_1377,N_924);
or U5363 (N_5363,N_804,N_93);
and U5364 (N_5364,N_3974,N_3679);
or U5365 (N_5365,N_1665,N_2271);
and U5366 (N_5366,N_384,N_1725);
xnor U5367 (N_5367,N_134,N_3122);
nor U5368 (N_5368,N_684,N_2665);
nor U5369 (N_5369,N_1185,N_941);
or U5370 (N_5370,N_2678,N_3079);
nor U5371 (N_5371,N_3425,N_312);
or U5372 (N_5372,N_1544,N_2396);
nor U5373 (N_5373,N_796,N_523);
nor U5374 (N_5374,N_2190,N_272);
nor U5375 (N_5375,N_1241,N_1978);
nor U5376 (N_5376,N_1237,N_12);
xor U5377 (N_5377,N_1184,N_3278);
or U5378 (N_5378,N_1712,N_277);
nor U5379 (N_5379,N_3265,N_1391);
xnor U5380 (N_5380,N_2966,N_2988);
and U5381 (N_5381,N_2791,N_3998);
nand U5382 (N_5382,N_2786,N_2360);
and U5383 (N_5383,N_2037,N_3068);
or U5384 (N_5384,N_3866,N_3178);
nor U5385 (N_5385,N_2548,N_462);
nand U5386 (N_5386,N_1789,N_1433);
nor U5387 (N_5387,N_2805,N_1992);
nand U5388 (N_5388,N_3405,N_2613);
nor U5389 (N_5389,N_2573,N_3100);
and U5390 (N_5390,N_2171,N_749);
or U5391 (N_5391,N_3837,N_3961);
and U5392 (N_5392,N_344,N_3535);
and U5393 (N_5393,N_1568,N_1649);
and U5394 (N_5394,N_3627,N_798);
xor U5395 (N_5395,N_646,N_2371);
nor U5396 (N_5396,N_2667,N_3591);
or U5397 (N_5397,N_1757,N_3560);
or U5398 (N_5398,N_2342,N_1338);
or U5399 (N_5399,N_3349,N_3175);
or U5400 (N_5400,N_2647,N_1667);
nand U5401 (N_5401,N_2485,N_1637);
nor U5402 (N_5402,N_1138,N_2158);
xnor U5403 (N_5403,N_2198,N_1024);
or U5404 (N_5404,N_1698,N_248);
nand U5405 (N_5405,N_869,N_3702);
nand U5406 (N_5406,N_2729,N_3222);
and U5407 (N_5407,N_784,N_3565);
and U5408 (N_5408,N_3848,N_3986);
or U5409 (N_5409,N_570,N_322);
nor U5410 (N_5410,N_1569,N_3381);
xor U5411 (N_5411,N_2187,N_3282);
nand U5412 (N_5412,N_3926,N_1426);
and U5413 (N_5413,N_409,N_1166);
xnor U5414 (N_5414,N_1427,N_3708);
nor U5415 (N_5415,N_1141,N_2632);
nand U5416 (N_5416,N_297,N_88);
and U5417 (N_5417,N_2016,N_2010);
xor U5418 (N_5418,N_1765,N_2624);
nand U5419 (N_5419,N_2201,N_2378);
and U5420 (N_5420,N_3665,N_3705);
nand U5421 (N_5421,N_1440,N_475);
nor U5422 (N_5422,N_3488,N_3030);
or U5423 (N_5423,N_3067,N_2837);
and U5424 (N_5424,N_1857,N_1806);
nand U5425 (N_5425,N_2376,N_1809);
nor U5426 (N_5426,N_2609,N_1633);
nor U5427 (N_5427,N_3165,N_502);
nand U5428 (N_5428,N_85,N_2018);
nand U5429 (N_5429,N_2968,N_3881);
xnor U5430 (N_5430,N_712,N_824);
xor U5431 (N_5431,N_3334,N_3228);
xnor U5432 (N_5432,N_3142,N_1434);
xnor U5433 (N_5433,N_86,N_408);
and U5434 (N_5434,N_1251,N_2309);
and U5435 (N_5435,N_514,N_1819);
xor U5436 (N_5436,N_2118,N_1921);
nand U5437 (N_5437,N_3149,N_1984);
or U5438 (N_5438,N_3154,N_2660);
xor U5439 (N_5439,N_727,N_3291);
or U5440 (N_5440,N_520,N_1348);
xnor U5441 (N_5441,N_3446,N_2717);
xor U5442 (N_5442,N_618,N_3731);
nand U5443 (N_5443,N_3773,N_933);
or U5444 (N_5444,N_2231,N_3106);
and U5445 (N_5445,N_3831,N_2716);
xor U5446 (N_5446,N_2818,N_1447);
nor U5447 (N_5447,N_2103,N_2386);
or U5448 (N_5448,N_501,N_1779);
xnor U5449 (N_5449,N_518,N_220);
and U5450 (N_5450,N_3143,N_20);
or U5451 (N_5451,N_1140,N_3024);
and U5452 (N_5452,N_3548,N_1365);
or U5453 (N_5453,N_2808,N_553);
nor U5454 (N_5454,N_3276,N_197);
nor U5455 (N_5455,N_3720,N_3571);
or U5456 (N_5456,N_3551,N_1149);
and U5457 (N_5457,N_2914,N_2562);
nor U5458 (N_5458,N_2554,N_2413);
or U5459 (N_5459,N_1105,N_483);
nor U5460 (N_5460,N_2681,N_2216);
and U5461 (N_5461,N_1586,N_2391);
nand U5462 (N_5462,N_2414,N_3424);
xor U5463 (N_5463,N_306,N_2827);
nor U5464 (N_5464,N_1736,N_302);
nand U5465 (N_5465,N_1213,N_2131);
nand U5466 (N_5466,N_1163,N_802);
or U5467 (N_5467,N_2129,N_2140);
or U5468 (N_5468,N_3655,N_168);
xor U5469 (N_5469,N_555,N_2719);
and U5470 (N_5470,N_536,N_2151);
nand U5471 (N_5471,N_883,N_3065);
xnor U5472 (N_5472,N_1486,N_3772);
xnor U5473 (N_5473,N_2875,N_3786);
and U5474 (N_5474,N_430,N_1980);
or U5475 (N_5475,N_1443,N_992);
nor U5476 (N_5476,N_840,N_2781);
nor U5477 (N_5477,N_973,N_1206);
nor U5478 (N_5478,N_1270,N_675);
xor U5479 (N_5479,N_1379,N_1155);
or U5480 (N_5480,N_994,N_3970);
xnor U5481 (N_5481,N_2113,N_739);
and U5482 (N_5482,N_181,N_3914);
or U5483 (N_5483,N_2908,N_3335);
and U5484 (N_5484,N_2568,N_2558);
nor U5485 (N_5485,N_1701,N_2168);
and U5486 (N_5486,N_95,N_418);
xnor U5487 (N_5487,N_3976,N_573);
nor U5488 (N_5488,N_699,N_2577);
or U5489 (N_5489,N_3799,N_262);
nor U5490 (N_5490,N_3189,N_3204);
nand U5491 (N_5491,N_1792,N_3437);
or U5492 (N_5492,N_2377,N_3520);
nand U5493 (N_5493,N_1610,N_3987);
or U5494 (N_5494,N_2447,N_2992);
or U5495 (N_5495,N_1551,N_3114);
or U5496 (N_5496,N_1416,N_3808);
nor U5497 (N_5497,N_2552,N_104);
nor U5498 (N_5498,N_2280,N_157);
nand U5499 (N_5499,N_976,N_1831);
and U5500 (N_5500,N_3811,N_431);
nor U5501 (N_5501,N_1451,N_575);
and U5502 (N_5502,N_918,N_50);
and U5503 (N_5503,N_1399,N_3119);
xnor U5504 (N_5504,N_610,N_1990);
xnor U5505 (N_5505,N_2672,N_2352);
xnor U5506 (N_5506,N_1827,N_2779);
xnor U5507 (N_5507,N_2096,N_1817);
xor U5508 (N_5508,N_2611,N_2242);
xnor U5509 (N_5509,N_2328,N_3163);
nand U5510 (N_5510,N_1640,N_1394);
xor U5511 (N_5511,N_3388,N_3351);
nand U5512 (N_5512,N_515,N_1401);
nor U5513 (N_5513,N_2876,N_2438);
xnor U5514 (N_5514,N_1390,N_2527);
nor U5515 (N_5515,N_1584,N_2508);
or U5516 (N_5516,N_508,N_380);
and U5517 (N_5517,N_658,N_295);
and U5518 (N_5518,N_347,N_2516);
nand U5519 (N_5519,N_1393,N_261);
and U5520 (N_5520,N_2226,N_2641);
nor U5521 (N_5521,N_3486,N_1880);
xnor U5522 (N_5522,N_3950,N_2424);
nand U5523 (N_5523,N_3085,N_2962);
nor U5524 (N_5524,N_211,N_1769);
and U5525 (N_5525,N_3418,N_2874);
or U5526 (N_5526,N_2223,N_1290);
nand U5527 (N_5527,N_850,N_2828);
xor U5528 (N_5528,N_1332,N_2519);
xor U5529 (N_5529,N_1956,N_1802);
nand U5530 (N_5530,N_3082,N_3434);
nand U5531 (N_5531,N_1382,N_2658);
and U5532 (N_5532,N_3793,N_1146);
xnor U5533 (N_5533,N_3578,N_3136);
or U5534 (N_5534,N_1823,N_1976);
or U5535 (N_5535,N_2760,N_1787);
or U5536 (N_5536,N_3448,N_1614);
and U5537 (N_5537,N_630,N_908);
nor U5538 (N_5538,N_3895,N_1240);
nor U5539 (N_5539,N_3707,N_3475);
and U5540 (N_5540,N_3971,N_1215);
xor U5541 (N_5541,N_3897,N_2440);
and U5542 (N_5542,N_1743,N_1812);
and U5543 (N_5543,N_1245,N_2500);
nand U5544 (N_5544,N_611,N_962);
and U5545 (N_5545,N_3911,N_3056);
or U5546 (N_5546,N_3505,N_808);
xnor U5547 (N_5547,N_3542,N_2934);
nor U5548 (N_5548,N_1187,N_706);
xor U5549 (N_5549,N_2599,N_1174);
nor U5550 (N_5550,N_315,N_2533);
or U5551 (N_5551,N_1670,N_2351);
and U5552 (N_5552,N_2230,N_3605);
or U5553 (N_5553,N_66,N_3660);
xnor U5554 (N_5554,N_237,N_3997);
xnor U5555 (N_5555,N_1248,N_1303);
nand U5556 (N_5556,N_612,N_39);
nor U5557 (N_5557,N_3201,N_3110);
nor U5558 (N_5558,N_2167,N_3176);
nand U5559 (N_5559,N_3280,N_1983);
nor U5560 (N_5560,N_156,N_3635);
nand U5561 (N_5561,N_3541,N_1908);
nor U5562 (N_5562,N_3070,N_1521);
nand U5563 (N_5563,N_2955,N_980);
xnor U5564 (N_5564,N_470,N_577);
xor U5565 (N_5565,N_786,N_972);
nor U5566 (N_5566,N_348,N_44);
and U5567 (N_5567,N_760,N_1459);
nor U5568 (N_5568,N_3310,N_3867);
nor U5569 (N_5569,N_3225,N_141);
and U5570 (N_5570,N_3346,N_3979);
nand U5571 (N_5571,N_3929,N_2446);
nand U5572 (N_5572,N_2304,N_598);
xor U5573 (N_5573,N_3760,N_3294);
and U5574 (N_5574,N_775,N_1526);
nor U5575 (N_5575,N_3685,N_2049);
nand U5576 (N_5576,N_1355,N_281);
nor U5577 (N_5577,N_126,N_674);
and U5578 (N_5578,N_2071,N_3116);
xor U5579 (N_5579,N_1997,N_1875);
and U5580 (N_5580,N_873,N_3366);
nand U5581 (N_5581,N_2551,N_574);
nand U5582 (N_5582,N_2237,N_193);
xnor U5583 (N_5583,N_357,N_2964);
nor U5584 (N_5584,N_1904,N_3332);
nand U5585 (N_5585,N_2490,N_2451);
nand U5586 (N_5586,N_997,N_492);
or U5587 (N_5587,N_320,N_2422);
or U5588 (N_5588,N_1718,N_715);
nand U5589 (N_5589,N_1423,N_2258);
nor U5590 (N_5590,N_2545,N_49);
nor U5591 (N_5591,N_2892,N_537);
nor U5592 (N_5592,N_813,N_2950);
or U5593 (N_5593,N_3958,N_1217);
or U5594 (N_5594,N_2942,N_1378);
or U5595 (N_5595,N_90,N_3285);
or U5596 (N_5596,N_1928,N_3497);
nand U5597 (N_5597,N_1080,N_2442);
xor U5598 (N_5598,N_754,N_1117);
xor U5599 (N_5599,N_1453,N_1608);
xor U5600 (N_5600,N_1834,N_1474);
nand U5601 (N_5601,N_3558,N_1214);
and U5602 (N_5602,N_832,N_3331);
nor U5603 (N_5603,N_1039,N_130);
and U5604 (N_5604,N_3324,N_2359);
nand U5605 (N_5605,N_2195,N_2430);
or U5606 (N_5606,N_1418,N_3242);
or U5607 (N_5607,N_755,N_2904);
or U5608 (N_5608,N_3622,N_3883);
nor U5609 (N_5609,N_2811,N_1099);
xnor U5610 (N_5610,N_1069,N_1894);
and U5611 (N_5611,N_2087,N_3882);
or U5612 (N_5612,N_3559,N_1878);
nand U5613 (N_5613,N_2836,N_3744);
nor U5614 (N_5614,N_593,N_3267);
nand U5615 (N_5615,N_2703,N_1420);
nand U5616 (N_5616,N_2468,N_1347);
nor U5617 (N_5617,N_1652,N_276);
and U5618 (N_5618,N_436,N_2963);
xor U5619 (N_5619,N_2571,N_1624);
xnor U5620 (N_5620,N_3245,N_3787);
or U5621 (N_5621,N_1600,N_554);
or U5622 (N_5622,N_707,N_1598);
and U5623 (N_5623,N_1783,N_564);
xor U5624 (N_5624,N_1636,N_985);
and U5625 (N_5625,N_1639,N_1160);
nand U5626 (N_5626,N_1462,N_1729);
or U5627 (N_5627,N_1560,N_3447);
nor U5628 (N_5628,N_733,N_2772);
nor U5629 (N_5629,N_1492,N_2104);
nand U5630 (N_5630,N_3180,N_3783);
xor U5631 (N_5631,N_829,N_3830);
xor U5632 (N_5632,N_1808,N_77);
nand U5633 (N_5633,N_3477,N_1630);
nand U5634 (N_5634,N_1830,N_817);
xnor U5635 (N_5635,N_2207,N_46);
nor U5636 (N_5636,N_1304,N_2028);
xor U5637 (N_5637,N_486,N_3305);
nor U5638 (N_5638,N_2602,N_1829);
or U5639 (N_5639,N_3449,N_3031);
and U5640 (N_5640,N_1172,N_3006);
or U5641 (N_5641,N_3003,N_2299);
nor U5642 (N_5642,N_3303,N_3227);
nor U5643 (N_5643,N_1750,N_2116);
or U5644 (N_5644,N_1690,N_2851);
or U5645 (N_5645,N_2134,N_3016);
nor U5646 (N_5646,N_723,N_1602);
or U5647 (N_5647,N_3514,N_2083);
or U5648 (N_5648,N_3922,N_776);
xor U5649 (N_5649,N_1530,N_375);
nand U5650 (N_5650,N_30,N_3429);
or U5651 (N_5651,N_3833,N_1042);
or U5652 (N_5652,N_679,N_2984);
and U5653 (N_5653,N_1498,N_171);
nand U5654 (N_5654,N_1320,N_1786);
nor U5655 (N_5655,N_967,N_1484);
and U5656 (N_5656,N_2909,N_1628);
nand U5657 (N_5657,N_1731,N_3316);
xor U5658 (N_5658,N_1607,N_3304);
xor U5659 (N_5659,N_1087,N_3614);
nor U5660 (N_5660,N_3767,N_268);
and U5661 (N_5661,N_3743,N_1030);
xor U5662 (N_5662,N_3647,N_1239);
xor U5663 (N_5663,N_639,N_3483);
or U5664 (N_5664,N_1859,N_55);
nand U5665 (N_5665,N_625,N_926);
nand U5666 (N_5666,N_916,N_2593);
xnor U5667 (N_5667,N_1811,N_3654);
nor U5668 (N_5668,N_153,N_2126);
and U5669 (N_5669,N_3872,N_3372);
and U5670 (N_5670,N_716,N_3751);
nor U5671 (N_5671,N_2522,N_3680);
xnor U5672 (N_5672,N_3798,N_3522);
xnor U5673 (N_5673,N_1917,N_2945);
nand U5674 (N_5674,N_835,N_3308);
nand U5675 (N_5675,N_2324,N_458);
nor U5676 (N_5676,N_1941,N_698);
nand U5677 (N_5677,N_623,N_2916);
or U5678 (N_5678,N_3826,N_1896);
and U5679 (N_5679,N_730,N_353);
xnor U5680 (N_5680,N_2561,N_2757);
and U5681 (N_5681,N_363,N_336);
nand U5682 (N_5682,N_1740,N_3864);
xor U5683 (N_5683,N_1373,N_3846);
and U5684 (N_5684,N_814,N_3423);
or U5685 (N_5685,N_367,N_2702);
or U5686 (N_5686,N_1173,N_1265);
or U5687 (N_5687,N_2980,N_1534);
xor U5688 (N_5688,N_1536,N_3363);
or U5689 (N_5689,N_3011,N_1093);
nor U5690 (N_5690,N_2022,N_647);
nand U5691 (N_5691,N_2905,N_1702);
nor U5692 (N_5692,N_2150,N_3525);
nand U5693 (N_5693,N_1839,N_2033);
or U5694 (N_5694,N_2614,N_3126);
xnor U5695 (N_5695,N_1518,N_2375);
nand U5696 (N_5696,N_1354,N_2282);
and U5697 (N_5697,N_0,N_460);
or U5698 (N_5698,N_2215,N_1678);
and U5699 (N_5699,N_2462,N_2124);
and U5700 (N_5700,N_1257,N_3315);
xnor U5701 (N_5701,N_3376,N_1502);
xor U5702 (N_5702,N_2264,N_1481);
nand U5703 (N_5703,N_2803,N_1576);
and U5704 (N_5704,N_880,N_3940);
nor U5705 (N_5705,N_3454,N_1142);
or U5706 (N_5706,N_362,N_2619);
xor U5707 (N_5707,N_3150,N_2687);
xnor U5708 (N_5708,N_1225,N_2959);
nor U5709 (N_5709,N_3755,N_1432);
nor U5710 (N_5710,N_2327,N_3877);
xor U5711 (N_5711,N_1996,N_3894);
nor U5712 (N_5712,N_654,N_2175);
nor U5713 (N_5713,N_2300,N_1258);
nor U5714 (N_5714,N_950,N_2967);
nor U5715 (N_5715,N_2246,N_865);
or U5716 (N_5716,N_3164,N_2100);
or U5717 (N_5717,N_1728,N_1437);
xnor U5718 (N_5718,N_3782,N_2797);
xor U5719 (N_5719,N_3784,N_1685);
or U5720 (N_5720,N_719,N_3820);
and U5721 (N_5721,N_2704,N_791);
nand U5722 (N_5722,N_1406,N_3517);
nand U5723 (N_5723,N_3932,N_653);
nor U5724 (N_5724,N_1920,N_558);
or U5725 (N_5725,N_3991,N_381);
or U5726 (N_5726,N_1565,N_2186);
and U5727 (N_5727,N_1682,N_1058);
nor U5728 (N_5728,N_1108,N_3631);
xnor U5729 (N_5729,N_3080,N_2753);
and U5730 (N_5730,N_1960,N_1019);
nand U5731 (N_5731,N_3794,N_1656);
xnor U5732 (N_5732,N_424,N_2912);
xnor U5733 (N_5733,N_1219,N_2400);
nand U5734 (N_5734,N_2542,N_1076);
nor U5735 (N_5735,N_3098,N_1919);
xor U5736 (N_5736,N_839,N_2350);
nand U5737 (N_5737,N_3933,N_2074);
or U5738 (N_5738,N_279,N_3481);
nor U5739 (N_5739,N_287,N_2373);
xor U5740 (N_5740,N_2633,N_87);
nand U5741 (N_5741,N_1601,N_1653);
xnor U5742 (N_5742,N_3935,N_854);
and U5743 (N_5743,N_3944,N_119);
nor U5744 (N_5744,N_3250,N_3402);
or U5745 (N_5745,N_400,N_2853);
xor U5746 (N_5746,N_3668,N_953);
xnor U5747 (N_5747,N_1592,N_2929);
xor U5748 (N_5748,N_410,N_954);
xor U5749 (N_5749,N_3646,N_3339);
and U5750 (N_5750,N_1547,N_2675);
nand U5751 (N_5751,N_1705,N_3506);
xor U5752 (N_5752,N_3156,N_3608);
and U5753 (N_5753,N_3824,N_1351);
nor U5754 (N_5754,N_105,N_3948);
nand U5755 (N_5755,N_2502,N_2848);
nor U5756 (N_5756,N_1961,N_957);
nand U5757 (N_5757,N_2590,N_2162);
and U5758 (N_5758,N_1144,N_3917);
xor U5759 (N_5759,N_128,N_542);
or U5760 (N_5760,N_959,N_3692);
and U5761 (N_5761,N_688,N_3099);
and U5762 (N_5762,N_1371,N_757);
and U5763 (N_5763,N_3155,N_3900);
nor U5764 (N_5764,N_2993,N_825);
nand U5765 (N_5765,N_3134,N_2872);
and U5766 (N_5766,N_1913,N_861);
or U5767 (N_5767,N_2778,N_806);
or U5768 (N_5768,N_1884,N_3599);
nand U5769 (N_5769,N_1397,N_440);
nor U5770 (N_5770,N_3999,N_1056);
or U5771 (N_5771,N_1722,N_350);
xor U5772 (N_5772,N_2913,N_1818);
nand U5773 (N_5773,N_1645,N_2708);
and U5774 (N_5774,N_1554,N_27);
and U5775 (N_5775,N_1065,N_3066);
and U5776 (N_5776,N_1483,N_2459);
xnor U5777 (N_5777,N_3819,N_2085);
or U5778 (N_5778,N_3107,N_1942);
xor U5779 (N_5779,N_159,N_327);
and U5780 (N_5780,N_2005,N_2125);
and U5781 (N_5781,N_213,N_2799);
and U5782 (N_5782,N_1771,N_1719);
and U5783 (N_5783,N_3886,N_2322);
nor U5784 (N_5784,N_3309,N_3101);
or U5785 (N_5785,N_2733,N_452);
xor U5786 (N_5786,N_3723,N_438);
and U5787 (N_5787,N_1143,N_3103);
and U5788 (N_5788,N_1321,N_3072);
and U5789 (N_5789,N_48,N_3643);
or U5790 (N_5790,N_3015,N_201);
nor U5791 (N_5791,N_354,N_3810);
nor U5792 (N_5792,N_3564,N_1387);
xor U5793 (N_5793,N_2117,N_3943);
xnor U5794 (N_5794,N_3224,N_2834);
and U5795 (N_5795,N_3859,N_902);
or U5796 (N_5796,N_823,N_3613);
or U5797 (N_5797,N_396,N_3411);
nand U5798 (N_5798,N_2965,N_2706);
nor U5799 (N_5799,N_710,N_3141);
nor U5800 (N_5800,N_3590,N_3377);
nand U5801 (N_5801,N_3060,N_1307);
and U5802 (N_5802,N_756,N_3996);
or U5803 (N_5803,N_645,N_3766);
and U5804 (N_5804,N_3460,N_2202);
nand U5805 (N_5805,N_3828,N_2463);
xnor U5806 (N_5806,N_463,N_2007);
xor U5807 (N_5807,N_830,N_1940);
xor U5808 (N_5808,N_1201,N_3190);
nand U5809 (N_5809,N_1836,N_929);
and U5810 (N_5810,N_2003,N_1059);
and U5811 (N_5811,N_3286,N_2358);
or U5812 (N_5812,N_859,N_960);
or U5813 (N_5813,N_1764,N_3112);
or U5814 (N_5814,N_1590,N_58);
nand U5815 (N_5815,N_3052,N_204);
nor U5816 (N_5816,N_1843,N_621);
nor U5817 (N_5817,N_2013,N_2238);
nand U5818 (N_5818,N_1046,N_2854);
nand U5819 (N_5819,N_3584,N_1968);
nor U5820 (N_5820,N_2800,N_479);
and U5821 (N_5821,N_3358,N_1);
nor U5822 (N_5822,N_2115,N_1766);
xnor U5823 (N_5823,N_3538,N_3673);
nor U5824 (N_5824,N_3050,N_697);
nand U5825 (N_5825,N_1822,N_2718);
nor U5826 (N_5826,N_64,N_3084);
nand U5827 (N_5827,N_1658,N_3850);
nand U5828 (N_5828,N_3233,N_3927);
and U5829 (N_5829,N_2385,N_1228);
xor U5830 (N_5830,N_3841,N_1935);
or U5831 (N_5831,N_505,N_3021);
or U5832 (N_5832,N_3879,N_2855);
nand U5833 (N_5833,N_3796,N_195);
xnor U5834 (N_5834,N_190,N_2936);
or U5835 (N_5835,N_3965,N_2147);
and U5836 (N_5836,N_2820,N_990);
nand U5837 (N_5837,N_365,N_2038);
and U5838 (N_5838,N_2218,N_1045);
xor U5839 (N_5839,N_1482,N_1150);
xnor U5840 (N_5840,N_422,N_2343);
nand U5841 (N_5841,N_3387,N_1876);
xor U5842 (N_5842,N_877,N_1037);
nor U5843 (N_5843,N_3618,N_1063);
nand U5844 (N_5844,N_2505,N_2407);
xnor U5845 (N_5845,N_3386,N_1835);
nor U5846 (N_5846,N_949,N_1363);
nand U5847 (N_5847,N_3899,N_229);
or U5848 (N_5848,N_443,N_745);
and U5849 (N_5849,N_1677,N_3984);
and U5850 (N_5850,N_2715,N_2762);
or U5851 (N_5851,N_1295,N_2105);
nand U5852 (N_5852,N_1376,N_98);
or U5853 (N_5853,N_1567,N_3420);
and U5854 (N_5854,N_2616,N_2178);
or U5855 (N_5855,N_2209,N_1293);
nor U5856 (N_5856,N_2369,N_2630);
nor U5857 (N_5857,N_3177,N_2506);
or U5858 (N_5858,N_2651,N_2642);
nand U5859 (N_5859,N_1090,N_3117);
and U5860 (N_5860,N_255,N_355);
nand U5861 (N_5861,N_2287,N_3047);
xnor U5862 (N_5862,N_3147,N_1052);
xor U5863 (N_5863,N_3816,N_3237);
and U5864 (N_5864,N_2939,N_672);
xor U5865 (N_5865,N_3789,N_1621);
or U5866 (N_5866,N_1977,N_3817);
and U5867 (N_5867,N_945,N_886);
nor U5868 (N_5868,N_655,N_1641);
xor U5869 (N_5869,N_2245,N_2259);
xnor U5870 (N_5870,N_3096,N_1855);
nand U5871 (N_5871,N_1579,N_1881);
xor U5872 (N_5872,N_3269,N_1755);
and U5873 (N_5873,N_3397,N_3078);
or U5874 (N_5874,N_846,N_927);
and U5875 (N_5875,N_591,N_2976);
xor U5876 (N_5876,N_921,N_607);
or U5877 (N_5877,N_1198,N_1506);
and U5878 (N_5878,N_3902,N_1323);
nor U5879 (N_5879,N_2042,N_1454);
nand U5880 (N_5880,N_3583,N_1832);
and U5881 (N_5881,N_907,N_2133);
nand U5882 (N_5882,N_2713,N_3105);
and U5883 (N_5883,N_1538,N_2741);
and U5884 (N_5884,N_1074,N_1053);
xor U5885 (N_5885,N_2419,N_1067);
nand U5886 (N_5886,N_398,N_1003);
nand U5887 (N_5887,N_2262,N_1098);
xnor U5888 (N_5888,N_1455,N_136);
nor U5889 (N_5889,N_2366,N_1269);
or U5890 (N_5890,N_137,N_969);
nor U5891 (N_5891,N_1158,N_402);
nor U5892 (N_5892,N_819,N_1211);
nand U5893 (N_5893,N_1436,N_687);
nor U5894 (N_5894,N_1680,N_3218);
nand U5895 (N_5895,N_18,N_1874);
xor U5896 (N_5896,N_1742,N_2923);
nand U5897 (N_5897,N_3022,N_781);
or U5898 (N_5898,N_300,N_2054);
nor U5899 (N_5899,N_3990,N_887);
and U5900 (N_5900,N_3809,N_328);
nand U5901 (N_5901,N_485,N_1285);
and U5902 (N_5902,N_2411,N_3217);
nor U5903 (N_5903,N_1924,N_2093);
xor U5904 (N_5904,N_1097,N_1905);
xnor U5905 (N_5905,N_818,N_1450);
nand U5906 (N_5906,N_3959,N_2025);
or U5907 (N_5907,N_397,N_3495);
xor U5908 (N_5908,N_259,N_1606);
nor U5909 (N_5909,N_3891,N_3272);
and U5910 (N_5910,N_3102,N_2249);
xor U5911 (N_5911,N_377,N_3671);
nor U5912 (N_5912,N_931,N_310);
nor U5913 (N_5913,N_3617,N_3501);
or U5914 (N_5914,N_3391,N_1566);
nand U5915 (N_5915,N_3205,N_401);
and U5916 (N_5916,N_928,N_84);
and U5917 (N_5917,N_1993,N_1148);
or U5918 (N_5918,N_1071,N_3185);
and U5919 (N_5919,N_1923,N_1259);
nor U5920 (N_5920,N_2268,N_3158);
xor U5921 (N_5921,N_2792,N_3682);
nor U5922 (N_5922,N_2991,N_1548);
xnor U5923 (N_5923,N_1306,N_2119);
nand U5924 (N_5924,N_1871,N_3858);
nand U5925 (N_5925,N_1388,N_3716);
and U5926 (N_5926,N_3825,N_2771);
nand U5927 (N_5927,N_2211,N_581);
nand U5928 (N_5928,N_3903,N_890);
and U5929 (N_5929,N_837,N_987);
nand U5930 (N_5930,N_1949,N_2824);
nor U5931 (N_5931,N_1675,N_3211);
xor U5932 (N_5932,N_2806,N_2917);
xnor U5933 (N_5933,N_2457,N_2497);
or U5934 (N_5934,N_2275,N_26);
nand U5935 (N_5935,N_3528,N_1103);
or U5936 (N_5936,N_2453,N_662);
nand U5937 (N_5937,N_2444,N_147);
xor U5938 (N_5938,N_1845,N_3737);
and U5939 (N_5939,N_608,N_3461);
and U5940 (N_5940,N_3513,N_335);
nor U5941 (N_5941,N_509,N_1013);
or U5942 (N_5942,N_1021,N_2197);
or U5943 (N_5943,N_797,N_3529);
and U5944 (N_5944,N_2591,N_1805);
xnor U5945 (N_5945,N_2480,N_2272);
xor U5946 (N_5946,N_592,N_2312);
or U5947 (N_5947,N_2204,N_3889);
nand U5948 (N_5948,N_2525,N_17);
and U5949 (N_5949,N_264,N_1659);
nor U5950 (N_5950,N_1124,N_3184);
nand U5951 (N_5951,N_2663,N_152);
nand U5952 (N_5952,N_3235,N_1448);
nand U5953 (N_5953,N_2144,N_2906);
nor U5954 (N_5954,N_3470,N_2055);
or U5955 (N_5955,N_3721,N_2723);
and U5956 (N_5956,N_2810,N_2766);
and U5957 (N_5957,N_2790,N_345);
nor U5958 (N_5958,N_3380,N_2709);
nor U5959 (N_5959,N_3504,N_1999);
nand U5960 (N_5960,N_1230,N_1233);
nor U5961 (N_5961,N_3088,N_2635);
nand U5962 (N_5962,N_516,N_3385);
nand U5963 (N_5963,N_2288,N_242);
nand U5964 (N_5964,N_1478,N_895);
xor U5965 (N_5965,N_3485,N_1023);
nor U5966 (N_5966,N_2515,N_2958);
xnor U5967 (N_5967,N_319,N_1558);
nor U5968 (N_5968,N_3284,N_496);
xnor U5969 (N_5969,N_2765,N_47);
nand U5970 (N_5970,N_2476,N_2090);
or U5971 (N_5971,N_149,N_2428);
nand U5972 (N_5972,N_179,N_1210);
or U5973 (N_5973,N_474,N_2897);
or U5974 (N_5974,N_244,N_2122);
or U5975 (N_5975,N_3035,N_412);
and U5976 (N_5976,N_1330,N_2353);
nor U5977 (N_5977,N_2572,N_3290);
and U5978 (N_5978,N_550,N_3777);
and U5979 (N_5979,N_133,N_3153);
nor U5980 (N_5980,N_1249,N_3081);
or U5981 (N_5981,N_2412,N_3815);
nand U5982 (N_5982,N_2283,N_3361);
nand U5983 (N_5983,N_3747,N_596);
or U5984 (N_5984,N_2132,N_3455);
and U5985 (N_5985,N_1570,N_2756);
nor U5986 (N_5986,N_1500,N_627);
nand U5987 (N_5987,N_2873,N_3856);
or U5988 (N_5988,N_1954,N_633);
xor U5989 (N_5989,N_226,N_2996);
or U5990 (N_5990,N_2227,N_9);
and U5991 (N_5991,N_394,N_2636);
or U5992 (N_5992,N_1442,N_1612);
nor U5993 (N_5993,N_3546,N_998);
nor U5994 (N_5994,N_810,N_1191);
nor U5995 (N_5995,N_421,N_2325);
or U5996 (N_5996,N_2731,N_2423);
xor U5997 (N_5997,N_2278,N_874);
and U5998 (N_5998,N_3689,N_2816);
nand U5999 (N_5999,N_1001,N_693);
xnor U6000 (N_6000,N_1691,N_1844);
nand U6001 (N_6001,N_672,N_619);
and U6002 (N_6002,N_1643,N_135);
xor U6003 (N_6003,N_807,N_2327);
and U6004 (N_6004,N_2081,N_929);
and U6005 (N_6005,N_3892,N_874);
nor U6006 (N_6006,N_2406,N_2768);
xnor U6007 (N_6007,N_3842,N_3211);
and U6008 (N_6008,N_1486,N_261);
nor U6009 (N_6009,N_492,N_268);
or U6010 (N_6010,N_824,N_2021);
nor U6011 (N_6011,N_172,N_2089);
nor U6012 (N_6012,N_1595,N_536);
or U6013 (N_6013,N_2019,N_428);
xor U6014 (N_6014,N_1805,N_3353);
nor U6015 (N_6015,N_3007,N_3607);
xor U6016 (N_6016,N_3634,N_309);
nand U6017 (N_6017,N_2529,N_451);
nand U6018 (N_6018,N_2661,N_1768);
nand U6019 (N_6019,N_1472,N_905);
and U6020 (N_6020,N_976,N_1471);
and U6021 (N_6021,N_3457,N_2459);
xor U6022 (N_6022,N_3517,N_1436);
or U6023 (N_6023,N_2057,N_3907);
nand U6024 (N_6024,N_688,N_1180);
and U6025 (N_6025,N_1936,N_1199);
nand U6026 (N_6026,N_699,N_3997);
nor U6027 (N_6027,N_2939,N_3341);
xor U6028 (N_6028,N_2812,N_3556);
nand U6029 (N_6029,N_3899,N_2461);
and U6030 (N_6030,N_2424,N_3898);
or U6031 (N_6031,N_1598,N_2220);
nand U6032 (N_6032,N_326,N_2103);
nor U6033 (N_6033,N_2331,N_2458);
xnor U6034 (N_6034,N_2607,N_1051);
and U6035 (N_6035,N_3318,N_276);
xnor U6036 (N_6036,N_1580,N_3888);
nand U6037 (N_6037,N_3742,N_3675);
nor U6038 (N_6038,N_3533,N_2898);
nor U6039 (N_6039,N_74,N_967);
nand U6040 (N_6040,N_242,N_1049);
and U6041 (N_6041,N_2109,N_2190);
xnor U6042 (N_6042,N_1334,N_2724);
or U6043 (N_6043,N_3124,N_3119);
and U6044 (N_6044,N_3959,N_3582);
xnor U6045 (N_6045,N_1537,N_301);
nor U6046 (N_6046,N_1674,N_1703);
nand U6047 (N_6047,N_2267,N_100);
or U6048 (N_6048,N_3101,N_2949);
nand U6049 (N_6049,N_1531,N_660);
nand U6050 (N_6050,N_1866,N_3657);
xor U6051 (N_6051,N_1160,N_3891);
nand U6052 (N_6052,N_2980,N_682);
xor U6053 (N_6053,N_1522,N_2634);
or U6054 (N_6054,N_2868,N_3375);
nand U6055 (N_6055,N_1601,N_2329);
nor U6056 (N_6056,N_790,N_3650);
xnor U6057 (N_6057,N_3819,N_2404);
xor U6058 (N_6058,N_2144,N_3291);
nor U6059 (N_6059,N_3767,N_1137);
nand U6060 (N_6060,N_3524,N_1472);
or U6061 (N_6061,N_2426,N_2070);
nand U6062 (N_6062,N_229,N_1154);
nor U6063 (N_6063,N_303,N_3849);
nor U6064 (N_6064,N_1301,N_1727);
and U6065 (N_6065,N_1155,N_1183);
nand U6066 (N_6066,N_3548,N_3505);
nor U6067 (N_6067,N_3027,N_3841);
nor U6068 (N_6068,N_2891,N_435);
or U6069 (N_6069,N_2546,N_3962);
nor U6070 (N_6070,N_664,N_951);
or U6071 (N_6071,N_2024,N_3030);
or U6072 (N_6072,N_643,N_2173);
or U6073 (N_6073,N_1231,N_2953);
xnor U6074 (N_6074,N_1589,N_1931);
xnor U6075 (N_6075,N_1241,N_2445);
nand U6076 (N_6076,N_206,N_573);
and U6077 (N_6077,N_2419,N_1911);
nor U6078 (N_6078,N_2558,N_1742);
nand U6079 (N_6079,N_1935,N_3731);
nand U6080 (N_6080,N_3319,N_1733);
xnor U6081 (N_6081,N_2379,N_19);
and U6082 (N_6082,N_1032,N_587);
nand U6083 (N_6083,N_3795,N_2764);
nor U6084 (N_6084,N_1173,N_792);
xnor U6085 (N_6085,N_121,N_286);
nor U6086 (N_6086,N_592,N_2859);
nor U6087 (N_6087,N_2534,N_1189);
nor U6088 (N_6088,N_3523,N_908);
nand U6089 (N_6089,N_1815,N_3814);
or U6090 (N_6090,N_1193,N_1004);
and U6091 (N_6091,N_3659,N_3542);
nand U6092 (N_6092,N_3831,N_3631);
nand U6093 (N_6093,N_2516,N_2754);
xnor U6094 (N_6094,N_2391,N_3646);
xor U6095 (N_6095,N_697,N_3804);
nand U6096 (N_6096,N_91,N_3946);
nand U6097 (N_6097,N_2302,N_2487);
and U6098 (N_6098,N_1025,N_2850);
nand U6099 (N_6099,N_3097,N_3911);
nor U6100 (N_6100,N_2132,N_711);
xor U6101 (N_6101,N_1037,N_3104);
nor U6102 (N_6102,N_3290,N_2467);
and U6103 (N_6103,N_2259,N_3898);
or U6104 (N_6104,N_455,N_88);
nand U6105 (N_6105,N_3918,N_1486);
xnor U6106 (N_6106,N_1853,N_3582);
or U6107 (N_6107,N_2150,N_1294);
and U6108 (N_6108,N_1776,N_272);
xnor U6109 (N_6109,N_2956,N_3667);
or U6110 (N_6110,N_3995,N_3502);
or U6111 (N_6111,N_1515,N_3424);
nor U6112 (N_6112,N_3096,N_3039);
or U6113 (N_6113,N_2741,N_2461);
and U6114 (N_6114,N_3454,N_885);
nand U6115 (N_6115,N_1317,N_1023);
and U6116 (N_6116,N_3742,N_1218);
nor U6117 (N_6117,N_129,N_2363);
nand U6118 (N_6118,N_3150,N_2396);
nand U6119 (N_6119,N_2144,N_3067);
xnor U6120 (N_6120,N_1610,N_1871);
nand U6121 (N_6121,N_283,N_612);
or U6122 (N_6122,N_1782,N_3112);
or U6123 (N_6123,N_302,N_1554);
xor U6124 (N_6124,N_3784,N_3878);
and U6125 (N_6125,N_891,N_500);
or U6126 (N_6126,N_183,N_1044);
nor U6127 (N_6127,N_2678,N_689);
and U6128 (N_6128,N_2030,N_754);
or U6129 (N_6129,N_1534,N_539);
nor U6130 (N_6130,N_3308,N_1624);
xnor U6131 (N_6131,N_688,N_2452);
xnor U6132 (N_6132,N_374,N_3327);
nand U6133 (N_6133,N_2869,N_250);
or U6134 (N_6134,N_3692,N_3906);
and U6135 (N_6135,N_1539,N_1434);
nand U6136 (N_6136,N_476,N_1980);
or U6137 (N_6137,N_3984,N_3040);
nand U6138 (N_6138,N_2522,N_3803);
and U6139 (N_6139,N_1264,N_3826);
and U6140 (N_6140,N_1649,N_1540);
or U6141 (N_6141,N_1592,N_2685);
nand U6142 (N_6142,N_1977,N_1605);
nand U6143 (N_6143,N_1232,N_1416);
nor U6144 (N_6144,N_560,N_2760);
and U6145 (N_6145,N_2146,N_640);
xnor U6146 (N_6146,N_2409,N_480);
and U6147 (N_6147,N_2088,N_589);
and U6148 (N_6148,N_3845,N_1231);
xnor U6149 (N_6149,N_493,N_3614);
nor U6150 (N_6150,N_511,N_1032);
xnor U6151 (N_6151,N_912,N_2009);
nand U6152 (N_6152,N_612,N_823);
and U6153 (N_6153,N_2895,N_2452);
and U6154 (N_6154,N_1113,N_2019);
nand U6155 (N_6155,N_1845,N_3093);
nor U6156 (N_6156,N_621,N_3230);
nand U6157 (N_6157,N_559,N_1738);
nand U6158 (N_6158,N_3382,N_3379);
or U6159 (N_6159,N_3033,N_1346);
and U6160 (N_6160,N_1670,N_847);
nand U6161 (N_6161,N_1161,N_3937);
and U6162 (N_6162,N_2776,N_661);
xnor U6163 (N_6163,N_3599,N_3086);
and U6164 (N_6164,N_1383,N_2845);
nand U6165 (N_6165,N_1635,N_186);
xor U6166 (N_6166,N_2242,N_3962);
or U6167 (N_6167,N_2487,N_1779);
nand U6168 (N_6168,N_3304,N_3429);
and U6169 (N_6169,N_868,N_53);
or U6170 (N_6170,N_1256,N_2614);
xor U6171 (N_6171,N_3389,N_328);
xor U6172 (N_6172,N_1430,N_653);
or U6173 (N_6173,N_1770,N_3858);
or U6174 (N_6174,N_2654,N_2933);
xnor U6175 (N_6175,N_1031,N_3406);
or U6176 (N_6176,N_1465,N_3177);
nor U6177 (N_6177,N_3579,N_425);
nor U6178 (N_6178,N_3882,N_3104);
nor U6179 (N_6179,N_2309,N_3960);
nand U6180 (N_6180,N_88,N_3457);
and U6181 (N_6181,N_3208,N_152);
or U6182 (N_6182,N_2391,N_3968);
xnor U6183 (N_6183,N_965,N_1549);
nor U6184 (N_6184,N_1944,N_3808);
xor U6185 (N_6185,N_2710,N_2289);
or U6186 (N_6186,N_3149,N_3235);
nor U6187 (N_6187,N_91,N_523);
nor U6188 (N_6188,N_1661,N_958);
nand U6189 (N_6189,N_1810,N_894);
xor U6190 (N_6190,N_229,N_3179);
nor U6191 (N_6191,N_2638,N_663);
nor U6192 (N_6192,N_339,N_2102);
nand U6193 (N_6193,N_1561,N_2756);
and U6194 (N_6194,N_2500,N_2320);
or U6195 (N_6195,N_2378,N_3035);
xnor U6196 (N_6196,N_3191,N_1644);
xor U6197 (N_6197,N_1396,N_3087);
xnor U6198 (N_6198,N_2478,N_3168);
or U6199 (N_6199,N_1924,N_2503);
nand U6200 (N_6200,N_3682,N_2037);
or U6201 (N_6201,N_1767,N_861);
and U6202 (N_6202,N_3226,N_3230);
xor U6203 (N_6203,N_230,N_1527);
nand U6204 (N_6204,N_1927,N_12);
or U6205 (N_6205,N_81,N_2167);
and U6206 (N_6206,N_2048,N_2737);
xor U6207 (N_6207,N_2870,N_937);
nand U6208 (N_6208,N_1466,N_2736);
or U6209 (N_6209,N_1405,N_3332);
xnor U6210 (N_6210,N_2369,N_1529);
nand U6211 (N_6211,N_3289,N_1942);
nor U6212 (N_6212,N_2983,N_3274);
and U6213 (N_6213,N_1824,N_1746);
nor U6214 (N_6214,N_1812,N_688);
or U6215 (N_6215,N_518,N_347);
and U6216 (N_6216,N_381,N_2439);
xnor U6217 (N_6217,N_331,N_839);
xnor U6218 (N_6218,N_562,N_2374);
and U6219 (N_6219,N_1003,N_805);
or U6220 (N_6220,N_280,N_3702);
xnor U6221 (N_6221,N_3905,N_230);
nor U6222 (N_6222,N_1055,N_611);
nor U6223 (N_6223,N_3673,N_656);
and U6224 (N_6224,N_528,N_1951);
and U6225 (N_6225,N_2248,N_2651);
xnor U6226 (N_6226,N_3410,N_2194);
xnor U6227 (N_6227,N_2060,N_3991);
and U6228 (N_6228,N_3647,N_1464);
or U6229 (N_6229,N_1874,N_2119);
or U6230 (N_6230,N_479,N_1089);
nor U6231 (N_6231,N_3128,N_495);
nand U6232 (N_6232,N_3019,N_2501);
and U6233 (N_6233,N_1105,N_2332);
xnor U6234 (N_6234,N_3186,N_2954);
nand U6235 (N_6235,N_2111,N_2420);
and U6236 (N_6236,N_282,N_2409);
nand U6237 (N_6237,N_3620,N_2664);
or U6238 (N_6238,N_2126,N_3246);
xnor U6239 (N_6239,N_1183,N_800);
nand U6240 (N_6240,N_3179,N_3037);
xnor U6241 (N_6241,N_2260,N_3946);
xnor U6242 (N_6242,N_2872,N_1718);
or U6243 (N_6243,N_3834,N_2722);
nand U6244 (N_6244,N_610,N_76);
nand U6245 (N_6245,N_317,N_2223);
nor U6246 (N_6246,N_2570,N_378);
nand U6247 (N_6247,N_931,N_1879);
nand U6248 (N_6248,N_2498,N_3683);
nand U6249 (N_6249,N_173,N_2443);
nand U6250 (N_6250,N_654,N_1600);
or U6251 (N_6251,N_2212,N_3737);
xor U6252 (N_6252,N_811,N_2014);
xnor U6253 (N_6253,N_322,N_3987);
and U6254 (N_6254,N_2744,N_1753);
nor U6255 (N_6255,N_541,N_3650);
nand U6256 (N_6256,N_3854,N_2994);
or U6257 (N_6257,N_789,N_146);
or U6258 (N_6258,N_3901,N_1233);
and U6259 (N_6259,N_1783,N_3984);
nand U6260 (N_6260,N_3667,N_3604);
xnor U6261 (N_6261,N_3493,N_2456);
or U6262 (N_6262,N_3894,N_3812);
and U6263 (N_6263,N_1001,N_3685);
nand U6264 (N_6264,N_3385,N_3038);
nor U6265 (N_6265,N_3538,N_3900);
nand U6266 (N_6266,N_807,N_1950);
or U6267 (N_6267,N_2085,N_2800);
and U6268 (N_6268,N_1220,N_3132);
nor U6269 (N_6269,N_712,N_3507);
xor U6270 (N_6270,N_2817,N_3525);
and U6271 (N_6271,N_3419,N_2558);
xnor U6272 (N_6272,N_2626,N_2193);
nand U6273 (N_6273,N_1889,N_809);
xnor U6274 (N_6274,N_3582,N_829);
nand U6275 (N_6275,N_1035,N_2011);
xor U6276 (N_6276,N_3959,N_1614);
and U6277 (N_6277,N_2091,N_449);
xnor U6278 (N_6278,N_1964,N_2342);
and U6279 (N_6279,N_2083,N_3782);
nand U6280 (N_6280,N_3993,N_2611);
xor U6281 (N_6281,N_1003,N_1084);
xor U6282 (N_6282,N_2957,N_942);
nor U6283 (N_6283,N_3086,N_2438);
xnor U6284 (N_6284,N_282,N_1385);
and U6285 (N_6285,N_3527,N_2177);
and U6286 (N_6286,N_384,N_2273);
and U6287 (N_6287,N_2683,N_2120);
nor U6288 (N_6288,N_2847,N_3755);
and U6289 (N_6289,N_286,N_756);
xor U6290 (N_6290,N_71,N_2592);
xor U6291 (N_6291,N_1088,N_3490);
or U6292 (N_6292,N_170,N_3435);
nand U6293 (N_6293,N_614,N_2183);
or U6294 (N_6294,N_2737,N_3494);
nand U6295 (N_6295,N_1334,N_2560);
nand U6296 (N_6296,N_588,N_3310);
and U6297 (N_6297,N_2197,N_2749);
xnor U6298 (N_6298,N_2352,N_649);
nand U6299 (N_6299,N_1565,N_3277);
nand U6300 (N_6300,N_1187,N_1787);
or U6301 (N_6301,N_1583,N_346);
xnor U6302 (N_6302,N_2170,N_3015);
nand U6303 (N_6303,N_735,N_2702);
nor U6304 (N_6304,N_656,N_230);
nand U6305 (N_6305,N_3488,N_2665);
xor U6306 (N_6306,N_395,N_655);
nand U6307 (N_6307,N_2509,N_592);
nand U6308 (N_6308,N_3359,N_3548);
xnor U6309 (N_6309,N_536,N_3398);
nor U6310 (N_6310,N_1051,N_3804);
nor U6311 (N_6311,N_2215,N_1526);
and U6312 (N_6312,N_3088,N_3438);
nand U6313 (N_6313,N_234,N_1702);
xnor U6314 (N_6314,N_2427,N_2281);
xnor U6315 (N_6315,N_3484,N_3680);
and U6316 (N_6316,N_1737,N_2364);
or U6317 (N_6317,N_3598,N_8);
and U6318 (N_6318,N_1119,N_20);
or U6319 (N_6319,N_2247,N_966);
xor U6320 (N_6320,N_2502,N_2676);
or U6321 (N_6321,N_3688,N_138);
xnor U6322 (N_6322,N_3281,N_2413);
or U6323 (N_6323,N_523,N_825);
or U6324 (N_6324,N_3303,N_2803);
nor U6325 (N_6325,N_472,N_1469);
nand U6326 (N_6326,N_1404,N_1752);
or U6327 (N_6327,N_49,N_2450);
nand U6328 (N_6328,N_2758,N_1192);
or U6329 (N_6329,N_2768,N_1524);
nand U6330 (N_6330,N_2304,N_3275);
nor U6331 (N_6331,N_3976,N_2448);
and U6332 (N_6332,N_2185,N_585);
nor U6333 (N_6333,N_3804,N_2822);
xnor U6334 (N_6334,N_38,N_3091);
nand U6335 (N_6335,N_311,N_3682);
nor U6336 (N_6336,N_2819,N_2466);
xor U6337 (N_6337,N_3885,N_83);
or U6338 (N_6338,N_13,N_2041);
nand U6339 (N_6339,N_2087,N_1706);
nand U6340 (N_6340,N_1516,N_2569);
and U6341 (N_6341,N_2313,N_744);
nand U6342 (N_6342,N_3339,N_750);
or U6343 (N_6343,N_3793,N_512);
nand U6344 (N_6344,N_1146,N_2376);
and U6345 (N_6345,N_1123,N_616);
nand U6346 (N_6346,N_2768,N_3340);
xor U6347 (N_6347,N_2855,N_1841);
xor U6348 (N_6348,N_1493,N_1019);
xnor U6349 (N_6349,N_1698,N_1795);
or U6350 (N_6350,N_1906,N_3943);
or U6351 (N_6351,N_922,N_1442);
or U6352 (N_6352,N_674,N_2530);
nor U6353 (N_6353,N_3026,N_2145);
nor U6354 (N_6354,N_2825,N_899);
nand U6355 (N_6355,N_1580,N_1640);
xnor U6356 (N_6356,N_3078,N_1509);
and U6357 (N_6357,N_2791,N_851);
xnor U6358 (N_6358,N_3079,N_2278);
or U6359 (N_6359,N_3745,N_333);
or U6360 (N_6360,N_1993,N_3251);
nor U6361 (N_6361,N_2537,N_100);
nand U6362 (N_6362,N_686,N_1411);
nand U6363 (N_6363,N_339,N_682);
and U6364 (N_6364,N_402,N_3557);
nand U6365 (N_6365,N_1177,N_2671);
and U6366 (N_6366,N_202,N_2498);
and U6367 (N_6367,N_1510,N_2497);
and U6368 (N_6368,N_3507,N_397);
xnor U6369 (N_6369,N_2794,N_123);
or U6370 (N_6370,N_1599,N_146);
or U6371 (N_6371,N_721,N_1587);
nand U6372 (N_6372,N_1790,N_623);
xor U6373 (N_6373,N_285,N_3710);
xnor U6374 (N_6374,N_243,N_257);
nor U6375 (N_6375,N_1359,N_3642);
nand U6376 (N_6376,N_2474,N_3705);
nand U6377 (N_6377,N_3420,N_772);
and U6378 (N_6378,N_2884,N_2627);
xnor U6379 (N_6379,N_3769,N_2370);
nand U6380 (N_6380,N_71,N_3395);
nor U6381 (N_6381,N_250,N_2085);
or U6382 (N_6382,N_174,N_3508);
xor U6383 (N_6383,N_3327,N_283);
or U6384 (N_6384,N_1397,N_2857);
and U6385 (N_6385,N_1024,N_1087);
nor U6386 (N_6386,N_2855,N_3023);
nor U6387 (N_6387,N_99,N_1828);
or U6388 (N_6388,N_1982,N_3211);
and U6389 (N_6389,N_3475,N_3964);
nand U6390 (N_6390,N_433,N_1196);
nor U6391 (N_6391,N_1433,N_1702);
or U6392 (N_6392,N_3077,N_1044);
nor U6393 (N_6393,N_837,N_716);
and U6394 (N_6394,N_1904,N_645);
and U6395 (N_6395,N_1029,N_730);
xor U6396 (N_6396,N_1532,N_146);
or U6397 (N_6397,N_195,N_2415);
and U6398 (N_6398,N_360,N_3566);
and U6399 (N_6399,N_3800,N_229);
nand U6400 (N_6400,N_1029,N_1486);
nor U6401 (N_6401,N_1885,N_1839);
or U6402 (N_6402,N_2993,N_2413);
and U6403 (N_6403,N_1290,N_866);
nor U6404 (N_6404,N_1782,N_1209);
nand U6405 (N_6405,N_1609,N_150);
or U6406 (N_6406,N_2221,N_2222);
xor U6407 (N_6407,N_2655,N_2547);
nor U6408 (N_6408,N_564,N_3813);
nor U6409 (N_6409,N_3930,N_1256);
xnor U6410 (N_6410,N_2041,N_2129);
xor U6411 (N_6411,N_3766,N_2934);
nor U6412 (N_6412,N_2694,N_3243);
and U6413 (N_6413,N_549,N_2584);
nand U6414 (N_6414,N_849,N_647);
or U6415 (N_6415,N_588,N_2142);
and U6416 (N_6416,N_599,N_248);
or U6417 (N_6417,N_3553,N_2718);
xnor U6418 (N_6418,N_3482,N_3435);
nor U6419 (N_6419,N_3407,N_2735);
or U6420 (N_6420,N_2694,N_1607);
nor U6421 (N_6421,N_30,N_3699);
xor U6422 (N_6422,N_472,N_596);
xnor U6423 (N_6423,N_1708,N_1566);
nand U6424 (N_6424,N_3842,N_3358);
xnor U6425 (N_6425,N_881,N_3785);
nand U6426 (N_6426,N_152,N_2708);
and U6427 (N_6427,N_222,N_2102);
or U6428 (N_6428,N_3588,N_2871);
xnor U6429 (N_6429,N_2089,N_2387);
and U6430 (N_6430,N_2801,N_1757);
xor U6431 (N_6431,N_979,N_1335);
nand U6432 (N_6432,N_3933,N_1015);
nor U6433 (N_6433,N_2418,N_1633);
nor U6434 (N_6434,N_3744,N_2895);
nor U6435 (N_6435,N_3492,N_2458);
or U6436 (N_6436,N_1774,N_100);
nor U6437 (N_6437,N_2771,N_3432);
nand U6438 (N_6438,N_2433,N_3686);
xor U6439 (N_6439,N_935,N_2999);
nand U6440 (N_6440,N_2451,N_75);
nor U6441 (N_6441,N_2672,N_929);
and U6442 (N_6442,N_1271,N_3206);
xor U6443 (N_6443,N_1885,N_530);
nand U6444 (N_6444,N_1213,N_3587);
xnor U6445 (N_6445,N_3463,N_1096);
or U6446 (N_6446,N_299,N_2758);
nand U6447 (N_6447,N_2678,N_473);
or U6448 (N_6448,N_1474,N_1736);
xnor U6449 (N_6449,N_2449,N_348);
nand U6450 (N_6450,N_3042,N_2744);
and U6451 (N_6451,N_363,N_721);
or U6452 (N_6452,N_3513,N_3675);
or U6453 (N_6453,N_3585,N_58);
nand U6454 (N_6454,N_2737,N_3135);
and U6455 (N_6455,N_2973,N_1303);
nor U6456 (N_6456,N_513,N_1592);
nor U6457 (N_6457,N_524,N_3055);
nand U6458 (N_6458,N_3954,N_3603);
or U6459 (N_6459,N_171,N_3017);
nor U6460 (N_6460,N_702,N_859);
nor U6461 (N_6461,N_1881,N_380);
xor U6462 (N_6462,N_3334,N_1188);
nand U6463 (N_6463,N_673,N_1160);
nor U6464 (N_6464,N_1456,N_3676);
or U6465 (N_6465,N_3804,N_288);
xnor U6466 (N_6466,N_2405,N_2124);
nand U6467 (N_6467,N_737,N_568);
and U6468 (N_6468,N_422,N_3831);
nor U6469 (N_6469,N_2538,N_1565);
xnor U6470 (N_6470,N_1333,N_2252);
nand U6471 (N_6471,N_3658,N_3641);
xnor U6472 (N_6472,N_1267,N_1938);
xor U6473 (N_6473,N_1289,N_2067);
xnor U6474 (N_6474,N_1202,N_1632);
nor U6475 (N_6475,N_2640,N_1404);
or U6476 (N_6476,N_1478,N_1764);
or U6477 (N_6477,N_247,N_2524);
nand U6478 (N_6478,N_1438,N_2167);
nor U6479 (N_6479,N_2204,N_3454);
nand U6480 (N_6480,N_3992,N_1198);
and U6481 (N_6481,N_1838,N_2527);
nand U6482 (N_6482,N_578,N_1591);
nand U6483 (N_6483,N_35,N_1905);
xor U6484 (N_6484,N_2297,N_767);
and U6485 (N_6485,N_1452,N_899);
and U6486 (N_6486,N_213,N_2782);
nand U6487 (N_6487,N_3823,N_2082);
nor U6488 (N_6488,N_3777,N_905);
nand U6489 (N_6489,N_2530,N_898);
and U6490 (N_6490,N_52,N_2265);
xnor U6491 (N_6491,N_260,N_3243);
xor U6492 (N_6492,N_2926,N_1863);
nor U6493 (N_6493,N_280,N_1155);
or U6494 (N_6494,N_277,N_2060);
nand U6495 (N_6495,N_3447,N_3671);
nor U6496 (N_6496,N_89,N_3987);
and U6497 (N_6497,N_754,N_1413);
xnor U6498 (N_6498,N_2351,N_3852);
and U6499 (N_6499,N_3650,N_3713);
nand U6500 (N_6500,N_2842,N_279);
xnor U6501 (N_6501,N_2379,N_1088);
nor U6502 (N_6502,N_1331,N_2885);
and U6503 (N_6503,N_3032,N_1754);
nand U6504 (N_6504,N_1498,N_2014);
or U6505 (N_6505,N_492,N_3859);
nand U6506 (N_6506,N_2140,N_3406);
nand U6507 (N_6507,N_3245,N_3494);
xnor U6508 (N_6508,N_3112,N_1110);
or U6509 (N_6509,N_864,N_3125);
xor U6510 (N_6510,N_2427,N_3808);
xor U6511 (N_6511,N_3817,N_1823);
and U6512 (N_6512,N_3406,N_3033);
or U6513 (N_6513,N_2691,N_826);
or U6514 (N_6514,N_697,N_2704);
or U6515 (N_6515,N_2031,N_1339);
nand U6516 (N_6516,N_1115,N_2331);
nor U6517 (N_6517,N_1261,N_2563);
xnor U6518 (N_6518,N_4,N_1992);
or U6519 (N_6519,N_1350,N_2194);
and U6520 (N_6520,N_3052,N_3478);
nand U6521 (N_6521,N_2842,N_584);
and U6522 (N_6522,N_2986,N_2246);
xor U6523 (N_6523,N_1625,N_2670);
nor U6524 (N_6524,N_3848,N_3434);
nor U6525 (N_6525,N_775,N_1686);
nor U6526 (N_6526,N_2351,N_760);
and U6527 (N_6527,N_3651,N_1256);
nor U6528 (N_6528,N_2451,N_3432);
nand U6529 (N_6529,N_3454,N_3723);
nor U6530 (N_6530,N_1062,N_2373);
nor U6531 (N_6531,N_363,N_3761);
nand U6532 (N_6532,N_3178,N_652);
nor U6533 (N_6533,N_188,N_915);
xor U6534 (N_6534,N_3855,N_1415);
or U6535 (N_6535,N_2128,N_448);
and U6536 (N_6536,N_3461,N_667);
or U6537 (N_6537,N_2408,N_300);
or U6538 (N_6538,N_909,N_1674);
or U6539 (N_6539,N_2579,N_1995);
xor U6540 (N_6540,N_415,N_3748);
nand U6541 (N_6541,N_3172,N_2326);
or U6542 (N_6542,N_619,N_60);
nor U6543 (N_6543,N_1772,N_1697);
xnor U6544 (N_6544,N_2363,N_2689);
and U6545 (N_6545,N_535,N_173);
xnor U6546 (N_6546,N_1299,N_3513);
and U6547 (N_6547,N_2625,N_2786);
or U6548 (N_6548,N_1865,N_196);
and U6549 (N_6549,N_3215,N_2383);
xnor U6550 (N_6550,N_2290,N_3123);
nor U6551 (N_6551,N_2843,N_3435);
xor U6552 (N_6552,N_2125,N_2940);
and U6553 (N_6553,N_3852,N_2648);
or U6554 (N_6554,N_543,N_871);
xor U6555 (N_6555,N_542,N_3529);
and U6556 (N_6556,N_1336,N_3840);
nand U6557 (N_6557,N_1957,N_805);
and U6558 (N_6558,N_573,N_3045);
nand U6559 (N_6559,N_1331,N_3190);
and U6560 (N_6560,N_1870,N_1386);
nand U6561 (N_6561,N_49,N_2140);
or U6562 (N_6562,N_1861,N_826);
and U6563 (N_6563,N_3030,N_2643);
xnor U6564 (N_6564,N_1357,N_2797);
nor U6565 (N_6565,N_1250,N_3572);
nand U6566 (N_6566,N_168,N_434);
xnor U6567 (N_6567,N_178,N_992);
xnor U6568 (N_6568,N_2484,N_3935);
xor U6569 (N_6569,N_2967,N_2889);
or U6570 (N_6570,N_1469,N_3011);
or U6571 (N_6571,N_1172,N_513);
and U6572 (N_6572,N_3400,N_3068);
nand U6573 (N_6573,N_3623,N_102);
or U6574 (N_6574,N_639,N_563);
and U6575 (N_6575,N_1358,N_126);
nand U6576 (N_6576,N_618,N_2292);
xnor U6577 (N_6577,N_2709,N_173);
or U6578 (N_6578,N_453,N_1208);
nor U6579 (N_6579,N_73,N_3814);
or U6580 (N_6580,N_3050,N_3398);
or U6581 (N_6581,N_1846,N_531);
or U6582 (N_6582,N_143,N_2620);
and U6583 (N_6583,N_144,N_3145);
xnor U6584 (N_6584,N_3739,N_3268);
nor U6585 (N_6585,N_959,N_3665);
xor U6586 (N_6586,N_842,N_3781);
nand U6587 (N_6587,N_1101,N_560);
xnor U6588 (N_6588,N_1130,N_3432);
nand U6589 (N_6589,N_473,N_1527);
nand U6590 (N_6590,N_2447,N_2235);
or U6591 (N_6591,N_2278,N_1532);
or U6592 (N_6592,N_2775,N_3706);
nor U6593 (N_6593,N_3987,N_586);
and U6594 (N_6594,N_1131,N_754);
nand U6595 (N_6595,N_1245,N_1818);
or U6596 (N_6596,N_856,N_3550);
nor U6597 (N_6597,N_990,N_1933);
or U6598 (N_6598,N_134,N_2311);
nand U6599 (N_6599,N_1202,N_1838);
nor U6600 (N_6600,N_2293,N_1367);
and U6601 (N_6601,N_325,N_3271);
nor U6602 (N_6602,N_3723,N_2786);
and U6603 (N_6603,N_3563,N_3914);
xnor U6604 (N_6604,N_1153,N_1488);
nand U6605 (N_6605,N_1568,N_1617);
xor U6606 (N_6606,N_1894,N_108);
nand U6607 (N_6607,N_3772,N_1960);
nor U6608 (N_6608,N_3845,N_3629);
and U6609 (N_6609,N_3428,N_962);
nor U6610 (N_6610,N_1635,N_899);
nor U6611 (N_6611,N_1165,N_386);
nor U6612 (N_6612,N_1610,N_1079);
xnor U6613 (N_6613,N_792,N_3198);
nand U6614 (N_6614,N_364,N_3396);
or U6615 (N_6615,N_2898,N_445);
and U6616 (N_6616,N_2015,N_3435);
and U6617 (N_6617,N_601,N_3519);
or U6618 (N_6618,N_682,N_3903);
and U6619 (N_6619,N_1342,N_3553);
or U6620 (N_6620,N_1002,N_3625);
and U6621 (N_6621,N_3699,N_3738);
nor U6622 (N_6622,N_1405,N_1178);
and U6623 (N_6623,N_1995,N_1883);
xnor U6624 (N_6624,N_1814,N_2356);
nor U6625 (N_6625,N_630,N_126);
and U6626 (N_6626,N_610,N_3658);
nand U6627 (N_6627,N_3875,N_405);
or U6628 (N_6628,N_3245,N_228);
nor U6629 (N_6629,N_703,N_427);
or U6630 (N_6630,N_684,N_10);
or U6631 (N_6631,N_2535,N_1240);
and U6632 (N_6632,N_3543,N_2292);
and U6633 (N_6633,N_2715,N_3975);
and U6634 (N_6634,N_544,N_2939);
or U6635 (N_6635,N_3318,N_3346);
and U6636 (N_6636,N_3458,N_866);
or U6637 (N_6637,N_1941,N_866);
or U6638 (N_6638,N_2811,N_2223);
and U6639 (N_6639,N_527,N_485);
nor U6640 (N_6640,N_3383,N_3631);
xor U6641 (N_6641,N_1664,N_3556);
nand U6642 (N_6642,N_726,N_501);
nand U6643 (N_6643,N_1495,N_1831);
xnor U6644 (N_6644,N_918,N_1722);
nor U6645 (N_6645,N_3458,N_3923);
xnor U6646 (N_6646,N_984,N_334);
nand U6647 (N_6647,N_3099,N_1775);
nor U6648 (N_6648,N_948,N_2910);
xnor U6649 (N_6649,N_1235,N_2827);
nor U6650 (N_6650,N_2725,N_461);
xor U6651 (N_6651,N_485,N_869);
xor U6652 (N_6652,N_2535,N_772);
nand U6653 (N_6653,N_3660,N_2308);
xnor U6654 (N_6654,N_1478,N_3767);
nand U6655 (N_6655,N_400,N_445);
nor U6656 (N_6656,N_701,N_932);
nand U6657 (N_6657,N_2861,N_860);
or U6658 (N_6658,N_1206,N_2342);
or U6659 (N_6659,N_3855,N_1612);
nor U6660 (N_6660,N_570,N_3617);
and U6661 (N_6661,N_210,N_1761);
or U6662 (N_6662,N_1658,N_340);
nand U6663 (N_6663,N_2986,N_1280);
or U6664 (N_6664,N_3927,N_2443);
xnor U6665 (N_6665,N_1285,N_2226);
or U6666 (N_6666,N_2494,N_3511);
nand U6667 (N_6667,N_664,N_610);
or U6668 (N_6668,N_3689,N_590);
and U6669 (N_6669,N_225,N_3223);
nand U6670 (N_6670,N_2568,N_3258);
xor U6671 (N_6671,N_3788,N_905);
nand U6672 (N_6672,N_2100,N_2218);
nor U6673 (N_6673,N_1573,N_3810);
and U6674 (N_6674,N_3328,N_1363);
or U6675 (N_6675,N_3851,N_3592);
nand U6676 (N_6676,N_293,N_2196);
nand U6677 (N_6677,N_721,N_898);
and U6678 (N_6678,N_2393,N_2072);
or U6679 (N_6679,N_3053,N_538);
xor U6680 (N_6680,N_3049,N_1477);
nor U6681 (N_6681,N_3144,N_1929);
or U6682 (N_6682,N_1863,N_759);
nor U6683 (N_6683,N_1599,N_1705);
nand U6684 (N_6684,N_1634,N_1495);
or U6685 (N_6685,N_1725,N_1408);
and U6686 (N_6686,N_2507,N_3346);
nor U6687 (N_6687,N_3394,N_598);
and U6688 (N_6688,N_2843,N_2804);
or U6689 (N_6689,N_130,N_70);
xor U6690 (N_6690,N_697,N_636);
nand U6691 (N_6691,N_1778,N_2692);
or U6692 (N_6692,N_3285,N_3141);
or U6693 (N_6693,N_3165,N_2772);
xnor U6694 (N_6694,N_2307,N_1261);
nor U6695 (N_6695,N_3429,N_2134);
or U6696 (N_6696,N_3159,N_1631);
nand U6697 (N_6697,N_733,N_1662);
or U6698 (N_6698,N_2117,N_3637);
nor U6699 (N_6699,N_1337,N_886);
xor U6700 (N_6700,N_3692,N_2964);
nand U6701 (N_6701,N_1522,N_617);
and U6702 (N_6702,N_1477,N_2662);
nand U6703 (N_6703,N_2290,N_235);
and U6704 (N_6704,N_1462,N_1625);
nor U6705 (N_6705,N_589,N_1172);
nor U6706 (N_6706,N_2676,N_1941);
xnor U6707 (N_6707,N_3353,N_2299);
nand U6708 (N_6708,N_2366,N_2113);
xnor U6709 (N_6709,N_3647,N_89);
nand U6710 (N_6710,N_2563,N_2608);
and U6711 (N_6711,N_3063,N_3915);
xnor U6712 (N_6712,N_1877,N_1860);
xor U6713 (N_6713,N_2145,N_3099);
nand U6714 (N_6714,N_1915,N_3137);
or U6715 (N_6715,N_1523,N_3686);
xor U6716 (N_6716,N_46,N_3407);
and U6717 (N_6717,N_3560,N_2906);
or U6718 (N_6718,N_1830,N_3622);
or U6719 (N_6719,N_1953,N_1152);
and U6720 (N_6720,N_904,N_1487);
or U6721 (N_6721,N_2433,N_1133);
xor U6722 (N_6722,N_2059,N_3464);
nor U6723 (N_6723,N_1266,N_3008);
nor U6724 (N_6724,N_3028,N_1985);
and U6725 (N_6725,N_1853,N_3223);
nand U6726 (N_6726,N_490,N_3660);
nor U6727 (N_6727,N_3816,N_35);
xor U6728 (N_6728,N_3838,N_2586);
or U6729 (N_6729,N_2885,N_2432);
nor U6730 (N_6730,N_3707,N_1608);
xor U6731 (N_6731,N_3485,N_1716);
nor U6732 (N_6732,N_3274,N_2912);
or U6733 (N_6733,N_119,N_3802);
nand U6734 (N_6734,N_894,N_2237);
xnor U6735 (N_6735,N_2867,N_2905);
nor U6736 (N_6736,N_77,N_1459);
nor U6737 (N_6737,N_432,N_3923);
xor U6738 (N_6738,N_840,N_566);
or U6739 (N_6739,N_2383,N_2755);
nand U6740 (N_6740,N_13,N_914);
or U6741 (N_6741,N_2977,N_1983);
nand U6742 (N_6742,N_897,N_2515);
or U6743 (N_6743,N_22,N_2974);
or U6744 (N_6744,N_2854,N_3743);
xor U6745 (N_6745,N_578,N_2769);
nor U6746 (N_6746,N_3925,N_3651);
nand U6747 (N_6747,N_1524,N_3802);
xor U6748 (N_6748,N_333,N_1718);
nor U6749 (N_6749,N_2908,N_2084);
xnor U6750 (N_6750,N_1794,N_619);
nand U6751 (N_6751,N_3765,N_1759);
or U6752 (N_6752,N_3975,N_156);
xor U6753 (N_6753,N_2715,N_3575);
or U6754 (N_6754,N_2286,N_1243);
nor U6755 (N_6755,N_2190,N_1354);
nor U6756 (N_6756,N_3663,N_3944);
nand U6757 (N_6757,N_1246,N_2333);
or U6758 (N_6758,N_2109,N_3001);
or U6759 (N_6759,N_2823,N_2947);
nand U6760 (N_6760,N_3318,N_1792);
nand U6761 (N_6761,N_3678,N_1749);
or U6762 (N_6762,N_1206,N_2482);
nor U6763 (N_6763,N_281,N_3255);
xor U6764 (N_6764,N_2845,N_1662);
and U6765 (N_6765,N_761,N_2662);
nand U6766 (N_6766,N_691,N_2324);
nor U6767 (N_6767,N_3221,N_1042);
nor U6768 (N_6768,N_1995,N_647);
xor U6769 (N_6769,N_3144,N_1053);
nand U6770 (N_6770,N_827,N_2729);
nor U6771 (N_6771,N_872,N_2751);
and U6772 (N_6772,N_414,N_1426);
and U6773 (N_6773,N_1360,N_18);
nor U6774 (N_6774,N_3384,N_3933);
or U6775 (N_6775,N_3164,N_2659);
nor U6776 (N_6776,N_1469,N_3990);
nor U6777 (N_6777,N_2150,N_457);
nor U6778 (N_6778,N_3143,N_3960);
xnor U6779 (N_6779,N_2486,N_2233);
or U6780 (N_6780,N_1221,N_2642);
nand U6781 (N_6781,N_2282,N_1723);
nor U6782 (N_6782,N_1863,N_3559);
and U6783 (N_6783,N_650,N_1880);
nor U6784 (N_6784,N_2800,N_2176);
nand U6785 (N_6785,N_456,N_545);
xor U6786 (N_6786,N_3618,N_3009);
nor U6787 (N_6787,N_1933,N_1202);
nor U6788 (N_6788,N_2875,N_3345);
xor U6789 (N_6789,N_69,N_3110);
or U6790 (N_6790,N_3966,N_2259);
nand U6791 (N_6791,N_2385,N_2892);
nor U6792 (N_6792,N_3951,N_727);
or U6793 (N_6793,N_1986,N_2101);
nand U6794 (N_6794,N_355,N_327);
or U6795 (N_6795,N_1254,N_3892);
or U6796 (N_6796,N_545,N_2145);
xnor U6797 (N_6797,N_489,N_923);
or U6798 (N_6798,N_3501,N_348);
nor U6799 (N_6799,N_2778,N_388);
nand U6800 (N_6800,N_2562,N_1209);
nor U6801 (N_6801,N_398,N_1190);
nand U6802 (N_6802,N_3492,N_1032);
or U6803 (N_6803,N_520,N_678);
nand U6804 (N_6804,N_1693,N_3295);
or U6805 (N_6805,N_3324,N_2880);
nor U6806 (N_6806,N_359,N_736);
xnor U6807 (N_6807,N_3706,N_948);
xor U6808 (N_6808,N_3093,N_2755);
nor U6809 (N_6809,N_254,N_3425);
xor U6810 (N_6810,N_1266,N_79);
nor U6811 (N_6811,N_3028,N_1412);
nor U6812 (N_6812,N_3059,N_1740);
or U6813 (N_6813,N_740,N_1772);
and U6814 (N_6814,N_2767,N_1358);
nand U6815 (N_6815,N_2525,N_2376);
nor U6816 (N_6816,N_2792,N_286);
or U6817 (N_6817,N_1946,N_1239);
nand U6818 (N_6818,N_1652,N_2848);
nand U6819 (N_6819,N_962,N_2627);
xnor U6820 (N_6820,N_2698,N_2809);
nand U6821 (N_6821,N_727,N_2097);
xnor U6822 (N_6822,N_437,N_3926);
xnor U6823 (N_6823,N_1500,N_1493);
nand U6824 (N_6824,N_1048,N_2860);
and U6825 (N_6825,N_798,N_2543);
xnor U6826 (N_6826,N_2454,N_1705);
nor U6827 (N_6827,N_3932,N_3626);
or U6828 (N_6828,N_3645,N_243);
and U6829 (N_6829,N_3292,N_2709);
nand U6830 (N_6830,N_493,N_3724);
xor U6831 (N_6831,N_2357,N_1953);
and U6832 (N_6832,N_154,N_3198);
nand U6833 (N_6833,N_3483,N_3398);
nand U6834 (N_6834,N_1148,N_3884);
xnor U6835 (N_6835,N_2703,N_271);
xnor U6836 (N_6836,N_1902,N_452);
and U6837 (N_6837,N_1482,N_242);
or U6838 (N_6838,N_3308,N_1035);
nor U6839 (N_6839,N_3317,N_2865);
nor U6840 (N_6840,N_2793,N_1026);
or U6841 (N_6841,N_3453,N_2321);
nor U6842 (N_6842,N_3378,N_1011);
xor U6843 (N_6843,N_218,N_951);
or U6844 (N_6844,N_2504,N_2637);
or U6845 (N_6845,N_945,N_3615);
and U6846 (N_6846,N_1556,N_3580);
or U6847 (N_6847,N_3130,N_3996);
and U6848 (N_6848,N_1874,N_3781);
xor U6849 (N_6849,N_981,N_3543);
xnor U6850 (N_6850,N_3555,N_2330);
and U6851 (N_6851,N_1203,N_2680);
or U6852 (N_6852,N_290,N_154);
nand U6853 (N_6853,N_1150,N_2753);
nor U6854 (N_6854,N_1436,N_3453);
nor U6855 (N_6855,N_785,N_419);
and U6856 (N_6856,N_3386,N_1893);
xor U6857 (N_6857,N_3639,N_481);
nand U6858 (N_6858,N_1732,N_3261);
xor U6859 (N_6859,N_3803,N_1640);
nand U6860 (N_6860,N_2150,N_2017);
or U6861 (N_6861,N_1375,N_2014);
nor U6862 (N_6862,N_3632,N_1693);
and U6863 (N_6863,N_1605,N_3482);
xor U6864 (N_6864,N_410,N_2256);
and U6865 (N_6865,N_1293,N_1827);
nor U6866 (N_6866,N_2293,N_2123);
xnor U6867 (N_6867,N_2148,N_3133);
nor U6868 (N_6868,N_3445,N_348);
nor U6869 (N_6869,N_139,N_3042);
nor U6870 (N_6870,N_1146,N_2476);
nand U6871 (N_6871,N_1825,N_322);
xor U6872 (N_6872,N_675,N_2632);
or U6873 (N_6873,N_2687,N_2638);
or U6874 (N_6874,N_3010,N_655);
nand U6875 (N_6875,N_3402,N_3619);
nor U6876 (N_6876,N_316,N_2737);
and U6877 (N_6877,N_1720,N_1435);
nor U6878 (N_6878,N_1927,N_254);
nand U6879 (N_6879,N_1640,N_3759);
or U6880 (N_6880,N_2101,N_3464);
nor U6881 (N_6881,N_1739,N_2244);
nor U6882 (N_6882,N_3651,N_3165);
xor U6883 (N_6883,N_2401,N_3748);
or U6884 (N_6884,N_3287,N_2768);
xnor U6885 (N_6885,N_118,N_3597);
nand U6886 (N_6886,N_1316,N_3228);
xnor U6887 (N_6887,N_961,N_263);
or U6888 (N_6888,N_3763,N_3212);
nand U6889 (N_6889,N_1724,N_1533);
nor U6890 (N_6890,N_1886,N_3091);
or U6891 (N_6891,N_2919,N_3361);
xor U6892 (N_6892,N_1600,N_2491);
nand U6893 (N_6893,N_1099,N_3516);
and U6894 (N_6894,N_1191,N_777);
nand U6895 (N_6895,N_593,N_396);
or U6896 (N_6896,N_775,N_3247);
nor U6897 (N_6897,N_3339,N_2987);
nor U6898 (N_6898,N_2864,N_3789);
nor U6899 (N_6899,N_513,N_761);
nor U6900 (N_6900,N_971,N_3708);
xnor U6901 (N_6901,N_3624,N_998);
nand U6902 (N_6902,N_639,N_171);
nor U6903 (N_6903,N_3292,N_1447);
xnor U6904 (N_6904,N_571,N_3389);
nand U6905 (N_6905,N_56,N_856);
nor U6906 (N_6906,N_165,N_2818);
or U6907 (N_6907,N_3249,N_995);
or U6908 (N_6908,N_3997,N_2406);
nand U6909 (N_6909,N_1926,N_3834);
nor U6910 (N_6910,N_2854,N_915);
and U6911 (N_6911,N_1635,N_1881);
xor U6912 (N_6912,N_2097,N_2699);
nand U6913 (N_6913,N_3737,N_1766);
or U6914 (N_6914,N_3628,N_947);
and U6915 (N_6915,N_401,N_313);
and U6916 (N_6916,N_1810,N_1231);
or U6917 (N_6917,N_133,N_2745);
and U6918 (N_6918,N_2475,N_113);
nand U6919 (N_6919,N_866,N_3607);
or U6920 (N_6920,N_3538,N_803);
and U6921 (N_6921,N_2246,N_3691);
and U6922 (N_6922,N_1702,N_477);
xor U6923 (N_6923,N_2628,N_3819);
nor U6924 (N_6924,N_2054,N_366);
xor U6925 (N_6925,N_1788,N_837);
and U6926 (N_6926,N_1924,N_3261);
nor U6927 (N_6927,N_1535,N_725);
nand U6928 (N_6928,N_3592,N_2917);
nor U6929 (N_6929,N_1753,N_832);
xnor U6930 (N_6930,N_1858,N_2020);
and U6931 (N_6931,N_262,N_1420);
and U6932 (N_6932,N_2048,N_2645);
xor U6933 (N_6933,N_1362,N_1287);
xnor U6934 (N_6934,N_3843,N_3652);
nand U6935 (N_6935,N_3542,N_2892);
xor U6936 (N_6936,N_3288,N_3268);
and U6937 (N_6937,N_3964,N_977);
nor U6938 (N_6938,N_2417,N_3582);
nor U6939 (N_6939,N_2227,N_1980);
nand U6940 (N_6940,N_2261,N_3025);
or U6941 (N_6941,N_1198,N_982);
or U6942 (N_6942,N_1682,N_3584);
xnor U6943 (N_6943,N_3471,N_543);
xor U6944 (N_6944,N_2352,N_3943);
xor U6945 (N_6945,N_1974,N_971);
nor U6946 (N_6946,N_3434,N_3687);
nand U6947 (N_6947,N_2790,N_3604);
xor U6948 (N_6948,N_768,N_2717);
xnor U6949 (N_6949,N_22,N_620);
nor U6950 (N_6950,N_2674,N_1024);
nor U6951 (N_6951,N_1135,N_2310);
and U6952 (N_6952,N_1535,N_3171);
nand U6953 (N_6953,N_3577,N_688);
or U6954 (N_6954,N_3603,N_3861);
xor U6955 (N_6955,N_3467,N_2020);
and U6956 (N_6956,N_3966,N_2888);
nor U6957 (N_6957,N_3909,N_2967);
nand U6958 (N_6958,N_1654,N_997);
nand U6959 (N_6959,N_3861,N_438);
xor U6960 (N_6960,N_3629,N_1799);
and U6961 (N_6961,N_3019,N_1403);
and U6962 (N_6962,N_278,N_2605);
nor U6963 (N_6963,N_3447,N_3951);
xnor U6964 (N_6964,N_1343,N_3155);
nand U6965 (N_6965,N_247,N_1648);
or U6966 (N_6966,N_1460,N_719);
or U6967 (N_6967,N_3777,N_3679);
xnor U6968 (N_6968,N_979,N_1354);
nor U6969 (N_6969,N_1891,N_1920);
nor U6970 (N_6970,N_3190,N_1612);
or U6971 (N_6971,N_1802,N_903);
nor U6972 (N_6972,N_3378,N_2936);
xor U6973 (N_6973,N_3452,N_596);
and U6974 (N_6974,N_2150,N_2607);
nor U6975 (N_6975,N_3301,N_1943);
and U6976 (N_6976,N_286,N_2477);
and U6977 (N_6977,N_1357,N_2765);
xor U6978 (N_6978,N_2600,N_503);
nand U6979 (N_6979,N_530,N_2856);
nand U6980 (N_6980,N_3542,N_281);
nor U6981 (N_6981,N_833,N_1671);
or U6982 (N_6982,N_1864,N_416);
nor U6983 (N_6983,N_1937,N_3145);
nand U6984 (N_6984,N_896,N_277);
nor U6985 (N_6985,N_3209,N_1403);
nand U6986 (N_6986,N_2973,N_1051);
and U6987 (N_6987,N_1548,N_1871);
and U6988 (N_6988,N_1475,N_550);
xor U6989 (N_6989,N_764,N_3043);
xor U6990 (N_6990,N_2290,N_3152);
nand U6991 (N_6991,N_3579,N_151);
nor U6992 (N_6992,N_604,N_1749);
or U6993 (N_6993,N_3832,N_1279);
and U6994 (N_6994,N_2760,N_465);
nor U6995 (N_6995,N_1432,N_1631);
nor U6996 (N_6996,N_2027,N_1547);
nor U6997 (N_6997,N_2713,N_321);
and U6998 (N_6998,N_1549,N_370);
nand U6999 (N_6999,N_3936,N_2557);
xor U7000 (N_7000,N_1347,N_1028);
nand U7001 (N_7001,N_1557,N_482);
nand U7002 (N_7002,N_38,N_2149);
xnor U7003 (N_7003,N_366,N_2027);
or U7004 (N_7004,N_1282,N_2307);
nor U7005 (N_7005,N_488,N_2428);
xnor U7006 (N_7006,N_749,N_1470);
or U7007 (N_7007,N_205,N_3403);
nor U7008 (N_7008,N_785,N_2382);
nor U7009 (N_7009,N_3368,N_1495);
nand U7010 (N_7010,N_257,N_2656);
nand U7011 (N_7011,N_914,N_2661);
nand U7012 (N_7012,N_3488,N_1970);
nor U7013 (N_7013,N_3573,N_2248);
or U7014 (N_7014,N_3809,N_3507);
xor U7015 (N_7015,N_514,N_840);
nor U7016 (N_7016,N_3219,N_964);
nor U7017 (N_7017,N_2389,N_1918);
xnor U7018 (N_7018,N_1477,N_2078);
and U7019 (N_7019,N_2081,N_80);
and U7020 (N_7020,N_319,N_610);
xor U7021 (N_7021,N_1177,N_630);
nor U7022 (N_7022,N_123,N_1701);
nor U7023 (N_7023,N_3493,N_1004);
xnor U7024 (N_7024,N_1887,N_1005);
nand U7025 (N_7025,N_2858,N_3411);
xor U7026 (N_7026,N_1313,N_2378);
xnor U7027 (N_7027,N_1146,N_3902);
xnor U7028 (N_7028,N_649,N_1881);
or U7029 (N_7029,N_283,N_1718);
nand U7030 (N_7030,N_1861,N_3486);
or U7031 (N_7031,N_1745,N_1239);
nor U7032 (N_7032,N_3534,N_2085);
and U7033 (N_7033,N_978,N_46);
or U7034 (N_7034,N_98,N_2829);
and U7035 (N_7035,N_3383,N_1554);
nor U7036 (N_7036,N_3308,N_1920);
or U7037 (N_7037,N_89,N_3102);
and U7038 (N_7038,N_3493,N_2958);
xnor U7039 (N_7039,N_2104,N_30);
nand U7040 (N_7040,N_1237,N_3705);
nor U7041 (N_7041,N_634,N_597);
or U7042 (N_7042,N_144,N_937);
and U7043 (N_7043,N_2575,N_1832);
and U7044 (N_7044,N_803,N_1858);
nor U7045 (N_7045,N_1830,N_486);
nand U7046 (N_7046,N_400,N_1099);
or U7047 (N_7047,N_1076,N_1549);
xnor U7048 (N_7048,N_3094,N_827);
and U7049 (N_7049,N_1032,N_2682);
nand U7050 (N_7050,N_692,N_1072);
nor U7051 (N_7051,N_2597,N_3274);
nor U7052 (N_7052,N_1552,N_1916);
and U7053 (N_7053,N_2071,N_1136);
nor U7054 (N_7054,N_827,N_1362);
or U7055 (N_7055,N_3774,N_2936);
or U7056 (N_7056,N_1103,N_1356);
and U7057 (N_7057,N_2819,N_47);
and U7058 (N_7058,N_2858,N_2689);
xor U7059 (N_7059,N_1139,N_1612);
xor U7060 (N_7060,N_712,N_3995);
and U7061 (N_7061,N_321,N_602);
or U7062 (N_7062,N_3791,N_808);
nand U7063 (N_7063,N_2348,N_3708);
xor U7064 (N_7064,N_1478,N_3342);
xor U7065 (N_7065,N_267,N_187);
nor U7066 (N_7066,N_3852,N_703);
and U7067 (N_7067,N_1372,N_3134);
or U7068 (N_7068,N_3254,N_5);
nor U7069 (N_7069,N_624,N_2749);
xnor U7070 (N_7070,N_1510,N_2727);
or U7071 (N_7071,N_3661,N_870);
nand U7072 (N_7072,N_2837,N_2291);
and U7073 (N_7073,N_162,N_487);
nor U7074 (N_7074,N_991,N_3625);
or U7075 (N_7075,N_3237,N_2218);
or U7076 (N_7076,N_2029,N_755);
or U7077 (N_7077,N_527,N_3913);
or U7078 (N_7078,N_3867,N_2579);
xnor U7079 (N_7079,N_2513,N_1668);
and U7080 (N_7080,N_2040,N_2850);
xnor U7081 (N_7081,N_2037,N_2555);
or U7082 (N_7082,N_382,N_2247);
nor U7083 (N_7083,N_2192,N_1798);
nand U7084 (N_7084,N_1310,N_657);
xnor U7085 (N_7085,N_590,N_1481);
and U7086 (N_7086,N_1046,N_2676);
or U7087 (N_7087,N_1961,N_2827);
xor U7088 (N_7088,N_1471,N_1532);
or U7089 (N_7089,N_377,N_1103);
nand U7090 (N_7090,N_2707,N_2382);
xor U7091 (N_7091,N_366,N_1247);
or U7092 (N_7092,N_2751,N_2969);
nand U7093 (N_7093,N_880,N_2568);
nand U7094 (N_7094,N_2879,N_2332);
xnor U7095 (N_7095,N_2329,N_2941);
or U7096 (N_7096,N_3723,N_1628);
nand U7097 (N_7097,N_2319,N_880);
or U7098 (N_7098,N_3401,N_249);
nor U7099 (N_7099,N_427,N_2501);
and U7100 (N_7100,N_1497,N_637);
nand U7101 (N_7101,N_2931,N_550);
nand U7102 (N_7102,N_3461,N_2855);
xor U7103 (N_7103,N_1420,N_3716);
xor U7104 (N_7104,N_2275,N_1175);
nor U7105 (N_7105,N_194,N_1830);
nand U7106 (N_7106,N_1294,N_1081);
nand U7107 (N_7107,N_268,N_3054);
nor U7108 (N_7108,N_3332,N_1969);
nor U7109 (N_7109,N_2047,N_873);
nor U7110 (N_7110,N_1488,N_1113);
xnor U7111 (N_7111,N_434,N_1333);
or U7112 (N_7112,N_2196,N_1926);
xnor U7113 (N_7113,N_1224,N_2427);
xor U7114 (N_7114,N_768,N_480);
nor U7115 (N_7115,N_3549,N_570);
nand U7116 (N_7116,N_564,N_2273);
nor U7117 (N_7117,N_3122,N_3298);
or U7118 (N_7118,N_1799,N_1547);
or U7119 (N_7119,N_1144,N_2522);
or U7120 (N_7120,N_1813,N_1208);
nor U7121 (N_7121,N_3686,N_623);
xnor U7122 (N_7122,N_2474,N_31);
or U7123 (N_7123,N_2948,N_3921);
and U7124 (N_7124,N_3408,N_2707);
or U7125 (N_7125,N_2419,N_2389);
nor U7126 (N_7126,N_1005,N_1555);
or U7127 (N_7127,N_3514,N_3076);
xor U7128 (N_7128,N_2426,N_1839);
xor U7129 (N_7129,N_3308,N_1443);
nand U7130 (N_7130,N_1254,N_2570);
or U7131 (N_7131,N_664,N_3348);
xnor U7132 (N_7132,N_1855,N_2482);
or U7133 (N_7133,N_2864,N_2516);
and U7134 (N_7134,N_3135,N_372);
xnor U7135 (N_7135,N_2035,N_1747);
and U7136 (N_7136,N_2207,N_672);
or U7137 (N_7137,N_3937,N_157);
nor U7138 (N_7138,N_1005,N_2925);
nor U7139 (N_7139,N_1409,N_935);
xnor U7140 (N_7140,N_1439,N_2217);
or U7141 (N_7141,N_1888,N_161);
xnor U7142 (N_7142,N_3253,N_2324);
nor U7143 (N_7143,N_270,N_155);
nand U7144 (N_7144,N_1071,N_337);
nand U7145 (N_7145,N_2537,N_2535);
nand U7146 (N_7146,N_1971,N_2514);
nand U7147 (N_7147,N_1709,N_230);
nor U7148 (N_7148,N_3652,N_3190);
nand U7149 (N_7149,N_1530,N_354);
nand U7150 (N_7150,N_3732,N_3377);
xnor U7151 (N_7151,N_3752,N_26);
xor U7152 (N_7152,N_943,N_3789);
nor U7153 (N_7153,N_839,N_3172);
xor U7154 (N_7154,N_3611,N_758);
and U7155 (N_7155,N_3731,N_3748);
nand U7156 (N_7156,N_583,N_1808);
and U7157 (N_7157,N_3489,N_1245);
and U7158 (N_7158,N_1973,N_3946);
or U7159 (N_7159,N_777,N_3169);
nand U7160 (N_7160,N_622,N_995);
or U7161 (N_7161,N_1015,N_932);
or U7162 (N_7162,N_131,N_3061);
nor U7163 (N_7163,N_2847,N_894);
nand U7164 (N_7164,N_2076,N_1678);
nand U7165 (N_7165,N_1379,N_1376);
nand U7166 (N_7166,N_775,N_1180);
nand U7167 (N_7167,N_3370,N_3687);
and U7168 (N_7168,N_2341,N_706);
and U7169 (N_7169,N_1979,N_1270);
xor U7170 (N_7170,N_2420,N_1847);
nor U7171 (N_7171,N_1988,N_3172);
nand U7172 (N_7172,N_2974,N_3355);
xnor U7173 (N_7173,N_2581,N_3754);
nor U7174 (N_7174,N_3449,N_1021);
nor U7175 (N_7175,N_3765,N_3634);
nor U7176 (N_7176,N_239,N_3228);
or U7177 (N_7177,N_2171,N_3863);
nor U7178 (N_7178,N_2625,N_2671);
nor U7179 (N_7179,N_2790,N_1238);
nand U7180 (N_7180,N_2451,N_2724);
or U7181 (N_7181,N_2550,N_3608);
nor U7182 (N_7182,N_2429,N_2759);
or U7183 (N_7183,N_1577,N_1389);
or U7184 (N_7184,N_825,N_3396);
or U7185 (N_7185,N_3349,N_751);
and U7186 (N_7186,N_1237,N_239);
nand U7187 (N_7187,N_949,N_3136);
nor U7188 (N_7188,N_3691,N_28);
nand U7189 (N_7189,N_2902,N_823);
nor U7190 (N_7190,N_3686,N_2018);
nand U7191 (N_7191,N_2216,N_1651);
nor U7192 (N_7192,N_3354,N_3151);
nor U7193 (N_7193,N_1675,N_1462);
nand U7194 (N_7194,N_639,N_3948);
or U7195 (N_7195,N_566,N_2808);
xnor U7196 (N_7196,N_1734,N_3641);
nor U7197 (N_7197,N_904,N_574);
nor U7198 (N_7198,N_3649,N_529);
nor U7199 (N_7199,N_2723,N_466);
nand U7200 (N_7200,N_1488,N_2163);
nor U7201 (N_7201,N_3813,N_3090);
xor U7202 (N_7202,N_0,N_2687);
or U7203 (N_7203,N_3714,N_235);
or U7204 (N_7204,N_1256,N_1891);
nand U7205 (N_7205,N_1841,N_1070);
and U7206 (N_7206,N_952,N_3498);
nor U7207 (N_7207,N_246,N_3344);
and U7208 (N_7208,N_2002,N_3415);
nand U7209 (N_7209,N_612,N_645);
nand U7210 (N_7210,N_656,N_3362);
nand U7211 (N_7211,N_949,N_2609);
and U7212 (N_7212,N_171,N_3607);
nand U7213 (N_7213,N_3463,N_1755);
nor U7214 (N_7214,N_2674,N_2942);
nor U7215 (N_7215,N_3986,N_2893);
nand U7216 (N_7216,N_2938,N_457);
or U7217 (N_7217,N_2142,N_124);
or U7218 (N_7218,N_2553,N_1819);
xor U7219 (N_7219,N_857,N_2017);
and U7220 (N_7220,N_198,N_2281);
xor U7221 (N_7221,N_1381,N_3023);
xnor U7222 (N_7222,N_2345,N_1399);
nor U7223 (N_7223,N_3429,N_1126);
nand U7224 (N_7224,N_3716,N_2308);
and U7225 (N_7225,N_3783,N_3236);
xor U7226 (N_7226,N_905,N_1734);
and U7227 (N_7227,N_3624,N_3659);
and U7228 (N_7228,N_905,N_3387);
nor U7229 (N_7229,N_3847,N_3017);
and U7230 (N_7230,N_2456,N_436);
nor U7231 (N_7231,N_174,N_1929);
nor U7232 (N_7232,N_3727,N_3502);
xnor U7233 (N_7233,N_2881,N_1882);
nor U7234 (N_7234,N_2539,N_3879);
or U7235 (N_7235,N_1332,N_1522);
nand U7236 (N_7236,N_338,N_3745);
or U7237 (N_7237,N_1631,N_3553);
nand U7238 (N_7238,N_700,N_2018);
and U7239 (N_7239,N_1488,N_3454);
xnor U7240 (N_7240,N_3432,N_3813);
nor U7241 (N_7241,N_2884,N_896);
xnor U7242 (N_7242,N_188,N_783);
xnor U7243 (N_7243,N_1105,N_3278);
xnor U7244 (N_7244,N_3190,N_933);
and U7245 (N_7245,N_1968,N_529);
and U7246 (N_7246,N_1116,N_2181);
xor U7247 (N_7247,N_3224,N_3025);
xor U7248 (N_7248,N_2979,N_681);
nor U7249 (N_7249,N_3022,N_2357);
nor U7250 (N_7250,N_2051,N_2265);
nor U7251 (N_7251,N_682,N_2528);
and U7252 (N_7252,N_2714,N_1979);
or U7253 (N_7253,N_2588,N_1626);
nor U7254 (N_7254,N_1620,N_808);
or U7255 (N_7255,N_1934,N_3965);
or U7256 (N_7256,N_2102,N_2219);
or U7257 (N_7257,N_679,N_2388);
nand U7258 (N_7258,N_3433,N_3662);
xor U7259 (N_7259,N_1002,N_649);
nor U7260 (N_7260,N_1703,N_2050);
xor U7261 (N_7261,N_1081,N_3013);
nand U7262 (N_7262,N_1242,N_699);
or U7263 (N_7263,N_1716,N_1757);
and U7264 (N_7264,N_3948,N_2797);
xnor U7265 (N_7265,N_3230,N_3328);
nor U7266 (N_7266,N_3874,N_2813);
nand U7267 (N_7267,N_407,N_965);
and U7268 (N_7268,N_360,N_3791);
nor U7269 (N_7269,N_410,N_1922);
or U7270 (N_7270,N_469,N_3711);
or U7271 (N_7271,N_3076,N_3128);
nor U7272 (N_7272,N_1354,N_1579);
xor U7273 (N_7273,N_2457,N_21);
and U7274 (N_7274,N_3253,N_821);
or U7275 (N_7275,N_3633,N_17);
nor U7276 (N_7276,N_3235,N_3273);
nand U7277 (N_7277,N_657,N_3049);
nor U7278 (N_7278,N_1943,N_1597);
nor U7279 (N_7279,N_1401,N_1001);
or U7280 (N_7280,N_2441,N_3523);
nor U7281 (N_7281,N_246,N_1668);
nand U7282 (N_7282,N_408,N_2498);
nand U7283 (N_7283,N_3045,N_377);
nor U7284 (N_7284,N_506,N_1354);
or U7285 (N_7285,N_20,N_2767);
nor U7286 (N_7286,N_1421,N_2015);
and U7287 (N_7287,N_674,N_13);
xor U7288 (N_7288,N_160,N_3710);
nor U7289 (N_7289,N_2453,N_1203);
or U7290 (N_7290,N_3887,N_2237);
nor U7291 (N_7291,N_3893,N_3488);
and U7292 (N_7292,N_48,N_1436);
xnor U7293 (N_7293,N_2737,N_1095);
nand U7294 (N_7294,N_841,N_3027);
and U7295 (N_7295,N_2614,N_2982);
and U7296 (N_7296,N_1744,N_3859);
or U7297 (N_7297,N_1966,N_3617);
xnor U7298 (N_7298,N_565,N_3865);
xnor U7299 (N_7299,N_3025,N_2499);
nand U7300 (N_7300,N_689,N_406);
or U7301 (N_7301,N_2455,N_1984);
xnor U7302 (N_7302,N_1306,N_3560);
xnor U7303 (N_7303,N_2772,N_600);
nor U7304 (N_7304,N_326,N_2354);
and U7305 (N_7305,N_1235,N_1137);
xnor U7306 (N_7306,N_3019,N_1023);
or U7307 (N_7307,N_3004,N_714);
and U7308 (N_7308,N_2299,N_1158);
and U7309 (N_7309,N_3669,N_83);
or U7310 (N_7310,N_563,N_1545);
or U7311 (N_7311,N_2281,N_2689);
xor U7312 (N_7312,N_1000,N_817);
nor U7313 (N_7313,N_2771,N_608);
and U7314 (N_7314,N_3417,N_3795);
nand U7315 (N_7315,N_3378,N_559);
and U7316 (N_7316,N_292,N_2979);
nor U7317 (N_7317,N_3096,N_944);
nor U7318 (N_7318,N_2277,N_2598);
nor U7319 (N_7319,N_2163,N_1853);
nand U7320 (N_7320,N_3950,N_3697);
and U7321 (N_7321,N_851,N_3703);
or U7322 (N_7322,N_78,N_2444);
nand U7323 (N_7323,N_719,N_1452);
xnor U7324 (N_7324,N_1518,N_1716);
and U7325 (N_7325,N_3852,N_1153);
nor U7326 (N_7326,N_2394,N_372);
xnor U7327 (N_7327,N_1204,N_3920);
nor U7328 (N_7328,N_3583,N_2291);
nand U7329 (N_7329,N_3303,N_3616);
xor U7330 (N_7330,N_1750,N_2620);
nor U7331 (N_7331,N_3454,N_3466);
xor U7332 (N_7332,N_3963,N_997);
nor U7333 (N_7333,N_398,N_2066);
and U7334 (N_7334,N_1740,N_3807);
xnor U7335 (N_7335,N_749,N_3889);
nand U7336 (N_7336,N_2814,N_1994);
nor U7337 (N_7337,N_2692,N_1465);
xor U7338 (N_7338,N_1231,N_3045);
or U7339 (N_7339,N_319,N_2616);
xnor U7340 (N_7340,N_1308,N_2494);
nor U7341 (N_7341,N_3090,N_2453);
xor U7342 (N_7342,N_1096,N_2263);
and U7343 (N_7343,N_3421,N_393);
or U7344 (N_7344,N_3168,N_2168);
xor U7345 (N_7345,N_3020,N_3888);
xnor U7346 (N_7346,N_3596,N_329);
or U7347 (N_7347,N_3794,N_3092);
nand U7348 (N_7348,N_3795,N_3334);
and U7349 (N_7349,N_1839,N_1186);
nand U7350 (N_7350,N_3591,N_2065);
nand U7351 (N_7351,N_2250,N_2212);
nor U7352 (N_7352,N_1590,N_2811);
nor U7353 (N_7353,N_3832,N_81);
xor U7354 (N_7354,N_689,N_2803);
or U7355 (N_7355,N_32,N_3014);
nand U7356 (N_7356,N_1232,N_1435);
and U7357 (N_7357,N_817,N_1748);
nor U7358 (N_7358,N_3234,N_1998);
xnor U7359 (N_7359,N_1172,N_795);
and U7360 (N_7360,N_2907,N_51);
and U7361 (N_7361,N_2332,N_383);
nand U7362 (N_7362,N_119,N_3958);
nor U7363 (N_7363,N_3552,N_3073);
xor U7364 (N_7364,N_680,N_1121);
nand U7365 (N_7365,N_588,N_5);
nand U7366 (N_7366,N_3021,N_1397);
and U7367 (N_7367,N_3628,N_2373);
xor U7368 (N_7368,N_2283,N_595);
and U7369 (N_7369,N_1234,N_236);
and U7370 (N_7370,N_1708,N_1147);
or U7371 (N_7371,N_1968,N_342);
nand U7372 (N_7372,N_3074,N_2797);
nor U7373 (N_7373,N_2711,N_718);
and U7374 (N_7374,N_3342,N_2282);
and U7375 (N_7375,N_2399,N_605);
nor U7376 (N_7376,N_661,N_301);
or U7377 (N_7377,N_3794,N_3720);
and U7378 (N_7378,N_3214,N_2934);
nand U7379 (N_7379,N_3598,N_2112);
or U7380 (N_7380,N_3035,N_1306);
nor U7381 (N_7381,N_3045,N_1758);
or U7382 (N_7382,N_1067,N_3093);
xnor U7383 (N_7383,N_3038,N_1634);
nor U7384 (N_7384,N_369,N_355);
xor U7385 (N_7385,N_1880,N_490);
and U7386 (N_7386,N_1908,N_1462);
xor U7387 (N_7387,N_1025,N_3136);
nor U7388 (N_7388,N_181,N_3167);
or U7389 (N_7389,N_322,N_3356);
nand U7390 (N_7390,N_3075,N_0);
or U7391 (N_7391,N_3534,N_862);
and U7392 (N_7392,N_3682,N_1483);
or U7393 (N_7393,N_3843,N_1898);
xnor U7394 (N_7394,N_3085,N_1964);
xnor U7395 (N_7395,N_2779,N_2511);
xor U7396 (N_7396,N_1153,N_776);
nor U7397 (N_7397,N_268,N_2621);
xnor U7398 (N_7398,N_1120,N_2805);
nand U7399 (N_7399,N_1522,N_265);
or U7400 (N_7400,N_317,N_1230);
nor U7401 (N_7401,N_3582,N_3801);
or U7402 (N_7402,N_416,N_146);
or U7403 (N_7403,N_3551,N_1371);
and U7404 (N_7404,N_2404,N_242);
or U7405 (N_7405,N_2459,N_1380);
xor U7406 (N_7406,N_1948,N_3652);
xor U7407 (N_7407,N_2536,N_3084);
or U7408 (N_7408,N_2248,N_1969);
nor U7409 (N_7409,N_1040,N_496);
xor U7410 (N_7410,N_1970,N_1644);
nand U7411 (N_7411,N_3838,N_2866);
or U7412 (N_7412,N_3826,N_2092);
nand U7413 (N_7413,N_1172,N_114);
nand U7414 (N_7414,N_135,N_2038);
nand U7415 (N_7415,N_303,N_301);
and U7416 (N_7416,N_3337,N_2477);
nand U7417 (N_7417,N_3898,N_3572);
xnor U7418 (N_7418,N_3186,N_1723);
or U7419 (N_7419,N_1549,N_2652);
xnor U7420 (N_7420,N_3760,N_3708);
nand U7421 (N_7421,N_3092,N_2010);
nor U7422 (N_7422,N_3819,N_2523);
nand U7423 (N_7423,N_2090,N_2300);
nand U7424 (N_7424,N_437,N_2015);
nor U7425 (N_7425,N_2714,N_2857);
and U7426 (N_7426,N_2944,N_3901);
nor U7427 (N_7427,N_3687,N_3361);
and U7428 (N_7428,N_2846,N_2631);
nor U7429 (N_7429,N_890,N_2831);
nor U7430 (N_7430,N_3874,N_3940);
and U7431 (N_7431,N_1793,N_3057);
nand U7432 (N_7432,N_1558,N_303);
or U7433 (N_7433,N_1673,N_2160);
and U7434 (N_7434,N_1366,N_3235);
or U7435 (N_7435,N_3071,N_1396);
and U7436 (N_7436,N_500,N_1701);
nand U7437 (N_7437,N_306,N_2016);
nand U7438 (N_7438,N_37,N_1386);
xor U7439 (N_7439,N_3518,N_1494);
nor U7440 (N_7440,N_877,N_1715);
nor U7441 (N_7441,N_1827,N_3856);
and U7442 (N_7442,N_775,N_2582);
and U7443 (N_7443,N_1079,N_2164);
nor U7444 (N_7444,N_1676,N_899);
and U7445 (N_7445,N_3797,N_2829);
and U7446 (N_7446,N_1601,N_1853);
and U7447 (N_7447,N_2049,N_128);
and U7448 (N_7448,N_3874,N_2301);
nor U7449 (N_7449,N_1433,N_324);
nor U7450 (N_7450,N_2848,N_482);
or U7451 (N_7451,N_3200,N_129);
nor U7452 (N_7452,N_1078,N_1745);
or U7453 (N_7453,N_751,N_3987);
nand U7454 (N_7454,N_1863,N_2688);
nor U7455 (N_7455,N_3340,N_3741);
xor U7456 (N_7456,N_1258,N_3345);
nand U7457 (N_7457,N_3481,N_1188);
nor U7458 (N_7458,N_3140,N_1779);
nand U7459 (N_7459,N_457,N_2871);
and U7460 (N_7460,N_1683,N_1645);
xor U7461 (N_7461,N_2677,N_1265);
nor U7462 (N_7462,N_1086,N_433);
xor U7463 (N_7463,N_1313,N_2797);
nor U7464 (N_7464,N_1787,N_1843);
xnor U7465 (N_7465,N_1951,N_3813);
nor U7466 (N_7466,N_2328,N_3650);
xor U7467 (N_7467,N_1468,N_3663);
nor U7468 (N_7468,N_1474,N_2609);
and U7469 (N_7469,N_3524,N_2526);
xor U7470 (N_7470,N_642,N_467);
and U7471 (N_7471,N_1392,N_3279);
nand U7472 (N_7472,N_1257,N_379);
nor U7473 (N_7473,N_1363,N_1685);
xor U7474 (N_7474,N_3831,N_6);
or U7475 (N_7475,N_2020,N_1206);
or U7476 (N_7476,N_1529,N_1377);
and U7477 (N_7477,N_2364,N_2794);
and U7478 (N_7478,N_1895,N_1675);
and U7479 (N_7479,N_3627,N_1049);
or U7480 (N_7480,N_3595,N_1480);
xor U7481 (N_7481,N_1172,N_2053);
or U7482 (N_7482,N_540,N_2821);
xnor U7483 (N_7483,N_2342,N_730);
or U7484 (N_7484,N_1547,N_506);
nand U7485 (N_7485,N_725,N_1887);
or U7486 (N_7486,N_3234,N_147);
xnor U7487 (N_7487,N_1536,N_3517);
and U7488 (N_7488,N_2565,N_3747);
nand U7489 (N_7489,N_2370,N_1674);
nor U7490 (N_7490,N_3824,N_1363);
or U7491 (N_7491,N_2859,N_1554);
xor U7492 (N_7492,N_1202,N_248);
and U7493 (N_7493,N_454,N_1908);
xnor U7494 (N_7494,N_3793,N_3288);
or U7495 (N_7495,N_3247,N_2337);
nor U7496 (N_7496,N_1976,N_264);
nor U7497 (N_7497,N_1018,N_2651);
or U7498 (N_7498,N_2882,N_372);
nand U7499 (N_7499,N_83,N_1302);
nand U7500 (N_7500,N_2556,N_753);
xor U7501 (N_7501,N_556,N_1098);
nor U7502 (N_7502,N_1180,N_593);
nand U7503 (N_7503,N_1415,N_1769);
nor U7504 (N_7504,N_2861,N_1054);
xnor U7505 (N_7505,N_1283,N_2355);
or U7506 (N_7506,N_744,N_1171);
xnor U7507 (N_7507,N_256,N_3707);
nor U7508 (N_7508,N_643,N_3733);
nand U7509 (N_7509,N_1970,N_3757);
nand U7510 (N_7510,N_2210,N_519);
xor U7511 (N_7511,N_560,N_3082);
nand U7512 (N_7512,N_276,N_1171);
nand U7513 (N_7513,N_1616,N_3761);
nand U7514 (N_7514,N_1064,N_3680);
nor U7515 (N_7515,N_3537,N_1404);
nor U7516 (N_7516,N_3511,N_2779);
and U7517 (N_7517,N_558,N_81);
nor U7518 (N_7518,N_898,N_1575);
and U7519 (N_7519,N_3373,N_2545);
xor U7520 (N_7520,N_2699,N_2419);
xnor U7521 (N_7521,N_2945,N_2345);
and U7522 (N_7522,N_2556,N_2476);
nor U7523 (N_7523,N_574,N_100);
xnor U7524 (N_7524,N_198,N_2621);
nor U7525 (N_7525,N_3390,N_3992);
nor U7526 (N_7526,N_2018,N_3824);
and U7527 (N_7527,N_3485,N_293);
or U7528 (N_7528,N_2827,N_1569);
nand U7529 (N_7529,N_1053,N_3176);
nand U7530 (N_7530,N_1262,N_3029);
and U7531 (N_7531,N_291,N_959);
nor U7532 (N_7532,N_2874,N_3898);
nor U7533 (N_7533,N_542,N_1516);
nand U7534 (N_7534,N_848,N_714);
nor U7535 (N_7535,N_2297,N_3615);
and U7536 (N_7536,N_450,N_3725);
or U7537 (N_7537,N_846,N_2067);
and U7538 (N_7538,N_1521,N_2652);
and U7539 (N_7539,N_1979,N_1500);
or U7540 (N_7540,N_1984,N_214);
and U7541 (N_7541,N_2541,N_1584);
nor U7542 (N_7542,N_479,N_929);
or U7543 (N_7543,N_1766,N_1025);
and U7544 (N_7544,N_526,N_3697);
and U7545 (N_7545,N_1670,N_884);
nor U7546 (N_7546,N_2293,N_423);
xnor U7547 (N_7547,N_332,N_1345);
or U7548 (N_7548,N_3506,N_2933);
and U7549 (N_7549,N_1006,N_3547);
and U7550 (N_7550,N_818,N_3270);
nor U7551 (N_7551,N_643,N_890);
xor U7552 (N_7552,N_1908,N_3567);
and U7553 (N_7553,N_1868,N_2455);
nor U7554 (N_7554,N_1703,N_1241);
nand U7555 (N_7555,N_1495,N_2265);
xor U7556 (N_7556,N_666,N_330);
xor U7557 (N_7557,N_3969,N_619);
or U7558 (N_7558,N_3342,N_1653);
and U7559 (N_7559,N_3185,N_1047);
xor U7560 (N_7560,N_2431,N_3669);
and U7561 (N_7561,N_355,N_1656);
nor U7562 (N_7562,N_352,N_3375);
and U7563 (N_7563,N_2534,N_2002);
xor U7564 (N_7564,N_181,N_1058);
xor U7565 (N_7565,N_2669,N_2150);
nor U7566 (N_7566,N_1479,N_1952);
xnor U7567 (N_7567,N_2010,N_2603);
and U7568 (N_7568,N_598,N_1632);
xor U7569 (N_7569,N_2453,N_91);
or U7570 (N_7570,N_142,N_3975);
and U7571 (N_7571,N_282,N_3476);
and U7572 (N_7572,N_858,N_2284);
xor U7573 (N_7573,N_3382,N_1803);
nor U7574 (N_7574,N_330,N_2748);
or U7575 (N_7575,N_2053,N_1833);
and U7576 (N_7576,N_841,N_3226);
nand U7577 (N_7577,N_859,N_1881);
or U7578 (N_7578,N_910,N_3646);
xnor U7579 (N_7579,N_2926,N_2325);
nor U7580 (N_7580,N_1257,N_1768);
or U7581 (N_7581,N_1312,N_2771);
xnor U7582 (N_7582,N_538,N_3355);
nand U7583 (N_7583,N_3731,N_1631);
xor U7584 (N_7584,N_2796,N_3640);
nor U7585 (N_7585,N_2094,N_2913);
and U7586 (N_7586,N_646,N_2723);
xor U7587 (N_7587,N_3748,N_3786);
and U7588 (N_7588,N_3677,N_1535);
xnor U7589 (N_7589,N_1958,N_2774);
or U7590 (N_7590,N_571,N_1685);
or U7591 (N_7591,N_1851,N_3994);
xnor U7592 (N_7592,N_241,N_591);
xnor U7593 (N_7593,N_3251,N_674);
or U7594 (N_7594,N_671,N_1802);
nor U7595 (N_7595,N_1397,N_3497);
nand U7596 (N_7596,N_786,N_2223);
nand U7597 (N_7597,N_3595,N_2434);
nor U7598 (N_7598,N_2220,N_2370);
and U7599 (N_7599,N_1052,N_15);
xnor U7600 (N_7600,N_3555,N_2288);
nor U7601 (N_7601,N_2008,N_2588);
nand U7602 (N_7602,N_2902,N_901);
xor U7603 (N_7603,N_1098,N_549);
xnor U7604 (N_7604,N_459,N_1245);
and U7605 (N_7605,N_3922,N_1141);
or U7606 (N_7606,N_2788,N_1505);
or U7607 (N_7607,N_1119,N_1717);
xnor U7608 (N_7608,N_489,N_446);
xor U7609 (N_7609,N_2877,N_1398);
and U7610 (N_7610,N_1382,N_1495);
nand U7611 (N_7611,N_2251,N_1124);
or U7612 (N_7612,N_1843,N_1581);
xor U7613 (N_7613,N_3948,N_2949);
nand U7614 (N_7614,N_184,N_2649);
nor U7615 (N_7615,N_2862,N_2116);
xnor U7616 (N_7616,N_975,N_2069);
and U7617 (N_7617,N_1930,N_2985);
or U7618 (N_7618,N_2142,N_74);
nor U7619 (N_7619,N_2782,N_3618);
and U7620 (N_7620,N_2265,N_1139);
or U7621 (N_7621,N_1948,N_2440);
or U7622 (N_7622,N_2862,N_2700);
xor U7623 (N_7623,N_2312,N_3485);
nor U7624 (N_7624,N_2379,N_648);
or U7625 (N_7625,N_1418,N_2511);
xnor U7626 (N_7626,N_3266,N_3949);
and U7627 (N_7627,N_1450,N_3603);
xnor U7628 (N_7628,N_3718,N_1704);
nor U7629 (N_7629,N_3505,N_3969);
nor U7630 (N_7630,N_2289,N_2887);
nor U7631 (N_7631,N_2592,N_2799);
or U7632 (N_7632,N_2747,N_3263);
xor U7633 (N_7633,N_2308,N_1130);
and U7634 (N_7634,N_891,N_1812);
and U7635 (N_7635,N_3709,N_1739);
nand U7636 (N_7636,N_1050,N_2598);
xnor U7637 (N_7637,N_1733,N_1444);
and U7638 (N_7638,N_2102,N_475);
and U7639 (N_7639,N_1403,N_2708);
xnor U7640 (N_7640,N_1082,N_2305);
nand U7641 (N_7641,N_2054,N_1848);
and U7642 (N_7642,N_3128,N_3466);
or U7643 (N_7643,N_3261,N_2216);
xor U7644 (N_7644,N_69,N_2619);
and U7645 (N_7645,N_1969,N_677);
and U7646 (N_7646,N_1522,N_1724);
or U7647 (N_7647,N_2303,N_2109);
nand U7648 (N_7648,N_874,N_3748);
nand U7649 (N_7649,N_2169,N_2638);
xor U7650 (N_7650,N_2396,N_1573);
and U7651 (N_7651,N_87,N_2584);
nand U7652 (N_7652,N_1639,N_3529);
and U7653 (N_7653,N_2270,N_374);
or U7654 (N_7654,N_1019,N_1934);
nand U7655 (N_7655,N_2504,N_730);
or U7656 (N_7656,N_37,N_3813);
and U7657 (N_7657,N_1614,N_2430);
nand U7658 (N_7658,N_3356,N_163);
nor U7659 (N_7659,N_2942,N_3380);
nand U7660 (N_7660,N_1516,N_2740);
and U7661 (N_7661,N_1364,N_1974);
nand U7662 (N_7662,N_658,N_2266);
and U7663 (N_7663,N_2859,N_3850);
nand U7664 (N_7664,N_636,N_1507);
and U7665 (N_7665,N_2098,N_2510);
and U7666 (N_7666,N_527,N_3229);
nor U7667 (N_7667,N_259,N_548);
nor U7668 (N_7668,N_722,N_2924);
nand U7669 (N_7669,N_1853,N_3693);
xnor U7670 (N_7670,N_595,N_741);
xnor U7671 (N_7671,N_796,N_713);
xnor U7672 (N_7672,N_3515,N_382);
and U7673 (N_7673,N_2218,N_1261);
xor U7674 (N_7674,N_3110,N_3775);
nand U7675 (N_7675,N_3524,N_1983);
or U7676 (N_7676,N_1848,N_566);
nor U7677 (N_7677,N_2061,N_2218);
and U7678 (N_7678,N_925,N_603);
nor U7679 (N_7679,N_2395,N_409);
or U7680 (N_7680,N_498,N_855);
nand U7681 (N_7681,N_1851,N_217);
nor U7682 (N_7682,N_3766,N_2293);
and U7683 (N_7683,N_1008,N_976);
or U7684 (N_7684,N_2716,N_1429);
nand U7685 (N_7685,N_2928,N_1860);
and U7686 (N_7686,N_980,N_1266);
or U7687 (N_7687,N_3448,N_26);
xnor U7688 (N_7688,N_1339,N_1445);
or U7689 (N_7689,N_2446,N_1023);
nand U7690 (N_7690,N_1911,N_699);
or U7691 (N_7691,N_755,N_2828);
xnor U7692 (N_7692,N_370,N_2552);
xnor U7693 (N_7693,N_319,N_1465);
xnor U7694 (N_7694,N_1149,N_3719);
or U7695 (N_7695,N_3053,N_3042);
or U7696 (N_7696,N_1267,N_1082);
xnor U7697 (N_7697,N_1675,N_3655);
nor U7698 (N_7698,N_808,N_2963);
xor U7699 (N_7699,N_932,N_2384);
or U7700 (N_7700,N_154,N_3616);
or U7701 (N_7701,N_3849,N_2598);
or U7702 (N_7702,N_737,N_732);
nor U7703 (N_7703,N_1344,N_2237);
nand U7704 (N_7704,N_2406,N_1371);
xor U7705 (N_7705,N_869,N_2069);
or U7706 (N_7706,N_3907,N_2245);
nand U7707 (N_7707,N_716,N_241);
xnor U7708 (N_7708,N_2649,N_3318);
nor U7709 (N_7709,N_1146,N_755);
nor U7710 (N_7710,N_2197,N_583);
xor U7711 (N_7711,N_2034,N_224);
or U7712 (N_7712,N_2098,N_1328);
nand U7713 (N_7713,N_259,N_2871);
nor U7714 (N_7714,N_1635,N_3728);
xor U7715 (N_7715,N_920,N_2906);
nand U7716 (N_7716,N_3979,N_3438);
or U7717 (N_7717,N_3936,N_328);
xor U7718 (N_7718,N_672,N_2279);
xor U7719 (N_7719,N_3798,N_19);
and U7720 (N_7720,N_3466,N_2991);
and U7721 (N_7721,N_3363,N_691);
and U7722 (N_7722,N_3966,N_929);
nor U7723 (N_7723,N_3080,N_474);
nand U7724 (N_7724,N_2694,N_1355);
nor U7725 (N_7725,N_590,N_2449);
nor U7726 (N_7726,N_2732,N_3131);
xnor U7727 (N_7727,N_1988,N_2933);
nand U7728 (N_7728,N_3524,N_229);
or U7729 (N_7729,N_1094,N_3143);
and U7730 (N_7730,N_1469,N_1428);
nor U7731 (N_7731,N_2304,N_2441);
nor U7732 (N_7732,N_1286,N_1302);
xor U7733 (N_7733,N_1089,N_1568);
xnor U7734 (N_7734,N_535,N_1775);
and U7735 (N_7735,N_3382,N_2417);
or U7736 (N_7736,N_1301,N_405);
nor U7737 (N_7737,N_2414,N_1030);
nor U7738 (N_7738,N_3828,N_3318);
nor U7739 (N_7739,N_2741,N_2981);
nor U7740 (N_7740,N_3834,N_2516);
nand U7741 (N_7741,N_3611,N_618);
xor U7742 (N_7742,N_585,N_3461);
xor U7743 (N_7743,N_357,N_2701);
or U7744 (N_7744,N_103,N_2733);
nor U7745 (N_7745,N_433,N_2226);
and U7746 (N_7746,N_492,N_2198);
xor U7747 (N_7747,N_2883,N_472);
or U7748 (N_7748,N_2875,N_752);
or U7749 (N_7749,N_1371,N_3928);
and U7750 (N_7750,N_1467,N_3145);
xnor U7751 (N_7751,N_782,N_2847);
and U7752 (N_7752,N_1288,N_2351);
nor U7753 (N_7753,N_1352,N_2388);
xor U7754 (N_7754,N_3035,N_1513);
xnor U7755 (N_7755,N_2095,N_3682);
nand U7756 (N_7756,N_1681,N_1225);
and U7757 (N_7757,N_2436,N_3201);
and U7758 (N_7758,N_1959,N_449);
nand U7759 (N_7759,N_303,N_2803);
or U7760 (N_7760,N_2598,N_1116);
xor U7761 (N_7761,N_3637,N_937);
xor U7762 (N_7762,N_1021,N_1557);
and U7763 (N_7763,N_775,N_1420);
nor U7764 (N_7764,N_1328,N_3628);
or U7765 (N_7765,N_276,N_2322);
nor U7766 (N_7766,N_3073,N_2846);
xnor U7767 (N_7767,N_2293,N_2409);
or U7768 (N_7768,N_1210,N_2500);
nand U7769 (N_7769,N_2475,N_3987);
nor U7770 (N_7770,N_2428,N_1908);
or U7771 (N_7771,N_585,N_814);
nand U7772 (N_7772,N_3552,N_1351);
xnor U7773 (N_7773,N_249,N_3287);
or U7774 (N_7774,N_259,N_3011);
or U7775 (N_7775,N_28,N_3395);
nand U7776 (N_7776,N_3579,N_1084);
or U7777 (N_7777,N_2185,N_2340);
nand U7778 (N_7778,N_349,N_2655);
nor U7779 (N_7779,N_590,N_3137);
nor U7780 (N_7780,N_2436,N_2555);
nand U7781 (N_7781,N_933,N_1113);
and U7782 (N_7782,N_2916,N_1951);
nand U7783 (N_7783,N_2732,N_1451);
nor U7784 (N_7784,N_3166,N_1658);
nand U7785 (N_7785,N_1639,N_2889);
nand U7786 (N_7786,N_1183,N_2626);
xor U7787 (N_7787,N_2087,N_999);
and U7788 (N_7788,N_1767,N_3843);
or U7789 (N_7789,N_3960,N_758);
and U7790 (N_7790,N_3246,N_1355);
nand U7791 (N_7791,N_3088,N_587);
and U7792 (N_7792,N_1518,N_3728);
and U7793 (N_7793,N_3989,N_2260);
or U7794 (N_7794,N_1432,N_2807);
nor U7795 (N_7795,N_1043,N_683);
or U7796 (N_7796,N_1397,N_2537);
xor U7797 (N_7797,N_195,N_1673);
and U7798 (N_7798,N_1330,N_2142);
xnor U7799 (N_7799,N_3347,N_3605);
nand U7800 (N_7800,N_2468,N_2938);
or U7801 (N_7801,N_1844,N_2578);
and U7802 (N_7802,N_983,N_1344);
xnor U7803 (N_7803,N_391,N_295);
nand U7804 (N_7804,N_473,N_1400);
nor U7805 (N_7805,N_3866,N_873);
or U7806 (N_7806,N_3133,N_3770);
xnor U7807 (N_7807,N_2646,N_2139);
and U7808 (N_7808,N_3595,N_2307);
and U7809 (N_7809,N_2473,N_1131);
nor U7810 (N_7810,N_1750,N_1017);
nand U7811 (N_7811,N_1415,N_3131);
and U7812 (N_7812,N_280,N_421);
or U7813 (N_7813,N_2700,N_2618);
nand U7814 (N_7814,N_876,N_3374);
nand U7815 (N_7815,N_1236,N_2896);
nor U7816 (N_7816,N_862,N_2535);
or U7817 (N_7817,N_156,N_726);
nand U7818 (N_7818,N_1611,N_3320);
nor U7819 (N_7819,N_1880,N_3817);
and U7820 (N_7820,N_1656,N_951);
or U7821 (N_7821,N_940,N_2084);
or U7822 (N_7822,N_1271,N_3169);
or U7823 (N_7823,N_2660,N_2534);
xnor U7824 (N_7824,N_487,N_2035);
or U7825 (N_7825,N_1091,N_401);
xor U7826 (N_7826,N_1149,N_3124);
xor U7827 (N_7827,N_3195,N_2640);
or U7828 (N_7828,N_3352,N_1590);
xnor U7829 (N_7829,N_3041,N_2992);
and U7830 (N_7830,N_2809,N_1673);
and U7831 (N_7831,N_697,N_2362);
or U7832 (N_7832,N_1747,N_3226);
nand U7833 (N_7833,N_3894,N_2595);
nor U7834 (N_7834,N_568,N_3915);
xor U7835 (N_7835,N_1986,N_3669);
nor U7836 (N_7836,N_3579,N_1090);
nor U7837 (N_7837,N_1276,N_3048);
or U7838 (N_7838,N_3913,N_3463);
xor U7839 (N_7839,N_3183,N_51);
and U7840 (N_7840,N_1110,N_3295);
and U7841 (N_7841,N_1086,N_2036);
and U7842 (N_7842,N_3009,N_2173);
or U7843 (N_7843,N_3204,N_2602);
xor U7844 (N_7844,N_554,N_1800);
nor U7845 (N_7845,N_3452,N_3479);
nand U7846 (N_7846,N_2452,N_2323);
or U7847 (N_7847,N_1199,N_2322);
and U7848 (N_7848,N_3639,N_3511);
nor U7849 (N_7849,N_642,N_3209);
or U7850 (N_7850,N_3324,N_49);
and U7851 (N_7851,N_3074,N_1471);
or U7852 (N_7852,N_43,N_1964);
or U7853 (N_7853,N_3075,N_202);
or U7854 (N_7854,N_1706,N_665);
and U7855 (N_7855,N_860,N_2911);
and U7856 (N_7856,N_1487,N_2592);
and U7857 (N_7857,N_1708,N_1527);
xnor U7858 (N_7858,N_3104,N_2909);
nor U7859 (N_7859,N_3274,N_2854);
and U7860 (N_7860,N_43,N_2479);
or U7861 (N_7861,N_1665,N_2260);
or U7862 (N_7862,N_679,N_977);
nand U7863 (N_7863,N_243,N_1464);
nor U7864 (N_7864,N_456,N_3314);
xor U7865 (N_7865,N_2894,N_2867);
nor U7866 (N_7866,N_1712,N_379);
nand U7867 (N_7867,N_26,N_3504);
nor U7868 (N_7868,N_690,N_364);
or U7869 (N_7869,N_3409,N_1387);
and U7870 (N_7870,N_2041,N_3461);
and U7871 (N_7871,N_2342,N_1879);
nor U7872 (N_7872,N_3272,N_3907);
xor U7873 (N_7873,N_311,N_2072);
xnor U7874 (N_7874,N_3246,N_1070);
nor U7875 (N_7875,N_1371,N_498);
nand U7876 (N_7876,N_2777,N_3998);
nor U7877 (N_7877,N_3315,N_1226);
nand U7878 (N_7878,N_3841,N_3323);
or U7879 (N_7879,N_1885,N_813);
nor U7880 (N_7880,N_1089,N_2859);
nor U7881 (N_7881,N_2721,N_437);
xnor U7882 (N_7882,N_2681,N_1430);
nand U7883 (N_7883,N_149,N_889);
xor U7884 (N_7884,N_1587,N_729);
or U7885 (N_7885,N_1847,N_941);
or U7886 (N_7886,N_836,N_801);
and U7887 (N_7887,N_2824,N_1610);
and U7888 (N_7888,N_280,N_3897);
xnor U7889 (N_7889,N_544,N_1134);
nor U7890 (N_7890,N_3284,N_3449);
or U7891 (N_7891,N_535,N_2293);
nand U7892 (N_7892,N_2599,N_2023);
nor U7893 (N_7893,N_1401,N_2367);
nor U7894 (N_7894,N_1187,N_1779);
nor U7895 (N_7895,N_533,N_3216);
or U7896 (N_7896,N_3349,N_3158);
or U7897 (N_7897,N_968,N_2303);
and U7898 (N_7898,N_1352,N_2610);
nand U7899 (N_7899,N_724,N_1993);
and U7900 (N_7900,N_998,N_3208);
xnor U7901 (N_7901,N_3770,N_2731);
or U7902 (N_7902,N_2489,N_2705);
xor U7903 (N_7903,N_490,N_1902);
or U7904 (N_7904,N_1115,N_2471);
nand U7905 (N_7905,N_728,N_308);
and U7906 (N_7906,N_3972,N_376);
nand U7907 (N_7907,N_559,N_3716);
and U7908 (N_7908,N_3679,N_1075);
xnor U7909 (N_7909,N_1554,N_2569);
nand U7910 (N_7910,N_1082,N_2447);
nand U7911 (N_7911,N_594,N_3928);
or U7912 (N_7912,N_1015,N_1990);
nand U7913 (N_7913,N_1141,N_2685);
nand U7914 (N_7914,N_337,N_802);
xnor U7915 (N_7915,N_2174,N_2843);
or U7916 (N_7916,N_1707,N_255);
nor U7917 (N_7917,N_1295,N_1349);
and U7918 (N_7918,N_110,N_3550);
nor U7919 (N_7919,N_2081,N_511);
and U7920 (N_7920,N_2762,N_2027);
xor U7921 (N_7921,N_660,N_434);
nor U7922 (N_7922,N_2546,N_3317);
nand U7923 (N_7923,N_2679,N_3169);
nor U7924 (N_7924,N_1314,N_910);
xor U7925 (N_7925,N_3178,N_391);
or U7926 (N_7926,N_2801,N_1885);
nor U7927 (N_7927,N_3316,N_666);
nand U7928 (N_7928,N_2696,N_3297);
and U7929 (N_7929,N_3828,N_2919);
and U7930 (N_7930,N_2881,N_650);
xnor U7931 (N_7931,N_7,N_32);
or U7932 (N_7932,N_1985,N_2300);
nor U7933 (N_7933,N_2096,N_1595);
nand U7934 (N_7934,N_3155,N_236);
or U7935 (N_7935,N_3344,N_1815);
nand U7936 (N_7936,N_1314,N_168);
xnor U7937 (N_7937,N_637,N_2168);
or U7938 (N_7938,N_802,N_445);
or U7939 (N_7939,N_1580,N_2319);
xnor U7940 (N_7940,N_62,N_420);
or U7941 (N_7941,N_630,N_3729);
nand U7942 (N_7942,N_347,N_3395);
and U7943 (N_7943,N_2497,N_2769);
nand U7944 (N_7944,N_417,N_2095);
or U7945 (N_7945,N_2175,N_255);
and U7946 (N_7946,N_187,N_2293);
xor U7947 (N_7947,N_3014,N_252);
nand U7948 (N_7948,N_21,N_1317);
nand U7949 (N_7949,N_444,N_1756);
nand U7950 (N_7950,N_44,N_3198);
nor U7951 (N_7951,N_906,N_1535);
or U7952 (N_7952,N_1998,N_1057);
nor U7953 (N_7953,N_1465,N_1794);
or U7954 (N_7954,N_900,N_2240);
nor U7955 (N_7955,N_3744,N_1968);
and U7956 (N_7956,N_1610,N_3530);
xnor U7957 (N_7957,N_3919,N_2421);
nand U7958 (N_7958,N_2870,N_1682);
xor U7959 (N_7959,N_3876,N_2951);
or U7960 (N_7960,N_621,N_2850);
xor U7961 (N_7961,N_3877,N_1416);
nand U7962 (N_7962,N_2696,N_2521);
or U7963 (N_7963,N_675,N_1146);
nor U7964 (N_7964,N_3001,N_3752);
nor U7965 (N_7965,N_3402,N_2167);
nor U7966 (N_7966,N_1534,N_1518);
and U7967 (N_7967,N_498,N_2672);
or U7968 (N_7968,N_1819,N_3037);
nand U7969 (N_7969,N_1413,N_2344);
and U7970 (N_7970,N_2035,N_483);
nor U7971 (N_7971,N_161,N_579);
and U7972 (N_7972,N_3885,N_90);
or U7973 (N_7973,N_2284,N_3054);
nor U7974 (N_7974,N_1428,N_1319);
nand U7975 (N_7975,N_3974,N_2816);
nor U7976 (N_7976,N_851,N_3096);
nor U7977 (N_7977,N_3643,N_1944);
or U7978 (N_7978,N_1315,N_1154);
nand U7979 (N_7979,N_3666,N_2569);
and U7980 (N_7980,N_3871,N_2718);
or U7981 (N_7981,N_814,N_3557);
or U7982 (N_7982,N_3587,N_1482);
nand U7983 (N_7983,N_3371,N_3818);
or U7984 (N_7984,N_2317,N_2419);
xnor U7985 (N_7985,N_213,N_3791);
nand U7986 (N_7986,N_322,N_1179);
nand U7987 (N_7987,N_1977,N_580);
xor U7988 (N_7988,N_2899,N_1429);
nor U7989 (N_7989,N_2286,N_844);
or U7990 (N_7990,N_2206,N_592);
nor U7991 (N_7991,N_2436,N_398);
nor U7992 (N_7992,N_2997,N_1856);
nor U7993 (N_7993,N_690,N_1189);
xnor U7994 (N_7994,N_1400,N_1208);
and U7995 (N_7995,N_2689,N_17);
or U7996 (N_7996,N_122,N_810);
nor U7997 (N_7997,N_375,N_1769);
nand U7998 (N_7998,N_1103,N_718);
nand U7999 (N_7999,N_1139,N_1954);
or U8000 (N_8000,N_6013,N_7080);
nand U8001 (N_8001,N_7775,N_4356);
or U8002 (N_8002,N_4502,N_6156);
or U8003 (N_8003,N_4376,N_4565);
nand U8004 (N_8004,N_5681,N_7674);
nand U8005 (N_8005,N_5424,N_5583);
xnor U8006 (N_8006,N_7028,N_6250);
nor U8007 (N_8007,N_7008,N_6432);
nor U8008 (N_8008,N_6678,N_5794);
xor U8009 (N_8009,N_5767,N_6100);
nand U8010 (N_8010,N_5477,N_6442);
and U8011 (N_8011,N_6585,N_5735);
and U8012 (N_8012,N_5361,N_5574);
or U8013 (N_8013,N_6344,N_6727);
or U8014 (N_8014,N_4115,N_6473);
nor U8015 (N_8015,N_4351,N_5578);
xnor U8016 (N_8016,N_7742,N_5799);
or U8017 (N_8017,N_7535,N_7689);
nor U8018 (N_8018,N_7533,N_7122);
xor U8019 (N_8019,N_4674,N_5149);
xor U8020 (N_8020,N_4558,N_6812);
or U8021 (N_8021,N_4863,N_4839);
nand U8022 (N_8022,N_7400,N_5093);
nor U8023 (N_8023,N_7646,N_4668);
and U8024 (N_8024,N_5970,N_6909);
nand U8025 (N_8025,N_4231,N_6019);
xor U8026 (N_8026,N_5363,N_6178);
xor U8027 (N_8027,N_4452,N_6641);
nor U8028 (N_8028,N_6653,N_4746);
and U8029 (N_8029,N_4461,N_4190);
nor U8030 (N_8030,N_5816,N_5516);
or U8031 (N_8031,N_6881,N_6425);
nor U8032 (N_8032,N_7229,N_6203);
or U8033 (N_8033,N_4197,N_6785);
xnor U8034 (N_8034,N_7837,N_7587);
nor U8035 (N_8035,N_7138,N_6333);
or U8036 (N_8036,N_7499,N_6628);
xor U8037 (N_8037,N_6599,N_4894);
and U8038 (N_8038,N_5994,N_4369);
nand U8039 (N_8039,N_4793,N_5371);
xor U8040 (N_8040,N_5848,N_5895);
xor U8041 (N_8041,N_6774,N_6088);
nand U8042 (N_8042,N_7590,N_7137);
or U8043 (N_8043,N_4174,N_7757);
or U8044 (N_8044,N_5060,N_6128);
xnor U8045 (N_8045,N_4717,N_5193);
or U8046 (N_8046,N_7176,N_7382);
and U8047 (N_8047,N_5148,N_7253);
nor U8048 (N_8048,N_7687,N_4968);
nand U8049 (N_8049,N_6371,N_5854);
or U8050 (N_8050,N_5438,N_6457);
and U8051 (N_8051,N_5980,N_6916);
or U8052 (N_8052,N_6948,N_4990);
or U8053 (N_8053,N_5039,N_7723);
and U8054 (N_8054,N_6900,N_6361);
and U8055 (N_8055,N_6502,N_4037);
and U8056 (N_8056,N_6142,N_7476);
nand U8057 (N_8057,N_7384,N_4886);
xor U8058 (N_8058,N_4074,N_5935);
and U8059 (N_8059,N_5270,N_4339);
nand U8060 (N_8060,N_6720,N_4344);
or U8061 (N_8061,N_6841,N_5126);
nor U8062 (N_8062,N_5421,N_5308);
or U8063 (N_8063,N_7230,N_6665);
nand U8064 (N_8064,N_7112,N_7811);
or U8065 (N_8065,N_7691,N_6805);
and U8066 (N_8066,N_6219,N_6509);
xor U8067 (N_8067,N_6077,N_7490);
nand U8068 (N_8068,N_6747,N_5910);
nand U8069 (N_8069,N_4959,N_5731);
nand U8070 (N_8070,N_5032,N_6707);
nor U8071 (N_8071,N_5224,N_5598);
xnor U8072 (N_8072,N_7399,N_7795);
xnor U8073 (N_8073,N_7185,N_5792);
xor U8074 (N_8074,N_6410,N_6086);
or U8075 (N_8075,N_6043,N_5857);
xor U8076 (N_8076,N_7900,N_7810);
nor U8077 (N_8077,N_6436,N_6122);
nor U8078 (N_8078,N_5919,N_7644);
and U8079 (N_8079,N_6474,N_7487);
nand U8080 (N_8080,N_5601,N_5163);
or U8081 (N_8081,N_7680,N_5011);
nand U8082 (N_8082,N_4872,N_4666);
nand U8083 (N_8083,N_6381,N_7827);
and U8084 (N_8084,N_7525,N_6397);
or U8085 (N_8085,N_6376,N_4543);
or U8086 (N_8086,N_5461,N_7302);
xnor U8087 (N_8087,N_4146,N_4789);
nor U8088 (N_8088,N_4679,N_6946);
nor U8089 (N_8089,N_7505,N_6701);
xnor U8090 (N_8090,N_7061,N_6065);
nor U8091 (N_8091,N_4070,N_4229);
xnor U8092 (N_8092,N_4887,N_7193);
nor U8093 (N_8093,N_7958,N_5652);
nand U8094 (N_8094,N_4470,N_5441);
nor U8095 (N_8095,N_6238,N_7031);
xnor U8096 (N_8096,N_4498,N_6637);
nand U8097 (N_8097,N_7312,N_7600);
xnor U8098 (N_8098,N_5947,N_6406);
xor U8099 (N_8099,N_6192,N_7840);
nor U8100 (N_8100,N_6363,N_6117);
and U8101 (N_8101,N_4049,N_7026);
xnor U8102 (N_8102,N_5991,N_7602);
or U8103 (N_8103,N_5688,N_7359);
nor U8104 (N_8104,N_7580,N_5013);
nand U8105 (N_8105,N_7783,N_5633);
nand U8106 (N_8106,N_4606,N_4203);
and U8107 (N_8107,N_7162,N_7376);
and U8108 (N_8108,N_6405,N_7098);
and U8109 (N_8109,N_4172,N_6233);
xor U8110 (N_8110,N_6882,N_5266);
xnor U8111 (N_8111,N_5973,N_7632);
or U8112 (N_8112,N_7362,N_5218);
nor U8113 (N_8113,N_4426,N_6109);
nand U8114 (N_8114,N_7497,N_7621);
nand U8115 (N_8115,N_4370,N_6115);
nand U8116 (N_8116,N_5143,N_7921);
and U8117 (N_8117,N_5339,N_4248);
nor U8118 (N_8118,N_4308,N_5462);
or U8119 (N_8119,N_4664,N_5705);
nand U8120 (N_8120,N_5996,N_7336);
and U8121 (N_8121,N_7892,N_6658);
xor U8122 (N_8122,N_6736,N_4034);
and U8123 (N_8123,N_6022,N_6412);
nand U8124 (N_8124,N_4327,N_6280);
xnor U8125 (N_8125,N_5096,N_4041);
nor U8126 (N_8126,N_4384,N_7240);
or U8127 (N_8127,N_4734,N_7576);
or U8128 (N_8128,N_5064,N_6551);
and U8129 (N_8129,N_4023,N_4224);
nand U8130 (N_8130,N_5599,N_4320);
xnor U8131 (N_8131,N_7287,N_6932);
nand U8132 (N_8132,N_5426,N_4216);
nand U8133 (N_8133,N_4552,N_5117);
and U8134 (N_8134,N_6159,N_4812);
and U8135 (N_8135,N_7044,N_7539);
or U8136 (N_8136,N_6708,N_6012);
xor U8137 (N_8137,N_6721,N_7804);
and U8138 (N_8138,N_7430,N_7984);
and U8139 (N_8139,N_5539,N_4529);
and U8140 (N_8140,N_5999,N_7421);
nor U8141 (N_8141,N_6617,N_6190);
nand U8142 (N_8142,N_4360,N_6400);
nor U8143 (N_8143,N_5328,N_7702);
nand U8144 (N_8144,N_6781,N_6503);
or U8145 (N_8145,N_7348,N_4992);
and U8146 (N_8146,N_7378,N_6582);
nand U8147 (N_8147,N_7995,N_6464);
nor U8148 (N_8148,N_6673,N_5326);
and U8149 (N_8149,N_7924,N_4016);
nand U8150 (N_8150,N_5928,N_7994);
xor U8151 (N_8151,N_7938,N_7531);
nor U8152 (N_8152,N_6271,N_7196);
xor U8153 (N_8153,N_6015,N_7506);
or U8154 (N_8154,N_6155,N_4391);
and U8155 (N_8155,N_4245,N_5151);
or U8156 (N_8156,N_5275,N_5906);
xnor U8157 (N_8157,N_4177,N_5787);
nor U8158 (N_8158,N_6912,N_7781);
nand U8159 (N_8159,N_4333,N_5136);
nor U8160 (N_8160,N_6667,N_6931);
nor U8161 (N_8161,N_7522,N_5563);
or U8162 (N_8162,N_7290,N_5536);
nor U8163 (N_8163,N_5548,N_5391);
or U8164 (N_8164,N_5923,N_6231);
and U8165 (N_8165,N_6698,N_6668);
or U8166 (N_8166,N_4388,N_4732);
xnor U8167 (N_8167,N_5432,N_5034);
xor U8168 (N_8168,N_5868,N_4846);
nor U8169 (N_8169,N_4154,N_7953);
nor U8170 (N_8170,N_4591,N_6516);
nand U8171 (N_8171,N_7179,N_7456);
xor U8172 (N_8172,N_5142,N_6028);
nand U8173 (N_8173,N_7609,N_6073);
xor U8174 (N_8174,N_6869,N_6740);
and U8175 (N_8175,N_6259,N_7990);
xnor U8176 (N_8176,N_6385,N_5079);
and U8177 (N_8177,N_5028,N_6794);
xnor U8178 (N_8178,N_5227,N_7555);
xor U8179 (N_8179,N_7592,N_6205);
xor U8180 (N_8180,N_5492,N_6248);
nand U8181 (N_8181,N_7625,N_6601);
nand U8182 (N_8182,N_4214,N_4392);
xnor U8183 (N_8183,N_6640,N_6839);
or U8184 (N_8184,N_7013,N_5805);
and U8185 (N_8185,N_4755,N_4842);
and U8186 (N_8186,N_4701,N_5761);
and U8187 (N_8187,N_6246,N_5707);
xnor U8188 (N_8188,N_6697,N_5097);
nor U8189 (N_8189,N_5430,N_6369);
and U8190 (N_8190,N_5900,N_7259);
xnor U8191 (N_8191,N_4085,N_4551);
and U8192 (N_8192,N_4962,N_4466);
nor U8193 (N_8193,N_6004,N_4390);
nor U8194 (N_8194,N_7737,N_7982);
and U8195 (N_8195,N_6103,N_4366);
xor U8196 (N_8196,N_4646,N_4513);
nand U8197 (N_8197,N_4143,N_4865);
nor U8198 (N_8198,N_4446,N_6296);
xnor U8199 (N_8199,N_7326,N_7599);
or U8200 (N_8200,N_4970,N_5833);
and U8201 (N_8201,N_5873,N_7090);
nor U8202 (N_8202,N_4189,N_7719);
nor U8203 (N_8203,N_5116,N_7853);
nor U8204 (N_8204,N_7330,N_7432);
and U8205 (N_8205,N_6394,N_5304);
xnor U8206 (N_8206,N_6198,N_6561);
nor U8207 (N_8207,N_6168,N_5934);
nor U8208 (N_8208,N_6165,N_5544);
nand U8209 (N_8209,N_6976,N_7672);
or U8210 (N_8210,N_6763,N_7416);
and U8211 (N_8211,N_7860,N_5258);
nor U8212 (N_8212,N_7077,N_6594);
nand U8213 (N_8213,N_7886,N_6853);
nand U8214 (N_8214,N_6398,N_4110);
nand U8215 (N_8215,N_4548,N_6251);
xor U8216 (N_8216,N_6196,N_6386);
nor U8217 (N_8217,N_4159,N_4258);
xor U8218 (N_8218,N_4422,N_5954);
or U8219 (N_8219,N_6789,N_6281);
or U8220 (N_8220,N_4613,N_7466);
xor U8221 (N_8221,N_7793,N_4620);
nor U8222 (N_8222,N_7046,N_5734);
and U8223 (N_8223,N_4563,N_5770);
nor U8224 (N_8224,N_5090,N_4557);
nand U8225 (N_8225,N_7393,N_5621);
or U8226 (N_8226,N_4864,N_7548);
and U8227 (N_8227,N_6924,N_4240);
and U8228 (N_8228,N_4500,N_5213);
and U8229 (N_8229,N_4331,N_5405);
xor U8230 (N_8230,N_5993,N_4757);
or U8231 (N_8231,N_5831,N_6269);
xor U8232 (N_8232,N_4136,N_4031);
nand U8233 (N_8233,N_4379,N_7120);
nand U8234 (N_8234,N_4028,N_4241);
or U8235 (N_8235,N_6552,N_7504);
and U8236 (N_8236,N_7911,N_4766);
xnor U8237 (N_8237,N_7299,N_5184);
or U8238 (N_8238,N_6389,N_7079);
nor U8239 (N_8239,N_6954,N_7649);
nor U8240 (N_8240,N_7203,N_7927);
nor U8241 (N_8241,N_6663,N_4805);
or U8242 (N_8242,N_6603,N_6989);
and U8243 (N_8243,N_7469,N_4553);
xnor U8244 (N_8244,N_7666,N_4862);
and U8245 (N_8245,N_4799,N_5709);
nand U8246 (N_8246,N_6266,N_6120);
or U8247 (N_8247,N_4753,N_6961);
xnor U8248 (N_8248,N_6471,N_7475);
nor U8249 (N_8249,N_7059,N_4788);
or U8250 (N_8250,N_6630,N_5909);
xnor U8251 (N_8251,N_6513,N_6298);
nand U8252 (N_8252,N_6137,N_4627);
nor U8253 (N_8253,N_4103,N_4907);
or U8254 (N_8254,N_4955,N_6826);
nand U8255 (N_8255,N_6753,N_5966);
nor U8256 (N_8256,N_4087,N_6475);
nor U8257 (N_8257,N_6141,N_6230);
nor U8258 (N_8258,N_5692,N_4768);
nor U8259 (N_8259,N_5262,N_7463);
nor U8260 (N_8260,N_4210,N_7086);
or U8261 (N_8261,N_6879,N_6815);
nand U8262 (N_8262,N_4910,N_5879);
and U8263 (N_8263,N_4160,N_4610);
nor U8264 (N_8264,N_5535,N_7233);
xor U8265 (N_8265,N_4050,N_6758);
and U8266 (N_8266,N_5716,N_7100);
xor U8267 (N_8267,N_4129,N_7991);
and U8268 (N_8268,N_4100,N_5500);
nor U8269 (N_8269,N_7248,N_5656);
or U8270 (N_8270,N_4305,N_7740);
nand U8271 (N_8271,N_4938,N_5866);
nand U8272 (N_8272,N_4642,N_4059);
and U8273 (N_8273,N_4365,N_5051);
or U8274 (N_8274,N_6408,N_5239);
or U8275 (N_8275,N_6477,N_5964);
nand U8276 (N_8276,N_6144,N_5431);
xnor U8277 (N_8277,N_7738,N_4600);
nor U8278 (N_8278,N_4228,N_5031);
nor U8279 (N_8279,N_7244,N_6240);
xnor U8280 (N_8280,N_7882,N_7569);
or U8281 (N_8281,N_6487,N_6000);
or U8282 (N_8282,N_7198,N_4246);
or U8283 (N_8283,N_7934,N_5941);
xnor U8284 (N_8284,N_5518,N_4082);
xor U8285 (N_8285,N_6490,N_5261);
nor U8286 (N_8286,N_5596,N_6472);
nand U8287 (N_8287,N_6716,N_4684);
nand U8288 (N_8288,N_7055,N_4782);
nor U8289 (N_8289,N_7500,N_7067);
or U8290 (N_8290,N_7191,N_6510);
xor U8291 (N_8291,N_5501,N_4425);
nor U8292 (N_8292,N_7849,N_7231);
nand U8293 (N_8293,N_7129,N_7772);
nor U8294 (N_8294,N_5622,N_5394);
nor U8295 (N_8295,N_6466,N_4357);
and U8296 (N_8296,N_6959,N_4086);
nor U8297 (N_8297,N_5472,N_6878);
nor U8298 (N_8298,N_5524,N_4225);
or U8299 (N_8299,N_6044,N_5072);
nor U8300 (N_8300,N_4213,N_4437);
or U8301 (N_8301,N_6360,N_7307);
nand U8302 (N_8302,N_6664,N_6666);
nor U8303 (N_8303,N_6831,N_6237);
nand U8304 (N_8304,N_7647,N_4381);
nand U8305 (N_8305,N_4338,N_7972);
nand U8306 (N_8306,N_5154,N_4877);
nor U8307 (N_8307,N_6549,N_5454);
or U8308 (N_8308,N_7023,N_7441);
or U8309 (N_8309,N_4284,N_4869);
or U8310 (N_8310,N_7655,N_7216);
nor U8311 (N_8311,N_7693,N_7431);
nor U8312 (N_8312,N_7623,N_6352);
and U8313 (N_8313,N_7489,N_4407);
xnor U8314 (N_8314,N_7217,N_7513);
nand U8315 (N_8315,N_5134,N_4754);
nor U8316 (N_8316,N_6782,N_6530);
or U8317 (N_8317,N_5532,N_4608);
nand U8318 (N_8318,N_7752,N_5696);
nor U8319 (N_8319,N_5094,N_7797);
and U8320 (N_8320,N_5479,N_7607);
or U8321 (N_8321,N_4647,N_7438);
nand U8322 (N_8322,N_5570,N_7219);
xor U8323 (N_8323,N_6094,N_5939);
or U8324 (N_8324,N_7683,N_5365);
or U8325 (N_8325,N_6732,N_7803);
nand U8326 (N_8326,N_6330,N_6966);
and U8327 (N_8327,N_6301,N_5292);
xnor U8328 (N_8328,N_6645,N_5020);
xor U8329 (N_8329,N_5826,N_4525);
nand U8330 (N_8330,N_4816,N_5503);
and U8331 (N_8331,N_7186,N_4409);
xor U8332 (N_8332,N_6072,N_6903);
nor U8333 (N_8333,N_6705,N_4455);
nand U8334 (N_8334,N_7496,N_6814);
xor U8335 (N_8335,N_7769,N_5331);
or U8336 (N_8336,N_7825,N_4705);
nand U8337 (N_8337,N_6342,N_7610);
and U8338 (N_8338,N_6462,N_7532);
xor U8339 (N_8339,N_4111,N_4510);
xor U8340 (N_8340,N_6304,N_4811);
xor U8341 (N_8341,N_6880,N_6748);
nor U8342 (N_8342,N_6730,N_7885);
nand U8343 (N_8343,N_4429,N_7405);
nor U8344 (N_8344,N_5357,N_4982);
nor U8345 (N_8345,N_6070,N_5319);
or U8346 (N_8346,N_4221,N_6082);
xnor U8347 (N_8347,N_7733,N_6684);
or U8348 (N_8348,N_5443,N_5623);
and U8349 (N_8349,N_5089,N_7971);
or U8350 (N_8350,N_4697,N_6213);
or U8351 (N_8351,N_6169,N_6654);
nand U8352 (N_8352,N_7454,N_7916);
nor U8353 (N_8353,N_6195,N_4855);
or U8354 (N_8354,N_5087,N_6152);
or U8355 (N_8355,N_7778,N_6855);
nor U8356 (N_8356,N_4215,N_7690);
nand U8357 (N_8357,N_5335,N_5765);
xor U8358 (N_8358,N_6706,N_4514);
and U8359 (N_8359,N_7043,N_7942);
or U8360 (N_8360,N_7969,N_7817);
or U8361 (N_8361,N_6001,N_6309);
nand U8362 (N_8362,N_7836,N_5006);
xnor U8363 (N_8363,N_4279,N_6693);
nor U8364 (N_8364,N_4184,N_7643);
and U8365 (N_8365,N_6107,N_5471);
nand U8366 (N_8366,N_7746,N_4472);
nor U8367 (N_8367,N_5124,N_4921);
nand U8368 (N_8368,N_7225,N_7669);
nor U8369 (N_8369,N_6559,N_6484);
nand U8370 (N_8370,N_7876,N_6067);
nor U8371 (N_8371,N_5297,N_4899);
nand U8372 (N_8372,N_5250,N_4499);
nand U8373 (N_8373,N_7692,N_7327);
nor U8374 (N_8374,N_5358,N_4084);
xnor U8375 (N_8375,N_7104,N_5442);
nor U8376 (N_8376,N_7977,N_4092);
or U8377 (N_8377,N_6064,N_5068);
nor U8378 (N_8378,N_5246,N_7285);
xor U8379 (N_8379,N_4948,N_4904);
or U8380 (N_8380,N_7367,N_4763);
nor U8381 (N_8381,N_7020,N_4343);
nand U8382 (N_8382,N_5323,N_7874);
and U8383 (N_8383,N_4930,N_5661);
nand U8384 (N_8384,N_6886,N_5607);
or U8385 (N_8385,N_7767,N_6536);
and U8386 (N_8386,N_5670,N_4698);
nand U8387 (N_8387,N_4290,N_6501);
nand U8388 (N_8388,N_7980,N_7549);
nand U8389 (N_8389,N_4896,N_4532);
xor U8390 (N_8390,N_4434,N_6616);
or U8391 (N_8391,N_5377,N_6867);
xnor U8392 (N_8392,N_7851,N_6134);
nand U8393 (N_8393,N_7320,N_7800);
xor U8394 (N_8394,N_5401,N_4881);
xor U8395 (N_8395,N_4412,N_5385);
or U8396 (N_8396,N_4478,N_6085);
xor U8397 (N_8397,N_6467,N_4737);
nand U8398 (N_8398,N_6054,N_4432);
or U8399 (N_8399,N_6834,N_4994);
and U8400 (N_8400,N_5674,N_4878);
nand U8401 (N_8401,N_6925,N_7965);
and U8402 (N_8402,N_7736,N_7920);
xor U8403 (N_8403,N_5197,N_4544);
xnor U8404 (N_8404,N_4520,N_5478);
nand U8405 (N_8405,N_7758,N_7677);
or U8406 (N_8406,N_4194,N_7741);
or U8407 (N_8407,N_5368,N_4021);
or U8408 (N_8408,N_7612,N_5330);
or U8409 (N_8409,N_7147,N_5602);
nand U8410 (N_8410,N_5738,N_4662);
xor U8411 (N_8411,N_5965,N_4670);
or U8412 (N_8412,N_6816,N_5043);
or U8413 (N_8413,N_6928,N_6050);
or U8414 (N_8414,N_6556,N_4716);
nand U8415 (N_8415,N_4958,N_7952);
or U8416 (N_8416,N_4671,N_7234);
nand U8417 (N_8417,N_6988,N_7829);
nor U8418 (N_8418,N_4682,N_7585);
xor U8419 (N_8419,N_7973,N_4122);
nor U8420 (N_8420,N_6648,N_6135);
nand U8421 (N_8421,N_7355,N_5008);
or U8422 (N_8422,N_5714,N_5210);
and U8423 (N_8423,N_7863,N_6350);
xor U8424 (N_8424,N_4774,N_6861);
or U8425 (N_8425,N_4919,N_6367);
and U8426 (N_8426,N_5538,N_4927);
xor U8427 (N_8427,N_5676,N_6613);
nor U8428 (N_8428,N_4814,N_5931);
nand U8429 (N_8429,N_4348,N_7163);
nor U8430 (N_8430,N_6186,N_6624);
or U8431 (N_8431,N_6311,N_4148);
or U8432 (N_8432,N_5740,N_4905);
nand U8433 (N_8433,N_6393,N_7485);
nand U8434 (N_8434,N_5299,N_5915);
and U8435 (N_8435,N_4306,N_7664);
or U8436 (N_8436,N_5437,N_5384);
nor U8437 (N_8437,N_4775,N_5231);
nand U8438 (N_8438,N_4299,N_7651);
nand U8439 (N_8439,N_7053,N_4566);
nor U8440 (N_8440,N_4696,N_4139);
xnor U8441 (N_8441,N_5286,N_7016);
nand U8442 (N_8442,N_4106,N_7967);
nor U8443 (N_8443,N_6187,N_6023);
or U8444 (N_8444,N_5850,N_4556);
nand U8445 (N_8445,N_5170,N_7173);
and U8446 (N_8446,N_7880,N_5105);
nor U8447 (N_8447,N_4272,N_7679);
xor U8448 (N_8448,N_6353,N_6116);
xnor U8449 (N_8449,N_5427,N_5809);
and U8450 (N_8450,N_4202,N_6850);
nor U8451 (N_8451,N_6985,N_7512);
nand U8452 (N_8452,N_7192,N_7319);
or U8453 (N_8453,N_6683,N_6149);
nor U8454 (N_8454,N_6798,N_5214);
and U8455 (N_8455,N_6323,N_7184);
or U8456 (N_8456,N_4710,N_4024);
or U8457 (N_8457,N_7996,N_4007);
nand U8458 (N_8458,N_7865,N_5916);
xnor U8459 (N_8459,N_7905,N_4756);
or U8460 (N_8460,N_7389,N_7261);
xor U8461 (N_8461,N_4777,N_6680);
and U8462 (N_8462,N_5315,N_7774);
xnor U8463 (N_8463,N_4477,N_6537);
or U8464 (N_8464,N_7611,N_6769);
nand U8465 (N_8465,N_7989,N_6583);
or U8466 (N_8466,N_6292,N_5369);
nand U8467 (N_8467,N_7088,N_6262);
xnor U8468 (N_8468,N_5665,N_6750);
nand U8469 (N_8469,N_5891,N_7986);
xor U8470 (N_8470,N_7349,N_7749);
or U8471 (N_8471,N_7235,N_5751);
nand U8472 (N_8472,N_6136,N_5413);
xor U8473 (N_8473,N_7369,N_4095);
nor U8474 (N_8474,N_6810,N_7819);
xnor U8475 (N_8475,N_6066,N_7280);
or U8476 (N_8476,N_6914,N_4616);
nor U8477 (N_8477,N_4868,N_6779);
or U8478 (N_8478,N_5156,N_7418);
xor U8479 (N_8479,N_6532,N_7826);
nor U8480 (N_8480,N_6570,N_4932);
nor U8481 (N_8481,N_5648,N_5957);
xor U8482 (N_8482,N_7335,N_5415);
nand U8483 (N_8483,N_4694,N_6236);
nor U8484 (N_8484,N_5905,N_6153);
nand U8485 (N_8485,N_7332,N_7727);
and U8486 (N_8486,N_6799,N_7919);
or U8487 (N_8487,N_5509,N_7822);
and U8488 (N_8488,N_7241,N_7070);
or U8489 (N_8489,N_6453,N_5230);
and U8490 (N_8490,N_6539,N_5823);
nand U8491 (N_8491,N_4634,N_5961);
and U8492 (N_8492,N_4019,N_4821);
or U8493 (N_8493,N_6962,N_5309);
nand U8494 (N_8494,N_6545,N_5643);
nand U8495 (N_8495,N_6542,N_4656);
and U8496 (N_8496,N_5215,N_5445);
xnor U8497 (N_8497,N_5158,N_4198);
or U8498 (N_8498,N_7002,N_7410);
nor U8499 (N_8499,N_7642,N_7142);
xnor U8500 (N_8500,N_6145,N_4526);
xor U8501 (N_8501,N_5194,N_6669);
and U8502 (N_8502,N_4644,N_6254);
and U8503 (N_8503,N_5217,N_4924);
nor U8504 (N_8504,N_5933,N_7954);
nand U8505 (N_8505,N_5813,N_5414);
xnor U8506 (N_8506,N_4715,N_5929);
nor U8507 (N_8507,N_4005,N_5708);
and U8508 (N_8508,N_4964,N_4860);
xor U8509 (N_8509,N_4233,N_7862);
xor U8510 (N_8510,N_7588,N_7582);
xor U8511 (N_8511,N_6214,N_7218);
nor U8512 (N_8512,N_7484,N_7855);
or U8513 (N_8513,N_6918,N_4292);
and U8514 (N_8514,N_5924,N_4713);
and U8515 (N_8515,N_7745,N_5896);
nor U8516 (N_8516,N_7178,N_6862);
xor U8517 (N_8517,N_6897,N_4971);
nor U8518 (N_8518,N_5693,N_7204);
or U8519 (N_8519,N_6306,N_4829);
and U8520 (N_8520,N_7118,N_4624);
and U8521 (N_8521,N_4700,N_4131);
and U8522 (N_8522,N_7426,N_4107);
nand U8523 (N_8523,N_7988,N_6228);
nor U8524 (N_8524,N_5666,N_7258);
nand U8525 (N_8525,N_6679,N_4998);
nor U8526 (N_8526,N_7558,N_4564);
xor U8527 (N_8527,N_6600,N_5510);
nor U8528 (N_8528,N_7465,N_6795);
or U8529 (N_8529,N_4988,N_6982);
xor U8530 (N_8530,N_6026,N_6923);
or U8531 (N_8531,N_4650,N_7530);
xnor U8532 (N_8532,N_4588,N_6671);
xnor U8533 (N_8533,N_7269,N_4375);
and U8534 (N_8534,N_6081,N_7150);
nor U8535 (N_8535,N_5593,N_7902);
nand U8536 (N_8536,N_4469,N_6366);
nor U8537 (N_8537,N_4673,N_5914);
or U8538 (N_8538,N_7943,N_6483);
nor U8539 (N_8539,N_6661,N_4012);
or U8540 (N_8540,N_4685,N_6772);
and U8541 (N_8541,N_5412,N_7102);
nor U8542 (N_8542,N_4844,N_5689);
xor U8543 (N_8543,N_5101,N_4206);
or U8544 (N_8544,N_4722,N_5281);
nor U8545 (N_8545,N_4524,N_5710);
and U8546 (N_8546,N_4419,N_5284);
and U8547 (N_8547,N_4781,N_4835);
nor U8548 (N_8548,N_7848,N_5983);
nand U8549 (N_8549,N_7333,N_4677);
xnor U8550 (N_8550,N_6902,N_4505);
xor U8551 (N_8551,N_5836,N_5182);
xnor U8552 (N_8552,N_4386,N_5779);
xor U8553 (N_8553,N_6258,N_6964);
and U8554 (N_8554,N_7939,N_5141);
xnor U8555 (N_8555,N_6399,N_4871);
xnor U8556 (N_8556,N_7591,N_5588);
and U8557 (N_8557,N_7409,N_7615);
and U8558 (N_8558,N_5066,N_5575);
or U8559 (N_8559,N_4751,N_4180);
nor U8560 (N_8560,N_5366,N_7560);
nor U8561 (N_8561,N_5395,N_5969);
nand U8562 (N_8562,N_7445,N_5122);
nand U8563 (N_8563,N_7334,N_4771);
nand U8564 (N_8564,N_4792,N_5968);
nand U8565 (N_8565,N_6182,N_7676);
xor U8566 (N_8566,N_6199,N_4504);
and U8567 (N_8567,N_4665,N_5133);
nand U8568 (N_8568,N_5789,N_6127);
nand U8569 (N_8569,N_5650,N_5393);
or U8570 (N_8570,N_7520,N_4410);
nand U8571 (N_8571,N_4117,N_5436);
or U8572 (N_8572,N_7540,N_7557);
and U8573 (N_8573,N_6992,N_7718);
and U8574 (N_8574,N_6579,N_6950);
and U8575 (N_8575,N_4571,N_5756);
nand U8576 (N_8576,N_7833,N_6334);
or U8577 (N_8577,N_6283,N_7681);
nand U8578 (N_8578,N_7675,N_5336);
nor U8579 (N_8579,N_5383,N_7869);
or U8580 (N_8580,N_4185,N_4081);
nand U8581 (N_8581,N_4261,N_7375);
nor U8582 (N_8582,N_7776,N_5550);
and U8583 (N_8583,N_7437,N_5581);
nand U8584 (N_8584,N_5591,N_6560);
nor U8585 (N_8585,N_4067,N_6692);
xnor U8586 (N_8586,N_6092,N_5940);
nor U8587 (N_8587,N_7271,N_4803);
or U8588 (N_8588,N_7415,N_7717);
xnor U8589 (N_8589,N_5922,N_5360);
xor U8590 (N_8590,N_5819,N_6179);
and U8591 (N_8591,N_6619,N_5654);
or U8592 (N_8592,N_6002,N_4270);
and U8593 (N_8593,N_7117,N_5706);
nand U8594 (N_8594,N_6700,N_6215);
and U8595 (N_8595,N_6965,N_5296);
nand U8596 (N_8596,N_4873,N_6325);
xor U8597 (N_8597,N_6687,N_7239);
xor U8598 (N_8598,N_7823,N_4761);
nand U8599 (N_8599,N_6365,N_7834);
nand U8600 (N_8600,N_7893,N_6053);
xnor U8601 (N_8601,N_7018,N_4801);
xor U8602 (N_8602,N_7183,N_5342);
or U8603 (N_8603,N_7207,N_6076);
nand U8604 (N_8604,N_7981,N_4127);
or U8605 (N_8605,N_7597,N_4946);
xor U8606 (N_8606,N_5428,N_5174);
xnor U8607 (N_8607,N_4638,N_7725);
and U8608 (N_8608,N_6390,N_6910);
xor U8609 (N_8609,N_7347,N_5561);
and U8610 (N_8610,N_7806,N_6118);
or U8611 (N_8611,N_4884,N_4738);
or U8612 (N_8612,N_4066,N_4156);
or U8613 (N_8613,N_7564,N_5103);
and U8614 (N_8614,N_7297,N_7483);
xnor U8615 (N_8615,N_5624,N_6990);
and U8616 (N_8616,N_7627,N_4555);
nor U8617 (N_8617,N_6388,N_5860);
nand U8618 (N_8618,N_4486,N_6150);
nand U8619 (N_8619,N_4337,N_6057);
xor U8620 (N_8620,N_5264,N_7455);
xor U8621 (N_8621,N_5465,N_6191);
and U8622 (N_8622,N_7524,N_5632);
nor U8623 (N_8623,N_7386,N_7126);
and U8624 (N_8624,N_5159,N_6413);
nor U8625 (N_8625,N_7284,N_5178);
xor U8626 (N_8626,N_4997,N_4415);
nor U8627 (N_8627,N_6685,N_5029);
or U8628 (N_8628,N_4920,N_5012);
nor U8629 (N_8629,N_4212,N_6775);
and U8630 (N_8630,N_5743,N_5568);
and U8631 (N_8631,N_5499,N_5844);
xnor U8632 (N_8632,N_7937,N_6362);
nand U8633 (N_8633,N_6544,N_4138);
or U8634 (N_8634,N_7908,N_5989);
xnor U8635 (N_8635,N_5855,N_5301);
or U8636 (N_8636,N_4441,N_4018);
nand U8637 (N_8637,N_7652,N_7784);
xor U8638 (N_8638,N_5541,N_5549);
nand U8639 (N_8639,N_5995,N_4731);
or U8640 (N_8640,N_7923,N_4026);
and U8641 (N_8641,N_4527,N_4603);
xor U8642 (N_8642,N_5475,N_7033);
or U8643 (N_8643,N_6029,N_6373);
or U8644 (N_8644,N_6039,N_6580);
and U8645 (N_8645,N_5605,N_5613);
and U8646 (N_8646,N_4022,N_5979);
nor U8647 (N_8647,N_6377,N_4928);
and U8648 (N_8648,N_4661,N_4612);
or U8649 (N_8649,N_7787,N_5338);
and U8650 (N_8650,N_6895,N_6096);
and U8651 (N_8651,N_4961,N_7537);
xnor U8652 (N_8652,N_7699,N_4263);
nand U8653 (N_8653,N_4124,N_4947);
nor U8654 (N_8654,N_4237,N_6686);
or U8655 (N_8655,N_7068,N_7831);
or U8656 (N_8656,N_7789,N_4631);
nand U8657 (N_8657,N_4838,N_4791);
xnor U8658 (N_8658,N_5768,N_6338);
nand U8659 (N_8659,N_5379,N_6726);
or U8660 (N_8660,N_6439,N_6804);
and U8661 (N_8661,N_6253,N_6303);
xor U8662 (N_8662,N_7364,N_5373);
nor U8663 (N_8663,N_6584,N_7371);
or U8664 (N_8664,N_6368,N_6524);
xor U8665 (N_8665,N_4414,N_5533);
nand U8666 (N_8666,N_7124,N_6297);
nand U8667 (N_8667,N_7313,N_4825);
and U8668 (N_8668,N_6102,N_4503);
or U8669 (N_8669,N_5899,N_7314);
xnor U8670 (N_8670,N_6776,N_4332);
nor U8671 (N_8671,N_7922,N_6217);
xor U8672 (N_8672,N_6171,N_5824);
xor U8673 (N_8673,N_5750,N_7756);
nor U8674 (N_8674,N_4675,N_7422);
or U8675 (N_8675,N_7073,N_4394);
nor U8676 (N_8676,N_6564,N_5634);
nor U8677 (N_8677,N_6905,N_7429);
or U8678 (N_8678,N_5378,N_4813);
or U8679 (N_8679,N_4836,N_7556);
or U8680 (N_8680,N_4040,N_5829);
or U8681 (N_8681,N_7148,N_4362);
nor U8682 (N_8682,N_5482,N_7205);
or U8683 (N_8683,N_5747,N_5080);
xor U8684 (N_8684,N_5259,N_4218);
nand U8685 (N_8685,N_6284,N_6223);
nor U8686 (N_8686,N_5663,N_7573);
xnor U8687 (N_8687,N_7309,N_6387);
and U8688 (N_8688,N_6971,N_6454);
and U8689 (N_8689,N_4377,N_7365);
or U8690 (N_8690,N_5901,N_7562);
or U8691 (N_8691,N_5179,N_7606);
nand U8692 (N_8692,N_4017,N_4531);
xnor U8693 (N_8693,N_4222,N_4048);
nor U8694 (N_8694,N_5419,N_5452);
xnor U8695 (N_8695,N_5755,N_7698);
xor U8696 (N_8696,N_4062,N_6497);
and U8697 (N_8697,N_5067,N_7477);
and U8698 (N_8698,N_4423,N_7346);
or U8699 (N_8699,N_5589,N_6565);
and U8700 (N_8700,N_7385,N_7589);
nand U8701 (N_8701,N_4770,N_4265);
nor U8702 (N_8702,N_7001,N_6746);
or U8703 (N_8703,N_5382,N_6557);
nand U8704 (N_8704,N_7766,N_7747);
xnor U8705 (N_8705,N_5701,N_5444);
nor U8706 (N_8706,N_4010,N_4800);
and U8707 (N_8707,N_5838,N_6021);
nand U8708 (N_8708,N_5463,N_5932);
or U8709 (N_8709,N_7639,N_6904);
nand U8710 (N_8710,N_7278,N_7167);
xnor U8711 (N_8711,N_4659,N_6337);
or U8712 (N_8712,N_6974,N_7554);
nor U8713 (N_8713,N_7479,N_4155);
and U8714 (N_8714,N_6095,N_7166);
nor U8715 (N_8715,N_4678,N_5480);
and U8716 (N_8716,N_5843,N_4223);
nand U8717 (N_8717,N_6936,N_6224);
nor U8718 (N_8718,N_6162,N_4511);
nand U8719 (N_8719,N_7604,N_5307);
xnor U8720 (N_8720,N_7563,N_4105);
nor U8721 (N_8721,N_7807,N_4083);
xor U8722 (N_8722,N_4236,N_5257);
and U8723 (N_8723,N_6384,N_6622);
nand U8724 (N_8724,N_6016,N_4064);
nor U8725 (N_8725,N_6773,N_7502);
and U8726 (N_8726,N_6744,N_5121);
or U8727 (N_8727,N_7957,N_4572);
nor U8728 (N_8728,N_5033,N_5736);
and U8729 (N_8729,N_6105,N_4942);
nand U8730 (N_8730,N_5712,N_7412);
nand U8731 (N_8731,N_7157,N_6293);
nand U8732 (N_8732,N_5289,N_7103);
nand U8733 (N_8733,N_6891,N_6518);
and U8734 (N_8734,N_5311,N_6525);
xor U8735 (N_8735,N_5410,N_5769);
and U8736 (N_8736,N_6575,N_7598);
nor U8737 (N_8737,N_6681,N_7060);
or U8738 (N_8738,N_4523,N_6434);
xnor U8739 (N_8739,N_5677,N_5820);
xnor U8740 (N_8740,N_5113,N_7041);
and U8741 (N_8741,N_5841,N_5249);
and U8742 (N_8742,N_7559,N_5085);
or U8743 (N_8743,N_5595,N_4030);
or U8744 (N_8744,N_7411,N_6119);
or U8745 (N_8745,N_6970,N_6754);
and U8746 (N_8746,N_5943,N_7846);
nand U8747 (N_8747,N_7131,N_6140);
xnor U8748 (N_8748,N_4304,N_5293);
or U8749 (N_8749,N_7021,N_4209);
and U8750 (N_8750,N_5290,N_5955);
or U8751 (N_8751,N_7898,N_4519);
nor U8752 (N_8752,N_6784,N_4458);
nor U8753 (N_8753,N_5571,N_6504);
and U8754 (N_8754,N_5181,N_6341);
nand U8755 (N_8755,N_6531,N_6963);
or U8756 (N_8756,N_7006,N_6113);
nand U8757 (N_8757,N_4164,N_5686);
nand U8758 (N_8758,N_4055,N_6468);
nor U8759 (N_8759,N_7267,N_4451);
or U8760 (N_8760,N_5885,N_4667);
or U8761 (N_8761,N_4618,N_4517);
and U8762 (N_8762,N_5356,N_5035);
or U8763 (N_8763,N_4396,N_6335);
and U8764 (N_8764,N_7744,N_6148);
or U8765 (N_8765,N_5070,N_6177);
and U8766 (N_8766,N_6351,N_6894);
nor U8767 (N_8767,N_6414,N_5175);
nand U8768 (N_8768,N_6090,N_6991);
xor U8769 (N_8769,N_7448,N_5084);
nand U8770 (N_8770,N_4883,N_4706);
nor U8771 (N_8771,N_5017,N_5327);
and U8772 (N_8772,N_6702,N_6567);
nand U8773 (N_8773,N_7237,N_5668);
and U8774 (N_8774,N_4244,N_6357);
nand U8775 (N_8775,N_5889,N_6218);
nor U8776 (N_8776,N_7622,N_6999);
nand U8777 (N_8777,N_6183,N_7584);
nor U8778 (N_8778,N_5271,N_4895);
and U8779 (N_8779,N_7380,N_4776);
nor U8780 (N_8780,N_7883,N_6056);
xnor U8781 (N_8781,N_4235,N_4687);
and U8782 (N_8782,N_7731,N_5616);
or U8783 (N_8783,N_7815,N_5135);
nand U8784 (N_8784,N_4060,N_4125);
nand U8785 (N_8785,N_6308,N_6901);
nand U8786 (N_8786,N_7879,N_7553);
xnor U8787 (N_8787,N_6543,N_4045);
xor U8788 (N_8788,N_6540,N_4691);
nor U8789 (N_8789,N_5411,N_7620);
xnor U8790 (N_8790,N_7425,N_7720);
or U8791 (N_8791,N_5449,N_7636);
or U8792 (N_8792,N_5375,N_6741);
and U8793 (N_8793,N_6193,N_5147);
and U8794 (N_8794,N_4590,N_6097);
nand U8795 (N_8795,N_5053,N_6864);
nand U8796 (N_8796,N_7397,N_6174);
or U8797 (N_8797,N_5222,N_4851);
xnor U8798 (N_8798,N_5321,N_4619);
xnor U8799 (N_8799,N_6521,N_4853);
nor U8800 (N_8800,N_7914,N_4042);
or U8801 (N_8801,N_4984,N_7136);
xor U8802 (N_8802,N_5531,N_5263);
and U8803 (N_8803,N_4493,N_6327);
or U8804 (N_8804,N_7019,N_7743);
xor U8805 (N_8805,N_7839,N_7528);
nor U8806 (N_8806,N_4617,N_4914);
xnor U8807 (N_8807,N_7895,N_5274);
xnor U8808 (N_8808,N_4602,N_4573);
nor U8809 (N_8809,N_7273,N_5766);
and U8810 (N_8810,N_5195,N_5741);
nand U8811 (N_8811,N_4848,N_7661);
nor U8812 (N_8812,N_5007,N_7750);
or U8813 (N_8813,N_4876,N_5639);
nor U8814 (N_8814,N_5146,N_5399);
nor U8815 (N_8815,N_5638,N_7368);
xor U8816 (N_8816,N_4354,N_6857);
nand U8817 (N_8817,N_5021,N_7974);
nor U8818 (N_8818,N_7700,N_5100);
nand U8819 (N_8819,N_7036,N_5076);
nand U8820 (N_8820,N_4718,N_6586);
nor U8821 (N_8821,N_6951,N_4020);
or U8822 (N_8822,N_7404,N_6045);
xnor U8823 (N_8823,N_4039,N_6647);
or U8824 (N_8824,N_7838,N_5849);
or U8825 (N_8825,N_5106,N_7575);
nor U8826 (N_8826,N_6079,N_7867);
nand U8827 (N_8827,N_4965,N_5423);
xor U8828 (N_8828,N_5243,N_5256);
nand U8829 (N_8829,N_7710,N_4438);
nand U8830 (N_8830,N_5726,N_5904);
nor U8831 (N_8831,N_4622,N_7571);
nand U8832 (N_8832,N_7075,N_6060);
or U8833 (N_8833,N_4903,N_7480);
or U8834 (N_8834,N_5959,N_4481);
or U8835 (N_8835,N_6427,N_5952);
or U8836 (N_8836,N_5690,N_5306);
nor U8837 (N_8837,N_7351,N_5355);
xnor U8838 (N_8838,N_5206,N_7398);
or U8839 (N_8839,N_7667,N_4297);
or U8840 (N_8840,N_7978,N_6611);
and U8841 (N_8841,N_5265,N_4275);
xnor U8842 (N_8842,N_7703,N_7250);
nor U8843 (N_8843,N_5487,N_6597);
and U8844 (N_8844,N_5520,N_5782);
nand U8845 (N_8845,N_5123,N_7311);
xor U8846 (N_8846,N_5211,N_6438);
and U8847 (N_8847,N_6317,N_6278);
and U8848 (N_8848,N_5703,N_6263);
xor U8849 (N_8849,N_5821,N_4480);
nand U8850 (N_8850,N_6005,N_5667);
nor U8851 (N_8851,N_6709,N_7308);
or U8852 (N_8852,N_5642,N_7788);
nand U8853 (N_8853,N_6069,N_6494);
and U8854 (N_8854,N_7451,N_6621);
nand U8855 (N_8855,N_4257,N_4643);
nand U8856 (N_8856,N_6885,N_7868);
nand U8857 (N_8857,N_5842,N_6260);
xnor U8858 (N_8858,N_4818,N_7493);
xor U8859 (N_8859,N_5114,N_6378);
or U8860 (N_8860,N_5902,N_4852);
xor U8861 (N_8861,N_4416,N_6167);
xor U8862 (N_8862,N_5715,N_6972);
nor U8863 (N_8863,N_5881,N_7444);
and U8864 (N_8864,N_7705,N_6703);
nand U8865 (N_8865,N_6605,N_7095);
or U8866 (N_8866,N_5763,N_6485);
or U8867 (N_8867,N_4326,N_4114);
xnor U8868 (N_8868,N_6455,N_6670);
xor U8869 (N_8869,N_4750,N_7780);
nand U8870 (N_8870,N_7948,N_7288);
and U8871 (N_8871,N_5276,N_6290);
nand U8872 (N_8872,N_6899,N_6286);
and U8873 (N_8873,N_6660,N_4826);
or U8874 (N_8874,N_6558,N_7453);
nand U8875 (N_8875,N_7040,N_7631);
nor U8876 (N_8876,N_7232,N_6949);
nor U8877 (N_8877,N_6755,N_4204);
and U8878 (N_8878,N_5204,N_5491);
or U8879 (N_8879,N_5176,N_7903);
xnor U8880 (N_8880,N_6819,N_4892);
or U8881 (N_8881,N_5802,N_7315);
and U8882 (N_8882,N_5111,N_5791);
or U8883 (N_8883,N_6157,N_5972);
and U8884 (N_8884,N_4798,N_7896);
nor U8885 (N_8885,N_4253,N_5662);
nor U8886 (N_8886,N_7577,N_4823);
nor U8887 (N_8887,N_4785,N_7545);
nor U8888 (N_8888,N_4002,N_7089);
xor U8889 (N_8889,N_5903,N_6633);
xor U8890 (N_8890,N_4157,N_7706);
nand U8891 (N_8891,N_5978,N_6061);
or U8892 (N_8892,N_7037,N_7189);
nor U8893 (N_8893,N_6522,N_4708);
nor U8894 (N_8894,N_5523,N_4276);
nand U8895 (N_8895,N_6749,N_4870);
nor U8896 (N_8896,N_4522,N_7732);
xnor U8897 (N_8897,N_6623,N_7728);
xor U8898 (N_8898,N_5644,N_4546);
xor U8899 (N_8899,N_4547,N_5683);
and U8900 (N_8900,N_5488,N_7403);
xnor U8901 (N_8901,N_7045,N_6034);
xor U8902 (N_8902,N_6921,N_5493);
and U8903 (N_8903,N_5212,N_5260);
xor U8904 (N_8904,N_7277,N_7813);
nor U8905 (N_8905,N_6917,N_4495);
and U8906 (N_8906,N_4681,N_7790);
or U8907 (N_8907,N_5671,N_7085);
xnor U8908 (N_8908,N_4382,N_4875);
nor U8909 (N_8909,N_6239,N_4733);
nand U8910 (N_8910,N_6934,N_6059);
nand U8911 (N_8911,N_7966,N_5847);
or U8912 (N_8912,N_5073,N_6541);
and U8913 (N_8913,N_7875,N_4772);
xnor U8914 (N_8914,N_5723,N_5003);
xnor U8915 (N_8915,N_6553,N_7983);
nor U8916 (N_8916,N_7711,N_4453);
nand U8917 (N_8917,N_5115,N_5753);
and U8918 (N_8918,N_7751,N_5387);
or U8919 (N_8919,N_7133,N_5956);
xnor U8920 (N_8920,N_6835,N_5807);
and U8921 (N_8921,N_6953,N_7645);
and U8922 (N_8922,N_5945,N_5131);
nand U8923 (N_8923,N_5853,N_5234);
or U8924 (N_8924,N_6578,N_7704);
xor U8925 (N_8925,N_7381,N_4936);
or U8926 (N_8926,N_6620,N_7999);
nor U8927 (N_8927,N_6715,N_6517);
nor U8928 (N_8928,N_7214,N_4424);
nor U8929 (N_8929,N_5912,N_4334);
nand U8930 (N_8930,N_5537,N_4294);
xor U8931 (N_8931,N_6515,N_6287);
nor U8932 (N_8932,N_7158,N_5880);
nand U8933 (N_8933,N_5872,N_7910);
nor U8934 (N_8934,N_5988,N_4358);
or U8935 (N_8935,N_4038,N_4161);
nand U8936 (N_8936,N_6602,N_5014);
xor U8937 (N_8937,N_6614,N_4636);
nand U8938 (N_8938,N_6573,N_6143);
nand U8939 (N_8939,N_6347,N_7304);
nand U8940 (N_8940,N_4170,N_7887);
and U8941 (N_8941,N_7613,N_7383);
xor U8942 (N_8942,N_6593,N_4385);
nor U8943 (N_8943,N_4345,N_7594);
xnor U8944 (N_8944,N_6958,N_5225);
and U8945 (N_8945,N_5882,N_5627);
and U8946 (N_8946,N_5288,N_5062);
or U8947 (N_8947,N_5229,N_7464);
nand U8948 (N_8948,N_6112,N_4723);
nand U8949 (N_8949,N_4145,N_6802);
and U8950 (N_8950,N_4251,N_6783);
xor U8951 (N_8951,N_7407,N_5645);
and U8952 (N_8952,N_5167,N_4703);
nor U8953 (N_8953,N_4787,N_6933);
nand U8954 (N_8954,N_7873,N_5127);
nor U8955 (N_8955,N_4922,N_7926);
or U8956 (N_8956,N_5396,N_7066);
xor U8957 (N_8957,N_5757,N_6828);
or U8958 (N_8958,N_4318,N_5888);
nor U8959 (N_8959,N_6104,N_7935);
nand U8960 (N_8960,N_7828,N_7961);
xnor U8961 (N_8961,N_7424,N_4653);
nand U8962 (N_8962,N_7321,N_7940);
or U8963 (N_8963,N_5777,N_5272);
nand U8964 (N_8964,N_5235,N_5529);
nor U8965 (N_8965,N_5316,N_4625);
nand U8966 (N_8966,N_6419,N_6383);
nand U8967 (N_8967,N_6766,N_5725);
xnor U8968 (N_8968,N_4595,N_7361);
nand U8969 (N_8969,N_4321,N_7678);
nand U8970 (N_8970,N_4112,N_5015);
xor U8971 (N_8971,N_7195,N_6121);
and U8972 (N_8972,N_4689,N_7442);
nand U8973 (N_8973,N_7701,N_6194);
nand U8974 (N_8974,N_5019,N_7032);
nand U8975 (N_8975,N_6007,N_6639);
nor U8976 (N_8976,N_4317,N_7296);
and U8977 (N_8977,N_5637,N_4536);
and U8978 (N_8978,N_7339,N_6520);
and U8979 (N_8979,N_4188,N_6185);
or U8980 (N_8980,N_6256,N_4854);
and U8981 (N_8981,N_7527,N_7199);
nand U8982 (N_8982,N_4448,N_6245);
xor U8983 (N_8983,N_6125,N_6722);
nand U8984 (N_8984,N_4578,N_7458);
xor U8985 (N_8985,N_4956,N_4699);
or U8986 (N_8986,N_4283,N_5579);
nand U8987 (N_8987,N_5470,N_5926);
or U8988 (N_8988,N_4604,N_5102);
or U8989 (N_8989,N_7439,N_7128);
nand U8990 (N_8990,N_5056,N_6089);
nor U8991 (N_8991,N_7292,N_5279);
or U8992 (N_8992,N_4226,N_5352);
and U8993 (N_8993,N_6396,N_4940);
xnor U8994 (N_8994,N_5987,N_6030);
nor U8995 (N_8995,N_6505,N_6382);
nand U8996 (N_8996,N_5440,N_6915);
nor U8997 (N_8997,N_7175,N_6295);
xor U8998 (N_8998,N_6969,N_6941);
and U8999 (N_8999,N_7069,N_5386);
nand U9000 (N_9000,N_4280,N_4058);
or U9001 (N_9001,N_7567,N_6823);
nand U9002 (N_9002,N_5893,N_7668);
nor U9003 (N_9003,N_4439,N_4073);
or U9004 (N_9004,N_4807,N_4802);
and U9005 (N_9005,N_6587,N_7156);
and U9006 (N_9006,N_4714,N_7256);
nor U9007 (N_9007,N_6735,N_7266);
nor U9008 (N_9008,N_7579,N_6318);
and U9009 (N_9009,N_5191,N_7394);
nor U9010 (N_9010,N_6032,N_6206);
xnor U9011 (N_9011,N_6011,N_7242);
xnor U9012 (N_9012,N_5082,N_4580);
and U9013 (N_9013,N_4035,N_6204);
nand U9014 (N_9014,N_7153,N_4660);
or U9015 (N_9015,N_4815,N_4693);
and U9016 (N_9016,N_5504,N_6737);
nand U9017 (N_9017,N_7058,N_7395);
or U9018 (N_9018,N_7516,N_5138);
and U9019 (N_9019,N_5490,N_6273);
nor U9020 (N_9020,N_7065,N_6796);
or U9021 (N_9021,N_4859,N_4747);
or U9022 (N_9022,N_5647,N_5077);
nand U9023 (N_9023,N_4219,N_4267);
nor U9024 (N_9024,N_5244,N_6025);
or U9025 (N_9025,N_4882,N_5758);
nand U9026 (N_9026,N_5057,N_4047);
nor U9027 (N_9027,N_7946,N_4786);
nand U9028 (N_9028,N_4487,N_5422);
and U9029 (N_9029,N_7494,N_6947);
or U9030 (N_9030,N_6590,N_5207);
nand U9031 (N_9031,N_4911,N_5425);
nor U9032 (N_9032,N_4142,N_4827);
xor U9033 (N_9033,N_6312,N_7707);
nor U9034 (N_9034,N_5099,N_6672);
nor U9035 (N_9035,N_4707,N_5233);
nand U9036 (N_9036,N_4593,N_5201);
nor U9037 (N_9037,N_6876,N_7402);
or U9038 (N_9038,N_4421,N_5930);
or U9039 (N_9039,N_4582,N_4061);
nor U9040 (N_9040,N_4232,N_7039);
nand U9041 (N_9041,N_7072,N_5208);
nand U9042 (N_9042,N_4688,N_7709);
nand U9043 (N_9043,N_5606,N_4954);
nor U9044 (N_9044,N_7255,N_7634);
and U9045 (N_9045,N_5389,N_4999);
nand U9046 (N_9046,N_4075,N_7928);
nand U9047 (N_9047,N_4760,N_5564);
or U9048 (N_9048,N_5728,N_7447);
and U9049 (N_9049,N_6448,N_5720);
xor U9050 (N_9050,N_6160,N_6421);
nor U9051 (N_9051,N_5467,N_4837);
xor U9052 (N_9052,N_4046,N_6431);
or U9053 (N_9053,N_5162,N_6131);
or U9054 (N_9054,N_4949,N_5404);
nor U9055 (N_9055,N_6062,N_6760);
nand U9056 (N_9056,N_6930,N_5042);
xor U9057 (N_9057,N_7534,N_5646);
and U9058 (N_9058,N_5058,N_7962);
xor U9059 (N_9059,N_4346,N_4621);
or U9060 (N_9060,N_5376,N_7847);
or U9061 (N_9061,N_4427,N_4501);
nand U9062 (N_9062,N_5971,N_7660);
nor U9063 (N_9063,N_7282,N_4494);
and U9064 (N_9064,N_6402,N_4589);
or U9065 (N_9065,N_6456,N_6734);
xnor U9066 (N_9066,N_7816,N_6274);
nor U9067 (N_9067,N_4541,N_5317);
and U9068 (N_9068,N_7286,N_4742);
and U9069 (N_9069,N_5719,N_4986);
nand U9070 (N_9070,N_7891,N_5054);
nor U9071 (N_9071,N_5447,N_7245);
nand U9072 (N_9072,N_6042,N_5788);
and U9073 (N_9073,N_6898,N_5611);
xor U9074 (N_9074,N_5398,N_6460);
xnor U9075 (N_9075,N_6765,N_5700);
and U9076 (N_9076,N_6130,N_5631);
nand U9077 (N_9077,N_7478,N_5759);
nand U9078 (N_9078,N_4926,N_5586);
nor U9079 (N_9079,N_7015,N_4966);
nand U9080 (N_9080,N_5746,N_4611);
or U9081 (N_9081,N_6728,N_5268);
xnor U9082 (N_9082,N_5130,N_7945);
or U9083 (N_9083,N_7630,N_6461);
or U9084 (N_9084,N_4072,N_4485);
or U9085 (N_9085,N_5209,N_7884);
and U9086 (N_9086,N_7350,N_5458);
and U9087 (N_9087,N_5302,N_4521);
xnor U9088 (N_9088,N_4885,N_4372);
nand U9089 (N_9089,N_6151,N_5811);
nand U9090 (N_9090,N_6409,N_5269);
nor U9091 (N_9091,N_5617,N_4400);
nand U9092 (N_9092,N_6234,N_6550);
and U9093 (N_9093,N_4460,N_7523);
or U9094 (N_9094,N_7798,N_7614);
or U9095 (N_9095,N_7328,N_4004);
or U9096 (N_9096,N_5540,N_4840);
nor U9097 (N_9097,N_4633,N_6429);
or U9098 (N_9098,N_4052,N_6940);
nand U9099 (N_9099,N_4945,N_6908);
xor U9100 (N_9100,N_4833,N_6401);
nand U9101 (N_9101,N_6634,N_7985);
nand U9102 (N_9102,N_7017,N_5704);
and U9103 (N_9103,N_5852,N_7654);
xnor U9104 (N_9104,N_5320,N_4985);
xnor U9105 (N_9105,N_4476,N_6890);
nor U9106 (N_9106,N_6420,N_4467);
and U9107 (N_9107,N_7517,N_7236);
or U9108 (N_9108,N_4995,N_6529);
and U9109 (N_9109,N_4418,N_4277);
and U9110 (N_9110,N_6242,N_7024);
or U9111 (N_9111,N_4293,N_4147);
and U9112 (N_9112,N_7461,N_6657);
nor U9113 (N_9113,N_5016,N_4096);
nand U9114 (N_9114,N_6175,N_4676);
nand U9115 (N_9115,N_5862,N_5418);
xnor U9116 (N_9116,N_4130,N_4200);
nor U9117 (N_9117,N_6792,N_7474);
xnor U9118 (N_9118,N_6689,N_5196);
nand U9119 (N_9119,N_7501,N_6577);
or U9120 (N_9120,N_5827,N_5240);
nor U9121 (N_9121,N_5107,N_6676);
or U9122 (N_9122,N_4420,N_5825);
nor U9123 (N_9123,N_7714,N_4594);
nand U9124 (N_9124,N_4183,N_6710);
xor U9125 (N_9125,N_4652,N_4935);
xor U9126 (N_9126,N_4637,N_4054);
xor U9127 (N_9127,N_6718,N_5790);
nand U9128 (N_9128,N_7659,N_6998);
and U9129 (N_9129,N_4078,N_6644);
or U9130 (N_9130,N_4951,N_4889);
or U9131 (N_9131,N_7010,N_6052);
or U9132 (N_9132,N_5845,N_5615);
nor U9133 (N_9133,N_5894,N_4205);
or U9134 (N_9134,N_6282,N_4291);
and U9135 (N_9135,N_4473,N_4364);
nor U9136 (N_9136,N_6133,N_4335);
xor U9137 (N_9137,N_5869,N_7968);
or U9138 (N_9138,N_6569,N_4093);
xnor U9139 (N_9139,N_4483,N_6884);
nor U9140 (N_9140,N_7671,N_7353);
nor U9141 (N_9141,N_5241,N_7824);
or U9142 (N_9142,N_7915,N_7374);
nand U9143 (N_9143,N_6803,N_7063);
xor U9144 (N_9144,N_4916,N_7105);
and U9145 (N_9145,N_5545,N_6943);
nand U9146 (N_9146,N_4669,N_4535);
or U9147 (N_9147,N_7007,N_5618);
nand U9148 (N_9148,N_5526,N_4057);
or U9149 (N_9149,N_4692,N_7305);
xnor U9150 (N_9150,N_5507,N_6609);
nand U9151 (N_9151,N_5129,N_4402);
nand U9152 (N_9152,N_7515,N_5219);
and U9153 (N_9153,N_5112,N_4509);
nand U9154 (N_9154,N_6482,N_4874);
nand U9155 (N_9155,N_4794,N_5997);
and U9156 (N_9156,N_7856,N_4898);
nor U9157 (N_9157,N_6440,N_6927);
and U9158 (N_9158,N_5925,N_7301);
or U9159 (N_9159,N_4867,N_7174);
and U9160 (N_9160,N_5109,N_7172);
nand U9161 (N_9161,N_5691,N_7146);
nor U9162 (N_9162,N_7656,N_7115);
nand U9163 (N_9163,N_6255,N_5150);
nor U9164 (N_9164,N_6856,N_4303);
or U9165 (N_9165,N_5466,N_7143);
xnor U9166 (N_9166,N_6987,N_5713);
and U9167 (N_9167,N_4939,N_5451);
xor U9168 (N_9168,N_4917,N_4475);
and U9169 (N_9169,N_7570,N_5774);
xnor U9170 (N_9170,N_4285,N_7130);
nor U9171 (N_9171,N_7794,N_7805);
or U9172 (N_9172,N_4273,N_4195);
nor U9173 (N_9173,N_6243,N_7221);
xnor U9174 (N_9174,N_5110,N_7518);
and U9175 (N_9175,N_4967,N_4440);
xor U9176 (N_9176,N_5830,N_4539);
nor U9177 (N_9177,N_6751,N_4108);
nand U9178 (N_9178,N_5698,N_7373);
nor U9179 (N_9179,N_7574,N_5699);
and U9180 (N_9180,N_7224,N_6272);
xor U9181 (N_9181,N_7298,N_7109);
and U9182 (N_9182,N_4530,N_7243);
nor U9183 (N_9183,N_5344,N_5221);
and U9184 (N_9184,N_5742,N_4891);
or U9185 (N_9185,N_4405,N_6822);
nor U9186 (N_9186,N_6790,N_5010);
xor U9187 (N_9187,N_5783,N_4987);
or U9188 (N_9188,N_6591,N_5892);
nand U9189 (N_9189,N_7568,N_7091);
xnor U9190 (N_9190,N_7212,N_4512);
and U9191 (N_9191,N_4567,N_7029);
or U9192 (N_9192,N_5577,N_4249);
or U9193 (N_9193,N_4401,N_5406);
xor U9194 (N_9194,N_5576,N_6294);
nor U9195 (N_9195,N_7773,N_7356);
nor U9196 (N_9196,N_4069,N_6937);
nand U9197 (N_9197,N_5641,N_5046);
nor U9198 (N_9198,N_5834,N_6083);
nor U9199 (N_9199,N_4295,N_6827);
nand U9200 (N_9200,N_7763,N_5329);
nand U9201 (N_9201,N_7074,N_5155);
nor U9202 (N_9202,N_4234,N_4009);
xnor U9203 (N_9203,N_6008,N_6449);
or U9204 (N_9204,N_6488,N_5476);
and U9205 (N_9205,N_4759,N_7270);
or U9206 (N_9206,N_6922,N_7097);
xnor U9207 (N_9207,N_4118,N_6017);
and U9208 (N_9208,N_7801,N_4550);
and U9209 (N_9209,N_6825,N_4309);
nand U9210 (N_9210,N_5063,N_7341);
xnor U9211 (N_9211,N_4199,N_4720);
xor U9212 (N_9212,N_6349,N_7289);
xor U9213 (N_9213,N_5508,N_6837);
nand U9214 (N_9214,N_4690,N_7446);
nor U9215 (N_9215,N_5907,N_6791);
and U9216 (N_9216,N_5044,N_5388);
or U9217 (N_9217,N_5977,N_7265);
xor U9218 (N_9218,N_4013,N_5353);
nor U9219 (N_9219,N_6106,N_5190);
nor U9220 (N_9220,N_6315,N_5908);
xnor U9221 (N_9221,N_4311,N_4250);
and U9222 (N_9222,N_7608,N_7835);
nand U9223 (N_9223,N_7917,N_6548);
and U9224 (N_9224,N_4175,N_6328);
xor U9225 (N_9225,N_6848,N_6817);
or U9226 (N_9226,N_5762,N_7119);
nand U9227 (N_9227,N_7387,N_5921);
and U9228 (N_9228,N_7765,N_7194);
and U9229 (N_9229,N_4227,N_4918);
nor U9230 (N_9230,N_4960,N_4464);
nand U9231 (N_9231,N_7340,N_6870);
or U9232 (N_9232,N_4025,N_5513);
and U9233 (N_9233,N_4726,N_5313);
or U9234 (N_9234,N_4051,N_5004);
and U9235 (N_9235,N_4937,N_6662);
or U9236 (N_9236,N_6395,N_7096);
xor U9237 (N_9237,N_7786,N_5515);
or U9238 (N_9238,N_4036,N_6279);
or U9239 (N_9239,N_6780,N_7322);
or U9240 (N_9240,N_5187,N_7035);
and U9241 (N_9241,N_4179,N_7427);
or U9242 (N_9242,N_5733,N_6646);
or U9243 (N_9243,N_5030,N_6690);
xnor U9244 (N_9244,N_5695,N_6852);
nor U9245 (N_9245,N_5164,N_7909);
nand U9246 (N_9246,N_5781,N_6984);
or U9247 (N_9247,N_6632,N_4639);
and U9248 (N_9248,N_7959,N_5858);
xor U9249 (N_9249,N_4764,N_7011);
nor U9250 (N_9250,N_5732,N_7871);
nor U9251 (N_9251,N_5198,N_5649);
or U9252 (N_9252,N_7161,N_6221);
nand U9253 (N_9253,N_5629,N_5884);
nor U9254 (N_9254,N_6426,N_4658);
nor U9255 (N_9255,N_6872,N_7054);
nand U9256 (N_9256,N_5349,N_4941);
nand U9257 (N_9257,N_4537,N_7257);
xnor U9258 (N_9258,N_6533,N_6267);
nor U9259 (N_9259,N_6906,N_7648);
xnor U9260 (N_9260,N_5727,N_7401);
nand U9261 (N_9261,N_4167,N_5251);
xnor U9262 (N_9262,N_4607,N_4341);
nor U9263 (N_9263,N_4569,N_4053);
xnor U9264 (N_9264,N_5948,N_5635);
nand U9265 (N_9265,N_5381,N_7220);
or U9266 (N_9266,N_4134,N_4657);
nor U9267 (N_9267,N_7099,N_6801);
or U9268 (N_9268,N_4128,N_6403);
xnor U9269 (N_9269,N_7508,N_5865);
and U9270 (N_9270,N_7936,N_6919);
xnor U9271 (N_9271,N_6300,N_5803);
and U9272 (N_9272,N_6210,N_7949);
xnor U9273 (N_9273,N_5108,N_4135);
and U9274 (N_9274,N_6830,N_7947);
or U9275 (N_9275,N_7638,N_5950);
nand U9276 (N_9276,N_4492,N_7529);
or U9277 (N_9277,N_6320,N_5511);
nand U9278 (N_9278,N_6938,N_5140);
or U9279 (N_9279,N_7306,N_4033);
and U9280 (N_9280,N_4981,N_6027);
or U9281 (N_9281,N_5949,N_5050);
nand U9282 (N_9282,N_5242,N_4196);
nor U9283 (N_9283,N_5760,N_4599);
nand U9284 (N_9284,N_6778,N_7760);
xnor U9285 (N_9285,N_7684,N_7012);
nor U9286 (N_9286,N_6091,N_7997);
or U9287 (N_9287,N_7254,N_5542);
nand U9288 (N_9288,N_4417,N_4597);
nor U9289 (N_9289,N_4465,N_4353);
or U9290 (N_9290,N_7354,N_5333);
nor U9291 (N_9291,N_7722,N_5125);
xnor U9292 (N_9292,N_4474,N_7955);
xnor U9293 (N_9293,N_6724,N_5608);
or U9294 (N_9294,N_4454,N_5118);
xnor U9295 (N_9295,N_5347,N_5522);
nor U9296 (N_9296,N_5456,N_4913);
and U9297 (N_9297,N_4765,N_6020);
or U9298 (N_9298,N_4445,N_7640);
nor U9299 (N_9299,N_5337,N_5851);
nand U9300 (N_9300,N_7850,N_7730);
or U9301 (N_9301,N_4834,N_7360);
nor U9302 (N_9302,N_6444,N_6356);
and U9303 (N_9303,N_6554,N_4780);
or U9304 (N_9304,N_7177,N_6547);
nand U9305 (N_9305,N_5071,N_5173);
xor U9306 (N_9306,N_4262,N_5986);
nand U9307 (N_9307,N_4165,N_7227);
and U9308 (N_9308,N_4456,N_5944);
or U9309 (N_9309,N_7274,N_4797);
and U9310 (N_9310,N_7673,N_7633);
and U9311 (N_9311,N_7127,N_6652);
nand U9312 (N_9312,N_7281,N_6216);
nor U9313 (N_9313,N_5730,N_4561);
nand U9314 (N_9314,N_6469,N_6843);
nand U9315 (N_9315,N_4000,N_7498);
xnor U9316 (N_9316,N_7337,N_7753);
xor U9317 (N_9317,N_7832,N_7670);
nand U9318 (N_9318,N_7992,N_5354);
and U9319 (N_9319,N_6486,N_6581);
xor U9320 (N_9320,N_7941,N_7363);
nand U9321 (N_9321,N_4542,N_6821);
and U9322 (N_9322,N_6975,N_5059);
and U9323 (N_9323,N_4296,N_4133);
or U9324 (N_9324,N_7038,N_5796);
xnor U9325 (N_9325,N_7396,N_5512);
and U9326 (N_9326,N_6725,N_5183);
nand U9327 (N_9327,N_7025,N_6154);
xor U9328 (N_9328,N_4725,N_5128);
nor U9329 (N_9329,N_5609,N_7428);
xor U9330 (N_9330,N_5267,N_7171);
nor U9331 (N_9331,N_5484,N_7929);
or U9332 (N_9332,N_5505,N_7637);
nor U9333 (N_9333,N_4975,N_7688);
and U9334 (N_9334,N_7755,N_4560);
or U9335 (N_9335,N_4322,N_5569);
nand U9336 (N_9336,N_4841,N_5303);
or U9337 (N_9337,N_6201,N_5913);
and U9338 (N_9338,N_5859,N_4784);
and U9339 (N_9339,N_4686,N_5496);
or U9340 (N_9340,N_7443,N_6423);
xnor U9341 (N_9341,N_6465,N_4576);
xor U9342 (N_9342,N_6711,N_6197);
or U9343 (N_9343,N_5022,N_4822);
and U9344 (N_9344,N_7211,N_7841);
nor U9345 (N_9345,N_5248,N_7076);
nand U9346 (N_9346,N_4479,N_4371);
nor U9347 (N_9347,N_5808,N_7078);
nand U9348 (N_9348,N_6307,N_4015);
nand U9349 (N_9349,N_7519,N_4029);
and U9350 (N_9350,N_4508,N_4654);
nor U9351 (N_9351,N_7272,N_5380);
nor U9352 (N_9352,N_6288,N_7544);
xnor U9353 (N_9353,N_4367,N_6625);
nor U9354 (N_9354,N_4545,N_6944);
nand U9355 (N_9355,N_5047,N_6527);
xnor U9356 (N_9356,N_6211,N_7468);
nor U9357 (N_9357,N_7925,N_7785);
and U9358 (N_9358,N_7635,N_4655);
and U9359 (N_9359,N_4843,N_6046);
xnor U9360 (N_9360,N_5812,N_5778);
nand U9361 (N_9361,N_7357,N_6526);
or U9362 (N_9362,N_5189,N_6084);
nor U9363 (N_9363,N_6014,N_5572);
xnor U9364 (N_9364,N_5245,N_5408);
and U9365 (N_9365,N_5628,N_5573);
or U9366 (N_9366,N_6806,N_5660);
and U9367 (N_9367,N_5165,N_6514);
or U9368 (N_9368,N_7628,N_7964);
or U9369 (N_9369,N_6844,N_5636);
or U9370 (N_9370,N_5659,N_5620);
xor U9371 (N_9371,N_7536,N_4403);
nand U9372 (N_9372,N_7325,N_6913);
nor U9373 (N_9373,N_7881,N_6172);
nor U9374 (N_9374,N_6441,N_5282);
nand U9375 (N_9375,N_7913,N_6099);
xnor U9376 (N_9376,N_7603,N_5049);
xnor U9377 (N_9377,N_6694,N_4605);
or U9378 (N_9378,N_6392,N_6496);
nand U9379 (N_9379,N_5669,N_4831);
or U9380 (N_9380,N_6797,N_7460);
xnor U9381 (N_9381,N_7135,N_6445);
nor U9382 (N_9382,N_4744,N_6068);
or U9383 (N_9383,N_6973,N_7482);
nor U9384 (N_9384,N_4239,N_4363);
nor U9385 (N_9385,N_4230,N_7030);
nor U9386 (N_9386,N_6229,N_6595);
xnor U9387 (N_9387,N_4256,N_6481);
nand U9388 (N_9388,N_5495,N_7547);
nand U9389 (N_9389,N_7713,N_5679);
or U9390 (N_9390,N_6682,N_6111);
nor U9391 (N_9391,N_6877,N_4683);
and U9392 (N_9392,N_5364,N_5481);
or U9393 (N_9393,N_6875,N_7262);
or U9394 (N_9394,N_6261,N_6519);
nor U9395 (N_9395,N_5685,N_7858);
xnor U9396 (N_9396,N_5223,N_5502);
or U9397 (N_9397,N_6348,N_4264);
and U9398 (N_9398,N_5784,N_7716);
xor U9399 (N_9399,N_5390,N_4027);
or U9400 (N_9400,N_5506,N_7859);
nand U9401 (N_9401,N_7457,N_4983);
and U9402 (N_9402,N_7907,N_4314);
or U9403 (N_9403,N_6126,N_5519);
and U9404 (N_9404,N_6225,N_6277);
xor U9405 (N_9405,N_4579,N_7808);
and U9406 (N_9406,N_6942,N_4436);
and U9407 (N_9407,N_5527,N_4912);
xor U9408 (N_9408,N_6911,N_4739);
nor U9409 (N_9409,N_6809,N_4587);
or U9410 (N_9410,N_4856,N_4289);
or U9411 (N_9411,N_7201,N_4847);
or U9412 (N_9412,N_4398,N_6874);
nor U9413 (N_9413,N_6846,N_4399);
xor U9414 (N_9414,N_4890,N_5247);
xor U9415 (N_9415,N_7316,N_4201);
nand U9416 (N_9416,N_7215,N_6860);
nand U9417 (N_9417,N_5887,N_5351);
nand U9418 (N_9418,N_4319,N_6851);
and U9419 (N_9419,N_7616,N_5166);
xor U9420 (N_9420,N_4119,N_5457);
nor U9421 (N_9421,N_4162,N_6627);
xnor U9422 (N_9422,N_5717,N_7087);
nor U9423 (N_9423,N_6893,N_7004);
and U9424 (N_9424,N_6793,N_7210);
nor U9425 (N_9425,N_6391,N_4925);
nand U9426 (N_9426,N_7735,N_5252);
or U9427 (N_9427,N_7624,N_4991);
or U9428 (N_9428,N_6184,N_5332);
or U9429 (N_9429,N_5702,N_7413);
nor U9430 (N_9430,N_6275,N_5226);
or U9431 (N_9431,N_7503,N_5962);
or U9432 (N_9432,N_5002,N_4581);
or U9433 (N_9433,N_4097,N_4933);
or U9434 (N_9434,N_6604,N_5220);
and U9435 (N_9435,N_4704,N_5797);
nand U9436 (N_9436,N_7852,N_4449);
and U9437 (N_9437,N_6110,N_6093);
or U9438 (N_9438,N_4378,N_5585);
and U9439 (N_9439,N_4534,N_6935);
nor U9440 (N_9440,N_5967,N_6003);
nand U9441 (N_9441,N_6443,N_4979);
xnor U9442 (N_9442,N_6859,N_4389);
or U9443 (N_9443,N_6244,N_6643);
nand U9444 (N_9444,N_7082,N_6811);
nor U9445 (N_9445,N_6626,N_5237);
and U9446 (N_9446,N_6608,N_5514);
nand U9447 (N_9447,N_4098,N_7771);
xnor U9448 (N_9448,N_6476,N_6945);
xor U9449 (N_9449,N_4635,N_4044);
xnor U9450 (N_9450,N_4824,N_7663);
or U9451 (N_9451,N_6845,N_4540);
nand U9452 (N_9452,N_6305,N_5429);
or U9453 (N_9453,N_5817,N_7318);
nand U9454 (N_9454,N_5018,N_6818);
xnor U9455 (N_9455,N_4173,N_5160);
or U9456 (N_9456,N_7782,N_4373);
and U9457 (N_9457,N_6226,N_5065);
nand U9458 (N_9458,N_4144,N_6596);
nand U9459 (N_9459,N_5565,N_5975);
or U9460 (N_9460,N_7093,N_4515);
and U9461 (N_9461,N_5974,N_7552);
nor U9462 (N_9462,N_4076,N_7392);
and U9463 (N_9463,N_6321,N_7238);
and U9464 (N_9464,N_5917,N_4584);
and U9465 (N_9465,N_5584,N_7149);
xor U9466 (N_9466,N_6302,N_6768);
xnor U9467 (N_9467,N_7279,N_7165);
nor U9468 (N_9468,N_4442,N_5772);
xor U9469 (N_9469,N_7331,N_6829);
or U9470 (N_9470,N_4769,N_5038);
xor U9471 (N_9471,N_5960,N_4430);
xor U9472 (N_9472,N_6422,N_4302);
xor U9473 (N_9473,N_5721,N_5285);
xnor U9474 (N_9474,N_7844,N_5546);
and U9475 (N_9475,N_7792,N_5473);
xor U9476 (N_9476,N_6491,N_6952);
and U9477 (N_9477,N_6871,N_5567);
or U9478 (N_9478,N_7950,N_4301);
and U9479 (N_9479,N_7390,N_4342);
nand U9480 (N_9480,N_7514,N_6345);
nor U9481 (N_9481,N_5075,N_4287);
xor U9482 (N_9482,N_5186,N_6459);
nor U9483 (N_9483,N_7979,N_6555);
or U9484 (N_9484,N_4181,N_6907);
or U9485 (N_9485,N_4444,N_5283);
nor U9486 (N_9486,N_7507,N_6688);
xor U9487 (N_9487,N_4533,N_6299);
nor U9488 (N_9488,N_4601,N_5984);
nand U9489 (N_9489,N_7170,N_5773);
nor U9490 (N_9490,N_5739,N_7889);
nor U9491 (N_9491,N_7155,N_5392);
xnor U9492 (N_9492,N_7190,N_4313);
and U9493 (N_9493,N_5171,N_4374);
or U9494 (N_9494,N_6576,N_6642);
nand U9495 (N_9495,N_7956,N_4953);
nor U9496 (N_9496,N_7821,N_4641);
nor U9497 (N_9497,N_5664,N_7116);
and U9498 (N_9498,N_7695,N_5610);
nor U9499 (N_9499,N_6589,N_7721);
or U9500 (N_9500,N_6926,N_6208);
or U9501 (N_9501,N_4528,N_6712);
or U9502 (N_9502,N_7113,N_4549);
nor U9503 (N_9503,N_4740,N_4259);
nor U9504 (N_9504,N_5318,N_4120);
xor U9505 (N_9505,N_5580,N_7866);
xnor U9506 (N_9506,N_5998,N_4104);
nand U9507 (N_9507,N_6738,N_5026);
or U9508 (N_9508,N_5474,N_7391);
xnor U9509 (N_9509,N_6566,N_7121);
xnor U9510 (N_9510,N_7108,N_7657);
nor U9511 (N_9511,N_5559,N_6733);
and U9512 (N_9512,N_7543,N_4014);
nor U9513 (N_9513,N_7768,N_5202);
nand U9514 (N_9514,N_6418,N_6996);
nor U9515 (N_9515,N_6865,N_5000);
and U9516 (N_9516,N_4963,N_6209);
xor U9517 (N_9517,N_6375,N_7047);
and U9518 (N_9518,N_4307,N_4001);
and U9519 (N_9519,N_4562,N_6896);
and U9520 (N_9520,N_4957,N_6636);
nand U9521 (N_9521,N_5092,N_6873);
nand U9522 (N_9522,N_5045,N_5818);
nand U9523 (N_9523,N_5878,N_7770);
and U9524 (N_9524,N_4736,N_4413);
or U9525 (N_9525,N_5587,N_7578);
and U9526 (N_9526,N_4347,N_7062);
nor U9527 (N_9527,N_6598,N_5547);
or U9528 (N_9528,N_6158,N_4141);
and U9529 (N_9529,N_4260,N_7791);
or U9530 (N_9530,N_6719,N_5745);
and U9531 (N_9531,N_6372,N_4767);
nor U9532 (N_9532,N_7861,N_7601);
or U9533 (N_9533,N_4758,N_5169);
and U9534 (N_9534,N_6631,N_7697);
nand U9535 (N_9535,N_5483,N_7796);
nand U9536 (N_9536,N_5837,N_5839);
and U9537 (N_9537,N_7617,N_5672);
or U9538 (N_9538,N_7899,N_5785);
or U9539 (N_9539,N_7206,N_4238);
and U9540 (N_9540,N_4902,N_4457);
and U9541 (N_9541,N_6978,N_4749);
xnor U9542 (N_9542,N_5658,N_4255);
or U9543 (N_9543,N_6451,N_4773);
nor U9544 (N_9544,N_5104,N_4079);
nand U9545 (N_9545,N_5718,N_5086);
or U9546 (N_9546,N_7208,N_4151);
nand U9547 (N_9547,N_7014,N_7264);
nor U9548 (N_9548,N_6677,N_5278);
or U9549 (N_9549,N_4518,N_5216);
nor U9550 (N_9550,N_4711,N_7739);
and U9551 (N_9551,N_5655,N_6447);
nand U9552 (N_9552,N_5322,N_4663);
xnor U9553 (N_9553,N_6452,N_6264);
nor U9554 (N_9554,N_4615,N_4858);
xnor U9555 (N_9555,N_6359,N_5446);
and U9556 (N_9556,N_7114,N_7542);
xnor U9557 (N_9557,N_7366,N_5771);
nand U9558 (N_9558,N_6329,N_4506);
nor U9559 (N_9559,N_4944,N_7748);
xnor U9560 (N_9560,N_6854,N_5312);
nand U9561 (N_9561,N_6435,N_5786);
nor U9562 (N_9562,N_6731,N_6833);
xnor U9563 (N_9563,N_5450,N_4450);
nor U9564 (N_9564,N_4282,N_5199);
or U9565 (N_9565,N_7521,N_5776);
xnor U9566 (N_9566,N_7436,N_5942);
nand U9567 (N_9567,N_6071,N_7685);
and U9568 (N_9568,N_5177,N_5604);
or U9569 (N_9569,N_6696,N_6824);
and U9570 (N_9570,N_5469,N_4286);
xnor U9571 (N_9571,N_6180,N_5095);
xor U9572 (N_9572,N_4397,N_6592);
nor U9573 (N_9573,N_4003,N_6523);
and U9574 (N_9574,N_5340,N_6270);
nor U9575 (N_9575,N_4109,N_6695);
nand U9576 (N_9576,N_5614,N_7618);
and U9577 (N_9577,N_4931,N_4324);
nor U9578 (N_9578,N_5898,N_4796);
xor U9579 (N_9579,N_5041,N_7779);
xnor U9580 (N_9580,N_4217,N_5675);
xor U9581 (N_9581,N_7352,N_7084);
and U9582 (N_9582,N_6048,N_7488);
and U9583 (N_9583,N_7134,N_6212);
and U9584 (N_9584,N_6714,N_4496);
xnor U9585 (N_9585,N_5626,N_5594);
nor U9586 (N_9586,N_5856,N_4735);
nand U9587 (N_9587,N_4166,N_4538);
nand U9588 (N_9588,N_7042,N_4978);
nand U9589 (N_9589,N_7051,N_5558);
or U9590 (N_9590,N_5815,N_6268);
or U9591 (N_9591,N_4741,N_4915);
or U9592 (N_9592,N_7857,N_7417);
xor U9593 (N_9593,N_5091,N_5273);
nor U9594 (N_9594,N_6761,N_5822);
or U9595 (N_9595,N_7976,N_7586);
and U9596 (N_9596,N_7870,N_7818);
nor U9597 (N_9597,N_4094,N_6080);
and U9598 (N_9598,N_4252,N_7894);
xor U9599 (N_9599,N_7202,N_4614);
nor U9600 (N_9600,N_4089,N_4507);
and U9601 (N_9601,N_5005,N_4779);
nand U9602 (N_9602,N_5554,N_4178);
nand U9603 (N_9603,N_6615,N_7152);
or U9604 (N_9604,N_6358,N_7180);
nand U9605 (N_9605,N_7209,N_4192);
nand U9606 (N_9606,N_5697,N_4149);
and U9607 (N_9607,N_7083,N_7963);
nand U9608 (N_9608,N_5870,N_5682);
nor U9609 (N_9609,N_7140,N_7081);
nor U9610 (N_9610,N_6433,N_6147);
or U9611 (N_9611,N_7342,N_4795);
and U9612 (N_9612,N_4171,N_6332);
and U9613 (N_9613,N_5553,N_5294);
and U9614 (N_9614,N_5566,N_4247);
xnor U9615 (N_9615,N_6571,N_6993);
xor U9616 (N_9616,N_6075,N_4254);
nor U9617 (N_9617,N_4431,N_7123);
nor U9618 (N_9618,N_6892,N_4404);
nor U9619 (N_9619,N_7541,N_6767);
nor U9620 (N_9620,N_7888,N_7003);
and U9621 (N_9621,N_5871,N_5460);
nor U9622 (N_9622,N_6986,N_5074);
nand U9623 (N_9623,N_6656,N_4132);
nand U9624 (N_9624,N_4804,N_5552);
nand U9625 (N_9625,N_7729,N_6955);
or U9626 (N_9626,N_6610,N_6499);
and U9627 (N_9627,N_6939,N_4861);
and U9628 (N_9628,N_5612,N_7246);
and U9629 (N_9629,N_4323,N_5806);
nand U9630 (N_9630,N_4724,N_7408);
nand U9631 (N_9631,N_6024,N_7511);
nand U9632 (N_9632,N_5603,N_6164);
xor U9633 (N_9633,N_7151,N_5840);
xor U9634 (N_9634,N_5985,N_4554);
or U9635 (N_9635,N_6508,N_7641);
nand U9636 (N_9636,N_4102,N_5729);
and U9637 (N_9637,N_7486,N_4113);
nor U9638 (N_9638,N_6051,N_4137);
nand U9639 (N_9639,N_6129,N_6994);
xor U9640 (N_9640,N_5486,N_5875);
or U9641 (N_9641,N_6883,N_5439);
nand U9642 (N_9642,N_7761,N_4632);
or U9643 (N_9643,N_7619,N_6771);
nand U9644 (N_9644,N_6808,N_6463);
nand U9645 (N_9645,N_6428,N_4908);
nor U9646 (N_9646,N_7462,N_7509);
nand U9647 (N_9647,N_4809,N_6507);
nand U9648 (N_9648,N_7291,N_4640);
xnor U9649 (N_9649,N_6181,N_4490);
xor U9650 (N_9650,N_5069,N_6759);
xor U9651 (N_9651,N_6574,N_6495);
or U9652 (N_9652,N_5556,N_4383);
or U9653 (N_9653,N_6777,N_5562);
or U9654 (N_9654,N_5048,N_6606);
nand U9655 (N_9655,N_4609,N_6489);
nor U9656 (N_9656,N_5828,N_6957);
and U9657 (N_9657,N_5144,N_5651);
xnor U9658 (N_9658,N_6173,N_5024);
or U9659 (N_9659,N_7005,N_4832);
nor U9660 (N_9660,N_5192,N_6618);
nor U9661 (N_9661,N_4730,N_7762);
nand U9662 (N_9662,N_5346,N_7605);
or U9663 (N_9663,N_4182,N_7799);
nor U9664 (N_9664,N_4208,N_6820);
nor U9665 (N_9665,N_4428,N_7712);
and U9666 (N_9666,N_5810,N_6417);
xnor U9667 (N_9667,N_5370,N_5152);
xnor U9668 (N_9668,N_6354,N_6649);
or U9669 (N_9669,N_5325,N_6534);
and U9670 (N_9670,N_4888,N_4783);
and U9671 (N_9671,N_5180,N_6480);
nor U9672 (N_9672,N_5775,N_6235);
nand U9673 (N_9673,N_7252,N_6568);
nand U9674 (N_9674,N_4123,N_5078);
or U9675 (N_9675,N_4762,N_7057);
xor U9676 (N_9676,N_4934,N_4993);
and U9677 (N_9677,N_7223,N_7300);
xor U9678 (N_9678,N_4158,N_4176);
nor U9679 (N_9679,N_7144,N_6756);
or U9680 (N_9680,N_7050,N_5684);
xnor U9681 (N_9681,N_7440,N_7169);
nand U9682 (N_9682,N_6379,N_4315);
nand U9683 (N_9683,N_4340,N_6739);
and U9684 (N_9684,N_6479,N_4328);
xnor U9685 (N_9685,N_4952,N_5498);
nor U9686 (N_9686,N_7295,N_4443);
xor U9687 (N_9687,N_4056,N_7419);
xnor U9688 (N_9688,N_5409,N_4491);
and U9689 (N_9689,N_7141,N_7845);
nor U9690 (N_9690,N_5798,N_5433);
nor U9691 (N_9691,N_5937,N_7027);
or U9692 (N_9692,N_5139,N_5863);
and U9693 (N_9693,N_7918,N_5534);
nand U9694 (N_9694,N_5890,N_7188);
or U9695 (N_9695,N_7951,N_4628);
xnor U9696 (N_9696,N_7423,N_7890);
or U9697 (N_9697,N_6041,N_6374);
nor U9698 (N_9698,N_4349,N_7572);
or U9699 (N_9699,N_6723,N_5203);
or U9700 (N_9700,N_5953,N_6314);
nand U9701 (N_9701,N_4484,N_5600);
nand U9702 (N_9702,N_4300,N_5464);
nor U9703 (N_9703,N_4088,N_4828);
xor U9704 (N_9704,N_5153,N_6033);
xnor U9705 (N_9705,N_7998,N_6232);
xnor U9706 (N_9706,N_6458,N_5291);
and U9707 (N_9707,N_4068,N_6047);
xor U9708 (N_9708,N_4748,N_5287);
xor U9709 (N_9709,N_6786,N_4163);
or U9710 (N_9710,N_4830,N_6285);
nand U9711 (N_9711,N_7993,N_4950);
nand U9712 (N_9712,N_6968,N_4648);
and U9713 (N_9713,N_6842,N_4845);
nor U9714 (N_9714,N_4850,N_6037);
xor U9715 (N_9715,N_7759,N_6257);
xnor U9716 (N_9716,N_7379,N_4278);
nand U9717 (N_9717,N_4269,N_4901);
or U9718 (N_9718,N_6635,N_4352);
xor U9719 (N_9719,N_5435,N_4585);
and U9720 (N_9720,N_5861,N_4489);
nand U9721 (N_9721,N_6981,N_7275);
xor U9722 (N_9722,N_7715,N_7812);
xnor U9723 (N_9723,N_6074,N_4355);
and U9724 (N_9724,N_4989,N_4712);
and U9725 (N_9725,N_5254,N_5417);
xnor U9726 (N_9726,N_6324,N_5468);
xnor U9727 (N_9727,N_7682,N_7406);
nor U9728 (N_9728,N_7022,N_7764);
or U9729 (N_9729,N_5543,N_6018);
or U9730 (N_9730,N_7658,N_6176);
nor U9731 (N_9731,N_6404,N_5448);
or U9732 (N_9732,N_7106,N_5359);
nor U9733 (N_9733,N_4187,N_5832);
or U9734 (N_9734,N_5025,N_4281);
xor U9735 (N_9735,N_6336,N_4150);
and U9736 (N_9736,N_6424,N_5228);
nand U9737 (N_9737,N_5402,N_5453);
or U9738 (N_9738,N_4063,N_7294);
or U9739 (N_9739,N_4288,N_5625);
nand U9740 (N_9740,N_6370,N_4359);
nand U9741 (N_9741,N_5748,N_4977);
xor U9742 (N_9742,N_4336,N_4242);
nand U9743 (N_9743,N_5874,N_5098);
xor U9744 (N_9744,N_6289,N_7526);
nand U9745 (N_9745,N_6800,N_6967);
xnor U9746 (N_9746,N_5132,N_5081);
and U9747 (N_9747,N_5341,N_4411);
and U9748 (N_9748,N_4819,N_7686);
nor U9749 (N_9749,N_7370,N_7228);
xnor U9750 (N_9750,N_7071,N_6493);
nand U9751 (N_9751,N_6470,N_4368);
nand U9752 (N_9752,N_5801,N_4778);
nand U9753 (N_9753,N_7435,N_7906);
xnor U9754 (N_9754,N_6291,N_4752);
or U9755 (N_9755,N_4274,N_5749);
nor U9756 (N_9756,N_6161,N_4709);
or U9757 (N_9757,N_5653,N_5793);
xor U9758 (N_9758,N_5814,N_6055);
or U9759 (N_9759,N_5938,N_6858);
nand U9760 (N_9760,N_6498,N_7734);
nand U9761 (N_9761,N_7694,N_4191);
nand U9762 (N_9762,N_5555,N_5372);
nand U9763 (N_9763,N_4817,N_4471);
nand U9764 (N_9764,N_7247,N_6310);
or U9765 (N_9765,N_6252,N_7377);
nor U9766 (N_9766,N_5350,N_7310);
or U9767 (N_9767,N_7470,N_7471);
xnor U9768 (N_9768,N_7932,N_7708);
nor U9769 (N_9769,N_6170,N_7388);
xnor U9770 (N_9770,N_6340,N_6546);
nand U9771 (N_9771,N_4186,N_7125);
and U9772 (N_9772,N_5886,N_7139);
nor U9773 (N_9773,N_7064,N_6241);
nand U9774 (N_9774,N_7830,N_4568);
or U9775 (N_9775,N_7132,N_6956);
or U9776 (N_9776,N_7182,N_4329);
nor U9777 (N_9777,N_6764,N_4719);
or U9778 (N_9778,N_4623,N_5640);
nand U9779 (N_9779,N_5497,N_4152);
xor U9780 (N_9780,N_7372,N_5298);
nand U9781 (N_9781,N_6983,N_4645);
or U9782 (N_9782,N_7110,N_6035);
or U9783 (N_9783,N_5877,N_7696);
and U9784 (N_9784,N_7459,N_7187);
or U9785 (N_9785,N_6139,N_6078);
nand U9786 (N_9786,N_4043,N_7358);
nor U9787 (N_9787,N_7052,N_4721);
and U9788 (N_9788,N_5946,N_5897);
nand U9789 (N_9789,N_5009,N_6612);
nand U9790 (N_9790,N_5407,N_7877);
nor U9791 (N_9791,N_4574,N_5397);
or U9792 (N_9792,N_6500,N_7111);
or U9793 (N_9793,N_7159,N_4468);
nand U9794 (N_9794,N_6655,N_7094);
and U9795 (N_9795,N_7901,N_7653);
and U9796 (N_9796,N_6717,N_4140);
nor U9797 (N_9797,N_6840,N_6492);
xnor U9798 (N_9798,N_6929,N_4630);
or U9799 (N_9799,N_6346,N_5280);
nor U9800 (N_9800,N_4433,N_4974);
nand U9801 (N_9801,N_6979,N_5673);
nand U9802 (N_9802,N_5403,N_4972);
nor U9803 (N_9803,N_7872,N_7595);
nand U9804 (N_9804,N_6995,N_5119);
nand U9805 (N_9805,N_4497,N_4077);
or U9806 (N_9806,N_5120,N_6437);
nor U9807 (N_9807,N_6538,N_5680);
and U9808 (N_9808,N_6355,N_6607);
xor U9809 (N_9809,N_5990,N_4629);
and U9810 (N_9810,N_5314,N_5582);
nand U9811 (N_9811,N_5161,N_7283);
nand U9812 (N_9812,N_5876,N_7726);
or U9813 (N_9813,N_7565,N_6202);
or U9814 (N_9814,N_5434,N_6659);
or U9815 (N_9815,N_4575,N_7583);
and U9816 (N_9816,N_6562,N_5597);
xnor U9817 (N_9817,N_4032,N_4101);
nand U9818 (N_9818,N_7596,N_7303);
nor U9819 (N_9819,N_4361,N_6506);
nand U9820 (N_9820,N_5560,N_7814);
xor U9821 (N_9821,N_5345,N_5864);
xor U9822 (N_9822,N_4929,N_7260);
xor U9823 (N_9823,N_6380,N_7724);
xnor U9824 (N_9824,N_6188,N_6114);
nor U9825 (N_9825,N_6847,N_6752);
nor U9826 (N_9826,N_4900,N_4330);
xnor U9827 (N_9827,N_4298,N_7650);
and U9828 (N_9828,N_5927,N_4923);
nand U9829 (N_9829,N_4207,N_7933);
nor U9830 (N_9830,N_6063,N_5232);
or U9831 (N_9831,N_6036,N_4435);
nor U9832 (N_9832,N_4879,N_6960);
nor U9833 (N_9833,N_5724,N_6138);
and U9834 (N_9834,N_6101,N_7414);
nand U9835 (N_9835,N_7581,N_4516);
nand U9836 (N_9836,N_4169,N_4090);
xnor U9837 (N_9837,N_7145,N_5737);
nand U9838 (N_9838,N_7200,N_7213);
or U9839 (N_9839,N_5920,N_6313);
and U9840 (N_9840,N_5711,N_5694);
xnor U9841 (N_9841,N_6704,N_7324);
nor U9842 (N_9842,N_7450,N_4271);
nand U9843 (N_9843,N_4312,N_4126);
nor U9844 (N_9844,N_5976,N_7160);
and U9845 (N_9845,N_6838,N_5590);
nor U9846 (N_9846,N_6788,N_4071);
and U9847 (N_9847,N_5455,N_7854);
and U9848 (N_9848,N_6319,N_5992);
nand U9849 (N_9849,N_5027,N_7344);
and U9850 (N_9850,N_6108,N_6049);
nor U9851 (N_9851,N_4849,N_6189);
xor U9852 (N_9852,N_6166,N_4586);
nor U9853 (N_9853,N_5255,N_5145);
xor U9854 (N_9854,N_4598,N_5238);
nand U9855 (N_9855,N_5374,N_5981);
xnor U9856 (N_9856,N_6807,N_5936);
xnor U9857 (N_9857,N_7510,N_5416);
nor U9858 (N_9858,N_5172,N_4980);
nand U9859 (N_9859,N_4395,N_4406);
nor U9860 (N_9860,N_5521,N_6010);
and U9861 (N_9861,N_5494,N_7809);
and U9862 (N_9862,N_6863,N_7777);
or U9863 (N_9863,N_7472,N_6512);
and U9864 (N_9864,N_5185,N_4482);
nor U9865 (N_9865,N_7467,N_5485);
and U9866 (N_9866,N_6866,N_6762);
xnor U9867 (N_9867,N_4943,N_6997);
or U9868 (N_9868,N_5795,N_5911);
xor U9869 (N_9869,N_6511,N_4463);
xor U9870 (N_9870,N_7593,N_6132);
nor U9871 (N_9871,N_5023,N_7626);
nand U9872 (N_9872,N_6699,N_6207);
xor U9873 (N_9873,N_7338,N_5780);
and U9874 (N_9874,N_6836,N_5722);
xnor U9875 (N_9875,N_7561,N_6098);
nand U9876 (N_9876,N_5835,N_5348);
nand U9877 (N_9877,N_4790,N_5157);
xnor U9878 (N_9878,N_4820,N_6265);
nand U9879 (N_9879,N_5061,N_5592);
nand U9880 (N_9880,N_4065,N_7434);
nand U9881 (N_9881,N_6430,N_4570);
xor U9882 (N_9882,N_6326,N_6920);
and U9883 (N_9883,N_4808,N_5963);
or U9884 (N_9884,N_4268,N_6009);
or U9885 (N_9885,N_5362,N_6220);
nand U9886 (N_9886,N_5253,N_7930);
xnor U9887 (N_9887,N_5752,N_5052);
or U9888 (N_9888,N_5200,N_5764);
nor U9889 (N_9889,N_7481,N_7546);
nor U9890 (N_9890,N_7551,N_5459);
xnor U9891 (N_9891,N_5036,N_6249);
nand U9892 (N_9892,N_4008,N_4857);
and U9893 (N_9893,N_6849,N_6888);
nand U9894 (N_9894,N_6980,N_4408);
nor U9895 (N_9895,N_6450,N_4266);
nand U9896 (N_9896,N_6535,N_4727);
xor U9897 (N_9897,N_6146,N_4153);
nor U9898 (N_9898,N_5528,N_7107);
nor U9899 (N_9899,N_6675,N_7944);
xor U9900 (N_9900,N_6163,N_4168);
or U9901 (N_9901,N_4220,N_6563);
or U9902 (N_9902,N_4592,N_7433);
or U9903 (N_9903,N_7345,N_6650);
or U9904 (N_9904,N_4702,N_5236);
xnor U9905 (N_9905,N_7960,N_7864);
or U9906 (N_9906,N_4996,N_6087);
nand U9907 (N_9907,N_7473,N_7092);
nand U9908 (N_9908,N_6364,N_4080);
and U9909 (N_9909,N_5040,N_6674);
nand U9910 (N_9910,N_4596,N_7168);
and U9911 (N_9911,N_5800,N_4006);
xnor U9912 (N_9912,N_4243,N_4116);
nand U9913 (N_9913,N_4459,N_4316);
nand U9914 (N_9914,N_7629,N_7897);
xor U9915 (N_9915,N_7154,N_4387);
or U9916 (N_9916,N_5205,N_6729);
nand U9917 (N_9917,N_6276,N_6757);
and U9918 (N_9918,N_5277,N_7048);
and U9919 (N_9919,N_6887,N_4672);
or U9920 (N_9920,N_4649,N_6813);
xor U9921 (N_9921,N_5300,N_6040);
nor U9922 (N_9922,N_7538,N_4976);
or U9923 (N_9923,N_5804,N_7492);
xnor U9924 (N_9924,N_6832,N_5530);
nor U9925 (N_9925,N_5557,N_4973);
or U9926 (N_9926,N_4488,N_7276);
and U9927 (N_9927,N_6411,N_6743);
xor U9928 (N_9928,N_7987,N_7249);
nand U9929 (N_9929,N_5951,N_5420);
and U9930 (N_9930,N_4866,N_5551);
and U9931 (N_9931,N_4728,N_6572);
and U9932 (N_9932,N_5517,N_4909);
nand U9933 (N_9933,N_6031,N_5744);
nor U9934 (N_9934,N_7197,N_5334);
nand U9935 (N_9935,N_7662,N_5687);
or U9936 (N_9936,N_7226,N_5367);
or U9937 (N_9937,N_6247,N_5168);
or U9938 (N_9938,N_7000,N_6123);
nand U9939 (N_9939,N_7970,N_5846);
nand U9940 (N_9940,N_5137,N_6478);
or U9941 (N_9941,N_4906,N_5867);
xor U9942 (N_9942,N_7975,N_4577);
nand U9943 (N_9943,N_4880,N_7566);
nand U9944 (N_9944,N_5958,N_5310);
nor U9945 (N_9945,N_7263,N_7878);
and U9946 (N_9946,N_7491,N_7802);
xor U9947 (N_9947,N_6446,N_6331);
or U9948 (N_9948,N_4745,N_7049);
nand U9949 (N_9949,N_5188,N_6588);
or U9950 (N_9950,N_5037,N_4893);
xnor U9951 (N_9951,N_5343,N_6868);
or U9952 (N_9952,N_4447,N_7268);
or U9953 (N_9953,N_4121,N_6227);
or U9954 (N_9954,N_5083,N_7495);
nand U9955 (N_9955,N_4729,N_5525);
or U9956 (N_9956,N_7843,N_6528);
nand U9957 (N_9957,N_4310,N_4393);
nor U9958 (N_9958,N_5489,N_6415);
nor U9959 (N_9959,N_4583,N_6713);
and U9960 (N_9960,N_7904,N_5324);
nand U9961 (N_9961,N_5001,N_7842);
nor U9962 (N_9962,N_7164,N_5630);
xnor U9963 (N_9963,N_6124,N_7754);
and U9964 (N_9964,N_7101,N_4806);
and U9965 (N_9965,N_7293,N_4380);
or U9966 (N_9966,N_6339,N_7931);
and U9967 (N_9967,N_7449,N_4350);
and U9968 (N_9968,N_6638,N_6770);
or U9969 (N_9969,N_7251,N_4211);
xnor U9970 (N_9970,N_7452,N_4695);
nand U9971 (N_9971,N_4897,N_7222);
nor U9972 (N_9972,N_4559,N_5918);
and U9973 (N_9973,N_6200,N_4193);
nor U9974 (N_9974,N_7034,N_6745);
xnor U9975 (N_9975,N_6629,N_7665);
xnor U9976 (N_9976,N_4091,N_5400);
nor U9977 (N_9977,N_4626,N_7009);
xor U9978 (N_9978,N_6691,N_6222);
and U9979 (N_9979,N_6343,N_5295);
nor U9980 (N_9980,N_4011,N_6006);
nor U9981 (N_9981,N_4743,N_4099);
nand U9982 (N_9982,N_4462,N_4969);
xnor U9983 (N_9983,N_6407,N_6416);
nor U9984 (N_9984,N_6889,N_5982);
nand U9985 (N_9985,N_5657,N_6322);
nand U9986 (N_9986,N_5678,N_5088);
xnor U9987 (N_9987,N_4651,N_5055);
or U9988 (N_9988,N_7820,N_7181);
and U9989 (N_9989,N_6742,N_5305);
nor U9990 (N_9990,N_7343,N_6651);
nor U9991 (N_9991,N_5619,N_4325);
nor U9992 (N_9992,N_7056,N_7420);
nor U9993 (N_9993,N_6977,N_7912);
xnor U9994 (N_9994,N_7550,N_7323);
nor U9995 (N_9995,N_4810,N_5883);
nor U9996 (N_9996,N_7317,N_6787);
nor U9997 (N_9997,N_6316,N_4680);
or U9998 (N_9998,N_5754,N_7329);
nand U9999 (N_9999,N_6038,N_6058);
or U10000 (N_10000,N_7011,N_4651);
xnor U10001 (N_10001,N_7311,N_4569);
or U10002 (N_10002,N_4715,N_4939);
or U10003 (N_10003,N_6366,N_4191);
xnor U10004 (N_10004,N_5844,N_4777);
xor U10005 (N_10005,N_4634,N_6894);
xnor U10006 (N_10006,N_4253,N_4538);
nand U10007 (N_10007,N_4504,N_7681);
xor U10008 (N_10008,N_5607,N_5399);
and U10009 (N_10009,N_7893,N_5369);
nand U10010 (N_10010,N_7115,N_7516);
xnor U10011 (N_10011,N_5090,N_5691);
nor U10012 (N_10012,N_7222,N_4240);
nand U10013 (N_10013,N_4959,N_5156);
nand U10014 (N_10014,N_7329,N_4664);
and U10015 (N_10015,N_4481,N_4288);
nor U10016 (N_10016,N_6007,N_7784);
xor U10017 (N_10017,N_7024,N_4068);
and U10018 (N_10018,N_5332,N_6615);
and U10019 (N_10019,N_7502,N_4985);
and U10020 (N_10020,N_4677,N_5461);
xor U10021 (N_10021,N_5628,N_7888);
nor U10022 (N_10022,N_7117,N_5481);
and U10023 (N_10023,N_5255,N_7478);
xnor U10024 (N_10024,N_4789,N_7494);
and U10025 (N_10025,N_6586,N_4321);
xnor U10026 (N_10026,N_6401,N_7509);
or U10027 (N_10027,N_5874,N_6214);
and U10028 (N_10028,N_4123,N_4617);
nor U10029 (N_10029,N_5427,N_5806);
and U10030 (N_10030,N_7580,N_6751);
nor U10031 (N_10031,N_5015,N_5580);
nor U10032 (N_10032,N_4192,N_7214);
or U10033 (N_10033,N_7461,N_6156);
and U10034 (N_10034,N_5652,N_6643);
nand U10035 (N_10035,N_6397,N_6681);
xor U10036 (N_10036,N_6700,N_7751);
and U10037 (N_10037,N_7871,N_6933);
nor U10038 (N_10038,N_6132,N_7082);
or U10039 (N_10039,N_7927,N_5872);
nor U10040 (N_10040,N_4251,N_4932);
and U10041 (N_10041,N_4775,N_5287);
and U10042 (N_10042,N_4852,N_7307);
and U10043 (N_10043,N_4576,N_7104);
nand U10044 (N_10044,N_5909,N_7241);
nor U10045 (N_10045,N_5266,N_6202);
nand U10046 (N_10046,N_5596,N_5485);
xor U10047 (N_10047,N_4846,N_6849);
nor U10048 (N_10048,N_5923,N_5235);
xnor U10049 (N_10049,N_6774,N_4559);
and U10050 (N_10050,N_6275,N_7369);
and U10051 (N_10051,N_6570,N_6435);
xnor U10052 (N_10052,N_7799,N_6671);
nand U10053 (N_10053,N_6902,N_5648);
and U10054 (N_10054,N_7568,N_4074);
or U10055 (N_10055,N_7682,N_7434);
and U10056 (N_10056,N_5379,N_7417);
nand U10057 (N_10057,N_6010,N_7389);
nor U10058 (N_10058,N_6551,N_4406);
nand U10059 (N_10059,N_6043,N_7318);
nor U10060 (N_10060,N_5587,N_4725);
and U10061 (N_10061,N_5852,N_5654);
xor U10062 (N_10062,N_4605,N_7124);
and U10063 (N_10063,N_6728,N_4104);
or U10064 (N_10064,N_5847,N_7115);
and U10065 (N_10065,N_6463,N_4120);
and U10066 (N_10066,N_6079,N_6957);
nor U10067 (N_10067,N_4742,N_5869);
nand U10068 (N_10068,N_4660,N_5250);
nand U10069 (N_10069,N_5604,N_5749);
or U10070 (N_10070,N_4307,N_4182);
nand U10071 (N_10071,N_4863,N_7720);
nor U10072 (N_10072,N_5939,N_5232);
nor U10073 (N_10073,N_7553,N_5740);
nor U10074 (N_10074,N_7935,N_5878);
and U10075 (N_10075,N_7731,N_7047);
nor U10076 (N_10076,N_6224,N_7211);
and U10077 (N_10077,N_5788,N_5526);
xor U10078 (N_10078,N_6193,N_7773);
xor U10079 (N_10079,N_5789,N_5824);
nand U10080 (N_10080,N_6779,N_5185);
or U10081 (N_10081,N_7373,N_7986);
or U10082 (N_10082,N_5978,N_5575);
or U10083 (N_10083,N_5661,N_5550);
and U10084 (N_10084,N_5067,N_4727);
nand U10085 (N_10085,N_4662,N_4835);
and U10086 (N_10086,N_5293,N_4447);
nand U10087 (N_10087,N_4071,N_6853);
nand U10088 (N_10088,N_7264,N_5617);
and U10089 (N_10089,N_7107,N_6328);
nand U10090 (N_10090,N_7958,N_4853);
and U10091 (N_10091,N_7010,N_5984);
nor U10092 (N_10092,N_7202,N_5347);
nand U10093 (N_10093,N_4516,N_4621);
and U10094 (N_10094,N_4614,N_7574);
or U10095 (N_10095,N_7626,N_6992);
and U10096 (N_10096,N_5467,N_5058);
and U10097 (N_10097,N_5458,N_5803);
or U10098 (N_10098,N_4546,N_5029);
and U10099 (N_10099,N_5540,N_4486);
nor U10100 (N_10100,N_4175,N_7435);
or U10101 (N_10101,N_5105,N_7778);
nor U10102 (N_10102,N_5502,N_4894);
xnor U10103 (N_10103,N_6350,N_6381);
nand U10104 (N_10104,N_4848,N_4413);
nand U10105 (N_10105,N_5504,N_6574);
or U10106 (N_10106,N_6629,N_6495);
or U10107 (N_10107,N_6696,N_4936);
or U10108 (N_10108,N_7346,N_5278);
and U10109 (N_10109,N_5335,N_5084);
and U10110 (N_10110,N_4289,N_4570);
xnor U10111 (N_10111,N_7192,N_7111);
nand U10112 (N_10112,N_7403,N_6773);
xnor U10113 (N_10113,N_7016,N_4351);
or U10114 (N_10114,N_4161,N_7246);
or U10115 (N_10115,N_6992,N_4200);
nand U10116 (N_10116,N_4606,N_5368);
nand U10117 (N_10117,N_5846,N_7759);
nor U10118 (N_10118,N_5032,N_6328);
nand U10119 (N_10119,N_6899,N_4579);
and U10120 (N_10120,N_4616,N_4158);
nor U10121 (N_10121,N_4321,N_5437);
and U10122 (N_10122,N_4088,N_4385);
nor U10123 (N_10123,N_4313,N_7360);
nor U10124 (N_10124,N_7021,N_4625);
and U10125 (N_10125,N_5675,N_5466);
nor U10126 (N_10126,N_6602,N_5372);
or U10127 (N_10127,N_6653,N_7824);
or U10128 (N_10128,N_5145,N_5630);
nor U10129 (N_10129,N_5357,N_7292);
nor U10130 (N_10130,N_5162,N_5291);
or U10131 (N_10131,N_5822,N_4770);
and U10132 (N_10132,N_7307,N_5608);
xnor U10133 (N_10133,N_5809,N_6123);
nor U10134 (N_10134,N_6566,N_5375);
or U10135 (N_10135,N_4867,N_7390);
nor U10136 (N_10136,N_7775,N_4737);
or U10137 (N_10137,N_6457,N_5648);
and U10138 (N_10138,N_5142,N_5609);
and U10139 (N_10139,N_4494,N_5539);
nor U10140 (N_10140,N_7806,N_4327);
nand U10141 (N_10141,N_4610,N_6197);
or U10142 (N_10142,N_6769,N_4391);
xnor U10143 (N_10143,N_7237,N_7034);
or U10144 (N_10144,N_4567,N_6828);
xnor U10145 (N_10145,N_5399,N_5166);
or U10146 (N_10146,N_4887,N_5632);
and U10147 (N_10147,N_6160,N_6430);
and U10148 (N_10148,N_7671,N_7278);
nor U10149 (N_10149,N_4495,N_6514);
and U10150 (N_10150,N_5386,N_7914);
xor U10151 (N_10151,N_5319,N_6130);
nand U10152 (N_10152,N_7263,N_4766);
xor U10153 (N_10153,N_7349,N_6150);
xor U10154 (N_10154,N_4405,N_7147);
nor U10155 (N_10155,N_4627,N_5578);
xnor U10156 (N_10156,N_7323,N_5375);
or U10157 (N_10157,N_6839,N_4791);
or U10158 (N_10158,N_7198,N_6780);
and U10159 (N_10159,N_7260,N_5033);
nor U10160 (N_10160,N_6744,N_7962);
or U10161 (N_10161,N_5594,N_4754);
nor U10162 (N_10162,N_7627,N_7171);
xor U10163 (N_10163,N_5006,N_5862);
nand U10164 (N_10164,N_5093,N_4686);
and U10165 (N_10165,N_5519,N_4550);
nand U10166 (N_10166,N_6870,N_7771);
xor U10167 (N_10167,N_7655,N_4115);
nand U10168 (N_10168,N_5166,N_5703);
xnor U10169 (N_10169,N_7235,N_6544);
xnor U10170 (N_10170,N_7143,N_5286);
nand U10171 (N_10171,N_5408,N_5850);
or U10172 (N_10172,N_5268,N_5603);
nand U10173 (N_10173,N_6274,N_4334);
or U10174 (N_10174,N_7334,N_6013);
nand U10175 (N_10175,N_5040,N_4978);
or U10176 (N_10176,N_5813,N_7459);
nor U10177 (N_10177,N_6352,N_6562);
xor U10178 (N_10178,N_7248,N_7383);
nand U10179 (N_10179,N_4210,N_7593);
nor U10180 (N_10180,N_6612,N_6640);
and U10181 (N_10181,N_5719,N_5011);
and U10182 (N_10182,N_4676,N_4734);
and U10183 (N_10183,N_4578,N_6758);
nor U10184 (N_10184,N_4008,N_7147);
nor U10185 (N_10185,N_7781,N_4357);
xor U10186 (N_10186,N_6081,N_5509);
and U10187 (N_10187,N_7500,N_7540);
nand U10188 (N_10188,N_6448,N_5201);
nor U10189 (N_10189,N_5020,N_5550);
or U10190 (N_10190,N_4085,N_6894);
nand U10191 (N_10191,N_5953,N_7606);
and U10192 (N_10192,N_4007,N_7736);
nand U10193 (N_10193,N_4567,N_7354);
nor U10194 (N_10194,N_7962,N_4009);
nor U10195 (N_10195,N_6187,N_4006);
nand U10196 (N_10196,N_6017,N_5583);
nor U10197 (N_10197,N_5533,N_7823);
and U10198 (N_10198,N_4585,N_5954);
and U10199 (N_10199,N_5275,N_4424);
and U10200 (N_10200,N_5176,N_5112);
and U10201 (N_10201,N_5531,N_4921);
nand U10202 (N_10202,N_5310,N_7272);
and U10203 (N_10203,N_7325,N_4880);
nor U10204 (N_10204,N_4625,N_6364);
and U10205 (N_10205,N_6737,N_5158);
xnor U10206 (N_10206,N_7287,N_4481);
nand U10207 (N_10207,N_7535,N_5761);
nand U10208 (N_10208,N_5923,N_6270);
nand U10209 (N_10209,N_4933,N_7778);
nor U10210 (N_10210,N_7182,N_6662);
and U10211 (N_10211,N_7684,N_6441);
nor U10212 (N_10212,N_6938,N_4311);
and U10213 (N_10213,N_5889,N_6519);
and U10214 (N_10214,N_6636,N_5114);
xnor U10215 (N_10215,N_7176,N_6771);
nor U10216 (N_10216,N_6967,N_6460);
or U10217 (N_10217,N_6180,N_5397);
nor U10218 (N_10218,N_5255,N_4949);
and U10219 (N_10219,N_6464,N_5184);
xnor U10220 (N_10220,N_4681,N_6166);
or U10221 (N_10221,N_6080,N_7105);
or U10222 (N_10222,N_5941,N_5092);
nor U10223 (N_10223,N_7303,N_7992);
nor U10224 (N_10224,N_5117,N_5959);
nor U10225 (N_10225,N_5301,N_5158);
xnor U10226 (N_10226,N_5245,N_5573);
nor U10227 (N_10227,N_5026,N_6767);
nand U10228 (N_10228,N_6198,N_5059);
nor U10229 (N_10229,N_6084,N_6636);
or U10230 (N_10230,N_7584,N_5932);
and U10231 (N_10231,N_5056,N_4942);
nor U10232 (N_10232,N_4510,N_4241);
nor U10233 (N_10233,N_6010,N_5011);
nand U10234 (N_10234,N_6379,N_4691);
or U10235 (N_10235,N_5950,N_5322);
xnor U10236 (N_10236,N_6642,N_6271);
nor U10237 (N_10237,N_5904,N_4419);
nand U10238 (N_10238,N_4923,N_6649);
and U10239 (N_10239,N_7644,N_4846);
nand U10240 (N_10240,N_6118,N_6133);
and U10241 (N_10241,N_7473,N_6003);
nor U10242 (N_10242,N_4149,N_6599);
and U10243 (N_10243,N_6234,N_6297);
nand U10244 (N_10244,N_4741,N_5811);
nor U10245 (N_10245,N_7390,N_4975);
and U10246 (N_10246,N_6946,N_7990);
nand U10247 (N_10247,N_5553,N_5758);
and U10248 (N_10248,N_7478,N_7704);
and U10249 (N_10249,N_5007,N_7539);
or U10250 (N_10250,N_5129,N_6726);
and U10251 (N_10251,N_6964,N_4183);
xnor U10252 (N_10252,N_5729,N_4376);
or U10253 (N_10253,N_4570,N_5988);
or U10254 (N_10254,N_6433,N_6166);
nor U10255 (N_10255,N_4778,N_5196);
nand U10256 (N_10256,N_5081,N_5148);
or U10257 (N_10257,N_4541,N_4013);
and U10258 (N_10258,N_5803,N_6025);
or U10259 (N_10259,N_4964,N_5594);
nand U10260 (N_10260,N_5357,N_6519);
and U10261 (N_10261,N_6211,N_7874);
xor U10262 (N_10262,N_5754,N_6629);
xor U10263 (N_10263,N_7632,N_5252);
nand U10264 (N_10264,N_4552,N_4911);
and U10265 (N_10265,N_6616,N_6636);
nor U10266 (N_10266,N_4804,N_5353);
nand U10267 (N_10267,N_6380,N_4458);
or U10268 (N_10268,N_7720,N_7823);
xnor U10269 (N_10269,N_6357,N_5776);
xnor U10270 (N_10270,N_5395,N_6310);
xor U10271 (N_10271,N_5860,N_6137);
and U10272 (N_10272,N_7912,N_6835);
or U10273 (N_10273,N_4073,N_7559);
nor U10274 (N_10274,N_7327,N_5299);
or U10275 (N_10275,N_6683,N_4726);
nor U10276 (N_10276,N_7831,N_4068);
nand U10277 (N_10277,N_7610,N_4642);
and U10278 (N_10278,N_4600,N_7436);
or U10279 (N_10279,N_7837,N_6216);
xor U10280 (N_10280,N_6884,N_5916);
xnor U10281 (N_10281,N_5569,N_5067);
and U10282 (N_10282,N_5881,N_6222);
nor U10283 (N_10283,N_6873,N_6994);
and U10284 (N_10284,N_4516,N_6883);
nor U10285 (N_10285,N_6320,N_5230);
nand U10286 (N_10286,N_4027,N_5280);
xnor U10287 (N_10287,N_5927,N_6143);
nor U10288 (N_10288,N_7443,N_7604);
and U10289 (N_10289,N_5851,N_6635);
xor U10290 (N_10290,N_4868,N_6377);
and U10291 (N_10291,N_4074,N_6222);
and U10292 (N_10292,N_6367,N_4712);
and U10293 (N_10293,N_5638,N_7689);
and U10294 (N_10294,N_7199,N_7942);
xor U10295 (N_10295,N_5820,N_4270);
nand U10296 (N_10296,N_4816,N_7759);
nor U10297 (N_10297,N_4379,N_7594);
nor U10298 (N_10298,N_4207,N_7230);
or U10299 (N_10299,N_5180,N_5599);
nor U10300 (N_10300,N_5513,N_5766);
xor U10301 (N_10301,N_5062,N_4086);
nor U10302 (N_10302,N_7386,N_7149);
nand U10303 (N_10303,N_5340,N_7132);
xor U10304 (N_10304,N_6770,N_5902);
and U10305 (N_10305,N_6230,N_7539);
nor U10306 (N_10306,N_6296,N_6955);
and U10307 (N_10307,N_5787,N_6288);
nand U10308 (N_10308,N_7446,N_4097);
or U10309 (N_10309,N_4494,N_6221);
nor U10310 (N_10310,N_4521,N_7600);
nor U10311 (N_10311,N_6966,N_4118);
xor U10312 (N_10312,N_5719,N_5079);
nor U10313 (N_10313,N_6929,N_4068);
or U10314 (N_10314,N_4935,N_4789);
or U10315 (N_10315,N_6665,N_4566);
xnor U10316 (N_10316,N_5139,N_5617);
and U10317 (N_10317,N_7803,N_7184);
xnor U10318 (N_10318,N_4865,N_4503);
xnor U10319 (N_10319,N_5018,N_4133);
or U10320 (N_10320,N_6400,N_4969);
and U10321 (N_10321,N_7242,N_4383);
nor U10322 (N_10322,N_7051,N_7884);
xor U10323 (N_10323,N_7929,N_5879);
or U10324 (N_10324,N_7298,N_4237);
and U10325 (N_10325,N_7101,N_6293);
nand U10326 (N_10326,N_6185,N_5785);
nor U10327 (N_10327,N_5874,N_5515);
xor U10328 (N_10328,N_7104,N_5765);
or U10329 (N_10329,N_7111,N_5886);
xnor U10330 (N_10330,N_6943,N_4241);
or U10331 (N_10331,N_5143,N_6338);
and U10332 (N_10332,N_7544,N_6300);
nor U10333 (N_10333,N_5081,N_4561);
nor U10334 (N_10334,N_6554,N_4043);
xnor U10335 (N_10335,N_7722,N_4882);
xor U10336 (N_10336,N_6902,N_5413);
nand U10337 (N_10337,N_7893,N_7206);
or U10338 (N_10338,N_6070,N_5601);
or U10339 (N_10339,N_4873,N_4113);
xor U10340 (N_10340,N_6569,N_6356);
nor U10341 (N_10341,N_4945,N_6101);
or U10342 (N_10342,N_6782,N_5429);
or U10343 (N_10343,N_4612,N_6479);
nor U10344 (N_10344,N_5843,N_6560);
or U10345 (N_10345,N_7113,N_5108);
and U10346 (N_10346,N_5189,N_4044);
and U10347 (N_10347,N_6455,N_6263);
or U10348 (N_10348,N_5702,N_6821);
xnor U10349 (N_10349,N_7388,N_7773);
nor U10350 (N_10350,N_4167,N_7867);
and U10351 (N_10351,N_5219,N_7649);
and U10352 (N_10352,N_4504,N_5012);
xor U10353 (N_10353,N_6244,N_7899);
xor U10354 (N_10354,N_4365,N_4215);
or U10355 (N_10355,N_7443,N_5765);
xnor U10356 (N_10356,N_6251,N_4517);
nand U10357 (N_10357,N_5878,N_4513);
xor U10358 (N_10358,N_7944,N_6986);
nor U10359 (N_10359,N_7019,N_4081);
or U10360 (N_10360,N_7835,N_7697);
xnor U10361 (N_10361,N_5187,N_4969);
or U10362 (N_10362,N_5147,N_7247);
and U10363 (N_10363,N_4231,N_5886);
xor U10364 (N_10364,N_4626,N_4173);
xor U10365 (N_10365,N_6789,N_5078);
nor U10366 (N_10366,N_6896,N_6741);
nor U10367 (N_10367,N_4333,N_6848);
xor U10368 (N_10368,N_6771,N_4593);
nor U10369 (N_10369,N_4751,N_6390);
nand U10370 (N_10370,N_4282,N_4669);
and U10371 (N_10371,N_6170,N_7686);
or U10372 (N_10372,N_5659,N_4640);
xor U10373 (N_10373,N_6842,N_5412);
or U10374 (N_10374,N_5821,N_4768);
or U10375 (N_10375,N_5637,N_5727);
and U10376 (N_10376,N_6443,N_7639);
xor U10377 (N_10377,N_5750,N_5395);
or U10378 (N_10378,N_5185,N_6659);
nor U10379 (N_10379,N_7217,N_5271);
xnor U10380 (N_10380,N_5372,N_5428);
and U10381 (N_10381,N_5544,N_7070);
xnor U10382 (N_10382,N_6442,N_4983);
nor U10383 (N_10383,N_5434,N_5695);
nand U10384 (N_10384,N_7512,N_4551);
xor U10385 (N_10385,N_4302,N_6156);
nand U10386 (N_10386,N_5851,N_5096);
and U10387 (N_10387,N_6128,N_7022);
nor U10388 (N_10388,N_5449,N_7459);
nor U10389 (N_10389,N_7898,N_4030);
nand U10390 (N_10390,N_5269,N_4663);
nor U10391 (N_10391,N_6615,N_4102);
nor U10392 (N_10392,N_4328,N_5397);
nand U10393 (N_10393,N_4127,N_4753);
and U10394 (N_10394,N_6056,N_5106);
and U10395 (N_10395,N_6175,N_5649);
nand U10396 (N_10396,N_6294,N_6875);
xor U10397 (N_10397,N_4419,N_4289);
or U10398 (N_10398,N_6292,N_5179);
or U10399 (N_10399,N_6671,N_5626);
xor U10400 (N_10400,N_6230,N_4728);
nand U10401 (N_10401,N_4693,N_6600);
xnor U10402 (N_10402,N_4982,N_4518);
nor U10403 (N_10403,N_6617,N_4140);
and U10404 (N_10404,N_5645,N_4890);
xor U10405 (N_10405,N_4052,N_7990);
and U10406 (N_10406,N_6162,N_4167);
nand U10407 (N_10407,N_7896,N_6722);
nor U10408 (N_10408,N_6589,N_4982);
and U10409 (N_10409,N_7377,N_6413);
xnor U10410 (N_10410,N_5681,N_7104);
xor U10411 (N_10411,N_4492,N_6736);
xnor U10412 (N_10412,N_6273,N_5641);
or U10413 (N_10413,N_6769,N_6549);
nand U10414 (N_10414,N_6160,N_7605);
and U10415 (N_10415,N_4602,N_7660);
nor U10416 (N_10416,N_5539,N_7652);
nor U10417 (N_10417,N_5654,N_5903);
xnor U10418 (N_10418,N_6245,N_7553);
nor U10419 (N_10419,N_4693,N_6200);
nand U10420 (N_10420,N_5711,N_4218);
nand U10421 (N_10421,N_5755,N_7128);
nor U10422 (N_10422,N_6953,N_4287);
or U10423 (N_10423,N_6217,N_6264);
nand U10424 (N_10424,N_5776,N_5181);
nand U10425 (N_10425,N_5445,N_5877);
xnor U10426 (N_10426,N_4296,N_5205);
or U10427 (N_10427,N_4350,N_7048);
or U10428 (N_10428,N_6286,N_7374);
and U10429 (N_10429,N_4882,N_5243);
or U10430 (N_10430,N_7090,N_6507);
and U10431 (N_10431,N_4886,N_7713);
nor U10432 (N_10432,N_4143,N_7241);
or U10433 (N_10433,N_5158,N_4505);
or U10434 (N_10434,N_6605,N_7687);
or U10435 (N_10435,N_6916,N_7148);
and U10436 (N_10436,N_4874,N_4530);
xnor U10437 (N_10437,N_6560,N_6021);
nand U10438 (N_10438,N_6677,N_6126);
nand U10439 (N_10439,N_7028,N_6732);
xnor U10440 (N_10440,N_6103,N_6982);
or U10441 (N_10441,N_4189,N_4905);
nand U10442 (N_10442,N_5680,N_6182);
or U10443 (N_10443,N_4481,N_6364);
and U10444 (N_10444,N_5085,N_4230);
and U10445 (N_10445,N_4869,N_4246);
or U10446 (N_10446,N_4511,N_7639);
xnor U10447 (N_10447,N_5905,N_7856);
nand U10448 (N_10448,N_7135,N_4516);
xnor U10449 (N_10449,N_6453,N_5149);
nand U10450 (N_10450,N_7135,N_7125);
and U10451 (N_10451,N_4681,N_4542);
xnor U10452 (N_10452,N_7059,N_7021);
and U10453 (N_10453,N_6657,N_4722);
and U10454 (N_10454,N_5173,N_7723);
and U10455 (N_10455,N_5835,N_4544);
and U10456 (N_10456,N_6784,N_4321);
nand U10457 (N_10457,N_4608,N_7118);
nor U10458 (N_10458,N_7089,N_7519);
xor U10459 (N_10459,N_6693,N_4151);
or U10460 (N_10460,N_7734,N_4949);
nand U10461 (N_10461,N_4420,N_6452);
nand U10462 (N_10462,N_5873,N_4059);
nor U10463 (N_10463,N_6509,N_4045);
and U10464 (N_10464,N_6383,N_7589);
or U10465 (N_10465,N_5271,N_7442);
nand U10466 (N_10466,N_6887,N_6365);
and U10467 (N_10467,N_4697,N_4928);
and U10468 (N_10468,N_5368,N_5100);
nand U10469 (N_10469,N_4146,N_4375);
nor U10470 (N_10470,N_7403,N_5320);
nor U10471 (N_10471,N_6054,N_5308);
or U10472 (N_10472,N_5574,N_7984);
or U10473 (N_10473,N_5890,N_4667);
xnor U10474 (N_10474,N_5349,N_7596);
and U10475 (N_10475,N_6530,N_5938);
nor U10476 (N_10476,N_6992,N_6998);
and U10477 (N_10477,N_6819,N_6441);
and U10478 (N_10478,N_7670,N_6259);
and U10479 (N_10479,N_5753,N_5886);
and U10480 (N_10480,N_6293,N_4040);
xnor U10481 (N_10481,N_7857,N_6773);
or U10482 (N_10482,N_6602,N_4257);
and U10483 (N_10483,N_7759,N_6306);
or U10484 (N_10484,N_5904,N_7841);
nor U10485 (N_10485,N_4944,N_4458);
nand U10486 (N_10486,N_4517,N_6819);
and U10487 (N_10487,N_7225,N_7850);
nand U10488 (N_10488,N_6054,N_5813);
nor U10489 (N_10489,N_7590,N_6303);
or U10490 (N_10490,N_6279,N_7401);
nand U10491 (N_10491,N_6726,N_7948);
xnor U10492 (N_10492,N_5442,N_7179);
nand U10493 (N_10493,N_6052,N_4304);
or U10494 (N_10494,N_4116,N_7966);
xnor U10495 (N_10495,N_4844,N_7404);
and U10496 (N_10496,N_6450,N_6611);
nor U10497 (N_10497,N_7373,N_7010);
and U10498 (N_10498,N_6843,N_4079);
and U10499 (N_10499,N_6373,N_6628);
and U10500 (N_10500,N_7143,N_4738);
or U10501 (N_10501,N_7220,N_6726);
nand U10502 (N_10502,N_6765,N_4932);
and U10503 (N_10503,N_7072,N_7457);
nand U10504 (N_10504,N_5935,N_6024);
or U10505 (N_10505,N_7899,N_5957);
nor U10506 (N_10506,N_6187,N_7028);
nor U10507 (N_10507,N_6485,N_4967);
and U10508 (N_10508,N_4634,N_7921);
nor U10509 (N_10509,N_4601,N_6919);
xnor U10510 (N_10510,N_4002,N_6974);
and U10511 (N_10511,N_7367,N_6654);
and U10512 (N_10512,N_7599,N_6869);
xor U10513 (N_10513,N_7930,N_4105);
and U10514 (N_10514,N_4399,N_6302);
nor U10515 (N_10515,N_6302,N_4328);
and U10516 (N_10516,N_4209,N_4673);
nor U10517 (N_10517,N_5101,N_4825);
and U10518 (N_10518,N_6822,N_7289);
nand U10519 (N_10519,N_6855,N_4863);
and U10520 (N_10520,N_7433,N_5879);
nor U10521 (N_10521,N_4092,N_4067);
or U10522 (N_10522,N_6676,N_6032);
and U10523 (N_10523,N_7596,N_5611);
xnor U10524 (N_10524,N_4161,N_7830);
nand U10525 (N_10525,N_6737,N_6007);
xnor U10526 (N_10526,N_7505,N_6706);
xnor U10527 (N_10527,N_5640,N_7183);
nand U10528 (N_10528,N_7591,N_6807);
and U10529 (N_10529,N_5124,N_5911);
nor U10530 (N_10530,N_4698,N_4870);
nor U10531 (N_10531,N_6427,N_5748);
and U10532 (N_10532,N_7076,N_5959);
xor U10533 (N_10533,N_7425,N_5977);
nor U10534 (N_10534,N_5484,N_6935);
xnor U10535 (N_10535,N_7904,N_6622);
nor U10536 (N_10536,N_4006,N_6487);
nand U10537 (N_10537,N_6001,N_6064);
nor U10538 (N_10538,N_6729,N_7412);
xnor U10539 (N_10539,N_6342,N_6441);
xor U10540 (N_10540,N_7614,N_7873);
xor U10541 (N_10541,N_5814,N_7809);
nand U10542 (N_10542,N_4586,N_5559);
and U10543 (N_10543,N_7011,N_7368);
or U10544 (N_10544,N_7510,N_7037);
nand U10545 (N_10545,N_4168,N_7046);
and U10546 (N_10546,N_5079,N_4584);
or U10547 (N_10547,N_7274,N_6930);
and U10548 (N_10548,N_4949,N_6836);
xnor U10549 (N_10549,N_5697,N_7698);
nor U10550 (N_10550,N_6107,N_6252);
and U10551 (N_10551,N_5171,N_4779);
or U10552 (N_10552,N_6550,N_4668);
and U10553 (N_10553,N_4889,N_7587);
or U10554 (N_10554,N_5525,N_7128);
nand U10555 (N_10555,N_6523,N_6760);
xnor U10556 (N_10556,N_5712,N_5943);
xnor U10557 (N_10557,N_6119,N_7252);
nand U10558 (N_10558,N_5376,N_4327);
nor U10559 (N_10559,N_4606,N_5172);
nor U10560 (N_10560,N_4575,N_7447);
nor U10561 (N_10561,N_7555,N_4377);
xnor U10562 (N_10562,N_4518,N_7502);
and U10563 (N_10563,N_6105,N_6371);
and U10564 (N_10564,N_4744,N_7012);
nor U10565 (N_10565,N_7678,N_4281);
xnor U10566 (N_10566,N_6889,N_7392);
nor U10567 (N_10567,N_7097,N_7316);
xnor U10568 (N_10568,N_6363,N_7018);
or U10569 (N_10569,N_5379,N_6258);
nand U10570 (N_10570,N_7259,N_6693);
or U10571 (N_10571,N_6893,N_7473);
nor U10572 (N_10572,N_6202,N_5660);
or U10573 (N_10573,N_7546,N_7995);
nor U10574 (N_10574,N_5227,N_4070);
and U10575 (N_10575,N_4985,N_7625);
or U10576 (N_10576,N_7018,N_6458);
or U10577 (N_10577,N_5590,N_6278);
nand U10578 (N_10578,N_4912,N_5600);
xor U10579 (N_10579,N_6785,N_6682);
and U10580 (N_10580,N_4422,N_6739);
nor U10581 (N_10581,N_7014,N_7083);
xnor U10582 (N_10582,N_7060,N_5207);
nand U10583 (N_10583,N_6397,N_7622);
nor U10584 (N_10584,N_6097,N_6860);
xor U10585 (N_10585,N_6594,N_4830);
or U10586 (N_10586,N_6131,N_4475);
nor U10587 (N_10587,N_7829,N_6584);
and U10588 (N_10588,N_7319,N_6172);
or U10589 (N_10589,N_4971,N_5570);
xnor U10590 (N_10590,N_7355,N_5613);
or U10591 (N_10591,N_4418,N_5623);
nor U10592 (N_10592,N_4942,N_7237);
nand U10593 (N_10593,N_6075,N_6992);
and U10594 (N_10594,N_7394,N_7177);
nor U10595 (N_10595,N_5678,N_7797);
or U10596 (N_10596,N_6721,N_4713);
nand U10597 (N_10597,N_6725,N_7036);
nor U10598 (N_10598,N_4707,N_5306);
nor U10599 (N_10599,N_6000,N_6009);
xor U10600 (N_10600,N_4662,N_5693);
or U10601 (N_10601,N_7527,N_7320);
or U10602 (N_10602,N_4984,N_5698);
xor U10603 (N_10603,N_6624,N_5838);
and U10604 (N_10604,N_7314,N_7964);
and U10605 (N_10605,N_7859,N_6620);
and U10606 (N_10606,N_6903,N_7865);
and U10607 (N_10607,N_7575,N_4803);
or U10608 (N_10608,N_5554,N_7593);
and U10609 (N_10609,N_5954,N_6781);
xnor U10610 (N_10610,N_7499,N_4123);
and U10611 (N_10611,N_5191,N_4762);
nand U10612 (N_10612,N_5458,N_7334);
nor U10613 (N_10613,N_7004,N_5974);
and U10614 (N_10614,N_7161,N_6474);
nand U10615 (N_10615,N_6147,N_6396);
or U10616 (N_10616,N_6872,N_6686);
nand U10617 (N_10617,N_7889,N_5370);
or U10618 (N_10618,N_5418,N_6519);
and U10619 (N_10619,N_6931,N_7519);
nor U10620 (N_10620,N_6547,N_7529);
and U10621 (N_10621,N_6376,N_6940);
and U10622 (N_10622,N_4947,N_6567);
or U10623 (N_10623,N_6655,N_4129);
or U10624 (N_10624,N_7178,N_5359);
nand U10625 (N_10625,N_7038,N_5151);
nand U10626 (N_10626,N_7425,N_5281);
and U10627 (N_10627,N_6479,N_4434);
nor U10628 (N_10628,N_4688,N_5214);
nand U10629 (N_10629,N_7243,N_7029);
and U10630 (N_10630,N_5466,N_6518);
or U10631 (N_10631,N_6234,N_6637);
nand U10632 (N_10632,N_6515,N_5614);
nor U10633 (N_10633,N_7975,N_4634);
or U10634 (N_10634,N_6816,N_7674);
nor U10635 (N_10635,N_7416,N_5007);
xor U10636 (N_10636,N_4107,N_5068);
or U10637 (N_10637,N_7603,N_5306);
or U10638 (N_10638,N_4341,N_7040);
nand U10639 (N_10639,N_7190,N_6222);
or U10640 (N_10640,N_5935,N_7942);
or U10641 (N_10641,N_5730,N_4382);
or U10642 (N_10642,N_4525,N_7002);
and U10643 (N_10643,N_7518,N_6687);
or U10644 (N_10644,N_4854,N_6262);
and U10645 (N_10645,N_4362,N_7103);
xnor U10646 (N_10646,N_6353,N_7718);
or U10647 (N_10647,N_7715,N_5358);
nand U10648 (N_10648,N_4236,N_5380);
xnor U10649 (N_10649,N_5713,N_7839);
and U10650 (N_10650,N_5740,N_7443);
nand U10651 (N_10651,N_6286,N_6022);
or U10652 (N_10652,N_5974,N_6199);
and U10653 (N_10653,N_6736,N_5072);
nand U10654 (N_10654,N_7821,N_4106);
nor U10655 (N_10655,N_7839,N_6070);
or U10656 (N_10656,N_4290,N_7187);
and U10657 (N_10657,N_5473,N_5545);
and U10658 (N_10658,N_6214,N_4180);
nor U10659 (N_10659,N_4680,N_6790);
nor U10660 (N_10660,N_4364,N_4612);
xor U10661 (N_10661,N_6874,N_4825);
xnor U10662 (N_10662,N_5193,N_4971);
xnor U10663 (N_10663,N_5906,N_5453);
and U10664 (N_10664,N_7281,N_4917);
nor U10665 (N_10665,N_7240,N_7710);
xor U10666 (N_10666,N_6685,N_6465);
nor U10667 (N_10667,N_4921,N_7907);
nand U10668 (N_10668,N_4475,N_5437);
xor U10669 (N_10669,N_7604,N_5733);
nor U10670 (N_10670,N_4351,N_5775);
nand U10671 (N_10671,N_5834,N_6494);
nand U10672 (N_10672,N_4249,N_5735);
xor U10673 (N_10673,N_4462,N_7796);
nor U10674 (N_10674,N_4427,N_5379);
nand U10675 (N_10675,N_4539,N_4773);
and U10676 (N_10676,N_7518,N_5216);
or U10677 (N_10677,N_4774,N_6130);
and U10678 (N_10678,N_7674,N_4956);
and U10679 (N_10679,N_4147,N_7413);
nand U10680 (N_10680,N_7651,N_6534);
xor U10681 (N_10681,N_4679,N_5024);
or U10682 (N_10682,N_4083,N_5292);
and U10683 (N_10683,N_6521,N_7700);
or U10684 (N_10684,N_5280,N_5807);
and U10685 (N_10685,N_5213,N_7473);
nor U10686 (N_10686,N_4405,N_7958);
nand U10687 (N_10687,N_7987,N_5419);
xnor U10688 (N_10688,N_6914,N_7019);
or U10689 (N_10689,N_4095,N_4002);
and U10690 (N_10690,N_4770,N_5963);
or U10691 (N_10691,N_7677,N_6414);
or U10692 (N_10692,N_7221,N_4219);
nor U10693 (N_10693,N_6253,N_5465);
nor U10694 (N_10694,N_5766,N_5725);
and U10695 (N_10695,N_7516,N_6210);
xnor U10696 (N_10696,N_6971,N_6368);
nand U10697 (N_10697,N_5707,N_4135);
nand U10698 (N_10698,N_7685,N_4155);
and U10699 (N_10699,N_4279,N_7804);
xnor U10700 (N_10700,N_7676,N_5133);
or U10701 (N_10701,N_7136,N_7825);
nor U10702 (N_10702,N_7795,N_5500);
xnor U10703 (N_10703,N_7048,N_7154);
xnor U10704 (N_10704,N_7024,N_6333);
nor U10705 (N_10705,N_7364,N_7525);
or U10706 (N_10706,N_6429,N_4749);
or U10707 (N_10707,N_7584,N_7763);
xor U10708 (N_10708,N_5159,N_5993);
nor U10709 (N_10709,N_4327,N_6348);
xnor U10710 (N_10710,N_4544,N_7500);
nand U10711 (N_10711,N_7811,N_4620);
or U10712 (N_10712,N_4765,N_4224);
or U10713 (N_10713,N_4869,N_7289);
nor U10714 (N_10714,N_5889,N_6510);
or U10715 (N_10715,N_6693,N_4846);
xor U10716 (N_10716,N_6829,N_5033);
nand U10717 (N_10717,N_7339,N_4389);
nor U10718 (N_10718,N_6696,N_7502);
nor U10719 (N_10719,N_7049,N_4082);
or U10720 (N_10720,N_7181,N_4527);
or U10721 (N_10721,N_6228,N_4752);
xnor U10722 (N_10722,N_4489,N_5039);
nand U10723 (N_10723,N_7717,N_7525);
nor U10724 (N_10724,N_6140,N_4138);
or U10725 (N_10725,N_6934,N_7535);
and U10726 (N_10726,N_6190,N_4599);
and U10727 (N_10727,N_7879,N_5727);
xor U10728 (N_10728,N_6967,N_6309);
or U10729 (N_10729,N_5198,N_7924);
and U10730 (N_10730,N_7027,N_5764);
nand U10731 (N_10731,N_7528,N_5500);
and U10732 (N_10732,N_4702,N_7750);
and U10733 (N_10733,N_6069,N_5633);
or U10734 (N_10734,N_6729,N_5547);
and U10735 (N_10735,N_4932,N_6737);
nor U10736 (N_10736,N_5052,N_7443);
and U10737 (N_10737,N_7909,N_5417);
xnor U10738 (N_10738,N_5898,N_6075);
nor U10739 (N_10739,N_4845,N_7623);
or U10740 (N_10740,N_7611,N_7460);
nand U10741 (N_10741,N_6073,N_6982);
nand U10742 (N_10742,N_7585,N_7209);
nor U10743 (N_10743,N_7416,N_4665);
and U10744 (N_10744,N_6611,N_5827);
xor U10745 (N_10745,N_4340,N_7962);
xor U10746 (N_10746,N_5389,N_5311);
nand U10747 (N_10747,N_5154,N_5670);
nor U10748 (N_10748,N_7134,N_4495);
nand U10749 (N_10749,N_7835,N_5306);
nor U10750 (N_10750,N_5750,N_6410);
nand U10751 (N_10751,N_5847,N_7765);
nand U10752 (N_10752,N_4462,N_5758);
and U10753 (N_10753,N_6134,N_7775);
or U10754 (N_10754,N_7974,N_6934);
xnor U10755 (N_10755,N_5096,N_6518);
xnor U10756 (N_10756,N_4294,N_6771);
or U10757 (N_10757,N_4629,N_6545);
nand U10758 (N_10758,N_7313,N_6428);
nand U10759 (N_10759,N_4100,N_4800);
nor U10760 (N_10760,N_6543,N_6552);
and U10761 (N_10761,N_6056,N_5292);
and U10762 (N_10762,N_6417,N_7332);
xnor U10763 (N_10763,N_7215,N_6248);
or U10764 (N_10764,N_5929,N_6448);
nor U10765 (N_10765,N_7732,N_4912);
nand U10766 (N_10766,N_7541,N_5204);
or U10767 (N_10767,N_4308,N_6928);
or U10768 (N_10768,N_7243,N_6820);
or U10769 (N_10769,N_7920,N_5914);
nand U10770 (N_10770,N_6596,N_4596);
nor U10771 (N_10771,N_7150,N_7922);
nand U10772 (N_10772,N_5302,N_6040);
xnor U10773 (N_10773,N_6818,N_4964);
or U10774 (N_10774,N_5465,N_6316);
nor U10775 (N_10775,N_6352,N_5439);
and U10776 (N_10776,N_6312,N_4114);
nor U10777 (N_10777,N_6392,N_4248);
nor U10778 (N_10778,N_4346,N_6799);
and U10779 (N_10779,N_5389,N_4616);
xnor U10780 (N_10780,N_7523,N_5688);
and U10781 (N_10781,N_6921,N_4219);
xor U10782 (N_10782,N_6374,N_5016);
and U10783 (N_10783,N_4816,N_7373);
or U10784 (N_10784,N_5905,N_4364);
xnor U10785 (N_10785,N_5371,N_6353);
xnor U10786 (N_10786,N_7945,N_5812);
nor U10787 (N_10787,N_5393,N_7925);
xnor U10788 (N_10788,N_7319,N_5389);
xnor U10789 (N_10789,N_5828,N_7513);
and U10790 (N_10790,N_6990,N_7108);
or U10791 (N_10791,N_7505,N_6600);
or U10792 (N_10792,N_6440,N_6529);
and U10793 (N_10793,N_6635,N_4236);
or U10794 (N_10794,N_5825,N_7607);
xnor U10795 (N_10795,N_5601,N_4650);
and U10796 (N_10796,N_7334,N_7210);
or U10797 (N_10797,N_6126,N_7255);
nor U10798 (N_10798,N_7461,N_4109);
xor U10799 (N_10799,N_6700,N_7699);
or U10800 (N_10800,N_4066,N_6582);
and U10801 (N_10801,N_5094,N_6635);
xor U10802 (N_10802,N_6581,N_4113);
and U10803 (N_10803,N_4640,N_4232);
nor U10804 (N_10804,N_7205,N_4848);
xnor U10805 (N_10805,N_6343,N_6523);
xor U10806 (N_10806,N_5256,N_7922);
or U10807 (N_10807,N_6292,N_5669);
xnor U10808 (N_10808,N_5792,N_4394);
and U10809 (N_10809,N_5322,N_6154);
xor U10810 (N_10810,N_5544,N_6691);
nor U10811 (N_10811,N_4044,N_5472);
nand U10812 (N_10812,N_4038,N_5808);
and U10813 (N_10813,N_6615,N_4152);
xnor U10814 (N_10814,N_5620,N_4876);
nor U10815 (N_10815,N_7843,N_7476);
or U10816 (N_10816,N_5138,N_5396);
or U10817 (N_10817,N_6497,N_6884);
nor U10818 (N_10818,N_6570,N_6496);
nor U10819 (N_10819,N_7120,N_7099);
nor U10820 (N_10820,N_7377,N_5707);
nand U10821 (N_10821,N_5406,N_4410);
nor U10822 (N_10822,N_6455,N_7193);
xor U10823 (N_10823,N_7711,N_7332);
or U10824 (N_10824,N_6353,N_5929);
or U10825 (N_10825,N_4653,N_6901);
or U10826 (N_10826,N_7519,N_6960);
and U10827 (N_10827,N_6307,N_6880);
nand U10828 (N_10828,N_4054,N_5016);
and U10829 (N_10829,N_5125,N_4208);
nor U10830 (N_10830,N_4302,N_7521);
and U10831 (N_10831,N_7847,N_5766);
nor U10832 (N_10832,N_6058,N_7156);
xnor U10833 (N_10833,N_4405,N_5810);
and U10834 (N_10834,N_6812,N_6961);
nor U10835 (N_10835,N_5235,N_6782);
nand U10836 (N_10836,N_4673,N_6979);
and U10837 (N_10837,N_5793,N_5080);
xor U10838 (N_10838,N_5819,N_6373);
and U10839 (N_10839,N_6842,N_6756);
and U10840 (N_10840,N_4029,N_7794);
xor U10841 (N_10841,N_7346,N_4296);
or U10842 (N_10842,N_7339,N_4183);
and U10843 (N_10843,N_4744,N_6759);
and U10844 (N_10844,N_6851,N_4523);
nand U10845 (N_10845,N_7238,N_6143);
and U10846 (N_10846,N_7180,N_4280);
xnor U10847 (N_10847,N_5339,N_5821);
and U10848 (N_10848,N_4840,N_5024);
xnor U10849 (N_10849,N_6206,N_5997);
or U10850 (N_10850,N_5911,N_6679);
xnor U10851 (N_10851,N_7828,N_6369);
and U10852 (N_10852,N_5592,N_7528);
and U10853 (N_10853,N_7426,N_7471);
and U10854 (N_10854,N_7494,N_5993);
xor U10855 (N_10855,N_7762,N_7898);
xor U10856 (N_10856,N_6575,N_6347);
xnor U10857 (N_10857,N_5671,N_6261);
or U10858 (N_10858,N_6867,N_4088);
xnor U10859 (N_10859,N_4723,N_5237);
xor U10860 (N_10860,N_7155,N_5595);
or U10861 (N_10861,N_4090,N_7490);
or U10862 (N_10862,N_4514,N_5205);
and U10863 (N_10863,N_4126,N_4618);
nand U10864 (N_10864,N_5103,N_7665);
or U10865 (N_10865,N_5084,N_6912);
xnor U10866 (N_10866,N_4309,N_5924);
nand U10867 (N_10867,N_5424,N_6957);
or U10868 (N_10868,N_5851,N_6279);
and U10869 (N_10869,N_6797,N_6148);
nor U10870 (N_10870,N_6898,N_5486);
nor U10871 (N_10871,N_5997,N_4292);
or U10872 (N_10872,N_5930,N_6815);
nor U10873 (N_10873,N_5899,N_6145);
and U10874 (N_10874,N_4064,N_7438);
nor U10875 (N_10875,N_4426,N_6385);
xor U10876 (N_10876,N_7174,N_5068);
or U10877 (N_10877,N_7252,N_6822);
or U10878 (N_10878,N_5873,N_7265);
and U10879 (N_10879,N_4308,N_7549);
nand U10880 (N_10880,N_6844,N_7782);
nand U10881 (N_10881,N_6702,N_4699);
xor U10882 (N_10882,N_5631,N_5506);
nand U10883 (N_10883,N_7794,N_6865);
nor U10884 (N_10884,N_7792,N_7027);
nor U10885 (N_10885,N_5480,N_4655);
or U10886 (N_10886,N_7715,N_4656);
nand U10887 (N_10887,N_7548,N_4609);
xor U10888 (N_10888,N_5580,N_7886);
or U10889 (N_10889,N_6093,N_7162);
nand U10890 (N_10890,N_5785,N_4980);
and U10891 (N_10891,N_7791,N_7406);
or U10892 (N_10892,N_4403,N_7377);
nor U10893 (N_10893,N_4912,N_4656);
nand U10894 (N_10894,N_4173,N_5645);
xnor U10895 (N_10895,N_6640,N_4020);
nand U10896 (N_10896,N_7834,N_5820);
xnor U10897 (N_10897,N_4847,N_5492);
nor U10898 (N_10898,N_4219,N_4902);
and U10899 (N_10899,N_4149,N_5873);
nor U10900 (N_10900,N_4884,N_6609);
nand U10901 (N_10901,N_4379,N_7398);
nor U10902 (N_10902,N_7859,N_5197);
or U10903 (N_10903,N_7673,N_7605);
nor U10904 (N_10904,N_7926,N_5693);
nand U10905 (N_10905,N_4208,N_7952);
xnor U10906 (N_10906,N_4141,N_4082);
or U10907 (N_10907,N_6638,N_5344);
nand U10908 (N_10908,N_5604,N_6764);
nor U10909 (N_10909,N_7252,N_5561);
nor U10910 (N_10910,N_6348,N_4892);
or U10911 (N_10911,N_4410,N_7445);
and U10912 (N_10912,N_4437,N_7938);
nand U10913 (N_10913,N_5080,N_4747);
nand U10914 (N_10914,N_7742,N_5949);
xnor U10915 (N_10915,N_7201,N_4948);
or U10916 (N_10916,N_6261,N_4789);
or U10917 (N_10917,N_5925,N_6380);
or U10918 (N_10918,N_6788,N_7249);
and U10919 (N_10919,N_5495,N_4752);
and U10920 (N_10920,N_4573,N_7119);
nor U10921 (N_10921,N_5434,N_7374);
nand U10922 (N_10922,N_4648,N_5488);
or U10923 (N_10923,N_7161,N_5065);
and U10924 (N_10924,N_4525,N_4825);
nand U10925 (N_10925,N_5630,N_5212);
or U10926 (N_10926,N_7954,N_6718);
xor U10927 (N_10927,N_6369,N_7370);
nor U10928 (N_10928,N_6067,N_4675);
or U10929 (N_10929,N_5810,N_4917);
xnor U10930 (N_10930,N_4804,N_6440);
xor U10931 (N_10931,N_4721,N_5402);
and U10932 (N_10932,N_6291,N_7637);
nand U10933 (N_10933,N_5208,N_5478);
xnor U10934 (N_10934,N_6549,N_6066);
nand U10935 (N_10935,N_7349,N_7813);
xor U10936 (N_10936,N_4626,N_5609);
or U10937 (N_10937,N_6041,N_5272);
xnor U10938 (N_10938,N_6677,N_5916);
nand U10939 (N_10939,N_7735,N_6665);
nand U10940 (N_10940,N_7145,N_6117);
xnor U10941 (N_10941,N_6880,N_6799);
xnor U10942 (N_10942,N_4110,N_6076);
xor U10943 (N_10943,N_6833,N_7500);
xor U10944 (N_10944,N_4821,N_6765);
and U10945 (N_10945,N_5934,N_5318);
nand U10946 (N_10946,N_6987,N_7702);
nor U10947 (N_10947,N_5226,N_4327);
nand U10948 (N_10948,N_7920,N_5394);
and U10949 (N_10949,N_7280,N_4723);
xnor U10950 (N_10950,N_7437,N_6970);
and U10951 (N_10951,N_5444,N_6581);
and U10952 (N_10952,N_4714,N_7521);
nor U10953 (N_10953,N_5608,N_7998);
or U10954 (N_10954,N_5676,N_7597);
and U10955 (N_10955,N_6390,N_4478);
nor U10956 (N_10956,N_4824,N_4029);
xor U10957 (N_10957,N_5434,N_6929);
and U10958 (N_10958,N_7817,N_6324);
or U10959 (N_10959,N_6488,N_7069);
nand U10960 (N_10960,N_5345,N_7869);
or U10961 (N_10961,N_4555,N_4444);
and U10962 (N_10962,N_5313,N_5927);
nand U10963 (N_10963,N_6359,N_6707);
nor U10964 (N_10964,N_6598,N_7773);
nand U10965 (N_10965,N_5881,N_6388);
or U10966 (N_10966,N_6169,N_5525);
xnor U10967 (N_10967,N_5301,N_5040);
xor U10968 (N_10968,N_4409,N_7192);
nor U10969 (N_10969,N_4641,N_7323);
and U10970 (N_10970,N_7824,N_6215);
nor U10971 (N_10971,N_7271,N_4594);
nor U10972 (N_10972,N_7699,N_4363);
or U10973 (N_10973,N_5922,N_6686);
or U10974 (N_10974,N_6644,N_6647);
nor U10975 (N_10975,N_7768,N_6171);
nand U10976 (N_10976,N_5349,N_6708);
and U10977 (N_10977,N_6182,N_7997);
and U10978 (N_10978,N_5092,N_5231);
nor U10979 (N_10979,N_4991,N_6593);
or U10980 (N_10980,N_4147,N_6857);
and U10981 (N_10981,N_4250,N_6789);
and U10982 (N_10982,N_7593,N_5822);
or U10983 (N_10983,N_7015,N_4693);
or U10984 (N_10984,N_5697,N_4352);
nand U10985 (N_10985,N_7890,N_4005);
nand U10986 (N_10986,N_7723,N_5004);
nor U10987 (N_10987,N_6126,N_7681);
xor U10988 (N_10988,N_7021,N_4343);
and U10989 (N_10989,N_5199,N_7003);
and U10990 (N_10990,N_7507,N_7315);
or U10991 (N_10991,N_4888,N_7803);
and U10992 (N_10992,N_7533,N_4436);
or U10993 (N_10993,N_5973,N_5454);
xnor U10994 (N_10994,N_5492,N_5094);
or U10995 (N_10995,N_5215,N_6313);
nor U10996 (N_10996,N_5934,N_7773);
nor U10997 (N_10997,N_5531,N_5278);
xnor U10998 (N_10998,N_6316,N_7152);
nor U10999 (N_10999,N_7562,N_7466);
and U11000 (N_11000,N_4877,N_6937);
xnor U11001 (N_11001,N_5048,N_4095);
and U11002 (N_11002,N_4843,N_5562);
nand U11003 (N_11003,N_6063,N_4169);
xnor U11004 (N_11004,N_6057,N_7187);
or U11005 (N_11005,N_7086,N_5151);
xor U11006 (N_11006,N_6647,N_4350);
or U11007 (N_11007,N_4998,N_5026);
nand U11008 (N_11008,N_7313,N_6024);
nor U11009 (N_11009,N_4600,N_5141);
xnor U11010 (N_11010,N_6737,N_4552);
and U11011 (N_11011,N_5708,N_6064);
and U11012 (N_11012,N_6593,N_5314);
nor U11013 (N_11013,N_6616,N_5552);
and U11014 (N_11014,N_6982,N_5205);
or U11015 (N_11015,N_7128,N_4768);
and U11016 (N_11016,N_7466,N_7576);
or U11017 (N_11017,N_4673,N_5140);
nor U11018 (N_11018,N_6004,N_5372);
or U11019 (N_11019,N_7603,N_6626);
nor U11020 (N_11020,N_7194,N_6647);
xor U11021 (N_11021,N_7183,N_5660);
xor U11022 (N_11022,N_7792,N_6658);
nor U11023 (N_11023,N_4499,N_4343);
or U11024 (N_11024,N_6454,N_5859);
nand U11025 (N_11025,N_6887,N_5323);
or U11026 (N_11026,N_6132,N_4234);
and U11027 (N_11027,N_5322,N_4586);
or U11028 (N_11028,N_6176,N_6078);
and U11029 (N_11029,N_4349,N_4596);
nor U11030 (N_11030,N_6077,N_5099);
or U11031 (N_11031,N_4385,N_4701);
xor U11032 (N_11032,N_7436,N_5046);
and U11033 (N_11033,N_4358,N_7660);
and U11034 (N_11034,N_5612,N_4871);
and U11035 (N_11035,N_4912,N_5262);
xnor U11036 (N_11036,N_5337,N_7144);
nand U11037 (N_11037,N_4150,N_6349);
xnor U11038 (N_11038,N_4302,N_4229);
and U11039 (N_11039,N_7787,N_7792);
xnor U11040 (N_11040,N_6281,N_5322);
nand U11041 (N_11041,N_5557,N_6315);
nor U11042 (N_11042,N_5783,N_4409);
and U11043 (N_11043,N_7772,N_4158);
or U11044 (N_11044,N_6710,N_4480);
or U11045 (N_11045,N_5064,N_4365);
nor U11046 (N_11046,N_6270,N_5304);
xor U11047 (N_11047,N_4269,N_6047);
nand U11048 (N_11048,N_4173,N_4241);
nand U11049 (N_11049,N_5325,N_4461);
xnor U11050 (N_11050,N_5328,N_5191);
xor U11051 (N_11051,N_5061,N_4703);
and U11052 (N_11052,N_5085,N_4727);
nor U11053 (N_11053,N_6947,N_6428);
nor U11054 (N_11054,N_4293,N_5380);
or U11055 (N_11055,N_5590,N_7604);
nor U11056 (N_11056,N_6847,N_5052);
xnor U11057 (N_11057,N_4400,N_6412);
and U11058 (N_11058,N_4981,N_5093);
nand U11059 (N_11059,N_5706,N_5786);
or U11060 (N_11060,N_7380,N_7080);
and U11061 (N_11061,N_6722,N_5243);
nand U11062 (N_11062,N_4733,N_6727);
nand U11063 (N_11063,N_4578,N_4002);
or U11064 (N_11064,N_7844,N_4787);
xnor U11065 (N_11065,N_5427,N_6049);
nand U11066 (N_11066,N_5987,N_5428);
and U11067 (N_11067,N_7706,N_5150);
nand U11068 (N_11068,N_7873,N_7142);
nor U11069 (N_11069,N_7697,N_5576);
or U11070 (N_11070,N_6395,N_4127);
xor U11071 (N_11071,N_6902,N_6794);
nand U11072 (N_11072,N_5585,N_6621);
or U11073 (N_11073,N_4515,N_5411);
or U11074 (N_11074,N_6929,N_6710);
and U11075 (N_11075,N_6715,N_5888);
or U11076 (N_11076,N_4578,N_7153);
or U11077 (N_11077,N_4789,N_5223);
xnor U11078 (N_11078,N_4561,N_6468);
xor U11079 (N_11079,N_7219,N_5185);
nand U11080 (N_11080,N_7224,N_6260);
xnor U11081 (N_11081,N_7010,N_7116);
xnor U11082 (N_11082,N_6784,N_6625);
nor U11083 (N_11083,N_6839,N_5910);
nand U11084 (N_11084,N_7176,N_6152);
xnor U11085 (N_11085,N_6459,N_7404);
or U11086 (N_11086,N_5754,N_7961);
nor U11087 (N_11087,N_4520,N_6495);
and U11088 (N_11088,N_4327,N_5535);
xor U11089 (N_11089,N_7143,N_6436);
xnor U11090 (N_11090,N_4738,N_5741);
xnor U11091 (N_11091,N_6639,N_6171);
xnor U11092 (N_11092,N_5334,N_7034);
or U11093 (N_11093,N_5395,N_7524);
nand U11094 (N_11094,N_5848,N_7833);
xnor U11095 (N_11095,N_5758,N_4646);
or U11096 (N_11096,N_5637,N_6185);
nor U11097 (N_11097,N_6780,N_7018);
nand U11098 (N_11098,N_7627,N_4779);
xnor U11099 (N_11099,N_4632,N_6949);
or U11100 (N_11100,N_7905,N_7453);
or U11101 (N_11101,N_6981,N_6272);
nor U11102 (N_11102,N_5483,N_6067);
and U11103 (N_11103,N_7399,N_5606);
nor U11104 (N_11104,N_5894,N_6329);
nand U11105 (N_11105,N_7304,N_6183);
or U11106 (N_11106,N_6359,N_7570);
nand U11107 (N_11107,N_7818,N_6156);
xnor U11108 (N_11108,N_4380,N_5824);
or U11109 (N_11109,N_6292,N_6551);
nor U11110 (N_11110,N_5266,N_6451);
nand U11111 (N_11111,N_4287,N_7376);
and U11112 (N_11112,N_6976,N_7630);
nor U11113 (N_11113,N_4255,N_5449);
and U11114 (N_11114,N_4532,N_6291);
or U11115 (N_11115,N_5349,N_7479);
nor U11116 (N_11116,N_7193,N_7916);
xor U11117 (N_11117,N_4056,N_6830);
nand U11118 (N_11118,N_4601,N_5169);
nand U11119 (N_11119,N_6660,N_7861);
xnor U11120 (N_11120,N_6053,N_4684);
nand U11121 (N_11121,N_5475,N_7616);
nor U11122 (N_11122,N_4321,N_5236);
and U11123 (N_11123,N_6449,N_6330);
xnor U11124 (N_11124,N_5497,N_7190);
xnor U11125 (N_11125,N_7997,N_6031);
or U11126 (N_11126,N_6981,N_4043);
and U11127 (N_11127,N_6933,N_6076);
xnor U11128 (N_11128,N_5701,N_6256);
or U11129 (N_11129,N_5713,N_4916);
xnor U11130 (N_11130,N_5403,N_6818);
nor U11131 (N_11131,N_5761,N_6721);
nor U11132 (N_11132,N_4436,N_7653);
or U11133 (N_11133,N_4872,N_7446);
or U11134 (N_11134,N_4611,N_6436);
nor U11135 (N_11135,N_6585,N_5569);
nand U11136 (N_11136,N_7177,N_7808);
xnor U11137 (N_11137,N_7671,N_6201);
nand U11138 (N_11138,N_5300,N_7289);
xor U11139 (N_11139,N_5634,N_7663);
nand U11140 (N_11140,N_6414,N_4696);
nor U11141 (N_11141,N_4438,N_5278);
or U11142 (N_11142,N_4556,N_6642);
and U11143 (N_11143,N_4276,N_5164);
and U11144 (N_11144,N_5643,N_5774);
xor U11145 (N_11145,N_5840,N_5619);
xnor U11146 (N_11146,N_4375,N_7054);
and U11147 (N_11147,N_4149,N_7810);
xor U11148 (N_11148,N_5110,N_4670);
and U11149 (N_11149,N_6365,N_7049);
or U11150 (N_11150,N_4046,N_4940);
nor U11151 (N_11151,N_5561,N_7134);
nor U11152 (N_11152,N_6774,N_6249);
xnor U11153 (N_11153,N_6093,N_7102);
xnor U11154 (N_11154,N_5612,N_6609);
xor U11155 (N_11155,N_4801,N_5431);
nor U11156 (N_11156,N_6676,N_5904);
or U11157 (N_11157,N_7443,N_5923);
xor U11158 (N_11158,N_7666,N_4948);
or U11159 (N_11159,N_6146,N_6414);
nor U11160 (N_11160,N_6322,N_5469);
or U11161 (N_11161,N_7642,N_5352);
xnor U11162 (N_11162,N_5607,N_5237);
and U11163 (N_11163,N_5016,N_4700);
nor U11164 (N_11164,N_7510,N_7664);
nand U11165 (N_11165,N_7762,N_6857);
nand U11166 (N_11166,N_6296,N_7392);
or U11167 (N_11167,N_5203,N_5920);
or U11168 (N_11168,N_7078,N_7274);
nor U11169 (N_11169,N_7498,N_4949);
and U11170 (N_11170,N_6616,N_7293);
xor U11171 (N_11171,N_5704,N_6492);
nor U11172 (N_11172,N_6466,N_5496);
nand U11173 (N_11173,N_5831,N_6435);
nor U11174 (N_11174,N_6728,N_7970);
and U11175 (N_11175,N_5214,N_7353);
nand U11176 (N_11176,N_4889,N_6826);
xor U11177 (N_11177,N_5542,N_5048);
and U11178 (N_11178,N_6998,N_6016);
nor U11179 (N_11179,N_4662,N_5105);
xor U11180 (N_11180,N_6405,N_7420);
nand U11181 (N_11181,N_5927,N_6146);
or U11182 (N_11182,N_5962,N_6797);
xor U11183 (N_11183,N_4776,N_7748);
xnor U11184 (N_11184,N_5161,N_6177);
nor U11185 (N_11185,N_5201,N_7008);
and U11186 (N_11186,N_4752,N_6125);
xor U11187 (N_11187,N_6930,N_7265);
nand U11188 (N_11188,N_4735,N_4694);
or U11189 (N_11189,N_4106,N_6488);
nand U11190 (N_11190,N_5621,N_4163);
and U11191 (N_11191,N_5785,N_4557);
or U11192 (N_11192,N_6542,N_7581);
nand U11193 (N_11193,N_4312,N_6858);
nand U11194 (N_11194,N_5072,N_6117);
xor U11195 (N_11195,N_7352,N_5802);
or U11196 (N_11196,N_5019,N_7803);
nor U11197 (N_11197,N_5469,N_5787);
xor U11198 (N_11198,N_5689,N_4373);
or U11199 (N_11199,N_4564,N_5170);
xor U11200 (N_11200,N_7264,N_7854);
nor U11201 (N_11201,N_6533,N_4978);
nand U11202 (N_11202,N_4192,N_4485);
or U11203 (N_11203,N_5202,N_6753);
or U11204 (N_11204,N_7072,N_5336);
and U11205 (N_11205,N_5243,N_6271);
and U11206 (N_11206,N_5671,N_7881);
xnor U11207 (N_11207,N_4874,N_7461);
xnor U11208 (N_11208,N_4971,N_4868);
xnor U11209 (N_11209,N_5524,N_7853);
or U11210 (N_11210,N_5588,N_5595);
xor U11211 (N_11211,N_6035,N_5310);
and U11212 (N_11212,N_6709,N_7393);
and U11213 (N_11213,N_4927,N_7631);
xnor U11214 (N_11214,N_4821,N_5936);
xor U11215 (N_11215,N_5520,N_7570);
nor U11216 (N_11216,N_7530,N_6244);
xor U11217 (N_11217,N_7866,N_4359);
or U11218 (N_11218,N_4806,N_6196);
and U11219 (N_11219,N_7604,N_7754);
nand U11220 (N_11220,N_4911,N_4965);
xnor U11221 (N_11221,N_4243,N_4239);
nand U11222 (N_11222,N_7174,N_4802);
xor U11223 (N_11223,N_7230,N_6949);
nor U11224 (N_11224,N_7604,N_4454);
nor U11225 (N_11225,N_5233,N_6519);
nor U11226 (N_11226,N_7740,N_4042);
nor U11227 (N_11227,N_5475,N_7050);
or U11228 (N_11228,N_4044,N_4058);
nand U11229 (N_11229,N_4054,N_5628);
or U11230 (N_11230,N_7221,N_6282);
or U11231 (N_11231,N_4402,N_7173);
nor U11232 (N_11232,N_6065,N_6205);
or U11233 (N_11233,N_5906,N_6406);
nor U11234 (N_11234,N_6605,N_5851);
nand U11235 (N_11235,N_7430,N_7251);
xor U11236 (N_11236,N_7353,N_4639);
and U11237 (N_11237,N_4334,N_5431);
nor U11238 (N_11238,N_5004,N_5985);
and U11239 (N_11239,N_7046,N_5643);
xor U11240 (N_11240,N_5023,N_6654);
nand U11241 (N_11241,N_7340,N_4819);
and U11242 (N_11242,N_5149,N_5047);
nand U11243 (N_11243,N_6147,N_7635);
nand U11244 (N_11244,N_6137,N_5213);
or U11245 (N_11245,N_6511,N_7997);
nor U11246 (N_11246,N_6186,N_7202);
nor U11247 (N_11247,N_6657,N_6259);
xnor U11248 (N_11248,N_4576,N_6870);
nor U11249 (N_11249,N_5142,N_5089);
nand U11250 (N_11250,N_6488,N_7542);
and U11251 (N_11251,N_6350,N_6644);
or U11252 (N_11252,N_5785,N_4744);
or U11253 (N_11253,N_5729,N_4690);
or U11254 (N_11254,N_4953,N_7983);
nand U11255 (N_11255,N_4756,N_6882);
nand U11256 (N_11256,N_6967,N_7382);
and U11257 (N_11257,N_4191,N_7542);
nand U11258 (N_11258,N_7801,N_4814);
xnor U11259 (N_11259,N_4513,N_7842);
xor U11260 (N_11260,N_4311,N_6090);
and U11261 (N_11261,N_4338,N_4381);
nor U11262 (N_11262,N_7665,N_4258);
nand U11263 (N_11263,N_4767,N_4020);
nand U11264 (N_11264,N_6976,N_5501);
nand U11265 (N_11265,N_7670,N_5280);
xor U11266 (N_11266,N_4704,N_5960);
and U11267 (N_11267,N_6184,N_6690);
and U11268 (N_11268,N_4334,N_5509);
and U11269 (N_11269,N_4426,N_5482);
nand U11270 (N_11270,N_7819,N_7851);
nand U11271 (N_11271,N_4326,N_7532);
or U11272 (N_11272,N_7499,N_6215);
nor U11273 (N_11273,N_5631,N_7650);
nor U11274 (N_11274,N_7472,N_6345);
and U11275 (N_11275,N_5730,N_6643);
and U11276 (N_11276,N_7009,N_7409);
xnor U11277 (N_11277,N_7052,N_7501);
xor U11278 (N_11278,N_4841,N_4928);
and U11279 (N_11279,N_5255,N_4152);
xor U11280 (N_11280,N_6220,N_5085);
xnor U11281 (N_11281,N_7709,N_6034);
xor U11282 (N_11282,N_6818,N_4808);
and U11283 (N_11283,N_5739,N_5520);
nor U11284 (N_11284,N_5045,N_7299);
and U11285 (N_11285,N_7466,N_5127);
or U11286 (N_11286,N_4151,N_7112);
and U11287 (N_11287,N_7598,N_5133);
nor U11288 (N_11288,N_4059,N_5726);
nand U11289 (N_11289,N_4109,N_6994);
xor U11290 (N_11290,N_7157,N_4446);
nand U11291 (N_11291,N_7799,N_6684);
nand U11292 (N_11292,N_7060,N_6066);
nor U11293 (N_11293,N_4710,N_4183);
nand U11294 (N_11294,N_5006,N_6413);
nand U11295 (N_11295,N_7854,N_6331);
xnor U11296 (N_11296,N_6933,N_6727);
and U11297 (N_11297,N_7352,N_7492);
nor U11298 (N_11298,N_4657,N_7341);
nand U11299 (N_11299,N_4243,N_5041);
nand U11300 (N_11300,N_6763,N_6290);
or U11301 (N_11301,N_7596,N_7494);
or U11302 (N_11302,N_6181,N_4225);
nor U11303 (N_11303,N_6458,N_5252);
and U11304 (N_11304,N_6176,N_6674);
and U11305 (N_11305,N_5899,N_4395);
and U11306 (N_11306,N_6437,N_7297);
and U11307 (N_11307,N_4651,N_5394);
nor U11308 (N_11308,N_7795,N_5398);
nand U11309 (N_11309,N_7249,N_4654);
nand U11310 (N_11310,N_7021,N_5220);
and U11311 (N_11311,N_6220,N_6248);
and U11312 (N_11312,N_7236,N_5041);
or U11313 (N_11313,N_5907,N_5555);
nor U11314 (N_11314,N_5510,N_5471);
nand U11315 (N_11315,N_4062,N_4695);
xnor U11316 (N_11316,N_5255,N_6090);
and U11317 (N_11317,N_4321,N_5237);
nand U11318 (N_11318,N_4330,N_5268);
nand U11319 (N_11319,N_6822,N_4250);
or U11320 (N_11320,N_5279,N_5474);
xnor U11321 (N_11321,N_7288,N_7315);
xor U11322 (N_11322,N_7263,N_6649);
nor U11323 (N_11323,N_5612,N_4577);
nand U11324 (N_11324,N_4548,N_4655);
xor U11325 (N_11325,N_7979,N_5173);
and U11326 (N_11326,N_6665,N_4857);
or U11327 (N_11327,N_6581,N_4896);
or U11328 (N_11328,N_7964,N_7529);
and U11329 (N_11329,N_6662,N_4248);
or U11330 (N_11330,N_4764,N_7745);
and U11331 (N_11331,N_4035,N_5199);
xor U11332 (N_11332,N_4637,N_5718);
and U11333 (N_11333,N_6201,N_6558);
nand U11334 (N_11334,N_6592,N_7976);
nor U11335 (N_11335,N_7915,N_4116);
nand U11336 (N_11336,N_7196,N_4439);
and U11337 (N_11337,N_7897,N_7995);
nor U11338 (N_11338,N_7056,N_5578);
nand U11339 (N_11339,N_5270,N_4296);
nand U11340 (N_11340,N_6170,N_6772);
nor U11341 (N_11341,N_7878,N_7770);
or U11342 (N_11342,N_7927,N_7360);
nand U11343 (N_11343,N_4179,N_6907);
nor U11344 (N_11344,N_6325,N_4432);
nor U11345 (N_11345,N_5205,N_6431);
xnor U11346 (N_11346,N_4632,N_7613);
or U11347 (N_11347,N_7879,N_6721);
or U11348 (N_11348,N_6724,N_7261);
nor U11349 (N_11349,N_7489,N_7589);
nand U11350 (N_11350,N_6204,N_4075);
nor U11351 (N_11351,N_4169,N_4660);
and U11352 (N_11352,N_5305,N_6955);
nor U11353 (N_11353,N_6366,N_6743);
nand U11354 (N_11354,N_4824,N_7039);
or U11355 (N_11355,N_5469,N_7794);
and U11356 (N_11356,N_7329,N_4986);
nor U11357 (N_11357,N_6801,N_5406);
or U11358 (N_11358,N_5050,N_6301);
nand U11359 (N_11359,N_7619,N_7578);
nand U11360 (N_11360,N_7137,N_6919);
nand U11361 (N_11361,N_5189,N_5779);
xor U11362 (N_11362,N_6443,N_5612);
xor U11363 (N_11363,N_7072,N_6375);
or U11364 (N_11364,N_7532,N_4578);
nor U11365 (N_11365,N_5388,N_7047);
xor U11366 (N_11366,N_5750,N_5580);
and U11367 (N_11367,N_4416,N_4799);
nand U11368 (N_11368,N_6200,N_4035);
and U11369 (N_11369,N_4237,N_6442);
nor U11370 (N_11370,N_4901,N_5742);
or U11371 (N_11371,N_6980,N_6112);
xor U11372 (N_11372,N_6708,N_4200);
nor U11373 (N_11373,N_7926,N_6083);
and U11374 (N_11374,N_4503,N_5643);
xnor U11375 (N_11375,N_6711,N_4875);
xor U11376 (N_11376,N_6049,N_7422);
or U11377 (N_11377,N_7719,N_6739);
or U11378 (N_11378,N_5587,N_6482);
nand U11379 (N_11379,N_6442,N_4170);
nor U11380 (N_11380,N_4421,N_6291);
and U11381 (N_11381,N_4859,N_6935);
or U11382 (N_11382,N_5051,N_5602);
xor U11383 (N_11383,N_4103,N_4646);
nand U11384 (N_11384,N_6991,N_7709);
nand U11385 (N_11385,N_7677,N_6129);
xnor U11386 (N_11386,N_6944,N_5061);
nor U11387 (N_11387,N_7256,N_5080);
nor U11388 (N_11388,N_5773,N_7495);
xnor U11389 (N_11389,N_5665,N_4219);
nand U11390 (N_11390,N_5781,N_4672);
nor U11391 (N_11391,N_5334,N_7717);
nand U11392 (N_11392,N_5681,N_5366);
and U11393 (N_11393,N_6090,N_6080);
xnor U11394 (N_11394,N_7801,N_4900);
or U11395 (N_11395,N_4695,N_4057);
nor U11396 (N_11396,N_5726,N_4494);
xor U11397 (N_11397,N_4321,N_6134);
nand U11398 (N_11398,N_5141,N_6718);
and U11399 (N_11399,N_7480,N_6349);
nor U11400 (N_11400,N_6182,N_7670);
xor U11401 (N_11401,N_5626,N_6531);
and U11402 (N_11402,N_6843,N_6981);
nor U11403 (N_11403,N_6809,N_5177);
or U11404 (N_11404,N_6413,N_4925);
and U11405 (N_11405,N_6106,N_4715);
or U11406 (N_11406,N_7686,N_6744);
xor U11407 (N_11407,N_5122,N_5404);
or U11408 (N_11408,N_4907,N_5391);
nor U11409 (N_11409,N_4072,N_5401);
nand U11410 (N_11410,N_6266,N_7459);
nor U11411 (N_11411,N_5723,N_7184);
nand U11412 (N_11412,N_4376,N_7697);
and U11413 (N_11413,N_5350,N_6592);
xnor U11414 (N_11414,N_7504,N_7846);
nand U11415 (N_11415,N_7848,N_5364);
or U11416 (N_11416,N_6533,N_5243);
and U11417 (N_11417,N_6673,N_7217);
or U11418 (N_11418,N_4666,N_6319);
nor U11419 (N_11419,N_6995,N_5836);
or U11420 (N_11420,N_7929,N_7844);
nor U11421 (N_11421,N_7420,N_7566);
and U11422 (N_11422,N_6996,N_5260);
nor U11423 (N_11423,N_5227,N_4153);
nor U11424 (N_11424,N_4837,N_4611);
and U11425 (N_11425,N_4561,N_7308);
and U11426 (N_11426,N_5947,N_6034);
or U11427 (N_11427,N_4872,N_4149);
nand U11428 (N_11428,N_4070,N_4860);
xnor U11429 (N_11429,N_7037,N_4003);
xnor U11430 (N_11430,N_5493,N_5200);
nor U11431 (N_11431,N_7739,N_4051);
xor U11432 (N_11432,N_4856,N_4179);
and U11433 (N_11433,N_5011,N_5924);
xor U11434 (N_11434,N_6428,N_7940);
nor U11435 (N_11435,N_4726,N_6380);
or U11436 (N_11436,N_6471,N_7386);
xnor U11437 (N_11437,N_7810,N_7225);
nand U11438 (N_11438,N_7882,N_4471);
xor U11439 (N_11439,N_6597,N_5223);
xor U11440 (N_11440,N_5665,N_5055);
or U11441 (N_11441,N_6526,N_4311);
and U11442 (N_11442,N_6409,N_4893);
nand U11443 (N_11443,N_5096,N_7393);
and U11444 (N_11444,N_6184,N_6747);
xor U11445 (N_11445,N_7765,N_4974);
nor U11446 (N_11446,N_6675,N_5426);
nor U11447 (N_11447,N_6234,N_4774);
nor U11448 (N_11448,N_7323,N_7228);
xor U11449 (N_11449,N_5704,N_7768);
xnor U11450 (N_11450,N_7700,N_4859);
nor U11451 (N_11451,N_5785,N_4201);
nand U11452 (N_11452,N_7794,N_6665);
or U11453 (N_11453,N_7803,N_6444);
nor U11454 (N_11454,N_5546,N_6209);
or U11455 (N_11455,N_5640,N_5830);
nand U11456 (N_11456,N_5409,N_4877);
or U11457 (N_11457,N_5312,N_5180);
or U11458 (N_11458,N_5049,N_7734);
nor U11459 (N_11459,N_4046,N_5593);
or U11460 (N_11460,N_6546,N_5368);
or U11461 (N_11461,N_4525,N_7448);
nor U11462 (N_11462,N_6208,N_5067);
and U11463 (N_11463,N_6742,N_5828);
xor U11464 (N_11464,N_7826,N_6307);
nand U11465 (N_11465,N_5026,N_7349);
nor U11466 (N_11466,N_7857,N_7212);
nor U11467 (N_11467,N_7819,N_4438);
or U11468 (N_11468,N_5707,N_7949);
nor U11469 (N_11469,N_7865,N_5606);
nand U11470 (N_11470,N_4468,N_7707);
nand U11471 (N_11471,N_5067,N_4901);
nor U11472 (N_11472,N_6987,N_4246);
xnor U11473 (N_11473,N_5993,N_7017);
xnor U11474 (N_11474,N_4420,N_7068);
xnor U11475 (N_11475,N_7529,N_6710);
nor U11476 (N_11476,N_7034,N_5355);
xor U11477 (N_11477,N_7767,N_5561);
nor U11478 (N_11478,N_6943,N_6912);
nor U11479 (N_11479,N_6155,N_4733);
nand U11480 (N_11480,N_5221,N_6392);
nand U11481 (N_11481,N_5299,N_7113);
or U11482 (N_11482,N_6281,N_5336);
or U11483 (N_11483,N_6448,N_4766);
nor U11484 (N_11484,N_5122,N_6784);
or U11485 (N_11485,N_5987,N_6939);
xor U11486 (N_11486,N_4006,N_4752);
and U11487 (N_11487,N_6476,N_5344);
xnor U11488 (N_11488,N_5769,N_5020);
nand U11489 (N_11489,N_6741,N_4273);
xnor U11490 (N_11490,N_5273,N_5773);
xor U11491 (N_11491,N_5039,N_5657);
or U11492 (N_11492,N_7479,N_4935);
and U11493 (N_11493,N_6655,N_6155);
and U11494 (N_11494,N_5150,N_5974);
and U11495 (N_11495,N_4451,N_7855);
or U11496 (N_11496,N_4149,N_6717);
nand U11497 (N_11497,N_5562,N_4767);
xor U11498 (N_11498,N_7908,N_6132);
and U11499 (N_11499,N_6519,N_5626);
or U11500 (N_11500,N_4519,N_5655);
and U11501 (N_11501,N_5886,N_4186);
and U11502 (N_11502,N_6050,N_5664);
and U11503 (N_11503,N_5152,N_6692);
and U11504 (N_11504,N_7190,N_5115);
xor U11505 (N_11505,N_7440,N_6835);
nor U11506 (N_11506,N_6943,N_7444);
or U11507 (N_11507,N_6207,N_5342);
and U11508 (N_11508,N_7259,N_5340);
or U11509 (N_11509,N_7010,N_5001);
nand U11510 (N_11510,N_4879,N_6385);
xnor U11511 (N_11511,N_6033,N_7995);
and U11512 (N_11512,N_5812,N_6945);
and U11513 (N_11513,N_5432,N_5717);
nor U11514 (N_11514,N_6419,N_4402);
nor U11515 (N_11515,N_6950,N_5923);
or U11516 (N_11516,N_6667,N_6018);
nand U11517 (N_11517,N_5874,N_4684);
nand U11518 (N_11518,N_7529,N_6656);
nor U11519 (N_11519,N_7143,N_6379);
nor U11520 (N_11520,N_7165,N_6041);
nand U11521 (N_11521,N_6351,N_6178);
nor U11522 (N_11522,N_7228,N_6596);
nor U11523 (N_11523,N_7580,N_7857);
nand U11524 (N_11524,N_7151,N_6814);
nor U11525 (N_11525,N_6326,N_7847);
nand U11526 (N_11526,N_5098,N_6027);
nor U11527 (N_11527,N_4088,N_4785);
and U11528 (N_11528,N_6976,N_4142);
xor U11529 (N_11529,N_7073,N_6301);
xor U11530 (N_11530,N_7065,N_4510);
and U11531 (N_11531,N_7907,N_6005);
and U11532 (N_11532,N_6038,N_6559);
and U11533 (N_11533,N_4494,N_7507);
and U11534 (N_11534,N_4473,N_6273);
nor U11535 (N_11535,N_5317,N_4677);
nor U11536 (N_11536,N_7047,N_5083);
and U11537 (N_11537,N_6409,N_5815);
xnor U11538 (N_11538,N_6425,N_7419);
nor U11539 (N_11539,N_5337,N_4337);
nand U11540 (N_11540,N_7144,N_4209);
and U11541 (N_11541,N_6500,N_4365);
nand U11542 (N_11542,N_6471,N_5208);
nor U11543 (N_11543,N_4569,N_7162);
or U11544 (N_11544,N_7434,N_6807);
nor U11545 (N_11545,N_4709,N_7868);
or U11546 (N_11546,N_4751,N_6441);
and U11547 (N_11547,N_6472,N_6234);
nand U11548 (N_11548,N_7011,N_4833);
nand U11549 (N_11549,N_5928,N_5601);
or U11550 (N_11550,N_5649,N_7467);
and U11551 (N_11551,N_5264,N_6438);
or U11552 (N_11552,N_6295,N_6612);
nand U11553 (N_11553,N_7272,N_5583);
nor U11554 (N_11554,N_5809,N_5988);
xnor U11555 (N_11555,N_4658,N_4790);
or U11556 (N_11556,N_6479,N_5639);
nor U11557 (N_11557,N_6668,N_6655);
nor U11558 (N_11558,N_5978,N_5390);
nor U11559 (N_11559,N_4585,N_6502);
or U11560 (N_11560,N_6047,N_4107);
or U11561 (N_11561,N_4153,N_6339);
and U11562 (N_11562,N_7157,N_6763);
or U11563 (N_11563,N_7396,N_6653);
nor U11564 (N_11564,N_7335,N_7469);
or U11565 (N_11565,N_7042,N_5445);
xnor U11566 (N_11566,N_5251,N_7689);
or U11567 (N_11567,N_4954,N_5577);
nor U11568 (N_11568,N_4229,N_5290);
nor U11569 (N_11569,N_6393,N_7293);
xnor U11570 (N_11570,N_5557,N_7325);
or U11571 (N_11571,N_6692,N_6239);
xnor U11572 (N_11572,N_7269,N_6237);
or U11573 (N_11573,N_7856,N_4518);
or U11574 (N_11574,N_6583,N_5393);
xor U11575 (N_11575,N_6383,N_5357);
xor U11576 (N_11576,N_5773,N_4247);
and U11577 (N_11577,N_4879,N_5347);
or U11578 (N_11578,N_4745,N_4869);
and U11579 (N_11579,N_5004,N_5791);
nand U11580 (N_11580,N_5908,N_4594);
xnor U11581 (N_11581,N_4825,N_4617);
nand U11582 (N_11582,N_6204,N_5795);
nand U11583 (N_11583,N_5795,N_4992);
nand U11584 (N_11584,N_7229,N_7606);
xnor U11585 (N_11585,N_6636,N_7940);
or U11586 (N_11586,N_4218,N_6606);
nand U11587 (N_11587,N_4601,N_6335);
xor U11588 (N_11588,N_4248,N_7945);
nand U11589 (N_11589,N_5433,N_6244);
nand U11590 (N_11590,N_4741,N_5223);
or U11591 (N_11591,N_4768,N_5767);
or U11592 (N_11592,N_4473,N_4824);
nand U11593 (N_11593,N_5702,N_6948);
xor U11594 (N_11594,N_7596,N_7646);
and U11595 (N_11595,N_5333,N_6134);
and U11596 (N_11596,N_5243,N_7395);
and U11597 (N_11597,N_6538,N_5015);
nand U11598 (N_11598,N_6244,N_6281);
nand U11599 (N_11599,N_6034,N_5990);
xnor U11600 (N_11600,N_5220,N_4338);
nor U11601 (N_11601,N_4508,N_4468);
or U11602 (N_11602,N_4246,N_4802);
xor U11603 (N_11603,N_7248,N_7326);
nand U11604 (N_11604,N_4794,N_4710);
nor U11605 (N_11605,N_4834,N_7052);
xnor U11606 (N_11606,N_7942,N_6726);
nand U11607 (N_11607,N_4848,N_4808);
nand U11608 (N_11608,N_5495,N_4727);
or U11609 (N_11609,N_7363,N_4838);
and U11610 (N_11610,N_4287,N_7045);
nor U11611 (N_11611,N_7801,N_7148);
and U11612 (N_11612,N_5939,N_5534);
xor U11613 (N_11613,N_5278,N_4101);
xor U11614 (N_11614,N_7330,N_4497);
xnor U11615 (N_11615,N_4034,N_6552);
nand U11616 (N_11616,N_5814,N_5303);
or U11617 (N_11617,N_4853,N_4455);
xnor U11618 (N_11618,N_6025,N_5863);
and U11619 (N_11619,N_6059,N_6512);
or U11620 (N_11620,N_5569,N_4007);
xnor U11621 (N_11621,N_6243,N_6704);
nor U11622 (N_11622,N_5284,N_4581);
xnor U11623 (N_11623,N_7932,N_4519);
nand U11624 (N_11624,N_6444,N_5889);
and U11625 (N_11625,N_4909,N_6319);
xor U11626 (N_11626,N_5020,N_4575);
and U11627 (N_11627,N_7604,N_4393);
nor U11628 (N_11628,N_4049,N_5931);
xor U11629 (N_11629,N_5955,N_6977);
or U11630 (N_11630,N_6980,N_4347);
nand U11631 (N_11631,N_6784,N_4308);
xnor U11632 (N_11632,N_6694,N_5142);
xnor U11633 (N_11633,N_7219,N_5153);
or U11634 (N_11634,N_5835,N_7897);
nand U11635 (N_11635,N_7799,N_7527);
nand U11636 (N_11636,N_7362,N_7818);
or U11637 (N_11637,N_7921,N_6006);
nor U11638 (N_11638,N_5288,N_5471);
nor U11639 (N_11639,N_7175,N_5169);
nand U11640 (N_11640,N_7866,N_4980);
and U11641 (N_11641,N_4673,N_5871);
and U11642 (N_11642,N_6628,N_4976);
nor U11643 (N_11643,N_6777,N_7528);
or U11644 (N_11644,N_7876,N_6610);
nor U11645 (N_11645,N_5431,N_7132);
xnor U11646 (N_11646,N_6725,N_6240);
and U11647 (N_11647,N_4367,N_6393);
nor U11648 (N_11648,N_6939,N_7127);
and U11649 (N_11649,N_4006,N_6574);
and U11650 (N_11650,N_5313,N_4574);
and U11651 (N_11651,N_5098,N_5965);
and U11652 (N_11652,N_7251,N_4062);
or U11653 (N_11653,N_6969,N_6936);
nand U11654 (N_11654,N_4850,N_5121);
nand U11655 (N_11655,N_4747,N_5468);
xor U11656 (N_11656,N_7876,N_7433);
xor U11657 (N_11657,N_4709,N_6042);
or U11658 (N_11658,N_4900,N_6297);
nor U11659 (N_11659,N_5453,N_6253);
nand U11660 (N_11660,N_4246,N_7797);
and U11661 (N_11661,N_6139,N_6436);
nand U11662 (N_11662,N_6605,N_6017);
nor U11663 (N_11663,N_4775,N_7020);
or U11664 (N_11664,N_7618,N_6464);
nor U11665 (N_11665,N_5927,N_7084);
nand U11666 (N_11666,N_5350,N_6439);
nor U11667 (N_11667,N_5719,N_4496);
xor U11668 (N_11668,N_4699,N_4518);
nand U11669 (N_11669,N_4148,N_6923);
or U11670 (N_11670,N_7469,N_6858);
or U11671 (N_11671,N_4172,N_5072);
and U11672 (N_11672,N_4955,N_7073);
or U11673 (N_11673,N_5435,N_7779);
nand U11674 (N_11674,N_5640,N_6848);
and U11675 (N_11675,N_5457,N_6693);
xnor U11676 (N_11676,N_6138,N_6573);
or U11677 (N_11677,N_6486,N_4971);
xor U11678 (N_11678,N_5088,N_4772);
nor U11679 (N_11679,N_7098,N_7920);
xor U11680 (N_11680,N_6154,N_4537);
xor U11681 (N_11681,N_4820,N_5591);
and U11682 (N_11682,N_7433,N_5769);
nor U11683 (N_11683,N_5160,N_5861);
nor U11684 (N_11684,N_5963,N_6236);
xnor U11685 (N_11685,N_5651,N_4174);
or U11686 (N_11686,N_4164,N_7946);
nor U11687 (N_11687,N_6426,N_6528);
nor U11688 (N_11688,N_6362,N_5697);
xnor U11689 (N_11689,N_4799,N_5311);
and U11690 (N_11690,N_6791,N_6685);
xor U11691 (N_11691,N_6895,N_6175);
nor U11692 (N_11692,N_7752,N_5306);
and U11693 (N_11693,N_5910,N_6553);
nand U11694 (N_11694,N_7451,N_5707);
or U11695 (N_11695,N_6969,N_5241);
and U11696 (N_11696,N_5455,N_7492);
xnor U11697 (N_11697,N_4915,N_7833);
nand U11698 (N_11698,N_4639,N_4799);
or U11699 (N_11699,N_5134,N_6192);
or U11700 (N_11700,N_5350,N_7344);
or U11701 (N_11701,N_7426,N_6708);
nand U11702 (N_11702,N_6480,N_7919);
nand U11703 (N_11703,N_7940,N_6988);
or U11704 (N_11704,N_5345,N_6095);
and U11705 (N_11705,N_6427,N_5167);
or U11706 (N_11706,N_5944,N_7586);
and U11707 (N_11707,N_4592,N_6995);
nor U11708 (N_11708,N_7636,N_6160);
xnor U11709 (N_11709,N_7399,N_7498);
or U11710 (N_11710,N_4738,N_5031);
xnor U11711 (N_11711,N_5674,N_6551);
or U11712 (N_11712,N_5879,N_7504);
xnor U11713 (N_11713,N_7839,N_6619);
xor U11714 (N_11714,N_4965,N_4301);
and U11715 (N_11715,N_4995,N_5557);
and U11716 (N_11716,N_5527,N_6125);
or U11717 (N_11717,N_4662,N_5730);
and U11718 (N_11718,N_7963,N_6150);
nor U11719 (N_11719,N_5929,N_4379);
xor U11720 (N_11720,N_5669,N_4869);
and U11721 (N_11721,N_5583,N_5642);
nand U11722 (N_11722,N_7435,N_4285);
nand U11723 (N_11723,N_5730,N_4396);
or U11724 (N_11724,N_7026,N_5722);
nor U11725 (N_11725,N_7687,N_7911);
nand U11726 (N_11726,N_7517,N_6124);
xor U11727 (N_11727,N_6349,N_6852);
xnor U11728 (N_11728,N_4320,N_4532);
nor U11729 (N_11729,N_7475,N_6163);
nor U11730 (N_11730,N_6191,N_7971);
and U11731 (N_11731,N_5521,N_5986);
nand U11732 (N_11732,N_6526,N_6432);
xor U11733 (N_11733,N_7924,N_5568);
xnor U11734 (N_11734,N_5351,N_4233);
xnor U11735 (N_11735,N_7724,N_7050);
or U11736 (N_11736,N_5724,N_7071);
and U11737 (N_11737,N_7930,N_7422);
or U11738 (N_11738,N_4451,N_7176);
or U11739 (N_11739,N_6678,N_5256);
or U11740 (N_11740,N_6878,N_4373);
nor U11741 (N_11741,N_4523,N_4960);
and U11742 (N_11742,N_4807,N_6741);
and U11743 (N_11743,N_7296,N_6690);
nor U11744 (N_11744,N_7599,N_4269);
nand U11745 (N_11745,N_4136,N_6112);
and U11746 (N_11746,N_7581,N_4284);
nand U11747 (N_11747,N_5508,N_6108);
xor U11748 (N_11748,N_4040,N_7589);
xor U11749 (N_11749,N_6153,N_7291);
xnor U11750 (N_11750,N_5926,N_7424);
nand U11751 (N_11751,N_6329,N_7230);
or U11752 (N_11752,N_7625,N_6177);
and U11753 (N_11753,N_6421,N_5890);
xnor U11754 (N_11754,N_7969,N_4102);
nand U11755 (N_11755,N_7183,N_4293);
nor U11756 (N_11756,N_5194,N_5994);
and U11757 (N_11757,N_5729,N_7387);
or U11758 (N_11758,N_4085,N_4169);
nand U11759 (N_11759,N_7081,N_5776);
nor U11760 (N_11760,N_7831,N_4280);
and U11761 (N_11761,N_4195,N_7704);
nand U11762 (N_11762,N_4786,N_4624);
nor U11763 (N_11763,N_7896,N_4725);
nor U11764 (N_11764,N_5922,N_6286);
xnor U11765 (N_11765,N_4135,N_4151);
nor U11766 (N_11766,N_4295,N_5256);
nand U11767 (N_11767,N_5195,N_5389);
nand U11768 (N_11768,N_6459,N_7932);
and U11769 (N_11769,N_5888,N_7588);
nand U11770 (N_11770,N_7734,N_5481);
xor U11771 (N_11771,N_7157,N_5969);
nor U11772 (N_11772,N_4041,N_5895);
nand U11773 (N_11773,N_5030,N_7561);
nand U11774 (N_11774,N_5510,N_6825);
xnor U11775 (N_11775,N_5603,N_4067);
or U11776 (N_11776,N_5664,N_6687);
nand U11777 (N_11777,N_5164,N_4594);
nor U11778 (N_11778,N_6661,N_7368);
xnor U11779 (N_11779,N_6878,N_7739);
and U11780 (N_11780,N_4752,N_6795);
xnor U11781 (N_11781,N_5762,N_5907);
or U11782 (N_11782,N_7315,N_5426);
xnor U11783 (N_11783,N_7231,N_5490);
nor U11784 (N_11784,N_4924,N_6313);
nand U11785 (N_11785,N_5049,N_7489);
nor U11786 (N_11786,N_7065,N_6318);
nor U11787 (N_11787,N_5385,N_5155);
and U11788 (N_11788,N_7812,N_4811);
nor U11789 (N_11789,N_4316,N_4662);
and U11790 (N_11790,N_5867,N_5324);
and U11791 (N_11791,N_4992,N_5512);
nand U11792 (N_11792,N_6741,N_6827);
or U11793 (N_11793,N_6231,N_7485);
xor U11794 (N_11794,N_7860,N_4870);
nor U11795 (N_11795,N_6286,N_7328);
nand U11796 (N_11796,N_4544,N_4307);
nand U11797 (N_11797,N_5169,N_5034);
nor U11798 (N_11798,N_6199,N_7884);
xnor U11799 (N_11799,N_5333,N_5372);
nor U11800 (N_11800,N_6252,N_5249);
and U11801 (N_11801,N_7481,N_5246);
nor U11802 (N_11802,N_6679,N_6121);
nand U11803 (N_11803,N_7276,N_4567);
xor U11804 (N_11804,N_4338,N_5164);
xnor U11805 (N_11805,N_5543,N_7650);
or U11806 (N_11806,N_6340,N_7219);
nor U11807 (N_11807,N_6270,N_7559);
nor U11808 (N_11808,N_6712,N_7247);
xor U11809 (N_11809,N_4686,N_6890);
nor U11810 (N_11810,N_6943,N_7476);
nor U11811 (N_11811,N_7436,N_5902);
and U11812 (N_11812,N_4631,N_7994);
and U11813 (N_11813,N_5358,N_7098);
and U11814 (N_11814,N_4910,N_6463);
nor U11815 (N_11815,N_5120,N_5272);
nand U11816 (N_11816,N_6722,N_6954);
and U11817 (N_11817,N_5020,N_5997);
nor U11818 (N_11818,N_4197,N_4328);
nand U11819 (N_11819,N_7390,N_7807);
xor U11820 (N_11820,N_5450,N_7203);
nor U11821 (N_11821,N_6225,N_4352);
or U11822 (N_11822,N_7688,N_5400);
or U11823 (N_11823,N_4366,N_7454);
nor U11824 (N_11824,N_4324,N_6652);
nor U11825 (N_11825,N_5266,N_5389);
nand U11826 (N_11826,N_4445,N_6470);
xor U11827 (N_11827,N_4490,N_6193);
nor U11828 (N_11828,N_6630,N_7346);
xnor U11829 (N_11829,N_7247,N_4658);
or U11830 (N_11830,N_6797,N_4034);
xor U11831 (N_11831,N_4825,N_6135);
or U11832 (N_11832,N_5897,N_5391);
or U11833 (N_11833,N_4017,N_6686);
nand U11834 (N_11834,N_4771,N_5439);
nand U11835 (N_11835,N_5990,N_5534);
nor U11836 (N_11836,N_4114,N_5619);
nor U11837 (N_11837,N_5911,N_4110);
nor U11838 (N_11838,N_4896,N_4451);
or U11839 (N_11839,N_7908,N_7066);
and U11840 (N_11840,N_6591,N_7579);
nand U11841 (N_11841,N_6236,N_4017);
and U11842 (N_11842,N_4638,N_5632);
and U11843 (N_11843,N_7594,N_6114);
nand U11844 (N_11844,N_4696,N_7262);
nand U11845 (N_11845,N_6543,N_5949);
nor U11846 (N_11846,N_5987,N_6935);
and U11847 (N_11847,N_5902,N_7453);
nand U11848 (N_11848,N_4062,N_7088);
and U11849 (N_11849,N_5446,N_6727);
nor U11850 (N_11850,N_5581,N_5644);
nor U11851 (N_11851,N_6168,N_5532);
nand U11852 (N_11852,N_6847,N_6041);
and U11853 (N_11853,N_6966,N_6206);
nor U11854 (N_11854,N_4606,N_7370);
and U11855 (N_11855,N_5218,N_6720);
and U11856 (N_11856,N_6664,N_7626);
nor U11857 (N_11857,N_4261,N_6348);
and U11858 (N_11858,N_7796,N_7970);
and U11859 (N_11859,N_7453,N_7625);
nor U11860 (N_11860,N_5810,N_7824);
or U11861 (N_11861,N_4133,N_7655);
nor U11862 (N_11862,N_6131,N_5355);
nor U11863 (N_11863,N_5086,N_7643);
nor U11864 (N_11864,N_5222,N_7829);
and U11865 (N_11865,N_4060,N_4031);
and U11866 (N_11866,N_6582,N_4750);
nor U11867 (N_11867,N_7323,N_7721);
nand U11868 (N_11868,N_6741,N_5969);
or U11869 (N_11869,N_4980,N_7554);
nand U11870 (N_11870,N_7943,N_7140);
nand U11871 (N_11871,N_6852,N_6533);
xor U11872 (N_11872,N_5144,N_5117);
nor U11873 (N_11873,N_4415,N_6707);
and U11874 (N_11874,N_7372,N_7227);
and U11875 (N_11875,N_7253,N_7513);
or U11876 (N_11876,N_7552,N_5718);
and U11877 (N_11877,N_6309,N_6038);
xor U11878 (N_11878,N_5545,N_7549);
and U11879 (N_11879,N_6405,N_4272);
nand U11880 (N_11880,N_6379,N_5238);
xor U11881 (N_11881,N_4985,N_7356);
or U11882 (N_11882,N_7703,N_7589);
nand U11883 (N_11883,N_7315,N_7506);
and U11884 (N_11884,N_6621,N_4071);
nand U11885 (N_11885,N_5382,N_5976);
or U11886 (N_11886,N_6639,N_7292);
or U11887 (N_11887,N_7421,N_5591);
xor U11888 (N_11888,N_7472,N_7232);
xor U11889 (N_11889,N_5387,N_7283);
and U11890 (N_11890,N_7164,N_4577);
nand U11891 (N_11891,N_4325,N_7121);
nor U11892 (N_11892,N_7923,N_6026);
nand U11893 (N_11893,N_6944,N_5890);
or U11894 (N_11894,N_7028,N_6382);
and U11895 (N_11895,N_4482,N_7149);
or U11896 (N_11896,N_6279,N_7926);
nor U11897 (N_11897,N_5182,N_5239);
xnor U11898 (N_11898,N_7007,N_7454);
and U11899 (N_11899,N_7451,N_6270);
nand U11900 (N_11900,N_5951,N_7003);
nand U11901 (N_11901,N_7479,N_4881);
and U11902 (N_11902,N_6345,N_6067);
or U11903 (N_11903,N_5779,N_4889);
xnor U11904 (N_11904,N_6774,N_5935);
or U11905 (N_11905,N_5540,N_4254);
or U11906 (N_11906,N_7830,N_6633);
or U11907 (N_11907,N_6767,N_6476);
or U11908 (N_11908,N_7601,N_6036);
nand U11909 (N_11909,N_7995,N_4375);
nand U11910 (N_11910,N_6355,N_6088);
nor U11911 (N_11911,N_5888,N_5589);
xor U11912 (N_11912,N_6499,N_5415);
and U11913 (N_11913,N_6722,N_5856);
nor U11914 (N_11914,N_5549,N_5059);
and U11915 (N_11915,N_4421,N_7269);
nand U11916 (N_11916,N_4213,N_6843);
or U11917 (N_11917,N_5306,N_4075);
and U11918 (N_11918,N_7371,N_6656);
xor U11919 (N_11919,N_4149,N_5966);
nand U11920 (N_11920,N_5810,N_6723);
or U11921 (N_11921,N_6053,N_6816);
nor U11922 (N_11922,N_7026,N_4231);
xnor U11923 (N_11923,N_7967,N_4413);
nor U11924 (N_11924,N_5535,N_7859);
nor U11925 (N_11925,N_5734,N_5392);
xor U11926 (N_11926,N_4388,N_5190);
nor U11927 (N_11927,N_6160,N_7101);
or U11928 (N_11928,N_5277,N_6759);
nor U11929 (N_11929,N_5591,N_7932);
xor U11930 (N_11930,N_5924,N_6254);
nand U11931 (N_11931,N_7439,N_7513);
nor U11932 (N_11932,N_5297,N_4974);
xor U11933 (N_11933,N_7780,N_6623);
and U11934 (N_11934,N_6679,N_5687);
or U11935 (N_11935,N_4344,N_4924);
or U11936 (N_11936,N_7152,N_6909);
and U11937 (N_11937,N_7084,N_4169);
nor U11938 (N_11938,N_7721,N_6203);
or U11939 (N_11939,N_6968,N_7547);
or U11940 (N_11940,N_5595,N_7986);
nand U11941 (N_11941,N_6164,N_4390);
nor U11942 (N_11942,N_7307,N_7534);
or U11943 (N_11943,N_5067,N_7101);
xnor U11944 (N_11944,N_6122,N_7386);
and U11945 (N_11945,N_5175,N_6585);
nor U11946 (N_11946,N_5626,N_7942);
xor U11947 (N_11947,N_4096,N_5737);
nand U11948 (N_11948,N_7335,N_6704);
nor U11949 (N_11949,N_4416,N_6319);
or U11950 (N_11950,N_4787,N_7483);
nand U11951 (N_11951,N_5892,N_7893);
and U11952 (N_11952,N_6165,N_7448);
nand U11953 (N_11953,N_4271,N_7536);
and U11954 (N_11954,N_4962,N_4058);
and U11955 (N_11955,N_6127,N_7672);
xor U11956 (N_11956,N_4458,N_7952);
or U11957 (N_11957,N_5494,N_7477);
xnor U11958 (N_11958,N_7128,N_5193);
nand U11959 (N_11959,N_5589,N_7401);
or U11960 (N_11960,N_4501,N_5938);
and U11961 (N_11961,N_6838,N_6464);
xnor U11962 (N_11962,N_7532,N_7854);
nor U11963 (N_11963,N_7805,N_4429);
xnor U11964 (N_11964,N_4580,N_6058);
and U11965 (N_11965,N_6685,N_6933);
nand U11966 (N_11966,N_7769,N_7512);
and U11967 (N_11967,N_7878,N_5759);
xor U11968 (N_11968,N_7381,N_7648);
nor U11969 (N_11969,N_4556,N_7516);
nand U11970 (N_11970,N_4808,N_6807);
or U11971 (N_11971,N_7500,N_6042);
xnor U11972 (N_11972,N_7852,N_7591);
or U11973 (N_11973,N_5010,N_5471);
xnor U11974 (N_11974,N_6289,N_6029);
and U11975 (N_11975,N_6846,N_4167);
nor U11976 (N_11976,N_4103,N_7688);
nor U11977 (N_11977,N_5519,N_4861);
nor U11978 (N_11978,N_6755,N_7493);
nor U11979 (N_11979,N_4010,N_6738);
xor U11980 (N_11980,N_4114,N_4934);
nor U11981 (N_11981,N_7292,N_6453);
or U11982 (N_11982,N_4275,N_7929);
nand U11983 (N_11983,N_4122,N_7239);
xor U11984 (N_11984,N_7962,N_6903);
or U11985 (N_11985,N_7271,N_7705);
nand U11986 (N_11986,N_5856,N_4119);
xnor U11987 (N_11987,N_5196,N_4676);
or U11988 (N_11988,N_4235,N_7658);
nand U11989 (N_11989,N_5464,N_6736);
nand U11990 (N_11990,N_6350,N_5027);
nand U11991 (N_11991,N_6950,N_6229);
and U11992 (N_11992,N_5709,N_4352);
xnor U11993 (N_11993,N_6935,N_5805);
nor U11994 (N_11994,N_7553,N_4495);
or U11995 (N_11995,N_4377,N_5193);
or U11996 (N_11996,N_7197,N_7223);
nor U11997 (N_11997,N_5984,N_6030);
nor U11998 (N_11998,N_4181,N_4897);
xnor U11999 (N_11999,N_6355,N_7969);
and U12000 (N_12000,N_9582,N_10589);
nand U12001 (N_12001,N_10201,N_8499);
nand U12002 (N_12002,N_9057,N_10274);
and U12003 (N_12003,N_11070,N_8032);
or U12004 (N_12004,N_8736,N_10971);
or U12005 (N_12005,N_9293,N_10503);
nor U12006 (N_12006,N_10179,N_11547);
and U12007 (N_12007,N_9774,N_10535);
nand U12008 (N_12008,N_9426,N_11530);
and U12009 (N_12009,N_10929,N_11678);
xnor U12010 (N_12010,N_10273,N_10432);
xor U12011 (N_12011,N_8903,N_11654);
nand U12012 (N_12012,N_8922,N_9607);
and U12013 (N_12013,N_10985,N_11603);
nand U12014 (N_12014,N_11364,N_11178);
and U12015 (N_12015,N_8967,N_8068);
xnor U12016 (N_12016,N_9417,N_11935);
xor U12017 (N_12017,N_8474,N_11323);
and U12018 (N_12018,N_11766,N_8777);
or U12019 (N_12019,N_10318,N_11642);
nand U12020 (N_12020,N_10964,N_9710);
or U12021 (N_12021,N_10252,N_11708);
or U12022 (N_12022,N_11199,N_10487);
nor U12023 (N_12023,N_8046,N_11007);
nand U12024 (N_12024,N_9126,N_10673);
or U12025 (N_12025,N_8061,N_9020);
nor U12026 (N_12026,N_8540,N_9427);
xnor U12027 (N_12027,N_10948,N_9890);
or U12028 (N_12028,N_8188,N_9198);
and U12029 (N_12029,N_11454,N_11952);
and U12030 (N_12030,N_10039,N_10213);
xnor U12031 (N_12031,N_10987,N_10307);
and U12032 (N_12032,N_8109,N_10603);
nand U12033 (N_12033,N_10458,N_8975);
or U12034 (N_12034,N_9546,N_9495);
nor U12035 (N_12035,N_9393,N_9153);
or U12036 (N_12036,N_10263,N_8079);
and U12037 (N_12037,N_8837,N_10141);
nor U12038 (N_12038,N_8521,N_9828);
and U12039 (N_12039,N_11962,N_11676);
nor U12040 (N_12040,N_10925,N_11153);
nor U12041 (N_12041,N_9610,N_11857);
nand U12042 (N_12042,N_11757,N_10214);
xor U12043 (N_12043,N_11033,N_8180);
xnor U12044 (N_12044,N_10643,N_11889);
or U12045 (N_12045,N_11414,N_11542);
xnor U12046 (N_12046,N_11856,N_10581);
nor U12047 (N_12047,N_11733,N_11800);
and U12048 (N_12048,N_10664,N_9056);
or U12049 (N_12049,N_11407,N_8944);
xor U12050 (N_12050,N_10628,N_8843);
nor U12051 (N_12051,N_11356,N_11329);
or U12052 (N_12052,N_9931,N_9058);
nor U12053 (N_12053,N_10712,N_10192);
nand U12054 (N_12054,N_9471,N_8639);
or U12055 (N_12055,N_8411,N_9540);
nor U12056 (N_12056,N_8451,N_10669);
or U12057 (N_12057,N_10129,N_8774);
nand U12058 (N_12058,N_10558,N_11671);
and U12059 (N_12059,N_8120,N_8013);
nand U12060 (N_12060,N_8164,N_10960);
or U12061 (N_12061,N_10716,N_9306);
nand U12062 (N_12062,N_9305,N_10498);
and U12063 (N_12063,N_11279,N_9978);
xor U12064 (N_12064,N_10687,N_9913);
and U12065 (N_12065,N_9968,N_11629);
nand U12066 (N_12066,N_11833,N_11220);
nand U12067 (N_12067,N_11493,N_10209);
xnor U12068 (N_12068,N_9278,N_9115);
nor U12069 (N_12069,N_9700,N_8218);
xor U12070 (N_12070,N_11755,N_8692);
nor U12071 (N_12071,N_10494,N_9037);
xor U12072 (N_12072,N_11382,N_9855);
nand U12073 (N_12073,N_8191,N_8492);
xnor U12074 (N_12074,N_10021,N_9672);
and U12075 (N_12075,N_11675,N_8604);
xor U12076 (N_12076,N_8089,N_11525);
nor U12077 (N_12077,N_11781,N_11036);
and U12078 (N_12078,N_9706,N_11185);
or U12079 (N_12079,N_11840,N_9491);
xor U12080 (N_12080,N_10732,N_11752);
or U12081 (N_12081,N_10738,N_11680);
or U12082 (N_12082,N_9813,N_10937);
and U12083 (N_12083,N_11424,N_9838);
and U12084 (N_12084,N_8189,N_9209);
nor U12085 (N_12085,N_8948,N_9681);
or U12086 (N_12086,N_10623,N_10060);
xnor U12087 (N_12087,N_8877,N_8569);
and U12088 (N_12088,N_10227,N_11221);
xor U12089 (N_12089,N_8332,N_11836);
nand U12090 (N_12090,N_9340,N_9212);
or U12091 (N_12091,N_9104,N_11148);
xnor U12092 (N_12092,N_8809,N_10768);
and U12093 (N_12093,N_9485,N_11795);
xnor U12094 (N_12094,N_9050,N_8848);
nand U12095 (N_12095,N_8437,N_11059);
nor U12096 (N_12096,N_8129,N_11050);
nor U12097 (N_12097,N_9390,N_8594);
and U12098 (N_12098,N_8351,N_8452);
or U12099 (N_12099,N_8512,N_8830);
nand U12100 (N_12100,N_11235,N_8005);
or U12101 (N_12101,N_8582,N_8573);
and U12102 (N_12102,N_11282,N_9450);
xnor U12103 (N_12103,N_11812,N_8516);
xor U12104 (N_12104,N_9785,N_11581);
xor U12105 (N_12105,N_8909,N_10430);
nor U12106 (N_12106,N_9523,N_10470);
and U12107 (N_12107,N_8447,N_11958);
and U12108 (N_12108,N_8530,N_11014);
nor U12109 (N_12109,N_10478,N_8235);
nor U12110 (N_12110,N_10629,N_9778);
xor U12111 (N_12111,N_10812,N_9142);
and U12112 (N_12112,N_11331,N_8298);
nand U12113 (N_12113,N_9704,N_10115);
nor U12114 (N_12114,N_8140,N_8552);
and U12115 (N_12115,N_11989,N_11154);
xor U12116 (N_12116,N_8181,N_8767);
or U12117 (N_12117,N_9203,N_10747);
nand U12118 (N_12118,N_10617,N_11947);
nor U12119 (N_12119,N_10431,N_9708);
nor U12120 (N_12120,N_9239,N_8864);
xnor U12121 (N_12121,N_11257,N_11724);
nand U12122 (N_12122,N_8003,N_10809);
nand U12123 (N_12123,N_11203,N_10187);
or U12124 (N_12124,N_10889,N_11880);
xor U12125 (N_12125,N_9157,N_11817);
and U12126 (N_12126,N_9361,N_8222);
xnor U12127 (N_12127,N_8456,N_10649);
xor U12128 (N_12128,N_10236,N_11118);
nor U12129 (N_12129,N_10941,N_10750);
nand U12130 (N_12130,N_9762,N_10407);
or U12131 (N_12131,N_10059,N_9698);
and U12132 (N_12132,N_10616,N_8566);
nand U12133 (N_12133,N_10707,N_8868);
xor U12134 (N_12134,N_9612,N_10098);
nand U12135 (N_12135,N_9385,N_11866);
or U12136 (N_12136,N_8312,N_8099);
nand U12137 (N_12137,N_10406,N_10901);
xnor U12138 (N_12138,N_8067,N_10740);
nand U12139 (N_12139,N_9812,N_10534);
xor U12140 (N_12140,N_8800,N_10438);
and U12141 (N_12141,N_11919,N_8750);
and U12142 (N_12142,N_8102,N_8136);
and U12143 (N_12143,N_8740,N_9516);
or U12144 (N_12144,N_10927,N_9645);
nor U12145 (N_12145,N_8647,N_11893);
nor U12146 (N_12146,N_11596,N_10315);
or U12147 (N_12147,N_9942,N_9566);
and U12148 (N_12148,N_11689,N_11379);
xor U12149 (N_12149,N_11318,N_9353);
or U12150 (N_12150,N_9169,N_11630);
nor U12151 (N_12151,N_11735,N_8618);
and U12152 (N_12152,N_9827,N_8953);
nor U12153 (N_12153,N_8963,N_11869);
and U12154 (N_12154,N_10167,N_11151);
xor U12155 (N_12155,N_11835,N_11745);
nor U12156 (N_12156,N_10600,N_10878);
or U12157 (N_12157,N_11219,N_8572);
nor U12158 (N_12158,N_10570,N_11823);
nor U12159 (N_12159,N_8232,N_10797);
nand U12160 (N_12160,N_10342,N_9188);
and U12161 (N_12161,N_8522,N_10101);
or U12162 (N_12162,N_10297,N_10011);
xor U12163 (N_12163,N_10147,N_8314);
and U12164 (N_12164,N_8434,N_9506);
and U12165 (N_12165,N_8444,N_11479);
nand U12166 (N_12166,N_8589,N_10991);
nand U12167 (N_12167,N_10977,N_10198);
nor U12168 (N_12168,N_9884,N_11861);
nor U12169 (N_12169,N_10823,N_9752);
xor U12170 (N_12170,N_11428,N_8477);
xnor U12171 (N_12171,N_8996,N_11000);
nand U12172 (N_12172,N_8838,N_11569);
or U12173 (N_12173,N_11066,N_8168);
nor U12174 (N_12174,N_10696,N_11432);
and U12175 (N_12175,N_11172,N_11419);
nand U12176 (N_12176,N_9837,N_8699);
or U12177 (N_12177,N_11370,N_9842);
nand U12178 (N_12178,N_9928,N_9027);
nor U12179 (N_12179,N_10266,N_8386);
or U12180 (N_12180,N_11820,N_10351);
xor U12181 (N_12181,N_10247,N_10408);
and U12182 (N_12182,N_9834,N_8727);
nor U12183 (N_12183,N_10818,N_11631);
and U12184 (N_12184,N_10569,N_9419);
xnor U12185 (N_12185,N_10719,N_9382);
nand U12186 (N_12186,N_9034,N_9745);
nor U12187 (N_12187,N_11982,N_10680);
nor U12188 (N_12188,N_11274,N_9897);
nand U12189 (N_12189,N_11799,N_8449);
and U12190 (N_12190,N_10435,N_9699);
nand U12191 (N_12191,N_9051,N_9605);
xnor U12192 (N_12192,N_8599,N_9149);
nand U12193 (N_12193,N_10068,N_8588);
or U12194 (N_12194,N_9729,N_9052);
nor U12195 (N_12195,N_8607,N_10757);
nor U12196 (N_12196,N_10362,N_11934);
xor U12197 (N_12197,N_11384,N_8501);
nor U12198 (N_12198,N_8743,N_11200);
nor U12199 (N_12199,N_8593,N_11848);
or U12200 (N_12200,N_10420,N_11402);
nor U12201 (N_12201,N_8128,N_9483);
nand U12202 (N_12202,N_9448,N_10921);
nor U12203 (N_12203,N_9476,N_11162);
nor U12204 (N_12204,N_10316,N_8725);
nor U12205 (N_12205,N_9323,N_8491);
nor U12206 (N_12206,N_11413,N_11195);
xor U12207 (N_12207,N_10820,N_10134);
nor U12208 (N_12208,N_9467,N_11386);
nor U12209 (N_12209,N_8342,N_8713);
or U12210 (N_12210,N_8598,N_9243);
or U12211 (N_12211,N_9696,N_8755);
xnor U12212 (N_12212,N_8721,N_10848);
nand U12213 (N_12213,N_10286,N_9287);
nor U12214 (N_12214,N_9286,N_8832);
xnor U12215 (N_12215,N_10621,N_10978);
nor U12216 (N_12216,N_10546,N_11756);
and U12217 (N_12217,N_9727,N_11863);
or U12218 (N_12218,N_10436,N_9422);
xor U12219 (N_12219,N_8786,N_9215);
and U12220 (N_12220,N_9715,N_8545);
xnor U12221 (N_12221,N_9714,N_11886);
nand U12222 (N_12222,N_8148,N_10804);
xnor U12223 (N_12223,N_11742,N_8293);
nor U12224 (N_12224,N_8428,N_11957);
or U12225 (N_12225,N_8365,N_9045);
nor U12226 (N_12226,N_9983,N_10374);
nand U12227 (N_12227,N_9849,N_11288);
nor U12228 (N_12228,N_8372,N_8949);
or U12229 (N_12229,N_9197,N_10332);
and U12230 (N_12230,N_11316,N_10468);
or U12231 (N_12231,N_9632,N_11684);
and U12232 (N_12232,N_8753,N_11566);
nand U12233 (N_12233,N_8898,N_11518);
nor U12234 (N_12234,N_9617,N_9141);
nor U12235 (N_12235,N_9830,N_11457);
or U12236 (N_12236,N_8419,N_9924);
nand U12237 (N_12237,N_10653,N_9761);
xnor U12238 (N_12238,N_8022,N_9481);
and U12239 (N_12239,N_10940,N_11262);
or U12240 (N_12240,N_11707,N_10841);
xor U12241 (N_12241,N_8883,N_8813);
nand U12242 (N_12242,N_9581,N_9132);
nor U12243 (N_12243,N_11739,N_8283);
and U12244 (N_12244,N_8033,N_11056);
or U12245 (N_12245,N_10996,N_8664);
or U12246 (N_12246,N_11805,N_11746);
nand U12247 (N_12247,N_9906,N_8870);
and U12248 (N_12248,N_10839,N_8684);
and U12249 (N_12249,N_8849,N_8973);
xor U12250 (N_12250,N_11074,N_11335);
xnor U12251 (N_12251,N_9967,N_10989);
nand U12252 (N_12252,N_11607,N_8336);
or U12253 (N_12253,N_11468,N_8887);
xnor U12254 (N_12254,N_11488,N_8968);
or U12255 (N_12255,N_9507,N_8483);
nand U12256 (N_12256,N_10052,N_10481);
nand U12257 (N_12257,N_10635,N_8073);
nand U12258 (N_12258,N_10693,N_8009);
nor U12259 (N_12259,N_8264,N_9786);
and U12260 (N_12260,N_11830,N_10763);
or U12261 (N_12261,N_9613,N_9357);
nor U12262 (N_12262,N_8867,N_9086);
nor U12263 (N_12263,N_11346,N_9438);
and U12264 (N_12264,N_8673,N_10658);
nand U12265 (N_12265,N_8912,N_8654);
xnor U12266 (N_12266,N_8791,N_10027);
and U12267 (N_12267,N_11878,N_9131);
nand U12268 (N_12268,N_9244,N_9962);
xor U12269 (N_12269,N_9437,N_9539);
xnor U12270 (N_12270,N_11164,N_10099);
nand U12271 (N_12271,N_9087,N_9098);
xor U12272 (N_12272,N_8651,N_9735);
xor U12273 (N_12273,N_9042,N_11946);
xor U12274 (N_12274,N_9811,N_9847);
nor U12275 (N_12275,N_10178,N_8693);
xor U12276 (N_12276,N_9737,N_11481);
and U12277 (N_12277,N_9592,N_10887);
nand U12278 (N_12278,N_10353,N_11433);
and U12279 (N_12279,N_9380,N_8108);
xor U12280 (N_12280,N_10279,N_8702);
and U12281 (N_12281,N_10338,N_10632);
nor U12282 (N_12282,N_9848,N_10473);
or U12283 (N_12283,N_10152,N_9776);
or U12284 (N_12284,N_10114,N_8507);
nand U12285 (N_12285,N_11804,N_10303);
xnor U12286 (N_12286,N_10942,N_8083);
xnor U12287 (N_12287,N_11146,N_10913);
and U12288 (N_12288,N_10548,N_10419);
nand U12289 (N_12289,N_9604,N_9492);
nand U12290 (N_12290,N_8257,N_11251);
and U12291 (N_12291,N_9109,N_8010);
nand U12292 (N_12292,N_11467,N_10947);
nor U12293 (N_12293,N_9334,N_11669);
xnor U12294 (N_12294,N_10410,N_8862);
xor U12295 (N_12295,N_9479,N_11324);
and U12296 (N_12296,N_10495,N_11234);
nor U12297 (N_12297,N_9145,N_10933);
xnor U12298 (N_12298,N_8955,N_10995);
and U12299 (N_12299,N_9392,N_10296);
and U12300 (N_12300,N_8587,N_9067);
nor U12301 (N_12301,N_9671,N_10111);
nand U12302 (N_12302,N_11932,N_8924);
nand U12303 (N_12303,N_8957,N_8827);
xnor U12304 (N_12304,N_8966,N_10601);
or U12305 (N_12305,N_9449,N_10701);
nor U12306 (N_12306,N_8747,N_8605);
nor U12307 (N_12307,N_11736,N_9736);
nand U12308 (N_12308,N_10908,N_11822);
xor U12309 (N_12309,N_10372,N_9277);
or U12310 (N_12310,N_11140,N_11030);
xor U12311 (N_12311,N_9128,N_10233);
or U12312 (N_12312,N_9826,N_11831);
and U12313 (N_12313,N_8233,N_10781);
or U12314 (N_12314,N_9019,N_8268);
or U12315 (N_12315,N_11929,N_8260);
or U12316 (N_12316,N_11954,N_8462);
and U12317 (N_12317,N_8124,N_11048);
and U12318 (N_12318,N_10250,N_10700);
nor U12319 (N_12319,N_10720,N_9886);
or U12320 (N_12320,N_8846,N_9015);
or U12321 (N_12321,N_9789,N_11672);
nand U12322 (N_12322,N_8193,N_8198);
xor U12323 (N_12323,N_10048,N_11729);
xor U12324 (N_12324,N_10242,N_11290);
and U12325 (N_12325,N_9846,N_11844);
xor U12326 (N_12326,N_10868,N_9013);
nand U12327 (N_12327,N_8247,N_11426);
and U12328 (N_12328,N_10241,N_8681);
xor U12329 (N_12329,N_8248,N_8050);
and U12330 (N_12330,N_8245,N_11911);
and U12331 (N_12331,N_9232,N_9724);
or U12332 (N_12332,N_9777,N_10737);
nand U12333 (N_12333,N_9375,N_8230);
nor U12334 (N_12334,N_9957,N_8689);
nor U12335 (N_12335,N_10517,N_9241);
nor U12336 (N_12336,N_11811,N_10071);
nor U12337 (N_12337,N_9014,N_8939);
nand U12338 (N_12338,N_8918,N_9654);
nor U12339 (N_12339,N_8687,N_9451);
nand U12340 (N_12340,N_8231,N_11979);
xor U12341 (N_12341,N_8900,N_9112);
xnor U12342 (N_12342,N_10780,N_10047);
or U12343 (N_12343,N_8431,N_9688);
nor U12344 (N_12344,N_9339,N_9869);
nor U12345 (N_12345,N_11691,N_10683);
and U12346 (N_12346,N_11604,N_8584);
and U12347 (N_12347,N_11305,N_11697);
nor U12348 (N_12348,N_9519,N_8258);
xnor U12349 (N_12349,N_9366,N_9093);
and U12350 (N_12350,N_9952,N_8363);
nor U12351 (N_12351,N_11080,N_11565);
and U12352 (N_12352,N_10008,N_11273);
xnor U12353 (N_12353,N_8701,N_9873);
xor U12354 (N_12354,N_11174,N_10865);
or U12355 (N_12355,N_8715,N_9183);
and U12356 (N_12356,N_10014,N_8306);
or U12357 (N_12357,N_10082,N_8236);
xor U12358 (N_12358,N_10912,N_8146);
and U12359 (N_12359,N_11650,N_8209);
nand U12360 (N_12360,N_8454,N_9821);
nor U12361 (N_12361,N_10672,N_10488);
and U12362 (N_12362,N_8591,N_8072);
nor U12363 (N_12363,N_8561,N_9084);
nand U12364 (N_12364,N_11108,N_11839);
xor U12365 (N_12365,N_9598,N_8608);
or U12366 (N_12366,N_9011,N_10541);
xor U12367 (N_12367,N_8871,N_10825);
or U12368 (N_12368,N_9077,N_10935);
nand U12369 (N_12369,N_8496,N_11321);
xor U12370 (N_12370,N_9114,N_8821);
nand U12371 (N_12371,N_11725,N_10699);
and U12372 (N_12372,N_11142,N_10657);
xnor U12373 (N_12373,N_8783,N_8398);
nor U12374 (N_12374,N_8631,N_10743);
nor U12375 (N_12375,N_8249,N_11602);
nor U12376 (N_12376,N_11380,N_8142);
and U12377 (N_12377,N_11060,N_9503);
nand U12378 (N_12378,N_9939,N_9370);
and U12379 (N_12379,N_11170,N_8118);
or U12380 (N_12380,N_11052,N_9489);
nand U12381 (N_12381,N_9354,N_8865);
nand U12382 (N_12382,N_10684,N_9460);
xnor U12383 (N_12383,N_10417,N_8352);
nand U12384 (N_12384,N_8538,N_10382);
xnor U12385 (N_12385,N_10529,N_11955);
and U12386 (N_12386,N_8954,N_10210);
nand U12387 (N_12387,N_11230,N_9927);
or U12388 (N_12388,N_9800,N_11921);
nand U12389 (N_12389,N_8560,N_8833);
nand U12390 (N_12390,N_10645,N_11423);
or U12391 (N_12391,N_9759,N_11881);
nand U12392 (N_12392,N_11342,N_10527);
nor U12393 (N_12393,N_8229,N_9505);
or U12394 (N_12394,N_10654,N_11436);
and U12395 (N_12395,N_8658,N_10451);
nor U12396 (N_12396,N_11367,N_11303);
and U12397 (N_12397,N_11285,N_10882);
and U12398 (N_12398,N_8446,N_11429);
and U12399 (N_12399,N_10862,N_9316);
nand U12400 (N_12400,N_10972,N_10872);
and U12401 (N_12401,N_8737,N_8779);
xor U12402 (N_12402,N_11560,N_10822);
nor U12403 (N_12403,N_10479,N_11039);
and U12404 (N_12404,N_10611,N_10585);
xor U12405 (N_12405,N_10393,N_9247);
nand U12406 (N_12406,N_10930,N_8993);
nand U12407 (N_12407,N_11543,N_8364);
and U12408 (N_12408,N_10900,N_11100);
and U12409 (N_12409,N_10708,N_11332);
nor U12410 (N_12410,N_11622,N_10462);
nand U12411 (N_12411,N_9860,N_10069);
nor U12412 (N_12412,N_10009,N_10994);
nand U12413 (N_12413,N_8346,N_10967);
and U12414 (N_12414,N_11345,N_10109);
xor U12415 (N_12415,N_10386,N_8952);
or U12416 (N_12416,N_8256,N_9537);
xor U12417 (N_12417,N_8207,N_10173);
nor U12418 (N_12418,N_9480,N_9032);
nor U12419 (N_12419,N_8376,N_8158);
and U12420 (N_12420,N_8595,N_11512);
xnor U12421 (N_12421,N_10910,N_9016);
nor U12422 (N_12422,N_10838,N_11431);
nor U12423 (N_12423,N_10127,N_10322);
nand U12424 (N_12424,N_8043,N_9458);
xnor U12425 (N_12425,N_8907,N_10217);
or U12426 (N_12426,N_10916,N_8237);
xnor U12427 (N_12427,N_11673,N_11701);
nand U12428 (N_12428,N_8389,N_11016);
or U12429 (N_12429,N_10168,N_8397);
xnor U12430 (N_12430,N_9527,N_10599);
and U12431 (N_12431,N_11349,N_11191);
and U12432 (N_12432,N_10320,N_11974);
nor U12433 (N_12433,N_9573,N_8976);
xor U12434 (N_12434,N_10656,N_11632);
xnor U12435 (N_12435,N_8058,N_9733);
and U12436 (N_12436,N_11860,N_11255);
nor U12437 (N_12437,N_8310,N_9602);
xor U12438 (N_12438,N_8718,N_10513);
or U12439 (N_12439,N_11006,N_9388);
or U12440 (N_12440,N_8334,N_11312);
nand U12441 (N_12441,N_9387,N_11127);
nand U12442 (N_12442,N_9958,N_10045);
xnor U12443 (N_12443,N_8484,N_11841);
nor U12444 (N_12444,N_9819,N_8469);
and U12445 (N_12445,N_9333,N_11988);
and U12446 (N_12446,N_8823,N_10923);
nor U12447 (N_12447,N_9973,N_9707);
and U12448 (N_12448,N_9857,N_10932);
nor U12449 (N_12449,N_9571,N_9965);
and U12450 (N_12450,N_10396,N_10999);
and U12451 (N_12451,N_11299,N_10723);
and U12452 (N_12452,N_10471,N_11605);
and U12453 (N_12453,N_10530,N_10063);
and U12454 (N_12454,N_8520,N_8765);
xnor U12455 (N_12455,N_9023,N_10260);
and U12456 (N_12456,N_9269,N_10171);
and U12457 (N_12457,N_10113,N_10840);
nor U12458 (N_12458,N_9046,N_10955);
nor U12459 (N_12459,N_9676,N_9631);
nand U12460 (N_12460,N_9469,N_8919);
and U12461 (N_12461,N_9229,N_10143);
nand U12462 (N_12462,N_8070,N_10560);
or U12463 (N_12463,N_10031,N_10120);
nor U12464 (N_12464,N_8616,N_11598);
nand U12465 (N_12465,N_11459,N_8891);
nor U12466 (N_12466,N_10028,N_11229);
nand U12467 (N_12467,N_8175,N_11727);
nor U12468 (N_12468,N_8455,N_8254);
nand U12469 (N_12469,N_8262,N_9069);
nor U12470 (N_12470,N_8206,N_11107);
xor U12471 (N_12471,N_9242,N_10182);
and U12472 (N_12472,N_8368,N_8675);
and U12473 (N_12473,N_9719,N_8819);
and U12474 (N_12474,N_10218,N_10255);
nand U12475 (N_12475,N_9946,N_11904);
xor U12476 (N_12476,N_11403,N_11845);
xor U12477 (N_12477,N_9120,N_9615);
or U12478 (N_12478,N_9085,N_11851);
and U12479 (N_12479,N_8730,N_11797);
nor U12480 (N_12480,N_11824,N_8267);
or U12481 (N_12481,N_11063,N_9841);
nor U12482 (N_12482,N_10365,N_9144);
nor U12483 (N_12483,N_8728,N_11450);
nand U12484 (N_12484,N_9943,N_11284);
nor U12485 (N_12485,N_9265,N_9439);
and U12486 (N_12486,N_8869,N_8650);
or U12487 (N_12487,N_9755,N_11046);
and U12488 (N_12488,N_11325,N_10145);
xor U12489 (N_12489,N_9525,N_8778);
nand U12490 (N_12490,N_10549,N_8932);
nor U12491 (N_12491,N_11420,N_9139);
nand U12492 (N_12492,N_10538,N_10238);
and U12493 (N_12493,N_9337,N_8601);
and U12494 (N_12494,N_10671,N_8575);
nand U12495 (N_12495,N_9044,N_10758);
nor U12496 (N_12496,N_8350,N_10590);
xnor U12497 (N_12497,N_8984,N_10497);
xor U12498 (N_12498,N_9428,N_10425);
or U12499 (N_12499,N_8513,N_9675);
and U12500 (N_12500,N_11638,N_11976);
xor U12501 (N_12501,N_9634,N_8795);
or U12502 (N_12502,N_9726,N_11731);
or U12503 (N_12503,N_10741,N_11326);
nand U12504 (N_12504,N_8787,N_9992);
nor U12505 (N_12505,N_9720,N_8305);
and U12506 (N_12506,N_11609,N_8858);
or U12507 (N_12507,N_9805,N_10149);
or U12508 (N_12508,N_9803,N_8759);
or U12509 (N_12509,N_9308,N_11181);
nand U12510 (N_12510,N_11586,N_11864);
nand U12511 (N_12511,N_10939,N_10554);
nor U12512 (N_12512,N_10944,N_11771);
nor U12513 (N_12513,N_8307,N_10576);
and U12514 (N_12514,N_11716,N_11899);
and U12515 (N_12515,N_10258,N_10276);
nand U12516 (N_12516,N_9892,N_8850);
xnor U12517 (N_12517,N_10083,N_8416);
or U12518 (N_12518,N_10695,N_9871);
xnor U12519 (N_12519,N_11589,N_8686);
nor U12520 (N_12520,N_8304,N_9579);
xor U12521 (N_12521,N_11238,N_8921);
nand U12522 (N_12522,N_8135,N_10013);
and U12523 (N_12523,N_10774,N_11416);
and U12524 (N_12524,N_9630,N_10375);
or U12525 (N_12525,N_11617,N_9063);
nor U12526 (N_12526,N_11295,N_9964);
nand U12527 (N_12527,N_11570,N_11944);
or U12528 (N_12528,N_9143,N_10559);
and U12529 (N_12529,N_10291,N_11798);
and U12530 (N_12530,N_9856,N_11116);
and U12531 (N_12531,N_9095,N_11849);
or U12532 (N_12532,N_11842,N_8942);
or U12533 (N_12533,N_11173,N_9711);
xnor U12534 (N_12534,N_8913,N_11855);
nand U12535 (N_12535,N_8597,N_11511);
nor U12536 (N_12536,N_10811,N_9140);
xnor U12537 (N_12537,N_10974,N_9167);
xor U12538 (N_12538,N_9423,N_10212);
or U12539 (N_12539,N_10514,N_11726);
or U12540 (N_12540,N_9911,N_11306);
or U12541 (N_12541,N_10169,N_9553);
and U12542 (N_12542,N_11491,N_8947);
nand U12543 (N_12543,N_8671,N_8410);
nor U12544 (N_12544,N_8523,N_11205);
or U12545 (N_12545,N_9768,N_10506);
xor U12546 (N_12546,N_10799,N_9940);
or U12547 (N_12547,N_9059,N_8316);
nor U12548 (N_12548,N_11615,N_9725);
and U12549 (N_12549,N_9608,N_10816);
xnor U12550 (N_12550,N_9377,N_10172);
or U12551 (N_12551,N_11015,N_8078);
nor U12552 (N_12552,N_11500,N_9709);
nor U12553 (N_12553,N_8666,N_11027);
and U12554 (N_12554,N_10520,N_9330);
xor U12555 (N_12555,N_11738,N_8008);
nand U12556 (N_12556,N_9723,N_9905);
and U12557 (N_12557,N_8872,N_8156);
nor U12558 (N_12558,N_8754,N_9921);
nand U12559 (N_12559,N_10230,N_10786);
nand U12560 (N_12560,N_8426,N_9403);
nand U12561 (N_12561,N_11557,N_8035);
or U12562 (N_12562,N_10107,N_9961);
xnor U12563 (N_12563,N_11711,N_10032);
and U12564 (N_12564,N_10272,N_9996);
xnor U12565 (N_12565,N_8204,N_10054);
and U12566 (N_12566,N_10926,N_9739);
nand U12567 (N_12567,N_9893,N_8882);
or U12568 (N_12568,N_8653,N_9235);
nor U12569 (N_12569,N_11194,N_9146);
or U12570 (N_12570,N_8840,N_11101);
xor U12571 (N_12571,N_8402,N_8355);
xor U12572 (N_12572,N_10540,N_11289);
nor U12573 (N_12573,N_9251,N_11043);
or U12574 (N_12574,N_9272,N_9872);
and U12575 (N_12575,N_9342,N_11834);
and U12576 (N_12576,N_8333,N_9275);
nand U12577 (N_12577,N_11344,N_8744);
and U12578 (N_12578,N_9294,N_8678);
xor U12579 (N_12579,N_8329,N_11175);
or U12580 (N_12580,N_11081,N_10057);
or U12581 (N_12581,N_9746,N_9637);
nor U12582 (N_12582,N_8611,N_10379);
and U12583 (N_12583,N_10697,N_10313);
nor U12584 (N_12584,N_8546,N_10354);
or U12585 (N_12585,N_9162,N_9008);
nor U12586 (N_12586,N_11554,N_9482);
xor U12587 (N_12587,N_9618,N_8828);
nand U12588 (N_12588,N_9397,N_8399);
and U12589 (N_12589,N_11217,N_10472);
and U12590 (N_12590,N_8781,N_10346);
nand U12591 (N_12591,N_10137,N_11160);
xnor U12592 (N_12592,N_11940,N_9291);
nor U12593 (N_12593,N_11102,N_9929);
or U12594 (N_12594,N_8279,N_10952);
or U12595 (N_12595,N_8571,N_10662);
nand U12596 (N_12596,N_10077,N_9465);
or U12597 (N_12597,N_11505,N_9552);
nand U12598 (N_12598,N_8606,N_9932);
or U12599 (N_12599,N_9782,N_10748);
nand U12600 (N_12600,N_9496,N_9718);
and U12601 (N_12601,N_9470,N_10033);
or U12602 (N_12602,N_11774,N_11028);
or U12603 (N_12603,N_10443,N_8979);
nor U12604 (N_12604,N_9092,N_8296);
nor U12605 (N_12605,N_9862,N_9989);
nor U12606 (N_12606,N_9665,N_10892);
or U12607 (N_12607,N_10489,N_10074);
or U12608 (N_12608,N_8792,N_9875);
xnor U12609 (N_12609,N_10567,N_11308);
nand U12610 (N_12610,N_11544,N_9374);
or U12611 (N_12611,N_8373,N_11760);
xor U12612 (N_12612,N_11020,N_9386);
or U12613 (N_12613,N_8723,N_9292);
xnor U12614 (N_12614,N_8122,N_11361);
and U12615 (N_12615,N_11667,N_9629);
xor U12616 (N_12616,N_10440,N_11591);
nand U12617 (N_12617,N_11992,N_11640);
nor U12618 (N_12618,N_10220,N_9901);
nand U12619 (N_12619,N_9237,N_10906);
nand U12620 (N_12620,N_10859,N_10174);
nand U12621 (N_12621,N_8432,N_11456);
or U12622 (N_12622,N_8366,N_11610);
nand U12623 (N_12623,N_9937,N_8059);
xnor U12624 (N_12624,N_10998,N_9053);
xnor U12625 (N_12625,N_9521,N_9766);
nor U12626 (N_12626,N_9569,N_10641);
nand U12627 (N_12627,N_11509,N_9025);
nor U12628 (N_12628,N_11145,N_10001);
and U12629 (N_12629,N_11398,N_9659);
xor U12630 (N_12630,N_9285,N_8391);
nor U12631 (N_12631,N_11263,N_9210);
or U12632 (N_12632,N_8698,N_8662);
nand U12633 (N_12633,N_10249,N_8517);
or U12634 (N_12634,N_8902,N_10771);
and U12635 (N_12635,N_11267,N_10920);
nor U12636 (N_12636,N_9648,N_11577);
or U12637 (N_12637,N_9657,N_10181);
or U12638 (N_12638,N_9040,N_10135);
xor U12639 (N_12639,N_8945,N_9224);
nand U12640 (N_12640,N_11470,N_9515);
or U12641 (N_12641,N_9369,N_9520);
and U12642 (N_12642,N_11941,N_10605);
xnor U12643 (N_12643,N_9781,N_10528);
xnor U12644 (N_12644,N_8532,N_8526);
xor U12645 (N_12645,N_8804,N_8748);
nor U12646 (N_12646,N_10349,N_8485);
xnor U12647 (N_12647,N_11653,N_11327);
and U12648 (N_12648,N_9321,N_8674);
xor U12649 (N_12649,N_11259,N_8563);
xor U12650 (N_12650,N_8278,N_10670);
xor U12651 (N_12651,N_10787,N_11114);
xnor U12652 (N_12652,N_10833,N_10856);
and U12653 (N_12653,N_10836,N_8087);
nand U12654 (N_12654,N_9117,N_10485);
and U12655 (N_12655,N_9792,N_11540);
and U12656 (N_12656,N_10943,N_8548);
or U12657 (N_12657,N_11497,N_8731);
and U12658 (N_12658,N_10563,N_10634);
or U12659 (N_12659,N_9561,N_8361);
nand U12660 (N_12660,N_10277,N_9963);
nor U12661 (N_12661,N_8062,N_10132);
or U12662 (N_12662,N_11453,N_9909);
and U12663 (N_12663,N_10301,N_11336);
xor U12664 (N_12664,N_8667,N_11319);
or U12665 (N_12665,N_10773,N_10512);
and U12666 (N_12666,N_8358,N_10079);
and U12667 (N_12667,N_8829,N_9920);
nor U12668 (N_12668,N_8570,N_9653);
nor U12669 (N_12669,N_9824,N_8092);
and U12670 (N_12670,N_10064,N_9288);
nor U12671 (N_12671,N_8514,N_10660);
xor U12672 (N_12672,N_8145,N_9784);
or U12673 (N_12673,N_9445,N_8478);
and U12674 (N_12674,N_9378,N_11157);
or U12675 (N_12675,N_11643,N_9740);
or U12676 (N_12676,N_11269,N_11847);
nor U12677 (N_12677,N_11784,N_11787);
xnor U12678 (N_12678,N_9497,N_10154);
nor U12679 (N_12679,N_8564,N_9267);
nand U12680 (N_12680,N_11585,N_10744);
xor U12681 (N_12681,N_8383,N_9760);
xor U12682 (N_12682,N_8270,N_9756);
or U12683 (N_12683,N_9747,N_11406);
and U12684 (N_12684,N_9226,N_11239);
or U12685 (N_12685,N_9158,N_9651);
nor U12686 (N_12686,N_11013,N_10287);
or U12687 (N_12687,N_10564,N_10395);
nor U12688 (N_12688,N_10499,N_11776);
and U12689 (N_12689,N_8150,N_10543);
and U12690 (N_12690,N_9835,N_8242);
or U12691 (N_12691,N_11124,N_8214);
and U12692 (N_12692,N_8746,N_8205);
nor U12693 (N_12693,N_11430,N_11167);
xor U12694 (N_12694,N_10483,N_8244);
xnor U12695 (N_12695,N_11715,N_8104);
xor U12696 (N_12696,N_8335,N_11951);
or U12697 (N_12697,N_8814,N_8165);
and U12698 (N_12698,N_9988,N_8007);
nor U12699 (N_12699,N_8659,N_8941);
or U12700 (N_12700,N_8018,N_8133);
xnor U12701 (N_12701,N_8212,N_8036);
nor U12702 (N_12702,N_9395,N_9908);
and U12703 (N_12703,N_11244,N_11963);
nand U12704 (N_12704,N_11905,N_8722);
xnor U12705 (N_12705,N_10176,N_11754);
nand U12706 (N_12706,N_8369,N_11469);
nor U12707 (N_12707,N_11360,N_8185);
nand U12708 (N_12708,N_10025,N_9329);
nand U12709 (N_12709,N_10356,N_9512);
and U12710 (N_12710,N_10579,N_11184);
nor U12711 (N_12711,N_11803,N_10416);
nand U12712 (N_12712,N_8384,N_9678);
nand U12713 (N_12713,N_10663,N_10078);
or U12714 (N_12714,N_11832,N_8380);
xor U12715 (N_12715,N_8002,N_8130);
nor U12716 (N_12716,N_10953,N_11903);
or U12717 (N_12717,N_8637,N_11226);
and U12718 (N_12718,N_10131,N_9594);
xor U12719 (N_12719,N_10085,N_11785);
or U12720 (N_12720,N_9843,N_10861);
nor U12721 (N_12721,N_8438,N_10121);
nand U12722 (N_12722,N_11373,N_9882);
nor U12723 (N_12723,N_10208,N_11521);
nor U12724 (N_12724,N_9668,N_8509);
and U12725 (N_12725,N_10950,N_11668);
and U12726 (N_12726,N_8379,N_11750);
and U12727 (N_12727,N_10091,N_9955);
or U12728 (N_12728,N_11690,N_9176);
nor U12729 (N_12729,N_8053,N_9754);
and U12730 (N_12730,N_8636,N_9550);
nor U12731 (N_12731,N_10294,N_8669);
nand U12732 (N_12732,N_8610,N_10519);
or U12733 (N_12733,N_8387,N_10326);
or U12734 (N_12734,N_9850,N_9547);
nand U12735 (N_12735,N_10651,N_8812);
xnor U12736 (N_12736,N_11106,N_8404);
nor U12737 (N_12737,N_9297,N_10456);
nand U12738 (N_12738,N_8057,N_9111);
or U12739 (N_12739,N_8660,N_10165);
and U12740 (N_12740,N_8972,N_10837);
nor U12741 (N_12741,N_9624,N_10288);
nand U12742 (N_12742,N_10177,N_10450);
or U12743 (N_12743,N_10949,N_8836);
nor U12744 (N_12744,N_9891,N_8412);
xor U12745 (N_12745,N_10434,N_8853);
nand U12746 (N_12746,N_10961,N_8377);
xor U12747 (N_12747,N_11999,N_8300);
nor U12748 (N_12748,N_8717,N_11058);
or U12749 (N_12749,N_8969,N_8458);
or U12750 (N_12750,N_10205,N_11906);
nor U12751 (N_12751,N_8489,N_10779);
and U12752 (N_12752,N_11396,N_10447);
nand U12753 (N_12753,N_8132,N_9184);
or U12754 (N_12754,N_11582,N_8703);
nand U12755 (N_12755,N_11210,N_11813);
xor U12756 (N_12756,N_11232,N_10185);
nand U12757 (N_12757,N_10061,N_11062);
or U12758 (N_12758,N_11369,N_9368);
xnor U12759 (N_12759,N_8178,N_8881);
xnor U12760 (N_12760,N_9508,N_9545);
and U12761 (N_12761,N_8048,N_10140);
nor U12762 (N_12762,N_8159,N_8958);
and U12763 (N_12763,N_10100,N_10842);
xor U12764 (N_12764,N_9199,N_10533);
or U12765 (N_12765,N_11623,N_8199);
xor U12766 (N_12766,N_11158,N_8986);
xnor U12767 (N_12767,N_10992,N_11189);
nor U12768 (N_12768,N_8147,N_10502);
and U12769 (N_12769,N_10919,N_8418);
xor U12770 (N_12770,N_11619,N_8488);
xnor U12771 (N_12771,N_8210,N_11599);
xnor U12772 (N_12772,N_10222,N_10055);
nand U12773 (N_12773,N_11821,N_9748);
nor U12774 (N_12774,N_8602,N_9902);
xnor U12775 (N_12775,N_9960,N_8630);
nor U12776 (N_12776,N_8382,N_8498);
xnor U12777 (N_12777,N_11096,N_9170);
xor U12778 (N_12778,N_8773,N_8541);
nand U12779 (N_12779,N_9809,N_10815);
or U12780 (N_12780,N_9424,N_11490);
and U12781 (N_12781,N_8055,N_8506);
nor U12782 (N_12782,N_8327,N_10924);
nor U12783 (N_12783,N_11348,N_9301);
nand U12784 (N_12784,N_11093,N_8824);
and U12785 (N_12785,N_9261,N_9236);
or U12786 (N_12786,N_10612,N_11538);
nor U12787 (N_12787,N_10360,N_9461);
nor U12788 (N_12788,N_10310,N_11452);
or U12789 (N_12789,N_10459,N_11159);
nand U12790 (N_12790,N_11440,N_9454);
nand U12791 (N_12791,N_10056,N_9580);
xnor U12792 (N_12792,N_9974,N_11180);
xor U12793 (N_12793,N_10464,N_10980);
xnor U12794 (N_12794,N_9641,N_11218);
nand U12795 (N_12795,N_10975,N_9462);
and U12796 (N_12796,N_10557,N_11924);
or U12797 (N_12797,N_10993,N_10253);
and U12798 (N_12798,N_8770,N_9234);
and U12799 (N_12799,N_10679,N_8768);
nand U12800 (N_12800,N_9919,N_10398);
nor U12801 (N_12801,N_8543,N_9326);
xor U12802 (N_12802,N_11664,N_9271);
nor U12803 (N_12803,N_11123,N_10202);
or U12804 (N_12804,N_9572,N_8341);
and U12805 (N_12805,N_8311,N_11665);
and U12806 (N_12806,N_9325,N_10714);
or U12807 (N_12807,N_9356,N_11183);
xnor U12808 (N_12808,N_10945,N_10586);
nand U12809 (N_12809,N_8112,N_11718);
nand U12810 (N_12810,N_11359,N_11292);
nand U12811 (N_12811,N_10223,N_11186);
nand U12812 (N_12812,N_11815,N_8051);
nor U12813 (N_12813,N_11768,N_9734);
xor U12814 (N_12814,N_11247,N_9412);
nand U12815 (N_12815,N_10973,N_11972);
and U12816 (N_12816,N_9246,N_9881);
nor U12817 (N_12817,N_8286,N_11010);
or U12818 (N_12818,N_11053,N_8162);
and U12819 (N_12819,N_8634,N_9071);
xor U12820 (N_12820,N_9036,N_9765);
xnor U12821 (N_12821,N_11258,N_9914);
nand U12822 (N_12822,N_11656,N_10088);
nor U12823 (N_12823,N_11868,N_8238);
nor U12824 (N_12824,N_10733,N_8567);
nand U12825 (N_12825,N_10979,N_10879);
and U12826 (N_12826,N_10523,N_8302);
xnor U12827 (N_12827,N_10423,N_9201);
nor U12828 (N_12828,N_9418,N_11177);
nor U12829 (N_12829,N_11399,N_8201);
or U12830 (N_12830,N_11385,N_11545);
nand U12831 (N_12831,N_8998,N_11910);
xor U12832 (N_12832,N_8213,N_11625);
nand U12833 (N_12833,N_9182,N_10962);
nor U12834 (N_12834,N_11168,N_9652);
nor U12835 (N_12835,N_10364,N_8551);
nand U12836 (N_12836,N_9060,N_10010);
nand U12837 (N_12837,N_9773,N_8354);
nor U12838 (N_12838,N_10963,N_8652);
or U12839 (N_12839,N_9900,N_9794);
or U12840 (N_12840,N_11788,N_9094);
xnor U12841 (N_12841,N_11519,N_11829);
and U12842 (N_12842,N_11487,N_10123);
nor U12843 (N_12843,N_8166,N_11858);
or U12844 (N_12844,N_11130,N_11143);
xor U12845 (N_12845,N_9640,N_9425);
nor U12846 (N_12846,N_11807,N_9986);
nor U12847 (N_12847,N_11655,N_10728);
xor U12848 (N_12848,N_11437,N_9870);
xnor U12849 (N_12849,N_9066,N_11641);
nand U12850 (N_12850,N_9560,N_8401);
nor U12851 (N_12851,N_9823,N_8225);
xor U12852 (N_12852,N_11037,N_9941);
and U12853 (N_12853,N_11132,N_8580);
and U12854 (N_12854,N_11001,N_8126);
and U12855 (N_12855,N_8084,N_8851);
or U12856 (N_12856,N_10587,N_9252);
nand U12857 (N_12857,N_9064,N_10090);
nor U12858 (N_12858,N_11097,N_10461);
xnor U12859 (N_12859,N_10116,N_9528);
or U12860 (N_12860,N_11573,N_11475);
nor U12861 (N_12861,N_11294,N_8510);
or U12862 (N_12862,N_10097,N_9738);
xor U12863 (N_12863,N_11256,N_8289);
nor U12864 (N_12864,N_8161,N_9276);
nor U12865 (N_12865,N_10170,N_10620);
xor U12866 (N_12866,N_10317,N_11534);
xnor U12867 (N_12867,N_8889,N_8220);
and U12868 (N_12868,N_10041,N_10855);
or U12869 (N_12869,N_9840,N_11993);
or U12870 (N_12870,N_8134,N_8885);
xor U12871 (N_12871,N_9096,N_8672);
nand U12872 (N_12872,N_11983,N_10688);
xnor U12873 (N_12873,N_8090,N_10437);
nand U12874 (N_12874,N_9003,N_11888);
nor U12875 (N_12875,N_10358,N_10299);
xor U12876 (N_12876,N_9880,N_8859);
nand U12877 (N_12877,N_8528,N_10102);
or U12878 (N_12878,N_10655,N_9851);
nand U12879 (N_12879,N_9959,N_9355);
nand U12880 (N_12880,N_10244,N_9078);
nand U12881 (N_12881,N_10880,N_9435);
nor U12882 (N_12882,N_8024,N_10463);
xnor U12883 (N_12883,N_8026,N_10849);
nor U12884 (N_12884,N_8448,N_11859);
and U12885 (N_12885,N_10475,N_9938);
xor U12886 (N_12886,N_9638,N_8683);
or U12887 (N_12887,N_10894,N_8282);
nand U12888 (N_12888,N_9544,N_8959);
xnor U12889 (N_12889,N_8482,N_8101);
and U12890 (N_12890,N_8874,N_9463);
and U12891 (N_12891,N_11064,N_10267);
nor U12892 (N_12892,N_11083,N_11524);
nor U12893 (N_12893,N_11966,N_8518);
nand U12894 (N_12894,N_10080,N_9818);
xor U12895 (N_12895,N_9352,N_11706);
nand U12896 (N_12896,N_8901,N_9543);
or U12897 (N_12897,N_8028,N_9101);
nand U12898 (N_12898,N_9029,N_10981);
or U12899 (N_12899,N_11197,N_10765);
or U12900 (N_12900,N_10268,N_11019);
or U12901 (N_12901,N_9670,N_11427);
xor U12902 (N_12902,N_9038,N_9065);
or U12903 (N_12903,N_10232,N_11945);
nand U12904 (N_12904,N_8676,N_8056);
and U12905 (N_12905,N_11968,N_10783);
xor U12906 (N_12906,N_9100,N_11283);
or U12907 (N_12907,N_9173,N_10761);
or U12908 (N_12908,N_11352,N_11404);
nor U12909 (N_12909,N_11388,N_9536);
nand U12910 (N_12910,N_9693,N_11997);
nand U12911 (N_12911,N_8811,N_10966);
and U12912 (N_12912,N_10608,N_9116);
and U12913 (N_12913,N_11994,N_11417);
nor U12914 (N_12914,N_10661,N_11818);
nor U12915 (N_12915,N_11620,N_9193);
and U12916 (N_12916,N_10847,N_11695);
and U12917 (N_12917,N_8121,N_10851);
nand U12918 (N_12918,N_10846,N_9861);
nor U12919 (N_12919,N_10857,N_9799);
xnor U12920 (N_12920,N_9200,N_9565);
xnor U12921 (N_12921,N_10957,N_9466);
and U12922 (N_12922,N_8761,N_11884);
nor U12923 (N_12923,N_11389,N_11686);
and U12924 (N_12924,N_9757,N_9152);
and U12925 (N_12925,N_10248,N_9625);
and U12926 (N_12926,N_10094,N_10753);
xnor U12927 (N_12927,N_9371,N_11748);
nand U12928 (N_12928,N_11464,N_8116);
or U12929 (N_12929,N_11120,N_8172);
nand U12930 (N_12930,N_9567,N_9614);
and U12931 (N_12931,N_10424,N_8123);
nand U12932 (N_12932,N_8015,N_8490);
and U12933 (N_12933,N_10159,N_8127);
or U12934 (N_12934,N_8360,N_11917);
or U12935 (N_12935,N_11600,N_10504);
xnor U12936 (N_12936,N_8890,N_11302);
or U12937 (N_12937,N_8424,N_8508);
nand U12938 (N_12938,N_9953,N_11937);
or U12939 (N_12939,N_11187,N_9314);
nor U12940 (N_12940,N_8556,N_8790);
xnor U12941 (N_12941,N_10164,N_8930);
nor U12942 (N_12942,N_10281,N_10525);
and U12943 (N_12943,N_9744,N_8030);
and U12944 (N_12944,N_9549,N_9522);
xor U12945 (N_12945,N_9319,N_10228);
xnor U12946 (N_12946,N_8422,N_11002);
nand U12947 (N_12947,N_10721,N_9351);
or U12948 (N_12948,N_11809,N_8844);
and U12949 (N_12949,N_9583,N_8645);
and U12950 (N_12950,N_11446,N_9874);
nand U12951 (N_12951,N_11041,N_10226);
nor U12952 (N_12952,N_9682,N_8103);
and U12953 (N_12953,N_9302,N_11801);
nor U12954 (N_12954,N_8691,N_11462);
xor U12955 (N_12955,N_11734,N_11442);
nor U12956 (N_12956,N_11278,N_8794);
nor U12957 (N_12957,N_11264,N_11721);
or U12958 (N_12958,N_11122,N_10216);
nand U12959 (N_12959,N_11580,N_9833);
and U12960 (N_12960,N_8098,N_11161);
nand U12961 (N_12961,N_10639,N_10883);
nor U12962 (N_12962,N_9877,N_9933);
nor U12963 (N_12963,N_11722,N_9175);
and U12964 (N_12964,N_9168,N_8716);
nand U12965 (N_12965,N_11862,N_11131);
or U12966 (N_12966,N_11068,N_8295);
or U12967 (N_12967,N_11018,N_10875);
xor U12968 (N_12968,N_10053,N_11357);
or U12969 (N_12969,N_11761,N_10449);
or U12970 (N_12970,N_11212,N_8640);
nor U12971 (N_12971,N_9205,N_9054);
and U12972 (N_12972,N_11943,N_8613);
nand U12973 (N_12973,N_8697,N_9102);
or U12974 (N_12974,N_8374,N_9593);
and U12975 (N_12975,N_10507,N_8343);
xor U12976 (N_12976,N_9384,N_11683);
nand U12977 (N_12977,N_10017,N_9151);
and U12978 (N_12978,N_8855,N_8388);
or U12979 (N_12979,N_8529,N_10160);
nor U12980 (N_12980,N_11314,N_8995);
nor U12981 (N_12981,N_10588,N_8082);
or U12982 (N_12982,N_9538,N_8668);
and U12983 (N_12983,N_8978,N_8280);
nand U12984 (N_12984,N_11381,N_10760);
and U12985 (N_12985,N_10547,N_11991);
nor U12986 (N_12986,N_10850,N_9253);
nor U12987 (N_12987,N_11871,N_11144);
nor U12988 (N_12988,N_9853,N_11347);
and U12989 (N_12989,N_11874,N_10035);
and U12990 (N_12990,N_11031,N_8536);
nor U12991 (N_12991,N_9910,N_10871);
or U12992 (N_12992,N_8396,N_8685);
and U12993 (N_12993,N_10845,N_10460);
or U12994 (N_12994,N_8757,N_11339);
nor U12995 (N_12995,N_9804,N_10526);
xnor U12996 (N_12996,N_10282,N_9331);
nor U12997 (N_12997,N_11091,N_10397);
nor U12998 (N_12998,N_8285,N_8502);
and U12999 (N_12999,N_11465,N_8586);
or U13000 (N_13000,N_9926,N_10199);
and U13001 (N_13001,N_10155,N_8839);
nor U13002 (N_13002,N_10982,N_11645);
xnor U13003 (N_13003,N_9473,N_8184);
nand U13004 (N_13004,N_11126,N_9763);
xor U13005 (N_13005,N_10300,N_8980);
xor U13006 (N_13006,N_9262,N_10433);
xnor U13007 (N_13007,N_10442,N_8290);
or U13008 (N_13008,N_11732,N_11208);
nand U13009 (N_13009,N_9876,N_9000);
nor U13010 (N_13010,N_9298,N_10262);
nor U13011 (N_13011,N_10911,N_11915);
nor U13012 (N_13012,N_9486,N_11828);
nor U13013 (N_13013,N_10246,N_11350);
and U13014 (N_13014,N_8378,N_8331);
nor U13015 (N_13015,N_11201,N_10764);
nor U13016 (N_13016,N_10650,N_8933);
nand U13017 (N_13017,N_9105,N_10036);
or U13018 (N_13018,N_8782,N_9110);
nor U13019 (N_13019,N_9810,N_8504);
and U13020 (N_13020,N_10685,N_11737);
and U13021 (N_13021,N_9981,N_8705);
or U13022 (N_13022,N_11009,N_11236);
nand U13023 (N_13023,N_8784,N_10637);
and U13024 (N_13024,N_11594,N_9622);
xnor U13025 (N_13025,N_9616,N_9477);
or U13026 (N_13026,N_11507,N_11483);
or U13027 (N_13027,N_8780,N_9118);
nand U13028 (N_13028,N_9012,N_9815);
or U13029 (N_13029,N_11681,N_8323);
xnor U13030 (N_13030,N_11090,N_11297);
or U13031 (N_13031,N_10142,N_10886);
nor U13032 (N_13032,N_11779,N_11476);
xor U13033 (N_13033,N_9091,N_10371);
or U13034 (N_13034,N_10298,N_9172);
and U13035 (N_13035,N_11109,N_11421);
or U13036 (N_13036,N_8196,N_9807);
xor U13037 (N_13037,N_9021,N_11646);
xor U13038 (N_13038,N_8642,N_10652);
and U13039 (N_13039,N_10752,N_11110);
nand U13040 (N_13040,N_9320,N_9327);
and U13041 (N_13041,N_8899,N_8905);
or U13042 (N_13042,N_10331,N_9588);
xor U13043 (N_13043,N_9255,N_10808);
or U13044 (N_13044,N_10788,N_11613);
and U13045 (N_13045,N_9222,N_9177);
and U13046 (N_13046,N_11551,N_10128);
or U13047 (N_13047,N_8203,N_11266);
nand U13048 (N_13048,N_8910,N_9661);
and U13049 (N_13049,N_11633,N_11568);
or U13050 (N_13050,N_11280,N_8917);
xor U13051 (N_13051,N_9231,N_9514);
nor U13052 (N_13052,N_10474,N_9062);
nand U13053 (N_13053,N_8732,N_9160);
xnor U13054 (N_13054,N_10508,N_9969);
and U13055 (N_13055,N_11928,N_9007);
nor U13056 (N_13056,N_8275,N_11578);
and U13057 (N_13057,N_8149,N_10415);
and U13058 (N_13058,N_11065,N_10638);
nor U13059 (N_13059,N_9447,N_11012);
nand U13060 (N_13060,N_8742,N_9230);
xnor U13061 (N_13061,N_10308,N_11666);
xnor U13062 (N_13062,N_11981,N_8096);
and U13063 (N_13063,N_10157,N_11317);
nand U13064 (N_13064,N_10703,N_9137);
nor U13065 (N_13065,N_8621,N_8107);
nand U13066 (N_13066,N_11035,N_9487);
and U13067 (N_13067,N_11529,N_10352);
nor U13068 (N_13068,N_11202,N_8453);
xnor U13069 (N_13069,N_9076,N_10357);
and U13070 (N_13070,N_10675,N_11152);
nor U13071 (N_13071,N_10043,N_10103);
nor U13072 (N_13072,N_11624,N_10867);
or U13073 (N_13073,N_8550,N_10524);
nor U13074 (N_13074,N_11498,N_8515);
xor U13075 (N_13075,N_8060,N_11635);
nor U13076 (N_13076,N_11343,N_10633);
nand U13077 (N_13077,N_11076,N_8200);
or U13078 (N_13078,N_8226,N_10843);
and U13079 (N_13079,N_9970,N_10792);
xnor U13080 (N_13080,N_11885,N_9663);
xnor U13081 (N_13081,N_9429,N_9945);
nand U13082 (N_13082,N_11137,N_8927);
nor U13083 (N_13083,N_9533,N_10844);
nand U13084 (N_13084,N_9664,N_8415);
xor U13085 (N_13085,N_9296,N_11564);
nand U13086 (N_13086,N_9689,N_9742);
xnor U13087 (N_13087,N_11073,N_10754);
or U13088 (N_13088,N_11182,N_8250);
and U13089 (N_13089,N_11301,N_10341);
nor U13090 (N_13090,N_10782,N_8857);
or U13091 (N_13091,N_10928,N_9510);
nor U13092 (N_13092,N_10081,N_9407);
xor U13093 (N_13093,N_8074,N_9795);
nand U13094 (N_13094,N_8183,N_11696);
xnor U13095 (N_13095,N_11663,N_8297);
nor U13096 (N_13096,N_10834,N_9245);
nor U13097 (N_13097,N_10093,N_11528);
nor U13098 (N_13098,N_8086,N_9420);
nor U13099 (N_13099,N_10339,N_11587);
xnor U13100 (N_13100,N_8531,N_9865);
or U13101 (N_13101,N_8143,N_10627);
xnor U13102 (N_13102,N_11719,N_8287);
and U13103 (N_13103,N_11246,N_11243);
and U13104 (N_13104,N_8435,N_9806);
nand U13105 (N_13105,N_8308,N_9591);
xor U13106 (N_13106,N_8001,N_10592);
nor U13107 (N_13107,N_11092,N_11658);
xor U13108 (N_13108,N_9430,N_8359);
nand U13109 (N_13109,N_8724,N_10619);
xnor U13110 (N_13110,N_10122,N_10521);
or U13111 (N_13111,N_11506,N_10931);
or U13112 (N_13112,N_10275,N_11231);
xnor U13113 (N_13113,N_11927,N_10445);
and U13114 (N_13114,N_8884,N_8994);
nand U13115 (N_13115,N_9282,N_11789);
or U13116 (N_13116,N_8367,N_10624);
xor U13117 (N_13117,N_11365,N_9845);
nand U13118 (N_13118,N_8537,N_11198);
or U13119 (N_13119,N_10958,N_9122);
and U13120 (N_13120,N_8461,N_8239);
nor U13121 (N_13121,N_10951,N_11710);
nand U13122 (N_13122,N_10578,N_10368);
or U13123 (N_13123,N_10854,N_11003);
xor U13124 (N_13124,N_9511,N_8299);
nor U13125 (N_13125,N_11597,N_11873);
nor U13126 (N_13126,N_10562,N_11550);
nand U13127 (N_13127,N_11827,N_8745);
xnor U13128 (N_13128,N_11925,N_10092);
nand U13129 (N_13129,N_11890,N_8054);
nor U13130 (N_13130,N_10936,N_10050);
or U13131 (N_13131,N_9214,N_10724);
nand U13132 (N_13132,N_10510,N_11793);
or U13133 (N_13133,N_11155,N_8695);
or U13134 (N_13134,N_11907,N_9490);
or U13135 (N_13135,N_10647,N_9431);
and U13136 (N_13136,N_11499,N_10402);
or U13137 (N_13137,N_11328,N_9204);
and U13138 (N_13138,N_11852,N_10224);
or U13139 (N_13139,N_8261,N_11527);
nor U13140 (N_13140,N_10545,N_10161);
and U13141 (N_13141,N_9048,N_9233);
nand U13142 (N_13142,N_9123,N_9716);
or U13143 (N_13143,N_10613,N_10591);
or U13144 (N_13144,N_11533,N_9925);
nand U13145 (N_13145,N_11393,N_9717);
or U13146 (N_13146,N_8115,N_10745);
or U13147 (N_13147,N_11764,N_9535);
nor U13148 (N_13148,N_11094,N_9728);
xor U13149 (N_13149,N_8841,N_11494);
xnor U13150 (N_13150,N_8815,N_11477);
nand U13151 (N_13151,N_8294,N_8047);
or U13152 (N_13152,N_11535,N_10666);
and U13153 (N_13153,N_10832,N_8624);
nor U13154 (N_13154,N_11883,N_10791);
xnor U13155 (N_13155,N_11163,N_9499);
and U13156 (N_13156,N_10239,N_9801);
or U13157 (N_13157,N_10200,N_10902);
and U13158 (N_13158,N_10189,N_8417);
nand U13159 (N_13159,N_10087,N_10361);
nor U13160 (N_13160,N_11298,N_8153);
nand U13161 (N_13161,N_8117,N_9312);
and U13162 (N_13162,N_10439,N_8617);
and U13163 (N_13163,N_11484,N_10075);
or U13164 (N_13164,N_8741,N_11353);
nor U13165 (N_13165,N_10727,N_10040);
xnor U13166 (N_13166,N_9350,N_11796);
and U13167 (N_13167,N_11139,N_10188);
nor U13168 (N_13168,N_8272,N_10726);
or U13169 (N_13169,N_10166,N_10694);
nand U13170 (N_13170,N_11023,N_11495);
or U13171 (N_13171,N_10584,N_8427);
or U13172 (N_13172,N_10903,N_10283);
nand U13173 (N_13173,N_8596,N_8776);
or U13174 (N_13174,N_11651,N_8934);
nand U13175 (N_13175,N_8915,N_8442);
or U13176 (N_13176,N_9195,N_10674);
nor U13177 (N_13177,N_9820,N_9916);
nand U13178 (N_13178,N_9359,N_9997);
nand U13179 (N_13179,N_11892,N_10038);
nand U13180 (N_13180,N_8625,N_10465);
xor U13181 (N_13181,N_11517,N_9290);
xor U13182 (N_13182,N_9564,N_9030);
nand U13183 (N_13183,N_11749,N_8665);
and U13184 (N_13184,N_10730,N_9433);
nor U13185 (N_13185,N_8080,N_11104);
xnor U13186 (N_13186,N_11392,N_11485);
xor U13187 (N_13187,N_9186,N_10986);
nor U13188 (N_13188,N_10610,N_11112);
nand U13189 (N_13189,N_9702,N_8171);
or U13190 (N_13190,N_9644,N_9586);
nand U13191 (N_13191,N_11895,N_10259);
or U13192 (N_13192,N_10492,N_10235);
or U13193 (N_13193,N_10706,N_10767);
nor U13194 (N_13194,N_8574,N_9106);
nor U13195 (N_13195,N_10144,N_10742);
and U13196 (N_13196,N_11938,N_8711);
xnor U13197 (N_13197,N_11778,N_9394);
and U13198 (N_13198,N_10826,N_10118);
or U13199 (N_13199,N_10234,N_11843);
nand U13200 (N_13200,N_9075,N_10221);
nor U13201 (N_13201,N_8069,N_11769);
or U13202 (N_13202,N_9041,N_10756);
or U13203 (N_13203,N_9694,N_10677);
or U13204 (N_13204,N_9228,N_8394);
and U13205 (N_13205,N_11395,N_9621);
nor U13206 (N_13206,N_8592,N_9859);
and U13207 (N_13207,N_11960,N_8860);
or U13208 (N_13208,N_11659,N_9187);
or U13209 (N_13209,N_11171,N_9797);
xnor U13210 (N_13210,N_10058,N_9626);
nor U13211 (N_13211,N_8714,N_8385);
and U13212 (N_13212,N_11434,N_9028);
or U13213 (N_13213,N_11950,N_9894);
or U13214 (N_13214,N_9683,N_10573);
or U13215 (N_13215,N_8114,N_8738);
nor U13216 (N_13216,N_9338,N_10515);
nor U13217 (N_13217,N_11400,N_9332);
and U13218 (N_13218,N_11703,N_9121);
xnor U13219 (N_13219,N_11042,N_8337);
and U13220 (N_13220,N_8985,N_8981);
or U13221 (N_13221,N_8734,N_10381);
xnor U13222 (N_13222,N_8284,N_10225);
or U13223 (N_13223,N_9303,N_9898);
and U13224 (N_13224,N_11901,N_10542);
or U13225 (N_13225,N_9135,N_10705);
xor U13226 (N_13226,N_8407,N_10000);
or U13227 (N_13227,N_9345,N_9896);
xnor U13228 (N_13228,N_8174,N_10229);
nand U13229 (N_13229,N_10405,N_10858);
nor U13230 (N_13230,N_11079,N_9930);
nor U13231 (N_13231,N_9328,N_8708);
or U13232 (N_13232,N_11786,N_11121);
and U13233 (N_13233,N_11215,N_10817);
nand U13234 (N_13234,N_9701,N_10853);
nor U13235 (N_13235,N_11913,N_11281);
or U13236 (N_13236,N_8252,N_10197);
xor U13237 (N_13237,N_8494,N_10877);
and U13238 (N_13238,N_11792,N_9524);
nand U13239 (N_13239,N_9472,N_9364);
nand U13240 (N_13240,N_8982,N_10355);
and U13241 (N_13241,N_8663,N_9266);
nor U13242 (N_13242,N_9787,N_9596);
or U13243 (N_13243,N_8152,N_8016);
xor U13244 (N_13244,N_10736,N_11644);
or U13245 (N_13245,N_11942,N_8524);
and U13246 (N_13246,N_10729,N_9478);
or U13247 (N_13247,N_9405,N_9972);
xor U13248 (N_13248,N_11546,N_11204);
and U13249 (N_13249,N_8471,N_9559);
and U13250 (N_13250,N_8169,N_10819);
xnor U13251 (N_13251,N_10441,N_11826);
and U13252 (N_13252,N_11502,N_8990);
xor U13253 (N_13253,N_10678,N_11953);
xnor U13254 (N_13254,N_10411,N_8861);
or U13255 (N_13255,N_8241,N_8429);
xnor U13256 (N_13256,N_11448,N_9322);
or U13257 (N_13257,N_10204,N_10163);
nor U13258 (N_13258,N_11998,N_9576);
or U13259 (N_13259,N_10412,N_8646);
xnor U13260 (N_13260,N_8818,N_8344);
nand U13261 (N_13261,N_9976,N_9599);
and U13262 (N_13262,N_10890,N_10158);
and U13263 (N_13263,N_11637,N_11977);
xnor U13264 (N_13264,N_9381,N_8886);
nor U13265 (N_13265,N_9831,N_8420);
nor U13266 (N_13266,N_9948,N_11846);
xnor U13267 (N_13267,N_10373,N_8049);
nor U13268 (N_13268,N_11700,N_8246);
nor U13269 (N_13269,N_10860,N_9068);
nand U13270 (N_13270,N_8956,N_11765);
nand U13271 (N_13271,N_11926,N_10539);
or U13272 (N_13272,N_9179,N_9685);
or U13273 (N_13273,N_10467,N_11922);
and U13274 (N_13274,N_8878,N_9258);
nand U13275 (N_13275,N_11636,N_11296);
or U13276 (N_13276,N_11986,N_11270);
or U13277 (N_13277,N_8326,N_11503);
xor U13278 (N_13278,N_11271,N_8340);
xnor U13279 (N_13279,N_8357,N_10934);
nand U13280 (N_13280,N_9751,N_9864);
nand U13281 (N_13281,N_11741,N_9679);
nor U13282 (N_13282,N_10256,N_11806);
xor U13283 (N_13283,N_9531,N_9647);
and U13284 (N_13284,N_11933,N_9923);
or U13285 (N_13285,N_8706,N_9611);
nand U13286 (N_13286,N_10922,N_10709);
and U13287 (N_13287,N_8847,N_10156);
and U13288 (N_13288,N_9829,N_9410);
xnor U13289 (N_13289,N_10917,N_10305);
or U13290 (N_13290,N_10550,N_10112);
and U13291 (N_13291,N_10125,N_9347);
nor U13292 (N_13292,N_9879,N_10895);
nor U13293 (N_13293,N_11802,N_10304);
or U13294 (N_13294,N_11415,N_9585);
nand U13295 (N_13295,N_9680,N_11872);
nand U13296 (N_13296,N_11287,N_10309);
and U13297 (N_13297,N_11085,N_8789);
and U13298 (N_13298,N_11320,N_11095);
nand U13299 (N_13299,N_11647,N_9082);
nor U13300 (N_13300,N_10686,N_9601);
nor U13301 (N_13301,N_11129,N_8806);
nand U13302 (N_13302,N_10946,N_9494);
nor U13303 (N_13303,N_10340,N_9413);
or U13304 (N_13304,N_9703,N_8906);
nor U13305 (N_13305,N_10271,N_10555);
and U13306 (N_13306,N_11751,N_11378);
or U13307 (N_13307,N_11593,N_9793);
or U13308 (N_13308,N_8463,N_8066);
and U13309 (N_13309,N_8324,N_9250);
and U13310 (N_13310,N_8831,N_10873);
and U13311 (N_13311,N_10335,N_10343);
nor U13312 (N_13312,N_10350,N_10005);
or U13313 (N_13313,N_10049,N_8682);
nor U13314 (N_13314,N_9335,N_8585);
nor U13315 (N_13315,N_11762,N_10067);
or U13316 (N_13316,N_8590,N_11439);
nor U13317 (N_13317,N_10896,N_11985);
xor U13318 (N_13318,N_9568,N_10667);
and U13319 (N_13319,N_11693,N_9741);
nand U13320 (N_13320,N_11948,N_11034);
nor U13321 (N_13321,N_11541,N_8151);
or U13322 (N_13322,N_9072,N_11188);
or U13323 (N_13323,N_11510,N_11627);
xnor U13324 (N_13324,N_11473,N_11808);
nand U13325 (N_13325,N_9619,N_10566);
xnor U13326 (N_13326,N_8221,N_11410);
nor U13327 (N_13327,N_8071,N_11051);
or U13328 (N_13328,N_8583,N_10835);
nor U13329 (N_13329,N_10806,N_9284);
xnor U13330 (N_13330,N_11515,N_9155);
or U13331 (N_13331,N_8144,N_10190);
and U13332 (N_13332,N_9775,N_9440);
nor U13333 (N_13333,N_9798,N_8562);
nand U13334 (N_13334,N_11252,N_9264);
and U13335 (N_13335,N_11661,N_10086);
and U13336 (N_13336,N_11875,N_11670);
nand U13337 (N_13337,N_8771,N_9667);
nor U13338 (N_13338,N_8177,N_9895);
xor U13339 (N_13339,N_11662,N_11918);
and U13340 (N_13340,N_11965,N_9223);
and U13341 (N_13341,N_8390,N_9103);
or U13342 (N_13342,N_10284,N_8807);
xnor U13343 (N_13343,N_8464,N_9220);
and U13344 (N_13344,N_8623,N_11657);
nor U13345 (N_13345,N_9691,N_8421);
nand U13346 (N_13346,N_11176,N_8749);
xnor U13347 (N_13347,N_9769,N_9587);
xnor U13348 (N_13348,N_11614,N_9814);
and U13349 (N_13349,N_8255,N_8160);
nor U13350 (N_13350,N_11984,N_8042);
and U13351 (N_13351,N_8936,N_9658);
nand U13352 (N_13352,N_9304,N_11021);
or U13353 (N_13353,N_8875,N_8119);
and U13354 (N_13354,N_11412,N_9401);
xor U13355 (N_13355,N_9001,N_10072);
nor U13356 (N_13356,N_8021,N_11969);
nor U13357 (N_13357,N_9017,N_8796);
and U13358 (N_13358,N_10295,N_9031);
nor U13359 (N_13359,N_10219,N_10784);
or U13360 (N_13360,N_9107,N_11222);
nand U13361 (N_13361,N_11558,N_8274);
nand U13362 (N_13362,N_9309,N_10126);
or U13363 (N_13363,N_8603,N_11783);
nand U13364 (N_13364,N_11649,N_9934);
xnor U13365 (N_13365,N_10821,N_9690);
nor U13366 (N_13366,N_9903,N_8801);
and U13367 (N_13367,N_8321,N_10702);
nand U13368 (N_13368,N_10366,N_9367);
nand U13369 (N_13369,N_8170,N_11334);
and U13370 (N_13370,N_10251,N_10391);
and U13371 (N_13371,N_9191,N_8031);
or U13372 (N_13372,N_8338,N_9771);
or U13373 (N_13373,N_11333,N_8991);
nand U13374 (N_13374,N_10775,N_8330);
and U13375 (N_13375,N_9501,N_11837);
nand U13376 (N_13376,N_9764,N_11914);
and U13377 (N_13377,N_8834,N_8709);
nand U13378 (N_13378,N_9502,N_8679);
or U13379 (N_13379,N_8288,N_9498);
nand U13380 (N_13380,N_11612,N_9548);
xor U13381 (N_13381,N_8763,N_10186);
and U13382 (N_13382,N_9240,N_9400);
xnor U13383 (N_13383,N_11375,N_9452);
and U13384 (N_13384,N_11777,N_11418);
and U13385 (N_13385,N_11763,N_10243);
nand U13386 (N_13386,N_9421,N_11254);
and U13387 (N_13387,N_11838,N_9987);
nand U13388 (N_13388,N_10893,N_8187);
and U13389 (N_13389,N_11891,N_11909);
and U13390 (N_13390,N_8511,N_11449);
xor U13391 (N_13391,N_10766,N_9033);
nor U13392 (N_13392,N_9839,N_8925);
nand U13393 (N_13393,N_8052,N_8940);
and U13394 (N_13394,N_10571,N_10333);
nor U13395 (N_13395,N_11508,N_11376);
or U13396 (N_13396,N_9971,N_11445);
and U13397 (N_13397,N_9402,N_11584);
xnor U13398 (N_13398,N_10606,N_11770);
nand U13399 (N_13399,N_8578,N_9655);
and U13400 (N_13400,N_9722,N_8106);
and U13401 (N_13401,N_11626,N_8014);
and U13402 (N_13402,N_8803,N_8277);
and U13403 (N_13403,N_10051,N_9904);
nor U13404 (N_13404,N_8762,N_10968);
xnor U13405 (N_13405,N_11444,N_11260);
nand U13406 (N_13406,N_10990,N_9147);
or U13407 (N_13407,N_8802,N_8405);
nor U13408 (N_13408,N_9570,N_10698);
xor U13409 (N_13409,N_8240,N_10984);
xor U13410 (N_13410,N_9509,N_11209);
or U13411 (N_13411,N_10044,N_9912);
or U13412 (N_13412,N_11354,N_8926);
or U13413 (N_13413,N_9249,N_8983);
and U13414 (N_13414,N_10184,N_9185);
and U13415 (N_13415,N_8764,N_9600);
nor U13416 (N_13416,N_9558,N_10476);
or U13417 (N_13417,N_8167,N_11310);
nand U13418 (N_13418,N_10444,N_10195);
and U13419 (N_13419,N_11374,N_8224);
or U13420 (N_13420,N_9156,N_9273);
xnor U13421 (N_13421,N_9885,N_9311);
or U13422 (N_13422,N_9999,N_10367);
or U13423 (N_13423,N_9178,N_10755);
xor U13424 (N_13424,N_11411,N_10022);
xnor U13425 (N_13425,N_9791,N_11961);
nand U13426 (N_13426,N_10480,N_10012);
or U13427 (N_13427,N_11555,N_8320);
nand U13428 (N_13428,N_11995,N_10622);
or U13429 (N_13429,N_10749,N_10378);
or U13430 (N_13430,N_8766,N_11639);
xor U13431 (N_13431,N_10426,N_10336);
xor U13432 (N_13432,N_10715,N_9416);
or U13433 (N_13433,N_10089,N_11471);
and U13434 (N_13434,N_8805,N_8349);
nand U13435 (N_13435,N_10874,N_8892);
nand U13436 (N_13436,N_11045,N_10614);
and U13437 (N_13437,N_11964,N_9216);
nor U13438 (N_13438,N_11387,N_10644);
nand U13439 (N_13439,N_9313,N_9192);
or U13440 (N_13440,N_9049,N_9977);
xnor U13441 (N_13441,N_10731,N_9995);
and U13442 (N_13442,N_8904,N_11717);
xnor U13443 (N_13443,N_9363,N_11987);
nand U13444 (N_13444,N_11242,N_8555);
and U13445 (N_13445,N_8137,N_11478);
nor U13446 (N_13446,N_9889,N_11682);
and U13447 (N_13447,N_10421,N_11561);
or U13448 (N_13448,N_11562,N_8935);
or U13449 (N_13449,N_11608,N_8194);
nand U13450 (N_13450,N_10501,N_11026);
nand U13451 (N_13451,N_9280,N_9854);
nand U13452 (N_13452,N_10457,N_8291);
xnor U13453 (N_13453,N_9530,N_8999);
or U13454 (N_13454,N_10626,N_11117);
xnor U13455 (N_13455,N_9979,N_9649);
nand U13456 (N_13456,N_9597,N_11687);
xor U13457 (N_13457,N_8527,N_8317);
nand U13458 (N_13458,N_8863,N_9362);
or U13459 (N_13459,N_8423,N_8190);
or U13460 (N_13460,N_8544,N_10359);
and U13461 (N_13461,N_11087,N_11583);
or U13462 (N_13462,N_9697,N_11207);
xor U13463 (N_13463,N_8479,N_10084);
or U13464 (N_13464,N_11850,N_8228);
nand U13465 (N_13465,N_8873,N_9190);
nor U13466 (N_13466,N_9749,N_11213);
xnor U13467 (N_13467,N_11652,N_8436);
xor U13468 (N_13468,N_11537,N_8468);
and U13469 (N_13469,N_8077,N_8345);
nor U13470 (N_13470,N_8735,N_10552);
nand U13471 (N_13471,N_8076,N_8758);
nand U13472 (N_13472,N_11458,N_10490);
or U13473 (N_13473,N_8263,N_8433);
or U13474 (N_13474,N_8495,N_10153);
or U13475 (N_13475,N_9956,N_9225);
and U13476 (N_13476,N_11466,N_9684);
nor U13477 (N_13477,N_9888,N_9899);
xor U13478 (N_13478,N_10312,N_9907);
or U13479 (N_13479,N_8888,N_11128);
and U13480 (N_13480,N_8176,N_11747);
nor U13481 (N_13481,N_11248,N_9951);
nand U13482 (N_13482,N_9730,N_11245);
nand U13483 (N_13483,N_9562,N_11819);
and U13484 (N_13484,N_10280,N_10870);
nor U13485 (N_13485,N_10446,N_11261);
or U13486 (N_13486,N_10148,N_11674);
xnor U13487 (N_13487,N_10006,N_11660);
nor U13488 (N_13488,N_11553,N_9254);
xnor U13489 (N_13489,N_8656,N_8219);
nand U13490 (N_13490,N_9464,N_11237);
or U13491 (N_13491,N_9108,N_8614);
or U13492 (N_13492,N_11709,N_8612);
xor U13493 (N_13493,N_11363,N_8626);
or U13494 (N_13494,N_8775,N_9635);
nand U13495 (N_13495,N_8879,N_8318);
or U13496 (N_13496,N_9318,N_10751);
or U13497 (N_13497,N_11455,N_9080);
nand U13498 (N_13498,N_8450,N_11366);
xnor U13499 (N_13499,N_9289,N_10802);
and U13500 (N_13500,N_10385,N_10615);
and U13501 (N_13501,N_11040,N_11304);
and U13502 (N_13502,N_9526,N_10796);
nand U13503 (N_13503,N_10399,N_8403);
or U13504 (N_13504,N_8281,N_8997);
xnor U13505 (N_13505,N_9994,N_8641);
nand U13506 (N_13506,N_11078,N_11621);
and U13507 (N_13507,N_8356,N_11179);
or U13508 (N_13508,N_10537,N_11268);
or U13509 (N_13509,N_11383,N_10136);
and U13510 (N_13510,N_8347,N_11409);
or U13511 (N_13511,N_11061,N_11579);
nor U13512 (N_13512,N_10240,N_11147);
and U13513 (N_13513,N_9083,N_10785);
and U13514 (N_13514,N_10183,N_11685);
nor U13515 (N_13515,N_10681,N_11338);
nand U13516 (N_13516,N_10789,N_9808);
nor U13517 (N_13517,N_9966,N_11115);
or U13518 (N_13518,N_10418,N_11854);
nand U13519 (N_13519,N_11930,N_11782);
or U13520 (N_13520,N_10409,N_8739);
xnor U13521 (N_13521,N_11293,N_9743);
nand U13522 (N_13522,N_8897,N_11029);
xor U13523 (N_13523,N_9922,N_10876);
xor U13524 (N_13524,N_8234,N_8125);
nand U13525 (N_13525,N_11214,N_10493);
or U13526 (N_13526,N_11712,N_11368);
and U13527 (N_13527,N_8752,N_10711);
nand U13528 (N_13528,N_8251,N_10034);
nor U13529 (N_13529,N_11438,N_9770);
xor U13530 (N_13530,N_10191,N_10609);
or U13531 (N_13531,N_9211,N_8085);
nor U13532 (N_13532,N_11390,N_11377);
and U13533 (N_13533,N_8154,N_10790);
nor U13534 (N_13534,N_10565,N_10325);
nand U13535 (N_13535,N_9434,N_10983);
or U13536 (N_13536,N_9161,N_9221);
and U13537 (N_13537,N_10676,N_11276);
nor U13538 (N_13538,N_10824,N_9274);
nor U13539 (N_13539,N_11959,N_10394);
xor U13540 (N_13540,N_10759,N_8315);
nand U13541 (N_13541,N_10427,N_8657);
nor U13542 (N_13542,N_10023,N_8470);
or U13543 (N_13543,N_9061,N_10595);
and U13544 (N_13544,N_8643,N_8719);
or U13545 (N_13545,N_9026,N_11193);
and U13546 (N_13546,N_11887,N_10692);
and U13547 (N_13547,N_10659,N_8600);
nand U13548 (N_13548,N_8856,N_8648);
xor U13549 (N_13549,N_10561,N_9705);
nor U13550 (N_13550,N_11075,N_9595);
xor U13551 (N_13551,N_10810,N_10518);
and U13552 (N_13552,N_9534,N_9206);
and U13553 (N_13553,N_11723,N_8694);
or U13554 (N_13554,N_8259,N_11939);
nor U13555 (N_13555,N_10344,N_9299);
nand U13556 (N_13556,N_10015,N_8381);
nand U13557 (N_13557,N_11894,N_11425);
nor U13558 (N_13558,N_8943,N_9767);
or U13559 (N_13559,N_9529,N_10801);
xor U13560 (N_13560,N_10466,N_11307);
xnor U13561 (N_13561,N_10066,N_8269);
and U13562 (N_13562,N_8243,N_11931);
and U13563 (N_13563,N_8565,N_9039);
nor U13564 (N_13564,N_8534,N_10482);
xor U13565 (N_13565,N_11286,N_11265);
xnor U13566 (N_13566,N_9004,N_10602);
xor U13567 (N_13567,N_10323,N_8989);
xnor U13568 (N_13568,N_8414,N_8393);
nand U13569 (N_13569,N_8040,N_10596);
nand U13570 (N_13570,N_10130,N_11004);
or U13571 (N_13571,N_8670,N_8914);
and U13572 (N_13572,N_9283,N_9518);
xnor U13573 (N_13573,N_8707,N_11548);
xor U13574 (N_13574,N_10150,N_10891);
nand U13575 (N_13575,N_11677,N_8131);
xor U13576 (N_13576,N_8020,N_11532);
nand U13577 (N_13577,N_10866,N_10327);
nand U13578 (N_13578,N_8441,N_10648);
and U13579 (N_13579,N_11775,N_10110);
nor U13580 (N_13580,N_8696,N_10769);
or U13581 (N_13581,N_8408,N_11313);
or U13582 (N_13582,N_10401,N_11814);
nand U13583 (N_13583,N_9174,N_8785);
or U13584 (N_13584,N_11233,N_8503);
nand U13585 (N_13585,N_8920,N_10881);
or U13586 (N_13586,N_11391,N_10448);
and U13587 (N_13587,N_11119,N_9557);
nand U13588 (N_13588,N_8045,N_9606);
nand U13589 (N_13589,N_11240,N_11949);
nor U13590 (N_13590,N_11241,N_10970);
xor U13591 (N_13591,N_11250,N_8970);
or U13592 (N_13592,N_11980,N_9772);
nor U13593 (N_13593,N_9024,N_10146);
xnor U13594 (N_13594,N_11024,N_9202);
or U13595 (N_13595,N_11549,N_10311);
nor U13596 (N_13596,N_9005,N_8974);
nor U13597 (N_13597,N_8619,N_11362);
and U13598 (N_13598,N_8577,N_9656);
nor U13599 (N_13599,N_9279,N_11156);
and U13600 (N_13600,N_8208,N_10646);
or U13601 (N_13601,N_9484,N_10020);
nand U13602 (N_13602,N_8497,N_10076);
or U13603 (N_13603,N_8313,N_10414);
nor U13604 (N_13604,N_11522,N_9208);
nand U13605 (N_13605,N_8216,N_9018);
or U13606 (N_13606,N_10827,N_8923);
nand U13607 (N_13607,N_8353,N_10211);
nand U13608 (N_13608,N_10422,N_9207);
or U13609 (N_13609,N_10193,N_11249);
xor U13610 (N_13610,N_9817,N_10965);
or U13611 (N_13611,N_10897,N_9627);
nor U13612 (N_13612,N_11032,N_9436);
xor U13613 (N_13613,N_8309,N_11688);
and U13614 (N_13614,N_10290,N_11025);
and U13615 (N_13615,N_10734,N_9500);
xor U13616 (N_13616,N_11224,N_8445);
and U13617 (N_13617,N_8622,N_8609);
nand U13618 (N_13618,N_10004,N_9113);
or U13619 (N_13619,N_11441,N_8000);
or U13620 (N_13620,N_10532,N_10348);
and U13621 (N_13621,N_9836,N_8370);
xor U13622 (N_13622,N_8011,N_9383);
and U13623 (N_13623,N_8493,N_9868);
xor U13624 (N_13624,N_10046,N_9867);
xnor U13625 (N_13625,N_9603,N_8173);
xor U13626 (N_13626,N_10007,N_10690);
xor U13627 (N_13627,N_8946,N_9666);
and U13628 (N_13628,N_8916,N_10988);
and U13629 (N_13629,N_8480,N_11422);
xnor U13630 (N_13630,N_11897,N_9073);
or U13631 (N_13631,N_10869,N_9006);
nand U13632 (N_13632,N_8576,N_10270);
and U13633 (N_13633,N_10347,N_10636);
and U13634 (N_13634,N_10292,N_9985);
nand U13635 (N_13635,N_10175,N_10380);
and U13636 (N_13636,N_8105,N_11054);
nor U13637 (N_13637,N_9878,N_10625);
and U13638 (N_13638,N_8542,N_9936);
and U13639 (N_13639,N_8025,N_10429);
or U13640 (N_13640,N_9642,N_10400);
or U13641 (N_13641,N_10511,N_8620);
and U13642 (N_13642,N_8992,N_11149);
nor U13643 (N_13643,N_9731,N_11405);
or U13644 (N_13644,N_11223,N_10885);
nor U13645 (N_13645,N_11916,N_10725);
nor U13646 (N_13646,N_10582,N_11253);
and U13647 (N_13647,N_10376,N_11480);
nand U13648 (N_13648,N_11595,N_11351);
nand U13649 (N_13649,N_10914,N_11790);
and U13650 (N_13650,N_10813,N_10884);
or U13651 (N_13651,N_11501,N_9136);
xnor U13652 (N_13652,N_10106,N_8635);
and U13653 (N_13653,N_8519,N_11322);
nand U13654 (N_13654,N_10778,N_11634);
and U13655 (N_13655,N_10793,N_11098);
xnor U13656 (N_13656,N_11486,N_9554);
xor U13657 (N_13657,N_9780,N_8253);
or U13658 (N_13658,N_10553,N_10956);
xnor U13659 (N_13659,N_11017,N_10607);
nand U13660 (N_13660,N_10138,N_11067);
and U13661 (N_13661,N_10289,N_11618);
or U13662 (N_13662,N_9399,N_11867);
nor U13663 (N_13663,N_9917,N_10264);
and U13664 (N_13664,N_11216,N_9887);
nand U13665 (N_13665,N_10206,N_9695);
nand U13666 (N_13666,N_9324,N_11559);
nand U13667 (N_13667,N_8951,N_10105);
nor U13668 (N_13668,N_10954,N_10018);
nand U13669 (N_13669,N_11099,N_11920);
and U13670 (N_13670,N_9260,N_8964);
xor U13671 (N_13671,N_10907,N_9379);
nand U13672 (N_13672,N_10334,N_9409);
xor U13673 (N_13673,N_10030,N_10117);
nor U13674 (N_13674,N_9998,N_9035);
nor U13675 (N_13675,N_9165,N_8931);
and U13676 (N_13676,N_11898,N_10257);
and U13677 (N_13677,N_10800,N_8553);
nor U13678 (N_13678,N_10551,N_11590);
nor U13679 (N_13679,N_9488,N_9650);
xnor U13680 (N_13680,N_9669,N_9343);
nand U13681 (N_13681,N_11592,N_10598);
and U13682 (N_13682,N_8822,N_9732);
or U13683 (N_13683,N_10413,N_8473);
and U13684 (N_13684,N_8292,N_11967);
nor U13685 (N_13685,N_10577,N_11825);
xor U13686 (N_13686,N_10133,N_10631);
xnor U13687 (N_13687,N_10486,N_8064);
or U13688 (N_13688,N_10969,N_8937);
xor U13689 (N_13689,N_9218,N_9348);
and U13690 (N_13690,N_8273,N_9089);
nand U13691 (N_13691,N_11125,N_9074);
xnor U13692 (N_13692,N_11134,N_8095);
and U13693 (N_13693,N_10070,N_10665);
and U13694 (N_13694,N_9259,N_8409);
or U13695 (N_13695,N_8733,N_11337);
nor U13696 (N_13696,N_8547,N_11571);
xor U13697 (N_13697,N_10469,N_9129);
nand U13698 (N_13698,N_11572,N_9662);
nor U13699 (N_13699,N_8704,N_8962);
nor U13700 (N_13700,N_11055,N_9415);
xnor U13701 (N_13701,N_9687,N_9196);
nor U13702 (N_13702,N_9365,N_9317);
and U13703 (N_13703,N_11896,N_9219);
and U13704 (N_13704,N_11341,N_10261);
and U13705 (N_13705,N_11141,N_11113);
nand U13706 (N_13706,N_10306,N_11192);
nor U13707 (N_13707,N_10477,N_8549);
and U13708 (N_13708,N_10324,N_8440);
or U13709 (N_13709,N_8097,N_8559);
or U13710 (N_13710,N_8328,N_10713);
xnor U13711 (N_13711,N_9825,N_10583);
and U13712 (N_13712,N_10387,N_10500);
or U13713 (N_13713,N_9796,N_8325);
nand U13714 (N_13714,N_11692,N_8533);
and U13715 (N_13715,N_11397,N_11275);
xnor U13716 (N_13716,N_8688,N_10124);
xor U13717 (N_13717,N_8466,N_10389);
xnor U13718 (N_13718,N_8139,N_8475);
nand U13719 (N_13719,N_8680,N_8760);
xnor U13720 (N_13720,N_9574,N_9341);
or U13721 (N_13721,N_11970,N_8459);
nand U13722 (N_13722,N_8406,N_8568);
and U13723 (N_13723,N_11870,N_10522);
nand U13724 (N_13724,N_10899,N_8211);
nand U13725 (N_13725,N_8649,N_8322);
nand U13726 (N_13726,N_10909,N_10604);
and U13727 (N_13727,N_8227,N_10319);
and U13728 (N_13728,N_8192,N_9133);
nand U13729 (N_13729,N_8911,N_9408);
nor U13730 (N_13730,N_9459,N_8628);
nand U13731 (N_13731,N_11516,N_11103);
or U13732 (N_13732,N_11699,N_9360);
nor U13733 (N_13733,N_11514,N_9858);
or U13734 (N_13734,N_8339,N_8371);
and U13735 (N_13735,N_9398,N_8798);
xnor U13736 (N_13736,N_8029,N_11489);
nor U13737 (N_13737,N_11882,N_8987);
nand U13738 (N_13738,N_11461,N_8677);
nand U13739 (N_13739,N_8217,N_8895);
or U13740 (N_13740,N_8044,N_9643);
and U13741 (N_13741,N_8751,N_10710);
and U13742 (N_13742,N_11702,N_9674);
or U13743 (N_13743,N_9099,N_10777);
nand U13744 (N_13744,N_8266,N_9504);
nand U13745 (N_13745,N_11574,N_8644);
nand U13746 (N_13746,N_11563,N_9336);
and U13747 (N_13747,N_11228,N_9349);
or U13748 (N_13748,N_9712,N_9389);
xor U13749 (N_13749,N_11539,N_9009);
and U13750 (N_13750,N_11900,N_11277);
and U13751 (N_13751,N_11865,N_11169);
and U13752 (N_13752,N_11330,N_8039);
and U13753 (N_13753,N_11816,N_11720);
xnor U13754 (N_13754,N_10831,N_10976);
or U13755 (N_13755,N_8027,N_8579);
or U13756 (N_13756,N_8197,N_9633);
nor U13757 (N_13757,N_8632,N_9180);
nand U13758 (N_13758,N_8690,N_10704);
and U13759 (N_13759,N_8726,N_8443);
nor U13760 (N_13760,N_11135,N_9713);
or U13761 (N_13761,N_11526,N_9406);
nand U13762 (N_13762,N_10245,N_10689);
xnor U13763 (N_13763,N_10630,N_9542);
or U13764 (N_13764,N_9268,N_9456);
nand U13765 (N_13765,N_9256,N_8157);
nor U13766 (N_13766,N_11311,N_11936);
or U13767 (N_13767,N_10798,N_9376);
nand U13768 (N_13768,N_8081,N_9088);
or U13769 (N_13769,N_8988,N_11435);
and U13770 (N_13770,N_9411,N_8186);
and U13771 (N_13771,N_11616,N_10597);
and U13772 (N_13772,N_11089,N_11978);
nand U13773 (N_13773,N_9866,N_9982);
nand U13774 (N_13774,N_11082,N_11780);
xor U13775 (N_13775,N_9950,N_10330);
nand U13776 (N_13776,N_9248,N_8182);
and U13777 (N_13777,N_8038,N_9532);
nor U13778 (N_13778,N_9081,N_9453);
and U13779 (N_13779,N_9677,N_11956);
nand U13780 (N_13780,N_9984,N_9043);
and U13781 (N_13781,N_10162,N_8581);
and U13782 (N_13782,N_10516,N_8535);
and U13783 (N_13783,N_11853,N_10997);
and U13784 (N_13784,N_10002,N_11492);
or U13785 (N_13785,N_8141,N_11996);
and U13786 (N_13786,N_11451,N_11923);
or U13787 (N_13787,N_10026,N_8557);
or U13788 (N_13788,N_9541,N_9779);
xor U13789 (N_13789,N_9852,N_11472);
nor U13790 (N_13790,N_11759,N_9551);
xnor U13791 (N_13791,N_9148,N_10390);
xor U13792 (N_13792,N_9119,N_9758);
nor U13793 (N_13793,N_9475,N_9270);
nor U13794 (N_13794,N_9159,N_8075);
xnor U13795 (N_13795,N_10104,N_8457);
xnor U13796 (N_13796,N_8845,N_11876);
nand U13797 (N_13797,N_11713,N_8929);
nor U13798 (N_13798,N_8896,N_10668);
nand U13799 (N_13799,N_9138,N_8842);
or U13800 (N_13800,N_9443,N_8348);
nand U13801 (N_13801,N_9949,N_10369);
nor U13802 (N_13802,N_11300,N_8500);
nand U13803 (N_13803,N_10196,N_10575);
xor U13804 (N_13804,N_11165,N_8100);
nand U13805 (N_13805,N_9832,N_10852);
or U13806 (N_13806,N_11523,N_9227);
nand U13807 (N_13807,N_10370,N_9134);
nand U13808 (N_13808,N_11394,N_11575);
xnor U13809 (N_13809,N_8265,N_11072);
xnor U13810 (N_13810,N_8810,N_8797);
or U13811 (N_13811,N_11084,N_11447);
nand U13812 (N_13812,N_11531,N_11773);
and U13813 (N_13813,N_9446,N_10404);
nand U13814 (N_13814,N_11628,N_8615);
and U13815 (N_13815,N_9590,N_11912);
and U13816 (N_13816,N_9125,N_9391);
nor U13817 (N_13817,N_8558,N_10805);
and U13818 (N_13818,N_9295,N_11077);
xor U13819 (N_13819,N_8486,N_11648);
nor U13820 (N_13820,N_9788,N_11758);
xnor U13821 (N_13821,N_8395,N_11047);
nand U13822 (N_13822,N_8756,N_9358);
xor U13823 (N_13823,N_11150,N_10491);
nor U13824 (N_13824,N_11443,N_9589);
nand U13825 (N_13825,N_8094,N_8629);
nand U13826 (N_13826,N_9802,N_8835);
and U13827 (N_13827,N_8487,N_11057);
xor U13828 (N_13828,N_8113,N_10718);
nor U13829 (N_13829,N_11810,N_11744);
nor U13830 (N_13830,N_9883,N_10618);
nor U13831 (N_13831,N_8505,N_9639);
nand U13832 (N_13832,N_10594,N_11071);
xnor U13833 (N_13833,N_8799,N_11225);
or U13834 (N_13834,N_11340,N_10682);
xnor U13835 (N_13835,N_10139,N_10888);
nand U13836 (N_13836,N_11011,N_11879);
xor U13837 (N_13837,N_9124,N_11482);
nor U13838 (N_13838,N_10337,N_11196);
nand U13839 (N_13839,N_8476,N_8825);
and U13840 (N_13840,N_10905,N_11902);
xnor U13841 (N_13841,N_9090,N_8392);
and U13842 (N_13842,N_8539,N_10265);
and U13843 (N_13843,N_8195,N_10505);
nor U13844 (N_13844,N_10904,N_9944);
or U13845 (N_13845,N_9022,N_10019);
or U13846 (N_13846,N_10151,N_8375);
nand U13847 (N_13847,N_10898,N_9315);
nor U13848 (N_13848,N_10453,N_8700);
nor U13849 (N_13849,N_10254,N_10484);
or U13850 (N_13850,N_9577,N_11136);
xnor U13851 (N_13851,N_9620,N_10328);
and U13852 (N_13852,N_11371,N_10642);
nor U13853 (N_13853,N_11166,N_11552);
xnor U13854 (N_13854,N_9213,N_10215);
nand U13855 (N_13855,N_8425,N_10717);
nand U13856 (N_13856,N_10037,N_10231);
xnor U13857 (N_13857,N_9079,N_8138);
nor U13858 (N_13858,N_10194,N_9947);
or U13859 (N_13859,N_9660,N_8023);
nand U13860 (N_13860,N_10454,N_9455);
or U13861 (N_13861,N_10807,N_9822);
or U13862 (N_13862,N_9980,N_9750);
nand U13863 (N_13863,N_8655,N_10302);
xor U13864 (N_13864,N_11133,N_9344);
nor U13865 (N_13865,N_8413,N_8467);
nor U13866 (N_13866,N_8481,N_8816);
and U13867 (N_13867,N_10556,N_10180);
nor U13868 (N_13868,N_9609,N_9300);
nor U13869 (N_13869,N_8400,N_10029);
or U13870 (N_13870,N_10863,N_11291);
nand U13871 (N_13871,N_8638,N_9404);
nand U13872 (N_13872,N_9154,N_9783);
nand U13873 (N_13873,N_9584,N_10269);
nand U13874 (N_13874,N_10531,N_10739);
xor U13875 (N_13875,N_11520,N_11772);
or U13876 (N_13876,N_10237,N_8472);
xnor U13877 (N_13877,N_10203,N_9686);
xor U13878 (N_13878,N_10794,N_9070);
nand U13879 (N_13879,N_9163,N_8303);
xor U13880 (N_13880,N_11211,N_10829);
nand U13881 (N_13881,N_10321,N_8854);
xnor U13882 (N_13882,N_8820,N_8091);
xnor U13883 (N_13883,N_10574,N_11588);
nand U13884 (N_13884,N_9441,N_8866);
nand U13885 (N_13885,N_8817,N_10580);
nand U13886 (N_13886,N_8826,N_9993);
or U13887 (N_13887,N_8894,N_8006);
nor U13888 (N_13888,N_11069,N_11460);
nand U13889 (N_13889,N_11606,N_8971);
and U13890 (N_13890,N_10377,N_8163);
xor U13891 (N_13891,N_10814,N_9010);
nor U13892 (N_13892,N_10383,N_11791);
nor U13893 (N_13893,N_11556,N_10640);
nor U13894 (N_13894,N_9753,N_8271);
nand U13895 (N_13895,N_9636,N_11358);
nor U13896 (N_13896,N_8223,N_9474);
nor U13897 (N_13897,N_8808,N_10509);
nand U13898 (N_13898,N_8012,N_8460);
nand U13899 (N_13899,N_11372,N_11990);
nor U13900 (N_13900,N_9373,N_10329);
nor U13901 (N_13901,N_10544,N_10285);
or U13902 (N_13902,N_9563,N_11105);
nand U13903 (N_13903,N_10455,N_11309);
xor U13904 (N_13904,N_10363,N_9918);
nand U13905 (N_13905,N_8362,N_11567);
xor U13906 (N_13906,N_10776,N_9444);
or U13907 (N_13907,N_8017,N_8793);
or U13908 (N_13908,N_9646,N_11740);
nand U13909 (N_13909,N_10024,N_10746);
and U13910 (N_13910,N_8065,N_11705);
nand U13911 (N_13911,N_9493,N_11536);
nor U13912 (N_13912,N_11044,N_8465);
and U13913 (N_13913,N_8041,N_8977);
nor U13914 (N_13914,N_8965,N_10536);
and U13915 (N_13915,N_11138,N_11767);
xor U13916 (N_13916,N_9171,N_11730);
and U13917 (N_13917,N_11576,N_11504);
and U13918 (N_13918,N_8179,N_10568);
nand U13919 (N_13919,N_10428,N_8215);
nand U13920 (N_13920,N_10735,N_11005);
xnor U13921 (N_13921,N_11401,N_11496);
and U13922 (N_13922,N_10959,N_9047);
nand U13923 (N_13923,N_9432,N_11190);
xor U13924 (N_13924,N_8633,N_11513);
nor U13925 (N_13925,N_9442,N_10795);
xor U13926 (N_13926,N_8938,N_10388);
xor U13927 (N_13927,N_11111,N_11908);
nor U13928 (N_13928,N_10593,N_9238);
nor U13929 (N_13929,N_9150,N_11049);
nand U13930 (N_13930,N_10062,N_8729);
nand U13931 (N_13931,N_8772,N_9217);
and U13932 (N_13932,N_8037,N_11975);
xnor U13933 (N_13933,N_9556,N_10918);
or U13934 (N_13934,N_11704,N_9346);
or U13935 (N_13935,N_11973,N_11088);
xor U13936 (N_13936,N_10108,N_8202);
and U13937 (N_13937,N_10042,N_9721);
nand U13938 (N_13938,N_8720,N_9990);
nor U13939 (N_13939,N_9263,N_11463);
and U13940 (N_13940,N_9181,N_8019);
or U13941 (N_13941,N_9055,N_10065);
xor U13942 (N_13942,N_11355,N_11714);
nand U13943 (N_13943,N_8525,N_8769);
and U13944 (N_13944,N_9396,N_9307);
or U13945 (N_13945,N_10345,N_9863);
nand U13946 (N_13946,N_8004,N_11694);
nand U13947 (N_13947,N_9097,N_9628);
or U13948 (N_13948,N_10392,N_11753);
nor U13949 (N_13949,N_11038,N_10293);
and U13950 (N_13950,N_10828,N_9468);
xnor U13951 (N_13951,N_9844,N_9513);
nor U13952 (N_13952,N_9002,N_11474);
nand U13953 (N_13953,N_11601,N_10572);
and U13954 (N_13954,N_9194,N_8880);
and U13955 (N_13955,N_8063,N_8110);
nand U13956 (N_13956,N_9281,N_8034);
nand U13957 (N_13957,N_10073,N_11679);
nor U13958 (N_13958,N_8301,N_10384);
and U13959 (N_13959,N_9790,N_10403);
nor U13960 (N_13960,N_10314,N_8627);
xor U13961 (N_13961,N_9991,N_10830);
xor U13962 (N_13962,N_9623,N_9578);
or U13963 (N_13963,N_11315,N_11794);
and U13964 (N_13964,N_8710,N_9166);
xor U13965 (N_13965,N_10003,N_11008);
or U13966 (N_13966,N_11272,N_10770);
or U13967 (N_13967,N_9692,N_9575);
nor U13968 (N_13968,N_8788,N_9954);
nor U13969 (N_13969,N_8155,N_11877);
nand U13970 (N_13970,N_9257,N_10095);
nand U13971 (N_13971,N_9673,N_9189);
nor U13972 (N_13972,N_11743,N_8093);
nand U13973 (N_13973,N_8661,N_9130);
or U13974 (N_13974,N_9816,N_10119);
nor U13975 (N_13975,N_8088,N_8276);
nor U13976 (N_13976,N_10207,N_10938);
nor U13977 (N_13977,N_8712,N_9372);
xor U13978 (N_13978,N_9517,N_9414);
or U13979 (N_13979,N_11971,N_10016);
nor U13980 (N_13980,N_11611,N_11227);
or U13981 (N_13981,N_9975,N_8893);
nand U13982 (N_13982,N_8960,N_10762);
and U13983 (N_13983,N_11728,N_11206);
nor U13984 (N_13984,N_9555,N_8319);
nand U13985 (N_13985,N_10722,N_9164);
and U13986 (N_13986,N_10803,N_8908);
and U13987 (N_13987,N_10496,N_8430);
nand U13988 (N_13988,N_9457,N_8111);
nand U13989 (N_13989,N_9915,N_8950);
xnor U13990 (N_13990,N_11408,N_10864);
and U13991 (N_13991,N_10772,N_8554);
or U13992 (N_13992,N_11022,N_10691);
xnor U13993 (N_13993,N_9935,N_11698);
nor U13994 (N_13994,N_11086,N_10452);
nand U13995 (N_13995,N_8439,N_8852);
nand U13996 (N_13996,N_8876,N_8928);
xnor U13997 (N_13997,N_9310,N_8961);
and U13998 (N_13998,N_10096,N_10915);
nand U13999 (N_13999,N_10278,N_9127);
and U14000 (N_14000,N_10008,N_9068);
nor U14001 (N_14001,N_8747,N_11851);
and U14002 (N_14002,N_9080,N_11013);
and U14003 (N_14003,N_10189,N_10615);
or U14004 (N_14004,N_10717,N_8605);
xnor U14005 (N_14005,N_11394,N_9705);
nor U14006 (N_14006,N_11487,N_11192);
or U14007 (N_14007,N_10338,N_9944);
or U14008 (N_14008,N_8364,N_11201);
or U14009 (N_14009,N_8844,N_9226);
or U14010 (N_14010,N_10754,N_11529);
and U14011 (N_14011,N_8976,N_10428);
xor U14012 (N_14012,N_9893,N_9780);
nor U14013 (N_14013,N_10281,N_8220);
xor U14014 (N_14014,N_8353,N_11475);
nor U14015 (N_14015,N_10283,N_9576);
and U14016 (N_14016,N_8394,N_8170);
or U14017 (N_14017,N_8614,N_8961);
nor U14018 (N_14018,N_10300,N_8400);
nor U14019 (N_14019,N_10770,N_9491);
nor U14020 (N_14020,N_11226,N_9053);
or U14021 (N_14021,N_11969,N_9151);
xnor U14022 (N_14022,N_11169,N_9349);
nand U14023 (N_14023,N_8121,N_9199);
nand U14024 (N_14024,N_8148,N_8255);
xor U14025 (N_14025,N_10849,N_10745);
nand U14026 (N_14026,N_8240,N_11001);
nor U14027 (N_14027,N_10458,N_10434);
nand U14028 (N_14028,N_8584,N_11128);
or U14029 (N_14029,N_9855,N_10982);
or U14030 (N_14030,N_10986,N_8946);
nand U14031 (N_14031,N_9045,N_9338);
and U14032 (N_14032,N_8414,N_11932);
nor U14033 (N_14033,N_8235,N_10473);
nor U14034 (N_14034,N_8929,N_10163);
nor U14035 (N_14035,N_11547,N_11943);
nand U14036 (N_14036,N_8865,N_11823);
xnor U14037 (N_14037,N_11614,N_11044);
nand U14038 (N_14038,N_9743,N_9838);
or U14039 (N_14039,N_9959,N_11218);
nor U14040 (N_14040,N_9104,N_8905);
or U14041 (N_14041,N_8577,N_11152);
or U14042 (N_14042,N_10257,N_9198);
xor U14043 (N_14043,N_9041,N_9825);
nor U14044 (N_14044,N_8265,N_9351);
or U14045 (N_14045,N_8063,N_8126);
nand U14046 (N_14046,N_11477,N_10291);
or U14047 (N_14047,N_10075,N_11298);
or U14048 (N_14048,N_10543,N_11551);
xnor U14049 (N_14049,N_10620,N_11083);
nand U14050 (N_14050,N_9187,N_11007);
and U14051 (N_14051,N_10077,N_11905);
or U14052 (N_14052,N_11407,N_11318);
nor U14053 (N_14053,N_9706,N_8742);
xnor U14054 (N_14054,N_11919,N_9871);
nand U14055 (N_14055,N_9605,N_11200);
xnor U14056 (N_14056,N_8565,N_8985);
nand U14057 (N_14057,N_9155,N_11341);
and U14058 (N_14058,N_9670,N_11352);
xnor U14059 (N_14059,N_9511,N_9770);
and U14060 (N_14060,N_10957,N_11697);
nor U14061 (N_14061,N_10917,N_10074);
and U14062 (N_14062,N_9106,N_11067);
xor U14063 (N_14063,N_11238,N_11996);
and U14064 (N_14064,N_10764,N_9019);
xor U14065 (N_14065,N_10115,N_9492);
nand U14066 (N_14066,N_10439,N_8739);
and U14067 (N_14067,N_8503,N_9597);
nor U14068 (N_14068,N_11233,N_11696);
or U14069 (N_14069,N_8287,N_8916);
nor U14070 (N_14070,N_11423,N_11256);
and U14071 (N_14071,N_11223,N_11230);
nor U14072 (N_14072,N_10366,N_8280);
or U14073 (N_14073,N_10517,N_10864);
nand U14074 (N_14074,N_8288,N_10064);
nand U14075 (N_14075,N_9434,N_8365);
xnor U14076 (N_14076,N_9910,N_11342);
xor U14077 (N_14077,N_10840,N_9359);
or U14078 (N_14078,N_11585,N_11041);
xor U14079 (N_14079,N_9716,N_10201);
and U14080 (N_14080,N_8132,N_11725);
nor U14081 (N_14081,N_8824,N_8469);
xor U14082 (N_14082,N_11318,N_10263);
xor U14083 (N_14083,N_11710,N_11606);
nand U14084 (N_14084,N_8840,N_9951);
xnor U14085 (N_14085,N_11603,N_11719);
nand U14086 (N_14086,N_9655,N_8714);
xnor U14087 (N_14087,N_9022,N_9255);
nor U14088 (N_14088,N_11539,N_9146);
xnor U14089 (N_14089,N_11734,N_11157);
nand U14090 (N_14090,N_10861,N_8035);
nor U14091 (N_14091,N_11701,N_8025);
nor U14092 (N_14092,N_8341,N_11400);
nor U14093 (N_14093,N_11039,N_10914);
and U14094 (N_14094,N_8858,N_9126);
nand U14095 (N_14095,N_11954,N_11290);
nand U14096 (N_14096,N_9849,N_10533);
and U14097 (N_14097,N_9898,N_10336);
and U14098 (N_14098,N_8190,N_11923);
and U14099 (N_14099,N_10903,N_8099);
or U14100 (N_14100,N_8818,N_10996);
xnor U14101 (N_14101,N_8258,N_10432);
nor U14102 (N_14102,N_11067,N_9083);
or U14103 (N_14103,N_11746,N_11748);
nor U14104 (N_14104,N_10969,N_10608);
xor U14105 (N_14105,N_8845,N_9376);
and U14106 (N_14106,N_11364,N_10293);
nor U14107 (N_14107,N_10714,N_8743);
nand U14108 (N_14108,N_11368,N_8162);
nor U14109 (N_14109,N_9294,N_10324);
nand U14110 (N_14110,N_9940,N_10925);
xnor U14111 (N_14111,N_8743,N_11066);
or U14112 (N_14112,N_10482,N_11984);
or U14113 (N_14113,N_11400,N_8232);
nor U14114 (N_14114,N_9483,N_10648);
nand U14115 (N_14115,N_9542,N_11761);
or U14116 (N_14116,N_8539,N_8184);
nand U14117 (N_14117,N_11219,N_10757);
or U14118 (N_14118,N_10656,N_9557);
or U14119 (N_14119,N_10685,N_8118);
or U14120 (N_14120,N_9594,N_11476);
and U14121 (N_14121,N_10890,N_11116);
nand U14122 (N_14122,N_9007,N_11189);
xnor U14123 (N_14123,N_9107,N_10226);
or U14124 (N_14124,N_8093,N_10493);
nand U14125 (N_14125,N_9988,N_10730);
and U14126 (N_14126,N_9637,N_10329);
xnor U14127 (N_14127,N_10635,N_11597);
nor U14128 (N_14128,N_9517,N_8081);
nor U14129 (N_14129,N_9223,N_10802);
nor U14130 (N_14130,N_10871,N_8028);
xnor U14131 (N_14131,N_10116,N_9294);
or U14132 (N_14132,N_11369,N_8433);
and U14133 (N_14133,N_8738,N_10806);
xor U14134 (N_14134,N_8914,N_10174);
or U14135 (N_14135,N_8181,N_8373);
or U14136 (N_14136,N_10794,N_9619);
or U14137 (N_14137,N_10632,N_10958);
nor U14138 (N_14138,N_11769,N_8040);
nand U14139 (N_14139,N_9927,N_8853);
and U14140 (N_14140,N_10722,N_8048);
nor U14141 (N_14141,N_9261,N_10437);
nor U14142 (N_14142,N_8839,N_9158);
or U14143 (N_14143,N_10361,N_11545);
and U14144 (N_14144,N_10717,N_9629);
nand U14145 (N_14145,N_8649,N_11886);
nand U14146 (N_14146,N_9220,N_11859);
or U14147 (N_14147,N_10663,N_8703);
xor U14148 (N_14148,N_11850,N_9284);
nand U14149 (N_14149,N_8241,N_11441);
or U14150 (N_14150,N_9222,N_10819);
xnor U14151 (N_14151,N_10990,N_8030);
and U14152 (N_14152,N_11631,N_11357);
nor U14153 (N_14153,N_11925,N_9372);
nor U14154 (N_14154,N_8877,N_11866);
or U14155 (N_14155,N_9846,N_9340);
xnor U14156 (N_14156,N_11608,N_9808);
xor U14157 (N_14157,N_10786,N_11823);
xor U14158 (N_14158,N_8283,N_11059);
and U14159 (N_14159,N_8078,N_9258);
or U14160 (N_14160,N_9166,N_11996);
and U14161 (N_14161,N_9851,N_11564);
nand U14162 (N_14162,N_8511,N_10978);
nor U14163 (N_14163,N_10010,N_9160);
nand U14164 (N_14164,N_11791,N_10122);
xnor U14165 (N_14165,N_11035,N_11539);
or U14166 (N_14166,N_11933,N_11001);
xnor U14167 (N_14167,N_9976,N_10621);
nor U14168 (N_14168,N_9465,N_8588);
nand U14169 (N_14169,N_10640,N_9481);
nand U14170 (N_14170,N_10687,N_10684);
xnor U14171 (N_14171,N_10560,N_8299);
xor U14172 (N_14172,N_10867,N_10030);
xnor U14173 (N_14173,N_10064,N_10536);
nand U14174 (N_14174,N_11479,N_8333);
xor U14175 (N_14175,N_10475,N_10295);
nand U14176 (N_14176,N_10354,N_10735);
or U14177 (N_14177,N_9093,N_8225);
and U14178 (N_14178,N_10001,N_8896);
nor U14179 (N_14179,N_8055,N_11490);
or U14180 (N_14180,N_8644,N_10123);
and U14181 (N_14181,N_9962,N_11022);
xor U14182 (N_14182,N_11408,N_9028);
or U14183 (N_14183,N_10764,N_11771);
nand U14184 (N_14184,N_9688,N_11901);
or U14185 (N_14185,N_10769,N_10211);
and U14186 (N_14186,N_11931,N_8946);
nand U14187 (N_14187,N_8035,N_10249);
and U14188 (N_14188,N_11791,N_8430);
xor U14189 (N_14189,N_10290,N_11119);
nor U14190 (N_14190,N_8020,N_8094);
nor U14191 (N_14191,N_11640,N_10245);
or U14192 (N_14192,N_8622,N_11492);
and U14193 (N_14193,N_10270,N_11163);
and U14194 (N_14194,N_10233,N_11826);
or U14195 (N_14195,N_8824,N_9005);
nor U14196 (N_14196,N_9768,N_8778);
nand U14197 (N_14197,N_9766,N_9441);
or U14198 (N_14198,N_10745,N_9101);
or U14199 (N_14199,N_11864,N_8511);
or U14200 (N_14200,N_9363,N_9750);
and U14201 (N_14201,N_8389,N_10276);
or U14202 (N_14202,N_10891,N_9017);
or U14203 (N_14203,N_9024,N_8905);
nor U14204 (N_14204,N_11922,N_10749);
and U14205 (N_14205,N_9028,N_10007);
nand U14206 (N_14206,N_10032,N_11014);
nand U14207 (N_14207,N_9568,N_8892);
nand U14208 (N_14208,N_10024,N_10298);
and U14209 (N_14209,N_10901,N_8126);
xor U14210 (N_14210,N_9616,N_10503);
xnor U14211 (N_14211,N_11462,N_9755);
nor U14212 (N_14212,N_11650,N_8397);
and U14213 (N_14213,N_8350,N_9931);
and U14214 (N_14214,N_8730,N_8909);
nor U14215 (N_14215,N_8334,N_9589);
and U14216 (N_14216,N_8572,N_9640);
nor U14217 (N_14217,N_9352,N_8949);
or U14218 (N_14218,N_11335,N_10160);
or U14219 (N_14219,N_9885,N_8075);
nor U14220 (N_14220,N_10938,N_9629);
nor U14221 (N_14221,N_8884,N_11000);
nor U14222 (N_14222,N_11603,N_11332);
or U14223 (N_14223,N_11763,N_9295);
nand U14224 (N_14224,N_10916,N_11353);
nor U14225 (N_14225,N_8840,N_9018);
xor U14226 (N_14226,N_8306,N_11462);
or U14227 (N_14227,N_9918,N_10569);
nand U14228 (N_14228,N_9600,N_11325);
and U14229 (N_14229,N_9874,N_9986);
nand U14230 (N_14230,N_9037,N_9951);
xor U14231 (N_14231,N_11812,N_9400);
or U14232 (N_14232,N_10558,N_11433);
and U14233 (N_14233,N_11026,N_8515);
or U14234 (N_14234,N_9975,N_8413);
and U14235 (N_14235,N_9281,N_9524);
or U14236 (N_14236,N_10471,N_9002);
and U14237 (N_14237,N_8404,N_9035);
or U14238 (N_14238,N_8024,N_11451);
or U14239 (N_14239,N_8046,N_9631);
or U14240 (N_14240,N_9694,N_10518);
and U14241 (N_14241,N_9932,N_9402);
and U14242 (N_14242,N_10274,N_10738);
nand U14243 (N_14243,N_9212,N_9045);
and U14244 (N_14244,N_8101,N_8490);
and U14245 (N_14245,N_9419,N_10606);
and U14246 (N_14246,N_11223,N_11736);
and U14247 (N_14247,N_9525,N_9480);
nor U14248 (N_14248,N_11094,N_11230);
nand U14249 (N_14249,N_10141,N_8910);
xor U14250 (N_14250,N_9617,N_11321);
xnor U14251 (N_14251,N_8327,N_10455);
and U14252 (N_14252,N_10220,N_9402);
nand U14253 (N_14253,N_10771,N_11225);
nor U14254 (N_14254,N_10202,N_8487);
and U14255 (N_14255,N_11975,N_8591);
and U14256 (N_14256,N_11419,N_10207);
or U14257 (N_14257,N_9950,N_10826);
nor U14258 (N_14258,N_10960,N_11505);
or U14259 (N_14259,N_11829,N_8308);
nor U14260 (N_14260,N_11356,N_11193);
xnor U14261 (N_14261,N_10662,N_10766);
and U14262 (N_14262,N_11257,N_11587);
nand U14263 (N_14263,N_11426,N_9844);
or U14264 (N_14264,N_8917,N_10004);
nor U14265 (N_14265,N_9377,N_11751);
and U14266 (N_14266,N_10903,N_11011);
or U14267 (N_14267,N_10407,N_10606);
nor U14268 (N_14268,N_11975,N_8541);
and U14269 (N_14269,N_11927,N_10730);
nor U14270 (N_14270,N_9368,N_11850);
nor U14271 (N_14271,N_8277,N_8081);
and U14272 (N_14272,N_11323,N_11980);
nand U14273 (N_14273,N_10996,N_10214);
nand U14274 (N_14274,N_10091,N_11558);
or U14275 (N_14275,N_10296,N_9554);
xnor U14276 (N_14276,N_10736,N_9040);
nor U14277 (N_14277,N_9367,N_8181);
nand U14278 (N_14278,N_8325,N_10928);
nor U14279 (N_14279,N_9843,N_10831);
nand U14280 (N_14280,N_11186,N_9954);
and U14281 (N_14281,N_10321,N_8567);
or U14282 (N_14282,N_11929,N_9113);
nor U14283 (N_14283,N_9971,N_9732);
and U14284 (N_14284,N_9059,N_10337);
and U14285 (N_14285,N_8221,N_11716);
xor U14286 (N_14286,N_10199,N_11060);
or U14287 (N_14287,N_9689,N_11174);
nand U14288 (N_14288,N_10286,N_8279);
and U14289 (N_14289,N_10475,N_8347);
nand U14290 (N_14290,N_11459,N_10715);
xnor U14291 (N_14291,N_9935,N_11314);
and U14292 (N_14292,N_11873,N_11569);
and U14293 (N_14293,N_8532,N_11140);
xnor U14294 (N_14294,N_8608,N_10216);
nand U14295 (N_14295,N_11387,N_9409);
xnor U14296 (N_14296,N_10379,N_10958);
nor U14297 (N_14297,N_10834,N_8388);
nor U14298 (N_14298,N_11865,N_11391);
nor U14299 (N_14299,N_11948,N_8545);
and U14300 (N_14300,N_11325,N_9114);
nor U14301 (N_14301,N_11313,N_8076);
xnor U14302 (N_14302,N_8069,N_10109);
nand U14303 (N_14303,N_8351,N_9929);
nand U14304 (N_14304,N_8040,N_9445);
nand U14305 (N_14305,N_8556,N_8262);
or U14306 (N_14306,N_8719,N_8656);
and U14307 (N_14307,N_9909,N_8850);
and U14308 (N_14308,N_10231,N_11811);
nor U14309 (N_14309,N_9472,N_10931);
or U14310 (N_14310,N_10966,N_10011);
xnor U14311 (N_14311,N_10355,N_8869);
nor U14312 (N_14312,N_10275,N_10099);
and U14313 (N_14313,N_9687,N_8883);
nand U14314 (N_14314,N_9924,N_8298);
nor U14315 (N_14315,N_9689,N_11056);
or U14316 (N_14316,N_8867,N_9427);
xnor U14317 (N_14317,N_8189,N_11067);
nand U14318 (N_14318,N_8059,N_11948);
xnor U14319 (N_14319,N_8104,N_10795);
and U14320 (N_14320,N_9272,N_9792);
and U14321 (N_14321,N_8952,N_11069);
or U14322 (N_14322,N_8164,N_8664);
and U14323 (N_14323,N_11541,N_9241);
xnor U14324 (N_14324,N_8929,N_9425);
and U14325 (N_14325,N_9565,N_10156);
nor U14326 (N_14326,N_10171,N_11816);
nor U14327 (N_14327,N_11928,N_11239);
or U14328 (N_14328,N_9928,N_11666);
and U14329 (N_14329,N_8122,N_11135);
or U14330 (N_14330,N_8890,N_11911);
nor U14331 (N_14331,N_9849,N_10716);
nand U14332 (N_14332,N_9817,N_9024);
xor U14333 (N_14333,N_9503,N_11045);
and U14334 (N_14334,N_10081,N_8925);
and U14335 (N_14335,N_9555,N_9761);
nor U14336 (N_14336,N_9966,N_11727);
nor U14337 (N_14337,N_9372,N_8193);
or U14338 (N_14338,N_11941,N_8068);
nand U14339 (N_14339,N_10363,N_10035);
nand U14340 (N_14340,N_8541,N_9861);
and U14341 (N_14341,N_10957,N_9962);
and U14342 (N_14342,N_8174,N_9858);
or U14343 (N_14343,N_9985,N_10906);
nor U14344 (N_14344,N_9607,N_9847);
nand U14345 (N_14345,N_10380,N_11356);
or U14346 (N_14346,N_8908,N_10923);
nand U14347 (N_14347,N_9390,N_10523);
xnor U14348 (N_14348,N_9893,N_8967);
xor U14349 (N_14349,N_11908,N_9082);
nor U14350 (N_14350,N_9416,N_10174);
xnor U14351 (N_14351,N_8297,N_10798);
nand U14352 (N_14352,N_8968,N_8988);
and U14353 (N_14353,N_10617,N_10256);
or U14354 (N_14354,N_10842,N_8379);
nand U14355 (N_14355,N_10524,N_10098);
nand U14356 (N_14356,N_9997,N_9097);
nor U14357 (N_14357,N_10194,N_9808);
xor U14358 (N_14358,N_9848,N_9019);
nor U14359 (N_14359,N_9156,N_10782);
nor U14360 (N_14360,N_11584,N_11023);
nor U14361 (N_14361,N_11651,N_11626);
and U14362 (N_14362,N_8462,N_10491);
nor U14363 (N_14363,N_8187,N_9431);
and U14364 (N_14364,N_11575,N_10314);
nand U14365 (N_14365,N_11330,N_10207);
nor U14366 (N_14366,N_11692,N_8753);
or U14367 (N_14367,N_11413,N_11591);
xor U14368 (N_14368,N_8345,N_11902);
or U14369 (N_14369,N_9319,N_9067);
or U14370 (N_14370,N_9202,N_9142);
nor U14371 (N_14371,N_10085,N_8870);
or U14372 (N_14372,N_11383,N_10451);
nand U14373 (N_14373,N_10418,N_9259);
or U14374 (N_14374,N_9331,N_10052);
nor U14375 (N_14375,N_8574,N_9865);
xor U14376 (N_14376,N_8564,N_8298);
xor U14377 (N_14377,N_9527,N_9291);
nand U14378 (N_14378,N_11916,N_10352);
or U14379 (N_14379,N_8338,N_11165);
and U14380 (N_14380,N_8294,N_9558);
xor U14381 (N_14381,N_8799,N_9727);
nand U14382 (N_14382,N_9216,N_11431);
or U14383 (N_14383,N_10436,N_10229);
nand U14384 (N_14384,N_10191,N_11189);
nand U14385 (N_14385,N_8322,N_9920);
nand U14386 (N_14386,N_9187,N_8184);
nand U14387 (N_14387,N_9340,N_11800);
or U14388 (N_14388,N_8600,N_8803);
or U14389 (N_14389,N_11731,N_11059);
and U14390 (N_14390,N_10059,N_11824);
xor U14391 (N_14391,N_8478,N_10268);
or U14392 (N_14392,N_10099,N_11130);
nand U14393 (N_14393,N_10093,N_11855);
nor U14394 (N_14394,N_11281,N_10116);
nand U14395 (N_14395,N_8661,N_10729);
xor U14396 (N_14396,N_10612,N_10663);
nor U14397 (N_14397,N_8912,N_8011);
nor U14398 (N_14398,N_9019,N_10356);
nand U14399 (N_14399,N_9791,N_9143);
or U14400 (N_14400,N_10388,N_8821);
nor U14401 (N_14401,N_11812,N_11816);
nand U14402 (N_14402,N_9788,N_11913);
or U14403 (N_14403,N_10337,N_11280);
nand U14404 (N_14404,N_11592,N_11999);
nand U14405 (N_14405,N_10114,N_10693);
nor U14406 (N_14406,N_11874,N_9332);
nand U14407 (N_14407,N_9727,N_8324);
nand U14408 (N_14408,N_9847,N_9017);
nor U14409 (N_14409,N_9611,N_11290);
nor U14410 (N_14410,N_10257,N_10652);
or U14411 (N_14411,N_9162,N_9644);
xnor U14412 (N_14412,N_11885,N_9013);
nand U14413 (N_14413,N_8675,N_10902);
or U14414 (N_14414,N_8060,N_10073);
nand U14415 (N_14415,N_10790,N_11671);
or U14416 (N_14416,N_11857,N_9638);
and U14417 (N_14417,N_10277,N_9248);
xor U14418 (N_14418,N_9664,N_11825);
nor U14419 (N_14419,N_9845,N_8703);
and U14420 (N_14420,N_8385,N_9897);
or U14421 (N_14421,N_10521,N_9037);
nand U14422 (N_14422,N_9837,N_9815);
nand U14423 (N_14423,N_10318,N_10361);
and U14424 (N_14424,N_9191,N_8475);
nor U14425 (N_14425,N_9684,N_10791);
nor U14426 (N_14426,N_11297,N_8948);
or U14427 (N_14427,N_8578,N_11014);
nand U14428 (N_14428,N_11061,N_11532);
or U14429 (N_14429,N_11317,N_8567);
xor U14430 (N_14430,N_9184,N_9716);
and U14431 (N_14431,N_8515,N_8133);
xor U14432 (N_14432,N_8642,N_11230);
or U14433 (N_14433,N_10864,N_11926);
and U14434 (N_14434,N_8579,N_8108);
nand U14435 (N_14435,N_11503,N_11814);
and U14436 (N_14436,N_11483,N_11050);
or U14437 (N_14437,N_8240,N_8079);
xnor U14438 (N_14438,N_8804,N_8755);
and U14439 (N_14439,N_9126,N_11377);
or U14440 (N_14440,N_8134,N_10791);
xor U14441 (N_14441,N_8032,N_9314);
nor U14442 (N_14442,N_10742,N_9815);
nand U14443 (N_14443,N_9013,N_8855);
and U14444 (N_14444,N_11820,N_8202);
nor U14445 (N_14445,N_8741,N_9489);
nor U14446 (N_14446,N_10157,N_8309);
and U14447 (N_14447,N_10611,N_9958);
nor U14448 (N_14448,N_9914,N_11060);
nand U14449 (N_14449,N_9536,N_9695);
nor U14450 (N_14450,N_8235,N_11690);
nor U14451 (N_14451,N_11565,N_10931);
nand U14452 (N_14452,N_8689,N_9860);
xnor U14453 (N_14453,N_8745,N_9337);
and U14454 (N_14454,N_11252,N_10120);
and U14455 (N_14455,N_9703,N_8903);
and U14456 (N_14456,N_10921,N_9595);
or U14457 (N_14457,N_10256,N_8358);
xnor U14458 (N_14458,N_8431,N_11760);
and U14459 (N_14459,N_8933,N_10302);
and U14460 (N_14460,N_11149,N_11558);
nor U14461 (N_14461,N_8594,N_8772);
nor U14462 (N_14462,N_8948,N_10967);
xnor U14463 (N_14463,N_10446,N_10609);
xor U14464 (N_14464,N_10337,N_9453);
nand U14465 (N_14465,N_9095,N_10390);
or U14466 (N_14466,N_9895,N_9682);
nand U14467 (N_14467,N_10706,N_8812);
xnor U14468 (N_14468,N_9035,N_10618);
nand U14469 (N_14469,N_9582,N_8103);
xor U14470 (N_14470,N_9795,N_8080);
nand U14471 (N_14471,N_10853,N_8322);
and U14472 (N_14472,N_9375,N_9905);
and U14473 (N_14473,N_10401,N_10604);
nand U14474 (N_14474,N_10388,N_9919);
and U14475 (N_14475,N_9550,N_10263);
nand U14476 (N_14476,N_10605,N_9549);
or U14477 (N_14477,N_8475,N_8944);
and U14478 (N_14478,N_8250,N_9649);
nor U14479 (N_14479,N_11382,N_9607);
or U14480 (N_14480,N_10045,N_8391);
or U14481 (N_14481,N_9030,N_9987);
or U14482 (N_14482,N_10328,N_9999);
and U14483 (N_14483,N_8883,N_11199);
nand U14484 (N_14484,N_8540,N_11967);
xor U14485 (N_14485,N_10314,N_9499);
nor U14486 (N_14486,N_9427,N_8821);
or U14487 (N_14487,N_9393,N_9815);
nor U14488 (N_14488,N_9779,N_10581);
nor U14489 (N_14489,N_11068,N_8631);
and U14490 (N_14490,N_11183,N_9470);
nor U14491 (N_14491,N_9582,N_9762);
nor U14492 (N_14492,N_8497,N_11046);
and U14493 (N_14493,N_8933,N_11554);
or U14494 (N_14494,N_9744,N_8971);
or U14495 (N_14495,N_10756,N_10641);
xnor U14496 (N_14496,N_8320,N_9962);
nand U14497 (N_14497,N_10662,N_8932);
or U14498 (N_14498,N_8896,N_11947);
and U14499 (N_14499,N_10874,N_10740);
and U14500 (N_14500,N_9847,N_9318);
nor U14501 (N_14501,N_9466,N_9720);
xnor U14502 (N_14502,N_11379,N_10235);
nor U14503 (N_14503,N_11944,N_9651);
or U14504 (N_14504,N_8423,N_9034);
nand U14505 (N_14505,N_10370,N_8689);
nor U14506 (N_14506,N_9214,N_9987);
nand U14507 (N_14507,N_9360,N_8593);
xor U14508 (N_14508,N_10591,N_11715);
nand U14509 (N_14509,N_8248,N_11599);
or U14510 (N_14510,N_10647,N_9950);
xnor U14511 (N_14511,N_9277,N_10977);
and U14512 (N_14512,N_11056,N_8810);
nor U14513 (N_14513,N_9890,N_8379);
and U14514 (N_14514,N_8922,N_11767);
xor U14515 (N_14515,N_9713,N_9726);
or U14516 (N_14516,N_10188,N_10934);
xor U14517 (N_14517,N_9877,N_11536);
xnor U14518 (N_14518,N_10458,N_9896);
and U14519 (N_14519,N_11991,N_10963);
or U14520 (N_14520,N_8167,N_10884);
and U14521 (N_14521,N_9514,N_9815);
nor U14522 (N_14522,N_8765,N_9585);
xnor U14523 (N_14523,N_9293,N_11926);
xor U14524 (N_14524,N_11185,N_8326);
and U14525 (N_14525,N_9507,N_8273);
xor U14526 (N_14526,N_11909,N_11112);
or U14527 (N_14527,N_11974,N_9427);
and U14528 (N_14528,N_9503,N_9994);
nor U14529 (N_14529,N_11645,N_11191);
nand U14530 (N_14530,N_11433,N_10788);
nor U14531 (N_14531,N_11641,N_10594);
and U14532 (N_14532,N_8230,N_8171);
nand U14533 (N_14533,N_11526,N_11116);
nand U14534 (N_14534,N_11456,N_8910);
or U14535 (N_14535,N_8062,N_9897);
xnor U14536 (N_14536,N_8824,N_9322);
or U14537 (N_14537,N_9602,N_10465);
and U14538 (N_14538,N_11333,N_9550);
xnor U14539 (N_14539,N_8933,N_9309);
or U14540 (N_14540,N_11747,N_9835);
or U14541 (N_14541,N_8858,N_9414);
or U14542 (N_14542,N_9227,N_8243);
xor U14543 (N_14543,N_9510,N_11686);
nor U14544 (N_14544,N_11173,N_10746);
xor U14545 (N_14545,N_9598,N_9918);
xnor U14546 (N_14546,N_10485,N_8026);
nand U14547 (N_14547,N_10109,N_8972);
xor U14548 (N_14548,N_10736,N_9195);
xor U14549 (N_14549,N_11431,N_11198);
nor U14550 (N_14550,N_10496,N_8957);
nand U14551 (N_14551,N_11551,N_10389);
xnor U14552 (N_14552,N_9984,N_8523);
nor U14553 (N_14553,N_10196,N_10706);
xor U14554 (N_14554,N_10040,N_8033);
or U14555 (N_14555,N_11162,N_10951);
xor U14556 (N_14556,N_11434,N_8282);
and U14557 (N_14557,N_8142,N_9109);
nand U14558 (N_14558,N_11105,N_11205);
or U14559 (N_14559,N_11255,N_10976);
or U14560 (N_14560,N_8851,N_9289);
nor U14561 (N_14561,N_9833,N_8584);
nor U14562 (N_14562,N_9721,N_10135);
nor U14563 (N_14563,N_10120,N_11399);
or U14564 (N_14564,N_11708,N_9032);
xor U14565 (N_14565,N_9066,N_10809);
nor U14566 (N_14566,N_10256,N_10172);
or U14567 (N_14567,N_11683,N_10649);
or U14568 (N_14568,N_11050,N_8452);
nand U14569 (N_14569,N_11013,N_10292);
xor U14570 (N_14570,N_11539,N_8774);
or U14571 (N_14571,N_10523,N_10391);
xor U14572 (N_14572,N_8814,N_10202);
nand U14573 (N_14573,N_8795,N_9152);
nand U14574 (N_14574,N_11518,N_11808);
nor U14575 (N_14575,N_11706,N_8831);
xnor U14576 (N_14576,N_8565,N_10508);
nand U14577 (N_14577,N_10387,N_8806);
xnor U14578 (N_14578,N_9272,N_8215);
xor U14579 (N_14579,N_8657,N_11373);
nand U14580 (N_14580,N_8902,N_8453);
nand U14581 (N_14581,N_11626,N_9594);
or U14582 (N_14582,N_10198,N_10756);
xor U14583 (N_14583,N_10303,N_9364);
nor U14584 (N_14584,N_11498,N_11058);
nand U14585 (N_14585,N_9729,N_10586);
and U14586 (N_14586,N_9922,N_8226);
nand U14587 (N_14587,N_10231,N_11774);
nor U14588 (N_14588,N_11728,N_8584);
and U14589 (N_14589,N_8864,N_9167);
nand U14590 (N_14590,N_8277,N_11947);
nor U14591 (N_14591,N_9090,N_8319);
and U14592 (N_14592,N_11669,N_10852);
nor U14593 (N_14593,N_9480,N_11056);
nor U14594 (N_14594,N_10246,N_8579);
nor U14595 (N_14595,N_8481,N_10561);
or U14596 (N_14596,N_8092,N_9251);
nand U14597 (N_14597,N_9879,N_9113);
nand U14598 (N_14598,N_11027,N_10098);
and U14599 (N_14599,N_9323,N_9497);
or U14600 (N_14600,N_11312,N_8922);
or U14601 (N_14601,N_9687,N_10939);
nor U14602 (N_14602,N_9431,N_8656);
xnor U14603 (N_14603,N_8678,N_10025);
and U14604 (N_14604,N_9727,N_10211);
nor U14605 (N_14605,N_8773,N_10255);
and U14606 (N_14606,N_10887,N_9376);
nand U14607 (N_14607,N_9637,N_8034);
nor U14608 (N_14608,N_11634,N_8217);
xor U14609 (N_14609,N_11263,N_11746);
xnor U14610 (N_14610,N_8008,N_9262);
and U14611 (N_14611,N_11355,N_9539);
and U14612 (N_14612,N_10144,N_11166);
nor U14613 (N_14613,N_8831,N_10325);
and U14614 (N_14614,N_8936,N_8766);
nand U14615 (N_14615,N_8481,N_9044);
and U14616 (N_14616,N_8330,N_8808);
or U14617 (N_14617,N_10809,N_11782);
or U14618 (N_14618,N_10221,N_10326);
nor U14619 (N_14619,N_10588,N_9509);
nor U14620 (N_14620,N_8222,N_8416);
nor U14621 (N_14621,N_10161,N_10163);
nand U14622 (N_14622,N_10048,N_8701);
or U14623 (N_14623,N_8087,N_9244);
nor U14624 (N_14624,N_11047,N_8967);
nand U14625 (N_14625,N_8552,N_10245);
nor U14626 (N_14626,N_8393,N_8345);
xnor U14627 (N_14627,N_9097,N_9480);
or U14628 (N_14628,N_11310,N_9381);
or U14629 (N_14629,N_8698,N_11782);
or U14630 (N_14630,N_8277,N_11519);
xnor U14631 (N_14631,N_9873,N_8057);
nor U14632 (N_14632,N_8120,N_8066);
or U14633 (N_14633,N_10146,N_11437);
xor U14634 (N_14634,N_10427,N_8309);
xor U14635 (N_14635,N_9617,N_11530);
and U14636 (N_14636,N_10799,N_8376);
nand U14637 (N_14637,N_9818,N_11003);
or U14638 (N_14638,N_9065,N_9002);
nand U14639 (N_14639,N_8764,N_11233);
nor U14640 (N_14640,N_8814,N_8319);
or U14641 (N_14641,N_10090,N_10073);
nor U14642 (N_14642,N_10326,N_10344);
nor U14643 (N_14643,N_11819,N_9871);
xnor U14644 (N_14644,N_10393,N_10310);
xor U14645 (N_14645,N_8337,N_11713);
or U14646 (N_14646,N_9885,N_10066);
nand U14647 (N_14647,N_11158,N_9678);
nor U14648 (N_14648,N_10626,N_11615);
and U14649 (N_14649,N_11897,N_11052);
nand U14650 (N_14650,N_11642,N_10744);
nand U14651 (N_14651,N_10077,N_9522);
nand U14652 (N_14652,N_11776,N_10605);
and U14653 (N_14653,N_10894,N_9878);
xor U14654 (N_14654,N_11115,N_8559);
nand U14655 (N_14655,N_11590,N_8060);
or U14656 (N_14656,N_11235,N_10766);
nor U14657 (N_14657,N_9126,N_9744);
nand U14658 (N_14658,N_10783,N_8525);
or U14659 (N_14659,N_11380,N_11473);
nand U14660 (N_14660,N_9012,N_9266);
xor U14661 (N_14661,N_9453,N_8390);
nor U14662 (N_14662,N_8953,N_8522);
nor U14663 (N_14663,N_10896,N_9626);
xor U14664 (N_14664,N_11417,N_11507);
xor U14665 (N_14665,N_10753,N_10073);
and U14666 (N_14666,N_11889,N_9237);
or U14667 (N_14667,N_8997,N_9201);
xor U14668 (N_14668,N_8326,N_11049);
xor U14669 (N_14669,N_11539,N_9411);
nand U14670 (N_14670,N_10430,N_9861);
and U14671 (N_14671,N_9046,N_8013);
nand U14672 (N_14672,N_11755,N_10467);
and U14673 (N_14673,N_10725,N_10282);
and U14674 (N_14674,N_9739,N_10099);
and U14675 (N_14675,N_8558,N_9982);
xnor U14676 (N_14676,N_9064,N_8835);
and U14677 (N_14677,N_11705,N_10259);
nand U14678 (N_14678,N_10638,N_10038);
nor U14679 (N_14679,N_9739,N_10921);
or U14680 (N_14680,N_9208,N_9891);
nand U14681 (N_14681,N_11534,N_8498);
nor U14682 (N_14682,N_11904,N_10090);
and U14683 (N_14683,N_9406,N_10502);
xnor U14684 (N_14684,N_8085,N_11512);
xor U14685 (N_14685,N_11082,N_9261);
nand U14686 (N_14686,N_8023,N_9941);
nand U14687 (N_14687,N_8872,N_10968);
nand U14688 (N_14688,N_10760,N_11268);
nor U14689 (N_14689,N_8125,N_8481);
and U14690 (N_14690,N_10177,N_11102);
xnor U14691 (N_14691,N_10297,N_8206);
or U14692 (N_14692,N_9934,N_8362);
xor U14693 (N_14693,N_10771,N_8148);
and U14694 (N_14694,N_9370,N_9264);
xor U14695 (N_14695,N_11973,N_10504);
nand U14696 (N_14696,N_10167,N_8196);
nand U14697 (N_14697,N_10614,N_10813);
and U14698 (N_14698,N_8020,N_9564);
nor U14699 (N_14699,N_9368,N_9815);
nand U14700 (N_14700,N_10098,N_10011);
nand U14701 (N_14701,N_9752,N_8189);
or U14702 (N_14702,N_8274,N_8910);
nand U14703 (N_14703,N_8830,N_10611);
or U14704 (N_14704,N_9311,N_8859);
and U14705 (N_14705,N_10676,N_8145);
or U14706 (N_14706,N_8316,N_11913);
or U14707 (N_14707,N_8582,N_8628);
nand U14708 (N_14708,N_9383,N_10277);
or U14709 (N_14709,N_8735,N_8531);
and U14710 (N_14710,N_8307,N_10828);
nand U14711 (N_14711,N_10668,N_10889);
nor U14712 (N_14712,N_11264,N_9085);
and U14713 (N_14713,N_10434,N_10030);
and U14714 (N_14714,N_8394,N_11370);
nor U14715 (N_14715,N_11760,N_8393);
nand U14716 (N_14716,N_9344,N_9474);
or U14717 (N_14717,N_8576,N_9223);
or U14718 (N_14718,N_8504,N_10529);
xnor U14719 (N_14719,N_9721,N_9944);
nand U14720 (N_14720,N_8795,N_9544);
nor U14721 (N_14721,N_11176,N_11183);
and U14722 (N_14722,N_8545,N_10418);
xor U14723 (N_14723,N_8039,N_10468);
xnor U14724 (N_14724,N_10403,N_11147);
or U14725 (N_14725,N_8891,N_9745);
or U14726 (N_14726,N_11955,N_10576);
or U14727 (N_14727,N_8493,N_11798);
and U14728 (N_14728,N_9796,N_9888);
or U14729 (N_14729,N_9398,N_11683);
nand U14730 (N_14730,N_9873,N_11955);
or U14731 (N_14731,N_10004,N_9240);
nand U14732 (N_14732,N_11589,N_9853);
nor U14733 (N_14733,N_10232,N_9850);
nor U14734 (N_14734,N_9074,N_10571);
nor U14735 (N_14735,N_8476,N_10443);
and U14736 (N_14736,N_8819,N_10506);
nor U14737 (N_14737,N_9509,N_9182);
or U14738 (N_14738,N_10619,N_9273);
and U14739 (N_14739,N_11653,N_11193);
nand U14740 (N_14740,N_8459,N_11829);
nand U14741 (N_14741,N_10652,N_11901);
nor U14742 (N_14742,N_9213,N_11112);
nand U14743 (N_14743,N_8241,N_8331);
xor U14744 (N_14744,N_9618,N_9955);
and U14745 (N_14745,N_11436,N_10623);
and U14746 (N_14746,N_10729,N_10766);
and U14747 (N_14747,N_11410,N_8027);
and U14748 (N_14748,N_8346,N_10068);
nand U14749 (N_14749,N_9547,N_11064);
or U14750 (N_14750,N_9572,N_8070);
nand U14751 (N_14751,N_8914,N_8284);
and U14752 (N_14752,N_9309,N_11747);
and U14753 (N_14753,N_10231,N_8876);
or U14754 (N_14754,N_11668,N_8769);
xor U14755 (N_14755,N_9129,N_10864);
or U14756 (N_14756,N_11270,N_8724);
xnor U14757 (N_14757,N_11034,N_8408);
and U14758 (N_14758,N_10678,N_11264);
nor U14759 (N_14759,N_10647,N_10775);
or U14760 (N_14760,N_11312,N_8043);
or U14761 (N_14761,N_10913,N_11495);
or U14762 (N_14762,N_11990,N_10314);
and U14763 (N_14763,N_9828,N_11557);
nand U14764 (N_14764,N_9612,N_10291);
xor U14765 (N_14765,N_9008,N_9328);
or U14766 (N_14766,N_8471,N_10687);
xor U14767 (N_14767,N_8557,N_11780);
or U14768 (N_14768,N_10958,N_8834);
and U14769 (N_14769,N_11330,N_9849);
or U14770 (N_14770,N_10109,N_10526);
or U14771 (N_14771,N_11038,N_10427);
nor U14772 (N_14772,N_11510,N_9075);
and U14773 (N_14773,N_10531,N_9102);
and U14774 (N_14774,N_10834,N_8319);
nand U14775 (N_14775,N_11350,N_9093);
or U14776 (N_14776,N_11744,N_8283);
and U14777 (N_14777,N_9018,N_10479);
and U14778 (N_14778,N_10609,N_9620);
xnor U14779 (N_14779,N_9868,N_9054);
or U14780 (N_14780,N_9668,N_8681);
or U14781 (N_14781,N_11795,N_9339);
xor U14782 (N_14782,N_11666,N_9044);
xor U14783 (N_14783,N_8803,N_11647);
xnor U14784 (N_14784,N_11777,N_10034);
nand U14785 (N_14785,N_8589,N_10024);
or U14786 (N_14786,N_9987,N_9192);
nand U14787 (N_14787,N_10573,N_11091);
xnor U14788 (N_14788,N_11966,N_8812);
nand U14789 (N_14789,N_10519,N_8715);
nor U14790 (N_14790,N_9198,N_11240);
nor U14791 (N_14791,N_10334,N_8076);
or U14792 (N_14792,N_9712,N_10107);
nor U14793 (N_14793,N_9092,N_10913);
nand U14794 (N_14794,N_9445,N_8695);
or U14795 (N_14795,N_9982,N_11503);
xor U14796 (N_14796,N_9603,N_8299);
and U14797 (N_14797,N_8582,N_10701);
xor U14798 (N_14798,N_8916,N_10473);
or U14799 (N_14799,N_8309,N_9400);
nand U14800 (N_14800,N_10570,N_9327);
and U14801 (N_14801,N_10424,N_10242);
nand U14802 (N_14802,N_9273,N_10582);
xnor U14803 (N_14803,N_11246,N_10188);
and U14804 (N_14804,N_10164,N_8463);
nand U14805 (N_14805,N_10078,N_9540);
xnor U14806 (N_14806,N_9643,N_8696);
nand U14807 (N_14807,N_11399,N_8678);
xnor U14808 (N_14808,N_8154,N_10112);
nand U14809 (N_14809,N_11329,N_11717);
nor U14810 (N_14810,N_10321,N_10993);
nor U14811 (N_14811,N_9195,N_9349);
xor U14812 (N_14812,N_8231,N_11989);
nand U14813 (N_14813,N_9135,N_9095);
nor U14814 (N_14814,N_11137,N_9083);
nor U14815 (N_14815,N_8725,N_9666);
xor U14816 (N_14816,N_8601,N_10301);
or U14817 (N_14817,N_9568,N_8257);
and U14818 (N_14818,N_9873,N_8653);
or U14819 (N_14819,N_9447,N_9643);
nor U14820 (N_14820,N_11509,N_10030);
or U14821 (N_14821,N_9048,N_10099);
nand U14822 (N_14822,N_11634,N_8716);
nand U14823 (N_14823,N_10304,N_11403);
or U14824 (N_14824,N_8746,N_8713);
nor U14825 (N_14825,N_10695,N_9129);
nand U14826 (N_14826,N_8417,N_9884);
or U14827 (N_14827,N_9073,N_10178);
and U14828 (N_14828,N_10134,N_11445);
xnor U14829 (N_14829,N_8299,N_10200);
nor U14830 (N_14830,N_9358,N_10190);
or U14831 (N_14831,N_11836,N_11401);
xor U14832 (N_14832,N_10730,N_10468);
nor U14833 (N_14833,N_8957,N_11629);
or U14834 (N_14834,N_10469,N_8835);
xnor U14835 (N_14835,N_11398,N_9518);
nand U14836 (N_14836,N_8751,N_8396);
xor U14837 (N_14837,N_9517,N_11625);
and U14838 (N_14838,N_9036,N_10224);
nand U14839 (N_14839,N_8680,N_10638);
nand U14840 (N_14840,N_10331,N_11877);
and U14841 (N_14841,N_11583,N_11363);
nand U14842 (N_14842,N_10921,N_11929);
or U14843 (N_14843,N_9090,N_10275);
xnor U14844 (N_14844,N_10771,N_11040);
nor U14845 (N_14845,N_11527,N_9223);
nor U14846 (N_14846,N_11651,N_8455);
nor U14847 (N_14847,N_8843,N_9914);
and U14848 (N_14848,N_8867,N_10581);
nor U14849 (N_14849,N_9680,N_11577);
nor U14850 (N_14850,N_11815,N_10140);
xor U14851 (N_14851,N_8295,N_11354);
xor U14852 (N_14852,N_10856,N_8021);
and U14853 (N_14853,N_10425,N_8505);
or U14854 (N_14854,N_10951,N_10104);
or U14855 (N_14855,N_11063,N_9573);
xor U14856 (N_14856,N_9600,N_10318);
and U14857 (N_14857,N_11419,N_9683);
nand U14858 (N_14858,N_11730,N_11666);
or U14859 (N_14859,N_10835,N_9417);
or U14860 (N_14860,N_10249,N_9924);
nand U14861 (N_14861,N_9368,N_10990);
and U14862 (N_14862,N_10930,N_11484);
nor U14863 (N_14863,N_10678,N_11505);
nand U14864 (N_14864,N_11581,N_10486);
and U14865 (N_14865,N_11452,N_11728);
xor U14866 (N_14866,N_9945,N_8233);
nor U14867 (N_14867,N_10906,N_8224);
xor U14868 (N_14868,N_11563,N_9433);
and U14869 (N_14869,N_9253,N_9994);
nand U14870 (N_14870,N_9913,N_10096);
nand U14871 (N_14871,N_8520,N_8475);
nand U14872 (N_14872,N_11396,N_10576);
xor U14873 (N_14873,N_10300,N_9803);
and U14874 (N_14874,N_8281,N_9407);
nand U14875 (N_14875,N_9325,N_8128);
or U14876 (N_14876,N_11102,N_9342);
or U14877 (N_14877,N_10928,N_8903);
nand U14878 (N_14878,N_10173,N_9315);
or U14879 (N_14879,N_11388,N_10396);
xor U14880 (N_14880,N_8583,N_10924);
nor U14881 (N_14881,N_10709,N_11831);
xor U14882 (N_14882,N_11968,N_8867);
nor U14883 (N_14883,N_9900,N_11941);
nor U14884 (N_14884,N_10587,N_8037);
nor U14885 (N_14885,N_11456,N_8088);
or U14886 (N_14886,N_9318,N_8007);
xor U14887 (N_14887,N_10937,N_8086);
xnor U14888 (N_14888,N_10119,N_10286);
nand U14889 (N_14889,N_11277,N_9079);
xor U14890 (N_14890,N_10006,N_9860);
nand U14891 (N_14891,N_8759,N_10794);
nor U14892 (N_14892,N_10859,N_8764);
nor U14893 (N_14893,N_8180,N_9785);
or U14894 (N_14894,N_9638,N_8233);
xor U14895 (N_14895,N_10713,N_10067);
nor U14896 (N_14896,N_8451,N_10861);
and U14897 (N_14897,N_11352,N_10423);
or U14898 (N_14898,N_8519,N_8651);
nor U14899 (N_14899,N_9218,N_10666);
xnor U14900 (N_14900,N_11963,N_10268);
xor U14901 (N_14901,N_10308,N_11004);
nor U14902 (N_14902,N_8404,N_10375);
nor U14903 (N_14903,N_10753,N_11453);
nor U14904 (N_14904,N_10342,N_8059);
xnor U14905 (N_14905,N_11128,N_8031);
nor U14906 (N_14906,N_11708,N_10819);
xnor U14907 (N_14907,N_9496,N_9587);
and U14908 (N_14908,N_10868,N_11274);
nor U14909 (N_14909,N_11434,N_8674);
nor U14910 (N_14910,N_9067,N_9504);
nand U14911 (N_14911,N_11077,N_10786);
nor U14912 (N_14912,N_9156,N_10896);
or U14913 (N_14913,N_11736,N_11415);
nor U14914 (N_14914,N_11754,N_9086);
nor U14915 (N_14915,N_11757,N_9828);
nor U14916 (N_14916,N_11663,N_8330);
nor U14917 (N_14917,N_11643,N_8341);
and U14918 (N_14918,N_8835,N_8143);
nor U14919 (N_14919,N_10116,N_9790);
and U14920 (N_14920,N_9444,N_9547);
nor U14921 (N_14921,N_8929,N_8095);
or U14922 (N_14922,N_9926,N_11451);
and U14923 (N_14923,N_9169,N_9375);
xnor U14924 (N_14924,N_11169,N_11616);
nor U14925 (N_14925,N_11803,N_9936);
nand U14926 (N_14926,N_8144,N_8740);
and U14927 (N_14927,N_11027,N_11231);
and U14928 (N_14928,N_10677,N_8365);
and U14929 (N_14929,N_11266,N_8416);
and U14930 (N_14930,N_9189,N_10932);
and U14931 (N_14931,N_9366,N_8022);
nor U14932 (N_14932,N_10900,N_10485);
nand U14933 (N_14933,N_10399,N_10945);
and U14934 (N_14934,N_8048,N_9073);
and U14935 (N_14935,N_9094,N_9115);
and U14936 (N_14936,N_10362,N_11649);
xor U14937 (N_14937,N_10723,N_10350);
nand U14938 (N_14938,N_10275,N_8304);
or U14939 (N_14939,N_8044,N_9117);
xor U14940 (N_14940,N_10863,N_8443);
nor U14941 (N_14941,N_11441,N_11037);
nand U14942 (N_14942,N_10888,N_11364);
nor U14943 (N_14943,N_11308,N_9925);
nor U14944 (N_14944,N_10970,N_9549);
or U14945 (N_14945,N_9671,N_10071);
and U14946 (N_14946,N_10268,N_11316);
nor U14947 (N_14947,N_10491,N_9092);
xor U14948 (N_14948,N_8885,N_11520);
and U14949 (N_14949,N_9865,N_10666);
nand U14950 (N_14950,N_8990,N_8692);
xnor U14951 (N_14951,N_8193,N_10906);
or U14952 (N_14952,N_10446,N_10862);
or U14953 (N_14953,N_8811,N_11987);
and U14954 (N_14954,N_10684,N_10570);
xor U14955 (N_14955,N_8745,N_9833);
nand U14956 (N_14956,N_8363,N_8423);
and U14957 (N_14957,N_11481,N_8780);
nor U14958 (N_14958,N_10193,N_9284);
or U14959 (N_14959,N_11128,N_10561);
nor U14960 (N_14960,N_11212,N_11962);
xor U14961 (N_14961,N_11267,N_8267);
or U14962 (N_14962,N_10504,N_10698);
nand U14963 (N_14963,N_9522,N_8750);
or U14964 (N_14964,N_10358,N_8240);
xor U14965 (N_14965,N_10974,N_9168);
xnor U14966 (N_14966,N_8200,N_11451);
nand U14967 (N_14967,N_10260,N_11020);
nand U14968 (N_14968,N_8270,N_10244);
nor U14969 (N_14969,N_10179,N_10103);
nor U14970 (N_14970,N_10823,N_8696);
xor U14971 (N_14971,N_8522,N_8372);
nor U14972 (N_14972,N_11694,N_11048);
xor U14973 (N_14973,N_8764,N_8581);
nand U14974 (N_14974,N_9605,N_8656);
xnor U14975 (N_14975,N_10142,N_10751);
nand U14976 (N_14976,N_11548,N_11373);
and U14977 (N_14977,N_9802,N_11134);
xor U14978 (N_14978,N_8207,N_9904);
or U14979 (N_14979,N_11446,N_8371);
or U14980 (N_14980,N_9808,N_10479);
or U14981 (N_14981,N_11862,N_8431);
or U14982 (N_14982,N_9425,N_8676);
or U14983 (N_14983,N_9197,N_8312);
and U14984 (N_14984,N_11707,N_11423);
xor U14985 (N_14985,N_9717,N_9346);
or U14986 (N_14986,N_11020,N_10882);
and U14987 (N_14987,N_11508,N_11419);
xnor U14988 (N_14988,N_8557,N_11509);
nor U14989 (N_14989,N_10066,N_8816);
xor U14990 (N_14990,N_10312,N_8929);
xnor U14991 (N_14991,N_9489,N_8391);
nor U14992 (N_14992,N_9816,N_10366);
nand U14993 (N_14993,N_9877,N_10747);
xor U14994 (N_14994,N_8266,N_9197);
xnor U14995 (N_14995,N_8179,N_9985);
or U14996 (N_14996,N_11845,N_10551);
xor U14997 (N_14997,N_9279,N_8782);
xor U14998 (N_14998,N_10498,N_10233);
and U14999 (N_14999,N_11149,N_8755);
and U15000 (N_15000,N_9195,N_8012);
nor U15001 (N_15001,N_11025,N_9873);
nand U15002 (N_15002,N_8047,N_11055);
and U15003 (N_15003,N_11232,N_8518);
nand U15004 (N_15004,N_10223,N_9093);
or U15005 (N_15005,N_9694,N_9036);
nor U15006 (N_15006,N_8027,N_8020);
nor U15007 (N_15007,N_10217,N_9104);
and U15008 (N_15008,N_9134,N_11712);
nor U15009 (N_15009,N_9005,N_11193);
nand U15010 (N_15010,N_11693,N_8654);
nor U15011 (N_15011,N_11914,N_10990);
xnor U15012 (N_15012,N_11209,N_8343);
and U15013 (N_15013,N_11670,N_9778);
xor U15014 (N_15014,N_9810,N_10278);
xor U15015 (N_15015,N_8501,N_10224);
and U15016 (N_15016,N_11849,N_8895);
nand U15017 (N_15017,N_9287,N_9050);
xor U15018 (N_15018,N_8202,N_8904);
and U15019 (N_15019,N_11906,N_11104);
nand U15020 (N_15020,N_8195,N_10644);
or U15021 (N_15021,N_11115,N_11160);
nand U15022 (N_15022,N_11951,N_10330);
and U15023 (N_15023,N_10966,N_11700);
xnor U15024 (N_15024,N_9962,N_10166);
and U15025 (N_15025,N_10624,N_10199);
or U15026 (N_15026,N_10967,N_11134);
xor U15027 (N_15027,N_8809,N_9254);
nand U15028 (N_15028,N_8747,N_9886);
and U15029 (N_15029,N_9500,N_11005);
xor U15030 (N_15030,N_11753,N_8614);
and U15031 (N_15031,N_11742,N_9304);
nand U15032 (N_15032,N_8090,N_8518);
or U15033 (N_15033,N_8034,N_11244);
or U15034 (N_15034,N_10772,N_10756);
or U15035 (N_15035,N_11291,N_8773);
and U15036 (N_15036,N_10477,N_9726);
nand U15037 (N_15037,N_10045,N_10571);
or U15038 (N_15038,N_8798,N_10380);
xor U15039 (N_15039,N_11838,N_8388);
nand U15040 (N_15040,N_10763,N_9525);
or U15041 (N_15041,N_10049,N_9709);
nor U15042 (N_15042,N_11959,N_10736);
and U15043 (N_15043,N_9896,N_11288);
nor U15044 (N_15044,N_9186,N_11292);
nor U15045 (N_15045,N_8790,N_11526);
nand U15046 (N_15046,N_11407,N_10941);
nor U15047 (N_15047,N_10627,N_9510);
or U15048 (N_15048,N_10902,N_8050);
nor U15049 (N_15049,N_10311,N_8175);
nand U15050 (N_15050,N_8012,N_9229);
nand U15051 (N_15051,N_9494,N_9061);
and U15052 (N_15052,N_11747,N_11729);
xor U15053 (N_15053,N_11096,N_9663);
nand U15054 (N_15054,N_11086,N_9341);
or U15055 (N_15055,N_11336,N_10976);
or U15056 (N_15056,N_8691,N_8257);
nor U15057 (N_15057,N_8302,N_8756);
xnor U15058 (N_15058,N_11929,N_10434);
and U15059 (N_15059,N_11958,N_10937);
xnor U15060 (N_15060,N_10232,N_11727);
xor U15061 (N_15061,N_11966,N_8838);
nand U15062 (N_15062,N_8997,N_8009);
nand U15063 (N_15063,N_11686,N_8314);
or U15064 (N_15064,N_9812,N_11105);
nor U15065 (N_15065,N_10302,N_10090);
and U15066 (N_15066,N_8434,N_9630);
nand U15067 (N_15067,N_10326,N_9020);
and U15068 (N_15068,N_8187,N_9598);
nor U15069 (N_15069,N_8813,N_9319);
and U15070 (N_15070,N_9619,N_8753);
or U15071 (N_15071,N_8339,N_11424);
nor U15072 (N_15072,N_9360,N_8939);
and U15073 (N_15073,N_10883,N_8262);
or U15074 (N_15074,N_10750,N_11572);
nor U15075 (N_15075,N_11767,N_8172);
nand U15076 (N_15076,N_10953,N_11143);
xor U15077 (N_15077,N_9811,N_11735);
xor U15078 (N_15078,N_8603,N_11125);
nor U15079 (N_15079,N_9963,N_8825);
or U15080 (N_15080,N_9917,N_8668);
and U15081 (N_15081,N_8446,N_10959);
nand U15082 (N_15082,N_11898,N_11197);
nand U15083 (N_15083,N_9908,N_11305);
or U15084 (N_15084,N_11097,N_11942);
nor U15085 (N_15085,N_9410,N_8322);
xor U15086 (N_15086,N_9862,N_10355);
nand U15087 (N_15087,N_11070,N_11532);
nor U15088 (N_15088,N_9113,N_11454);
and U15089 (N_15089,N_10271,N_10471);
nor U15090 (N_15090,N_10768,N_8470);
xor U15091 (N_15091,N_8917,N_11650);
xnor U15092 (N_15092,N_10414,N_10452);
or U15093 (N_15093,N_10441,N_10723);
and U15094 (N_15094,N_8220,N_8419);
and U15095 (N_15095,N_10277,N_9232);
nand U15096 (N_15096,N_8805,N_8790);
nand U15097 (N_15097,N_8705,N_9479);
or U15098 (N_15098,N_11895,N_9782);
and U15099 (N_15099,N_8332,N_11678);
nor U15100 (N_15100,N_11802,N_10366);
nor U15101 (N_15101,N_8061,N_8487);
nor U15102 (N_15102,N_9910,N_11092);
nand U15103 (N_15103,N_11656,N_9070);
nand U15104 (N_15104,N_8014,N_9966);
nand U15105 (N_15105,N_10676,N_8769);
nor U15106 (N_15106,N_8536,N_9140);
nand U15107 (N_15107,N_11885,N_10224);
or U15108 (N_15108,N_8571,N_11509);
xor U15109 (N_15109,N_8235,N_8791);
nor U15110 (N_15110,N_8098,N_11287);
and U15111 (N_15111,N_8288,N_11272);
or U15112 (N_15112,N_8564,N_11554);
nor U15113 (N_15113,N_8093,N_10943);
nor U15114 (N_15114,N_10948,N_9099);
nor U15115 (N_15115,N_10549,N_8209);
or U15116 (N_15116,N_11811,N_8053);
xor U15117 (N_15117,N_8529,N_11871);
nor U15118 (N_15118,N_9393,N_11302);
xnor U15119 (N_15119,N_10364,N_8954);
xnor U15120 (N_15120,N_8861,N_11921);
nand U15121 (N_15121,N_8125,N_8326);
nand U15122 (N_15122,N_10070,N_11210);
xor U15123 (N_15123,N_10385,N_10357);
xor U15124 (N_15124,N_11565,N_9480);
xnor U15125 (N_15125,N_8984,N_10329);
xor U15126 (N_15126,N_11823,N_11293);
xnor U15127 (N_15127,N_9699,N_10113);
nor U15128 (N_15128,N_9766,N_11720);
nor U15129 (N_15129,N_8335,N_8075);
or U15130 (N_15130,N_11904,N_11782);
or U15131 (N_15131,N_11205,N_11708);
or U15132 (N_15132,N_8648,N_10543);
or U15133 (N_15133,N_8190,N_8022);
and U15134 (N_15134,N_9558,N_11602);
or U15135 (N_15135,N_11270,N_8472);
and U15136 (N_15136,N_8311,N_8193);
xnor U15137 (N_15137,N_8497,N_9499);
and U15138 (N_15138,N_8973,N_8810);
nand U15139 (N_15139,N_10227,N_11034);
nor U15140 (N_15140,N_11449,N_10886);
xnor U15141 (N_15141,N_11283,N_9783);
nand U15142 (N_15142,N_11631,N_10223);
nand U15143 (N_15143,N_9110,N_11675);
or U15144 (N_15144,N_10631,N_9609);
or U15145 (N_15145,N_10894,N_11309);
and U15146 (N_15146,N_9582,N_10484);
nand U15147 (N_15147,N_11972,N_10151);
and U15148 (N_15148,N_10060,N_11208);
xnor U15149 (N_15149,N_10581,N_8497);
and U15150 (N_15150,N_10971,N_8967);
nand U15151 (N_15151,N_10228,N_10487);
xor U15152 (N_15152,N_11119,N_8712);
xnor U15153 (N_15153,N_10075,N_8140);
nor U15154 (N_15154,N_11476,N_9663);
nor U15155 (N_15155,N_10115,N_10590);
or U15156 (N_15156,N_10826,N_9667);
or U15157 (N_15157,N_11312,N_11654);
xnor U15158 (N_15158,N_9402,N_9737);
xor U15159 (N_15159,N_10499,N_8325);
xor U15160 (N_15160,N_10493,N_11570);
xnor U15161 (N_15161,N_8648,N_11150);
nand U15162 (N_15162,N_8627,N_9001);
and U15163 (N_15163,N_10791,N_10932);
nor U15164 (N_15164,N_8791,N_8717);
nor U15165 (N_15165,N_10203,N_9403);
xnor U15166 (N_15166,N_8531,N_11099);
or U15167 (N_15167,N_8412,N_9784);
xnor U15168 (N_15168,N_10298,N_9080);
xor U15169 (N_15169,N_8169,N_10817);
nor U15170 (N_15170,N_8038,N_9702);
nor U15171 (N_15171,N_8185,N_11017);
nor U15172 (N_15172,N_9485,N_9832);
xnor U15173 (N_15173,N_11707,N_8009);
nor U15174 (N_15174,N_10885,N_8372);
or U15175 (N_15175,N_10063,N_8740);
and U15176 (N_15176,N_8841,N_8453);
nor U15177 (N_15177,N_11576,N_9870);
xor U15178 (N_15178,N_8323,N_11904);
xnor U15179 (N_15179,N_11906,N_10129);
xor U15180 (N_15180,N_10306,N_11956);
and U15181 (N_15181,N_9783,N_9000);
and U15182 (N_15182,N_9316,N_8296);
or U15183 (N_15183,N_11038,N_11803);
nand U15184 (N_15184,N_8449,N_11874);
and U15185 (N_15185,N_10084,N_10319);
and U15186 (N_15186,N_11839,N_8298);
nand U15187 (N_15187,N_9802,N_10818);
nand U15188 (N_15188,N_11260,N_10847);
and U15189 (N_15189,N_8284,N_8288);
nand U15190 (N_15190,N_9741,N_11876);
nand U15191 (N_15191,N_9534,N_10998);
and U15192 (N_15192,N_10226,N_10526);
or U15193 (N_15193,N_8270,N_10487);
nand U15194 (N_15194,N_11909,N_8774);
nor U15195 (N_15195,N_10925,N_11572);
nor U15196 (N_15196,N_8209,N_8881);
nand U15197 (N_15197,N_11060,N_11000);
xor U15198 (N_15198,N_8934,N_11421);
nand U15199 (N_15199,N_11481,N_8685);
xnor U15200 (N_15200,N_11613,N_8942);
xor U15201 (N_15201,N_11012,N_8112);
nor U15202 (N_15202,N_10158,N_11945);
and U15203 (N_15203,N_10254,N_11231);
xnor U15204 (N_15204,N_8331,N_8997);
or U15205 (N_15205,N_10370,N_11465);
or U15206 (N_15206,N_9420,N_8544);
nor U15207 (N_15207,N_10611,N_8051);
nor U15208 (N_15208,N_10416,N_9761);
xnor U15209 (N_15209,N_10454,N_10673);
xor U15210 (N_15210,N_10783,N_10310);
and U15211 (N_15211,N_9080,N_9307);
nor U15212 (N_15212,N_8561,N_10711);
nor U15213 (N_15213,N_8768,N_11574);
nand U15214 (N_15214,N_10213,N_11626);
or U15215 (N_15215,N_10079,N_8090);
or U15216 (N_15216,N_8702,N_10417);
and U15217 (N_15217,N_8158,N_9827);
xnor U15218 (N_15218,N_8393,N_10329);
nand U15219 (N_15219,N_10864,N_11482);
or U15220 (N_15220,N_10227,N_9807);
and U15221 (N_15221,N_11515,N_10690);
nand U15222 (N_15222,N_8606,N_10094);
nand U15223 (N_15223,N_10914,N_10262);
nand U15224 (N_15224,N_8751,N_11692);
or U15225 (N_15225,N_10606,N_8971);
xnor U15226 (N_15226,N_9538,N_8026);
nand U15227 (N_15227,N_8784,N_11048);
and U15228 (N_15228,N_8395,N_9839);
nor U15229 (N_15229,N_9949,N_8186);
and U15230 (N_15230,N_8036,N_9132);
or U15231 (N_15231,N_10457,N_10146);
xnor U15232 (N_15232,N_9363,N_8342);
nor U15233 (N_15233,N_10995,N_11629);
and U15234 (N_15234,N_8929,N_11034);
or U15235 (N_15235,N_10896,N_9922);
or U15236 (N_15236,N_10813,N_10632);
and U15237 (N_15237,N_10457,N_10207);
nand U15238 (N_15238,N_10378,N_11705);
nor U15239 (N_15239,N_8798,N_9148);
or U15240 (N_15240,N_9653,N_9694);
or U15241 (N_15241,N_11296,N_10276);
or U15242 (N_15242,N_9290,N_8436);
nor U15243 (N_15243,N_9959,N_10630);
nand U15244 (N_15244,N_11478,N_9457);
or U15245 (N_15245,N_10209,N_11755);
and U15246 (N_15246,N_10631,N_9859);
xor U15247 (N_15247,N_11669,N_8699);
and U15248 (N_15248,N_9579,N_10892);
or U15249 (N_15249,N_11390,N_10032);
xnor U15250 (N_15250,N_9250,N_9930);
or U15251 (N_15251,N_10332,N_11820);
nor U15252 (N_15252,N_10280,N_8780);
nor U15253 (N_15253,N_8668,N_8419);
xnor U15254 (N_15254,N_8974,N_11670);
or U15255 (N_15255,N_8410,N_11261);
or U15256 (N_15256,N_8242,N_8314);
or U15257 (N_15257,N_9430,N_11343);
nor U15258 (N_15258,N_11971,N_9353);
and U15259 (N_15259,N_11817,N_8201);
and U15260 (N_15260,N_10623,N_8638);
xnor U15261 (N_15261,N_8066,N_8835);
nor U15262 (N_15262,N_10711,N_11220);
nand U15263 (N_15263,N_8527,N_10647);
and U15264 (N_15264,N_11966,N_10863);
and U15265 (N_15265,N_10542,N_11181);
or U15266 (N_15266,N_8623,N_9430);
and U15267 (N_15267,N_10639,N_9993);
nand U15268 (N_15268,N_10638,N_10068);
or U15269 (N_15269,N_8317,N_10634);
or U15270 (N_15270,N_8425,N_11337);
and U15271 (N_15271,N_8245,N_11050);
xnor U15272 (N_15272,N_11240,N_11365);
and U15273 (N_15273,N_10709,N_8110);
nand U15274 (N_15274,N_11361,N_9386);
nand U15275 (N_15275,N_11256,N_11141);
and U15276 (N_15276,N_10068,N_8934);
nand U15277 (N_15277,N_11686,N_8466);
and U15278 (N_15278,N_11888,N_11040);
nand U15279 (N_15279,N_9763,N_9186);
xor U15280 (N_15280,N_10453,N_11526);
or U15281 (N_15281,N_9573,N_8574);
nor U15282 (N_15282,N_8217,N_10283);
and U15283 (N_15283,N_9840,N_9677);
xnor U15284 (N_15284,N_10121,N_11732);
or U15285 (N_15285,N_9838,N_9404);
nor U15286 (N_15286,N_9849,N_8522);
and U15287 (N_15287,N_9960,N_9665);
nand U15288 (N_15288,N_8263,N_9132);
and U15289 (N_15289,N_8063,N_11432);
and U15290 (N_15290,N_9442,N_10717);
and U15291 (N_15291,N_10027,N_10781);
nand U15292 (N_15292,N_9407,N_9995);
nor U15293 (N_15293,N_10731,N_9009);
nor U15294 (N_15294,N_9730,N_8179);
nor U15295 (N_15295,N_9841,N_9930);
nand U15296 (N_15296,N_10481,N_8815);
xnor U15297 (N_15297,N_9772,N_10356);
xor U15298 (N_15298,N_9367,N_9060);
xnor U15299 (N_15299,N_11346,N_11886);
nor U15300 (N_15300,N_10485,N_11286);
xnor U15301 (N_15301,N_11957,N_8805);
and U15302 (N_15302,N_11917,N_9552);
or U15303 (N_15303,N_11081,N_11998);
xor U15304 (N_15304,N_10558,N_9491);
or U15305 (N_15305,N_10371,N_11030);
or U15306 (N_15306,N_9896,N_9248);
and U15307 (N_15307,N_8849,N_10302);
and U15308 (N_15308,N_11840,N_8300);
and U15309 (N_15309,N_11234,N_10825);
xnor U15310 (N_15310,N_11015,N_10227);
nand U15311 (N_15311,N_10343,N_10873);
and U15312 (N_15312,N_10726,N_10464);
nand U15313 (N_15313,N_9307,N_9741);
nor U15314 (N_15314,N_11071,N_8955);
and U15315 (N_15315,N_11058,N_9447);
nand U15316 (N_15316,N_11499,N_11213);
and U15317 (N_15317,N_9928,N_10253);
and U15318 (N_15318,N_9931,N_9152);
and U15319 (N_15319,N_9734,N_10199);
xor U15320 (N_15320,N_10401,N_9418);
nor U15321 (N_15321,N_9115,N_9476);
or U15322 (N_15322,N_11960,N_9418);
nor U15323 (N_15323,N_11680,N_8313);
nand U15324 (N_15324,N_11025,N_11013);
or U15325 (N_15325,N_8844,N_10770);
xnor U15326 (N_15326,N_11297,N_11045);
nand U15327 (N_15327,N_9703,N_9942);
nor U15328 (N_15328,N_11442,N_8351);
or U15329 (N_15329,N_8558,N_9247);
xor U15330 (N_15330,N_10211,N_9287);
nand U15331 (N_15331,N_11875,N_9172);
nand U15332 (N_15332,N_11940,N_8110);
nor U15333 (N_15333,N_8903,N_9353);
and U15334 (N_15334,N_8528,N_9982);
and U15335 (N_15335,N_11022,N_8320);
xor U15336 (N_15336,N_8942,N_10917);
or U15337 (N_15337,N_10039,N_10527);
and U15338 (N_15338,N_10524,N_9451);
and U15339 (N_15339,N_11468,N_9454);
nand U15340 (N_15340,N_9666,N_10098);
nand U15341 (N_15341,N_10892,N_8533);
and U15342 (N_15342,N_10569,N_11960);
nand U15343 (N_15343,N_9317,N_11751);
nor U15344 (N_15344,N_11063,N_9418);
and U15345 (N_15345,N_10806,N_9083);
nor U15346 (N_15346,N_9599,N_9002);
xor U15347 (N_15347,N_11238,N_11205);
or U15348 (N_15348,N_10086,N_8439);
or U15349 (N_15349,N_11167,N_8923);
nand U15350 (N_15350,N_9938,N_11212);
and U15351 (N_15351,N_11813,N_10323);
and U15352 (N_15352,N_9427,N_11462);
and U15353 (N_15353,N_9968,N_8402);
nand U15354 (N_15354,N_10056,N_9540);
nand U15355 (N_15355,N_11200,N_10516);
nor U15356 (N_15356,N_8234,N_11000);
nand U15357 (N_15357,N_9036,N_10353);
nand U15358 (N_15358,N_9382,N_8968);
xnor U15359 (N_15359,N_11399,N_11132);
xor U15360 (N_15360,N_8521,N_8161);
or U15361 (N_15361,N_8870,N_11395);
nor U15362 (N_15362,N_11850,N_9177);
nor U15363 (N_15363,N_10137,N_8697);
xnor U15364 (N_15364,N_10741,N_9237);
or U15365 (N_15365,N_8410,N_11290);
nand U15366 (N_15366,N_10312,N_9434);
and U15367 (N_15367,N_10348,N_9780);
nor U15368 (N_15368,N_8645,N_11028);
nand U15369 (N_15369,N_10658,N_11335);
xnor U15370 (N_15370,N_8247,N_11648);
or U15371 (N_15371,N_9201,N_9727);
nand U15372 (N_15372,N_10626,N_8875);
or U15373 (N_15373,N_10435,N_11302);
or U15374 (N_15374,N_8026,N_8392);
nand U15375 (N_15375,N_9241,N_9232);
nor U15376 (N_15376,N_10323,N_8834);
or U15377 (N_15377,N_9693,N_11138);
xor U15378 (N_15378,N_9531,N_8881);
or U15379 (N_15379,N_8458,N_9926);
nand U15380 (N_15380,N_9318,N_10552);
nand U15381 (N_15381,N_11075,N_8197);
or U15382 (N_15382,N_11935,N_10008);
nand U15383 (N_15383,N_8657,N_9852);
nor U15384 (N_15384,N_10167,N_8327);
and U15385 (N_15385,N_10007,N_8163);
nand U15386 (N_15386,N_9129,N_8159);
xnor U15387 (N_15387,N_11967,N_11936);
nand U15388 (N_15388,N_9435,N_11426);
and U15389 (N_15389,N_10578,N_8823);
or U15390 (N_15390,N_11420,N_11055);
nand U15391 (N_15391,N_8011,N_9716);
or U15392 (N_15392,N_9464,N_10720);
nor U15393 (N_15393,N_10410,N_10572);
nor U15394 (N_15394,N_10684,N_9310);
and U15395 (N_15395,N_11608,N_11106);
nand U15396 (N_15396,N_9023,N_11959);
and U15397 (N_15397,N_8295,N_9348);
nor U15398 (N_15398,N_10940,N_10047);
xnor U15399 (N_15399,N_9641,N_8470);
and U15400 (N_15400,N_10811,N_10278);
xor U15401 (N_15401,N_10198,N_11885);
or U15402 (N_15402,N_8641,N_11671);
nand U15403 (N_15403,N_8110,N_11220);
and U15404 (N_15404,N_8192,N_10958);
or U15405 (N_15405,N_10790,N_10466);
and U15406 (N_15406,N_8384,N_11891);
or U15407 (N_15407,N_8429,N_9661);
nand U15408 (N_15408,N_10023,N_8478);
xor U15409 (N_15409,N_11621,N_11173);
xnor U15410 (N_15410,N_9295,N_10262);
or U15411 (N_15411,N_10401,N_8551);
nor U15412 (N_15412,N_11768,N_9806);
and U15413 (N_15413,N_11237,N_10137);
xnor U15414 (N_15414,N_9550,N_11809);
xnor U15415 (N_15415,N_9250,N_9842);
or U15416 (N_15416,N_10232,N_11397);
or U15417 (N_15417,N_8078,N_10453);
xor U15418 (N_15418,N_11832,N_10796);
nor U15419 (N_15419,N_9458,N_10630);
or U15420 (N_15420,N_10292,N_11183);
and U15421 (N_15421,N_11832,N_10561);
xnor U15422 (N_15422,N_11611,N_9951);
nor U15423 (N_15423,N_8038,N_8646);
or U15424 (N_15424,N_10711,N_10979);
nand U15425 (N_15425,N_10698,N_11030);
xnor U15426 (N_15426,N_8115,N_9042);
nand U15427 (N_15427,N_10698,N_8880);
xnor U15428 (N_15428,N_9395,N_10560);
xor U15429 (N_15429,N_9795,N_9791);
and U15430 (N_15430,N_8794,N_8324);
nand U15431 (N_15431,N_10460,N_8275);
and U15432 (N_15432,N_11613,N_8030);
nor U15433 (N_15433,N_9522,N_8275);
xnor U15434 (N_15434,N_10396,N_8293);
xor U15435 (N_15435,N_10403,N_8339);
xnor U15436 (N_15436,N_11180,N_9456);
xnor U15437 (N_15437,N_11480,N_8008);
xor U15438 (N_15438,N_10218,N_8040);
and U15439 (N_15439,N_9504,N_9278);
or U15440 (N_15440,N_11914,N_11447);
or U15441 (N_15441,N_11314,N_8220);
nand U15442 (N_15442,N_9571,N_10511);
and U15443 (N_15443,N_10217,N_9012);
nor U15444 (N_15444,N_9321,N_10013);
or U15445 (N_15445,N_11398,N_8864);
and U15446 (N_15446,N_8944,N_11759);
and U15447 (N_15447,N_8950,N_10296);
or U15448 (N_15448,N_9078,N_9954);
nor U15449 (N_15449,N_11489,N_8370);
nor U15450 (N_15450,N_8627,N_9903);
or U15451 (N_15451,N_8425,N_8419);
and U15452 (N_15452,N_9871,N_11037);
nand U15453 (N_15453,N_8485,N_8319);
and U15454 (N_15454,N_11013,N_8308);
nand U15455 (N_15455,N_9381,N_9923);
nand U15456 (N_15456,N_11083,N_8659);
xor U15457 (N_15457,N_11705,N_9815);
or U15458 (N_15458,N_8692,N_11138);
xnor U15459 (N_15459,N_9618,N_10550);
or U15460 (N_15460,N_9913,N_8119);
xor U15461 (N_15461,N_9919,N_9356);
and U15462 (N_15462,N_11544,N_8243);
or U15463 (N_15463,N_10216,N_8387);
or U15464 (N_15464,N_8087,N_11906);
nor U15465 (N_15465,N_9187,N_8261);
and U15466 (N_15466,N_8433,N_10501);
or U15467 (N_15467,N_8080,N_10716);
or U15468 (N_15468,N_11698,N_9750);
nor U15469 (N_15469,N_10266,N_10975);
and U15470 (N_15470,N_10748,N_8596);
xor U15471 (N_15471,N_10044,N_10838);
nand U15472 (N_15472,N_9522,N_9158);
nand U15473 (N_15473,N_8856,N_9390);
nand U15474 (N_15474,N_10857,N_10291);
or U15475 (N_15475,N_9283,N_8769);
nor U15476 (N_15476,N_11315,N_10368);
and U15477 (N_15477,N_11875,N_10529);
or U15478 (N_15478,N_11863,N_8220);
nor U15479 (N_15479,N_8342,N_9385);
nor U15480 (N_15480,N_8350,N_9074);
xor U15481 (N_15481,N_10781,N_11161);
or U15482 (N_15482,N_11220,N_8029);
nor U15483 (N_15483,N_10239,N_10495);
nor U15484 (N_15484,N_8681,N_8778);
nor U15485 (N_15485,N_10439,N_10263);
nand U15486 (N_15486,N_11717,N_11309);
nor U15487 (N_15487,N_11566,N_9947);
or U15488 (N_15488,N_10803,N_11617);
xnor U15489 (N_15489,N_10488,N_8074);
nor U15490 (N_15490,N_10763,N_10227);
or U15491 (N_15491,N_11202,N_10332);
nand U15492 (N_15492,N_10310,N_10941);
nand U15493 (N_15493,N_11202,N_11995);
xnor U15494 (N_15494,N_11783,N_8204);
nand U15495 (N_15495,N_9161,N_8091);
and U15496 (N_15496,N_9012,N_10340);
and U15497 (N_15497,N_8761,N_9825);
nand U15498 (N_15498,N_11286,N_8355);
nand U15499 (N_15499,N_11658,N_8196);
and U15500 (N_15500,N_8940,N_8656);
and U15501 (N_15501,N_8191,N_10276);
xnor U15502 (N_15502,N_11693,N_10824);
nor U15503 (N_15503,N_11847,N_11875);
nand U15504 (N_15504,N_10426,N_10969);
and U15505 (N_15505,N_9103,N_8893);
xor U15506 (N_15506,N_11160,N_10384);
nand U15507 (N_15507,N_11577,N_8695);
and U15508 (N_15508,N_8976,N_8911);
xnor U15509 (N_15509,N_10885,N_8654);
and U15510 (N_15510,N_8533,N_9849);
or U15511 (N_15511,N_10135,N_9063);
xnor U15512 (N_15512,N_11610,N_9754);
and U15513 (N_15513,N_10885,N_11527);
nand U15514 (N_15514,N_10057,N_11673);
or U15515 (N_15515,N_9537,N_10754);
nor U15516 (N_15516,N_8393,N_9308);
and U15517 (N_15517,N_10234,N_11110);
nor U15518 (N_15518,N_8774,N_11103);
xnor U15519 (N_15519,N_10474,N_9960);
nor U15520 (N_15520,N_10236,N_8770);
nor U15521 (N_15521,N_9644,N_10584);
nor U15522 (N_15522,N_9465,N_11437);
xor U15523 (N_15523,N_10467,N_10830);
nor U15524 (N_15524,N_10236,N_8894);
nor U15525 (N_15525,N_10507,N_11520);
xor U15526 (N_15526,N_11532,N_11958);
or U15527 (N_15527,N_10996,N_9451);
nand U15528 (N_15528,N_11504,N_9545);
nor U15529 (N_15529,N_11445,N_10280);
nor U15530 (N_15530,N_9403,N_10637);
nor U15531 (N_15531,N_8511,N_11234);
nor U15532 (N_15532,N_9472,N_10438);
and U15533 (N_15533,N_10901,N_11123);
nand U15534 (N_15534,N_9282,N_9763);
or U15535 (N_15535,N_11334,N_10634);
nand U15536 (N_15536,N_9068,N_10117);
xnor U15537 (N_15537,N_9920,N_9669);
nand U15538 (N_15538,N_11644,N_11610);
xor U15539 (N_15539,N_11554,N_11828);
and U15540 (N_15540,N_8999,N_11711);
and U15541 (N_15541,N_8284,N_10142);
nand U15542 (N_15542,N_10605,N_10093);
nand U15543 (N_15543,N_11683,N_10215);
xnor U15544 (N_15544,N_11159,N_10199);
nor U15545 (N_15545,N_11324,N_8125);
and U15546 (N_15546,N_11070,N_11779);
nand U15547 (N_15547,N_11427,N_10726);
nor U15548 (N_15548,N_11985,N_10929);
nand U15549 (N_15549,N_9451,N_9699);
xnor U15550 (N_15550,N_10990,N_11794);
or U15551 (N_15551,N_8241,N_8149);
and U15552 (N_15552,N_9823,N_9046);
or U15553 (N_15553,N_9144,N_10870);
nor U15554 (N_15554,N_8118,N_8513);
nor U15555 (N_15555,N_9391,N_10925);
nor U15556 (N_15556,N_11900,N_8100);
xnor U15557 (N_15557,N_11207,N_9354);
nor U15558 (N_15558,N_10504,N_9223);
nand U15559 (N_15559,N_10366,N_10044);
and U15560 (N_15560,N_10947,N_10297);
nand U15561 (N_15561,N_8428,N_11642);
nor U15562 (N_15562,N_9065,N_9116);
nand U15563 (N_15563,N_8766,N_11095);
nor U15564 (N_15564,N_10610,N_9762);
nor U15565 (N_15565,N_8752,N_9650);
and U15566 (N_15566,N_10128,N_9110);
nor U15567 (N_15567,N_10586,N_9828);
nor U15568 (N_15568,N_8998,N_9331);
nor U15569 (N_15569,N_11451,N_10724);
or U15570 (N_15570,N_8977,N_10519);
nor U15571 (N_15571,N_8454,N_11206);
and U15572 (N_15572,N_9398,N_11278);
and U15573 (N_15573,N_9787,N_8455);
or U15574 (N_15574,N_8919,N_8505);
nand U15575 (N_15575,N_9072,N_10389);
or U15576 (N_15576,N_11248,N_10746);
xor U15577 (N_15577,N_8842,N_10732);
and U15578 (N_15578,N_10011,N_11247);
xor U15579 (N_15579,N_9193,N_10164);
and U15580 (N_15580,N_11263,N_10226);
or U15581 (N_15581,N_9794,N_9111);
nor U15582 (N_15582,N_11797,N_10435);
and U15583 (N_15583,N_11609,N_11863);
nand U15584 (N_15584,N_8550,N_9876);
nor U15585 (N_15585,N_10549,N_9581);
nand U15586 (N_15586,N_8998,N_9350);
xor U15587 (N_15587,N_11475,N_9362);
nor U15588 (N_15588,N_8273,N_9666);
or U15589 (N_15589,N_8162,N_10982);
and U15590 (N_15590,N_8490,N_10108);
or U15591 (N_15591,N_8549,N_10409);
nor U15592 (N_15592,N_8259,N_8116);
xnor U15593 (N_15593,N_9960,N_8090);
nor U15594 (N_15594,N_11858,N_11268);
nor U15595 (N_15595,N_8985,N_9455);
xor U15596 (N_15596,N_11565,N_9159);
or U15597 (N_15597,N_9283,N_11183);
xor U15598 (N_15598,N_11521,N_9121);
and U15599 (N_15599,N_9485,N_10615);
nor U15600 (N_15600,N_11785,N_10468);
xnor U15601 (N_15601,N_8249,N_11244);
and U15602 (N_15602,N_10107,N_11265);
nand U15603 (N_15603,N_8609,N_9122);
xor U15604 (N_15604,N_11583,N_11965);
nand U15605 (N_15605,N_9882,N_8231);
and U15606 (N_15606,N_10707,N_10248);
nor U15607 (N_15607,N_8142,N_8510);
or U15608 (N_15608,N_11678,N_10658);
or U15609 (N_15609,N_10934,N_10411);
and U15610 (N_15610,N_8669,N_11104);
or U15611 (N_15611,N_11641,N_9019);
nor U15612 (N_15612,N_9429,N_8458);
nor U15613 (N_15613,N_11657,N_11712);
nand U15614 (N_15614,N_10704,N_9977);
or U15615 (N_15615,N_10901,N_11841);
nor U15616 (N_15616,N_9892,N_9593);
or U15617 (N_15617,N_9007,N_8784);
or U15618 (N_15618,N_9650,N_11625);
xor U15619 (N_15619,N_8846,N_8142);
nor U15620 (N_15620,N_9933,N_10304);
nand U15621 (N_15621,N_9371,N_8148);
nor U15622 (N_15622,N_9136,N_10801);
nor U15623 (N_15623,N_9904,N_10815);
and U15624 (N_15624,N_8763,N_8310);
or U15625 (N_15625,N_9198,N_8505);
or U15626 (N_15626,N_11465,N_9655);
nor U15627 (N_15627,N_10561,N_11133);
xnor U15628 (N_15628,N_10076,N_10690);
nand U15629 (N_15629,N_8601,N_11604);
and U15630 (N_15630,N_8465,N_10478);
nor U15631 (N_15631,N_8706,N_11104);
and U15632 (N_15632,N_11929,N_10378);
nand U15633 (N_15633,N_8237,N_8168);
nor U15634 (N_15634,N_11777,N_9208);
nand U15635 (N_15635,N_10789,N_11776);
xor U15636 (N_15636,N_8168,N_10154);
nor U15637 (N_15637,N_10693,N_8360);
nor U15638 (N_15638,N_8435,N_8224);
or U15639 (N_15639,N_8295,N_9533);
or U15640 (N_15640,N_9313,N_10264);
nor U15641 (N_15641,N_10706,N_10295);
or U15642 (N_15642,N_10582,N_10074);
nand U15643 (N_15643,N_8349,N_11457);
xor U15644 (N_15644,N_10877,N_11260);
or U15645 (N_15645,N_8843,N_9036);
xor U15646 (N_15646,N_11995,N_8149);
nor U15647 (N_15647,N_10826,N_10496);
and U15648 (N_15648,N_8301,N_10708);
or U15649 (N_15649,N_8662,N_8660);
xnor U15650 (N_15650,N_10591,N_11148);
nand U15651 (N_15651,N_10150,N_10552);
nand U15652 (N_15652,N_8061,N_11692);
xnor U15653 (N_15653,N_11035,N_11992);
nand U15654 (N_15654,N_10712,N_10942);
or U15655 (N_15655,N_8508,N_10455);
and U15656 (N_15656,N_9659,N_11327);
nor U15657 (N_15657,N_9642,N_11402);
nand U15658 (N_15658,N_10815,N_10313);
nand U15659 (N_15659,N_9199,N_10207);
nand U15660 (N_15660,N_9094,N_9597);
and U15661 (N_15661,N_10379,N_8000);
or U15662 (N_15662,N_9281,N_8287);
nor U15663 (N_15663,N_11331,N_8228);
nand U15664 (N_15664,N_9410,N_9350);
and U15665 (N_15665,N_10496,N_9372);
nor U15666 (N_15666,N_8452,N_11307);
and U15667 (N_15667,N_8860,N_9256);
or U15668 (N_15668,N_10715,N_9751);
nor U15669 (N_15669,N_11814,N_11455);
nand U15670 (N_15670,N_11242,N_10310);
nand U15671 (N_15671,N_8958,N_9274);
nor U15672 (N_15672,N_11702,N_10133);
or U15673 (N_15673,N_10975,N_11052);
xnor U15674 (N_15674,N_11183,N_11285);
nor U15675 (N_15675,N_8640,N_8041);
and U15676 (N_15676,N_8402,N_8716);
or U15677 (N_15677,N_9183,N_11050);
and U15678 (N_15678,N_11851,N_11350);
nand U15679 (N_15679,N_8192,N_9753);
and U15680 (N_15680,N_10030,N_8052);
and U15681 (N_15681,N_8138,N_9726);
nor U15682 (N_15682,N_11206,N_8213);
nand U15683 (N_15683,N_10614,N_8431);
nand U15684 (N_15684,N_10808,N_9684);
and U15685 (N_15685,N_8037,N_9726);
nor U15686 (N_15686,N_9563,N_10208);
and U15687 (N_15687,N_10220,N_11497);
xnor U15688 (N_15688,N_9506,N_11975);
xor U15689 (N_15689,N_11612,N_10901);
nand U15690 (N_15690,N_10929,N_9456);
nor U15691 (N_15691,N_10967,N_9436);
or U15692 (N_15692,N_9097,N_11906);
nor U15693 (N_15693,N_8160,N_10481);
or U15694 (N_15694,N_9708,N_11651);
and U15695 (N_15695,N_10952,N_9855);
or U15696 (N_15696,N_9438,N_11305);
nor U15697 (N_15697,N_8205,N_11660);
xor U15698 (N_15698,N_9901,N_8104);
nor U15699 (N_15699,N_11137,N_10158);
nor U15700 (N_15700,N_10846,N_11700);
xor U15701 (N_15701,N_11810,N_11337);
xor U15702 (N_15702,N_9996,N_8540);
nand U15703 (N_15703,N_11124,N_8446);
or U15704 (N_15704,N_9217,N_10037);
xnor U15705 (N_15705,N_8026,N_8714);
nor U15706 (N_15706,N_10405,N_10387);
nor U15707 (N_15707,N_11112,N_8487);
nor U15708 (N_15708,N_10128,N_11510);
and U15709 (N_15709,N_11978,N_9372);
nor U15710 (N_15710,N_8403,N_8151);
nor U15711 (N_15711,N_8967,N_10085);
and U15712 (N_15712,N_11751,N_9766);
nor U15713 (N_15713,N_9856,N_9085);
xor U15714 (N_15714,N_9550,N_9674);
xor U15715 (N_15715,N_11196,N_11763);
or U15716 (N_15716,N_10413,N_10393);
and U15717 (N_15717,N_8112,N_11526);
nor U15718 (N_15718,N_11363,N_10411);
and U15719 (N_15719,N_11429,N_10242);
xnor U15720 (N_15720,N_9839,N_8106);
and U15721 (N_15721,N_10306,N_9368);
nand U15722 (N_15722,N_10511,N_8693);
xor U15723 (N_15723,N_9769,N_9660);
xnor U15724 (N_15724,N_10658,N_8353);
or U15725 (N_15725,N_9974,N_9400);
nor U15726 (N_15726,N_9542,N_9471);
nor U15727 (N_15727,N_10957,N_11779);
xnor U15728 (N_15728,N_11803,N_8677);
xor U15729 (N_15729,N_8850,N_8385);
nor U15730 (N_15730,N_9995,N_10546);
nand U15731 (N_15731,N_11514,N_9337);
xor U15732 (N_15732,N_11059,N_11933);
xnor U15733 (N_15733,N_11806,N_10255);
or U15734 (N_15734,N_8665,N_9074);
nand U15735 (N_15735,N_8701,N_11057);
or U15736 (N_15736,N_10175,N_11187);
nand U15737 (N_15737,N_8023,N_11159);
and U15738 (N_15738,N_10444,N_8235);
xor U15739 (N_15739,N_10113,N_10368);
or U15740 (N_15740,N_11208,N_10588);
and U15741 (N_15741,N_11232,N_9152);
or U15742 (N_15742,N_10612,N_9991);
nor U15743 (N_15743,N_8710,N_9459);
xnor U15744 (N_15744,N_11067,N_11841);
nor U15745 (N_15745,N_10127,N_9364);
or U15746 (N_15746,N_8477,N_10193);
nor U15747 (N_15747,N_9984,N_10019);
or U15748 (N_15748,N_11441,N_9250);
nor U15749 (N_15749,N_9935,N_11646);
nand U15750 (N_15750,N_11668,N_10906);
and U15751 (N_15751,N_8201,N_11060);
nor U15752 (N_15752,N_9135,N_9078);
nor U15753 (N_15753,N_10956,N_9720);
or U15754 (N_15754,N_10719,N_11057);
or U15755 (N_15755,N_9309,N_11933);
nor U15756 (N_15756,N_9067,N_11356);
and U15757 (N_15757,N_9532,N_8239);
xor U15758 (N_15758,N_9526,N_8857);
and U15759 (N_15759,N_9026,N_9145);
and U15760 (N_15760,N_11598,N_11409);
xnor U15761 (N_15761,N_11298,N_11727);
nor U15762 (N_15762,N_8140,N_9820);
nor U15763 (N_15763,N_8581,N_11290);
nand U15764 (N_15764,N_8437,N_11972);
and U15765 (N_15765,N_10469,N_10865);
nor U15766 (N_15766,N_10249,N_10515);
xor U15767 (N_15767,N_9305,N_10931);
xnor U15768 (N_15768,N_8071,N_8410);
nor U15769 (N_15769,N_9982,N_11395);
and U15770 (N_15770,N_10530,N_9724);
nor U15771 (N_15771,N_10053,N_11587);
or U15772 (N_15772,N_8243,N_11974);
nand U15773 (N_15773,N_11806,N_10697);
nand U15774 (N_15774,N_9155,N_10748);
or U15775 (N_15775,N_8905,N_9111);
and U15776 (N_15776,N_10404,N_10351);
nor U15777 (N_15777,N_10924,N_11331);
and U15778 (N_15778,N_9212,N_10372);
nand U15779 (N_15779,N_8852,N_9735);
or U15780 (N_15780,N_8293,N_10623);
nand U15781 (N_15781,N_11411,N_10241);
xor U15782 (N_15782,N_8796,N_10141);
nor U15783 (N_15783,N_9650,N_8278);
xnor U15784 (N_15784,N_9119,N_11139);
nand U15785 (N_15785,N_9265,N_8166);
nand U15786 (N_15786,N_11244,N_10798);
or U15787 (N_15787,N_8624,N_8074);
nor U15788 (N_15788,N_8308,N_8214);
nor U15789 (N_15789,N_9251,N_9779);
nand U15790 (N_15790,N_8273,N_11253);
and U15791 (N_15791,N_11885,N_9604);
and U15792 (N_15792,N_11153,N_10944);
or U15793 (N_15793,N_9921,N_8922);
xnor U15794 (N_15794,N_10687,N_8277);
nand U15795 (N_15795,N_8011,N_8010);
xnor U15796 (N_15796,N_10526,N_11859);
and U15797 (N_15797,N_10326,N_9728);
or U15798 (N_15798,N_8531,N_11728);
nand U15799 (N_15799,N_8537,N_10393);
or U15800 (N_15800,N_9379,N_8391);
or U15801 (N_15801,N_11939,N_10778);
nand U15802 (N_15802,N_9794,N_11227);
and U15803 (N_15803,N_11239,N_10706);
or U15804 (N_15804,N_8358,N_9139);
and U15805 (N_15805,N_11924,N_8609);
and U15806 (N_15806,N_9544,N_11552);
and U15807 (N_15807,N_11200,N_10993);
nand U15808 (N_15808,N_10140,N_8735);
nor U15809 (N_15809,N_10568,N_11013);
nor U15810 (N_15810,N_10660,N_10055);
nor U15811 (N_15811,N_9560,N_10549);
nand U15812 (N_15812,N_9917,N_9175);
or U15813 (N_15813,N_9874,N_9074);
nand U15814 (N_15814,N_8248,N_9185);
nand U15815 (N_15815,N_9779,N_11492);
and U15816 (N_15816,N_8984,N_11556);
or U15817 (N_15817,N_9972,N_11703);
or U15818 (N_15818,N_11962,N_9128);
or U15819 (N_15819,N_10048,N_11702);
and U15820 (N_15820,N_10239,N_10218);
nand U15821 (N_15821,N_9228,N_8019);
nor U15822 (N_15822,N_10733,N_8454);
or U15823 (N_15823,N_9246,N_8699);
nor U15824 (N_15824,N_10962,N_11262);
xnor U15825 (N_15825,N_10623,N_11765);
nor U15826 (N_15826,N_8575,N_10133);
or U15827 (N_15827,N_10272,N_10017);
xor U15828 (N_15828,N_11515,N_11125);
and U15829 (N_15829,N_8353,N_8965);
and U15830 (N_15830,N_10662,N_9268);
xor U15831 (N_15831,N_10210,N_9277);
or U15832 (N_15832,N_10558,N_10248);
xor U15833 (N_15833,N_8169,N_10399);
or U15834 (N_15834,N_8456,N_11687);
or U15835 (N_15835,N_9653,N_11669);
nand U15836 (N_15836,N_8885,N_8607);
and U15837 (N_15837,N_10983,N_9076);
and U15838 (N_15838,N_10711,N_10608);
xnor U15839 (N_15839,N_10715,N_11785);
xnor U15840 (N_15840,N_8457,N_9229);
or U15841 (N_15841,N_9043,N_11428);
nor U15842 (N_15842,N_10335,N_8053);
nand U15843 (N_15843,N_8546,N_10464);
xor U15844 (N_15844,N_11587,N_8655);
xnor U15845 (N_15845,N_11309,N_8622);
nor U15846 (N_15846,N_10805,N_11729);
or U15847 (N_15847,N_8234,N_10409);
xnor U15848 (N_15848,N_10193,N_9635);
nor U15849 (N_15849,N_10657,N_10802);
xor U15850 (N_15850,N_9863,N_8976);
and U15851 (N_15851,N_10742,N_9664);
nand U15852 (N_15852,N_11839,N_8582);
or U15853 (N_15853,N_11673,N_8009);
nor U15854 (N_15854,N_10886,N_8320);
nor U15855 (N_15855,N_8585,N_9888);
or U15856 (N_15856,N_9080,N_8536);
or U15857 (N_15857,N_8868,N_11934);
nor U15858 (N_15858,N_9194,N_11177);
or U15859 (N_15859,N_9414,N_10641);
xnor U15860 (N_15860,N_10298,N_10466);
nand U15861 (N_15861,N_11166,N_11600);
xor U15862 (N_15862,N_8984,N_8908);
nand U15863 (N_15863,N_11362,N_10354);
nor U15864 (N_15864,N_11629,N_10445);
xor U15865 (N_15865,N_8501,N_9688);
nor U15866 (N_15866,N_11193,N_8075);
nor U15867 (N_15867,N_11985,N_9403);
nor U15868 (N_15868,N_11468,N_8549);
or U15869 (N_15869,N_8570,N_8144);
or U15870 (N_15870,N_10191,N_9475);
nor U15871 (N_15871,N_11685,N_9708);
nor U15872 (N_15872,N_11310,N_9294);
xnor U15873 (N_15873,N_9853,N_10415);
and U15874 (N_15874,N_11204,N_9855);
nand U15875 (N_15875,N_10703,N_10537);
xor U15876 (N_15876,N_11726,N_11642);
or U15877 (N_15877,N_8840,N_10693);
and U15878 (N_15878,N_9752,N_10990);
nor U15879 (N_15879,N_11639,N_9301);
or U15880 (N_15880,N_10156,N_10921);
nand U15881 (N_15881,N_9722,N_11720);
or U15882 (N_15882,N_9750,N_8175);
nor U15883 (N_15883,N_10649,N_9809);
xnor U15884 (N_15884,N_10937,N_8973);
or U15885 (N_15885,N_11330,N_9542);
and U15886 (N_15886,N_11883,N_8903);
nor U15887 (N_15887,N_11306,N_11492);
or U15888 (N_15888,N_10597,N_8143);
nor U15889 (N_15889,N_11156,N_10265);
and U15890 (N_15890,N_10529,N_11199);
xnor U15891 (N_15891,N_11581,N_8279);
xnor U15892 (N_15892,N_11908,N_11579);
nor U15893 (N_15893,N_8557,N_8748);
and U15894 (N_15894,N_10352,N_9406);
nand U15895 (N_15895,N_9127,N_11807);
nand U15896 (N_15896,N_9514,N_11272);
nand U15897 (N_15897,N_10656,N_10970);
and U15898 (N_15898,N_10867,N_10370);
or U15899 (N_15899,N_9651,N_9957);
nor U15900 (N_15900,N_11524,N_11112);
and U15901 (N_15901,N_9111,N_11778);
or U15902 (N_15902,N_10723,N_8733);
nand U15903 (N_15903,N_11532,N_9419);
nand U15904 (N_15904,N_11248,N_8547);
and U15905 (N_15905,N_9465,N_10099);
and U15906 (N_15906,N_8138,N_8552);
xnor U15907 (N_15907,N_8811,N_10771);
nor U15908 (N_15908,N_9691,N_10996);
or U15909 (N_15909,N_9552,N_11439);
nor U15910 (N_15910,N_10527,N_11091);
xnor U15911 (N_15911,N_10188,N_9635);
nand U15912 (N_15912,N_10620,N_11565);
and U15913 (N_15913,N_8121,N_9906);
nand U15914 (N_15914,N_10182,N_9761);
nor U15915 (N_15915,N_8887,N_8613);
and U15916 (N_15916,N_10935,N_9380);
xor U15917 (N_15917,N_11917,N_9743);
nor U15918 (N_15918,N_9368,N_8361);
and U15919 (N_15919,N_11760,N_9791);
xnor U15920 (N_15920,N_10105,N_11320);
and U15921 (N_15921,N_9065,N_8937);
and U15922 (N_15922,N_11560,N_10578);
nor U15923 (N_15923,N_9346,N_8881);
xor U15924 (N_15924,N_10571,N_9475);
or U15925 (N_15925,N_10584,N_9874);
or U15926 (N_15926,N_9534,N_11100);
and U15927 (N_15927,N_9942,N_8850);
or U15928 (N_15928,N_10772,N_9539);
or U15929 (N_15929,N_11994,N_11478);
xor U15930 (N_15930,N_9823,N_10284);
and U15931 (N_15931,N_10393,N_9205);
and U15932 (N_15932,N_8505,N_9737);
nor U15933 (N_15933,N_8791,N_11547);
and U15934 (N_15934,N_11310,N_11502);
nor U15935 (N_15935,N_10828,N_11331);
nor U15936 (N_15936,N_10115,N_11774);
nand U15937 (N_15937,N_10309,N_8367);
and U15938 (N_15938,N_11717,N_11877);
or U15939 (N_15939,N_11296,N_11385);
xnor U15940 (N_15940,N_10791,N_8884);
and U15941 (N_15941,N_11103,N_8497);
or U15942 (N_15942,N_10307,N_8102);
nand U15943 (N_15943,N_11936,N_11707);
nor U15944 (N_15944,N_10765,N_8941);
and U15945 (N_15945,N_10549,N_8415);
nor U15946 (N_15946,N_11567,N_11150);
xnor U15947 (N_15947,N_9283,N_8667);
or U15948 (N_15948,N_10085,N_10967);
xor U15949 (N_15949,N_11467,N_10509);
nor U15950 (N_15950,N_11753,N_10461);
nor U15951 (N_15951,N_8801,N_11176);
nand U15952 (N_15952,N_8327,N_9824);
nand U15953 (N_15953,N_9741,N_10535);
nand U15954 (N_15954,N_10726,N_9895);
or U15955 (N_15955,N_9574,N_8019);
xnor U15956 (N_15956,N_10617,N_10684);
and U15957 (N_15957,N_9330,N_10731);
or U15958 (N_15958,N_10630,N_10132);
nand U15959 (N_15959,N_10226,N_10866);
and U15960 (N_15960,N_10480,N_11054);
nor U15961 (N_15961,N_8355,N_11680);
and U15962 (N_15962,N_10111,N_11615);
nand U15963 (N_15963,N_9777,N_9417);
nand U15964 (N_15964,N_9531,N_10961);
and U15965 (N_15965,N_8521,N_10568);
xnor U15966 (N_15966,N_8296,N_9561);
and U15967 (N_15967,N_9607,N_11401);
nor U15968 (N_15968,N_10024,N_11604);
and U15969 (N_15969,N_11742,N_9377);
nand U15970 (N_15970,N_9224,N_9476);
xnor U15971 (N_15971,N_11618,N_9181);
and U15972 (N_15972,N_9525,N_9883);
xnor U15973 (N_15973,N_9722,N_10326);
or U15974 (N_15974,N_9335,N_9308);
xor U15975 (N_15975,N_8408,N_10740);
nor U15976 (N_15976,N_9071,N_11802);
nor U15977 (N_15977,N_10906,N_9822);
nand U15978 (N_15978,N_10800,N_9478);
or U15979 (N_15979,N_11733,N_8710);
and U15980 (N_15980,N_9855,N_10602);
nor U15981 (N_15981,N_10155,N_11911);
nor U15982 (N_15982,N_10900,N_10800);
nand U15983 (N_15983,N_11302,N_11984);
nand U15984 (N_15984,N_9815,N_9964);
or U15985 (N_15985,N_11231,N_11940);
or U15986 (N_15986,N_10709,N_9758);
and U15987 (N_15987,N_9228,N_9519);
nor U15988 (N_15988,N_8495,N_9438);
xnor U15989 (N_15989,N_8243,N_11783);
or U15990 (N_15990,N_8966,N_10281);
nand U15991 (N_15991,N_10863,N_8470);
xnor U15992 (N_15992,N_9852,N_10585);
nand U15993 (N_15993,N_11516,N_8467);
xor U15994 (N_15994,N_9437,N_10142);
xnor U15995 (N_15995,N_8830,N_9666);
xnor U15996 (N_15996,N_11446,N_11236);
nand U15997 (N_15997,N_10039,N_9341);
xor U15998 (N_15998,N_8360,N_9245);
xor U15999 (N_15999,N_10318,N_11171);
nand U16000 (N_16000,N_13892,N_13412);
and U16001 (N_16001,N_13978,N_15581);
or U16002 (N_16002,N_12904,N_13973);
and U16003 (N_16003,N_15989,N_12741);
and U16004 (N_16004,N_15206,N_14983);
nand U16005 (N_16005,N_14300,N_12479);
and U16006 (N_16006,N_15618,N_15228);
xnor U16007 (N_16007,N_12139,N_13212);
nand U16008 (N_16008,N_13602,N_12433);
xor U16009 (N_16009,N_13127,N_14391);
and U16010 (N_16010,N_12974,N_13494);
xor U16011 (N_16011,N_12030,N_13251);
nor U16012 (N_16012,N_14161,N_14304);
and U16013 (N_16013,N_13264,N_13630);
and U16014 (N_16014,N_13129,N_13324);
and U16015 (N_16015,N_14911,N_15844);
or U16016 (N_16016,N_12287,N_12873);
or U16017 (N_16017,N_13195,N_13760);
xor U16018 (N_16018,N_14477,N_12487);
or U16019 (N_16019,N_15922,N_13046);
and U16020 (N_16020,N_13047,N_12919);
or U16021 (N_16021,N_13719,N_12359);
and U16022 (N_16022,N_12209,N_14722);
nor U16023 (N_16023,N_12100,N_15147);
and U16024 (N_16024,N_13285,N_13036);
and U16025 (N_16025,N_14111,N_13987);
or U16026 (N_16026,N_14714,N_15873);
and U16027 (N_16027,N_12448,N_13140);
and U16028 (N_16028,N_12543,N_14982);
and U16029 (N_16029,N_12705,N_13540);
and U16030 (N_16030,N_12156,N_15127);
nor U16031 (N_16031,N_15010,N_14448);
or U16032 (N_16032,N_14016,N_15680);
or U16033 (N_16033,N_14057,N_13778);
and U16034 (N_16034,N_14277,N_14054);
or U16035 (N_16035,N_13015,N_15476);
nand U16036 (N_16036,N_15636,N_15863);
xor U16037 (N_16037,N_15980,N_13990);
and U16038 (N_16038,N_14893,N_15626);
and U16039 (N_16039,N_14798,N_14709);
nand U16040 (N_16040,N_13135,N_12596);
nand U16041 (N_16041,N_13656,N_13795);
nand U16042 (N_16042,N_13367,N_12679);
or U16043 (N_16043,N_15717,N_13054);
xnor U16044 (N_16044,N_15439,N_14322);
nand U16045 (N_16045,N_12285,N_14419);
nor U16046 (N_16046,N_15809,N_15464);
nor U16047 (N_16047,N_13049,N_12591);
or U16048 (N_16048,N_15929,N_13300);
and U16049 (N_16049,N_12746,N_15481);
nor U16050 (N_16050,N_15978,N_12770);
and U16051 (N_16051,N_15702,N_15693);
and U16052 (N_16052,N_13826,N_15577);
or U16053 (N_16053,N_12653,N_15383);
nand U16054 (N_16054,N_14620,N_12057);
xnor U16055 (N_16055,N_13851,N_12384);
nand U16056 (N_16056,N_12029,N_15241);
nand U16057 (N_16057,N_13016,N_13694);
nand U16058 (N_16058,N_12109,N_13974);
xor U16059 (N_16059,N_12240,N_12731);
xnor U16060 (N_16060,N_15645,N_13548);
and U16061 (N_16061,N_12925,N_14287);
nor U16062 (N_16062,N_12480,N_13202);
nor U16063 (N_16063,N_13669,N_15780);
nand U16064 (N_16064,N_13542,N_14811);
nor U16065 (N_16065,N_12718,N_12300);
nor U16066 (N_16066,N_13703,N_15415);
xnor U16067 (N_16067,N_13901,N_12097);
nand U16068 (N_16068,N_15991,N_12739);
and U16069 (N_16069,N_14717,N_14857);
nor U16070 (N_16070,N_15759,N_15771);
nand U16071 (N_16071,N_14110,N_13501);
nor U16072 (N_16072,N_13402,N_14467);
nand U16073 (N_16073,N_13690,N_15106);
or U16074 (N_16074,N_12115,N_15994);
and U16075 (N_16075,N_14913,N_13903);
and U16076 (N_16076,N_14416,N_13783);
nand U16077 (N_16077,N_15749,N_14774);
and U16078 (N_16078,N_13295,N_14818);
or U16079 (N_16079,N_14910,N_12588);
or U16080 (N_16080,N_15200,N_13192);
or U16081 (N_16081,N_13033,N_13169);
nor U16082 (N_16082,N_14083,N_13014);
or U16083 (N_16083,N_13335,N_14260);
nor U16084 (N_16084,N_14430,N_14427);
and U16085 (N_16085,N_15006,N_12875);
nor U16086 (N_16086,N_15907,N_14155);
nor U16087 (N_16087,N_12491,N_13699);
nor U16088 (N_16088,N_14286,N_14056);
xor U16089 (N_16089,N_15800,N_14623);
and U16090 (N_16090,N_13452,N_15840);
nand U16091 (N_16091,N_15421,N_14943);
nand U16092 (N_16092,N_12738,N_14332);
nand U16093 (N_16093,N_13546,N_12874);
or U16094 (N_16094,N_14696,N_12523);
nand U16095 (N_16095,N_15865,N_13789);
nor U16096 (N_16096,N_14432,N_13902);
nor U16097 (N_16097,N_13331,N_15242);
and U16098 (N_16098,N_14653,N_15979);
xnor U16099 (N_16099,N_15627,N_15117);
or U16100 (N_16100,N_15632,N_14951);
and U16101 (N_16101,N_12188,N_14815);
nor U16102 (N_16102,N_14704,N_13578);
and U16103 (N_16103,N_14514,N_15948);
nor U16104 (N_16104,N_13361,N_15278);
nor U16105 (N_16105,N_13244,N_15917);
nor U16106 (N_16106,N_15246,N_13675);
and U16107 (N_16107,N_12430,N_14906);
xnor U16108 (N_16108,N_14861,N_15190);
or U16109 (N_16109,N_14359,N_13609);
or U16110 (N_16110,N_15082,N_12550);
nand U16111 (N_16111,N_15177,N_12867);
or U16112 (N_16112,N_15723,N_12171);
nand U16113 (N_16113,N_13814,N_14999);
nor U16114 (N_16114,N_12497,N_13327);
or U16115 (N_16115,N_14450,N_12467);
nor U16116 (N_16116,N_14148,N_14768);
nor U16117 (N_16117,N_14400,N_14005);
nand U16118 (N_16118,N_14226,N_13203);
nand U16119 (N_16119,N_13372,N_13286);
or U16120 (N_16120,N_14449,N_13437);
xnor U16121 (N_16121,N_12839,N_13302);
nand U16122 (N_16122,N_12977,N_15855);
nor U16123 (N_16123,N_12759,N_14070);
nor U16124 (N_16124,N_15522,N_14905);
or U16125 (N_16125,N_13223,N_13048);
xnor U16126 (N_16126,N_12053,N_12119);
nand U16127 (N_16127,N_12437,N_14593);
nand U16128 (N_16128,N_15870,N_15957);
nor U16129 (N_16129,N_15208,N_14429);
or U16130 (N_16130,N_15672,N_13796);
nand U16131 (N_16131,N_12236,N_14525);
nor U16132 (N_16132,N_13822,N_15341);
or U16133 (N_16133,N_15696,N_13947);
xnor U16134 (N_16134,N_13770,N_12423);
xnor U16135 (N_16135,N_12899,N_14694);
nor U16136 (N_16136,N_13209,N_15361);
xor U16137 (N_16137,N_15395,N_13568);
and U16138 (N_16138,N_13252,N_12727);
xor U16139 (N_16139,N_15535,N_15732);
nor U16140 (N_16140,N_14371,N_15498);
and U16141 (N_16141,N_14784,N_12672);
and U16142 (N_16142,N_12647,N_15201);
and U16143 (N_16143,N_12734,N_12579);
nand U16144 (N_16144,N_15416,N_15451);
xnor U16145 (N_16145,N_15235,N_13842);
nand U16146 (N_16146,N_12829,N_13811);
nand U16147 (N_16147,N_13876,N_15417);
nand U16148 (N_16148,N_13599,N_15593);
nand U16149 (N_16149,N_14095,N_14840);
and U16150 (N_16150,N_12447,N_14828);
nand U16151 (N_16151,N_13788,N_14338);
nand U16152 (N_16152,N_15921,N_12312);
nor U16153 (N_16153,N_12354,N_12279);
nand U16154 (N_16154,N_14168,N_15324);
and U16155 (N_16155,N_12267,N_15370);
and U16156 (N_16156,N_12696,N_13891);
nor U16157 (N_16157,N_14045,N_14563);
nand U16158 (N_16158,N_13189,N_12199);
and U16159 (N_16159,N_15616,N_13344);
nor U16160 (N_16160,N_13512,N_15788);
nor U16161 (N_16161,N_14935,N_13627);
nand U16162 (N_16162,N_15144,N_14590);
nor U16163 (N_16163,N_14357,N_12931);
nor U16164 (N_16164,N_12706,N_12019);
nor U16165 (N_16165,N_14848,N_12182);
nand U16166 (N_16166,N_15765,N_15711);
nor U16167 (N_16167,N_14436,N_14843);
nand U16168 (N_16168,N_14132,N_15166);
nand U16169 (N_16169,N_15336,N_15047);
and U16170 (N_16170,N_12064,N_15996);
nor U16171 (N_16171,N_12783,N_15014);
xor U16172 (N_16172,N_14866,N_12861);
and U16173 (N_16173,N_14320,N_13066);
nand U16174 (N_16174,N_15032,N_13194);
nand U16175 (N_16175,N_12963,N_15815);
or U16176 (N_16176,N_12786,N_14059);
nand U16177 (N_16177,N_14502,N_12125);
and U16178 (N_16178,N_13874,N_13853);
nor U16179 (N_16179,N_14550,N_15783);
nand U16180 (N_16180,N_13387,N_15631);
and U16181 (N_16181,N_14124,N_15779);
and U16182 (N_16182,N_13311,N_13197);
nand U16183 (N_16183,N_15866,N_13174);
nand U16184 (N_16184,N_14692,N_15384);
xnor U16185 (N_16185,N_15879,N_12277);
and U16186 (N_16186,N_12206,N_12844);
and U16187 (N_16187,N_15443,N_14594);
or U16188 (N_16188,N_13716,N_12773);
or U16189 (N_16189,N_13185,N_15570);
or U16190 (N_16190,N_12996,N_15853);
and U16191 (N_16191,N_13371,N_13143);
nor U16192 (N_16192,N_15052,N_12490);
nor U16193 (N_16193,N_15191,N_13766);
or U16194 (N_16194,N_15269,N_15086);
or U16195 (N_16195,N_12344,N_12054);
or U16196 (N_16196,N_12386,N_13226);
or U16197 (N_16197,N_13918,N_15111);
nand U16198 (N_16198,N_13485,N_14298);
and U16199 (N_16199,N_14270,N_15952);
or U16200 (N_16200,N_14756,N_15161);
nand U16201 (N_16201,N_15130,N_14166);
or U16202 (N_16202,N_13722,N_14499);
or U16203 (N_16203,N_13895,N_13684);
xor U16204 (N_16204,N_15835,N_12035);
or U16205 (N_16205,N_15501,N_15735);
nor U16206 (N_16206,N_14962,N_14718);
and U16207 (N_16207,N_14081,N_14365);
xor U16208 (N_16208,N_14695,N_14702);
and U16209 (N_16209,N_14173,N_15679);
and U16210 (N_16210,N_14998,N_13279);
nor U16211 (N_16211,N_14330,N_12779);
nor U16212 (N_16212,N_13061,N_13291);
or U16213 (N_16213,N_12772,N_15905);
or U16214 (N_16214,N_15985,N_15475);
xnor U16215 (N_16215,N_14239,N_13827);
or U16216 (N_16216,N_13005,N_13089);
or U16217 (N_16217,N_14965,N_15318);
nor U16218 (N_16218,N_15126,N_15705);
nor U16219 (N_16219,N_14248,N_14625);
and U16220 (N_16220,N_13801,N_15364);
nand U16221 (N_16221,N_14823,N_15545);
nor U16222 (N_16222,N_13365,N_15251);
nor U16223 (N_16223,N_14790,N_13196);
xnor U16224 (N_16224,N_14602,N_15128);
nand U16225 (N_16225,N_12516,N_15002);
nand U16226 (N_16226,N_15926,N_12237);
nand U16227 (N_16227,N_13883,N_15592);
nand U16228 (N_16228,N_13071,N_14619);
nand U16229 (N_16229,N_15941,N_12548);
and U16230 (N_16230,N_15041,N_13262);
nor U16231 (N_16231,N_13498,N_12594);
and U16232 (N_16232,N_12618,N_13368);
and U16233 (N_16233,N_12699,N_13598);
xnor U16234 (N_16234,N_14308,N_12000);
or U16235 (N_16235,N_15659,N_13466);
or U16236 (N_16236,N_13607,N_13750);
xor U16237 (N_16237,N_12617,N_13704);
or U16238 (N_16238,N_13083,N_14881);
and U16239 (N_16239,N_12754,N_12113);
nand U16240 (N_16240,N_15834,N_12654);
or U16241 (N_16241,N_13771,N_13261);
nor U16242 (N_16242,N_12290,N_12173);
or U16243 (N_16243,N_14407,N_12584);
or U16244 (N_16244,N_14511,N_13507);
nor U16245 (N_16245,N_12634,N_13175);
xor U16246 (N_16246,N_14047,N_14180);
nor U16247 (N_16247,N_13081,N_14508);
and U16248 (N_16248,N_13097,N_15465);
xnor U16249 (N_16249,N_15213,N_14832);
or U16250 (N_16250,N_15359,N_12663);
or U16251 (N_16251,N_14367,N_15021);
and U16252 (N_16252,N_14312,N_14354);
and U16253 (N_16253,N_13687,N_15804);
nor U16254 (N_16254,N_15756,N_12367);
or U16255 (N_16255,N_15753,N_15268);
xnor U16256 (N_16256,N_15477,N_15848);
nand U16257 (N_16257,N_14479,N_15785);
or U16258 (N_16258,N_14442,N_14642);
nor U16259 (N_16259,N_13500,N_15141);
nor U16260 (N_16260,N_13405,N_12471);
nor U16261 (N_16261,N_12380,N_13531);
or U16262 (N_16262,N_14664,N_14437);
xor U16263 (N_16263,N_12078,N_15977);
and U16264 (N_16264,N_15039,N_14631);
or U16265 (N_16265,N_15293,N_13522);
and U16266 (N_16266,N_14720,N_13929);
nor U16267 (N_16267,N_14876,N_15775);
xor U16268 (N_16268,N_12278,N_15396);
nor U16269 (N_16269,N_15031,N_15463);
nor U16270 (N_16270,N_14188,N_12520);
nand U16271 (N_16271,N_13067,N_14099);
nor U16272 (N_16272,N_15916,N_15081);
and U16273 (N_16273,N_15874,N_15605);
and U16274 (N_16274,N_15868,N_13710);
xor U16275 (N_16275,N_15928,N_12259);
nor U16276 (N_16276,N_12216,N_14103);
nor U16277 (N_16277,N_14268,N_13931);
xnor U16278 (N_16278,N_12048,N_12638);
nor U16279 (N_16279,N_13142,N_12944);
or U16280 (N_16280,N_15966,N_15986);
nor U16281 (N_16281,N_15690,N_14898);
nand U16282 (N_16282,N_15656,N_12089);
nand U16283 (N_16283,N_13329,N_15113);
nor U16284 (N_16284,N_13044,N_13400);
and U16285 (N_16285,N_15387,N_12868);
nand U16286 (N_16286,N_15115,N_12703);
and U16287 (N_16287,N_12432,N_13856);
xnor U16288 (N_16288,N_12728,N_12508);
xnor U16289 (N_16289,N_15280,N_15940);
or U16290 (N_16290,N_14690,N_13167);
nand U16291 (N_16291,N_12052,N_14195);
nand U16292 (N_16292,N_13233,N_15319);
and U16293 (N_16293,N_12326,N_13063);
xnor U16294 (N_16294,N_13473,N_13744);
and U16295 (N_16295,N_13587,N_13552);
nand U16296 (N_16296,N_12789,N_12458);
and U16297 (N_16297,N_12541,N_12565);
or U16298 (N_16298,N_13949,N_12485);
and U16299 (N_16299,N_15492,N_12357);
nor U16300 (N_16300,N_13581,N_15369);
xor U16301 (N_16301,N_15248,N_15777);
nor U16302 (N_16302,N_15598,N_15900);
or U16303 (N_16303,N_13358,N_12655);
nor U16304 (N_16304,N_14093,N_15467);
xor U16305 (N_16305,N_12723,N_14739);
xor U16306 (N_16306,N_14725,N_13836);
xnor U16307 (N_16307,N_12559,N_13137);
xnor U16308 (N_16308,N_15628,N_14633);
or U16309 (N_16309,N_12832,N_14376);
nor U16310 (N_16310,N_15335,N_15438);
xnor U16311 (N_16311,N_14894,N_12145);
and U16312 (N_16312,N_15181,N_15488);
nand U16313 (N_16313,N_12489,N_15472);
nand U16314 (N_16314,N_12481,N_13734);
xnor U16315 (N_16315,N_14968,N_12842);
nor U16316 (N_16316,N_13276,N_12794);
xor U16317 (N_16317,N_12225,N_12218);
and U16318 (N_16318,N_13147,N_14397);
or U16319 (N_16319,N_12046,N_15580);
xor U16320 (N_16320,N_15017,N_13832);
nand U16321 (N_16321,N_13274,N_12602);
nor U16322 (N_16322,N_14141,N_12219);
or U16323 (N_16323,N_12972,N_15043);
xor U16324 (N_16324,N_14708,N_15386);
nor U16325 (N_16325,N_12722,N_14364);
and U16326 (N_16326,N_14204,N_14241);
nand U16327 (N_16327,N_14115,N_13667);
xnor U16328 (N_16328,N_14137,N_12247);
or U16329 (N_16329,N_14765,N_15778);
nand U16330 (N_16330,N_14542,N_15352);
nand U16331 (N_16331,N_13004,N_12691);
nand U16332 (N_16332,N_12304,N_15424);
xnor U16333 (N_16333,N_15608,N_14870);
nand U16334 (N_16334,N_13356,N_14939);
or U16335 (N_16335,N_14895,N_12778);
xor U16336 (N_16336,N_15595,N_12614);
nor U16337 (N_16337,N_15094,N_14516);
xnor U16338 (N_16338,N_12201,N_14107);
and U16339 (N_16339,N_15821,N_12499);
nor U16340 (N_16340,N_13439,N_13039);
nor U16341 (N_16341,N_13438,N_13395);
and U16342 (N_16342,N_12358,N_14920);
nand U16343 (N_16343,N_12866,N_13451);
nor U16344 (N_16344,N_12733,N_15088);
nor U16345 (N_16345,N_12311,N_15289);
nor U16346 (N_16346,N_15934,N_14738);
and U16347 (N_16347,N_14150,N_14776);
nor U16348 (N_16348,N_13511,N_15644);
xnor U16349 (N_16349,N_13413,N_15216);
nor U16350 (N_16350,N_15569,N_15737);
or U16351 (N_16351,N_13723,N_15987);
xnor U16352 (N_16352,N_12093,N_14865);
and U16353 (N_16353,N_12616,N_12760);
xor U16354 (N_16354,N_13379,N_12217);
xor U16355 (N_16355,N_15054,N_12853);
xnor U16356 (N_16356,N_14553,N_15262);
nand U16357 (N_16357,N_14766,N_14956);
and U16358 (N_16358,N_14335,N_13079);
nor U16359 (N_16359,N_12212,N_12845);
xor U16360 (N_16360,N_13236,N_13769);
or U16361 (N_16361,N_12066,N_14571);
or U16362 (N_16362,N_15053,N_13878);
or U16363 (N_16363,N_13339,N_14628);
or U16364 (N_16364,N_12645,N_12750);
nand U16365 (N_16365,N_15090,N_13380);
nand U16366 (N_16366,N_12270,N_15549);
nor U16367 (N_16367,N_15413,N_14804);
or U16368 (N_16368,N_14845,N_14849);
and U16369 (N_16369,N_15551,N_15282);
nor U16370 (N_16370,N_15349,N_14710);
nand U16371 (N_16371,N_12851,N_12393);
nand U16372 (N_16372,N_12708,N_12105);
xor U16373 (N_16373,N_13184,N_15093);
nand U16374 (N_16374,N_15305,N_14698);
or U16375 (N_16375,N_14246,N_12637);
and U16376 (N_16376,N_15585,N_12933);
nor U16377 (N_16377,N_13270,N_15588);
or U16378 (N_16378,N_13425,N_13007);
nand U16379 (N_16379,N_14624,N_15281);
nand U16380 (N_16380,N_14085,N_15642);
or U16381 (N_16381,N_15427,N_15483);
nor U16382 (N_16382,N_15441,N_13806);
nand U16383 (N_16383,N_13082,N_13867);
and U16384 (N_16384,N_12396,N_14880);
nand U16385 (N_16385,N_14570,N_12776);
or U16386 (N_16386,N_15565,N_15139);
or U16387 (N_16387,N_12365,N_13945);
and U16388 (N_16388,N_15303,N_15886);
nor U16389 (N_16389,N_14887,N_14039);
nand U16390 (N_16390,N_12379,N_14475);
nand U16391 (N_16391,N_14329,N_12863);
nand U16392 (N_16392,N_12020,N_12101);
and U16393 (N_16393,N_12902,N_14334);
nand U16394 (N_16394,N_13877,N_12039);
nor U16395 (N_16395,N_15403,N_14482);
nor U16396 (N_16396,N_12387,N_14979);
xnor U16397 (N_16397,N_12184,N_15652);
and U16398 (N_16398,N_14201,N_14807);
nor U16399 (N_16399,N_14460,N_14163);
or U16400 (N_16400,N_13421,N_12788);
nand U16401 (N_16401,N_12268,N_13539);
nor U16402 (N_16402,N_15160,N_12854);
or U16403 (N_16403,N_15715,N_13388);
nor U16404 (N_16404,N_14337,N_14066);
or U16405 (N_16405,N_15851,N_13064);
nor U16406 (N_16406,N_12678,N_15689);
nor U16407 (N_16407,N_13177,N_12427);
and U16408 (N_16408,N_13809,N_14087);
and U16409 (N_16409,N_14262,N_14902);
nand U16410 (N_16410,N_13316,N_12394);
xnor U16411 (N_16411,N_15007,N_14133);
or U16412 (N_16412,N_14000,N_12767);
nor U16413 (N_16413,N_15204,N_13784);
xor U16414 (N_16414,N_15400,N_12887);
nor U16415 (N_16415,N_12266,N_12568);
or U16416 (N_16416,N_12841,N_13923);
and U16417 (N_16417,N_12351,N_12674);
nor U16418 (N_16418,N_13622,N_15751);
nand U16419 (N_16419,N_13012,N_15018);
or U16420 (N_16420,N_15003,N_13056);
or U16421 (N_16421,N_15784,N_13596);
and U16422 (N_16422,N_14543,N_13724);
xnor U16423 (N_16423,N_12383,N_12466);
nand U16424 (N_16424,N_14612,N_12038);
nor U16425 (N_16425,N_14038,N_14750);
xnor U16426 (N_16426,N_13072,N_13366);
and U16427 (N_16427,N_15012,N_13757);
or U16428 (N_16428,N_12456,N_15304);
nor U16429 (N_16429,N_14547,N_13392);
nor U16430 (N_16430,N_13435,N_15739);
or U16431 (N_16431,N_13935,N_12987);
or U16432 (N_16432,N_14381,N_12272);
or U16433 (N_16433,N_14167,N_14523);
nor U16434 (N_16434,N_14517,N_14379);
or U16435 (N_16435,N_15096,N_12400);
and U16436 (N_16436,N_13686,N_13616);
nor U16437 (N_16437,N_15231,N_13653);
or U16438 (N_16438,N_13761,N_13764);
xnor U16439 (N_16439,N_12451,N_12833);
nand U16440 (N_16440,N_14575,N_13090);
or U16441 (N_16441,N_13709,N_13678);
and U16442 (N_16442,N_15954,N_13409);
xor U16443 (N_16443,N_13659,N_12293);
xor U16444 (N_16444,N_12228,N_15606);
xor U16445 (N_16445,N_12009,N_15153);
xnor U16446 (N_16446,N_14417,N_13266);
nand U16447 (N_16447,N_13965,N_12459);
xnor U16448 (N_16448,N_13643,N_14215);
nor U16449 (N_16449,N_12059,N_15512);
xnor U16450 (N_16450,N_12322,N_15230);
and U16451 (N_16451,N_12342,N_14558);
or U16452 (N_16452,N_14938,N_12371);
nand U16453 (N_16453,N_14190,N_15964);
or U16454 (N_16454,N_13674,N_12802);
nand U16455 (N_16455,N_14797,N_14799);
xnor U16456 (N_16456,N_13818,N_14626);
nor U16457 (N_16457,N_14996,N_13172);
and U16458 (N_16458,N_13559,N_15867);
or U16459 (N_16459,N_13620,N_15050);
and U16460 (N_16460,N_14859,N_13858);
xor U16461 (N_16461,N_14264,N_14787);
nand U16462 (N_16462,N_12527,N_14258);
and U16463 (N_16463,N_12421,N_12622);
nand U16464 (N_16464,N_13812,N_13182);
xor U16465 (N_16465,N_12503,N_13865);
or U16466 (N_16466,N_12368,N_15660);
xnor U16467 (N_16467,N_14443,N_15025);
xnor U16468 (N_16468,N_12855,N_12177);
or U16469 (N_16469,N_15892,N_15220);
nand U16470 (N_16470,N_12547,N_13134);
or U16471 (N_16471,N_13314,N_15380);
nor U16472 (N_16472,N_15773,N_13087);
nor U16473 (N_16473,N_12744,N_13807);
and U16474 (N_16474,N_14489,N_12238);
nor U16475 (N_16475,N_13802,N_15677);
nor U16476 (N_16476,N_14847,N_13427);
nor U16477 (N_16477,N_14842,N_12425);
xnor U16478 (N_16478,N_12318,N_14306);
nand U16479 (N_16479,N_12167,N_12824);
or U16480 (N_16480,N_15621,N_13162);
xor U16481 (N_16481,N_14869,N_14521);
and U16482 (N_16482,N_14515,N_13513);
xnor U16483 (N_16483,N_15292,N_15573);
nor U16484 (N_16484,N_15760,N_12542);
nand U16485 (N_16485,N_13608,N_13991);
nand U16486 (N_16486,N_15724,N_14961);
nor U16487 (N_16487,N_13852,N_15534);
nand U16488 (N_16488,N_15033,N_12410);
and U16489 (N_16489,N_12418,N_15706);
nor U16490 (N_16490,N_13484,N_12047);
or U16491 (N_16491,N_15752,N_13957);
nand U16492 (N_16492,N_12980,N_12338);
xor U16493 (N_16493,N_15210,N_13996);
xor U16494 (N_16494,N_13328,N_13943);
and U16495 (N_16495,N_14730,N_13100);
nor U16496 (N_16496,N_14089,N_13478);
nand U16497 (N_16497,N_15509,N_14757);
xor U16498 (N_16498,N_14522,N_14356);
and U16499 (N_16499,N_13355,N_15264);
nand U16500 (N_16500,N_13577,N_14323);
xnor U16501 (N_16501,N_12816,N_15158);
nor U16502 (N_16502,N_12281,N_13873);
nor U16503 (N_16503,N_15331,N_14297);
and U16504 (N_16504,N_14679,N_12872);
xor U16505 (N_16505,N_12325,N_12564);
and U16506 (N_16506,N_12040,N_14023);
nand U16507 (N_16507,N_12398,N_13964);
or U16508 (N_16508,N_14232,N_12292);
xor U16509 (N_16509,N_12667,N_14552);
nand U16510 (N_16510,N_14129,N_14014);
nand U16511 (N_16511,N_13346,N_14254);
nand U16512 (N_16512,N_15687,N_15741);
xnor U16513 (N_16513,N_15638,N_12592);
nand U16514 (N_16514,N_14819,N_13492);
nand U16515 (N_16515,N_13497,N_13325);
nor U16516 (N_16516,N_15532,N_12011);
or U16517 (N_16517,N_12659,N_13280);
and U16518 (N_16518,N_13429,N_13547);
or U16519 (N_16519,N_13523,N_13995);
and U16520 (N_16520,N_13493,N_14104);
nor U16521 (N_16521,N_15254,N_15899);
xor U16522 (N_16522,N_14969,N_13296);
or U16523 (N_16523,N_13749,N_12938);
nor U16524 (N_16524,N_13305,N_13352);
and U16525 (N_16525,N_13899,N_14358);
xor U16526 (N_16526,N_15301,N_15373);
xnor U16527 (N_16527,N_14636,N_15939);
or U16528 (N_16528,N_14537,N_15490);
xnor U16529 (N_16529,N_14324,N_13538);
xor U16530 (N_16530,N_12812,N_12693);
or U16531 (N_16531,N_12628,N_14891);
nand U16532 (N_16532,N_12544,N_14069);
xnor U16533 (N_16533,N_14135,N_15176);
and U16534 (N_16534,N_14705,N_12658);
nor U16535 (N_16535,N_12086,N_14856);
or U16536 (N_16536,N_12226,N_15883);
or U16537 (N_16537,N_12506,N_15221);
xnor U16538 (N_16538,N_13623,N_13272);
xor U16539 (N_16539,N_15502,N_15707);
or U16540 (N_16540,N_14128,N_15020);
and U16541 (N_16541,N_12352,N_14290);
xor U16542 (N_16542,N_13715,N_14614);
nand U16543 (N_16543,N_12023,N_14778);
xnor U16544 (N_16544,N_14406,N_13582);
nand U16545 (N_16545,N_14295,N_14924);
nor U16546 (N_16546,N_15321,N_15131);
nor U16547 (N_16547,N_15708,N_12941);
nand U16548 (N_16548,N_12108,N_15882);
xor U16549 (N_16549,N_12401,N_12174);
nor U16550 (N_16550,N_13489,N_14726);
xnor U16551 (N_16551,N_13461,N_14317);
or U16552 (N_16552,N_14368,N_15666);
nand U16553 (N_16553,N_13234,N_12598);
nand U16554 (N_16554,N_15197,N_12439);
xor U16555 (N_16555,N_15182,N_14812);
nor U16556 (N_16556,N_12979,N_15768);
nand U16557 (N_16557,N_15637,N_13791);
nand U16558 (N_16558,N_15445,N_13378);
and U16559 (N_16559,N_12959,N_14796);
nor U16560 (N_16560,N_15510,N_13820);
or U16561 (N_16561,N_13628,N_12211);
nand U16562 (N_16562,N_14402,N_13516);
and U16563 (N_16563,N_14027,N_12457);
nor U16564 (N_16564,N_12656,N_14122);
nand U16565 (N_16565,N_12422,N_13567);
and U16566 (N_16566,N_14583,N_14433);
nor U16567 (N_16567,N_15972,N_13971);
nand U16568 (N_16568,N_14918,N_15249);
and U16569 (N_16569,N_13790,N_15875);
nor U16570 (N_16570,N_13470,N_15664);
xor U16571 (N_16571,N_15613,N_13979);
nand U16572 (N_16572,N_14510,N_14572);
nand U16573 (N_16573,N_13341,N_15946);
nor U16574 (N_16574,N_13537,N_14316);
nand U16575 (N_16575,N_13364,N_12253);
or U16576 (N_16576,N_15789,N_15813);
and U16577 (N_16577,N_15663,N_13527);
nand U16578 (N_16578,N_14404,N_15346);
and U16579 (N_16579,N_13564,N_13794);
and U16580 (N_16580,N_15794,N_13403);
or U16581 (N_16581,N_15802,N_13925);
nor U16582 (N_16582,N_14294,N_15188);
nand U16583 (N_16583,N_15146,N_15185);
xnor U16584 (N_16584,N_14672,N_14278);
xor U16585 (N_16585,N_12126,N_14874);
and U16586 (N_16586,N_12298,N_15881);
or U16587 (N_16587,N_15850,N_14841);
or U16588 (N_16588,N_15808,N_14466);
nand U16589 (N_16589,N_15904,N_14839);
nor U16590 (N_16590,N_15528,N_15700);
or U16591 (N_16591,N_13154,N_15317);
nor U16592 (N_16592,N_13377,N_12954);
xor U16593 (N_16593,N_12835,N_12730);
nor U16594 (N_16594,N_12942,N_12557);
or U16595 (N_16595,N_12286,N_13938);
and U16596 (N_16596,N_12150,N_15920);
or U16597 (N_16597,N_12356,N_12103);
nand U16598 (N_16598,N_15484,N_13588);
xor U16599 (N_16599,N_15812,N_14131);
xnor U16600 (N_16600,N_14086,N_13849);
nand U16601 (N_16601,N_13752,N_14529);
or U16602 (N_16602,N_14393,N_13644);
and U16603 (N_16603,N_12571,N_12514);
and U16604 (N_16604,N_12815,N_15360);
xor U16605 (N_16605,N_13731,N_14719);
nor U16606 (N_16606,N_15065,N_12751);
or U16607 (N_16607,N_15822,N_12897);
xnor U16608 (N_16608,N_13505,N_15668);
or U16609 (N_16609,N_15470,N_12558);
nand U16610 (N_16610,N_13301,N_14011);
or U16611 (N_16611,N_13898,N_12695);
or U16612 (N_16612,N_14753,N_14897);
nor U16613 (N_16613,N_12347,N_14535);
xnor U16614 (N_16614,N_13835,N_13159);
nand U16615 (N_16615,N_13733,N_14703);
and U16616 (N_16616,N_15399,N_13128);
xnor U16617 (N_16617,N_14030,N_15138);
or U16618 (N_16618,N_13792,N_15530);
xnor U16619 (N_16619,N_14779,N_13845);
or U16620 (N_16620,N_15071,N_13188);
and U16621 (N_16621,N_12993,N_15738);
nand U16622 (N_16622,N_13070,N_15698);
and U16623 (N_16623,N_15733,N_15038);
and U16624 (N_16624,N_15048,N_12197);
and U16625 (N_16625,N_13886,N_15995);
and U16626 (N_16626,N_14281,N_12792);
or U16627 (N_16627,N_12151,N_15935);
nor U16628 (N_16628,N_14661,N_14862);
nand U16629 (N_16629,N_15155,N_13798);
nand U16630 (N_16630,N_12920,N_12283);
and U16631 (N_16631,N_13976,N_14805);
or U16632 (N_16632,N_13781,N_12194);
or U16633 (N_16633,N_13510,N_15365);
nor U16634 (N_16634,N_14227,N_12413);
xnor U16635 (N_16635,N_12136,N_12204);
nand U16636 (N_16636,N_12079,N_12399);
or U16637 (N_16637,N_12147,N_15423);
and U16638 (N_16638,N_14068,N_15970);
nor U16639 (N_16639,N_15328,N_14036);
nor U16640 (N_16640,N_14453,N_13170);
nand U16641 (N_16641,N_14347,N_13631);
and U16642 (N_16642,N_14205,N_14603);
and U16643 (N_16643,N_14527,N_15817);
nand U16644 (N_16644,N_12196,N_12683);
nand U16645 (N_16645,N_13774,N_12580);
nand U16646 (N_16646,N_14196,N_13846);
and U16647 (N_16647,N_13848,N_12526);
nand U16648 (N_16648,N_12880,N_14649);
and U16649 (N_16649,N_12373,N_13728);
xnor U16650 (N_16650,N_13386,N_13428);
or U16651 (N_16651,N_13269,N_14651);
nor U16652 (N_16652,N_15478,N_13805);
nand U16653 (N_16653,N_15993,N_12951);
nor U16654 (N_16654,N_12364,N_12595);
xnor U16655 (N_16655,N_15345,N_15397);
nand U16656 (N_16656,N_15552,N_13907);
or U16657 (N_16657,N_15168,N_12404);
xor U16658 (N_16658,N_12743,N_15793);
and U16659 (N_16659,N_12551,N_13859);
and U16660 (N_16660,N_12822,N_12484);
or U16661 (N_16661,N_12777,N_14864);
nor U16662 (N_16662,N_15447,N_14276);
nand U16663 (N_16663,N_12138,N_13362);
and U16664 (N_16664,N_12492,N_15938);
or U16665 (N_16665,N_13855,N_15960);
nand U16666 (N_16666,N_13453,N_12210);
nor U16667 (N_16667,N_13080,N_12026);
and U16668 (N_16668,N_12071,N_15260);
xor U16669 (N_16669,N_13893,N_12575);
nor U16670 (N_16670,N_12215,N_15625);
and U16671 (N_16671,N_14009,N_12791);
nand U16672 (N_16672,N_13661,N_13890);
nand U16673 (N_16673,N_13590,N_15713);
nand U16674 (N_16674,N_12134,N_15311);
xor U16675 (N_16675,N_12205,N_12798);
nand U16676 (N_16676,N_15604,N_14414);
or U16677 (N_16677,N_13755,N_12476);
or U16678 (N_16678,N_12895,N_15045);
xnor U16679 (N_16679,N_13913,N_12856);
nor U16680 (N_16680,N_14917,N_12032);
and U16681 (N_16681,N_13051,N_15747);
xor U16682 (N_16682,N_13166,N_15763);
or U16683 (N_16683,N_15243,N_12044);
nand U16684 (N_16684,N_15471,N_15600);
nor U16685 (N_16685,N_13157,N_14549);
or U16686 (N_16686,N_15872,N_12629);
nor U16687 (N_16687,N_13889,N_14462);
nor U16688 (N_16688,N_15901,N_13227);
and U16689 (N_16689,N_14064,N_14809);
and U16690 (N_16690,N_13062,N_15375);
or U16691 (N_16691,N_15211,N_14370);
xnor U16692 (N_16692,N_12806,N_14032);
nor U16693 (N_16693,N_14712,N_15283);
and U16694 (N_16694,N_12376,N_13514);
xor U16695 (N_16695,N_14885,N_13921);
nand U16696 (N_16696,N_15044,N_12091);
xnor U16697 (N_16697,N_12390,N_15036);
xnor U16698 (N_16698,N_15910,N_14284);
or U16699 (N_16699,N_15506,N_15564);
nor U16700 (N_16700,N_13714,N_12797);
nor U16701 (N_16701,N_14017,N_15560);
nor U16702 (N_16702,N_12611,N_12893);
nor U16703 (N_16703,N_15354,N_12860);
xnor U16704 (N_16704,N_14114,N_14072);
xor U16705 (N_16705,N_14401,N_14084);
nor U16706 (N_16706,N_14767,N_15832);
nand U16707 (N_16707,N_14257,N_13747);
nand U16708 (N_16708,N_14091,N_12665);
and U16709 (N_16709,N_12603,N_13271);
nand U16710 (N_16710,N_12507,N_13417);
and U16711 (N_16711,N_15758,N_15358);
nor U16712 (N_16712,N_13078,N_13446);
nor U16713 (N_16713,N_14478,N_14782);
and U16714 (N_16714,N_14598,N_15640);
or U16715 (N_16715,N_13250,N_12886);
and U16716 (N_16716,N_15179,N_12116);
xor U16717 (N_16717,N_14212,N_14206);
and U16718 (N_16718,N_13896,N_14744);
nor U16719 (N_16719,N_13635,N_12913);
and U16720 (N_16720,N_14492,N_12929);
nor U16721 (N_16721,N_13091,N_14816);
xnor U16722 (N_16722,N_15037,N_12412);
and U16723 (N_16723,N_15754,N_12524);
or U16724 (N_16724,N_15284,N_13111);
and U16725 (N_16725,N_14544,N_15487);
or U16726 (N_16726,N_15630,N_13476);
and U16727 (N_16727,N_14425,N_12018);
and U16728 (N_16728,N_12518,N_14130);
and U16729 (N_16729,N_15275,N_14662);
or U16730 (N_16730,N_15034,N_15889);
nand U16731 (N_16731,N_14451,N_14610);
nor U16732 (N_16732,N_15572,N_15500);
xor U16733 (N_16733,N_15955,N_13915);
and U16734 (N_16734,N_14972,N_15902);
nand U16735 (N_16735,N_15271,N_12709);
nand U16736 (N_16736,N_14904,N_13117);
nand U16737 (N_16737,N_12717,N_12682);
or U16738 (N_16738,N_12581,N_14240);
nand U16739 (N_16739,N_13011,N_15553);
xnor U16740 (N_16740,N_15140,N_13946);
or U16741 (N_16741,N_12843,N_13215);
nand U16742 (N_16742,N_13023,N_13375);
nand U16743 (N_16743,N_15801,N_14493);
and U16744 (N_16744,N_15704,N_15610);
nor U16745 (N_16745,N_14854,N_15442);
nor U16746 (N_16746,N_12962,N_12424);
nand U16747 (N_16747,N_13281,N_12303);
nand U16748 (N_16748,N_14934,N_12553);
nand U16749 (N_16749,N_13010,N_14344);
or U16750 (N_16750,N_12666,N_12690);
nand U16751 (N_16751,N_12114,N_13544);
nor U16752 (N_16752,N_14786,N_15225);
nand U16753 (N_16753,N_13611,N_12130);
nand U16754 (N_16754,N_14082,N_15273);
nor U16755 (N_16755,N_14458,N_15350);
xnor U16756 (N_16756,N_12910,N_14675);
nor U16757 (N_16757,N_14225,N_13994);
nor U16758 (N_16758,N_14658,N_13445);
nand U16759 (N_16759,N_15857,N_12360);
nor U16760 (N_16760,N_14251,N_14146);
nor U16761 (N_16761,N_13430,N_14736);
nor U16762 (N_16762,N_13257,N_12881);
xnor U16763 (N_16763,N_15026,N_13394);
xnor U16764 (N_16764,N_12083,N_12939);
nor U16765 (N_16765,N_12271,N_12224);
and U16766 (N_16766,N_13637,N_13385);
nand U16767 (N_16767,N_13436,N_13006);
xor U16768 (N_16768,N_15909,N_12475);
or U16769 (N_16769,N_15673,N_14513);
and U16770 (N_16770,N_12180,N_15250);
nand U16771 (N_16771,N_13939,N_14387);
xor U16772 (N_16772,N_14568,N_12961);
nand U16773 (N_16773,N_13954,N_13992);
and U16774 (N_16774,N_13163,N_13433);
nand U16775 (N_16775,N_14228,N_13662);
and U16776 (N_16776,N_14836,N_12309);
nor U16777 (N_16777,N_13586,N_14042);
and U16778 (N_16778,N_13563,N_12936);
xor U16779 (N_16779,N_15270,N_12095);
nor U16780 (N_16780,N_13057,N_15918);
or U16781 (N_16781,N_13222,N_13763);
xor U16782 (N_16782,N_15924,N_15504);
or U16783 (N_16783,N_12260,N_15137);
nand U16784 (N_16784,N_15234,N_15187);
and U16785 (N_16785,N_14975,N_13746);
xnor U16786 (N_16786,N_13758,N_14389);
nor U16787 (N_16787,N_15123,N_14200);
or U16788 (N_16788,N_15523,N_14834);
and U16789 (N_16789,N_14118,N_15184);
nand U16790 (N_16790,N_15836,N_13571);
or U16791 (N_16791,N_13554,N_12901);
nand U16792 (N_16792,N_13246,N_12058);
or U16793 (N_16793,N_15214,N_15721);
xnor U16794 (N_16794,N_15229,N_13292);
nor U16795 (N_16795,N_13972,N_15792);
and U16796 (N_16796,N_12249,N_14077);
and U16797 (N_16797,N_12428,N_14914);
or U16798 (N_16798,N_12072,N_13580);
nand U16799 (N_16799,N_15156,N_12274);
and U16800 (N_16800,N_15374,N_15887);
nand U16801 (N_16801,N_12335,N_15514);
and U16802 (N_16802,N_15653,N_14108);
nand U16803 (N_16803,N_14109,N_14193);
xor U16804 (N_16804,N_13824,N_14113);
or U16805 (N_16805,N_13732,N_14182);
xnor U16806 (N_16806,N_14456,N_15662);
and U16807 (N_16807,N_13638,N_13073);
xor U16808 (N_16808,N_13969,N_15408);
nand U16809 (N_16809,N_14564,N_15103);
and U16810 (N_16810,N_15297,N_13265);
and U16811 (N_16811,N_12120,N_12799);
nor U16812 (N_16812,N_12813,N_15893);
nor U16813 (N_16813,N_15388,N_14706);
or U16814 (N_16814,N_14817,N_15412);
nor U16815 (N_16815,N_15122,N_15694);
nand U16816 (N_16816,N_12736,N_14665);
or U16817 (N_16817,N_13614,N_13636);
and U16818 (N_16818,N_12619,N_15503);
nor U16819 (N_16819,N_13343,N_13503);
nand U16820 (N_16820,N_12891,N_12336);
xor U16821 (N_16821,N_14746,N_12753);
and U16822 (N_16822,N_13399,N_13960);
nor U16823 (N_16823,N_14480,N_14343);
or U16824 (N_16824,N_13799,N_15999);
xnor U16825 (N_16825,N_14713,N_15527);
xnor U16826 (N_16826,N_13666,N_15776);
or U16827 (N_16827,N_13245,N_14900);
and U16828 (N_16828,N_15407,N_13190);
and U16829 (N_16829,N_14551,N_14507);
xor U16830 (N_16830,N_15997,N_12593);
xor U16831 (N_16831,N_14667,N_14923);
or U16832 (N_16832,N_15120,N_13019);
and U16833 (N_16833,N_14233,N_14759);
nor U16834 (N_16834,N_13742,N_14878);
and U16835 (N_16835,N_14073,N_12641);
xnor U16836 (N_16836,N_15004,N_13854);
or U16837 (N_16837,N_12857,N_12406);
or U16838 (N_16838,N_13718,N_14994);
or U16839 (N_16839,N_14780,N_13739);
xnor U16840 (N_16840,N_14403,N_15634);
xor U16841 (N_16841,N_14309,N_13634);
or U16842 (N_16842,N_14995,N_14597);
and U16843 (N_16843,N_13668,N_15193);
nor U16844 (N_16844,N_15846,N_14966);
xnor U16845 (N_16845,N_12016,N_13058);
and U16846 (N_16846,N_15355,N_13076);
or U16847 (N_16847,N_14820,N_12563);
nand U16848 (N_16848,N_14399,N_14946);
or U16849 (N_16849,N_13431,N_13359);
and U16850 (N_16850,N_15529,N_13107);
or U16851 (N_16851,N_13242,N_15519);
or U16852 (N_16852,N_12320,N_13829);
or U16853 (N_16853,N_13029,N_15607);
and U16854 (N_16854,N_15314,N_13278);
nor U16855 (N_16855,N_15272,N_15343);
nor U16856 (N_16856,N_13570,N_14519);
or U16857 (N_16857,N_13583,N_15805);
xnor U16858 (N_16858,N_14431,N_13060);
xor U16859 (N_16859,N_12721,N_15351);
nand U16860 (N_16860,N_14410,N_15149);
and U16861 (N_16861,N_14987,N_12443);
xor U16862 (N_16862,N_15718,N_15425);
nor U16863 (N_16863,N_15937,N_13229);
nor U16864 (N_16864,N_14420,N_14288);
or U16865 (N_16865,N_12468,N_13228);
xor U16866 (N_16866,N_12947,N_12530);
xnor U16867 (N_16867,N_14903,N_14463);
and U16868 (N_16868,N_13743,N_14566);
or U16869 (N_16869,N_13651,N_13145);
nor U16870 (N_16870,N_15307,N_15209);
nand U16871 (N_16871,N_13740,N_14648);
and U16872 (N_16872,N_14325,N_12149);
or U16873 (N_16873,N_12950,N_15516);
nor U16874 (N_16874,N_13390,N_15452);
or U16875 (N_16875,N_12685,N_13624);
or U16876 (N_16876,N_13138,N_14172);
and U16877 (N_16877,N_14055,N_15173);
or U16878 (N_16878,N_15692,N_13629);
xor U16879 (N_16879,N_12633,N_13495);
or U16880 (N_16880,N_13124,N_13282);
nor U16881 (N_16881,N_14724,N_12441);
xnor U16882 (N_16882,N_13933,N_14940);
xnor U16883 (N_16883,N_12155,N_14785);
nor U16884 (N_16884,N_12607,N_15688);
nor U16885 (N_16885,N_12627,N_13434);
or U16886 (N_16886,N_14349,N_12203);
and U16887 (N_16887,N_13863,N_13831);
or U16888 (N_16888,N_15791,N_15828);
or U16889 (N_16889,N_12088,N_15537);
nand U16890 (N_16890,N_12317,N_14673);
or U16891 (N_16891,N_15049,N_12165);
xor U16892 (N_16892,N_13074,N_15109);
xnor U16893 (N_16893,N_13026,N_15450);
and U16894 (N_16894,N_13308,N_12402);
nor U16895 (N_16895,N_15726,N_12561);
and U16896 (N_16896,N_14271,N_14532);
and U16897 (N_16897,N_12092,N_12405);
nand U16898 (N_16898,N_14319,N_15334);
nand U16899 (N_16899,N_12050,N_14557);
xor U16900 (N_16900,N_12027,N_15609);
nor U16901 (N_16901,N_12988,N_12898);
xnor U16902 (N_16902,N_15798,N_15183);
and U16903 (N_16903,N_14139,N_15686);
nand U16904 (N_16904,N_12965,N_15965);
xnor U16905 (N_16905,N_14076,N_12296);
nand U16906 (N_16906,N_12850,N_15233);
xnor U16907 (N_16907,N_15665,N_12482);
nand U16908 (N_16908,N_12397,N_15119);
and U16909 (N_16909,N_12900,N_12075);
and U16910 (N_16910,N_13160,N_12033);
xnor U16911 (N_16911,N_14959,N_12820);
xnor U16912 (N_16912,N_15854,N_12597);
or U16913 (N_16913,N_13633,N_13721);
and U16914 (N_16914,N_13998,N_13767);
xor U16915 (N_16915,N_14307,N_13934);
nand U16916 (N_16916,N_13037,N_12185);
xor U16917 (N_16917,N_14145,N_15381);
nor U16918 (N_16918,N_14100,N_14112);
or U16919 (N_16919,N_12771,N_12202);
nand U16920 (N_16920,N_13952,N_14210);
or U16921 (N_16921,N_15040,N_14120);
xnor U16922 (N_16922,N_13369,N_12631);
nor U16923 (N_16923,N_13472,N_15539);
nand U16924 (N_16924,N_12889,N_15015);
and U16925 (N_16925,N_14976,N_15494);
nand U16926 (N_16926,N_12990,N_14031);
nand U16927 (N_16927,N_15430,N_13823);
or U16928 (N_16928,N_12008,N_12932);
xor U16929 (N_16929,N_13027,N_15895);
nand U16930 (N_16930,N_15685,N_14731);
and U16931 (N_16931,N_12230,N_13834);
or U16932 (N_16932,N_14948,N_12133);
xor U16933 (N_16933,N_15571,N_14230);
or U16934 (N_16934,N_13319,N_12455);
and U16935 (N_16935,N_15459,N_14160);
nand U16936 (N_16936,N_12346,N_13370);
or U16937 (N_16937,N_12774,N_14871);
nor U16938 (N_16938,N_12623,N_12284);
and U16939 (N_16939,N_14929,N_12823);
xnor U16940 (N_16940,N_12719,N_13594);
xor U16941 (N_16941,N_13841,N_12308);
nand U16942 (N_16942,N_12460,N_15574);
xnor U16943 (N_16943,N_12112,N_15479);
nor U16944 (N_16944,N_12276,N_12223);
xnor U16945 (N_16945,N_15073,N_13688);
or U16946 (N_16946,N_12143,N_13210);
xor U16947 (N_16947,N_13115,N_15393);
nand U16948 (N_16948,N_14363,N_15971);
and U16949 (N_16949,N_14803,N_12452);
nand U16950 (N_16950,N_12612,N_13573);
or U16951 (N_16951,N_12021,N_12585);
or U16952 (N_16952,N_13297,N_12043);
xor U16953 (N_16953,N_14388,N_12549);
and U16954 (N_16954,N_12545,N_15622);
xor U16955 (N_16955,N_15112,N_12846);
and U16956 (N_16956,N_13020,N_12273);
nand U16957 (N_16957,N_13002,N_14985);
or U16958 (N_16958,N_13391,N_13942);
nor U16959 (N_16959,N_13793,N_15238);
xor U16960 (N_16960,N_12689,N_15178);
and U16961 (N_16961,N_13866,N_14584);
xnor U16962 (N_16962,N_12251,N_15072);
and U16963 (N_16963,N_15750,N_15658);
and U16964 (N_16964,N_14580,N_12198);
and U16965 (N_16965,N_13401,N_12735);
xnor U16966 (N_16966,N_13253,N_13962);
xnor U16967 (N_16967,N_14781,N_14465);
nand U16968 (N_16968,N_12970,N_14280);
or U16969 (N_16969,N_13471,N_14273);
xor U16970 (N_16970,N_12669,N_15051);
xor U16971 (N_16971,N_15681,N_12574);
nand U16972 (N_16972,N_12190,N_14181);
nor U16973 (N_16973,N_12673,N_12207);
and U16974 (N_16974,N_13574,N_15614);
nor U16975 (N_16975,N_13555,N_14423);
xnor U16976 (N_16976,N_13720,N_14252);
nand U16977 (N_16977,N_15330,N_14468);
xnor U16978 (N_16978,N_14656,N_15332);
or U16979 (N_16979,N_12022,N_14471);
nand U16980 (N_16980,N_14772,N_14872);
nand U16981 (N_16981,N_13287,N_12014);
or U16982 (N_16982,N_12076,N_15402);
and U16983 (N_16983,N_12042,N_12494);
and U16984 (N_16984,N_14503,N_15974);
xnor U16985 (N_16985,N_12282,N_15655);
xor U16986 (N_16986,N_14875,N_14063);
nor U16987 (N_16987,N_15030,N_15437);
nand U16988 (N_16988,N_15772,N_15497);
or U16989 (N_16989,N_13442,N_13830);
xor U16990 (N_16990,N_13817,N_12742);
xnor U16991 (N_16991,N_15742,N_13810);
and U16992 (N_16992,N_13652,N_15142);
nand U16993 (N_16993,N_14922,N_12609);
nand U16994 (N_16994,N_14411,N_14860);
xor U16995 (N_16995,N_15419,N_13529);
or U16996 (N_16996,N_13022,N_12922);
nand U16997 (N_16997,N_13406,N_13705);
xor U16998 (N_16998,N_15761,N_12831);
or U16999 (N_16999,N_15489,N_15267);
xor U17000 (N_17000,N_14770,N_15584);
nor U17001 (N_17001,N_12056,N_12915);
and U17002 (N_17002,N_15810,N_13914);
xnor U17003 (N_17003,N_14669,N_15898);
and U17004 (N_17004,N_12324,N_14822);
nor U17005 (N_17005,N_14025,N_13150);
nand U17006 (N_17006,N_12964,N_12704);
nor U17007 (N_17007,N_12532,N_14674);
and U17008 (N_17008,N_14394,N_13642);
xor U17009 (N_17009,N_15285,N_12017);
nor U17010 (N_17010,N_12807,N_14238);
and U17011 (N_17011,N_13565,N_12555);
or U17012 (N_17012,N_14518,N_13665);
or U17013 (N_17013,N_14208,N_14646);
nand U17014 (N_17014,N_12998,N_12012);
or U17015 (N_17015,N_13785,N_15748);
nor U17016 (N_17016,N_15063,N_14313);
nor U17017 (N_17017,N_14191,N_13221);
nor U17018 (N_17018,N_12698,N_12462);
or U17019 (N_17019,N_12955,N_12257);
or U17020 (N_17020,N_13121,N_12613);
and U17021 (N_17021,N_12510,N_15556);
or U17022 (N_17022,N_13601,N_12768);
and U17023 (N_17023,N_12141,N_15499);
xor U17024 (N_17024,N_14678,N_15968);
xnor U17025 (N_17025,N_15027,N_15258);
xor U17026 (N_17026,N_12426,N_14029);
nor U17027 (N_17027,N_13950,N_15124);
or U17028 (N_17028,N_12301,N_13645);
nor U17029 (N_17029,N_13126,N_13102);
nor U17030 (N_17030,N_13569,N_13475);
xor U17031 (N_17031,N_13551,N_14078);
or U17032 (N_17032,N_14576,N_13288);
xor U17033 (N_17033,N_12626,N_13828);
xnor U17034 (N_17034,N_13671,N_13119);
xnor U17035 (N_17035,N_13647,N_15061);
nand U17036 (N_17036,N_12836,N_12763);
nand U17037 (N_17037,N_15555,N_15394);
or U17038 (N_17038,N_12805,N_12362);
nand U17039 (N_17039,N_12810,N_15295);
nand U17040 (N_17040,N_13920,N_14647);
and U17041 (N_17041,N_15382,N_14067);
and U17042 (N_17042,N_14538,N_12162);
and U17043 (N_17043,N_14217,N_14012);
or U17044 (N_17044,N_13116,N_12355);
or U17045 (N_17045,N_14749,N_14097);
xnor U17046 (N_17046,N_13632,N_13606);
or U17047 (N_17047,N_14153,N_14775);
and U17048 (N_17048,N_15826,N_14285);
xnor U17049 (N_17049,N_13096,N_15222);
and U17050 (N_17050,N_13207,N_14992);
or U17051 (N_17051,N_13910,N_13254);
or U17052 (N_17052,N_12315,N_13268);
or U17053 (N_17053,N_14140,N_15725);
or U17054 (N_17054,N_14158,N_15757);
and U17055 (N_17055,N_14827,N_12294);
nor U17056 (N_17056,N_14255,N_12407);
and U17057 (N_17057,N_13055,N_15876);
nand U17058 (N_17058,N_14990,N_13200);
nor U17059 (N_17059,N_15135,N_13104);
and U17060 (N_17060,N_13084,N_12461);
or U17061 (N_17061,N_14981,N_15009);
and U17062 (N_17062,N_12818,N_13028);
nor U17063 (N_17063,N_14793,N_12337);
and U17064 (N_17064,N_13986,N_13585);
and U17065 (N_17065,N_12649,N_13488);
nor U17066 (N_17066,N_14219,N_14004);
or U17067 (N_17067,N_13449,N_15744);
or U17068 (N_17068,N_12469,N_13455);
nand U17069 (N_17069,N_13487,N_12981);
nor U17070 (N_17070,N_12680,N_14826);
nor U17071 (N_17071,N_15462,N_12107);
and U17072 (N_17072,N_12796,N_12363);
xor U17073 (N_17073,N_13499,N_15849);
xor U17074 (N_17074,N_12388,N_14652);
and U17075 (N_17075,N_12940,N_12166);
nor U17076 (N_17076,N_13457,N_12725);
or U17077 (N_17077,N_15945,N_15180);
xor U17078 (N_17078,N_14398,N_14101);
nand U17079 (N_17079,N_15022,N_13717);
or U17080 (N_17080,N_15517,N_15440);
or U17081 (N_17081,N_14142,N_12906);
nand U17082 (N_17082,N_13619,N_14622);
or U17083 (N_17083,N_14742,N_15617);
nand U17084 (N_17084,N_12176,N_14378);
nand U17085 (N_17085,N_12142,N_12821);
xnor U17086 (N_17086,N_14020,N_14050);
and U17087 (N_17087,N_13284,N_15099);
and U17088 (N_17088,N_15406,N_15132);
xor U17089 (N_17089,N_13727,N_12036);
nor U17090 (N_17090,N_15148,N_15431);
xor U17091 (N_17091,N_12382,N_14792);
xnor U17092 (N_17092,N_14758,N_14606);
nand U17093 (N_17093,N_14138,N_14684);
or U17094 (N_17094,N_13179,N_15678);
xnor U17095 (N_17095,N_15448,N_12560);
nand U17096 (N_17096,N_13350,N_12828);
nor U17097 (N_17097,N_12552,N_12605);
or U17098 (N_17098,N_13576,N_14040);
or U17099 (N_17099,N_12323,N_15078);
nor U17100 (N_17100,N_15227,N_14808);
xor U17101 (N_17101,N_15461,N_15134);
xnor U17102 (N_17102,N_12540,N_14169);
nor U17103 (N_17103,N_12005,N_15101);
or U17104 (N_17104,N_13293,N_14604);
and U17105 (N_17105,N_14088,N_15864);
nand U17106 (N_17106,N_13306,N_14560);
and U17107 (N_17107,N_15342,N_13847);
nand U17108 (N_17108,N_15683,N_13158);
and U17109 (N_17109,N_12849,N_14486);
nand U17110 (N_17110,N_13738,N_15338);
and U17111 (N_17111,N_13605,N_12375);
and U17112 (N_17112,N_15769,N_14528);
nand U17113 (N_17113,N_12131,N_14327);
xnor U17114 (N_17114,N_14850,N_14657);
xor U17115 (N_17115,N_14562,N_13882);
nand U17116 (N_17116,N_14412,N_13450);
nor U17117 (N_17117,N_14051,N_15000);
xor U17118 (N_17118,N_15943,N_15795);
or U17119 (N_17119,N_14611,N_13217);
xnor U17120 (N_17120,N_14755,N_15410);
nor U17121 (N_17121,N_14873,N_12871);
or U17122 (N_17122,N_13131,N_15586);
xor U17123 (N_17123,N_12256,N_14339);
nor U17124 (N_17124,N_13787,N_14015);
nor U17125 (N_17125,N_13482,N_15562);
xor U17126 (N_17126,N_15511,N_13384);
nand U17127 (N_17127,N_15367,N_12995);
and U17128 (N_17128,N_12158,N_12556);
nor U17129 (N_17129,N_12067,N_15962);
nand U17130 (N_17130,N_12525,N_13342);
xnor U17131 (N_17131,N_15896,N_13900);
nand U17132 (N_17132,N_13021,N_12604);
nand U17133 (N_17133,N_14984,N_15056);
xnor U17134 (N_17134,N_15207,N_15596);
nand U17135 (N_17135,N_13017,N_14007);
or U17136 (N_17136,N_15411,N_13989);
nand U17137 (N_17137,N_12244,N_12884);
nor U17138 (N_17138,N_14728,N_12096);
xnor U17139 (N_17139,N_15219,N_12414);
nand U17140 (N_17140,N_15261,N_14435);
or U17141 (N_17141,N_12890,N_13298);
xnor U17142 (N_17142,N_13204,N_13911);
nor U17143 (N_17143,N_15507,N_15969);
nor U17144 (N_17144,N_14963,N_15302);
nand U17145 (N_17145,N_12615,N_12121);
nor U17146 (N_17146,N_14134,N_14291);
or U17147 (N_17147,N_13736,N_13773);
nand U17148 (N_17148,N_12473,N_14801);
nand U17149 (N_17149,N_15869,N_14613);
nand U17150 (N_17150,N_15587,N_15133);
or U17151 (N_17151,N_12389,N_14184);
and U17152 (N_17152,N_13139,N_12472);
nor U17153 (N_17153,N_12291,N_13148);
or U17154 (N_17154,N_14382,N_12740);
or U17155 (N_17155,N_14223,N_15803);
nor U17156 (N_17156,N_13869,N_15786);
or U17157 (N_17157,N_12509,N_14681);
xor U17158 (N_17158,N_13575,N_14858);
nor U17159 (N_17159,N_14348,N_14711);
and U17160 (N_17160,N_15016,N_12837);
nand U17161 (N_17161,N_14825,N_12978);
or U17162 (N_17162,N_13414,N_12957);
xor U17163 (N_17163,N_14810,N_15513);
and U17164 (N_17164,N_15390,N_12313);
nor U17165 (N_17165,N_14472,N_13237);
nor U17166 (N_17166,N_14654,N_14415);
xnor U17167 (N_17167,N_13650,N_15942);
nand U17168 (N_17168,N_15884,N_14019);
nor U17169 (N_17169,N_14677,N_13101);
and U17170 (N_17170,N_14058,N_15914);
or U17171 (N_17171,N_14178,N_14751);
xnor U17172 (N_17172,N_14380,N_15436);
xnor U17173 (N_17173,N_14540,N_14302);
xnor U17174 (N_17174,N_15457,N_12755);
or U17175 (N_17175,N_13777,N_15766);
or U17176 (N_17176,N_13698,N_12879);
and U17177 (N_17177,N_14003,N_12648);
nor U17178 (N_17178,N_14838,N_14740);
nor U17179 (N_17179,N_14600,N_12710);
xnor U17180 (N_17180,N_14748,N_15079);
xor U17181 (N_17181,N_15830,N_15256);
xor U17182 (N_17182,N_14591,N_13013);
or U17183 (N_17183,N_15897,N_13502);
and U17184 (N_17184,N_15422,N_15888);
and U17185 (N_17185,N_13696,N_14701);
nand U17186 (N_17186,N_14771,N_14033);
or U17187 (N_17187,N_14587,N_15799);
nor U17188 (N_17188,N_13009,N_14899);
nand U17189 (N_17189,N_14123,N_14955);
xor U17190 (N_17190,N_13708,N_12819);
xor U17191 (N_17191,N_12697,N_13968);
and U17192 (N_17192,N_13024,N_13407);
and U17193 (N_17193,N_15019,N_14342);
nand U17194 (N_17194,N_13330,N_15404);
or U17195 (N_17195,N_12784,N_12749);
nor U17196 (N_17196,N_13524,N_15818);
nand U17197 (N_17197,N_14634,N_14760);
nand U17198 (N_17198,N_12327,N_12949);
xnor U17199 (N_17199,N_13839,N_13003);
nor U17200 (N_17200,N_15880,N_14434);
or U17201 (N_17201,N_14901,N_14396);
xnor U17202 (N_17202,N_13905,N_12692);
xor U17203 (N_17203,N_14632,N_14582);
and U17204 (N_17204,N_15847,N_13088);
and U17205 (N_17205,N_13141,N_12385);
xnor U17206 (N_17206,N_14235,N_12715);
or U17207 (N_17207,N_13963,N_12168);
or U17208 (N_17208,N_12546,N_15743);
nor U17209 (N_17209,N_12140,N_13085);
nor U17210 (N_17210,N_12885,N_13528);
xor U17211 (N_17211,N_14272,N_12912);
nand U17212 (N_17212,N_13098,N_13468);
nand U17213 (N_17213,N_13095,N_13779);
nand U17214 (N_17214,N_12804,N_14533);
xor U17215 (N_17215,N_15145,N_12003);
and U17216 (N_17216,N_15567,N_12191);
and U17217 (N_17217,N_14127,N_12769);
nor U17218 (N_17218,N_15824,N_13550);
or U17219 (N_17219,N_15239,N_15312);
or U17220 (N_17220,N_12234,N_12302);
xnor U17221 (N_17221,N_12758,N_12681);
nand U17222 (N_17222,N_15468,N_12803);
and U17223 (N_17223,N_14863,N_13670);
and U17224 (N_17224,N_14541,N_12894);
and U17225 (N_17225,N_14353,N_12983);
xnor U17226 (N_17226,N_14090,N_14852);
and U17227 (N_17227,N_15557,N_15252);
or U17228 (N_17228,N_15418,N_15525);
or U17229 (N_17229,N_14315,N_14244);
and U17230 (N_17230,N_12924,N_13875);
and U17231 (N_17231,N_15859,N_13411);
and U17232 (N_17232,N_14074,N_14565);
nand U17233 (N_17233,N_14949,N_15165);
and U17234 (N_17234,N_13924,N_14328);
xnor U17235 (N_17235,N_14737,N_13726);
xnor U17236 (N_17236,N_15871,N_14151);
nand U17237 (N_17237,N_15237,N_13682);
xnor U17238 (N_17238,N_12305,N_12488);
nor U17239 (N_17239,N_15362,N_13881);
nor U17240 (N_17240,N_13422,N_14645);
nand U17241 (N_17241,N_13691,N_13173);
and U17242 (N_17242,N_13860,N_15819);
nand U17243 (N_17243,N_12960,N_15635);
xnor U17244 (N_17244,N_14668,N_14440);
nand U17245 (N_17245,N_14229,N_14682);
or U17246 (N_17246,N_13930,N_13680);
xnor U17247 (N_17247,N_14699,N_13404);
or U17248 (N_17248,N_13508,N_12606);
xnor U17249 (N_17249,N_12446,N_15930);
nor U17250 (N_17250,N_13053,N_15299);
nand U17251 (N_17251,N_13800,N_15531);
xor U17252 (N_17252,N_14890,N_12811);
nand U17253 (N_17253,N_15482,N_14833);
and U17254 (N_17254,N_13218,N_14231);
nor U17255 (N_17255,N_13463,N_13458);
and U17256 (N_17256,N_15426,N_13713);
or U17257 (N_17257,N_14457,N_15541);
nor U17258 (N_17258,N_13363,N_13208);
xnor U17259 (N_17259,N_15520,N_12245);
nor U17260 (N_17260,N_12077,N_13113);
xnor U17261 (N_17261,N_15518,N_13213);
or U17262 (N_17262,N_12676,N_15066);
nor U17263 (N_17263,N_13214,N_12310);
xor U17264 (N_17264,N_15309,N_13320);
and U17265 (N_17265,N_13506,N_12483);
nand U17266 (N_17266,N_13025,N_13283);
xor U17267 (N_17267,N_14971,N_12504);
xor U17268 (N_17268,N_13038,N_14663);
and U17269 (N_17269,N_14162,N_13481);
nor U17270 (N_17270,N_15860,N_14931);
or U17271 (N_17271,N_14555,N_13247);
nand U17272 (N_17272,N_13459,N_14256);
and U17273 (N_17273,N_12892,N_15657);
xor U17274 (N_17274,N_15933,N_13844);
and U17275 (N_17275,N_14484,N_13032);
or U17276 (N_17276,N_13850,N_14504);
nand U17277 (N_17277,N_15953,N_15845);
and U17278 (N_17278,N_14144,N_13034);
xnor U17279 (N_17279,N_15172,N_14879);
or U17280 (N_17280,N_14390,N_15546);
nand U17281 (N_17281,N_13383,N_15300);
nand U17282 (N_17282,N_12265,N_14588);
xnor U17283 (N_17283,N_15973,N_14927);
or U17284 (N_17284,N_14539,N_13701);
xor U17285 (N_17285,N_14536,N_13114);
and U17286 (N_17286,N_15508,N_14374);
nand U17287 (N_17287,N_12644,N_14500);
xnor U17288 (N_17288,N_14305,N_12025);
nor U17289 (N_17289,N_13748,N_14495);
or U17290 (N_17290,N_12187,N_12415);
nor U17291 (N_17291,N_15619,N_13456);
nor U17292 (N_17292,N_12263,N_15064);
nor U17293 (N_17293,N_12192,N_14889);
and U17294 (N_17294,N_13803,N_12366);
xnor U17295 (N_17295,N_14481,N_12737);
nand U17296 (N_17296,N_14345,N_13604);
xor U17297 (N_17297,N_13797,N_12031);
or U17298 (N_17298,N_12431,N_12061);
and U17299 (N_17299,N_15684,N_12534);
and U17300 (N_17300,N_13248,N_15578);
nor U17301 (N_17301,N_12869,N_13591);
and U17302 (N_17302,N_12208,N_13231);
xnor U17303 (N_17303,N_14596,N_15554);
xor U17304 (N_17304,N_15911,N_12170);
and U17305 (N_17305,N_12444,N_12024);
xnor U17306 (N_17306,N_14607,N_15831);
or U17307 (N_17307,N_14670,N_14892);
nor U17308 (N_17308,N_13312,N_14986);
or U17309 (N_17309,N_15745,N_13932);
or U17310 (N_17310,N_14630,N_14687);
nand U17311 (N_17311,N_14846,N_14395);
and U17312 (N_17312,N_13621,N_14886);
and U17313 (N_17313,N_15543,N_13326);
or U17314 (N_17314,N_14218,N_13353);
nand U17315 (N_17315,N_14688,N_12289);
nor U17316 (N_17316,N_13862,N_12409);
xnor U17317 (N_17317,N_13894,N_13193);
xnor U17318 (N_17318,N_12670,N_13106);
xnor U17319 (N_17319,N_14926,N_13349);
nand U17320 (N_17320,N_14024,N_14933);
xor U17321 (N_17321,N_12235,N_14117);
nand U17322 (N_17322,N_15583,N_15695);
or U17323 (N_17323,N_13191,N_13310);
and U17324 (N_17324,N_14121,N_12989);
and U17325 (N_17325,N_12438,N_12255);
xor U17326 (N_17326,N_12578,N_14945);
and U17327 (N_17327,N_13768,N_12154);
nor U17328 (N_17328,N_15192,N_13641);
and U17329 (N_17329,N_13259,N_15075);
or U17330 (N_17330,N_12328,N_14426);
or U17331 (N_17331,N_14853,N_15433);
xor U17332 (N_17332,N_15932,N_15055);
nand U17333 (N_17333,N_13999,N_15240);
and U17334 (N_17334,N_13765,N_14034);
and U17335 (N_17335,N_12661,N_13042);
or U17336 (N_17336,N_14908,N_13336);
nor U17337 (N_17337,N_14245,N_12826);
nor U17338 (N_17338,N_14501,N_12583);
or U17339 (N_17339,N_12341,N_12953);
and U17340 (N_17340,N_12262,N_12918);
nand U17341 (N_17341,N_15561,N_13872);
or U17342 (N_17342,N_14013,N_15624);
or U17343 (N_17343,N_15701,N_13416);
nor U17344 (N_17344,N_12517,N_15232);
xor U17345 (N_17345,N_14075,N_15550);
nand U17346 (N_17346,N_15245,N_15963);
xor U17347 (N_17347,N_15944,N_12982);
or U17348 (N_17348,N_15202,N_14261);
nand U17349 (N_17349,N_15568,N_14098);
nand U17350 (N_17350,N_12496,N_13338);
xnor U17351 (N_17351,N_14530,N_12411);
xor U17352 (N_17352,N_14476,N_12642);
xnor U17353 (N_17353,N_12908,N_14605);
nor U17354 (N_17354,N_15095,N_12748);
and U17355 (N_17355,N_12652,N_13625);
nand U17356 (N_17356,N_15008,N_13944);
and U17357 (N_17357,N_13480,N_13219);
nand U17358 (N_17358,N_14170,N_14470);
xor U17359 (N_17359,N_12227,N_14567);
and U17360 (N_17360,N_14366,N_13657);
or U17361 (N_17361,N_12110,N_15083);
and U17362 (N_17362,N_15286,N_13626);
nand U17363 (N_17363,N_13136,N_14243);
or U17364 (N_17364,N_15377,N_12144);
or U17365 (N_17365,N_15372,N_14187);
or U17366 (N_17366,N_12984,N_12577);
and U17367 (N_17367,N_13702,N_14921);
or U17368 (N_17368,N_13122,N_13813);
and U17369 (N_17369,N_12250,N_13125);
nor U17370 (N_17370,N_15919,N_14213);
nand U17371 (N_17371,N_14936,N_12686);
nand U17372 (N_17372,N_15391,N_12945);
and U17373 (N_17373,N_15521,N_14643);
nand U17374 (N_17374,N_13815,N_14043);
and U17375 (N_17375,N_15329,N_14164);
or U17376 (N_17376,N_13808,N_15152);
and U17377 (N_17377,N_14351,N_12716);
nand U17378 (N_17378,N_13906,N_15313);
nand U17379 (N_17379,N_13317,N_14126);
nor U17380 (N_17380,N_14392,N_15862);
or U17381 (N_17381,N_14008,N_12600);
nor U17382 (N_17382,N_13376,N_14520);
xor U17383 (N_17383,N_13176,N_15196);
nor U17384 (N_17384,N_12909,N_12554);
and U17385 (N_17385,N_14375,N_14052);
or U17386 (N_17386,N_13322,N_13646);
or U17387 (N_17387,N_12764,N_13068);
nor U17388 (N_17388,N_12069,N_13443);
and U17389 (N_17389,N_13099,N_15259);
and U17390 (N_17390,N_14311,N_12148);
nor U17391 (N_17391,N_12916,N_15189);
xor U17392 (N_17392,N_14409,N_14764);
nor U17393 (N_17393,N_14001,N_13566);
nor U17394 (N_17394,N_15163,N_14301);
nand U17395 (N_17395,N_14716,N_13870);
or U17396 (N_17396,N_15823,N_14743);
nand U17397 (N_17397,N_12434,N_13351);
nor U17398 (N_17398,N_14916,N_13235);
or U17399 (N_17399,N_13008,N_15674);
nor U17400 (N_17400,N_15199,N_12163);
nand U17401 (N_17401,N_12934,N_15175);
and U17402 (N_17402,N_15247,N_13360);
nor U17403 (N_17403,N_13230,N_13615);
and U17404 (N_17404,N_15121,N_12958);
and U17405 (N_17405,N_14640,N_12825);
nor U17406 (N_17406,N_12013,N_12852);
nand U17407 (N_17407,N_12229,N_15110);
xnor U17408 (N_17408,N_15903,N_13887);
xnor U17409 (N_17409,N_13603,N_14627);
xor U17410 (N_17410,N_15339,N_15912);
nand U17411 (N_17411,N_14002,N_14385);
nor U17412 (N_17412,N_12903,N_14049);
xor U17413 (N_17413,N_13819,N_15533);
nor U17414 (N_17414,N_12062,N_15116);
and U17415 (N_17415,N_13423,N_15378);
nand U17416 (N_17416,N_13525,N_13381);
or U17417 (N_17417,N_12010,N_12307);
and U17418 (N_17418,N_13118,N_12621);
xnor U17419 (N_17419,N_14314,N_13600);
and U17420 (N_17420,N_12464,N_14689);
and U17421 (N_17421,N_15651,N_14035);
nor U17422 (N_17422,N_12002,N_12757);
nand U17423 (N_17423,N_15323,N_15092);
nor U17424 (N_17424,N_15856,N_12539);
nand U17425 (N_17425,N_15599,N_14546);
and U17426 (N_17426,N_14474,N_14174);
xor U17427 (N_17427,N_12675,N_13897);
or U17428 (N_17428,N_14192,N_12416);
nor U17429 (N_17429,N_12070,N_15770);
and U17430 (N_17430,N_14942,N_13904);
nor U17431 (N_17431,N_12522,N_14802);
nand U17432 (N_17432,N_13420,N_13672);
nand U17433 (N_17433,N_15194,N_13689);
xnor U17434 (N_17434,N_14980,N_12766);
and U17435 (N_17435,N_15597,N_12651);
nand U17436 (N_17436,N_15975,N_15719);
or U17437 (N_17437,N_14806,N_12051);
nor U17438 (N_17438,N_13884,N_14194);
and U17439 (N_17439,N_14957,N_13123);
and U17440 (N_17440,N_14438,N_14455);
nor U17441 (N_17441,N_14577,N_13536);
or U17442 (N_17442,N_13927,N_13275);
nor U17443 (N_17443,N_15434,N_12200);
and U17444 (N_17444,N_13030,N_15276);
nand U17445 (N_17445,N_13465,N_14491);
nand U17446 (N_17446,N_14372,N_12474);
xnor U17447 (N_17447,N_13780,N_13043);
xnor U17448 (N_17448,N_15029,N_14947);
and U17449 (N_17449,N_12498,N_12834);
and U17450 (N_17450,N_14912,N_13454);
xor U17451 (N_17451,N_13804,N_15731);
nor U17452 (N_17452,N_12502,N_14928);
and U17453 (N_17453,N_12015,N_14105);
and U17454 (N_17454,N_13155,N_14960);
xnor U17455 (N_17455,N_13545,N_14683);
or U17456 (N_17456,N_13756,N_15143);
xor U17457 (N_17457,N_14729,N_13490);
nor U17458 (N_17458,N_12132,N_14247);
and U17459 (N_17459,N_12239,N_14293);
nand U17460 (N_17460,N_15727,N_14835);
nand U17461 (N_17461,N_12601,N_14010);
xnor U17462 (N_17462,N_12973,N_14615);
nor U17463 (N_17463,N_14159,N_14629);
or U17464 (N_17464,N_13693,N_13936);
nand U17465 (N_17465,N_15316,N_13309);
and U17466 (N_17466,N_12781,N_13864);
nor U17467 (N_17467,N_14909,N_15697);
or U17468 (N_17468,N_15005,N_13707);
or U17469 (N_17469,N_14490,N_13094);
nand U17470 (N_17470,N_15774,N_12440);
nand U17471 (N_17471,N_15667,N_12726);
nand U17472 (N_17472,N_13440,N_15326);
xor U17473 (N_17473,N_14282,N_14671);
nand U17474 (N_17474,N_15923,N_12883);
nand U17475 (N_17475,N_12864,N_13526);
or U17476 (N_17476,N_13267,N_14884);
and U17477 (N_17477,N_15236,N_14373);
xor U17478 (N_17478,N_13908,N_15136);
or U17479 (N_17479,N_13418,N_14197);
and U17480 (N_17480,N_14386,N_13843);
nor U17481 (N_17481,N_14559,N_13735);
xnor U17482 (N_17482,N_12343,N_15087);
or U17483 (N_17483,N_12429,N_15486);
and U17484 (N_17484,N_15890,N_14119);
nand U17485 (N_17485,N_12999,N_13290);
and U17486 (N_17486,N_15385,N_13103);
xor U17487 (N_17487,N_12269,N_12917);
and U17488 (N_17488,N_12146,N_13919);
or U17489 (N_17489,N_12129,N_14377);
and U17490 (N_17490,N_13711,N_14203);
xor U17491 (N_17491,N_15559,N_12662);
and U17492 (N_17492,N_13725,N_12037);
xnor U17493 (N_17493,N_13706,N_15347);
and U17494 (N_17494,N_12222,N_14237);
or U17495 (N_17495,N_15059,N_12636);
nand U17496 (N_17496,N_12159,N_15676);
or U17497 (N_17497,N_15458,N_14676);
or U17498 (N_17498,N_15811,N_13838);
and U17499 (N_17499,N_14974,N_12330);
and U17500 (N_17500,N_15720,N_12975);
nand U17501 (N_17501,N_13444,N_15074);
or U17502 (N_17502,N_12911,N_15787);
and U17503 (N_17503,N_14997,N_14686);
xor U17504 (N_17504,N_12671,N_15538);
xnor U17505 (N_17505,N_14844,N_14094);
nand U17506 (N_17506,N_13156,N_15837);
nand U17507 (N_17507,N_13562,N_13861);
and U17508 (N_17508,N_13572,N_13397);
and U17509 (N_17509,N_12098,N_13164);
nand U17510 (N_17510,N_12877,N_12074);
nor U17511 (N_17511,N_12349,N_15473);
nor U17512 (N_17512,N_12624,N_14106);
and U17513 (N_17513,N_12687,N_14531);
nor U17514 (N_17514,N_12321,N_14444);
xnor U17515 (N_17515,N_13825,N_14202);
and U17516 (N_17516,N_15420,N_15432);
and U17517 (N_17517,N_14198,N_13479);
and U17518 (N_17518,N_14355,N_15925);
nor U17519 (N_17519,N_14283,N_14732);
or U17520 (N_17520,N_14967,N_15164);
nand U17521 (N_17521,N_13415,N_13225);
or U17522 (N_17522,N_13432,N_13187);
or U17523 (N_17523,N_12528,N_12213);
xnor U17524 (N_17524,N_15601,N_14993);
and U17525 (N_17525,N_12632,N_12160);
or U17526 (N_17526,N_12775,N_12512);
nor U17527 (N_17527,N_12124,N_14915);
and U17528 (N_17528,N_15266,N_14524);
or U17529 (N_17529,N_15729,N_14310);
nor U17530 (N_17530,N_15485,N_12233);
and U17531 (N_17531,N_14548,N_12538);
xor U17532 (N_17532,N_14581,N_12232);
nor U17533 (N_17533,N_14350,N_15287);
xnor U17534 (N_17534,N_13654,N_13821);
nor U17535 (N_17535,N_12361,N_14165);
nor U17536 (N_17536,N_13557,N_13959);
nand U17537 (N_17537,N_13424,N_13149);
and U17538 (N_17538,N_15797,N_15852);
or U17539 (N_17539,N_14660,N_13426);
xor U17540 (N_17540,N_13239,N_14211);
and U17541 (N_17541,N_12220,N_12952);
and U17542 (N_17542,N_13885,N_13199);
nor U17543 (N_17543,N_14062,N_12801);
xnor U17544 (N_17544,N_13584,N_14383);
xnor U17545 (N_17545,N_13916,N_15288);
or U17546 (N_17546,N_15976,N_15558);
nand U17547 (N_17547,N_13161,N_15675);
or U17548 (N_17548,N_14579,N_12181);
nand U17549 (N_17549,N_12099,N_15540);
and U17550 (N_17550,N_14266,N_14149);
xnor U17551 (N_17551,N_15454,N_14469);
xnor U17552 (N_17552,N_13181,N_15449);
xnor U17553 (N_17553,N_14592,N_13967);
or U17554 (N_17554,N_13462,N_14333);
xnor U17555 (N_17555,N_12417,N_12306);
nor U17556 (N_17556,N_14259,N_15691);
xor U17557 (N_17557,N_14569,N_12765);
nand U17558 (N_17558,N_13180,N_13941);
or U17559 (N_17559,N_14154,N_13956);
and U17560 (N_17560,N_12065,N_15170);
xnor U17561 (N_17561,N_15959,N_14079);
xor U17562 (N_17562,N_14346,N_14428);
xor U17563 (N_17563,N_15389,N_14635);
and U17564 (N_17564,N_14046,N_14424);
or U17565 (N_17565,N_12586,N_15212);
xor U17566 (N_17566,N_14830,N_13648);
and U17567 (N_17567,N_13086,N_12465);
nand U17568 (N_17568,N_12436,N_15224);
and U17569 (N_17569,N_15042,N_14253);
nor U17570 (N_17570,N_12896,N_14269);
nor U17571 (N_17571,N_14882,N_12729);
nor U17572 (N_17572,N_14561,N_14788);
nor U17573 (N_17573,N_13315,N_14175);
xor U17574 (N_17574,N_14989,N_12041);
nor U17575 (N_17575,N_14209,N_14545);
nand U17576 (N_17576,N_15446,N_12034);
xor U17577 (N_17577,N_12817,N_14221);
or U17578 (N_17578,N_15255,N_13354);
xor U17579 (N_17579,N_14700,N_15102);
nand U17580 (N_17580,N_15089,N_15647);
and U17581 (N_17581,N_13655,N_13816);
xnor U17582 (N_17582,N_13018,N_12533);
or U17583 (N_17583,N_12567,N_13255);
or U17584 (N_17584,N_14136,N_12258);
xor U17585 (N_17585,N_14447,N_15505);
nor U17586 (N_17586,N_12127,N_12878);
xor U17587 (N_17587,N_12252,N_13348);
nor U17588 (N_17588,N_12694,N_15858);
xnor U17589 (N_17589,N_13926,N_15967);
xnor U17590 (N_17590,N_13549,N_15709);
nor U17591 (N_17591,N_12221,N_15582);
nor U17592 (N_17592,N_14907,N_13997);
xor U17593 (N_17593,N_13759,N_15159);
nor U17594 (N_17594,N_13130,N_14991);
or U17595 (N_17595,N_12707,N_13110);
or U17596 (N_17596,N_15927,N_15162);
xnor U17597 (N_17597,N_15474,N_15671);
nor U17598 (N_17598,N_15070,N_15306);
and U17599 (N_17599,N_13050,N_12582);
or U17600 (N_17600,N_15591,N_15878);
nor U17601 (N_17601,N_12454,N_14851);
nor U17602 (N_17602,N_12573,N_15398);
or U17603 (N_17603,N_12569,N_15982);
xnor U17604 (N_17604,N_12657,N_12536);
and U17605 (N_17605,N_15730,N_12752);
xor U17606 (N_17606,N_14950,N_15579);
nand U17607 (N_17607,N_14446,N_14954);
xnor U17608 (N_17608,N_12087,N_12847);
nor U17609 (N_17609,N_13618,N_14937);
nand U17610 (N_17610,N_15076,N_13612);
nor U17611 (N_17611,N_13595,N_14289);
xnor U17612 (N_17612,N_12643,N_14953);
nand U17613 (N_17613,N_12463,N_12084);
xor U17614 (N_17614,N_15806,N_14978);
nand U17615 (N_17615,N_15456,N_13077);
and U17616 (N_17616,N_12620,N_14487);
or U17617 (N_17617,N_12001,N_13151);
nand U17618 (N_17618,N_12519,N_13504);
nor U17619 (N_17619,N_15755,N_13243);
or U17620 (N_17620,N_13347,N_12501);
nor U17621 (N_17621,N_13937,N_15820);
xor U17622 (N_17622,N_15699,N_14762);
nand U17623 (N_17623,N_14733,N_14439);
nor U17624 (N_17624,N_13833,N_12926);
nand U17625 (N_17625,N_13496,N_15429);
and U17626 (N_17626,N_14821,N_13240);
nand U17627 (N_17627,N_14573,N_15217);
nand U17628 (N_17628,N_14952,N_12183);
nand U17629 (N_17629,N_15764,N_12350);
or U17630 (N_17630,N_13683,N_12369);
nor U17631 (N_17631,N_12700,N_13737);
nand U17632 (N_17632,N_12531,N_13289);
xnor U17633 (N_17633,N_14509,N_13530);
nand U17634 (N_17634,N_13260,N_13786);
nand U17635 (N_17635,N_13985,N_12677);
or U17636 (N_17636,N_15085,N_14464);
or U17637 (N_17637,N_15736,N_13983);
xor U17638 (N_17638,N_13685,N_13532);
nor U17639 (N_17639,N_14028,N_12189);
nor U17640 (N_17640,N_14408,N_12992);
or U17641 (N_17641,N_13345,N_13980);
or U17642 (N_17642,N_13871,N_15526);
nand U17643 (N_17643,N_15104,N_12809);
or U17644 (N_17644,N_13205,N_12295);
and U17645 (N_17645,N_15495,N_14177);
nand U17646 (N_17646,N_15265,N_13888);
nor U17647 (N_17647,N_15913,N_14616);
xor U17648 (N_17648,N_14970,N_13840);
xor U17649 (N_17649,N_13460,N_15215);
and U17650 (N_17650,N_14693,N_13410);
and U17651 (N_17651,N_14494,N_12261);
and U17652 (N_17652,N_12028,N_15167);
or U17653 (N_17653,N_13441,N_14497);
xnor U17654 (N_17654,N_12372,N_15223);
xnor U17655 (N_17655,N_14176,N_14932);
xor U17656 (N_17656,N_13961,N_14214);
nand U17657 (N_17657,N_12314,N_15714);
nand U17658 (N_17658,N_15455,N_14964);
and U17659 (N_17659,N_13069,N_12378);
or U17660 (N_17660,N_14554,N_13171);
or U17661 (N_17661,N_14265,N_15150);
or U17662 (N_17662,N_12800,N_12118);
nor U17663 (N_17663,N_13144,N_13120);
nand U17664 (N_17664,N_13132,N_15157);
and U17665 (N_17665,N_14263,N_14763);
nand U17666 (N_17666,N_12814,N_15091);
nor U17667 (N_17667,N_14973,N_14666);
nor U17668 (N_17668,N_15077,N_12186);
nand U17669 (N_17669,N_14199,N_14422);
and U17670 (N_17670,N_15992,N_15650);
and U17671 (N_17671,N_13216,N_15174);
and U17672 (N_17672,N_13535,N_14452);
or U17673 (N_17673,N_15169,N_15602);
or U17674 (N_17674,N_13152,N_12254);
or U17675 (N_17675,N_12625,N_12419);
nand U17676 (N_17676,N_12511,N_15363);
nor U17677 (N_17677,N_12175,N_14044);
nand U17678 (N_17678,N_13917,N_12214);
xnor U17679 (N_17679,N_15722,N_12599);
nor U17680 (N_17680,N_14715,N_14925);
xnor U17681 (N_17681,N_15796,N_12986);
or U17682 (N_17682,N_15279,N_15536);
and U17683 (N_17683,N_14988,N_12572);
and U17684 (N_17684,N_14207,N_13928);
nor U17685 (N_17685,N_15947,N_14116);
nor U17686 (N_17686,N_13186,N_12994);
and U17687 (N_17687,N_15084,N_14526);
xor U17688 (N_17688,N_12348,N_13396);
nand U17689 (N_17689,N_13206,N_12193);
or U17690 (N_17690,N_15315,N_15277);
nand U17691 (N_17691,N_12111,N_14369);
nor U17692 (N_17692,N_15612,N_13729);
nand U17693 (N_17693,N_12403,N_15195);
nor U17694 (N_17694,N_13273,N_15734);
nor U17695 (N_17695,N_15290,N_12870);
nand U17696 (N_17696,N_13745,N_15493);
and U17697 (N_17697,N_14222,N_14454);
nand U17698 (N_17698,N_15371,N_13303);
xnor U17699 (N_17699,N_14505,N_14156);
nor U17700 (N_17700,N_14267,N_12780);
xor U17701 (N_17701,N_15782,N_13610);
nand U17702 (N_17702,N_12907,N_15357);
nor U17703 (N_17703,N_14021,N_15983);
nand U17704 (N_17704,N_14637,N_15107);
nor U17705 (N_17705,N_13695,N_13953);
and U17706 (N_17706,N_15067,N_14026);
or U17707 (N_17707,N_15931,N_14326);
xor U17708 (N_17708,N_14362,N_12340);
nor U17709 (N_17709,N_15816,N_12063);
xor U17710 (N_17710,N_12720,N_13519);
and U17711 (N_17711,N_12164,N_14249);
nor U17712 (N_17712,N_13093,N_15984);
nand U17713 (N_17713,N_13993,N_14224);
nor U17714 (N_17714,N_13579,N_14589);
and U17715 (N_17715,N_12153,N_13541);
xnor U17716 (N_17716,N_14186,N_13059);
and U17717 (N_17717,N_12128,N_12178);
nor U17718 (N_17718,N_12243,N_15320);
and U17719 (N_17719,N_12231,N_12106);
and U17720 (N_17720,N_14944,N_15654);
xnor U17721 (N_17721,N_12157,N_14384);
xor U17722 (N_17722,N_12049,N_12152);
xnor U17723 (N_17723,N_13105,N_15961);
nor U17724 (N_17724,N_12976,N_12515);
nand U17725 (N_17725,N_12923,N_15833);
xnor U17726 (N_17726,N_15118,N_12838);
or U17727 (N_17727,N_15057,N_15046);
and U17728 (N_17728,N_13263,N_15337);
nand U17729 (N_17729,N_12280,N_15058);
or U17730 (N_17730,N_13031,N_14274);
xnor U17731 (N_17731,N_14769,N_14147);
xnor U17732 (N_17732,N_13520,N_12876);
xnor U17733 (N_17733,N_14318,N_12714);
nor U17734 (N_17734,N_13664,N_12971);
xnor U17735 (N_17735,N_15825,N_14048);
xor U17736 (N_17736,N_12377,N_12478);
nor U17737 (N_17737,N_13697,N_14795);
and U17738 (N_17738,N_14143,N_15633);
xnor U17739 (N_17739,N_13970,N_15098);
nand U17740 (N_17740,N_15643,N_13700);
xnor U17741 (N_17741,N_15936,N_15291);
and U17742 (N_17742,N_15781,N_13543);
nand U17743 (N_17743,N_12505,N_13679);
and U17744 (N_17744,N_13782,N_13660);
or U17745 (N_17745,N_14585,N_13332);
or U17746 (N_17746,N_14179,N_12449);
xnor U17747 (N_17747,N_14459,N_13065);
xnor U17748 (N_17748,N_13374,N_15125);
nand U17749 (N_17749,N_14888,N_13912);
or U17750 (N_17750,N_12650,N_15171);
nor U17751 (N_17751,N_12997,N_12493);
xnor U17752 (N_17752,N_13232,N_13448);
and U17753 (N_17753,N_13398,N_14608);
or U17754 (N_17754,N_13857,N_13382);
and U17755 (N_17755,N_13220,N_14680);
or U17756 (N_17756,N_15891,N_15218);
nor U17757 (N_17757,N_14707,N_14216);
and U17758 (N_17758,N_12712,N_14250);
xnor U17759 (N_17759,N_15544,N_12668);
or U17760 (N_17760,N_13955,N_12381);
or U17761 (N_17761,N_12435,N_15105);
and U17762 (N_17762,N_14096,N_12006);
nor U17763 (N_17763,N_14189,N_12135);
nand U17764 (N_17764,N_12610,N_13108);
nor U17765 (N_17765,N_13133,N_12117);
xor U17766 (N_17766,N_12713,N_13753);
or U17767 (N_17767,N_15001,N_14574);
xor U17768 (N_17768,N_15843,N_13340);
and U17769 (N_17769,N_12702,N_15154);
and U17770 (N_17770,N_15294,N_14065);
nand U17771 (N_17771,N_13533,N_13146);
nor U17772 (N_17772,N_14650,N_15894);
or U17773 (N_17773,N_13321,N_14741);
and U17774 (N_17774,N_15981,N_12529);
xnor U17775 (N_17775,N_12935,N_13515);
and U17776 (N_17776,N_12122,N_13592);
or U17777 (N_17777,N_14941,N_12827);
nor U17778 (N_17778,N_14794,N_13389);
nor U17779 (N_17779,N_15469,N_14092);
or U17780 (N_17780,N_15344,N_14883);
and U17781 (N_17781,N_12055,N_15024);
xor U17782 (N_17782,N_15670,N_12943);
and U17783 (N_17783,N_12905,N_14445);
xnor U17784 (N_17784,N_13211,N_14783);
and U17785 (N_17785,N_12333,N_12630);
and U17786 (N_17786,N_14341,N_15068);
and U17787 (N_17787,N_15069,N_12104);
xor U17788 (N_17788,N_14791,N_13597);
and U17789 (N_17789,N_13553,N_15186);
or U17790 (N_17790,N_12948,N_12082);
nor U17791 (N_17791,N_13977,N_15428);
or U17792 (N_17792,N_15401,N_13649);
nand U17793 (N_17793,N_13676,N_12608);
nor U17794 (N_17794,N_14556,N_12937);
nand U17795 (N_17795,N_14800,N_12711);
xnor U17796 (N_17796,N_13258,N_13663);
and U17797 (N_17797,N_12808,N_13658);
or U17798 (N_17798,N_12566,N_12576);
and U17799 (N_17799,N_13491,N_15716);
or U17800 (N_17800,N_15310,N_15080);
or U17801 (N_17801,N_15842,N_14773);
or U17802 (N_17802,N_13988,N_14930);
xor U17803 (N_17803,N_15298,N_12172);
nand U17804 (N_17804,N_14655,N_15100);
or U17805 (N_17805,N_15435,N_13951);
xnor U17806 (N_17806,N_13408,N_12635);
and U17807 (N_17807,N_15340,N_12445);
nor U17808 (N_17808,N_13168,N_12470);
nor U17809 (N_17809,N_15603,N_14361);
or U17810 (N_17810,N_12688,N_14185);
nand U17811 (N_17811,N_14639,N_14977);
nand U17812 (N_17812,N_12927,N_14360);
nand U17813 (N_17813,N_12495,N_13313);
and U17814 (N_17814,N_15244,N_12395);
nor U17815 (N_17815,N_12537,N_14761);
xnor U17816 (N_17816,N_14685,N_13238);
nor U17817 (N_17817,N_12450,N_14405);
or U17818 (N_17818,N_12684,N_12724);
nor U17819 (N_17819,N_14813,N_14723);
xor U17820 (N_17820,N_12334,N_13419);
nand U17821 (N_17821,N_12248,N_13593);
or U17822 (N_17822,N_15097,N_15515);
nor U17823 (N_17823,N_13518,N_15226);
xnor U17824 (N_17824,N_15576,N_15639);
xnor U17825 (N_17825,N_14275,N_13560);
and U17826 (N_17826,N_15861,N_13521);
xor U17827 (N_17827,N_15590,N_12080);
nand U17828 (N_17828,N_15325,N_13558);
or U17829 (N_17829,N_13249,N_12370);
or U17830 (N_17830,N_13464,N_13241);
and U17831 (N_17831,N_14102,N_13001);
xnor U17832 (N_17832,N_15480,N_15444);
nor U17833 (N_17833,N_15629,N_15035);
nand U17834 (N_17834,N_14418,N_12535);
xnor U17835 (N_17835,N_13256,N_12756);
xnor U17836 (N_17836,N_12392,N_13940);
nor U17837 (N_17837,N_13613,N_15524);
nor U17838 (N_17838,N_14022,N_13337);
or U17839 (N_17839,N_12408,N_14352);
xnor U17840 (N_17840,N_12169,N_12513);
nand U17841 (N_17841,N_13681,N_13692);
or U17842 (N_17842,N_13153,N_15405);
xnor U17843 (N_17843,N_13198,N_15542);
and U17844 (N_17844,N_13467,N_13673);
nand U17845 (N_17845,N_13041,N_12747);
or U17846 (N_17846,N_12888,N_15611);
or U17847 (N_17847,N_15129,N_12329);
nor U17848 (N_17848,N_13640,N_13775);
xor U17849 (N_17849,N_14171,N_15466);
xnor U17850 (N_17850,N_12332,N_14006);
xnor U17851 (N_17851,N_12319,N_12007);
nor U17852 (N_17852,N_12073,N_15356);
or U17853 (N_17853,N_12967,N_13561);
and U17854 (N_17854,N_14919,N_14236);
or U17855 (N_17855,N_14747,N_14831);
nand U17856 (N_17856,N_13035,N_15589);
xor U17857 (N_17857,N_13509,N_12477);
and U17858 (N_17858,N_13712,N_12969);
nand U17859 (N_17859,N_15877,N_15712);
nor U17860 (N_17860,N_13307,N_15906);
or U17861 (N_17861,N_15767,N_14053);
nand U17862 (N_17862,N_14829,N_15646);
and U17863 (N_17863,N_12790,N_13958);
or U17864 (N_17864,N_14242,N_12500);
and U17865 (N_17865,N_14331,N_15950);
nand U17866 (N_17866,N_14125,N_12299);
nand U17867 (N_17867,N_13879,N_15648);
nand U17868 (N_17868,N_15710,N_12858);
xnor U17869 (N_17869,N_12391,N_12068);
or U17870 (N_17870,N_12453,N_14336);
or U17871 (N_17871,N_12081,N_14659);
or U17872 (N_17872,N_15253,N_13201);
or U17873 (N_17873,N_12968,N_15703);
nand U17874 (N_17874,N_15575,N_14599);
nand U17875 (N_17875,N_13741,N_12570);
and U17876 (N_17876,N_13483,N_15885);
xnor U17877 (N_17877,N_13922,N_13178);
nor U17878 (N_17878,N_14220,N_12639);
xnor U17879 (N_17879,N_12486,N_15205);
nand U17880 (N_17880,N_12928,N_12241);
xnor U17881 (N_17881,N_13776,N_12761);
nor U17882 (N_17882,N_13318,N_14697);
nor U17883 (N_17883,N_14638,N_14506);
nor U17884 (N_17884,N_15453,N_12094);
nand U17885 (N_17885,N_15661,N_14578);
nor U17886 (N_17886,N_14292,N_14234);
xnor U17887 (N_17887,N_12701,N_13909);
nor U17888 (N_17888,N_14303,N_12589);
nor U17889 (N_17889,N_13183,N_14617);
nand U17890 (N_17890,N_15746,N_13294);
xor U17891 (N_17891,N_14473,N_15060);
and U17892 (N_17892,N_15956,N_13165);
nor U17893 (N_17893,N_15594,N_15839);
nor U17894 (N_17894,N_14485,N_15296);
nand U17895 (N_17895,N_15376,N_12787);
nor U17896 (N_17896,N_13837,N_12795);
nor U17897 (N_17897,N_14061,N_12085);
nand U17898 (N_17898,N_15114,N_13966);
nand U17899 (N_17899,N_13052,N_14824);
and U17900 (N_17900,N_14413,N_13975);
nor U17901 (N_17901,N_15998,N_14534);
or U17902 (N_17902,N_12640,N_13357);
and U17903 (N_17903,N_15990,N_13517);
and U17904 (N_17904,N_12732,N_15740);
xnor U17905 (N_17905,N_14512,N_13109);
nand U17906 (N_17906,N_12288,N_13981);
or U17907 (N_17907,N_15566,N_13075);
xnor U17908 (N_17908,N_12562,N_15274);
nand U17909 (N_17909,N_12297,N_14837);
nor U17910 (N_17910,N_14855,N_15548);
nand U17911 (N_17911,N_13304,N_14586);
or U17912 (N_17912,N_12374,N_15641);
xor U17913 (N_17913,N_13730,N_14752);
nor U17914 (N_17914,N_12745,N_15151);
nand U17915 (N_17915,N_12785,N_15366);
and U17916 (N_17916,N_14618,N_15649);
and U17917 (N_17917,N_15392,N_15011);
or U17918 (N_17918,N_12179,N_12353);
nand U17919 (N_17919,N_12991,N_14644);
or U17920 (N_17920,N_14498,N_13534);
and U17921 (N_17921,N_12848,N_14641);
xnor U17922 (N_17922,N_13982,N_12862);
xor U17923 (N_17923,N_15762,N_14488);
nor U17924 (N_17924,N_13984,N_14958);
nor U17925 (N_17925,N_13277,N_12793);
and U17926 (N_17926,N_12956,N_12966);
xor U17927 (N_17927,N_12840,N_14868);
nand U17928 (N_17928,N_14461,N_13447);
nor U17929 (N_17929,N_14060,N_13323);
or U17930 (N_17930,N_13772,N_14735);
nor U17931 (N_17931,N_13762,N_13000);
nand U17932 (N_17932,N_15790,N_12102);
xnor U17933 (N_17933,N_13477,N_14867);
nor U17934 (N_17934,N_14814,N_15682);
and U17935 (N_17935,N_15414,N_12123);
nor U17936 (N_17936,N_12914,N_15841);
and U17937 (N_17937,N_15728,N_12646);
and U17938 (N_17938,N_15257,N_14441);
or U17939 (N_17939,N_12882,N_15348);
nor U17940 (N_17940,N_12442,N_13333);
and U17941 (N_17941,N_13948,N_15838);
or U17942 (N_17942,N_12004,N_14777);
nor U17943 (N_17943,N_14721,N_13751);
nor U17944 (N_17944,N_12316,N_13880);
or U17945 (N_17945,N_14745,N_12762);
and U17946 (N_17946,N_13486,N_12660);
nand U17947 (N_17947,N_14789,N_12590);
nand U17948 (N_17948,N_13868,N_12161);
and U17949 (N_17949,N_15013,N_12060);
nand U17950 (N_17950,N_14037,N_13556);
or U17951 (N_17951,N_15308,N_15327);
nand U17952 (N_17952,N_13589,N_14018);
nor U17953 (N_17953,N_13393,N_15203);
xnor U17954 (N_17954,N_12930,N_14896);
or U17955 (N_17955,N_15958,N_14071);
nor U17956 (N_17956,N_12264,N_15023);
or U17957 (N_17957,N_12137,N_14727);
nand U17958 (N_17958,N_14621,N_15263);
and U17959 (N_17959,N_15563,N_12246);
xnor U17960 (N_17960,N_15949,N_14595);
and U17961 (N_17961,N_12664,N_13639);
and U17962 (N_17962,N_14279,N_13334);
and U17963 (N_17963,N_15669,N_14601);
xnor U17964 (N_17964,N_12587,N_14152);
nand U17965 (N_17965,N_12195,N_12090);
and U17966 (N_17966,N_14754,N_15623);
and U17967 (N_17967,N_12242,N_15460);
and U17968 (N_17968,N_14877,N_14734);
nand U17969 (N_17969,N_12521,N_15198);
nor U17970 (N_17970,N_14299,N_13617);
and U17971 (N_17971,N_15915,N_14321);
nand U17972 (N_17972,N_15620,N_15108);
and U17973 (N_17973,N_13045,N_13224);
nand U17974 (N_17974,N_14296,N_12345);
and U17975 (N_17975,N_14080,N_15353);
or U17976 (N_17976,N_15988,N_15827);
and U17977 (N_17977,N_13754,N_14183);
nor U17978 (N_17978,N_15409,N_14157);
and U17979 (N_17979,N_15333,N_15028);
or U17980 (N_17980,N_12830,N_12921);
xnor U17981 (N_17981,N_14421,N_13677);
nand U17982 (N_17982,N_15829,N_12865);
nand U17983 (N_17983,N_13299,N_15062);
nand U17984 (N_17984,N_14609,N_14340);
xnor U17985 (N_17985,N_12420,N_12946);
or U17986 (N_17986,N_13373,N_15807);
or U17987 (N_17987,N_12339,N_15368);
and U17988 (N_17988,N_15322,N_13112);
and U17989 (N_17989,N_14691,N_13092);
and U17990 (N_17990,N_15496,N_14496);
nand U17991 (N_17991,N_12331,N_12045);
nor U17992 (N_17992,N_12859,N_13474);
nor U17993 (N_17993,N_15814,N_12782);
and U17994 (N_17994,N_13040,N_12275);
xnor U17995 (N_17995,N_14041,N_15547);
nand U17996 (N_17996,N_15615,N_13469);
or U17997 (N_17997,N_15951,N_15491);
and U17998 (N_17998,N_12985,N_15908);
and U17999 (N_17999,N_14483,N_15379);
xnor U18000 (N_18000,N_14796,N_13227);
nand U18001 (N_18001,N_13158,N_12517);
nand U18002 (N_18002,N_12318,N_12539);
nor U18003 (N_18003,N_12472,N_12258);
and U18004 (N_18004,N_14830,N_12265);
xor U18005 (N_18005,N_14811,N_12210);
and U18006 (N_18006,N_15781,N_13447);
nand U18007 (N_18007,N_15739,N_12910);
nor U18008 (N_18008,N_15604,N_15403);
nand U18009 (N_18009,N_13685,N_15154);
and U18010 (N_18010,N_12494,N_15971);
nand U18011 (N_18011,N_13391,N_12225);
xor U18012 (N_18012,N_12415,N_14817);
nor U18013 (N_18013,N_13064,N_15133);
or U18014 (N_18014,N_14428,N_14417);
nor U18015 (N_18015,N_13673,N_13190);
xnor U18016 (N_18016,N_12278,N_14305);
xnor U18017 (N_18017,N_13448,N_12898);
and U18018 (N_18018,N_15576,N_13409);
xnor U18019 (N_18019,N_12143,N_15492);
or U18020 (N_18020,N_15560,N_12371);
and U18021 (N_18021,N_15005,N_14920);
and U18022 (N_18022,N_13165,N_13320);
xor U18023 (N_18023,N_13317,N_12918);
nor U18024 (N_18024,N_13335,N_12157);
or U18025 (N_18025,N_14277,N_12396);
and U18026 (N_18026,N_13962,N_13678);
xnor U18027 (N_18027,N_13489,N_12111);
or U18028 (N_18028,N_15935,N_13896);
and U18029 (N_18029,N_14345,N_15326);
or U18030 (N_18030,N_15780,N_12430);
nand U18031 (N_18031,N_13800,N_15428);
nor U18032 (N_18032,N_13812,N_12778);
xnor U18033 (N_18033,N_14201,N_12644);
and U18034 (N_18034,N_15080,N_14673);
xnor U18035 (N_18035,N_13341,N_13330);
nand U18036 (N_18036,N_12262,N_12846);
nand U18037 (N_18037,N_12168,N_13183);
xnor U18038 (N_18038,N_12731,N_14465);
nor U18039 (N_18039,N_15587,N_13963);
or U18040 (N_18040,N_12478,N_13125);
nor U18041 (N_18041,N_13823,N_12921);
xor U18042 (N_18042,N_15017,N_15942);
or U18043 (N_18043,N_15684,N_14389);
and U18044 (N_18044,N_15581,N_13637);
xnor U18045 (N_18045,N_15483,N_12439);
xnor U18046 (N_18046,N_15387,N_12226);
nor U18047 (N_18047,N_12695,N_14617);
and U18048 (N_18048,N_13955,N_14074);
and U18049 (N_18049,N_14948,N_12700);
xor U18050 (N_18050,N_14427,N_12579);
or U18051 (N_18051,N_12290,N_13516);
and U18052 (N_18052,N_13428,N_15924);
or U18053 (N_18053,N_12833,N_15621);
xnor U18054 (N_18054,N_12943,N_15936);
and U18055 (N_18055,N_12159,N_13476);
xor U18056 (N_18056,N_14412,N_15921);
nand U18057 (N_18057,N_14135,N_15146);
xor U18058 (N_18058,N_13659,N_13068);
nor U18059 (N_18059,N_12375,N_13418);
nand U18060 (N_18060,N_15245,N_13465);
nand U18061 (N_18061,N_14757,N_13640);
or U18062 (N_18062,N_13281,N_13927);
and U18063 (N_18063,N_12148,N_13864);
nor U18064 (N_18064,N_14226,N_15760);
nand U18065 (N_18065,N_12460,N_14479);
and U18066 (N_18066,N_13745,N_15129);
nand U18067 (N_18067,N_15757,N_15929);
xor U18068 (N_18068,N_15512,N_15596);
xor U18069 (N_18069,N_12129,N_14714);
and U18070 (N_18070,N_14246,N_14092);
nor U18071 (N_18071,N_12363,N_13475);
nor U18072 (N_18072,N_13913,N_15136);
nand U18073 (N_18073,N_14176,N_12103);
nand U18074 (N_18074,N_15233,N_15158);
nand U18075 (N_18075,N_13756,N_14754);
nor U18076 (N_18076,N_12253,N_12502);
and U18077 (N_18077,N_13497,N_15538);
nand U18078 (N_18078,N_12338,N_13066);
nand U18079 (N_18079,N_14954,N_13534);
nor U18080 (N_18080,N_12979,N_13639);
nor U18081 (N_18081,N_12313,N_13671);
and U18082 (N_18082,N_14369,N_14758);
and U18083 (N_18083,N_15470,N_15518);
or U18084 (N_18084,N_13237,N_15144);
nand U18085 (N_18085,N_14249,N_14492);
nand U18086 (N_18086,N_13142,N_14592);
nor U18087 (N_18087,N_15550,N_13551);
nand U18088 (N_18088,N_13469,N_13522);
and U18089 (N_18089,N_15116,N_12533);
or U18090 (N_18090,N_13801,N_12413);
or U18091 (N_18091,N_12368,N_15521);
xor U18092 (N_18092,N_13185,N_13324);
and U18093 (N_18093,N_13036,N_13623);
xnor U18094 (N_18094,N_14814,N_13864);
xor U18095 (N_18095,N_15176,N_13123);
and U18096 (N_18096,N_14312,N_14870);
nand U18097 (N_18097,N_14426,N_14268);
nand U18098 (N_18098,N_13486,N_13678);
nor U18099 (N_18099,N_14222,N_13060);
xnor U18100 (N_18100,N_15288,N_15576);
xnor U18101 (N_18101,N_12821,N_15295);
nand U18102 (N_18102,N_14613,N_15650);
nor U18103 (N_18103,N_15226,N_14366);
nor U18104 (N_18104,N_12409,N_15141);
and U18105 (N_18105,N_14127,N_14519);
or U18106 (N_18106,N_14560,N_12304);
and U18107 (N_18107,N_12606,N_13003);
nor U18108 (N_18108,N_14521,N_12052);
nand U18109 (N_18109,N_14618,N_12693);
nor U18110 (N_18110,N_13180,N_12028);
nand U18111 (N_18111,N_12391,N_14395);
nor U18112 (N_18112,N_12911,N_15263);
nand U18113 (N_18113,N_12016,N_12777);
nor U18114 (N_18114,N_13451,N_13245);
nor U18115 (N_18115,N_12786,N_12054);
or U18116 (N_18116,N_14501,N_13169);
xnor U18117 (N_18117,N_14634,N_14420);
and U18118 (N_18118,N_13408,N_15314);
nor U18119 (N_18119,N_12688,N_12859);
or U18120 (N_18120,N_12044,N_14488);
nor U18121 (N_18121,N_12935,N_13617);
nand U18122 (N_18122,N_15896,N_15145);
and U18123 (N_18123,N_15412,N_12763);
and U18124 (N_18124,N_15243,N_13467);
nand U18125 (N_18125,N_14721,N_15565);
and U18126 (N_18126,N_15597,N_15587);
or U18127 (N_18127,N_13594,N_14427);
or U18128 (N_18128,N_15230,N_12151);
and U18129 (N_18129,N_15365,N_14243);
or U18130 (N_18130,N_12209,N_15529);
nor U18131 (N_18131,N_12407,N_13075);
and U18132 (N_18132,N_14910,N_14723);
nor U18133 (N_18133,N_13993,N_14650);
or U18134 (N_18134,N_13102,N_13284);
nor U18135 (N_18135,N_12434,N_14478);
and U18136 (N_18136,N_14608,N_13710);
nor U18137 (N_18137,N_12942,N_12333);
nand U18138 (N_18138,N_14928,N_14634);
xor U18139 (N_18139,N_12175,N_14064);
or U18140 (N_18140,N_14861,N_13165);
and U18141 (N_18141,N_14189,N_13809);
nor U18142 (N_18142,N_13388,N_14958);
xnor U18143 (N_18143,N_13052,N_13254);
or U18144 (N_18144,N_13546,N_14016);
nand U18145 (N_18145,N_15107,N_12351);
nor U18146 (N_18146,N_12041,N_13186);
nand U18147 (N_18147,N_14528,N_14854);
nand U18148 (N_18148,N_14184,N_13239);
or U18149 (N_18149,N_13920,N_15019);
and U18150 (N_18150,N_12979,N_14271);
nand U18151 (N_18151,N_14821,N_13250);
nand U18152 (N_18152,N_12328,N_13653);
nand U18153 (N_18153,N_14323,N_13325);
nand U18154 (N_18154,N_13553,N_12773);
xnor U18155 (N_18155,N_13648,N_14679);
nand U18156 (N_18156,N_12750,N_13679);
xor U18157 (N_18157,N_13385,N_15540);
xnor U18158 (N_18158,N_13300,N_13008);
or U18159 (N_18159,N_15768,N_14579);
nand U18160 (N_18160,N_15093,N_13627);
xor U18161 (N_18161,N_15962,N_14019);
xnor U18162 (N_18162,N_13756,N_15783);
nand U18163 (N_18163,N_12521,N_14491);
or U18164 (N_18164,N_14130,N_14067);
or U18165 (N_18165,N_14224,N_15606);
and U18166 (N_18166,N_14682,N_12005);
or U18167 (N_18167,N_14808,N_15920);
and U18168 (N_18168,N_12620,N_15699);
xor U18169 (N_18169,N_12268,N_14548);
nand U18170 (N_18170,N_15531,N_13214);
xor U18171 (N_18171,N_15521,N_15192);
nor U18172 (N_18172,N_14123,N_12062);
xnor U18173 (N_18173,N_12166,N_15037);
nor U18174 (N_18174,N_14655,N_14942);
nor U18175 (N_18175,N_14511,N_15412);
nor U18176 (N_18176,N_13759,N_15126);
nor U18177 (N_18177,N_13376,N_15831);
and U18178 (N_18178,N_15934,N_13699);
nand U18179 (N_18179,N_15196,N_14009);
nand U18180 (N_18180,N_15210,N_12284);
nor U18181 (N_18181,N_14480,N_15958);
and U18182 (N_18182,N_15002,N_13362);
xor U18183 (N_18183,N_13489,N_13734);
xor U18184 (N_18184,N_12325,N_12040);
nand U18185 (N_18185,N_12947,N_13261);
nor U18186 (N_18186,N_12916,N_13633);
and U18187 (N_18187,N_12571,N_12363);
nand U18188 (N_18188,N_13350,N_14644);
nor U18189 (N_18189,N_14876,N_13196);
nor U18190 (N_18190,N_15792,N_12153);
xor U18191 (N_18191,N_12891,N_12985);
nand U18192 (N_18192,N_14407,N_15397);
or U18193 (N_18193,N_13014,N_15457);
nor U18194 (N_18194,N_12891,N_15660);
xnor U18195 (N_18195,N_14378,N_15936);
nand U18196 (N_18196,N_15511,N_14734);
xnor U18197 (N_18197,N_12951,N_15273);
nand U18198 (N_18198,N_13617,N_13056);
or U18199 (N_18199,N_13841,N_13298);
xor U18200 (N_18200,N_13443,N_13008);
nor U18201 (N_18201,N_12374,N_12130);
nor U18202 (N_18202,N_12002,N_12397);
and U18203 (N_18203,N_15175,N_15367);
xor U18204 (N_18204,N_15831,N_12830);
xor U18205 (N_18205,N_13155,N_13477);
nand U18206 (N_18206,N_12634,N_12701);
or U18207 (N_18207,N_14978,N_15985);
xor U18208 (N_18208,N_15307,N_12136);
xnor U18209 (N_18209,N_13546,N_12776);
or U18210 (N_18210,N_12867,N_15691);
nor U18211 (N_18211,N_12807,N_15563);
nor U18212 (N_18212,N_13773,N_14337);
nor U18213 (N_18213,N_13882,N_12118);
nand U18214 (N_18214,N_13579,N_12350);
xor U18215 (N_18215,N_14012,N_15686);
nor U18216 (N_18216,N_12002,N_14904);
xor U18217 (N_18217,N_13019,N_14736);
or U18218 (N_18218,N_14630,N_15063);
or U18219 (N_18219,N_13455,N_14206);
xor U18220 (N_18220,N_13600,N_12618);
or U18221 (N_18221,N_13983,N_14434);
or U18222 (N_18222,N_13508,N_14212);
xor U18223 (N_18223,N_12981,N_13606);
nor U18224 (N_18224,N_12720,N_13676);
or U18225 (N_18225,N_15122,N_15081);
nor U18226 (N_18226,N_14932,N_15043);
nor U18227 (N_18227,N_13098,N_13764);
or U18228 (N_18228,N_15843,N_14257);
or U18229 (N_18229,N_14685,N_15079);
nor U18230 (N_18230,N_14612,N_15935);
or U18231 (N_18231,N_14567,N_14982);
and U18232 (N_18232,N_12878,N_13611);
nor U18233 (N_18233,N_14312,N_15309);
nor U18234 (N_18234,N_14710,N_15440);
xnor U18235 (N_18235,N_12415,N_15770);
nor U18236 (N_18236,N_15019,N_14575);
and U18237 (N_18237,N_15877,N_15096);
nor U18238 (N_18238,N_13263,N_12092);
and U18239 (N_18239,N_13656,N_13660);
nand U18240 (N_18240,N_14676,N_15545);
nor U18241 (N_18241,N_13524,N_15339);
xnor U18242 (N_18242,N_15721,N_14954);
or U18243 (N_18243,N_14147,N_13485);
and U18244 (N_18244,N_12776,N_14885);
or U18245 (N_18245,N_14581,N_15070);
xnor U18246 (N_18246,N_15839,N_15253);
and U18247 (N_18247,N_13846,N_15643);
nand U18248 (N_18248,N_14519,N_12578);
and U18249 (N_18249,N_12865,N_15657);
xor U18250 (N_18250,N_13121,N_13397);
nand U18251 (N_18251,N_13952,N_13877);
and U18252 (N_18252,N_13326,N_14777);
or U18253 (N_18253,N_14055,N_15765);
and U18254 (N_18254,N_14867,N_13933);
nand U18255 (N_18255,N_14914,N_12587);
and U18256 (N_18256,N_13889,N_12592);
and U18257 (N_18257,N_13475,N_14210);
nor U18258 (N_18258,N_15963,N_14415);
or U18259 (N_18259,N_14234,N_15363);
nand U18260 (N_18260,N_13557,N_12206);
xor U18261 (N_18261,N_13066,N_15050);
and U18262 (N_18262,N_13832,N_14467);
nor U18263 (N_18263,N_14714,N_14481);
xor U18264 (N_18264,N_14493,N_14123);
or U18265 (N_18265,N_12059,N_15156);
and U18266 (N_18266,N_15917,N_13691);
nor U18267 (N_18267,N_14321,N_14466);
and U18268 (N_18268,N_15505,N_13485);
xor U18269 (N_18269,N_13114,N_12368);
xor U18270 (N_18270,N_12583,N_14587);
nand U18271 (N_18271,N_14720,N_13858);
or U18272 (N_18272,N_15715,N_13089);
xor U18273 (N_18273,N_12985,N_12526);
or U18274 (N_18274,N_13525,N_13214);
xnor U18275 (N_18275,N_13238,N_14716);
or U18276 (N_18276,N_12173,N_13923);
nor U18277 (N_18277,N_14541,N_12550);
or U18278 (N_18278,N_15348,N_12793);
or U18279 (N_18279,N_13249,N_15124);
nor U18280 (N_18280,N_14328,N_14720);
and U18281 (N_18281,N_15021,N_15109);
nor U18282 (N_18282,N_15028,N_15183);
nor U18283 (N_18283,N_13643,N_12211);
nor U18284 (N_18284,N_12283,N_14969);
nor U18285 (N_18285,N_12856,N_13672);
nand U18286 (N_18286,N_13574,N_12448);
nor U18287 (N_18287,N_15377,N_13064);
nand U18288 (N_18288,N_14315,N_14660);
and U18289 (N_18289,N_14447,N_13190);
nand U18290 (N_18290,N_14590,N_13374);
or U18291 (N_18291,N_15319,N_15199);
nor U18292 (N_18292,N_15625,N_15171);
nor U18293 (N_18293,N_15460,N_13286);
xor U18294 (N_18294,N_15106,N_14296);
nand U18295 (N_18295,N_12460,N_13409);
xnor U18296 (N_18296,N_12869,N_13347);
or U18297 (N_18297,N_12794,N_13738);
nand U18298 (N_18298,N_13572,N_14462);
xor U18299 (N_18299,N_13073,N_12700);
nor U18300 (N_18300,N_14638,N_12196);
xnor U18301 (N_18301,N_12184,N_12327);
and U18302 (N_18302,N_12080,N_13760);
nor U18303 (N_18303,N_12743,N_13462);
or U18304 (N_18304,N_14254,N_13451);
or U18305 (N_18305,N_15173,N_13859);
or U18306 (N_18306,N_14047,N_15568);
nor U18307 (N_18307,N_12423,N_15919);
nor U18308 (N_18308,N_13199,N_12057);
or U18309 (N_18309,N_15770,N_13193);
or U18310 (N_18310,N_14373,N_14968);
nand U18311 (N_18311,N_15526,N_15812);
or U18312 (N_18312,N_12098,N_12093);
nand U18313 (N_18313,N_12059,N_15029);
nand U18314 (N_18314,N_12847,N_14350);
nand U18315 (N_18315,N_13809,N_13664);
and U18316 (N_18316,N_12441,N_12591);
or U18317 (N_18317,N_12536,N_13937);
xor U18318 (N_18318,N_13735,N_12120);
nor U18319 (N_18319,N_14132,N_13896);
or U18320 (N_18320,N_15731,N_14555);
nand U18321 (N_18321,N_14863,N_15055);
or U18322 (N_18322,N_13410,N_14969);
nand U18323 (N_18323,N_13938,N_12565);
xnor U18324 (N_18324,N_13026,N_13241);
xor U18325 (N_18325,N_12349,N_13035);
nor U18326 (N_18326,N_12719,N_12156);
xor U18327 (N_18327,N_15980,N_13025);
or U18328 (N_18328,N_12608,N_15105);
xnor U18329 (N_18329,N_15507,N_15349);
nand U18330 (N_18330,N_12597,N_14224);
and U18331 (N_18331,N_14622,N_15196);
xnor U18332 (N_18332,N_12171,N_13883);
and U18333 (N_18333,N_12715,N_13954);
nor U18334 (N_18334,N_12600,N_12166);
or U18335 (N_18335,N_13569,N_15449);
and U18336 (N_18336,N_12167,N_14371);
and U18337 (N_18337,N_15096,N_15746);
nand U18338 (N_18338,N_13870,N_12467);
nor U18339 (N_18339,N_15583,N_14493);
xor U18340 (N_18340,N_15889,N_12652);
nand U18341 (N_18341,N_15937,N_14052);
xnor U18342 (N_18342,N_12882,N_15141);
or U18343 (N_18343,N_14131,N_14576);
and U18344 (N_18344,N_12927,N_14999);
and U18345 (N_18345,N_12361,N_14021);
nor U18346 (N_18346,N_12327,N_13706);
and U18347 (N_18347,N_14117,N_15135);
xnor U18348 (N_18348,N_14328,N_14999);
or U18349 (N_18349,N_13434,N_14625);
nor U18350 (N_18350,N_14362,N_14201);
nor U18351 (N_18351,N_14992,N_13902);
or U18352 (N_18352,N_13920,N_13799);
or U18353 (N_18353,N_13778,N_13275);
nor U18354 (N_18354,N_14883,N_14749);
or U18355 (N_18355,N_15253,N_14461);
nor U18356 (N_18356,N_15228,N_15580);
or U18357 (N_18357,N_13113,N_15027);
xnor U18358 (N_18358,N_12784,N_14770);
and U18359 (N_18359,N_13523,N_13516);
nor U18360 (N_18360,N_15257,N_15825);
and U18361 (N_18361,N_13274,N_12747);
and U18362 (N_18362,N_15635,N_12341);
xnor U18363 (N_18363,N_13766,N_15423);
xnor U18364 (N_18364,N_13021,N_14573);
and U18365 (N_18365,N_15964,N_14023);
nor U18366 (N_18366,N_14912,N_12577);
and U18367 (N_18367,N_15763,N_15173);
xnor U18368 (N_18368,N_12230,N_12030);
nand U18369 (N_18369,N_13642,N_12696);
xor U18370 (N_18370,N_15822,N_12281);
nor U18371 (N_18371,N_12878,N_15964);
or U18372 (N_18372,N_13898,N_12325);
xnor U18373 (N_18373,N_12013,N_13667);
nand U18374 (N_18374,N_14751,N_13270);
nand U18375 (N_18375,N_13873,N_14613);
nand U18376 (N_18376,N_15775,N_15011);
nor U18377 (N_18377,N_15759,N_12885);
nand U18378 (N_18378,N_14376,N_12075);
and U18379 (N_18379,N_14475,N_14954);
nand U18380 (N_18380,N_15727,N_15081);
or U18381 (N_18381,N_14322,N_12629);
nor U18382 (N_18382,N_13644,N_12766);
and U18383 (N_18383,N_15111,N_13574);
nor U18384 (N_18384,N_13657,N_15542);
nor U18385 (N_18385,N_12524,N_13247);
nor U18386 (N_18386,N_14136,N_12004);
xor U18387 (N_18387,N_12940,N_15555);
xnor U18388 (N_18388,N_13528,N_12988);
and U18389 (N_18389,N_13031,N_14700);
or U18390 (N_18390,N_15626,N_13166);
or U18391 (N_18391,N_13208,N_14271);
or U18392 (N_18392,N_15420,N_15897);
xor U18393 (N_18393,N_14311,N_15131);
xor U18394 (N_18394,N_15044,N_14505);
nand U18395 (N_18395,N_13769,N_13211);
nor U18396 (N_18396,N_12568,N_14040);
xor U18397 (N_18397,N_14368,N_13611);
nor U18398 (N_18398,N_12665,N_14029);
and U18399 (N_18399,N_15010,N_15817);
nor U18400 (N_18400,N_12542,N_15813);
nand U18401 (N_18401,N_15718,N_14714);
nand U18402 (N_18402,N_12970,N_12540);
nand U18403 (N_18403,N_14830,N_14123);
or U18404 (N_18404,N_12424,N_14401);
nor U18405 (N_18405,N_15896,N_15039);
and U18406 (N_18406,N_14775,N_14144);
xor U18407 (N_18407,N_14728,N_15759);
nand U18408 (N_18408,N_15016,N_14187);
and U18409 (N_18409,N_13254,N_12701);
or U18410 (N_18410,N_13300,N_12635);
nand U18411 (N_18411,N_12965,N_15509);
and U18412 (N_18412,N_13919,N_13072);
xnor U18413 (N_18413,N_12555,N_12624);
nand U18414 (N_18414,N_15240,N_13206);
or U18415 (N_18415,N_13503,N_15699);
nor U18416 (N_18416,N_12634,N_13549);
nand U18417 (N_18417,N_13100,N_12475);
or U18418 (N_18418,N_15257,N_12443);
or U18419 (N_18419,N_15794,N_12265);
or U18420 (N_18420,N_14847,N_13959);
or U18421 (N_18421,N_13299,N_14197);
and U18422 (N_18422,N_14453,N_12838);
nor U18423 (N_18423,N_15476,N_12670);
and U18424 (N_18424,N_14912,N_12839);
or U18425 (N_18425,N_15714,N_15605);
nor U18426 (N_18426,N_13346,N_12288);
nor U18427 (N_18427,N_15898,N_12348);
nand U18428 (N_18428,N_15891,N_13744);
and U18429 (N_18429,N_14576,N_14479);
nand U18430 (N_18430,N_13526,N_13107);
and U18431 (N_18431,N_13653,N_12504);
nand U18432 (N_18432,N_12935,N_12509);
nand U18433 (N_18433,N_14163,N_14019);
and U18434 (N_18434,N_12587,N_13789);
and U18435 (N_18435,N_15182,N_15335);
xnor U18436 (N_18436,N_13735,N_13344);
or U18437 (N_18437,N_13912,N_13035);
nor U18438 (N_18438,N_14560,N_12552);
nand U18439 (N_18439,N_14138,N_13108);
nor U18440 (N_18440,N_12662,N_15862);
nor U18441 (N_18441,N_12060,N_12058);
and U18442 (N_18442,N_13050,N_13953);
xnor U18443 (N_18443,N_13427,N_12314);
nor U18444 (N_18444,N_12341,N_13882);
and U18445 (N_18445,N_14485,N_14903);
xnor U18446 (N_18446,N_15211,N_12585);
xor U18447 (N_18447,N_13954,N_12049);
or U18448 (N_18448,N_12860,N_15959);
or U18449 (N_18449,N_12774,N_13557);
xnor U18450 (N_18450,N_12393,N_15635);
or U18451 (N_18451,N_15587,N_15900);
xnor U18452 (N_18452,N_15548,N_14709);
or U18453 (N_18453,N_13968,N_15040);
nor U18454 (N_18454,N_15233,N_13732);
nor U18455 (N_18455,N_13557,N_15437);
xnor U18456 (N_18456,N_13083,N_14854);
nor U18457 (N_18457,N_15140,N_13997);
or U18458 (N_18458,N_14136,N_15364);
or U18459 (N_18459,N_14573,N_12644);
and U18460 (N_18460,N_14102,N_13815);
xor U18461 (N_18461,N_12390,N_15922);
nand U18462 (N_18462,N_12649,N_12791);
nand U18463 (N_18463,N_15707,N_12303);
nand U18464 (N_18464,N_14500,N_13821);
and U18465 (N_18465,N_13493,N_12354);
nand U18466 (N_18466,N_13192,N_14601);
xor U18467 (N_18467,N_13046,N_13415);
and U18468 (N_18468,N_15842,N_12592);
and U18469 (N_18469,N_13128,N_14275);
or U18470 (N_18470,N_13824,N_15223);
and U18471 (N_18471,N_12662,N_13091);
or U18472 (N_18472,N_12088,N_14090);
or U18473 (N_18473,N_15793,N_12555);
nor U18474 (N_18474,N_14535,N_13058);
nand U18475 (N_18475,N_14006,N_12763);
xor U18476 (N_18476,N_13431,N_15397);
nand U18477 (N_18477,N_12005,N_15197);
and U18478 (N_18478,N_13442,N_12140);
nand U18479 (N_18479,N_14576,N_13646);
xor U18480 (N_18480,N_12597,N_14000);
or U18481 (N_18481,N_12054,N_15803);
xnor U18482 (N_18482,N_14720,N_12409);
nor U18483 (N_18483,N_15707,N_12345);
and U18484 (N_18484,N_14583,N_13172);
nand U18485 (N_18485,N_13850,N_13099);
nor U18486 (N_18486,N_15453,N_15927);
and U18487 (N_18487,N_15241,N_14138);
or U18488 (N_18488,N_12028,N_14004);
nand U18489 (N_18489,N_13335,N_12400);
and U18490 (N_18490,N_14403,N_15085);
nand U18491 (N_18491,N_15075,N_15008);
nand U18492 (N_18492,N_13833,N_14930);
nand U18493 (N_18493,N_15948,N_12298);
nor U18494 (N_18494,N_13469,N_15709);
or U18495 (N_18495,N_15894,N_14014);
nand U18496 (N_18496,N_15634,N_13807);
and U18497 (N_18497,N_12952,N_12271);
nor U18498 (N_18498,N_14777,N_13383);
xnor U18499 (N_18499,N_14572,N_12412);
nand U18500 (N_18500,N_12438,N_12825);
nor U18501 (N_18501,N_12694,N_13096);
nor U18502 (N_18502,N_15207,N_13451);
nand U18503 (N_18503,N_15364,N_15343);
and U18504 (N_18504,N_12565,N_15603);
and U18505 (N_18505,N_12994,N_15421);
and U18506 (N_18506,N_13825,N_13661);
nor U18507 (N_18507,N_12560,N_14948);
nand U18508 (N_18508,N_13499,N_14547);
and U18509 (N_18509,N_12102,N_13664);
nand U18510 (N_18510,N_13463,N_15417);
and U18511 (N_18511,N_15202,N_15464);
or U18512 (N_18512,N_15193,N_14204);
nor U18513 (N_18513,N_12971,N_15534);
nor U18514 (N_18514,N_12294,N_15161);
nor U18515 (N_18515,N_12346,N_14443);
xor U18516 (N_18516,N_14995,N_14765);
nor U18517 (N_18517,N_15062,N_14958);
nor U18518 (N_18518,N_12850,N_13477);
xnor U18519 (N_18519,N_14429,N_13969);
nand U18520 (N_18520,N_14421,N_13278);
xor U18521 (N_18521,N_15685,N_12988);
and U18522 (N_18522,N_13901,N_13776);
nor U18523 (N_18523,N_14502,N_15108);
or U18524 (N_18524,N_13751,N_14066);
nor U18525 (N_18525,N_13484,N_12757);
xnor U18526 (N_18526,N_14676,N_13485);
nor U18527 (N_18527,N_12387,N_14921);
nand U18528 (N_18528,N_15440,N_12980);
nor U18529 (N_18529,N_12746,N_15866);
nor U18530 (N_18530,N_14054,N_13674);
and U18531 (N_18531,N_15343,N_12572);
xnor U18532 (N_18532,N_15233,N_14934);
or U18533 (N_18533,N_14843,N_14093);
xnor U18534 (N_18534,N_15109,N_14766);
or U18535 (N_18535,N_13084,N_14047);
xnor U18536 (N_18536,N_13005,N_12796);
nand U18537 (N_18537,N_14215,N_15826);
nand U18538 (N_18538,N_14800,N_15082);
nand U18539 (N_18539,N_15827,N_12549);
xnor U18540 (N_18540,N_14734,N_14703);
nor U18541 (N_18541,N_15880,N_15017);
or U18542 (N_18542,N_14147,N_15065);
or U18543 (N_18543,N_12614,N_13169);
xor U18544 (N_18544,N_12433,N_14257);
nor U18545 (N_18545,N_13810,N_15356);
or U18546 (N_18546,N_13658,N_14836);
nor U18547 (N_18547,N_14447,N_14388);
xnor U18548 (N_18548,N_13634,N_15514);
nor U18549 (N_18549,N_12928,N_13511);
and U18550 (N_18550,N_14823,N_12001);
or U18551 (N_18551,N_13360,N_12243);
xnor U18552 (N_18552,N_15106,N_14222);
xor U18553 (N_18553,N_14864,N_15732);
or U18554 (N_18554,N_14206,N_14762);
nand U18555 (N_18555,N_13682,N_13393);
and U18556 (N_18556,N_14553,N_15509);
and U18557 (N_18557,N_13876,N_13978);
xnor U18558 (N_18558,N_15995,N_13025);
or U18559 (N_18559,N_15668,N_14052);
nor U18560 (N_18560,N_15913,N_12768);
nor U18561 (N_18561,N_13116,N_14493);
nor U18562 (N_18562,N_13833,N_12694);
xnor U18563 (N_18563,N_12824,N_15655);
and U18564 (N_18564,N_14999,N_12353);
or U18565 (N_18565,N_13243,N_13950);
nor U18566 (N_18566,N_15521,N_13638);
xor U18567 (N_18567,N_14157,N_12023);
or U18568 (N_18568,N_15535,N_12484);
nand U18569 (N_18569,N_12133,N_12147);
or U18570 (N_18570,N_13944,N_15543);
nand U18571 (N_18571,N_15308,N_14853);
and U18572 (N_18572,N_14182,N_13246);
nor U18573 (N_18573,N_14786,N_14498);
or U18574 (N_18574,N_14738,N_14044);
nand U18575 (N_18575,N_15434,N_12111);
nor U18576 (N_18576,N_12194,N_12389);
xor U18577 (N_18577,N_15536,N_12794);
xor U18578 (N_18578,N_13443,N_12939);
xor U18579 (N_18579,N_12759,N_13121);
and U18580 (N_18580,N_13143,N_15814);
or U18581 (N_18581,N_12436,N_12890);
or U18582 (N_18582,N_15083,N_13488);
xor U18583 (N_18583,N_12259,N_14335);
or U18584 (N_18584,N_15123,N_15518);
xor U18585 (N_18585,N_12808,N_15740);
nand U18586 (N_18586,N_12919,N_13764);
xnor U18587 (N_18587,N_15622,N_15652);
nand U18588 (N_18588,N_12178,N_15098);
or U18589 (N_18589,N_12758,N_13357);
or U18590 (N_18590,N_13552,N_14986);
nand U18591 (N_18591,N_15212,N_12445);
nor U18592 (N_18592,N_13726,N_12878);
nor U18593 (N_18593,N_14610,N_14894);
xnor U18594 (N_18594,N_13645,N_14594);
xor U18595 (N_18595,N_14057,N_15688);
and U18596 (N_18596,N_15488,N_13853);
or U18597 (N_18597,N_14888,N_12196);
nand U18598 (N_18598,N_12167,N_14191);
nand U18599 (N_18599,N_14896,N_13406);
xnor U18600 (N_18600,N_12671,N_14004);
or U18601 (N_18601,N_13084,N_13443);
and U18602 (N_18602,N_12938,N_12422);
nand U18603 (N_18603,N_14468,N_14104);
nor U18604 (N_18604,N_14430,N_15689);
nor U18605 (N_18605,N_14997,N_12843);
or U18606 (N_18606,N_15120,N_15250);
or U18607 (N_18607,N_14414,N_15731);
nor U18608 (N_18608,N_12432,N_14639);
nor U18609 (N_18609,N_14706,N_13304);
or U18610 (N_18610,N_12574,N_13824);
nor U18611 (N_18611,N_13538,N_15815);
xnor U18612 (N_18612,N_13977,N_14555);
nand U18613 (N_18613,N_12471,N_12951);
nand U18614 (N_18614,N_15950,N_14465);
nand U18615 (N_18615,N_12446,N_13162);
nor U18616 (N_18616,N_12702,N_13987);
nand U18617 (N_18617,N_14242,N_14209);
nand U18618 (N_18618,N_13561,N_12709);
and U18619 (N_18619,N_12340,N_15984);
nor U18620 (N_18620,N_15468,N_13429);
and U18621 (N_18621,N_14535,N_12742);
and U18622 (N_18622,N_13213,N_15853);
xor U18623 (N_18623,N_14145,N_14682);
nand U18624 (N_18624,N_14133,N_15072);
xnor U18625 (N_18625,N_14989,N_14284);
xor U18626 (N_18626,N_13873,N_14455);
and U18627 (N_18627,N_12004,N_12162);
and U18628 (N_18628,N_15897,N_15138);
nand U18629 (N_18629,N_12341,N_12776);
nor U18630 (N_18630,N_13898,N_13548);
nor U18631 (N_18631,N_14711,N_14392);
nor U18632 (N_18632,N_15307,N_13293);
xnor U18633 (N_18633,N_12125,N_12232);
or U18634 (N_18634,N_15006,N_14398);
xnor U18635 (N_18635,N_12587,N_15808);
or U18636 (N_18636,N_12980,N_12971);
or U18637 (N_18637,N_15438,N_14774);
nor U18638 (N_18638,N_13393,N_12989);
nor U18639 (N_18639,N_12684,N_13877);
or U18640 (N_18640,N_13204,N_12649);
and U18641 (N_18641,N_12969,N_15315);
nand U18642 (N_18642,N_13152,N_15324);
nand U18643 (N_18643,N_14617,N_14481);
xnor U18644 (N_18644,N_13307,N_15491);
xor U18645 (N_18645,N_12769,N_12154);
xor U18646 (N_18646,N_15313,N_13523);
nor U18647 (N_18647,N_12211,N_13903);
or U18648 (N_18648,N_13506,N_15973);
or U18649 (N_18649,N_15276,N_15941);
or U18650 (N_18650,N_12297,N_12834);
and U18651 (N_18651,N_13941,N_15523);
nor U18652 (N_18652,N_14626,N_15261);
nand U18653 (N_18653,N_13355,N_15132);
or U18654 (N_18654,N_15030,N_12253);
or U18655 (N_18655,N_15886,N_15240);
or U18656 (N_18656,N_14536,N_13735);
or U18657 (N_18657,N_12115,N_13763);
or U18658 (N_18658,N_12361,N_12722);
nor U18659 (N_18659,N_12747,N_15742);
xor U18660 (N_18660,N_12804,N_12901);
and U18661 (N_18661,N_13822,N_12508);
nand U18662 (N_18662,N_13801,N_15336);
nor U18663 (N_18663,N_15019,N_12966);
xor U18664 (N_18664,N_15503,N_15218);
or U18665 (N_18665,N_12658,N_15086);
nand U18666 (N_18666,N_13289,N_13612);
and U18667 (N_18667,N_13106,N_13600);
nor U18668 (N_18668,N_15807,N_13927);
or U18669 (N_18669,N_12695,N_12860);
nand U18670 (N_18670,N_12915,N_14520);
and U18671 (N_18671,N_12879,N_13384);
nor U18672 (N_18672,N_14566,N_15519);
nand U18673 (N_18673,N_15449,N_12935);
nand U18674 (N_18674,N_13225,N_13147);
xor U18675 (N_18675,N_14148,N_13209);
nand U18676 (N_18676,N_15318,N_14274);
nand U18677 (N_18677,N_12172,N_13023);
xor U18678 (N_18678,N_13726,N_14038);
xor U18679 (N_18679,N_13527,N_15283);
and U18680 (N_18680,N_15586,N_15422);
nand U18681 (N_18681,N_13138,N_12998);
xnor U18682 (N_18682,N_15634,N_15895);
xor U18683 (N_18683,N_12032,N_15596);
nor U18684 (N_18684,N_13640,N_13155);
nor U18685 (N_18685,N_15405,N_13894);
nor U18686 (N_18686,N_14250,N_12758);
xor U18687 (N_18687,N_14620,N_13104);
nand U18688 (N_18688,N_14912,N_12791);
nand U18689 (N_18689,N_15724,N_12390);
and U18690 (N_18690,N_14971,N_15278);
nor U18691 (N_18691,N_15484,N_13418);
and U18692 (N_18692,N_12515,N_12460);
nand U18693 (N_18693,N_12736,N_15578);
nand U18694 (N_18694,N_12355,N_12576);
and U18695 (N_18695,N_15997,N_14681);
nand U18696 (N_18696,N_14654,N_14126);
or U18697 (N_18697,N_14632,N_12146);
nor U18698 (N_18698,N_15482,N_15389);
or U18699 (N_18699,N_13585,N_15106);
or U18700 (N_18700,N_15787,N_15626);
or U18701 (N_18701,N_13744,N_15356);
nand U18702 (N_18702,N_13803,N_13587);
nand U18703 (N_18703,N_13167,N_12345);
xnor U18704 (N_18704,N_14525,N_15325);
nor U18705 (N_18705,N_13542,N_13521);
and U18706 (N_18706,N_12491,N_14201);
or U18707 (N_18707,N_14432,N_14861);
nor U18708 (N_18708,N_13853,N_13823);
nand U18709 (N_18709,N_12458,N_12625);
and U18710 (N_18710,N_15555,N_15147);
or U18711 (N_18711,N_14888,N_13489);
or U18712 (N_18712,N_13178,N_13006);
xor U18713 (N_18713,N_14118,N_13814);
nor U18714 (N_18714,N_12458,N_14884);
nand U18715 (N_18715,N_14616,N_12294);
and U18716 (N_18716,N_15703,N_15442);
and U18717 (N_18717,N_12879,N_15193);
nor U18718 (N_18718,N_14948,N_14877);
nor U18719 (N_18719,N_12072,N_15912);
or U18720 (N_18720,N_12459,N_13944);
and U18721 (N_18721,N_15034,N_13423);
xnor U18722 (N_18722,N_14306,N_14292);
nor U18723 (N_18723,N_15632,N_14126);
nor U18724 (N_18724,N_14525,N_13693);
or U18725 (N_18725,N_15340,N_15674);
xor U18726 (N_18726,N_15555,N_14146);
xnor U18727 (N_18727,N_13002,N_15441);
and U18728 (N_18728,N_14263,N_13986);
nor U18729 (N_18729,N_14914,N_15938);
nor U18730 (N_18730,N_13157,N_12749);
or U18731 (N_18731,N_14371,N_12364);
or U18732 (N_18732,N_12748,N_15787);
and U18733 (N_18733,N_13242,N_15025);
nor U18734 (N_18734,N_12430,N_13560);
or U18735 (N_18735,N_13900,N_14199);
nand U18736 (N_18736,N_14710,N_15088);
and U18737 (N_18737,N_12787,N_13142);
and U18738 (N_18738,N_13868,N_15721);
and U18739 (N_18739,N_13126,N_15352);
and U18740 (N_18740,N_13507,N_15543);
nor U18741 (N_18741,N_14740,N_14767);
nand U18742 (N_18742,N_14189,N_14051);
nor U18743 (N_18743,N_12329,N_15934);
xor U18744 (N_18744,N_13547,N_13749);
nand U18745 (N_18745,N_14862,N_14868);
nor U18746 (N_18746,N_13836,N_15797);
and U18747 (N_18747,N_14172,N_14627);
and U18748 (N_18748,N_14976,N_14071);
or U18749 (N_18749,N_12327,N_12896);
or U18750 (N_18750,N_13890,N_12742);
nand U18751 (N_18751,N_12900,N_14955);
and U18752 (N_18752,N_13079,N_14242);
nand U18753 (N_18753,N_15797,N_12468);
nor U18754 (N_18754,N_13878,N_12900);
nor U18755 (N_18755,N_12866,N_15168);
xor U18756 (N_18756,N_12154,N_15814);
nor U18757 (N_18757,N_15652,N_12285);
xor U18758 (N_18758,N_12003,N_14440);
nor U18759 (N_18759,N_15705,N_13206);
nand U18760 (N_18760,N_14403,N_15010);
nand U18761 (N_18761,N_12835,N_14645);
or U18762 (N_18762,N_14144,N_13065);
xnor U18763 (N_18763,N_13982,N_15710);
xnor U18764 (N_18764,N_14677,N_15398);
nor U18765 (N_18765,N_14186,N_15829);
nor U18766 (N_18766,N_14392,N_12372);
xor U18767 (N_18767,N_13831,N_12013);
nor U18768 (N_18768,N_14090,N_13341);
xnor U18769 (N_18769,N_15687,N_12279);
or U18770 (N_18770,N_15292,N_14153);
nor U18771 (N_18771,N_15102,N_14506);
and U18772 (N_18772,N_13247,N_14628);
nand U18773 (N_18773,N_14289,N_14224);
xnor U18774 (N_18774,N_13105,N_13990);
and U18775 (N_18775,N_15075,N_13863);
nand U18776 (N_18776,N_14163,N_15828);
xor U18777 (N_18777,N_13898,N_15555);
and U18778 (N_18778,N_15206,N_15258);
xnor U18779 (N_18779,N_13115,N_13504);
xor U18780 (N_18780,N_12817,N_13918);
or U18781 (N_18781,N_15904,N_13434);
and U18782 (N_18782,N_13505,N_15708);
nand U18783 (N_18783,N_15662,N_14958);
and U18784 (N_18784,N_15918,N_14131);
and U18785 (N_18785,N_15570,N_14510);
xnor U18786 (N_18786,N_13860,N_13783);
and U18787 (N_18787,N_13932,N_12411);
or U18788 (N_18788,N_13496,N_14798);
xor U18789 (N_18789,N_12945,N_14712);
nor U18790 (N_18790,N_15915,N_15614);
nor U18791 (N_18791,N_12870,N_14589);
and U18792 (N_18792,N_15828,N_14244);
nor U18793 (N_18793,N_14879,N_12601);
nand U18794 (N_18794,N_13088,N_15681);
xnor U18795 (N_18795,N_13767,N_15596);
nand U18796 (N_18796,N_13084,N_13061);
nor U18797 (N_18797,N_14641,N_14153);
and U18798 (N_18798,N_14132,N_15481);
nor U18799 (N_18799,N_13499,N_14824);
xor U18800 (N_18800,N_12222,N_13573);
and U18801 (N_18801,N_13065,N_14670);
or U18802 (N_18802,N_13517,N_14724);
nand U18803 (N_18803,N_12633,N_13877);
nor U18804 (N_18804,N_13449,N_14072);
or U18805 (N_18805,N_13216,N_15577);
nor U18806 (N_18806,N_15712,N_15441);
nand U18807 (N_18807,N_13812,N_14687);
and U18808 (N_18808,N_14117,N_14734);
xor U18809 (N_18809,N_15416,N_15276);
nand U18810 (N_18810,N_14687,N_14161);
nor U18811 (N_18811,N_14569,N_14938);
and U18812 (N_18812,N_13839,N_15472);
and U18813 (N_18813,N_13974,N_15822);
nand U18814 (N_18814,N_14198,N_15487);
xor U18815 (N_18815,N_13853,N_12433);
or U18816 (N_18816,N_12984,N_12404);
and U18817 (N_18817,N_12011,N_13317);
nand U18818 (N_18818,N_12918,N_12441);
nand U18819 (N_18819,N_14759,N_15822);
nand U18820 (N_18820,N_14213,N_12577);
nand U18821 (N_18821,N_15398,N_12718);
nand U18822 (N_18822,N_15622,N_12069);
xnor U18823 (N_18823,N_14022,N_12761);
xor U18824 (N_18824,N_15365,N_14698);
or U18825 (N_18825,N_12109,N_13872);
xnor U18826 (N_18826,N_14002,N_14758);
xnor U18827 (N_18827,N_14807,N_12615);
or U18828 (N_18828,N_12477,N_12405);
or U18829 (N_18829,N_12530,N_14994);
nand U18830 (N_18830,N_15631,N_14577);
nand U18831 (N_18831,N_15678,N_13211);
nand U18832 (N_18832,N_15906,N_15893);
or U18833 (N_18833,N_14563,N_13658);
nor U18834 (N_18834,N_14505,N_13757);
or U18835 (N_18835,N_13078,N_13697);
and U18836 (N_18836,N_14060,N_15486);
or U18837 (N_18837,N_13958,N_14780);
and U18838 (N_18838,N_14039,N_12483);
or U18839 (N_18839,N_14807,N_13259);
nand U18840 (N_18840,N_12325,N_13740);
or U18841 (N_18841,N_13544,N_12416);
and U18842 (N_18842,N_12904,N_13246);
nor U18843 (N_18843,N_14469,N_13645);
nor U18844 (N_18844,N_13020,N_12238);
and U18845 (N_18845,N_13228,N_15141);
nand U18846 (N_18846,N_13149,N_14388);
or U18847 (N_18847,N_12833,N_14270);
nand U18848 (N_18848,N_15762,N_15447);
nand U18849 (N_18849,N_15089,N_13784);
nor U18850 (N_18850,N_13240,N_15598);
nand U18851 (N_18851,N_14745,N_13238);
xor U18852 (N_18852,N_13998,N_15064);
nor U18853 (N_18853,N_15368,N_14476);
xnor U18854 (N_18854,N_12382,N_15620);
nand U18855 (N_18855,N_14079,N_12463);
or U18856 (N_18856,N_14540,N_12175);
or U18857 (N_18857,N_15128,N_13586);
xor U18858 (N_18858,N_14429,N_15464);
xor U18859 (N_18859,N_15161,N_15202);
and U18860 (N_18860,N_15624,N_13210);
xnor U18861 (N_18861,N_14967,N_13011);
nand U18862 (N_18862,N_15301,N_12536);
and U18863 (N_18863,N_12296,N_12184);
nor U18864 (N_18864,N_12510,N_14678);
or U18865 (N_18865,N_13708,N_14943);
xor U18866 (N_18866,N_12559,N_13261);
nor U18867 (N_18867,N_14934,N_15273);
nor U18868 (N_18868,N_13323,N_15417);
xnor U18869 (N_18869,N_14459,N_13072);
and U18870 (N_18870,N_15836,N_13357);
nand U18871 (N_18871,N_13927,N_13891);
nand U18872 (N_18872,N_14335,N_12913);
or U18873 (N_18873,N_14587,N_15674);
and U18874 (N_18874,N_12872,N_14328);
xor U18875 (N_18875,N_13338,N_15854);
nand U18876 (N_18876,N_12750,N_12511);
nand U18877 (N_18877,N_12769,N_15949);
nor U18878 (N_18878,N_13091,N_15793);
nand U18879 (N_18879,N_13602,N_12982);
nor U18880 (N_18880,N_13006,N_14063);
and U18881 (N_18881,N_15037,N_14749);
nor U18882 (N_18882,N_15995,N_12156);
nor U18883 (N_18883,N_14296,N_12239);
nor U18884 (N_18884,N_15348,N_15608);
and U18885 (N_18885,N_12348,N_13556);
or U18886 (N_18886,N_13128,N_15696);
nand U18887 (N_18887,N_15984,N_15167);
and U18888 (N_18888,N_13084,N_13360);
or U18889 (N_18889,N_14385,N_15948);
and U18890 (N_18890,N_13127,N_13798);
or U18891 (N_18891,N_15488,N_13409);
nand U18892 (N_18892,N_15108,N_14510);
nor U18893 (N_18893,N_15695,N_14462);
or U18894 (N_18894,N_14565,N_15604);
nor U18895 (N_18895,N_12731,N_15316);
nor U18896 (N_18896,N_14513,N_14898);
xnor U18897 (N_18897,N_14107,N_14924);
or U18898 (N_18898,N_13517,N_15751);
nand U18899 (N_18899,N_14762,N_14734);
and U18900 (N_18900,N_13255,N_14434);
nor U18901 (N_18901,N_12356,N_12288);
or U18902 (N_18902,N_14496,N_14539);
xor U18903 (N_18903,N_14046,N_14796);
xnor U18904 (N_18904,N_13547,N_15866);
nand U18905 (N_18905,N_14592,N_14814);
or U18906 (N_18906,N_14189,N_13874);
nand U18907 (N_18907,N_14291,N_12974);
and U18908 (N_18908,N_14866,N_14426);
nand U18909 (N_18909,N_15793,N_13658);
or U18910 (N_18910,N_13696,N_13562);
or U18911 (N_18911,N_13256,N_15726);
nand U18912 (N_18912,N_12093,N_13277);
xnor U18913 (N_18913,N_15775,N_12285);
and U18914 (N_18914,N_12343,N_13702);
nand U18915 (N_18915,N_15365,N_12263);
or U18916 (N_18916,N_13058,N_15514);
xnor U18917 (N_18917,N_13163,N_15194);
nor U18918 (N_18918,N_14160,N_15673);
xnor U18919 (N_18919,N_15061,N_15549);
nor U18920 (N_18920,N_15286,N_14739);
nor U18921 (N_18921,N_15469,N_13556);
nand U18922 (N_18922,N_13936,N_13429);
nand U18923 (N_18923,N_14359,N_12510);
xor U18924 (N_18924,N_12457,N_13085);
nand U18925 (N_18925,N_15010,N_15897);
or U18926 (N_18926,N_12377,N_13442);
and U18927 (N_18927,N_13360,N_13249);
and U18928 (N_18928,N_14807,N_12307);
and U18929 (N_18929,N_13000,N_14107);
and U18930 (N_18930,N_14828,N_14448);
or U18931 (N_18931,N_12850,N_12862);
and U18932 (N_18932,N_15520,N_15985);
and U18933 (N_18933,N_15998,N_15793);
and U18934 (N_18934,N_14099,N_15964);
nor U18935 (N_18935,N_12239,N_14958);
or U18936 (N_18936,N_13033,N_12372);
nand U18937 (N_18937,N_14352,N_14485);
nor U18938 (N_18938,N_14721,N_15678);
nor U18939 (N_18939,N_12501,N_15533);
or U18940 (N_18940,N_15837,N_12099);
and U18941 (N_18941,N_14299,N_15214);
nor U18942 (N_18942,N_15006,N_12273);
nand U18943 (N_18943,N_13221,N_13449);
xor U18944 (N_18944,N_15069,N_15530);
nor U18945 (N_18945,N_13693,N_13591);
or U18946 (N_18946,N_15151,N_15668);
xnor U18947 (N_18947,N_15506,N_12251);
or U18948 (N_18948,N_15702,N_14011);
xor U18949 (N_18949,N_12470,N_14707);
nor U18950 (N_18950,N_12724,N_13995);
and U18951 (N_18951,N_12024,N_15200);
nor U18952 (N_18952,N_13301,N_14761);
and U18953 (N_18953,N_14763,N_15703);
xnor U18954 (N_18954,N_15589,N_13839);
and U18955 (N_18955,N_14052,N_13454);
nor U18956 (N_18956,N_12466,N_14685);
xor U18957 (N_18957,N_15914,N_15484);
xor U18958 (N_18958,N_14341,N_12422);
or U18959 (N_18959,N_15409,N_13690);
and U18960 (N_18960,N_12611,N_13230);
nand U18961 (N_18961,N_13330,N_15782);
nand U18962 (N_18962,N_13536,N_12039);
nor U18963 (N_18963,N_13020,N_12127);
xnor U18964 (N_18964,N_12371,N_14545);
nand U18965 (N_18965,N_13643,N_15056);
xnor U18966 (N_18966,N_13511,N_14610);
and U18967 (N_18967,N_14713,N_12602);
nand U18968 (N_18968,N_15609,N_12893);
nor U18969 (N_18969,N_13237,N_13202);
nor U18970 (N_18970,N_14680,N_13272);
and U18971 (N_18971,N_12174,N_12926);
nor U18972 (N_18972,N_14517,N_15301);
and U18973 (N_18973,N_13968,N_14554);
nor U18974 (N_18974,N_12341,N_12698);
nor U18975 (N_18975,N_13335,N_14019);
nor U18976 (N_18976,N_15585,N_15500);
and U18977 (N_18977,N_14604,N_15210);
nand U18978 (N_18978,N_12638,N_12577);
or U18979 (N_18979,N_13796,N_14009);
xor U18980 (N_18980,N_13393,N_15857);
xnor U18981 (N_18981,N_15367,N_12096);
nand U18982 (N_18982,N_14448,N_14607);
or U18983 (N_18983,N_14267,N_13556);
nand U18984 (N_18984,N_15173,N_13519);
nand U18985 (N_18985,N_15428,N_15253);
or U18986 (N_18986,N_14279,N_13314);
nor U18987 (N_18987,N_15162,N_13614);
nand U18988 (N_18988,N_13137,N_15288);
xnor U18989 (N_18989,N_12230,N_12660);
or U18990 (N_18990,N_12812,N_14600);
xnor U18991 (N_18991,N_13578,N_15885);
nor U18992 (N_18992,N_13336,N_14933);
nor U18993 (N_18993,N_12365,N_14830);
nand U18994 (N_18994,N_14271,N_12036);
xnor U18995 (N_18995,N_13200,N_14047);
or U18996 (N_18996,N_13626,N_14374);
or U18997 (N_18997,N_13966,N_12388);
and U18998 (N_18998,N_13540,N_12044);
xnor U18999 (N_18999,N_13855,N_14232);
xor U19000 (N_19000,N_12278,N_14940);
nor U19001 (N_19001,N_14163,N_12558);
nand U19002 (N_19002,N_14811,N_15784);
xnor U19003 (N_19003,N_12330,N_14190);
and U19004 (N_19004,N_13092,N_15696);
nor U19005 (N_19005,N_12256,N_14363);
xor U19006 (N_19006,N_14544,N_12552);
and U19007 (N_19007,N_15926,N_12101);
nand U19008 (N_19008,N_14555,N_13985);
or U19009 (N_19009,N_12165,N_13514);
or U19010 (N_19010,N_13353,N_12673);
or U19011 (N_19011,N_12706,N_14509);
or U19012 (N_19012,N_13483,N_14633);
xor U19013 (N_19013,N_14503,N_13161);
and U19014 (N_19014,N_14741,N_14236);
nand U19015 (N_19015,N_15313,N_14429);
or U19016 (N_19016,N_15403,N_14027);
or U19017 (N_19017,N_14439,N_13361);
xor U19018 (N_19018,N_13568,N_12255);
or U19019 (N_19019,N_13537,N_15034);
xor U19020 (N_19020,N_13144,N_13850);
or U19021 (N_19021,N_14071,N_13667);
or U19022 (N_19022,N_14137,N_12148);
nor U19023 (N_19023,N_14732,N_14329);
nand U19024 (N_19024,N_14367,N_14864);
nor U19025 (N_19025,N_14115,N_12900);
or U19026 (N_19026,N_13153,N_13104);
xor U19027 (N_19027,N_15683,N_13764);
or U19028 (N_19028,N_13591,N_12807);
or U19029 (N_19029,N_12077,N_13999);
nor U19030 (N_19030,N_15240,N_13364);
and U19031 (N_19031,N_12821,N_14164);
nor U19032 (N_19032,N_15881,N_13062);
nand U19033 (N_19033,N_15170,N_12325);
nor U19034 (N_19034,N_13239,N_12547);
xor U19035 (N_19035,N_12323,N_12780);
or U19036 (N_19036,N_14275,N_13227);
xnor U19037 (N_19037,N_14324,N_13437);
nor U19038 (N_19038,N_12481,N_13585);
and U19039 (N_19039,N_13189,N_13334);
xnor U19040 (N_19040,N_12658,N_12579);
nand U19041 (N_19041,N_14375,N_13151);
xor U19042 (N_19042,N_13660,N_15045);
or U19043 (N_19043,N_14280,N_12533);
or U19044 (N_19044,N_12824,N_13497);
nand U19045 (N_19045,N_15061,N_14518);
xor U19046 (N_19046,N_12630,N_15499);
nor U19047 (N_19047,N_15513,N_14863);
and U19048 (N_19048,N_12694,N_14998);
and U19049 (N_19049,N_14800,N_15715);
and U19050 (N_19050,N_12238,N_12800);
and U19051 (N_19051,N_12210,N_14674);
nand U19052 (N_19052,N_15218,N_12606);
and U19053 (N_19053,N_13947,N_13804);
nand U19054 (N_19054,N_15040,N_13114);
and U19055 (N_19055,N_13457,N_15074);
or U19056 (N_19056,N_13000,N_15942);
xor U19057 (N_19057,N_15510,N_13850);
nand U19058 (N_19058,N_15084,N_15746);
nand U19059 (N_19059,N_15986,N_15375);
xnor U19060 (N_19060,N_12566,N_13973);
or U19061 (N_19061,N_14373,N_13226);
nor U19062 (N_19062,N_14852,N_15195);
and U19063 (N_19063,N_13283,N_14334);
and U19064 (N_19064,N_13909,N_14279);
or U19065 (N_19065,N_15963,N_13053);
and U19066 (N_19066,N_13322,N_13107);
or U19067 (N_19067,N_15959,N_15107);
and U19068 (N_19068,N_15358,N_14811);
xnor U19069 (N_19069,N_12123,N_14280);
and U19070 (N_19070,N_12276,N_12836);
nor U19071 (N_19071,N_12999,N_14880);
nand U19072 (N_19072,N_14923,N_13908);
and U19073 (N_19073,N_13678,N_14035);
and U19074 (N_19074,N_15918,N_15244);
nor U19075 (N_19075,N_13265,N_15019);
nand U19076 (N_19076,N_14058,N_13768);
nor U19077 (N_19077,N_13095,N_13591);
xnor U19078 (N_19078,N_14405,N_13571);
nand U19079 (N_19079,N_13340,N_15393);
xnor U19080 (N_19080,N_15405,N_15173);
xnor U19081 (N_19081,N_14545,N_13113);
or U19082 (N_19082,N_12550,N_12781);
nor U19083 (N_19083,N_14191,N_13225);
xor U19084 (N_19084,N_12508,N_13825);
xor U19085 (N_19085,N_12718,N_13459);
xnor U19086 (N_19086,N_12243,N_15508);
or U19087 (N_19087,N_13853,N_14122);
nand U19088 (N_19088,N_12970,N_13621);
and U19089 (N_19089,N_12912,N_13131);
xor U19090 (N_19090,N_14604,N_13088);
or U19091 (N_19091,N_14571,N_14036);
and U19092 (N_19092,N_13423,N_15816);
xor U19093 (N_19093,N_12132,N_14306);
xor U19094 (N_19094,N_14523,N_13046);
nand U19095 (N_19095,N_13584,N_15093);
nand U19096 (N_19096,N_15692,N_14756);
xor U19097 (N_19097,N_13038,N_15287);
xnor U19098 (N_19098,N_12948,N_14132);
nor U19099 (N_19099,N_12757,N_13371);
xor U19100 (N_19100,N_14704,N_12276);
xor U19101 (N_19101,N_12161,N_13906);
and U19102 (N_19102,N_13015,N_12348);
xnor U19103 (N_19103,N_15579,N_14538);
and U19104 (N_19104,N_15424,N_13552);
nor U19105 (N_19105,N_13326,N_14450);
or U19106 (N_19106,N_14806,N_13946);
and U19107 (N_19107,N_14890,N_15191);
nor U19108 (N_19108,N_12315,N_14659);
or U19109 (N_19109,N_12237,N_15369);
and U19110 (N_19110,N_12005,N_14974);
xnor U19111 (N_19111,N_15357,N_13420);
or U19112 (N_19112,N_14216,N_12968);
nor U19113 (N_19113,N_14549,N_15378);
xor U19114 (N_19114,N_14786,N_14837);
xor U19115 (N_19115,N_12285,N_14075);
nor U19116 (N_19116,N_15593,N_14768);
xnor U19117 (N_19117,N_13606,N_14714);
nor U19118 (N_19118,N_12187,N_13147);
xor U19119 (N_19119,N_14170,N_15549);
xnor U19120 (N_19120,N_15619,N_12474);
or U19121 (N_19121,N_14334,N_13450);
nor U19122 (N_19122,N_14728,N_12835);
and U19123 (N_19123,N_12986,N_14812);
xnor U19124 (N_19124,N_15871,N_12095);
and U19125 (N_19125,N_12798,N_13371);
nand U19126 (N_19126,N_14282,N_15435);
or U19127 (N_19127,N_12250,N_14655);
nor U19128 (N_19128,N_14619,N_12810);
nand U19129 (N_19129,N_13619,N_14505);
nor U19130 (N_19130,N_13045,N_14932);
xor U19131 (N_19131,N_13387,N_15472);
nand U19132 (N_19132,N_13900,N_12897);
nand U19133 (N_19133,N_13243,N_12870);
xor U19134 (N_19134,N_12275,N_15240);
nand U19135 (N_19135,N_15906,N_12795);
and U19136 (N_19136,N_14456,N_12778);
nor U19137 (N_19137,N_12368,N_14708);
xnor U19138 (N_19138,N_14004,N_15354);
nand U19139 (N_19139,N_12049,N_14108);
nor U19140 (N_19140,N_14664,N_13528);
nand U19141 (N_19141,N_15009,N_14965);
or U19142 (N_19142,N_12442,N_13064);
nor U19143 (N_19143,N_13938,N_14359);
nand U19144 (N_19144,N_12104,N_13081);
nand U19145 (N_19145,N_13487,N_14784);
or U19146 (N_19146,N_13803,N_14779);
and U19147 (N_19147,N_13905,N_12770);
or U19148 (N_19148,N_14960,N_13556);
nor U19149 (N_19149,N_12813,N_14097);
nand U19150 (N_19150,N_15116,N_13027);
nor U19151 (N_19151,N_14603,N_13606);
xor U19152 (N_19152,N_15034,N_12433);
nand U19153 (N_19153,N_12404,N_12272);
nor U19154 (N_19154,N_12323,N_12969);
xor U19155 (N_19155,N_13027,N_15095);
xor U19156 (N_19156,N_14931,N_13248);
or U19157 (N_19157,N_15374,N_12527);
or U19158 (N_19158,N_15213,N_12605);
nand U19159 (N_19159,N_14789,N_15303);
or U19160 (N_19160,N_15651,N_12771);
and U19161 (N_19161,N_12817,N_14558);
xnor U19162 (N_19162,N_13777,N_14633);
xor U19163 (N_19163,N_14538,N_12212);
or U19164 (N_19164,N_12095,N_15452);
nand U19165 (N_19165,N_14244,N_14006);
and U19166 (N_19166,N_13755,N_15153);
nor U19167 (N_19167,N_12366,N_13006);
nor U19168 (N_19168,N_13746,N_15664);
nor U19169 (N_19169,N_12927,N_12064);
nor U19170 (N_19170,N_15967,N_15545);
and U19171 (N_19171,N_13783,N_13246);
or U19172 (N_19172,N_15027,N_14389);
xnor U19173 (N_19173,N_13490,N_14831);
and U19174 (N_19174,N_12495,N_13010);
nor U19175 (N_19175,N_14645,N_15563);
and U19176 (N_19176,N_13671,N_13953);
nor U19177 (N_19177,N_13759,N_15554);
xor U19178 (N_19178,N_12138,N_12165);
or U19179 (N_19179,N_12331,N_12274);
or U19180 (N_19180,N_13301,N_12388);
nor U19181 (N_19181,N_15330,N_14441);
nand U19182 (N_19182,N_12713,N_15272);
xnor U19183 (N_19183,N_14535,N_14906);
and U19184 (N_19184,N_12186,N_14148);
nor U19185 (N_19185,N_14597,N_12851);
nor U19186 (N_19186,N_15699,N_14996);
and U19187 (N_19187,N_12993,N_14823);
nor U19188 (N_19188,N_13570,N_12354);
xnor U19189 (N_19189,N_12549,N_13598);
xor U19190 (N_19190,N_14029,N_14193);
or U19191 (N_19191,N_14543,N_13235);
xnor U19192 (N_19192,N_12782,N_15460);
nand U19193 (N_19193,N_15183,N_15503);
and U19194 (N_19194,N_14313,N_14523);
nand U19195 (N_19195,N_14115,N_12616);
xor U19196 (N_19196,N_12351,N_13926);
or U19197 (N_19197,N_13700,N_14354);
xor U19198 (N_19198,N_12915,N_12456);
or U19199 (N_19199,N_13589,N_15913);
or U19200 (N_19200,N_12447,N_15369);
nor U19201 (N_19201,N_15880,N_12651);
xnor U19202 (N_19202,N_15364,N_14724);
xor U19203 (N_19203,N_12437,N_13391);
or U19204 (N_19204,N_13217,N_14696);
and U19205 (N_19205,N_13274,N_13680);
xnor U19206 (N_19206,N_14756,N_13430);
nand U19207 (N_19207,N_14972,N_12329);
nor U19208 (N_19208,N_14162,N_15677);
nand U19209 (N_19209,N_12409,N_15151);
and U19210 (N_19210,N_13736,N_12665);
and U19211 (N_19211,N_13111,N_13311);
and U19212 (N_19212,N_15603,N_13624);
and U19213 (N_19213,N_12803,N_14594);
and U19214 (N_19214,N_12831,N_15229);
and U19215 (N_19215,N_12744,N_12180);
or U19216 (N_19216,N_13160,N_14451);
or U19217 (N_19217,N_13088,N_14908);
xnor U19218 (N_19218,N_15704,N_14993);
nor U19219 (N_19219,N_15760,N_14171);
nand U19220 (N_19220,N_15140,N_15001);
and U19221 (N_19221,N_13234,N_12064);
nand U19222 (N_19222,N_15710,N_15801);
xnor U19223 (N_19223,N_13368,N_13775);
and U19224 (N_19224,N_14762,N_13080);
nand U19225 (N_19225,N_13473,N_13350);
and U19226 (N_19226,N_13439,N_13013);
and U19227 (N_19227,N_14346,N_14681);
nand U19228 (N_19228,N_12818,N_13051);
and U19229 (N_19229,N_12042,N_15288);
nor U19230 (N_19230,N_12130,N_12988);
xor U19231 (N_19231,N_12947,N_12047);
and U19232 (N_19232,N_15321,N_12494);
nand U19233 (N_19233,N_14636,N_15377);
nand U19234 (N_19234,N_14648,N_12442);
nand U19235 (N_19235,N_12310,N_15906);
nor U19236 (N_19236,N_12579,N_15808);
and U19237 (N_19237,N_13026,N_12326);
nor U19238 (N_19238,N_15022,N_13479);
nor U19239 (N_19239,N_13991,N_14740);
nand U19240 (N_19240,N_13907,N_14594);
xnor U19241 (N_19241,N_13121,N_13623);
nand U19242 (N_19242,N_12844,N_15976);
nand U19243 (N_19243,N_15972,N_15278);
and U19244 (N_19244,N_12389,N_12704);
and U19245 (N_19245,N_15893,N_14506);
or U19246 (N_19246,N_15659,N_13527);
xnor U19247 (N_19247,N_12262,N_14192);
nand U19248 (N_19248,N_13431,N_15969);
nand U19249 (N_19249,N_13501,N_13296);
or U19250 (N_19250,N_12324,N_15865);
and U19251 (N_19251,N_15446,N_12149);
and U19252 (N_19252,N_12545,N_12810);
nor U19253 (N_19253,N_13454,N_15843);
and U19254 (N_19254,N_12755,N_12003);
nor U19255 (N_19255,N_15278,N_15090);
nand U19256 (N_19256,N_15777,N_12324);
nand U19257 (N_19257,N_12569,N_12807);
nor U19258 (N_19258,N_12986,N_13180);
xnor U19259 (N_19259,N_15871,N_14256);
nor U19260 (N_19260,N_14942,N_15855);
nand U19261 (N_19261,N_14895,N_15809);
nor U19262 (N_19262,N_14916,N_13072);
xnor U19263 (N_19263,N_14085,N_12508);
and U19264 (N_19264,N_15946,N_12746);
and U19265 (N_19265,N_15476,N_13337);
nand U19266 (N_19266,N_14166,N_15399);
nand U19267 (N_19267,N_12254,N_14120);
nor U19268 (N_19268,N_15682,N_13495);
xnor U19269 (N_19269,N_12556,N_15706);
nor U19270 (N_19270,N_15573,N_12792);
nand U19271 (N_19271,N_12924,N_14304);
xor U19272 (N_19272,N_14073,N_13294);
and U19273 (N_19273,N_14603,N_15055);
nor U19274 (N_19274,N_12266,N_12713);
xnor U19275 (N_19275,N_15987,N_14348);
nor U19276 (N_19276,N_13653,N_13298);
or U19277 (N_19277,N_13824,N_13282);
and U19278 (N_19278,N_13885,N_15944);
nor U19279 (N_19279,N_14312,N_12769);
or U19280 (N_19280,N_13578,N_15225);
xor U19281 (N_19281,N_13112,N_12407);
nand U19282 (N_19282,N_13274,N_15667);
nand U19283 (N_19283,N_14635,N_15319);
nor U19284 (N_19284,N_15537,N_14930);
nand U19285 (N_19285,N_12132,N_12410);
nor U19286 (N_19286,N_14861,N_13431);
or U19287 (N_19287,N_13697,N_12087);
nor U19288 (N_19288,N_15753,N_14708);
xor U19289 (N_19289,N_12933,N_15630);
or U19290 (N_19290,N_15811,N_13464);
and U19291 (N_19291,N_15066,N_14091);
nor U19292 (N_19292,N_14792,N_14324);
nor U19293 (N_19293,N_15723,N_15915);
and U19294 (N_19294,N_15756,N_12559);
nand U19295 (N_19295,N_14189,N_13756);
or U19296 (N_19296,N_15082,N_13551);
xor U19297 (N_19297,N_13028,N_12691);
or U19298 (N_19298,N_12223,N_12921);
nand U19299 (N_19299,N_12941,N_13335);
and U19300 (N_19300,N_13129,N_12065);
nor U19301 (N_19301,N_15609,N_12176);
or U19302 (N_19302,N_14335,N_14049);
nor U19303 (N_19303,N_14996,N_13623);
nor U19304 (N_19304,N_13838,N_15956);
nand U19305 (N_19305,N_14224,N_15854);
nor U19306 (N_19306,N_13885,N_15395);
nor U19307 (N_19307,N_15341,N_14339);
nand U19308 (N_19308,N_13181,N_12240);
xnor U19309 (N_19309,N_15249,N_15369);
nor U19310 (N_19310,N_15474,N_12246);
nand U19311 (N_19311,N_12814,N_13928);
nand U19312 (N_19312,N_14040,N_14599);
nor U19313 (N_19313,N_14270,N_13348);
nand U19314 (N_19314,N_14034,N_14795);
and U19315 (N_19315,N_15865,N_12010);
nand U19316 (N_19316,N_14623,N_15546);
nor U19317 (N_19317,N_15487,N_14981);
and U19318 (N_19318,N_14361,N_13346);
xor U19319 (N_19319,N_13177,N_13504);
or U19320 (N_19320,N_13154,N_13778);
and U19321 (N_19321,N_15246,N_13378);
nor U19322 (N_19322,N_12484,N_12988);
and U19323 (N_19323,N_15619,N_13189);
nor U19324 (N_19324,N_14589,N_12768);
or U19325 (N_19325,N_15002,N_15874);
and U19326 (N_19326,N_13486,N_15061);
nand U19327 (N_19327,N_15846,N_15736);
nor U19328 (N_19328,N_14152,N_13596);
and U19329 (N_19329,N_14872,N_13905);
nand U19330 (N_19330,N_15455,N_14420);
or U19331 (N_19331,N_14416,N_14765);
xnor U19332 (N_19332,N_12829,N_14361);
and U19333 (N_19333,N_14662,N_14962);
nand U19334 (N_19334,N_15540,N_14640);
and U19335 (N_19335,N_13970,N_12119);
xnor U19336 (N_19336,N_13808,N_12906);
or U19337 (N_19337,N_12106,N_13549);
nor U19338 (N_19338,N_14346,N_15411);
nand U19339 (N_19339,N_15720,N_14376);
or U19340 (N_19340,N_14782,N_12173);
xnor U19341 (N_19341,N_13846,N_14602);
or U19342 (N_19342,N_15442,N_12382);
and U19343 (N_19343,N_13155,N_15362);
xor U19344 (N_19344,N_15581,N_14381);
nor U19345 (N_19345,N_14574,N_13762);
xnor U19346 (N_19346,N_14141,N_12830);
and U19347 (N_19347,N_15695,N_15073);
nor U19348 (N_19348,N_13019,N_15039);
xor U19349 (N_19349,N_13286,N_15186);
nor U19350 (N_19350,N_13091,N_13002);
nor U19351 (N_19351,N_13035,N_13004);
nand U19352 (N_19352,N_14721,N_15129);
and U19353 (N_19353,N_15886,N_12424);
xor U19354 (N_19354,N_12768,N_15688);
nand U19355 (N_19355,N_12095,N_13398);
nand U19356 (N_19356,N_15279,N_13626);
or U19357 (N_19357,N_14504,N_13595);
nand U19358 (N_19358,N_14936,N_14016);
or U19359 (N_19359,N_14031,N_13600);
xnor U19360 (N_19360,N_14507,N_12618);
and U19361 (N_19361,N_13897,N_14874);
or U19362 (N_19362,N_15090,N_14926);
and U19363 (N_19363,N_12441,N_15647);
nor U19364 (N_19364,N_15284,N_14570);
and U19365 (N_19365,N_12642,N_15801);
nor U19366 (N_19366,N_13774,N_15075);
or U19367 (N_19367,N_14007,N_14817);
nand U19368 (N_19368,N_15250,N_15330);
nor U19369 (N_19369,N_15969,N_14347);
nor U19370 (N_19370,N_13287,N_14522);
and U19371 (N_19371,N_14164,N_12071);
nand U19372 (N_19372,N_14630,N_14268);
nor U19373 (N_19373,N_13263,N_14441);
nand U19374 (N_19374,N_13582,N_13192);
and U19375 (N_19375,N_15576,N_12927);
or U19376 (N_19376,N_14637,N_13980);
xor U19377 (N_19377,N_12278,N_15240);
nor U19378 (N_19378,N_12514,N_15477);
and U19379 (N_19379,N_12373,N_13263);
nand U19380 (N_19380,N_12462,N_14652);
or U19381 (N_19381,N_13595,N_12386);
nor U19382 (N_19382,N_14639,N_15200);
or U19383 (N_19383,N_12785,N_14344);
nand U19384 (N_19384,N_12970,N_15190);
or U19385 (N_19385,N_13243,N_14876);
and U19386 (N_19386,N_13639,N_14861);
nor U19387 (N_19387,N_12609,N_12493);
nor U19388 (N_19388,N_14539,N_14345);
xnor U19389 (N_19389,N_12005,N_14759);
xor U19390 (N_19390,N_14003,N_13735);
nor U19391 (N_19391,N_12587,N_14530);
xor U19392 (N_19392,N_12198,N_14826);
xnor U19393 (N_19393,N_13749,N_12034);
and U19394 (N_19394,N_13210,N_14009);
and U19395 (N_19395,N_13988,N_12126);
nor U19396 (N_19396,N_13680,N_14591);
nor U19397 (N_19397,N_14451,N_15743);
and U19398 (N_19398,N_15426,N_15568);
or U19399 (N_19399,N_14587,N_15432);
nand U19400 (N_19400,N_15935,N_12789);
and U19401 (N_19401,N_14955,N_15781);
or U19402 (N_19402,N_15090,N_12998);
or U19403 (N_19403,N_15563,N_14336);
nand U19404 (N_19404,N_12194,N_12449);
or U19405 (N_19405,N_13765,N_12881);
and U19406 (N_19406,N_13177,N_15400);
xnor U19407 (N_19407,N_13582,N_12751);
xor U19408 (N_19408,N_13372,N_12913);
xor U19409 (N_19409,N_12633,N_14258);
nand U19410 (N_19410,N_15613,N_12405);
nor U19411 (N_19411,N_15146,N_14110);
or U19412 (N_19412,N_14535,N_13120);
or U19413 (N_19413,N_15716,N_12131);
and U19414 (N_19414,N_12092,N_15495);
nor U19415 (N_19415,N_12549,N_13252);
nand U19416 (N_19416,N_13272,N_13510);
nand U19417 (N_19417,N_14772,N_15833);
and U19418 (N_19418,N_14784,N_14065);
and U19419 (N_19419,N_14955,N_15084);
and U19420 (N_19420,N_12115,N_12240);
or U19421 (N_19421,N_12180,N_13588);
or U19422 (N_19422,N_12349,N_15979);
nand U19423 (N_19423,N_14511,N_15349);
nor U19424 (N_19424,N_12958,N_15780);
nand U19425 (N_19425,N_12838,N_14815);
or U19426 (N_19426,N_12311,N_12257);
and U19427 (N_19427,N_13371,N_14295);
nor U19428 (N_19428,N_14655,N_13726);
and U19429 (N_19429,N_15171,N_12163);
or U19430 (N_19430,N_14248,N_14300);
and U19431 (N_19431,N_13951,N_12082);
nor U19432 (N_19432,N_13588,N_14186);
nor U19433 (N_19433,N_15772,N_14388);
nand U19434 (N_19434,N_15272,N_13066);
xor U19435 (N_19435,N_13622,N_14985);
or U19436 (N_19436,N_13800,N_14436);
nand U19437 (N_19437,N_12127,N_13361);
nand U19438 (N_19438,N_14324,N_13287);
or U19439 (N_19439,N_12974,N_15208);
or U19440 (N_19440,N_13039,N_15678);
nor U19441 (N_19441,N_15293,N_14997);
nand U19442 (N_19442,N_14755,N_14799);
nor U19443 (N_19443,N_15458,N_13195);
and U19444 (N_19444,N_15766,N_12451);
or U19445 (N_19445,N_13694,N_12050);
and U19446 (N_19446,N_12569,N_13886);
or U19447 (N_19447,N_15742,N_14942);
nand U19448 (N_19448,N_13623,N_12026);
and U19449 (N_19449,N_13674,N_14439);
xor U19450 (N_19450,N_15998,N_14972);
or U19451 (N_19451,N_15329,N_12998);
or U19452 (N_19452,N_14408,N_12941);
or U19453 (N_19453,N_14620,N_15657);
xor U19454 (N_19454,N_14779,N_14679);
xnor U19455 (N_19455,N_14103,N_15163);
or U19456 (N_19456,N_14058,N_14670);
and U19457 (N_19457,N_12312,N_15797);
and U19458 (N_19458,N_15376,N_14255);
or U19459 (N_19459,N_15409,N_15494);
or U19460 (N_19460,N_13696,N_15445);
or U19461 (N_19461,N_13947,N_14768);
and U19462 (N_19462,N_15643,N_15348);
and U19463 (N_19463,N_13686,N_14445);
and U19464 (N_19464,N_14698,N_13222);
nor U19465 (N_19465,N_12966,N_12631);
or U19466 (N_19466,N_15631,N_15480);
xor U19467 (N_19467,N_13936,N_14263);
and U19468 (N_19468,N_12607,N_13695);
or U19469 (N_19469,N_15827,N_14144);
or U19470 (N_19470,N_14449,N_13125);
and U19471 (N_19471,N_15437,N_14721);
and U19472 (N_19472,N_12225,N_14059);
nor U19473 (N_19473,N_12094,N_15053);
nor U19474 (N_19474,N_12715,N_12991);
nand U19475 (N_19475,N_13166,N_14857);
nand U19476 (N_19476,N_13007,N_13070);
nand U19477 (N_19477,N_13613,N_14724);
and U19478 (N_19478,N_14602,N_12930);
nand U19479 (N_19479,N_12634,N_13365);
nor U19480 (N_19480,N_14507,N_14410);
nand U19481 (N_19481,N_14882,N_13764);
xnor U19482 (N_19482,N_13183,N_14271);
or U19483 (N_19483,N_12238,N_15474);
or U19484 (N_19484,N_12551,N_12613);
nand U19485 (N_19485,N_14571,N_12281);
nor U19486 (N_19486,N_13502,N_13766);
and U19487 (N_19487,N_13784,N_15079);
or U19488 (N_19488,N_15778,N_14576);
nor U19489 (N_19489,N_13947,N_13257);
or U19490 (N_19490,N_14013,N_14437);
nor U19491 (N_19491,N_12900,N_14969);
or U19492 (N_19492,N_13048,N_13331);
and U19493 (N_19493,N_14692,N_12614);
nand U19494 (N_19494,N_12123,N_13313);
xor U19495 (N_19495,N_13071,N_12709);
xnor U19496 (N_19496,N_13952,N_14739);
nor U19497 (N_19497,N_12036,N_15049);
nand U19498 (N_19498,N_13164,N_14595);
nand U19499 (N_19499,N_13108,N_13804);
and U19500 (N_19500,N_14312,N_12478);
xor U19501 (N_19501,N_13496,N_13628);
and U19502 (N_19502,N_14103,N_12071);
and U19503 (N_19503,N_14419,N_15392);
and U19504 (N_19504,N_13728,N_13689);
or U19505 (N_19505,N_13635,N_12250);
nand U19506 (N_19506,N_12408,N_12855);
or U19507 (N_19507,N_14385,N_13531);
nand U19508 (N_19508,N_12098,N_13172);
nor U19509 (N_19509,N_13698,N_14942);
nand U19510 (N_19510,N_12921,N_12609);
nor U19511 (N_19511,N_13290,N_14586);
nor U19512 (N_19512,N_14958,N_14413);
nor U19513 (N_19513,N_13313,N_14977);
nor U19514 (N_19514,N_14967,N_15150);
or U19515 (N_19515,N_15876,N_15644);
xor U19516 (N_19516,N_15458,N_15758);
and U19517 (N_19517,N_15977,N_12723);
and U19518 (N_19518,N_13633,N_12627);
and U19519 (N_19519,N_13667,N_12663);
nor U19520 (N_19520,N_14547,N_13739);
or U19521 (N_19521,N_13203,N_13595);
nand U19522 (N_19522,N_14352,N_15082);
or U19523 (N_19523,N_14877,N_12395);
xnor U19524 (N_19524,N_12903,N_12105);
xnor U19525 (N_19525,N_13544,N_13988);
or U19526 (N_19526,N_12246,N_12222);
or U19527 (N_19527,N_12963,N_14165);
xor U19528 (N_19528,N_15097,N_12993);
xor U19529 (N_19529,N_14995,N_13819);
nor U19530 (N_19530,N_14034,N_12060);
nor U19531 (N_19531,N_14752,N_14573);
nand U19532 (N_19532,N_13749,N_12961);
xor U19533 (N_19533,N_14442,N_15730);
or U19534 (N_19534,N_13873,N_12988);
or U19535 (N_19535,N_15770,N_13923);
nand U19536 (N_19536,N_15994,N_15949);
or U19537 (N_19537,N_12438,N_15905);
nor U19538 (N_19538,N_15885,N_15478);
and U19539 (N_19539,N_12639,N_15359);
xnor U19540 (N_19540,N_15226,N_14700);
or U19541 (N_19541,N_13871,N_15304);
nand U19542 (N_19542,N_14599,N_14882);
nand U19543 (N_19543,N_15051,N_14436);
or U19544 (N_19544,N_14578,N_12736);
nor U19545 (N_19545,N_12115,N_15757);
xnor U19546 (N_19546,N_15303,N_14529);
nor U19547 (N_19547,N_15125,N_15222);
and U19548 (N_19548,N_15443,N_15863);
or U19549 (N_19549,N_14380,N_12223);
or U19550 (N_19550,N_15994,N_15894);
xnor U19551 (N_19551,N_14055,N_14447);
nor U19552 (N_19552,N_13501,N_12945);
nor U19553 (N_19553,N_12721,N_15646);
nand U19554 (N_19554,N_15528,N_13341);
nor U19555 (N_19555,N_13187,N_15592);
nor U19556 (N_19556,N_13248,N_12467);
xnor U19557 (N_19557,N_14061,N_12521);
nand U19558 (N_19558,N_14142,N_15409);
nand U19559 (N_19559,N_12024,N_13028);
xnor U19560 (N_19560,N_14459,N_13867);
or U19561 (N_19561,N_14509,N_13777);
xor U19562 (N_19562,N_13971,N_13821);
xor U19563 (N_19563,N_14228,N_14733);
nor U19564 (N_19564,N_15912,N_14342);
nand U19565 (N_19565,N_15564,N_15659);
and U19566 (N_19566,N_12777,N_13849);
xnor U19567 (N_19567,N_12317,N_15897);
and U19568 (N_19568,N_14240,N_15860);
and U19569 (N_19569,N_15140,N_15300);
nand U19570 (N_19570,N_15947,N_15637);
nand U19571 (N_19571,N_12283,N_12464);
xnor U19572 (N_19572,N_15953,N_15358);
and U19573 (N_19573,N_14143,N_12708);
nor U19574 (N_19574,N_12571,N_15459);
or U19575 (N_19575,N_13064,N_14967);
or U19576 (N_19576,N_12884,N_15513);
and U19577 (N_19577,N_15946,N_12574);
nor U19578 (N_19578,N_15800,N_14097);
nand U19579 (N_19579,N_15998,N_12039);
and U19580 (N_19580,N_14992,N_13025);
and U19581 (N_19581,N_12454,N_12159);
and U19582 (N_19582,N_14902,N_12204);
nand U19583 (N_19583,N_12103,N_15668);
nand U19584 (N_19584,N_13853,N_13126);
xor U19585 (N_19585,N_15305,N_12235);
nor U19586 (N_19586,N_13046,N_12737);
nand U19587 (N_19587,N_14145,N_14585);
xnor U19588 (N_19588,N_13285,N_14224);
nor U19589 (N_19589,N_14485,N_12228);
xor U19590 (N_19590,N_14910,N_15878);
and U19591 (N_19591,N_13272,N_13872);
or U19592 (N_19592,N_12461,N_15740);
nor U19593 (N_19593,N_14286,N_12863);
or U19594 (N_19594,N_14176,N_13824);
and U19595 (N_19595,N_14148,N_15592);
xor U19596 (N_19596,N_14393,N_15477);
or U19597 (N_19597,N_15241,N_13128);
nor U19598 (N_19598,N_13493,N_15945);
xor U19599 (N_19599,N_14373,N_12358);
xor U19600 (N_19600,N_13389,N_15596);
xor U19601 (N_19601,N_15525,N_13120);
xnor U19602 (N_19602,N_15108,N_15612);
or U19603 (N_19603,N_12403,N_13154);
xnor U19604 (N_19604,N_15396,N_14252);
and U19605 (N_19605,N_13785,N_12901);
or U19606 (N_19606,N_12587,N_12903);
or U19607 (N_19607,N_13978,N_13109);
nor U19608 (N_19608,N_14696,N_13530);
nor U19609 (N_19609,N_13754,N_12269);
nor U19610 (N_19610,N_14089,N_14245);
xnor U19611 (N_19611,N_12714,N_14930);
and U19612 (N_19612,N_15787,N_15602);
xnor U19613 (N_19613,N_13965,N_14261);
and U19614 (N_19614,N_13935,N_14025);
nand U19615 (N_19615,N_15230,N_13821);
nand U19616 (N_19616,N_12594,N_13849);
nand U19617 (N_19617,N_13129,N_15188);
nand U19618 (N_19618,N_12150,N_13212);
and U19619 (N_19619,N_12013,N_14650);
nand U19620 (N_19620,N_14956,N_15999);
and U19621 (N_19621,N_14064,N_12453);
nand U19622 (N_19622,N_13016,N_12815);
nor U19623 (N_19623,N_15653,N_13850);
nor U19624 (N_19624,N_12044,N_15130);
or U19625 (N_19625,N_14830,N_14607);
or U19626 (N_19626,N_15484,N_15536);
or U19627 (N_19627,N_12894,N_15316);
nor U19628 (N_19628,N_13594,N_13229);
nor U19629 (N_19629,N_12556,N_14537);
xor U19630 (N_19630,N_12292,N_13656);
nand U19631 (N_19631,N_12168,N_15308);
or U19632 (N_19632,N_14338,N_12604);
xnor U19633 (N_19633,N_15345,N_13881);
and U19634 (N_19634,N_13947,N_14865);
nand U19635 (N_19635,N_14184,N_15848);
nor U19636 (N_19636,N_14737,N_13529);
nor U19637 (N_19637,N_15779,N_13368);
nor U19638 (N_19638,N_13491,N_14630);
nand U19639 (N_19639,N_12350,N_13941);
nand U19640 (N_19640,N_12285,N_12074);
nor U19641 (N_19641,N_14348,N_15254);
nor U19642 (N_19642,N_14324,N_14863);
and U19643 (N_19643,N_15639,N_15787);
nor U19644 (N_19644,N_15866,N_14899);
nand U19645 (N_19645,N_13891,N_14587);
nor U19646 (N_19646,N_14314,N_15463);
or U19647 (N_19647,N_14852,N_14806);
and U19648 (N_19648,N_12398,N_13432);
nor U19649 (N_19649,N_13495,N_13213);
xnor U19650 (N_19650,N_12934,N_15919);
nand U19651 (N_19651,N_15106,N_13851);
and U19652 (N_19652,N_12983,N_15658);
xor U19653 (N_19653,N_14999,N_14674);
or U19654 (N_19654,N_13710,N_15850);
nor U19655 (N_19655,N_14186,N_12354);
and U19656 (N_19656,N_15780,N_15746);
nand U19657 (N_19657,N_15285,N_12462);
and U19658 (N_19658,N_14542,N_12650);
xor U19659 (N_19659,N_14965,N_14266);
or U19660 (N_19660,N_13047,N_13182);
and U19661 (N_19661,N_15441,N_15331);
and U19662 (N_19662,N_14273,N_14262);
nor U19663 (N_19663,N_12083,N_14222);
or U19664 (N_19664,N_14978,N_12060);
and U19665 (N_19665,N_12552,N_14832);
nand U19666 (N_19666,N_14670,N_14701);
or U19667 (N_19667,N_14338,N_14653);
or U19668 (N_19668,N_13010,N_12838);
nor U19669 (N_19669,N_15718,N_14480);
xnor U19670 (N_19670,N_12552,N_13587);
xnor U19671 (N_19671,N_15784,N_14211);
nand U19672 (N_19672,N_15989,N_13702);
nor U19673 (N_19673,N_14046,N_14631);
or U19674 (N_19674,N_13083,N_12713);
and U19675 (N_19675,N_12689,N_15792);
or U19676 (N_19676,N_13722,N_15080);
and U19677 (N_19677,N_13798,N_13076);
xor U19678 (N_19678,N_15669,N_15432);
and U19679 (N_19679,N_14744,N_15320);
nor U19680 (N_19680,N_15442,N_13291);
nand U19681 (N_19681,N_12862,N_14389);
nor U19682 (N_19682,N_14568,N_12189);
nor U19683 (N_19683,N_14809,N_12513);
nand U19684 (N_19684,N_15157,N_13321);
xnor U19685 (N_19685,N_14103,N_12292);
xor U19686 (N_19686,N_14215,N_12688);
nor U19687 (N_19687,N_13707,N_12504);
nand U19688 (N_19688,N_14700,N_15292);
nor U19689 (N_19689,N_12834,N_15869);
or U19690 (N_19690,N_15850,N_14563);
nor U19691 (N_19691,N_12897,N_15911);
or U19692 (N_19692,N_14505,N_14176);
nor U19693 (N_19693,N_14148,N_13220);
and U19694 (N_19694,N_14097,N_13918);
nand U19695 (N_19695,N_13070,N_14833);
xor U19696 (N_19696,N_15949,N_12404);
nor U19697 (N_19697,N_12278,N_15054);
nand U19698 (N_19698,N_14523,N_15012);
or U19699 (N_19699,N_12473,N_14460);
xnor U19700 (N_19700,N_14566,N_15068);
xor U19701 (N_19701,N_12720,N_13996);
or U19702 (N_19702,N_14285,N_12597);
nor U19703 (N_19703,N_14122,N_14309);
and U19704 (N_19704,N_13847,N_12035);
or U19705 (N_19705,N_13195,N_15932);
nor U19706 (N_19706,N_14277,N_14193);
and U19707 (N_19707,N_12900,N_13621);
nor U19708 (N_19708,N_13904,N_14614);
xor U19709 (N_19709,N_14581,N_14509);
or U19710 (N_19710,N_13939,N_15398);
and U19711 (N_19711,N_12218,N_14050);
nor U19712 (N_19712,N_12828,N_13854);
and U19713 (N_19713,N_15405,N_14403);
nor U19714 (N_19714,N_14595,N_12719);
xor U19715 (N_19715,N_12496,N_14929);
xnor U19716 (N_19716,N_12410,N_12052);
and U19717 (N_19717,N_13743,N_14264);
nand U19718 (N_19718,N_13022,N_14918);
xor U19719 (N_19719,N_12427,N_13866);
xor U19720 (N_19720,N_14101,N_12151);
nand U19721 (N_19721,N_13985,N_15367);
xor U19722 (N_19722,N_13879,N_13146);
xnor U19723 (N_19723,N_15076,N_13543);
xnor U19724 (N_19724,N_14534,N_12086);
nor U19725 (N_19725,N_13616,N_14373);
nand U19726 (N_19726,N_15252,N_12880);
nand U19727 (N_19727,N_15267,N_15991);
or U19728 (N_19728,N_15471,N_14974);
nand U19729 (N_19729,N_13322,N_13080);
nand U19730 (N_19730,N_13071,N_12346);
and U19731 (N_19731,N_15402,N_15201);
nand U19732 (N_19732,N_13787,N_12579);
nor U19733 (N_19733,N_12041,N_15941);
xor U19734 (N_19734,N_13168,N_13449);
nor U19735 (N_19735,N_14625,N_13249);
or U19736 (N_19736,N_15720,N_12692);
nor U19737 (N_19737,N_13450,N_12810);
and U19738 (N_19738,N_13466,N_12062);
or U19739 (N_19739,N_14482,N_15016);
nand U19740 (N_19740,N_12460,N_14006);
or U19741 (N_19741,N_14600,N_13937);
nor U19742 (N_19742,N_13249,N_12983);
or U19743 (N_19743,N_12525,N_15582);
nor U19744 (N_19744,N_13009,N_15358);
or U19745 (N_19745,N_14263,N_14256);
nand U19746 (N_19746,N_14736,N_13423);
nor U19747 (N_19747,N_15060,N_12919);
nand U19748 (N_19748,N_13342,N_12140);
nand U19749 (N_19749,N_14730,N_14947);
nor U19750 (N_19750,N_14170,N_12699);
nand U19751 (N_19751,N_14200,N_15977);
xor U19752 (N_19752,N_13131,N_13771);
or U19753 (N_19753,N_14714,N_15990);
or U19754 (N_19754,N_14462,N_14435);
xnor U19755 (N_19755,N_14969,N_13204);
or U19756 (N_19756,N_13989,N_12167);
or U19757 (N_19757,N_13639,N_14910);
and U19758 (N_19758,N_14601,N_13760);
nand U19759 (N_19759,N_15187,N_15764);
and U19760 (N_19760,N_13366,N_12523);
nor U19761 (N_19761,N_13699,N_14262);
nor U19762 (N_19762,N_13698,N_14324);
or U19763 (N_19763,N_15470,N_12098);
or U19764 (N_19764,N_12945,N_12399);
and U19765 (N_19765,N_12872,N_15874);
or U19766 (N_19766,N_14846,N_12655);
nand U19767 (N_19767,N_12711,N_12691);
or U19768 (N_19768,N_14792,N_14981);
xnor U19769 (N_19769,N_12337,N_12774);
nor U19770 (N_19770,N_15276,N_15502);
nor U19771 (N_19771,N_13371,N_13562);
or U19772 (N_19772,N_13362,N_15231);
nand U19773 (N_19773,N_15123,N_15479);
or U19774 (N_19774,N_12538,N_13985);
nor U19775 (N_19775,N_13805,N_15915);
xnor U19776 (N_19776,N_15249,N_14355);
xnor U19777 (N_19777,N_15858,N_15152);
nand U19778 (N_19778,N_14383,N_14586);
nor U19779 (N_19779,N_15504,N_15616);
nand U19780 (N_19780,N_15311,N_12457);
and U19781 (N_19781,N_13745,N_14013);
nor U19782 (N_19782,N_13271,N_14102);
nor U19783 (N_19783,N_13269,N_13676);
and U19784 (N_19784,N_13658,N_13970);
and U19785 (N_19785,N_12686,N_14985);
xnor U19786 (N_19786,N_12788,N_14579);
xnor U19787 (N_19787,N_12712,N_12354);
nand U19788 (N_19788,N_15369,N_12863);
nor U19789 (N_19789,N_15880,N_12507);
xnor U19790 (N_19790,N_15375,N_15002);
nor U19791 (N_19791,N_14293,N_15895);
xnor U19792 (N_19792,N_15626,N_15297);
nand U19793 (N_19793,N_14911,N_13463);
nand U19794 (N_19794,N_15875,N_14414);
xnor U19795 (N_19795,N_12556,N_14194);
and U19796 (N_19796,N_14907,N_13533);
or U19797 (N_19797,N_13545,N_15106);
nand U19798 (N_19798,N_14866,N_15364);
nand U19799 (N_19799,N_13757,N_12234);
nand U19800 (N_19800,N_13147,N_12609);
xor U19801 (N_19801,N_13014,N_13241);
nand U19802 (N_19802,N_14300,N_13939);
xor U19803 (N_19803,N_13480,N_12869);
nor U19804 (N_19804,N_13440,N_12333);
nand U19805 (N_19805,N_13441,N_15494);
nand U19806 (N_19806,N_12917,N_14405);
nand U19807 (N_19807,N_14771,N_12213);
and U19808 (N_19808,N_14506,N_12365);
xnor U19809 (N_19809,N_15731,N_15208);
or U19810 (N_19810,N_12139,N_14956);
xor U19811 (N_19811,N_14723,N_15253);
and U19812 (N_19812,N_12613,N_12178);
xnor U19813 (N_19813,N_13841,N_13759);
or U19814 (N_19814,N_15630,N_13421);
nor U19815 (N_19815,N_12397,N_13545);
nor U19816 (N_19816,N_14791,N_12718);
or U19817 (N_19817,N_13894,N_12191);
nor U19818 (N_19818,N_13489,N_15334);
xnor U19819 (N_19819,N_12671,N_12210);
or U19820 (N_19820,N_14433,N_15775);
and U19821 (N_19821,N_14094,N_13865);
nand U19822 (N_19822,N_12611,N_13524);
and U19823 (N_19823,N_15198,N_13070);
or U19824 (N_19824,N_15792,N_12646);
or U19825 (N_19825,N_14148,N_12990);
and U19826 (N_19826,N_15664,N_14907);
and U19827 (N_19827,N_14204,N_12525);
nand U19828 (N_19828,N_12582,N_13438);
or U19829 (N_19829,N_13187,N_12886);
nand U19830 (N_19830,N_12072,N_14179);
or U19831 (N_19831,N_12915,N_14523);
and U19832 (N_19832,N_13702,N_14624);
and U19833 (N_19833,N_13935,N_13444);
xnor U19834 (N_19834,N_14286,N_15489);
or U19835 (N_19835,N_12509,N_13931);
nand U19836 (N_19836,N_15010,N_13895);
or U19837 (N_19837,N_13786,N_15293);
and U19838 (N_19838,N_15693,N_15486);
xnor U19839 (N_19839,N_15706,N_15855);
nand U19840 (N_19840,N_15786,N_15495);
xnor U19841 (N_19841,N_14616,N_12823);
and U19842 (N_19842,N_14322,N_12065);
nand U19843 (N_19843,N_13106,N_13396);
nor U19844 (N_19844,N_14912,N_15455);
or U19845 (N_19845,N_12140,N_14032);
or U19846 (N_19846,N_13054,N_13961);
xor U19847 (N_19847,N_15540,N_14406);
xnor U19848 (N_19848,N_14984,N_14182);
and U19849 (N_19849,N_14412,N_13263);
or U19850 (N_19850,N_12162,N_14215);
xnor U19851 (N_19851,N_13932,N_14154);
xnor U19852 (N_19852,N_14686,N_15919);
nand U19853 (N_19853,N_15623,N_14010);
or U19854 (N_19854,N_15692,N_13659);
nor U19855 (N_19855,N_14380,N_13747);
xnor U19856 (N_19856,N_12701,N_13318);
xnor U19857 (N_19857,N_15923,N_14746);
nand U19858 (N_19858,N_14908,N_12875);
and U19859 (N_19859,N_13450,N_12541);
nand U19860 (N_19860,N_13501,N_15093);
nand U19861 (N_19861,N_13272,N_15640);
nand U19862 (N_19862,N_13990,N_15444);
nor U19863 (N_19863,N_15152,N_14348);
nor U19864 (N_19864,N_13628,N_12138);
nand U19865 (N_19865,N_13259,N_15863);
xor U19866 (N_19866,N_15873,N_15310);
nor U19867 (N_19867,N_15898,N_13815);
and U19868 (N_19868,N_14497,N_13502);
or U19869 (N_19869,N_14857,N_15922);
nor U19870 (N_19870,N_13065,N_15645);
xnor U19871 (N_19871,N_13925,N_13368);
xor U19872 (N_19872,N_13197,N_12359);
nand U19873 (N_19873,N_13665,N_12138);
nor U19874 (N_19874,N_14329,N_13664);
and U19875 (N_19875,N_14228,N_15988);
or U19876 (N_19876,N_13547,N_14160);
or U19877 (N_19877,N_13175,N_15107);
nand U19878 (N_19878,N_15163,N_14856);
xnor U19879 (N_19879,N_14318,N_14766);
nand U19880 (N_19880,N_12393,N_13418);
nand U19881 (N_19881,N_12564,N_12352);
or U19882 (N_19882,N_13460,N_14757);
and U19883 (N_19883,N_14420,N_15119);
nor U19884 (N_19884,N_13309,N_13171);
or U19885 (N_19885,N_15840,N_13480);
or U19886 (N_19886,N_12468,N_13968);
nand U19887 (N_19887,N_14445,N_13526);
and U19888 (N_19888,N_14176,N_15405);
nand U19889 (N_19889,N_14077,N_13396);
or U19890 (N_19890,N_13675,N_15826);
nor U19891 (N_19891,N_15184,N_13470);
nand U19892 (N_19892,N_12731,N_12025);
or U19893 (N_19893,N_14128,N_13816);
nor U19894 (N_19894,N_14570,N_13769);
and U19895 (N_19895,N_12059,N_14651);
xnor U19896 (N_19896,N_13322,N_15598);
nor U19897 (N_19897,N_15433,N_15572);
or U19898 (N_19898,N_12244,N_14657);
xnor U19899 (N_19899,N_13130,N_15409);
and U19900 (N_19900,N_15244,N_13092);
nand U19901 (N_19901,N_12431,N_14051);
or U19902 (N_19902,N_13829,N_14860);
xnor U19903 (N_19903,N_13764,N_15412);
or U19904 (N_19904,N_14507,N_12026);
and U19905 (N_19905,N_14596,N_14031);
nand U19906 (N_19906,N_14073,N_14650);
nor U19907 (N_19907,N_14913,N_13978);
or U19908 (N_19908,N_15104,N_14631);
nand U19909 (N_19909,N_14772,N_13123);
xnor U19910 (N_19910,N_15375,N_15062);
nor U19911 (N_19911,N_14043,N_13529);
and U19912 (N_19912,N_14096,N_14491);
nand U19913 (N_19913,N_15452,N_13580);
or U19914 (N_19914,N_15096,N_13973);
xnor U19915 (N_19915,N_13787,N_12010);
nand U19916 (N_19916,N_13325,N_15113);
or U19917 (N_19917,N_12676,N_15169);
nor U19918 (N_19918,N_13911,N_13444);
xor U19919 (N_19919,N_13473,N_12782);
nand U19920 (N_19920,N_15421,N_12388);
and U19921 (N_19921,N_15691,N_14272);
nand U19922 (N_19922,N_13019,N_14560);
or U19923 (N_19923,N_15046,N_14662);
nor U19924 (N_19924,N_12932,N_12045);
or U19925 (N_19925,N_13166,N_12423);
and U19926 (N_19926,N_12577,N_12498);
nor U19927 (N_19927,N_12672,N_13460);
nor U19928 (N_19928,N_15339,N_12929);
or U19929 (N_19929,N_14851,N_12948);
xnor U19930 (N_19930,N_14454,N_12673);
nand U19931 (N_19931,N_13101,N_13785);
xnor U19932 (N_19932,N_14033,N_14260);
or U19933 (N_19933,N_14938,N_13306);
and U19934 (N_19934,N_12418,N_14258);
nor U19935 (N_19935,N_15349,N_15027);
or U19936 (N_19936,N_13377,N_15186);
xnor U19937 (N_19937,N_13021,N_12523);
or U19938 (N_19938,N_14789,N_13193);
and U19939 (N_19939,N_12244,N_14615);
and U19940 (N_19940,N_14492,N_14951);
nand U19941 (N_19941,N_12069,N_12576);
nand U19942 (N_19942,N_14897,N_14394);
nand U19943 (N_19943,N_13280,N_15227);
or U19944 (N_19944,N_12968,N_13826);
and U19945 (N_19945,N_14289,N_12482);
and U19946 (N_19946,N_12258,N_12200);
or U19947 (N_19947,N_12140,N_14930);
nand U19948 (N_19948,N_13240,N_13346);
nand U19949 (N_19949,N_12931,N_12214);
and U19950 (N_19950,N_14114,N_13234);
xor U19951 (N_19951,N_12312,N_15630);
nand U19952 (N_19952,N_12161,N_13128);
nand U19953 (N_19953,N_14059,N_13655);
nor U19954 (N_19954,N_14262,N_12034);
or U19955 (N_19955,N_15524,N_14300);
nor U19956 (N_19956,N_12213,N_13716);
and U19957 (N_19957,N_14789,N_12134);
and U19958 (N_19958,N_13215,N_12852);
or U19959 (N_19959,N_14336,N_15501);
nor U19960 (N_19960,N_15222,N_13629);
or U19961 (N_19961,N_13438,N_12381);
or U19962 (N_19962,N_12960,N_12040);
xnor U19963 (N_19963,N_15558,N_14189);
nor U19964 (N_19964,N_14099,N_12222);
or U19965 (N_19965,N_15858,N_12768);
nor U19966 (N_19966,N_14790,N_15651);
or U19967 (N_19967,N_15343,N_12702);
xor U19968 (N_19968,N_13013,N_15600);
and U19969 (N_19969,N_14009,N_13852);
nand U19970 (N_19970,N_14394,N_13516);
or U19971 (N_19971,N_14510,N_14255);
or U19972 (N_19972,N_13926,N_14844);
or U19973 (N_19973,N_15278,N_14194);
or U19974 (N_19974,N_13633,N_15135);
nand U19975 (N_19975,N_12967,N_14525);
nand U19976 (N_19976,N_12091,N_14602);
nand U19977 (N_19977,N_13333,N_12494);
nand U19978 (N_19978,N_15087,N_15105);
nor U19979 (N_19979,N_12994,N_12499);
and U19980 (N_19980,N_15885,N_13614);
nand U19981 (N_19981,N_12529,N_12866);
nor U19982 (N_19982,N_14333,N_12550);
nor U19983 (N_19983,N_14741,N_15221);
or U19984 (N_19984,N_14012,N_13991);
or U19985 (N_19985,N_13446,N_15142);
xnor U19986 (N_19986,N_14214,N_14784);
and U19987 (N_19987,N_15625,N_12805);
and U19988 (N_19988,N_13079,N_14916);
nand U19989 (N_19989,N_15699,N_15286);
nand U19990 (N_19990,N_15184,N_13046);
xnor U19991 (N_19991,N_14084,N_15104);
nor U19992 (N_19992,N_12381,N_15650);
or U19993 (N_19993,N_12457,N_12097);
nor U19994 (N_19994,N_15872,N_13095);
xor U19995 (N_19995,N_12719,N_12258);
or U19996 (N_19996,N_13297,N_14333);
and U19997 (N_19997,N_15022,N_13952);
and U19998 (N_19998,N_13129,N_13806);
xnor U19999 (N_19999,N_12378,N_12833);
or UO_0 (O_0,N_16513,N_17427);
xnor UO_1 (O_1,N_16418,N_19851);
xnor UO_2 (O_2,N_16976,N_19781);
xor UO_3 (O_3,N_19409,N_16625);
xnor UO_4 (O_4,N_16721,N_16385);
nand UO_5 (O_5,N_16389,N_19741);
nand UO_6 (O_6,N_17514,N_18363);
xnor UO_7 (O_7,N_18071,N_18420);
nor UO_8 (O_8,N_19522,N_17088);
nand UO_9 (O_9,N_17506,N_19600);
or UO_10 (O_10,N_19029,N_16118);
or UO_11 (O_11,N_18725,N_17830);
and UO_12 (O_12,N_18964,N_16102);
xor UO_13 (O_13,N_17221,N_16877);
nor UO_14 (O_14,N_18489,N_16688);
xor UO_15 (O_15,N_18272,N_19474);
or UO_16 (O_16,N_18008,N_16152);
nand UO_17 (O_17,N_19449,N_18951);
nand UO_18 (O_18,N_16583,N_18395);
or UO_19 (O_19,N_18974,N_16277);
nor UO_20 (O_20,N_17770,N_18419);
xnor UO_21 (O_21,N_18193,N_18744);
and UO_22 (O_22,N_18219,N_17430);
or UO_23 (O_23,N_17069,N_16503);
or UO_24 (O_24,N_19613,N_18844);
nor UO_25 (O_25,N_16028,N_16391);
xor UO_26 (O_26,N_17433,N_19946);
nor UO_27 (O_27,N_19213,N_17455);
nor UO_28 (O_28,N_18471,N_18815);
or UO_29 (O_29,N_16049,N_19265);
nor UO_30 (O_30,N_17867,N_16082);
and UO_31 (O_31,N_16597,N_18559);
nor UO_32 (O_32,N_18973,N_19755);
xnor UO_33 (O_33,N_17763,N_17452);
nor UO_34 (O_34,N_19050,N_17762);
or UO_35 (O_35,N_18533,N_17731);
xnor UO_36 (O_36,N_17973,N_19709);
and UO_37 (O_37,N_16417,N_18274);
and UO_38 (O_38,N_16572,N_19128);
and UO_39 (O_39,N_19606,N_17085);
nand UO_40 (O_40,N_18083,N_16467);
and UO_41 (O_41,N_18125,N_17023);
xnor UO_42 (O_42,N_19266,N_17954);
xnor UO_43 (O_43,N_18215,N_16933);
nor UO_44 (O_44,N_18187,N_19072);
nor UO_45 (O_45,N_19350,N_16359);
nand UO_46 (O_46,N_16775,N_17424);
xnor UO_47 (O_47,N_18887,N_18062);
nand UO_48 (O_48,N_19419,N_16367);
nand UO_49 (O_49,N_19915,N_16630);
xnor UO_50 (O_50,N_18332,N_17493);
nand UO_51 (O_51,N_19322,N_19877);
nor UO_52 (O_52,N_19717,N_16160);
xor UO_53 (O_53,N_16217,N_18862);
or UO_54 (O_54,N_18446,N_16910);
nor UO_55 (O_55,N_19073,N_16654);
or UO_56 (O_56,N_17134,N_16593);
nor UO_57 (O_57,N_16500,N_18289);
or UO_58 (O_58,N_16619,N_19301);
nor UO_59 (O_59,N_16325,N_17858);
or UO_60 (O_60,N_18270,N_16097);
nor UO_61 (O_61,N_19428,N_19117);
nand UO_62 (O_62,N_19513,N_16661);
and UO_63 (O_63,N_17550,N_18113);
nor UO_64 (O_64,N_16626,N_16682);
xor UO_65 (O_65,N_16270,N_18040);
xnor UO_66 (O_66,N_18701,N_16282);
or UO_67 (O_67,N_18799,N_18797);
nand UO_68 (O_68,N_19179,N_19499);
or UO_69 (O_69,N_19664,N_17951);
or UO_70 (O_70,N_17462,N_16816);
or UO_71 (O_71,N_19818,N_18144);
nand UO_72 (O_72,N_19054,N_17137);
or UO_73 (O_73,N_16382,N_18339);
nor UO_74 (O_74,N_16960,N_17817);
nand UO_75 (O_75,N_19302,N_16579);
and UO_76 (O_76,N_17190,N_16739);
nand UO_77 (O_77,N_17511,N_19342);
and UO_78 (O_78,N_16128,N_18285);
xnor UO_79 (O_79,N_18400,N_16698);
nand UO_80 (O_80,N_19510,N_17875);
and UO_81 (O_81,N_17124,N_18880);
nand UO_82 (O_82,N_16293,N_18947);
or UO_83 (O_83,N_18535,N_16237);
xor UO_84 (O_84,N_19662,N_17984);
and UO_85 (O_85,N_19477,N_17479);
xnor UO_86 (O_86,N_16923,N_19896);
nand UO_87 (O_87,N_19379,N_19246);
nand UO_88 (O_88,N_18127,N_19401);
and UO_89 (O_89,N_16837,N_18095);
nor UO_90 (O_90,N_16618,N_18952);
or UO_91 (O_91,N_19794,N_17755);
nor UO_92 (O_92,N_17420,N_16413);
and UO_93 (O_93,N_17135,N_16471);
nand UO_94 (O_94,N_16156,N_19198);
nand UO_95 (O_95,N_16198,N_19922);
and UO_96 (O_96,N_19337,N_16675);
xor UO_97 (O_97,N_18307,N_16348);
nor UO_98 (O_98,N_17172,N_19874);
nand UO_99 (O_99,N_19586,N_17055);
and UO_100 (O_100,N_18229,N_17429);
or UO_101 (O_101,N_19888,N_17997);
xnor UO_102 (O_102,N_19320,N_17696);
and UO_103 (O_103,N_17100,N_17434);
nand UO_104 (O_104,N_18935,N_18809);
or UO_105 (O_105,N_17760,N_16064);
and UO_106 (O_106,N_17197,N_18385);
and UO_107 (O_107,N_19905,N_17224);
and UO_108 (O_108,N_18741,N_19514);
or UO_109 (O_109,N_19677,N_16221);
or UO_110 (O_110,N_16006,N_19566);
nor UO_111 (O_111,N_16261,N_16748);
and UO_112 (O_112,N_19464,N_17451);
nor UO_113 (O_113,N_16704,N_17527);
and UO_114 (O_114,N_19753,N_16719);
xor UO_115 (O_115,N_19212,N_16290);
xor UO_116 (O_116,N_19207,N_16294);
nor UO_117 (O_117,N_18722,N_17320);
and UO_118 (O_118,N_18764,N_18825);
nand UO_119 (O_119,N_18146,N_19253);
nand UO_120 (O_120,N_19804,N_18734);
nand UO_121 (O_121,N_16818,N_17574);
and UO_122 (O_122,N_19775,N_17811);
nor UO_123 (O_123,N_19454,N_19567);
nor UO_124 (O_124,N_17708,N_19288);
or UO_125 (O_125,N_18247,N_19046);
nand UO_126 (O_126,N_18654,N_17611);
nand UO_127 (O_127,N_19036,N_18837);
or UO_128 (O_128,N_19112,N_17250);
nor UO_129 (O_129,N_17295,N_17482);
nor UO_130 (O_130,N_17421,N_17233);
nor UO_131 (O_131,N_18949,N_19822);
xor UO_132 (O_132,N_16875,N_17729);
nand UO_133 (O_133,N_16959,N_19007);
xor UO_134 (O_134,N_16756,N_18852);
and UO_135 (O_135,N_19258,N_18706);
or UO_136 (O_136,N_19704,N_17651);
or UO_137 (O_137,N_16078,N_17089);
xnor UO_138 (O_138,N_18528,N_16361);
or UO_139 (O_139,N_19745,N_17662);
or UO_140 (O_140,N_19434,N_16558);
or UO_141 (O_141,N_16977,N_17710);
xnor UO_142 (O_142,N_18908,N_18622);
nor UO_143 (O_143,N_18991,N_16125);
and UO_144 (O_144,N_19906,N_19810);
nand UO_145 (O_145,N_18064,N_19585);
nor UO_146 (O_146,N_17630,N_19359);
and UO_147 (O_147,N_18282,N_16208);
and UO_148 (O_148,N_17046,N_19427);
and UO_149 (O_149,N_16038,N_18733);
xor UO_150 (O_150,N_16200,N_18579);
nor UO_151 (O_151,N_19899,N_16355);
and UO_152 (O_152,N_17910,N_19172);
or UO_153 (O_153,N_16077,N_18896);
xnor UO_154 (O_154,N_17877,N_16055);
nor UO_155 (O_155,N_19319,N_16252);
nor UO_156 (O_156,N_17570,N_17258);
xnor UO_157 (O_157,N_19996,N_17075);
and UO_158 (O_158,N_18718,N_19307);
and UO_159 (O_159,N_17736,N_17854);
nor UO_160 (O_160,N_18865,N_16044);
xnor UO_161 (O_161,N_19315,N_18213);
and UO_162 (O_162,N_17423,N_17780);
or UO_163 (O_163,N_18618,N_17679);
and UO_164 (O_164,N_18473,N_19979);
and UO_165 (O_165,N_17706,N_16600);
nor UO_166 (O_166,N_18140,N_18814);
and UO_167 (O_167,N_17881,N_17924);
xor UO_168 (O_168,N_19402,N_16581);
nor UO_169 (O_169,N_19856,N_18931);
and UO_170 (O_170,N_16122,N_19821);
and UO_171 (O_171,N_19715,N_16984);
nor UO_172 (O_172,N_19913,N_17966);
nor UO_173 (O_173,N_18834,N_16142);
nand UO_174 (O_174,N_19332,N_18261);
nand UO_175 (O_175,N_19184,N_16114);
nor UO_176 (O_176,N_18665,N_18875);
or UO_177 (O_177,N_19750,N_18640);
nor UO_178 (O_178,N_17523,N_17602);
xnor UO_179 (O_179,N_16248,N_17412);
xor UO_180 (O_180,N_17562,N_19352);
xnor UO_181 (O_181,N_16988,N_16435);
and UO_182 (O_182,N_17983,N_18231);
xor UO_183 (O_183,N_18136,N_16819);
or UO_184 (O_184,N_18671,N_17834);
nor UO_185 (O_185,N_18027,N_17143);
or UO_186 (O_186,N_18675,N_17961);
and UO_187 (O_187,N_17388,N_16398);
nor UO_188 (O_188,N_19360,N_19440);
xor UO_189 (O_189,N_19958,N_16390);
or UO_190 (O_190,N_16281,N_18819);
nand UO_191 (O_191,N_19666,N_18178);
nand UO_192 (O_192,N_18917,N_18239);
xnor UO_193 (O_193,N_16475,N_19938);
nor UO_194 (O_194,N_16576,N_16342);
and UO_195 (O_195,N_16338,N_16950);
or UO_196 (O_196,N_16036,N_19059);
nand UO_197 (O_197,N_18101,N_19278);
nand UO_198 (O_198,N_18341,N_17601);
nand UO_199 (O_199,N_18266,N_17339);
and UO_200 (O_200,N_18905,N_16865);
nor UO_201 (O_201,N_18041,N_19578);
nand UO_202 (O_202,N_17119,N_17816);
nand UO_203 (O_203,N_19189,N_16147);
nor UO_204 (O_204,N_16166,N_19201);
nand UO_205 (O_205,N_18646,N_19960);
nor UO_206 (O_206,N_19767,N_16083);
or UO_207 (O_207,N_18070,N_19008);
xnor UO_208 (O_208,N_16955,N_17164);
or UO_209 (O_209,N_18333,N_16781);
and UO_210 (O_210,N_19948,N_18963);
or UO_211 (O_211,N_19972,N_16745);
or UO_212 (O_212,N_17664,N_16821);
and UO_213 (O_213,N_19752,N_17558);
xor UO_214 (O_214,N_19724,N_19761);
nand UO_215 (O_215,N_17363,N_17014);
nor UO_216 (O_216,N_16729,N_19837);
nand UO_217 (O_217,N_19762,N_19356);
xor UO_218 (O_218,N_16269,N_17489);
or UO_219 (O_219,N_18783,N_17317);
and UO_220 (O_220,N_16387,N_16673);
nor UO_221 (O_221,N_18563,N_19871);
or UO_222 (O_222,N_17199,N_17245);
or UO_223 (O_223,N_19030,N_17526);
xnor UO_224 (O_224,N_19230,N_19384);
xor UO_225 (O_225,N_17311,N_19543);
xor UO_226 (O_226,N_16770,N_17828);
and UO_227 (O_227,N_16250,N_18813);
and UO_228 (O_228,N_16872,N_18388);
nor UO_229 (O_229,N_17692,N_19719);
xnor UO_230 (O_230,N_16318,N_18707);
nor UO_231 (O_231,N_17605,N_16997);
nor UO_232 (O_232,N_16140,N_17627);
and UO_233 (O_233,N_17787,N_18780);
and UO_234 (O_234,N_17782,N_16645);
nand UO_235 (O_235,N_19568,N_16880);
xnor UO_236 (O_236,N_18796,N_17887);
or UO_237 (O_237,N_19475,N_18588);
nor UO_238 (O_238,N_17517,N_18773);
nor UO_239 (O_239,N_18141,N_18561);
xnor UO_240 (O_240,N_16468,N_16982);
or UO_241 (O_241,N_17348,N_18645);
nor UO_242 (O_242,N_16333,N_17458);
nor UO_243 (O_243,N_19718,N_19870);
nand UO_244 (O_244,N_16437,N_16498);
nand UO_245 (O_245,N_19701,N_19653);
xor UO_246 (O_246,N_17248,N_18928);
nor UO_247 (O_247,N_16920,N_17883);
xnor UO_248 (O_248,N_19492,N_18345);
xnor UO_249 (O_249,N_19261,N_16566);
xor UO_250 (O_250,N_17902,N_16515);
xnor UO_251 (O_251,N_16123,N_19576);
or UO_252 (O_252,N_18872,N_16194);
or UO_253 (O_253,N_17594,N_18445);
or UO_254 (O_254,N_16327,N_19965);
nor UO_255 (O_255,N_19303,N_18566);
or UO_256 (O_256,N_17112,N_19582);
xor UO_257 (O_257,N_16022,N_17370);
nor UO_258 (O_258,N_19010,N_17447);
nor UO_259 (O_259,N_19828,N_19618);
nand UO_260 (O_260,N_17730,N_18776);
xnor UO_261 (O_261,N_17196,N_17242);
or UO_262 (O_262,N_18444,N_18207);
nand UO_263 (O_263,N_16854,N_18740);
xor UO_264 (O_264,N_18135,N_19236);
nor UO_265 (O_265,N_16668,N_17278);
xnor UO_266 (O_266,N_18674,N_18256);
or UO_267 (O_267,N_19658,N_19150);
and UO_268 (O_268,N_16530,N_19561);
nand UO_269 (O_269,N_18382,N_19270);
xnor UO_270 (O_270,N_17147,N_17975);
nor UO_271 (O_271,N_18977,N_16922);
nand UO_272 (O_272,N_16518,N_17767);
xor UO_273 (O_273,N_18553,N_17425);
nor UO_274 (O_274,N_17484,N_16724);
xnor UO_275 (O_275,N_17025,N_19037);
xor UO_276 (O_276,N_17156,N_16430);
nand UO_277 (O_277,N_16953,N_19195);
and UO_278 (O_278,N_17290,N_17443);
xnor UO_279 (O_279,N_17274,N_17646);
nor UO_280 (O_280,N_16224,N_16786);
and UO_281 (O_281,N_16067,N_18903);
and UO_282 (O_282,N_19254,N_19945);
xor UO_283 (O_283,N_19846,N_19465);
nor UO_284 (O_284,N_17628,N_18591);
nand UO_285 (O_285,N_17437,N_18832);
nor UO_286 (O_286,N_17744,N_16007);
nand UO_287 (O_287,N_19646,N_17449);
nor UO_288 (O_288,N_17718,N_19408);
xor UO_289 (O_289,N_19487,N_18584);
or UO_290 (O_290,N_16278,N_17074);
nand UO_291 (O_291,N_19732,N_19305);
or UO_292 (O_292,N_16832,N_16642);
nor UO_293 (O_293,N_19854,N_19109);
xor UO_294 (O_294,N_18237,N_16732);
nor UO_295 (O_295,N_17230,N_16436);
nor UO_296 (O_296,N_18848,N_17827);
or UO_297 (O_297,N_17658,N_19101);
xor UO_298 (O_298,N_18606,N_19295);
nand UO_299 (O_299,N_19272,N_17486);
or UO_300 (O_300,N_19623,N_19389);
nor UO_301 (O_301,N_17386,N_18781);
or UO_302 (O_302,N_18719,N_17943);
or UO_303 (O_303,N_16517,N_18075);
xnor UO_304 (O_304,N_18004,N_17560);
nor UO_305 (O_305,N_18853,N_17715);
or UO_306 (O_306,N_17261,N_19610);
xor UO_307 (O_307,N_16415,N_16559);
xnor UO_308 (O_308,N_16641,N_19624);
xnor UO_309 (O_309,N_19240,N_19726);
nand UO_310 (O_310,N_18251,N_16439);
xnor UO_311 (O_311,N_19841,N_19622);
xor UO_312 (O_312,N_18313,N_16936);
nand UO_313 (O_313,N_18623,N_16629);
xnor UO_314 (O_314,N_16979,N_18936);
xnor UO_315 (O_315,N_16350,N_18620);
or UO_316 (O_316,N_17971,N_16890);
nand UO_317 (O_317,N_19100,N_17937);
nand UO_318 (O_318,N_16331,N_17537);
nand UO_319 (O_319,N_17422,N_19306);
xor UO_320 (O_320,N_19604,N_18396);
or UO_321 (O_321,N_19148,N_17071);
or UO_322 (O_322,N_17163,N_19080);
nor UO_323 (O_323,N_19262,N_19040);
and UO_324 (O_324,N_18463,N_16951);
or UO_325 (O_325,N_18731,N_17191);
and UO_326 (O_326,N_17592,N_16717);
nand UO_327 (O_327,N_16029,N_16551);
or UO_328 (O_328,N_16053,N_17192);
nor UO_329 (O_329,N_19633,N_19552);
xnor UO_330 (O_330,N_18192,N_17237);
xor UO_331 (O_331,N_16065,N_19006);
nand UO_332 (O_332,N_19243,N_19928);
nor UO_333 (O_333,N_16138,N_16608);
and UO_334 (O_334,N_17539,N_17144);
nand UO_335 (O_335,N_16042,N_16295);
nand UO_336 (O_336,N_16206,N_16349);
and UO_337 (O_337,N_18002,N_19636);
nor UO_338 (O_338,N_19489,N_16400);
nor UO_339 (O_339,N_18988,N_16190);
and UO_340 (O_340,N_17389,N_19515);
or UO_341 (O_341,N_19503,N_16279);
nor UO_342 (O_342,N_17205,N_18669);
xnor UO_343 (O_343,N_16856,N_17781);
and UO_344 (O_344,N_18039,N_19211);
nand UO_345 (O_345,N_16879,N_18715);
or UO_346 (O_346,N_16299,N_18200);
nand UO_347 (O_347,N_17958,N_18739);
nand UO_348 (O_348,N_18006,N_18211);
or UO_349 (O_349,N_16906,N_16560);
and UO_350 (O_350,N_18263,N_19819);
nor UO_351 (O_351,N_18492,N_17945);
nor UO_352 (O_352,N_19308,N_16392);
nand UO_353 (O_353,N_18937,N_16425);
nand UO_354 (O_354,N_17380,N_17228);
and UO_355 (O_355,N_17254,N_18594);
or UO_356 (O_356,N_17373,N_16362);
nor UO_357 (O_357,N_19770,N_19136);
or UO_358 (O_358,N_16481,N_18349);
xor UO_359 (O_359,N_16337,N_16738);
nor UO_360 (O_360,N_17035,N_17798);
nand UO_361 (O_361,N_19169,N_18712);
xnor UO_362 (O_362,N_19146,N_18688);
nand UO_363 (O_363,N_19500,N_18804);
xnor UO_364 (O_364,N_17117,N_17461);
or UO_365 (O_365,N_17717,N_17946);
nand UO_366 (O_366,N_17998,N_16179);
nor UO_367 (O_367,N_17207,N_19348);
xnor UO_368 (O_368,N_19480,N_16824);
and UO_369 (O_369,N_17917,N_16777);
xnor UO_370 (O_370,N_17243,N_16202);
xor UO_371 (O_371,N_19989,N_19197);
and UO_372 (O_372,N_19962,N_16961);
and UO_373 (O_373,N_16782,N_16864);
nand UO_374 (O_374,N_16374,N_16372);
nand UO_375 (O_375,N_16886,N_17822);
or UO_376 (O_376,N_16501,N_18012);
nand UO_377 (O_377,N_16177,N_18761);
nor UO_378 (O_378,N_16607,N_19868);
nand UO_379 (O_379,N_19678,N_17491);
nand UO_380 (O_380,N_19255,N_18507);
and UO_381 (O_381,N_17499,N_16148);
nor UO_382 (O_382,N_16182,N_18913);
nand UO_383 (O_383,N_16871,N_17530);
and UO_384 (O_384,N_17154,N_19882);
xor UO_385 (O_385,N_16175,N_18129);
and UO_386 (O_386,N_16954,N_18763);
xor UO_387 (O_387,N_16615,N_16525);
nor UO_388 (O_388,N_19079,N_17864);
nand UO_389 (O_389,N_17841,N_16469);
and UO_390 (O_390,N_19880,N_19035);
nand UO_391 (O_391,N_18234,N_18076);
nor UO_392 (O_392,N_17359,N_17857);
nor UO_393 (O_393,N_19759,N_19720);
and UO_394 (O_394,N_18369,N_16452);
and UO_395 (O_395,N_17302,N_18479);
nand UO_396 (O_396,N_19377,N_17528);
xor UO_397 (O_397,N_17064,N_19644);
nand UO_398 (O_398,N_19460,N_18241);
nor UO_399 (O_399,N_19092,N_16310);
nor UO_400 (O_400,N_19144,N_16344);
nand UO_401 (O_401,N_16754,N_16573);
and UO_402 (O_402,N_16227,N_18415);
xnor UO_403 (O_403,N_19527,N_16808);
nor UO_404 (O_404,N_16883,N_16456);
or UO_405 (O_405,N_19508,N_19923);
nand UO_406 (O_406,N_17923,N_18442);
nor UO_407 (O_407,N_16693,N_19991);
xnor UO_408 (O_408,N_18314,N_18893);
or UO_409 (O_409,N_19206,N_19438);
xnor UO_410 (O_410,N_19707,N_16284);
xnor UO_411 (O_411,N_18067,N_17698);
or UO_412 (O_412,N_18371,N_19312);
xor UO_413 (O_413,N_17474,N_16846);
xnor UO_414 (O_414,N_16575,N_17956);
nor UO_415 (O_415,N_18944,N_18421);
nand UO_416 (O_416,N_17897,N_16666);
nor UO_417 (O_417,N_18053,N_16080);
nand UO_418 (O_418,N_16800,N_19632);
or UO_419 (O_419,N_17500,N_17660);
or UO_420 (O_420,N_18166,N_19385);
nand UO_421 (O_421,N_19426,N_17603);
and UO_422 (O_422,N_18538,N_17070);
or UO_423 (O_423,N_18529,N_18704);
nor UO_424 (O_424,N_17695,N_17815);
xor UO_425 (O_425,N_17246,N_16408);
nand UO_426 (O_426,N_17765,N_18779);
and UO_427 (O_427,N_16924,N_18727);
and UO_428 (O_428,N_17073,N_16720);
nor UO_429 (O_429,N_16131,N_17039);
nand UO_430 (O_430,N_16655,N_19133);
nand UO_431 (O_431,N_18082,N_19069);
xor UO_432 (O_432,N_19713,N_19645);
nor UO_433 (O_433,N_18690,N_19479);
and UO_434 (O_434,N_19382,N_19192);
xnor UO_435 (O_435,N_17783,N_18248);
and UO_436 (O_436,N_16831,N_17195);
and UO_437 (O_437,N_16728,N_17079);
or UO_438 (O_438,N_18480,N_16368);
and UO_439 (O_439,N_17683,N_17082);
nand UO_440 (O_440,N_19075,N_18299);
and UO_441 (O_441,N_16111,N_16132);
nand UO_442 (O_442,N_18860,N_19990);
nand UO_443 (O_443,N_19224,N_18537);
nand UO_444 (O_444,N_16780,N_17145);
xnor UO_445 (O_445,N_19505,N_16921);
xor UO_446 (O_446,N_16519,N_17341);
nand UO_447 (O_447,N_18120,N_16448);
nor UO_448 (O_448,N_17271,N_16743);
or UO_449 (O_449,N_18593,N_19941);
nor UO_450 (O_450,N_19812,N_17059);
nand UO_451 (O_451,N_19534,N_16752);
nand UO_452 (O_452,N_16076,N_17090);
xnor UO_453 (O_453,N_18598,N_18162);
or UO_454 (O_454,N_19977,N_18985);
nand UO_455 (O_455,N_16366,N_19866);
nor UO_456 (O_456,N_16586,N_19916);
and UO_457 (O_457,N_19982,N_16894);
nor UO_458 (O_458,N_17553,N_16637);
xnor UO_459 (O_459,N_17688,N_19873);
or UO_460 (O_460,N_16735,N_19787);
xor UO_461 (O_461,N_18072,N_18115);
nand UO_462 (O_462,N_18504,N_17566);
nand UO_463 (O_463,N_18061,N_19765);
nand UO_464 (O_464,N_17991,N_17031);
nor UO_465 (O_465,N_16090,N_17356);
or UO_466 (O_466,N_18037,N_16426);
or UO_467 (O_467,N_18615,N_19226);
nand UO_468 (O_468,N_17432,N_16918);
or UO_469 (O_469,N_17616,N_18770);
and UO_470 (O_470,N_16696,N_16120);
xnor UO_471 (O_471,N_17166,N_17383);
and UO_472 (O_472,N_18794,N_18257);
nand UO_473 (O_473,N_18116,N_17277);
or UO_474 (O_474,N_19190,N_17175);
nor UO_475 (O_475,N_18871,N_17702);
xnor UO_476 (O_476,N_17534,N_19572);
xnor UO_477 (O_477,N_18567,N_16723);
or UO_478 (O_478,N_18544,N_16827);
xnor UO_479 (O_479,N_18922,N_18817);
xor UO_480 (O_480,N_16609,N_19691);
or UO_481 (O_481,N_18227,N_19797);
or UO_482 (O_482,N_16736,N_19956);
xor UO_483 (O_483,N_17315,N_18347);
or UO_484 (O_484,N_17270,N_18406);
xnor UO_485 (O_485,N_17149,N_17694);
and UO_486 (O_486,N_18830,N_17522);
or UO_487 (O_487,N_19242,N_18503);
or UO_488 (O_488,N_18753,N_16611);
or UO_489 (O_489,N_19887,N_18312);
nor UO_490 (O_490,N_19094,N_16940);
or UO_491 (O_491,N_17665,N_18452);
xor UO_492 (O_492,N_16676,N_18042);
nand UO_493 (O_493,N_17494,N_16971);
nor UO_494 (O_494,N_19672,N_19655);
or UO_495 (O_495,N_19469,N_19349);
nand UO_496 (O_496,N_18460,N_16058);
nand UO_497 (O_497,N_18110,N_18767);
nor UO_498 (O_498,N_16220,N_16590);
xor UO_499 (O_499,N_17814,N_19939);
nor UO_500 (O_500,N_16858,N_18447);
nand UO_501 (O_501,N_18358,N_16016);
nor UO_502 (O_502,N_17332,N_18549);
nor UO_503 (O_503,N_19039,N_16947);
and UO_504 (O_504,N_16761,N_17509);
or UO_505 (O_505,N_16212,N_18755);
nor UO_506 (O_506,N_17703,N_16725);
nand UO_507 (O_507,N_17818,N_19123);
nand UO_508 (O_508,N_17481,N_17467);
nand UO_509 (O_509,N_17298,N_19857);
or UO_510 (O_510,N_16601,N_19607);
nand UO_511 (O_511,N_17159,N_18630);
or UO_512 (O_512,N_19443,N_17774);
and UO_513 (O_513,N_19083,N_18164);
nand UO_514 (O_514,N_19921,N_17569);
and UO_515 (O_515,N_19931,N_17264);
xnor UO_516 (O_516,N_17282,N_17580);
nor UO_517 (O_517,N_18895,N_17789);
nor UO_518 (O_518,N_17641,N_19656);
and UO_519 (O_519,N_18353,N_16963);
xor UO_520 (O_520,N_19018,N_19187);
or UO_521 (O_521,N_18290,N_16215);
xor UO_522 (O_522,N_18610,N_19276);
and UO_523 (O_523,N_17027,N_19222);
or UO_524 (O_524,N_19642,N_19740);
nor UO_525 (O_525,N_17086,N_18225);
nor UO_526 (O_526,N_18417,N_16242);
xnor UO_527 (O_527,N_18010,N_19674);
nor UO_528 (O_528,N_19353,N_18425);
nand UO_529 (O_529,N_17889,N_17653);
or UO_530 (O_530,N_19626,N_19175);
or UO_531 (O_531,N_17846,N_17742);
and UO_532 (O_532,N_16214,N_18950);
xnor UO_533 (O_533,N_19089,N_16867);
nand UO_534 (O_534,N_19859,N_16839);
and UO_535 (O_535,N_17644,N_18490);
or UO_536 (O_536,N_19843,N_17165);
nor UO_537 (O_537,N_16035,N_18994);
and UO_538 (O_538,N_19327,N_19806);
or UO_539 (O_539,N_19194,N_16860);
or UO_540 (O_540,N_16153,N_19249);
nand UO_541 (O_541,N_19328,N_17726);
nor UO_542 (O_542,N_18638,N_16632);
nor UO_543 (O_543,N_19330,N_18250);
and UO_544 (O_544,N_16033,N_17426);
nand UO_545 (O_545,N_16779,N_17352);
nor UO_546 (O_546,N_18642,N_19529);
xnor UO_547 (O_547,N_18321,N_18291);
nor UO_548 (O_548,N_19934,N_18876);
and UO_549 (O_549,N_19217,N_19282);
nand UO_550 (O_550,N_19798,N_17680);
or UO_551 (O_551,N_17788,N_19612);
xor UO_552 (O_552,N_16239,N_17013);
and UO_553 (O_553,N_18016,N_17548);
xnor UO_554 (O_554,N_17138,N_17707);
nand UO_555 (O_555,N_18562,N_18293);
nand UO_556 (O_556,N_18468,N_17153);
xnor UO_557 (O_557,N_19394,N_17099);
nand UO_558 (O_558,N_16052,N_17049);
xnor UO_559 (O_559,N_16866,N_16185);
xor UO_560 (O_560,N_19901,N_19667);
nand UO_561 (O_561,N_18941,N_16695);
nand UO_562 (O_562,N_18574,N_17985);
nand UO_563 (O_563,N_18279,N_19894);
and UO_564 (O_564,N_19903,N_16913);
nand UO_565 (O_565,N_19041,N_19340);
and UO_566 (O_566,N_16434,N_19565);
nand UO_567 (O_567,N_18575,N_16323);
xor UO_568 (O_568,N_18081,N_18746);
nand UO_569 (O_569,N_17790,N_19984);
xor UO_570 (O_570,N_18278,N_16797);
or UO_571 (O_571,N_16291,N_19227);
xor UO_572 (O_572,N_17078,N_17127);
nand UO_573 (O_573,N_19453,N_17676);
nand UO_574 (O_574,N_19693,N_17588);
nor UO_575 (O_575,N_18769,N_19285);
nand UO_576 (O_576,N_17417,N_17371);
nand UO_577 (O_577,N_18978,N_17456);
and UO_578 (O_578,N_18451,N_18511);
or UO_579 (O_579,N_17252,N_19824);
xor UO_580 (O_580,N_18502,N_18975);
and UO_581 (O_581,N_17047,N_16211);
xor UO_582 (O_582,N_17850,N_19355);
nor UO_583 (O_583,N_18737,N_17612);
nand UO_584 (O_584,N_17606,N_16332);
and UO_585 (O_585,N_16130,N_16840);
and UO_586 (O_586,N_16550,N_19463);
and UO_587 (O_587,N_18856,N_16946);
nand UO_588 (O_588,N_18536,N_16714);
and UO_589 (O_589,N_16479,N_17871);
and UO_590 (O_590,N_19174,N_17992);
or UO_591 (O_591,N_18808,N_18703);
nand UO_592 (O_592,N_18326,N_17344);
xnor UO_593 (O_593,N_18276,N_17856);
and UO_594 (O_594,N_17610,N_18861);
nand UO_595 (O_595,N_18121,N_17459);
xor UO_596 (O_596,N_17336,N_17216);
and UO_597 (O_597,N_16183,N_17416);
or UO_598 (O_598,N_16127,N_18467);
and UO_599 (O_599,N_19685,N_16987);
or UO_600 (O_600,N_16934,N_17711);
nand UO_601 (O_601,N_18487,N_18132);
nand UO_602 (O_602,N_19605,N_18628);
nand UO_603 (O_603,N_17786,N_16021);
xnor UO_604 (O_604,N_19573,N_17977);
or UO_605 (O_605,N_17792,N_16911);
xor UO_606 (O_606,N_18288,N_18150);
nor UO_607 (O_607,N_19338,N_18629);
nor UO_608 (O_608,N_18017,N_19983);
and UO_609 (O_609,N_18992,N_16013);
xor UO_610 (O_610,N_16168,N_16313);
and UO_611 (O_611,N_19661,N_18891);
nand UO_612 (O_612,N_18375,N_18495);
and UO_613 (O_613,N_17648,N_19455);
nand UO_614 (O_614,N_16459,N_18676);
nand UO_615 (O_615,N_17880,N_17888);
or UO_616 (O_616,N_19879,N_19852);
or UO_617 (O_617,N_18028,N_18643);
nor UO_618 (O_618,N_19518,N_19738);
nor UO_619 (O_619,N_17269,N_18986);
or UO_620 (O_620,N_17549,N_17771);
or UO_621 (O_621,N_19466,N_17939);
nand UO_622 (O_622,N_16395,N_18998);
nand UO_623 (O_623,N_17777,N_18325);
or UO_624 (O_624,N_18366,N_16107);
nand UO_625 (O_625,N_18523,N_18683);
or UO_626 (O_626,N_18238,N_19629);
nand UO_627 (O_627,N_18580,N_16859);
xnor UO_628 (O_628,N_18906,N_17773);
and UO_629 (O_629,N_19925,N_16336);
or UO_630 (O_630,N_18934,N_16635);
xor UO_631 (O_631,N_17309,N_18864);
nor UO_632 (O_632,N_17360,N_18576);
or UO_633 (O_633,N_17043,N_17305);
nor UO_634 (O_634,N_19005,N_16765);
or UO_635 (O_635,N_18221,N_19009);
nand UO_636 (O_636,N_16945,N_19432);
nor UO_637 (O_637,N_17669,N_19373);
and UO_638 (O_638,N_17533,N_18641);
or UO_639 (O_639,N_19641,N_19801);
or UO_640 (O_640,N_19271,N_19875);
nor UO_641 (O_641,N_19292,N_17019);
nor UO_642 (O_642,N_16126,N_17041);
nand UO_643 (O_643,N_17395,N_16788);
nand UO_644 (O_644,N_17929,N_19814);
nand UO_645 (O_645,N_19025,N_16397);
nand UO_646 (O_646,N_17044,N_19178);
nor UO_647 (O_647,N_16589,N_16730);
nand UO_648 (O_648,N_18253,N_17620);
nand UO_649 (O_649,N_17919,N_16210);
or UO_650 (O_650,N_19688,N_19933);
nand UO_651 (O_651,N_16431,N_19289);
and UO_652 (O_652,N_16778,N_17675);
nor UO_653 (O_653,N_18438,N_18659);
nor UO_654 (O_654,N_19097,N_19748);
xor UO_655 (O_655,N_17684,N_17564);
and UO_656 (O_656,N_18590,N_18923);
and UO_657 (O_657,N_18569,N_16539);
nand UO_658 (O_658,N_17775,N_16553);
or UO_659 (O_659,N_16050,N_17376);
nor UO_660 (O_660,N_17624,N_17621);
nand UO_661 (O_661,N_19002,N_18577);
and UO_662 (O_662,N_19530,N_17281);
and UO_663 (O_663,N_16917,N_17345);
xor UO_664 (O_664,N_16223,N_19853);
and UO_665 (O_665,N_16843,N_16810);
nor UO_666 (O_666,N_19722,N_16944);
nor UO_667 (O_667,N_17812,N_17287);
xnor UO_668 (O_668,N_19725,N_19537);
and UO_669 (O_669,N_16300,N_16203);
or UO_670 (O_670,N_16137,N_17745);
nor UO_671 (O_671,N_19531,N_18664);
or UO_672 (O_672,N_16432,N_16699);
xnor UO_673 (O_673,N_17239,N_16238);
and UO_674 (O_674,N_17565,N_18499);
and UO_675 (O_675,N_19751,N_18143);
or UO_676 (O_676,N_18160,N_18034);
xor UO_677 (O_677,N_19670,N_19878);
xor UO_678 (O_678,N_17931,N_16081);
nand UO_679 (O_679,N_17844,N_17327);
xnor UO_680 (O_680,N_16549,N_17949);
nand UO_681 (O_681,N_16893,N_18699);
xnor UO_682 (O_682,N_18106,N_17903);
or UO_683 (O_683,N_18653,N_16297);
nor UO_684 (O_684,N_18692,N_17795);
nor UO_685 (O_685,N_19838,N_16633);
nor UO_686 (O_686,N_16254,N_19176);
xor UO_687 (O_687,N_16257,N_17503);
nand UO_688 (O_688,N_16674,N_16529);
or UO_689 (O_689,N_19032,N_17979);
nor UO_690 (O_690,N_19202,N_17623);
nor UO_691 (O_691,N_16667,N_17353);
nand UO_692 (O_692,N_17608,N_18652);
nor UO_693 (O_693,N_16445,N_18525);
nand UO_694 (O_694,N_17797,N_19203);
nor UO_695 (O_695,N_18328,N_16353);
xor UO_696 (O_696,N_17920,N_17993);
or UO_697 (O_697,N_17194,N_17567);
nand UO_698 (O_698,N_19056,N_18810);
and UO_699 (O_699,N_17512,N_16188);
xnor UO_700 (O_700,N_19119,N_18782);
and UO_701 (O_701,N_16186,N_17379);
nand UO_702 (O_702,N_17415,N_16079);
or UO_703 (O_703,N_16030,N_18365);
or UO_704 (O_704,N_16707,N_16195);
nand UO_705 (O_705,N_16545,N_19540);
nand UO_706 (O_706,N_18940,N_18329);
xor UO_707 (O_707,N_19022,N_18530);
xnor UO_708 (O_708,N_17712,N_18305);
nand UO_709 (O_709,N_17544,N_16213);
xnor UO_710 (O_710,N_17994,N_17211);
or UO_711 (O_711,N_18777,N_19162);
nor UO_712 (O_712,N_19391,N_17738);
xor UO_713 (O_713,N_19140,N_18874);
or UO_714 (O_714,N_19027,N_16454);
or UO_715 (O_715,N_17105,N_17377);
xor UO_716 (O_716,N_17151,N_18398);
nor UO_717 (O_717,N_16621,N_18020);
or UO_718 (O_718,N_19949,N_17735);
or UO_719 (O_719,N_19232,N_17328);
xnor UO_720 (O_720,N_16204,N_18748);
xor UO_721 (O_721,N_19742,N_19538);
nand UO_722 (O_722,N_17036,N_19425);
or UO_723 (O_723,N_18156,N_17334);
or UO_724 (O_724,N_17898,N_19017);
nand UO_725 (O_725,N_19012,N_19157);
xnor UO_726 (O_726,N_18175,N_18043);
and UO_727 (O_727,N_18286,N_17338);
xor UO_728 (O_728,N_19105,N_19850);
and UO_729 (O_729,N_19548,N_18682);
and UO_730 (O_730,N_19114,N_19219);
xnor UO_731 (O_731,N_18392,N_17419);
nand UO_732 (O_732,N_18431,N_17092);
and UO_733 (O_733,N_17823,N_19214);
or UO_734 (O_734,N_17468,N_19665);
or UO_735 (O_735,N_19652,N_19544);
xor UO_736 (O_736,N_17106,N_17142);
xor UO_737 (O_737,N_19731,N_19439);
nand UO_738 (O_738,N_16105,N_16027);
and UO_739 (O_739,N_18194,N_16230);
or UO_740 (O_740,N_19608,N_18785);
or UO_741 (O_741,N_18693,N_18159);
nand UO_742 (O_742,N_18139,N_16656);
nor UO_743 (O_743,N_17123,N_16993);
nor UO_744 (O_744,N_18203,N_18190);
xor UO_745 (O_745,N_18472,N_17870);
and UO_746 (O_746,N_16341,N_18724);
nand UO_747 (O_747,N_17693,N_19216);
nand UO_748 (O_748,N_18252,N_16315);
or UO_749 (O_749,N_16312,N_17859);
or UO_750 (O_750,N_17942,N_17837);
and UO_751 (O_751,N_16427,N_17475);
xor UO_752 (O_752,N_18306,N_18605);
xnor UO_753 (O_753,N_17617,N_18259);
or UO_754 (O_754,N_17582,N_19525);
nand UO_755 (O_755,N_17541,N_16822);
and UO_756 (O_756,N_18055,N_19339);
nand UO_757 (O_757,N_16952,N_18210);
xnor UO_758 (O_758,N_19397,N_18344);
nand UO_759 (O_759,N_16370,N_17705);
nor UO_760 (O_760,N_16897,N_19260);
nand UO_761 (O_761,N_19867,N_16989);
nor UO_762 (O_762,N_17972,N_16264);
nor UO_763 (O_763,N_18077,N_19690);
nand UO_764 (O_764,N_17759,N_19924);
or UO_765 (O_765,N_18901,N_19792);
nand UO_766 (O_766,N_17508,N_16749);
and UO_767 (O_767,N_17847,N_19603);
xor UO_768 (O_768,N_16892,N_18768);
nand UO_769 (O_769,N_19834,N_17869);
nand UO_770 (O_770,N_19003,N_17179);
nand UO_771 (O_771,N_16753,N_18021);
xor UO_772 (O_772,N_16000,N_19526);
or UO_773 (O_773,N_17739,N_18283);
nand UO_774 (O_774,N_19329,N_16196);
nand UO_775 (O_775,N_17095,N_17026);
or UO_776 (O_776,N_16412,N_16552);
nor UO_777 (O_777,N_19829,N_16610);
xor UO_778 (O_778,N_19844,N_17136);
or UO_779 (O_779,N_17203,N_18619);
xor UO_780 (O_780,N_17586,N_16145);
nor UO_781 (O_781,N_18368,N_16904);
nor UO_782 (O_782,N_17982,N_17368);
nor UO_783 (O_783,N_17853,N_17178);
nor UO_784 (O_784,N_18754,N_16565);
nand UO_785 (O_785,N_16173,N_19619);
and UO_786 (O_786,N_17051,N_17185);
or UO_787 (O_787,N_16708,N_17120);
nand UO_788 (O_788,N_18705,N_19196);
and UO_789 (O_789,N_19864,N_17146);
nor UO_790 (O_790,N_17155,N_16862);
xor UO_791 (O_791,N_17749,N_18352);
nor UO_792 (O_792,N_19199,N_16014);
and UO_793 (O_793,N_18510,N_16491);
xor UO_794 (O_794,N_16497,N_18054);
and UO_795 (O_795,N_17643,N_17758);
nor UO_796 (O_796,N_19815,N_18868);
xnor UO_797 (O_797,N_16228,N_19121);
xor UO_798 (O_798,N_17672,N_19365);
or UO_799 (O_799,N_18596,N_18802);
or UO_800 (O_800,N_16722,N_18614);
and UO_801 (O_801,N_19154,N_16170);
and UO_802 (O_802,N_18050,N_19237);
or UO_803 (O_803,N_19997,N_16889);
or UO_804 (O_804,N_16460,N_16371);
and UO_805 (O_805,N_17184,N_18459);
or UO_806 (O_806,N_19793,N_16978);
nand UO_807 (O_807,N_16373,N_19145);
nand UO_808 (O_808,N_16931,N_19647);
nand UO_809 (O_809,N_16419,N_17935);
nand UO_810 (O_810,N_17122,N_19430);
and UO_811 (O_811,N_16935,N_19457);
or UO_812 (O_812,N_16829,N_18242);
nor UO_813 (O_813,N_16825,N_17953);
nand UO_814 (O_814,N_19895,N_16259);
or UO_815 (O_815,N_18240,N_17657);
or UO_816 (O_816,N_16181,N_17914);
nand UO_817 (O_817,N_18246,N_16512);
nor UO_818 (O_818,N_16158,N_17303);
nand UO_819 (O_819,N_18501,N_19433);
nand UO_820 (O_820,N_16260,N_18532);
or UO_821 (O_821,N_18617,N_19115);
nand UO_822 (O_822,N_16602,N_19218);
xnor UO_823 (O_823,N_18713,N_19836);
nor UO_824 (O_824,N_16303,N_16751);
nor UO_825 (O_825,N_18354,N_17232);
nand UO_826 (O_826,N_17206,N_17034);
or UO_827 (O_827,N_17408,N_17714);
xor UO_828 (O_828,N_17125,N_19366);
and UO_829 (O_829,N_16820,N_19914);
or UO_830 (O_830,N_16874,N_18205);
xnor UO_831 (O_831,N_16804,N_17001);
xnor UO_832 (O_832,N_16234,N_17825);
and UO_833 (O_833,N_16174,N_18414);
nor UO_834 (O_834,N_19648,N_17810);
or UO_835 (O_835,N_18486,N_16791);
xnor UO_836 (O_836,N_16772,N_17289);
nand UO_837 (O_837,N_19418,N_17600);
or UO_838 (O_838,N_16991,N_18822);
or UO_839 (O_839,N_17959,N_17634);
nand UO_840 (O_840,N_16154,N_17860);
nor UO_841 (O_841,N_19141,N_19737);
nand UO_842 (O_842,N_18989,N_18338);
and UO_843 (O_843,N_17284,N_19287);
and UO_844 (O_844,N_19085,N_18334);
nand UO_845 (O_845,N_19456,N_18811);
or UO_846 (O_846,N_16161,N_17091);
xor UO_847 (O_847,N_19951,N_19595);
xor UO_848 (O_848,N_17162,N_19331);
xnor UO_849 (O_849,N_17193,N_16841);
xnor UO_850 (O_850,N_17892,N_16354);
nand UO_851 (O_851,N_16746,N_17724);
or UO_852 (O_852,N_17504,N_19679);
and UO_853 (O_853,N_17396,N_17335);
or UO_854 (O_854,N_18886,N_16329);
nor UO_855 (O_855,N_17448,N_19346);
nor UO_856 (O_856,N_16759,N_19476);
and UO_857 (O_857,N_19351,N_16251);
nor UO_858 (O_858,N_19723,N_17776);
and UO_859 (O_859,N_17746,N_17351);
or UO_860 (O_860,N_16143,N_16162);
xnor UO_861 (O_861,N_19926,N_16657);
and UO_862 (O_862,N_16863,N_19733);
nand UO_863 (O_863,N_16851,N_19152);
nand UO_864 (O_864,N_18104,N_16084);
or UO_865 (O_865,N_18957,N_16253);
nor UO_866 (O_866,N_18331,N_19504);
xor UO_867 (O_867,N_19889,N_17655);
xor UO_868 (O_868,N_17909,N_19885);
and UO_869 (O_869,N_18087,N_16998);
or UO_870 (O_870,N_18910,N_17032);
nand UO_871 (O_871,N_17756,N_18478);
or UO_872 (O_872,N_19630,N_18543);
or UO_873 (O_873,N_18176,N_19992);
xnor UO_874 (O_874,N_16702,N_16358);
xnor UO_875 (O_875,N_18735,N_18264);
nand UO_876 (O_876,N_19378,N_18778);
and UO_877 (O_877,N_19961,N_19291);
or UO_878 (O_878,N_18476,N_16010);
nand UO_879 (O_879,N_16606,N_17670);
nor UO_880 (O_880,N_17097,N_16243);
nand UO_881 (O_881,N_18838,N_19985);
nand UO_882 (O_882,N_18046,N_18484);
and UO_883 (O_883,N_17839,N_19754);
or UO_884 (O_884,N_17210,N_16690);
or UO_885 (O_885,N_16533,N_18114);
nand UO_886 (O_886,N_17563,N_19865);
xnor UO_887 (O_887,N_19728,N_16442);
or UO_888 (O_888,N_17952,N_16218);
nor UO_889 (O_889,N_18546,N_17213);
xor UO_890 (O_890,N_18117,N_18840);
xnor UO_891 (O_891,N_16784,N_19311);
or UO_892 (O_892,N_17171,N_19193);
nor UO_893 (O_893,N_17940,N_17573);
or UO_894 (O_894,N_16246,N_17219);
xnor UO_895 (O_895,N_19516,N_18806);
xnor UO_896 (O_896,N_17081,N_17470);
and UO_897 (O_897,N_19170,N_18774);
xnor UO_898 (O_898,N_16396,N_16965);
nor UO_899 (O_899,N_19575,N_16034);
nand UO_900 (O_900,N_16726,N_16658);
and UO_901 (O_901,N_16510,N_16104);
nor UO_902 (O_902,N_17296,N_19234);
nor UO_903 (O_903,N_18520,N_19393);
or UO_904 (O_904,N_19068,N_18686);
nand UO_905 (O_905,N_16915,N_16085);
and UO_906 (O_906,N_16473,N_18943);
or UO_907 (O_907,N_18926,N_19028);
or UO_908 (O_908,N_17599,N_16731);
or UO_909 (O_909,N_16496,N_17632);
or UO_910 (O_910,N_17804,N_16477);
nor UO_911 (O_911,N_18235,N_16015);
nand UO_912 (O_912,N_17325,N_17686);
nor UO_913 (O_913,N_19406,N_17899);
or UO_914 (O_914,N_17990,N_19833);
xnor UO_915 (O_915,N_16937,N_19876);
or UO_916 (O_916,N_19519,N_16285);
or UO_917 (O_917,N_17280,N_17240);
nand UO_918 (O_918,N_17244,N_17331);
or UO_919 (O_919,N_16705,N_19478);
and UO_920 (O_920,N_18599,N_19238);
xor UO_921 (O_921,N_19051,N_16180);
nor UO_922 (O_922,N_19367,N_19545);
xnor UO_923 (O_923,N_16830,N_17806);
nand UO_924 (O_924,N_16681,N_18539);
and UO_925 (O_925,N_19138,N_16793);
and UO_926 (O_926,N_17989,N_19256);
nand UO_927 (O_927,N_19422,N_18587);
nand UO_928 (O_928,N_18929,N_19768);
and UO_929 (O_929,N_17614,N_19459);
and UO_930 (O_930,N_17852,N_17831);
and UO_931 (O_931,N_18695,N_16899);
nand UO_932 (O_932,N_17513,N_16541);
and UO_933 (O_933,N_16263,N_19317);
nor UO_934 (O_934,N_19564,N_17501);
and UO_935 (O_935,N_16178,N_19786);
nor UO_936 (O_936,N_19437,N_19580);
or UO_937 (O_937,N_17687,N_18982);
or UO_938 (O_938,N_19103,N_17631);
and UO_939 (O_939,N_16402,N_16288);
or UO_940 (O_940,N_18416,N_16429);
and UO_941 (O_941,N_18854,N_19462);
and UO_942 (O_942,N_19120,N_18255);
nor UO_943 (O_943,N_17366,N_17540);
nand UO_944 (O_944,N_18968,N_17008);
nor UO_945 (O_945,N_18531,N_18609);
nor UO_946 (O_946,N_19592,N_18829);
nand UO_947 (O_947,N_17796,N_16669);
and UO_948 (O_948,N_16634,N_17042);
xor UO_949 (O_949,N_19182,N_16046);
or UO_950 (O_950,N_19886,N_16789);
nor UO_951 (O_951,N_17087,N_19596);
nor UO_952 (O_952,N_19869,N_19163);
or UO_953 (O_953,N_16847,N_19695);
nand UO_954 (O_954,N_19049,N_18558);
nand UO_955 (O_955,N_17260,N_16919);
xnor UO_956 (O_956,N_19727,N_18346);
nor UO_957 (O_957,N_19987,N_16592);
nor UO_958 (O_958,N_19791,N_16405);
nand UO_959 (O_959,N_16941,N_18049);
or UO_960 (O_960,N_17807,N_16741);
or UO_961 (O_961,N_18795,N_17364);
and UO_962 (O_962,N_16149,N_16713);
and UO_963 (O_963,N_19493,N_18066);
or UO_964 (O_964,N_16433,N_16464);
nand UO_965 (O_965,N_16591,N_18138);
nand UO_966 (O_966,N_17571,N_19813);
nor UO_967 (O_967,N_16271,N_17446);
or UO_968 (O_968,N_18336,N_19057);
nor UO_969 (O_969,N_18647,N_16176);
or UO_970 (O_970,N_18743,N_18350);
or UO_971 (O_971,N_19597,N_16199);
nor UO_972 (O_972,N_17842,N_18919);
xnor UO_973 (O_973,N_19344,N_17052);
or UO_974 (O_974,N_19563,N_17161);
nor UO_975 (O_975,N_17590,N_17401);
and UO_976 (O_976,N_17908,N_18634);
or UO_977 (O_977,N_17697,N_16031);
xor UO_978 (O_978,N_16470,N_17109);
xnor UO_979 (O_979,N_18663,N_17699);
or UO_980 (O_980,N_16636,N_19047);
and UO_981 (O_981,N_17598,N_18925);
nor UO_982 (O_982,N_18031,N_19065);
or UO_983 (O_983,N_18033,N_16680);
and UO_984 (O_984,N_17128,N_17800);
or UO_985 (O_985,N_18666,N_16144);
and UO_986 (O_986,N_18262,N_16828);
nor UO_987 (O_987,N_18044,N_18884);
nor UO_988 (O_988,N_18086,N_17668);
nor UO_989 (O_989,N_18624,N_16562);
and UO_990 (O_990,N_18927,N_19142);
and UO_991 (O_991,N_18668,N_16535);
nand UO_992 (O_992,N_18541,N_17673);
or UO_993 (O_993,N_17283,N_16386);
nand UO_994 (O_994,N_18820,N_17113);
or UO_995 (O_995,N_16833,N_16683);
xnor UO_996 (O_996,N_17445,N_17033);
and UO_997 (O_997,N_17868,N_18003);
and UO_998 (O_998,N_19490,N_19920);
xor UO_999 (O_999,N_16888,N_17932);
nand UO_1000 (O_1000,N_18602,N_17394);
and UO_1001 (O_1001,N_16375,N_16805);
and UO_1002 (O_1002,N_16556,N_19705);
and UO_1003 (O_1003,N_18245,N_19964);
nor UO_1004 (O_1004,N_16106,N_18024);
xor UO_1005 (O_1005,N_18157,N_16785);
xnor UO_1006 (O_1006,N_19204,N_16506);
nand UO_1007 (O_1007,N_18454,N_18681);
or UO_1008 (O_1008,N_17374,N_17532);
xor UO_1009 (O_1009,N_19802,N_17126);
or UO_1010 (O_1010,N_19364,N_18660);
nor UO_1011 (O_1011,N_17876,N_18920);
xor UO_1012 (O_1012,N_19407,N_18191);
xnor UO_1013 (O_1013,N_18470,N_18716);
xnor UO_1014 (O_1014,N_19250,N_18090);
nor UO_1015 (O_1015,N_19957,N_19808);
nor UO_1016 (O_1016,N_19774,N_17413);
nand UO_1017 (O_1017,N_18677,N_17300);
nor UO_1018 (O_1018,N_16340,N_19269);
nand UO_1019 (O_1019,N_19078,N_17633);
or UO_1020 (O_1020,N_19975,N_16438);
nor UO_1021 (O_1021,N_19782,N_16848);
and UO_1022 (O_1022,N_18397,N_17346);
and UO_1023 (O_1023,N_16852,N_17176);
and UO_1024 (O_1024,N_18035,N_17257);
or UO_1025 (O_1025,N_18001,N_18885);
or UO_1026 (O_1026,N_17682,N_17157);
nor UO_1027 (O_1027,N_16887,N_16538);
or UO_1028 (O_1028,N_18174,N_17618);
nor UO_1029 (O_1029,N_18373,N_18409);
or UO_1030 (O_1030,N_19106,N_16458);
nand UO_1031 (O_1031,N_18651,N_17649);
nor UO_1032 (O_1032,N_18009,N_17160);
xnor UO_1033 (O_1033,N_16171,N_19790);
or UO_1034 (O_1034,N_19000,N_19682);
or UO_1035 (O_1035,N_18993,N_19412);
and UO_1036 (O_1036,N_16399,N_19014);
or UO_1037 (O_1037,N_18457,N_17535);
xor UO_1038 (O_1038,N_18866,N_19533);
xnor UO_1039 (O_1039,N_18980,N_18635);
nor UO_1040 (O_1040,N_18303,N_18226);
nor UO_1041 (O_1041,N_17251,N_19669);
nor UO_1042 (O_1042,N_18514,N_18327);
or UO_1043 (O_1043,N_18534,N_19313);
nand UO_1044 (O_1044,N_18984,N_17733);
nand UO_1045 (O_1045,N_16505,N_16764);
nor UO_1046 (O_1046,N_17799,N_17716);
nand UO_1047 (O_1047,N_17555,N_16546);
xor UO_1048 (O_1048,N_16973,N_16554);
xnor UO_1049 (O_1049,N_18163,N_18124);
nor UO_1050 (O_1050,N_18233,N_17480);
and UO_1051 (O_1051,N_19832,N_17222);
xor UO_1052 (O_1052,N_16466,N_18137);
nor UO_1053 (O_1053,N_16139,N_17202);
nor UO_1054 (O_1054,N_18185,N_17721);
or UO_1055 (O_1055,N_19274,N_16074);
xnor UO_1056 (O_1056,N_17821,N_19074);
and UO_1057 (O_1057,N_19796,N_17701);
nor UO_1058 (O_1058,N_19343,N_19372);
and UO_1059 (O_1059,N_17967,N_17150);
nor UO_1060 (O_1060,N_16706,N_18933);
nor UO_1061 (O_1061,N_16092,N_16073);
or UO_1062 (O_1062,N_17319,N_16037);
and UO_1063 (O_1063,N_18381,N_17167);
xor UO_1064 (O_1064,N_16424,N_17988);
xnor UO_1065 (O_1065,N_16141,N_16388);
or UO_1066 (O_1066,N_17659,N_16564);
xnor UO_1067 (O_1067,N_19033,N_19708);
xnor UO_1068 (O_1068,N_18873,N_16222);
and UO_1069 (O_1069,N_16060,N_17652);
or UO_1070 (O_1070,N_17441,N_19341);
nor UO_1071 (O_1071,N_17297,N_16603);
xnor UO_1072 (O_1072,N_16209,N_16742);
or UO_1073 (O_1073,N_16845,N_19588);
and UO_1074 (O_1074,N_17879,N_17262);
nor UO_1075 (O_1075,N_17543,N_19011);
nor UO_1076 (O_1076,N_16157,N_19692);
xnor UO_1077 (O_1077,N_19347,N_16440);
xor UO_1078 (O_1078,N_16100,N_16110);
xnor UO_1079 (O_1079,N_18556,N_18360);
xnor UO_1080 (O_1080,N_19910,N_18912);
nand UO_1081 (O_1081,N_19835,N_19823);
nand UO_1082 (O_1082,N_19358,N_16612);
nand UO_1083 (O_1083,N_16363,N_19942);
and UO_1084 (O_1084,N_18005,N_19706);
and UO_1085 (O_1085,N_16051,N_16975);
nor UO_1086 (O_1086,N_19228,N_18505);
xnor UO_1087 (O_1087,N_16346,N_18655);
or UO_1088 (O_1088,N_19416,N_17204);
nand UO_1089 (O_1089,N_18224,N_19651);
xor UO_1090 (O_1090,N_18209,N_18843);
nor UO_1091 (O_1091,N_19370,N_18377);
nand UO_1092 (O_1092,N_16811,N_16651);
xor UO_1093 (O_1093,N_17750,N_16309);
nor UO_1094 (O_1094,N_16001,N_17813);
and UO_1095 (O_1095,N_19998,N_17546);
nor UO_1096 (O_1096,N_19686,N_16514);
nor UO_1097 (O_1097,N_16908,N_17866);
and UO_1098 (O_1098,N_16787,N_19281);
xnor UO_1099 (O_1099,N_19988,N_17053);
xor UO_1100 (O_1100,N_16351,N_19800);
nor UO_1101 (O_1101,N_18060,N_17554);
xor UO_1102 (O_1102,N_19273,N_18384);
nor UO_1103 (O_1103,N_16275,N_17720);
xnor UO_1104 (O_1104,N_16929,N_19244);
and UO_1105 (O_1105,N_18702,N_18842);
or UO_1106 (O_1106,N_18608,N_16472);
nor UO_1107 (O_1107,N_17515,N_17904);
nor UO_1108 (O_1108,N_18218,N_18171);
and UO_1109 (O_1109,N_18551,N_17116);
nor UO_1110 (O_1110,N_18603,N_17350);
or UO_1111 (O_1111,N_17102,N_19569);
or UO_1112 (O_1112,N_18845,N_19293);
or UO_1113 (O_1113,N_17018,N_16694);
and UO_1114 (O_1114,N_17609,N_16484);
or UO_1115 (O_1115,N_19799,N_19590);
xnor UO_1116 (O_1116,N_18023,N_17385);
nand UO_1117 (O_1117,N_16462,N_19777);
and UO_1118 (O_1118,N_16002,N_18222);
and UO_1119 (O_1119,N_16849,N_18889);
nand UO_1120 (O_1120,N_16733,N_18775);
and UO_1121 (O_1121,N_19936,N_18869);
or UO_1122 (O_1122,N_18310,N_19264);
or UO_1123 (O_1123,N_19550,N_16317);
xnor UO_1124 (O_1124,N_16870,N_18199);
or UO_1125 (O_1125,N_17476,N_17901);
and UO_1126 (O_1126,N_16306,N_16595);
and UO_1127 (O_1127,N_19820,N_16968);
nor UO_1128 (O_1128,N_18111,N_17174);
nand UO_1129 (O_1129,N_19093,N_16983);
nor UO_1130 (O_1130,N_18679,N_18496);
xnor UO_1131 (O_1131,N_18542,N_17058);
or UO_1132 (O_1132,N_17483,N_17182);
nand UO_1133 (O_1133,N_16684,N_18254);
or UO_1134 (O_1134,N_18038,N_19334);
and UO_1135 (O_1135,N_17354,N_17030);
nor UO_1136 (O_1136,N_18877,N_18742);
and UO_1137 (O_1137,N_19435,N_17557);
and UO_1138 (O_1138,N_18721,N_16643);
xnor UO_1139 (O_1139,N_16189,N_16796);
nand UO_1140 (O_1140,N_18098,N_19413);
nor UO_1141 (O_1141,N_19165,N_17186);
and UO_1142 (O_1142,N_16962,N_18122);
xnor UO_1143 (O_1143,N_19898,N_19918);
xnor UO_1144 (O_1144,N_16457,N_19700);
nand UO_1145 (O_1145,N_16534,N_16094);
nor UO_1146 (O_1146,N_16853,N_16191);
nor UO_1147 (O_1147,N_19491,N_18841);
or UO_1148 (O_1148,N_17531,N_19076);
nand UO_1149 (O_1149,N_18330,N_17832);
and UO_1150 (O_1150,N_17265,N_18045);
xnor UO_1151 (O_1151,N_18571,N_17893);
nand UO_1152 (O_1152,N_17576,N_17613);
xnor UO_1153 (O_1153,N_16403,N_16274);
and UO_1154 (O_1154,N_19268,N_17238);
nand UO_1155 (O_1155,N_18626,N_16755);
xor UO_1156 (O_1156,N_18942,N_18342);
xnor UO_1157 (O_1157,N_18402,N_16536);
nor UO_1158 (O_1158,N_18308,N_18759);
xor UO_1159 (O_1159,N_16776,N_17622);
xor UO_1160 (O_1160,N_16734,N_16072);
xnor UO_1161 (O_1161,N_18161,N_18548);
or UO_1162 (O_1162,N_16101,N_17212);
nor UO_1163 (O_1163,N_16009,N_18394);
and UO_1164 (O_1164,N_19004,N_18188);
and UO_1165 (O_1165,N_19712,N_19721);
xor UO_1166 (O_1166,N_16596,N_16134);
xnor UO_1167 (O_1167,N_16305,N_19599);
xor UO_1168 (O_1168,N_18198,N_16794);
nand UO_1169 (O_1169,N_16411,N_19486);
nor UO_1170 (O_1170,N_19969,N_17748);
nand UO_1171 (O_1171,N_18186,N_16769);
xor UO_1172 (O_1172,N_19286,N_16011);
nor UO_1173 (O_1173,N_16262,N_17259);
and UO_1174 (O_1174,N_18430,N_16061);
nor UO_1175 (O_1175,N_16994,N_18757);
or UO_1176 (O_1176,N_17820,N_16115);
xor UO_1177 (O_1177,N_18196,N_17478);
nor UO_1178 (O_1178,N_18109,N_16823);
nor UO_1179 (O_1179,N_16451,N_18340);
nor UO_1180 (O_1180,N_19116,N_18999);
xor UO_1181 (O_1181,N_17589,N_19498);
xor UO_1182 (O_1182,N_16716,N_16062);
and UO_1183 (O_1183,N_19045,N_19323);
nor UO_1184 (O_1184,N_17878,N_16328);
or UO_1185 (O_1185,N_19591,N_17329);
xnor UO_1186 (O_1186,N_18720,N_18595);
or UO_1187 (O_1187,N_19055,N_19052);
xnor UO_1188 (O_1188,N_17365,N_18958);
xor UO_1189 (O_1189,N_19209,N_19634);
nor UO_1190 (O_1190,N_17824,N_19019);
and UO_1191 (O_1191,N_18230,N_16381);
xnor UO_1192 (O_1192,N_18597,N_18154);
or UO_1193 (O_1193,N_18079,N_19697);
or UO_1194 (O_1194,N_16492,N_16567);
nor UO_1195 (O_1195,N_19483,N_16524);
nor UO_1196 (O_1196,N_19363,N_19137);
nand UO_1197 (O_1197,N_16256,N_18970);
and UO_1198 (O_1198,N_16247,N_17519);
xor UO_1199 (O_1199,N_16521,N_19640);
and UO_1200 (O_1200,N_16771,N_18987);
or UO_1201 (O_1201,N_17152,N_16508);
nor UO_1202 (O_1202,N_18962,N_16686);
xnor UO_1203 (O_1203,N_19424,N_17886);
and UO_1204 (O_1204,N_19555,N_17347);
or UO_1205 (O_1205,N_17148,N_19558);
xnor UO_1206 (O_1206,N_18268,N_18448);
or UO_1207 (O_1207,N_17835,N_18030);
nand UO_1208 (O_1208,N_17737,N_18184);
or UO_1209 (O_1209,N_19929,N_19277);
or UO_1210 (O_1210,N_17469,N_17323);
or UO_1211 (O_1211,N_16838,N_19769);
nor UO_1212 (O_1212,N_19845,N_16869);
or UO_1213 (O_1213,N_16024,N_16476);
and UO_1214 (O_1214,N_16003,N_18859);
and UO_1215 (O_1215,N_18466,N_17115);
nor UO_1216 (O_1216,N_16543,N_18552);
xor UO_1217 (O_1217,N_18123,N_17358);
or UO_1218 (O_1218,N_16184,N_19034);
nand UO_1219 (O_1219,N_19023,N_17022);
nor UO_1220 (O_1220,N_16700,N_17861);
nand UO_1221 (O_1221,N_17473,N_17671);
nand UO_1222 (O_1222,N_17793,N_16004);
nor UO_1223 (O_1223,N_18214,N_17595);
and UO_1224 (O_1224,N_19900,N_19048);
nor UO_1225 (O_1225,N_17181,N_18378);
nor UO_1226 (O_1226,N_19587,N_18059);
and UO_1227 (O_1227,N_19660,N_17045);
and UO_1228 (O_1228,N_19689,N_19013);
nor UO_1229 (O_1229,N_19294,N_19511);
nand UO_1230 (O_1230,N_17236,N_18846);
nand UO_1231 (O_1231,N_18805,N_19251);
and UO_1232 (O_1232,N_18399,N_17307);
and UO_1233 (O_1233,N_16980,N_18730);
nand UO_1234 (O_1234,N_19579,N_16135);
nor UO_1235 (O_1235,N_16912,N_19071);
nand UO_1236 (O_1236,N_18684,N_19643);
nor UO_1237 (O_1237,N_18180,N_17077);
or UO_1238 (O_1238,N_17247,N_16814);
and UO_1239 (O_1239,N_19139,N_18148);
nor UO_1240 (O_1240,N_19861,N_16544);
and UO_1241 (O_1241,N_18465,N_17556);
and UO_1242 (O_1242,N_18961,N_16896);
and UO_1243 (O_1243,N_16930,N_19448);
and UO_1244 (O_1244,N_19577,N_18789);
nor UO_1245 (O_1245,N_16025,N_19090);
and UO_1246 (O_1246,N_19156,N_16569);
xnor UO_1247 (O_1247,N_17896,N_17321);
nor UO_1248 (O_1248,N_19081,N_16490);
nor UO_1249 (O_1249,N_17050,N_19099);
nand UO_1250 (O_1250,N_16799,N_16423);
xnor UO_1251 (O_1251,N_18092,N_17907);
and UO_1252 (O_1252,N_18433,N_18673);
xor UO_1253 (O_1253,N_16096,N_19986);
or UO_1254 (O_1254,N_16219,N_18099);
and UO_1255 (O_1255,N_17111,N_16289);
or UO_1256 (O_1256,N_19556,N_17637);
nor UO_1257 (O_1257,N_19239,N_18485);
and UO_1258 (O_1258,N_18946,N_18177);
and UO_1259 (O_1259,N_19159,N_17572);
nor UO_1260 (O_1260,N_16616,N_16404);
nand UO_1261 (O_1261,N_18945,N_16861);
or UO_1262 (O_1262,N_16008,N_18201);
nand UO_1263 (O_1263,N_19410,N_16441);
nand UO_1264 (O_1264,N_18168,N_17882);
or UO_1265 (O_1265,N_16570,N_17292);
and UO_1266 (O_1266,N_19153,N_17007);
xor UO_1267 (O_1267,N_18954,N_19309);
nand UO_1268 (O_1268,N_17355,N_18758);
nand UO_1269 (O_1269,N_16665,N_19663);
or UO_1270 (O_1270,N_18026,N_19160);
or UO_1271 (O_1271,N_17012,N_16928);
and UO_1272 (O_1272,N_19520,N_17938);
nor UO_1273 (O_1273,N_18022,N_19817);
nand UO_1274 (O_1274,N_18821,N_17410);
xor UO_1275 (O_1275,N_16205,N_16740);
and UO_1276 (O_1276,N_16582,N_18518);
nand UO_1277 (O_1277,N_18142,N_19883);
and UO_1278 (O_1278,N_17337,N_18747);
xnor UO_1279 (O_1279,N_17094,N_18818);
nand UO_1280 (O_1280,N_17098,N_18172);
nor UO_1281 (O_1281,N_19383,N_18494);
xnor UO_1282 (O_1282,N_16652,N_18839);
and UO_1283 (O_1283,N_17110,N_19739);
nor UO_1284 (O_1284,N_16231,N_18296);
or UO_1285 (O_1285,N_19581,N_18236);
and UO_1286 (O_1286,N_18658,N_18437);
nor UO_1287 (O_1287,N_16737,N_16766);
and UO_1288 (O_1288,N_18197,N_19557);
and UO_1289 (O_1289,N_18540,N_16356);
nand UO_1290 (O_1290,N_18493,N_19830);
nand UO_1291 (O_1291,N_18408,N_18167);
nand UO_1292 (O_1292,N_19155,N_19135);
nor UO_1293 (O_1293,N_16895,N_19496);
nor UO_1294 (O_1294,N_16043,N_16627);
and UO_1295 (O_1295,N_19431,N_19361);
xor UO_1296 (O_1296,N_18000,N_18389);
nor UO_1297 (O_1297,N_16172,N_16383);
and UO_1298 (O_1298,N_18428,N_19458);
or UO_1299 (O_1299,N_19912,N_17129);
and UO_1300 (O_1300,N_16150,N_17585);
nand UO_1301 (O_1301,N_19863,N_16485);
nand UO_1302 (O_1302,N_16807,N_19917);
xnor UO_1303 (O_1303,N_18616,N_16443);
xor UO_1304 (O_1304,N_18560,N_17873);
nor UO_1305 (O_1305,N_16628,N_18474);
nand UO_1306 (O_1306,N_17656,N_16817);
nor UO_1307 (O_1307,N_16970,N_16308);
nor UO_1308 (O_1308,N_17072,N_16197);
and UO_1309 (O_1309,N_16677,N_16364);
and UO_1310 (O_1310,N_16806,N_19955);
xor UO_1311 (O_1311,N_17619,N_18625);
or UO_1312 (O_1312,N_17414,N_19067);
and UO_1313 (O_1313,N_18729,N_18367);
xor UO_1314 (O_1314,N_17987,N_19396);
xor UO_1315 (O_1315,N_16834,N_19971);
and UO_1316 (O_1316,N_17650,N_19357);
xor UO_1317 (O_1317,N_17017,N_18972);
or UO_1318 (O_1318,N_17974,N_18524);
nand UO_1319 (O_1319,N_18522,N_19698);
xnor UO_1320 (O_1320,N_18667,N_17103);
nand UO_1321 (O_1321,N_18916,N_19795);
nand UO_1322 (O_1322,N_18981,N_18107);
nor UO_1323 (O_1323,N_19087,N_18311);
or UO_1324 (O_1324,N_16302,N_17403);
and UO_1325 (O_1325,N_17201,N_17934);
nor UO_1326 (O_1326,N_16233,N_17402);
nor UO_1327 (O_1327,N_17444,N_16747);
nand UO_1328 (O_1328,N_16835,N_18058);
xnor UO_1329 (O_1329,N_17922,N_19467);
xor UO_1330 (O_1330,N_19324,N_19862);
nor UO_1331 (O_1331,N_16045,N_16245);
and UO_1332 (O_1332,N_16969,N_17487);
nand UO_1333 (O_1333,N_19756,N_16360);
xor UO_1334 (O_1334,N_19441,N_17390);
xnor UO_1335 (O_1335,N_18458,N_17068);
nand UO_1336 (O_1336,N_18915,N_16089);
nor UO_1337 (O_1337,N_16523,N_18662);
xnor UO_1338 (O_1338,N_18697,N_18894);
and UO_1339 (O_1339,N_16335,N_16957);
or UO_1340 (O_1340,N_18025,N_16005);
nand UO_1341 (O_1341,N_16985,N_17003);
nor UO_1342 (O_1342,N_19181,N_19375);
nand UO_1343 (O_1343,N_18223,N_19060);
nand UO_1344 (O_1344,N_17442,N_19064);
or UO_1345 (O_1345,N_16201,N_17996);
or UO_1346 (O_1346,N_18823,N_17304);
and UO_1347 (O_1347,N_18565,N_17301);
nand UO_1348 (O_1348,N_18793,N_19730);
nor UO_1349 (O_1349,N_17915,N_19129);
and UO_1350 (O_1350,N_18294,N_19993);
and UO_1351 (O_1351,N_18689,N_17545);
nand UO_1352 (O_1352,N_17067,N_16286);
nand UO_1353 (O_1353,N_17006,N_17674);
and UO_1354 (O_1354,N_17158,N_17547);
and UO_1355 (O_1355,N_19963,N_16622);
and UO_1356 (O_1356,N_17318,N_19380);
or UO_1357 (O_1357,N_17791,N_16939);
nor UO_1358 (O_1358,N_18355,N_16258);
or UO_1359 (O_1359,N_17477,N_16557);
nand UO_1360 (O_1360,N_16727,N_19336);
nand UO_1361 (O_1361,N_17704,N_17021);
or UO_1362 (O_1362,N_18738,N_17751);
xor UO_1363 (O_1363,N_19495,N_16613);
and UO_1364 (O_1364,N_16087,N_17460);
and UO_1365 (O_1365,N_17950,N_17108);
and UO_1366 (O_1366,N_18145,N_18481);
nand UO_1367 (O_1367,N_19601,N_16750);
nor UO_1368 (O_1368,N_19944,N_16914);
nand UO_1369 (O_1369,N_16334,N_18650);
or UO_1370 (O_1370,N_16292,N_19177);
xnor UO_1371 (O_1371,N_16563,N_18052);
nand UO_1372 (O_1372,N_16207,N_19300);
nor UO_1373 (O_1373,N_18527,N_18791);
xnor UO_1374 (O_1374,N_16453,N_17577);
and UO_1375 (O_1375,N_17968,N_19890);
nand UO_1376 (O_1376,N_19171,N_19684);
or UO_1377 (O_1377,N_17663,N_16943);
xor UO_1378 (O_1378,N_19257,N_17225);
xnor UO_1379 (O_1379,N_18708,N_18267);
xor UO_1380 (O_1380,N_17217,N_18069);
and UO_1381 (O_1381,N_18078,N_19611);
nand UO_1382 (O_1382,N_18749,N_18637);
nor UO_1383 (O_1383,N_18831,N_18456);
xor UO_1384 (O_1384,N_18710,N_19031);
nor UO_1385 (O_1385,N_18315,N_16587);
nand UO_1386 (O_1386,N_19044,N_16697);
xnor UO_1387 (O_1387,N_19952,N_17604);
and UO_1388 (O_1388,N_17485,N_16319);
and UO_1389 (O_1389,N_19063,N_18801);
nor UO_1390 (O_1390,N_18589,N_19930);
nand UO_1391 (O_1391,N_19130,N_19151);
nand UO_1392 (O_1392,N_16809,N_19444);
or UO_1393 (O_1393,N_16701,N_18404);
and UO_1394 (O_1394,N_18613,N_19562);
xnor UO_1395 (O_1395,N_16604,N_17220);
or UO_1396 (O_1396,N_18036,N_18890);
nor UO_1397 (O_1397,N_16416,N_17016);
nor UO_1398 (O_1398,N_17957,N_17525);
nand UO_1399 (O_1399,N_16304,N_17784);
nor UO_1400 (O_1400,N_18585,N_18469);
and UO_1401 (O_1401,N_17226,N_17076);
nor UO_1402 (O_1402,N_17313,N_18824);
and UO_1403 (O_1403,N_17667,N_19763);
or UO_1404 (O_1404,N_16063,N_19584);
nor UO_1405 (O_1405,N_17208,N_16511);
nand UO_1406 (O_1406,N_18924,N_16679);
and UO_1407 (O_1407,N_18422,N_17728);
or UO_1408 (O_1408,N_16981,N_17865);
nand UO_1409 (O_1409,N_18449,N_17083);
xnor UO_1410 (O_1410,N_18784,N_17454);
xor UO_1411 (O_1411,N_19404,N_18220);
or UO_1412 (O_1412,N_17130,N_19411);
or UO_1413 (O_1413,N_16907,N_17492);
xnor UO_1414 (O_1414,N_18386,N_17779);
xor UO_1415 (O_1415,N_18554,N_19594);
xor UO_1416 (O_1416,N_18275,N_16298);
nand UO_1417 (O_1417,N_18093,N_18300);
and UO_1418 (O_1418,N_17970,N_16026);
or UO_1419 (O_1419,N_17393,N_19621);
or UO_1420 (O_1420,N_19892,N_19947);
nor UO_1421 (O_1421,N_17215,N_19959);
nand UO_1422 (O_1422,N_17009,N_17743);
xnor UO_1423 (O_1423,N_19620,N_17029);
nand UO_1424 (O_1424,N_16972,N_19296);
nand UO_1425 (O_1425,N_18687,N_16343);
xnor UO_1426 (O_1426,N_18265,N_19369);
and UO_1427 (O_1427,N_17911,N_18063);
nand UO_1428 (O_1428,N_18048,N_18672);
xnor UO_1429 (O_1429,N_18863,N_19445);
or UO_1430 (O_1430,N_16249,N_16352);
xor UO_1431 (O_1431,N_19447,N_16812);
xnor UO_1432 (O_1432,N_17930,N_18407);
nand UO_1433 (O_1433,N_16905,N_16792);
nor UO_1434 (O_1434,N_18029,N_19980);
nand UO_1435 (O_1435,N_17843,N_17584);
nand UO_1436 (O_1436,N_18644,N_17918);
xnor UO_1437 (O_1437,N_17272,N_16660);
nor UO_1438 (O_1438,N_17439,N_17256);
xnor UO_1439 (O_1439,N_19637,N_17170);
nor UO_1440 (O_1440,N_18280,N_16365);
and UO_1441 (O_1441,N_19668,N_18393);
nor UO_1442 (O_1442,N_19077,N_16032);
xnor UO_1443 (O_1443,N_18068,N_16066);
xnor UO_1444 (O_1444,N_18765,N_16744);
nand UO_1445 (O_1445,N_19839,N_19058);
and UO_1446 (O_1446,N_18997,N_17285);
and UO_1447 (O_1447,N_18153,N_18089);
or UO_1448 (O_1448,N_18586,N_17944);
xnor UO_1449 (O_1449,N_18450,N_17276);
nor UO_1450 (O_1450,N_19911,N_18649);
xnor UO_1451 (O_1451,N_18904,N_17677);
nand UO_1452 (O_1452,N_16054,N_17288);
nand UO_1453 (O_1453,N_19473,N_19932);
nand UO_1454 (O_1454,N_16757,N_17407);
and UO_1455 (O_1455,N_16966,N_17140);
and UO_1456 (O_1456,N_18506,N_16495);
nand UO_1457 (O_1457,N_19088,N_18126);
or UO_1458 (O_1458,N_18189,N_19310);
nand UO_1459 (O_1459,N_18426,N_17096);
nand UO_1460 (O_1460,N_19388,N_16578);
nand UO_1461 (O_1461,N_18183,N_18335);
xnor UO_1462 (O_1462,N_17496,N_19614);
nand UO_1463 (O_1463,N_19966,N_17826);
or UO_1464 (O_1464,N_18317,N_18097);
and UO_1465 (O_1465,N_16377,N_16229);
nand UO_1466 (O_1466,N_18996,N_18316);
nor UO_1467 (O_1467,N_19849,N_16802);
or UO_1468 (O_1468,N_19967,N_16499);
or UO_1469 (O_1469,N_17761,N_19539);
nand UO_1470 (O_1470,N_18085,N_18512);
xor UO_1471 (O_1471,N_19694,N_16898);
or UO_1472 (O_1472,N_16502,N_19183);
nor UO_1473 (O_1473,N_18812,N_17435);
nor UO_1474 (O_1474,N_17249,N_17340);
xor UO_1475 (O_1475,N_18243,N_18976);
nor UO_1476 (O_1476,N_18440,N_17681);
xor UO_1477 (O_1477,N_16916,N_16909);
and UO_1478 (O_1478,N_18351,N_16903);
xor UO_1479 (O_1479,N_19927,N_17056);
or UO_1480 (O_1480,N_18828,N_17231);
nor UO_1481 (O_1481,N_17139,N_19973);
xor UO_1482 (O_1482,N_17727,N_18578);
nor UO_1483 (O_1483,N_19161,N_17625);
nor UO_1484 (O_1484,N_16647,N_17801);
or UO_1485 (O_1485,N_18582,N_16240);
nand UO_1486 (O_1486,N_18179,N_17267);
or UO_1487 (O_1487,N_19771,N_17552);
and UO_1488 (O_1488,N_16671,N_18014);
xnor UO_1489 (O_1489,N_18990,N_18967);
xnor UO_1490 (O_1490,N_17709,N_16715);
and UO_1491 (O_1491,N_18752,N_18128);
xor UO_1492 (O_1492,N_19535,N_16948);
nand UO_1493 (O_1493,N_18728,N_19371);
xnor UO_1494 (O_1494,N_18297,N_19523);
or UO_1495 (O_1495,N_17840,N_19354);
xor UO_1496 (O_1496,N_16631,N_17615);
nor UO_1497 (O_1497,N_17010,N_18482);
and UO_1498 (O_1498,N_19825,N_19284);
nor UO_1499 (O_1499,N_16902,N_17431);
or UO_1500 (O_1500,N_19507,N_19847);
or UO_1501 (O_1501,N_19086,N_16685);
xor UO_1502 (O_1502,N_17995,N_18858);
xnor UO_1503 (O_1503,N_18826,N_19118);
and UO_1504 (O_1504,N_16709,N_19488);
or UO_1505 (O_1505,N_19210,N_19570);
nand UO_1506 (O_1506,N_16480,N_17369);
nor UO_1507 (O_1507,N_16790,N_17980);
nor UO_1508 (O_1508,N_18995,N_17754);
xor UO_1509 (O_1509,N_19042,N_19772);
or UO_1510 (O_1510,N_18387,N_17471);
xor UO_1511 (O_1511,N_19994,N_17024);
and UO_1512 (O_1512,N_18118,N_18204);
xnor UO_1513 (O_1513,N_18217,N_19783);
xnor UO_1514 (O_1514,N_19472,N_19345);
nor UO_1515 (O_1515,N_18847,N_18581);
or UO_1516 (O_1516,N_19208,N_16958);
or UO_1517 (O_1517,N_18102,N_19680);
nor UO_1518 (O_1518,N_16193,N_19571);
or UO_1519 (O_1519,N_19547,N_16056);
and UO_1520 (O_1520,N_18800,N_16850);
nand UO_1521 (O_1521,N_17418,N_17409);
or UO_1522 (O_1522,N_19275,N_18119);
and UO_1523 (O_1523,N_19970,N_17906);
or UO_1524 (O_1524,N_17362,N_17833);
nand UO_1525 (O_1525,N_18914,N_17927);
nor UO_1526 (O_1526,N_16767,N_17381);
and UO_1527 (O_1527,N_17732,N_19125);
or UO_1528 (O_1528,N_16710,N_18572);
xnor UO_1529 (O_1529,N_18545,N_17851);
or UO_1530 (O_1530,N_16324,N_18372);
or UO_1531 (O_1531,N_16884,N_18879);
nor UO_1532 (O_1532,N_18436,N_16121);
nand UO_1533 (O_1533,N_19872,N_16146);
nand UO_1534 (O_1534,N_19231,N_18921);
or UO_1535 (O_1535,N_17294,N_18100);
or UO_1536 (O_1536,N_18636,N_18461);
xnor UO_1537 (O_1537,N_19485,N_19166);
xor UO_1538 (O_1538,N_18897,N_17855);
nand UO_1539 (O_1539,N_18938,N_18604);
nor UO_1540 (O_1540,N_19855,N_19252);
or UO_1541 (O_1541,N_16040,N_17689);
xor UO_1542 (O_1542,N_16956,N_16842);
and UO_1543 (O_1543,N_18930,N_17286);
and UO_1544 (O_1544,N_16644,N_19395);
nor UO_1545 (O_1545,N_19687,N_16406);
xnor UO_1546 (O_1546,N_17060,N_19168);
and UO_1547 (O_1547,N_16017,N_17955);
and UO_1548 (O_1548,N_19673,N_18324);
xnor UO_1549 (O_1549,N_18497,N_17529);
and UO_1550 (O_1550,N_16380,N_16347);
xor UO_1551 (O_1551,N_16662,N_17722);
nand UO_1552 (O_1552,N_19860,N_16992);
nor UO_1553 (O_1553,N_17654,N_16878);
nor UO_1554 (O_1554,N_18094,N_19893);
nand UO_1555 (O_1555,N_19884,N_19481);
nor UO_1556 (O_1556,N_16421,N_17936);
nand UO_1557 (O_1557,N_18202,N_19185);
xnor UO_1558 (O_1558,N_17291,N_19082);
or UO_1559 (O_1559,N_16996,N_18418);
and UO_1560 (O_1560,N_18726,N_19333);
and UO_1561 (O_1561,N_17040,N_16494);
or UO_1562 (O_1562,N_16129,N_16455);
and UO_1563 (O_1563,N_17912,N_17849);
nor UO_1564 (O_1564,N_18019,N_18516);
nor UO_1565 (O_1565,N_18678,N_18851);
nand UO_1566 (O_1566,N_18091,N_17322);
xnor UO_1567 (O_1567,N_17638,N_17005);
or UO_1568 (O_1568,N_18359,N_18508);
or UO_1569 (O_1569,N_19220,N_17183);
xnor UO_1570 (O_1570,N_16532,N_18878);
xor UO_1571 (O_1571,N_19657,N_18370);
and UO_1572 (O_1572,N_16718,N_18281);
xor UO_1573 (O_1573,N_16967,N_17361);
and UO_1574 (O_1574,N_16422,N_17384);
or UO_1575 (O_1575,N_16483,N_16369);
nand UO_1576 (O_1576,N_19374,N_18948);
xnor UO_1577 (O_1577,N_19826,N_18287);
nor UO_1578 (O_1578,N_19747,N_17838);
and UO_1579 (O_1579,N_19415,N_17177);
nand UO_1580 (O_1580,N_16048,N_17463);
or UO_1581 (O_1581,N_19180,N_16446);
nor UO_1582 (O_1582,N_19711,N_19554);
nand UO_1583 (O_1583,N_16273,N_18698);
nand UO_1584 (O_1584,N_16648,N_17084);
and UO_1585 (O_1585,N_16465,N_17642);
xor UO_1586 (O_1586,N_18423,N_19559);
nand UO_1587 (O_1587,N_19628,N_19807);
or UO_1588 (O_1588,N_17061,N_18429);
or UO_1589 (O_1589,N_18955,N_16520);
xor UO_1590 (O_1590,N_18745,N_17015);
nor UO_1591 (O_1591,N_19602,N_16932);
nor UO_1592 (O_1592,N_17372,N_16594);
nand UO_1593 (O_1593,N_16815,N_16540);
or UO_1594 (O_1594,N_19502,N_19167);
and UO_1595 (O_1595,N_17752,N_19593);
nand UO_1596 (O_1596,N_18273,N_17764);
and UO_1597 (O_1597,N_18772,N_17900);
xor UO_1598 (O_1598,N_18960,N_16345);
xnor UO_1599 (O_1599,N_17497,N_19541);
nor UO_1600 (O_1600,N_19517,N_18443);
and UO_1601 (O_1601,N_18260,N_18966);
or UO_1602 (O_1602,N_16531,N_19778);
xor UO_1603 (O_1603,N_16528,N_17472);
or UO_1604 (O_1604,N_17778,N_19736);
nor UO_1605 (O_1605,N_17188,N_19907);
or UO_1606 (O_1606,N_17453,N_16326);
and UO_1607 (O_1607,N_16826,N_16925);
nor UO_1608 (O_1608,N_16882,N_17639);
xor UO_1609 (O_1609,N_19127,N_16113);
and UO_1610 (O_1610,N_17107,N_17808);
nor UO_1611 (O_1611,N_19943,N_16103);
nor UO_1612 (O_1612,N_18057,N_18322);
nand UO_1613 (O_1613,N_17392,N_19497);
nor UO_1614 (O_1614,N_18228,N_16639);
nand UO_1615 (O_1615,N_19696,N_17209);
nand UO_1616 (O_1616,N_16461,N_19368);
nor UO_1617 (O_1617,N_17803,N_18427);
xnor UO_1618 (O_1618,N_19981,N_19451);
nor UO_1619 (O_1619,N_16311,N_18357);
and UO_1620 (O_1620,N_17885,N_18519);
xnor UO_1621 (O_1621,N_18304,N_19729);
xor UO_1622 (O_1622,N_17141,N_16974);
xnor UO_1623 (O_1623,N_19776,N_18284);
nor UO_1624 (O_1624,N_19471,N_19436);
nand UO_1625 (O_1625,N_19546,N_19043);
nor UO_1626 (O_1626,N_16649,N_17976);
nor UO_1627 (O_1627,N_19615,N_16774);
or UO_1628 (O_1628,N_18103,N_16169);
or UO_1629 (O_1629,N_17863,N_18760);
nor UO_1630 (O_1630,N_19414,N_16379);
nand UO_1631 (O_1631,N_19616,N_18965);
xnor UO_1632 (O_1632,N_17114,N_17234);
nor UO_1633 (O_1633,N_17568,N_16938);
nor UO_1634 (O_1634,N_17591,N_18583);
and UO_1635 (O_1635,N_16763,N_16276);
nand UO_1636 (O_1636,N_17404,N_16482);
or UO_1637 (O_1637,N_19757,N_18627);
and UO_1638 (O_1638,N_17198,N_19124);
xnor UO_1639 (O_1639,N_17187,N_18892);
nor UO_1640 (O_1640,N_16187,N_18112);
xnor UO_1641 (O_1641,N_18694,N_18612);
nand UO_1642 (O_1642,N_16039,N_17965);
or UO_1643 (O_1643,N_17947,N_16588);
nor UO_1644 (O_1644,N_17316,N_18714);
nand UO_1645 (O_1645,N_18383,N_18867);
nor UO_1646 (O_1646,N_17397,N_19743);
nor UO_1647 (O_1647,N_19321,N_17342);
and UO_1648 (O_1648,N_18515,N_19205);
and UO_1649 (O_1649,N_17011,N_18550);
and UO_1650 (O_1650,N_18786,N_17000);
xor UO_1651 (O_1651,N_18979,N_16659);
nor UO_1652 (O_1652,N_18656,N_17575);
or UO_1653 (O_1653,N_19442,N_19143);
nand UO_1654 (O_1654,N_19066,N_18517);
nand UO_1655 (O_1655,N_19283,N_17768);
nor UO_1656 (O_1656,N_17330,N_16047);
or UO_1657 (O_1657,N_19703,N_16301);
xor UO_1658 (O_1658,N_18732,N_19095);
and UO_1659 (O_1659,N_18751,N_16493);
or UO_1660 (O_1660,N_16646,N_19583);
or UO_1661 (O_1661,N_16949,N_19318);
xor UO_1662 (O_1662,N_16478,N_18696);
and UO_1663 (O_1663,N_16069,N_17926);
xor UO_1664 (O_1664,N_16561,N_17629);
nor UO_1665 (O_1665,N_19024,N_17275);
nand UO_1666 (O_1666,N_19200,N_17428);
or UO_1667 (O_1667,N_17104,N_16420);
and UO_1668 (O_1668,N_17054,N_18657);
and UO_1669 (O_1669,N_16265,N_18390);
or UO_1670 (O_1670,N_18424,N_17753);
and UO_1671 (O_1671,N_18149,N_19290);
or UO_1672 (O_1672,N_16255,N_16760);
nand UO_1673 (O_1673,N_16320,N_18907);
xnor UO_1674 (O_1674,N_19999,N_19779);
and UO_1675 (O_1675,N_17450,N_16235);
nor UO_1676 (O_1676,N_16268,N_19104);
nor UO_1677 (O_1677,N_19102,N_17093);
and UO_1678 (O_1678,N_17020,N_18882);
xnor UO_1679 (O_1679,N_17636,N_17581);
nor UO_1680 (O_1680,N_16598,N_18633);
nor UO_1681 (O_1681,N_17133,N_18271);
nand UO_1682 (O_1682,N_16401,N_18073);
nor UO_1683 (O_1683,N_19551,N_18918);
nor UO_1684 (O_1684,N_17391,N_18181);
or UO_1685 (O_1685,N_19897,N_18971);
xnor UO_1686 (O_1686,N_17872,N_18816);
and UO_1687 (O_1687,N_19229,N_17719);
nor UO_1688 (O_1688,N_17314,N_19376);
and UO_1689 (O_1689,N_19528,N_18573);
and UO_1690 (O_1690,N_16267,N_19827);
nand UO_1691 (O_1691,N_16376,N_18547);
and UO_1692 (O_1692,N_19609,N_19542);
nor UO_1693 (O_1693,N_19937,N_18337);
and UO_1694 (O_1694,N_19107,N_18570);
and UO_1695 (O_1695,N_19891,N_16855);
and UO_1696 (O_1696,N_19233,N_16407);
or UO_1697 (O_1697,N_19512,N_19974);
or UO_1698 (O_1698,N_16614,N_16901);
xnor UO_1699 (O_1699,N_18074,N_18212);
or UO_1700 (O_1700,N_19020,N_17118);
nor UO_1701 (O_1701,N_17597,N_17266);
and UO_1702 (O_1702,N_18680,N_16108);
xor UO_1703 (O_1703,N_16409,N_18491);
xor UO_1704 (O_1704,N_16585,N_17542);
nor UO_1705 (O_1705,N_17343,N_17279);
nor UO_1706 (O_1706,N_18380,N_18592);
xnor UO_1707 (O_1707,N_16526,N_16133);
and UO_1708 (O_1708,N_17387,N_18909);
nor UO_1709 (O_1709,N_16577,N_18391);
or UO_1710 (O_1710,N_17524,N_19639);
and UO_1711 (O_1711,N_18096,N_17502);
nor UO_1712 (O_1712,N_18498,N_16287);
nand UO_1713 (O_1713,N_17583,N_19248);
nand UO_1714 (O_1714,N_17062,N_19259);
and UO_1715 (O_1715,N_18348,N_17367);
xor UO_1716 (O_1716,N_18051,N_16167);
or UO_1717 (O_1717,N_17080,N_19699);
and UO_1718 (O_1718,N_18771,N_19749);
xor UO_1719 (O_1719,N_18632,N_17490);
nand UO_1720 (O_1720,N_16620,N_18639);
nand UO_1721 (O_1721,N_19509,N_16873);
xnor UO_1722 (O_1722,N_19131,N_16322);
nor UO_1723 (O_1723,N_19976,N_18788);
xor UO_1724 (O_1724,N_19805,N_17438);
and UO_1725 (O_1725,N_16927,N_17626);
xnor UO_1726 (O_1726,N_19625,N_18723);
xor UO_1727 (O_1727,N_17713,N_19147);
xor UO_1728 (O_1728,N_16071,N_17700);
nand UO_1729 (O_1729,N_19681,N_17596);
nand UO_1730 (O_1730,N_19122,N_19840);
or UO_1731 (O_1731,N_16192,N_17464);
nor UO_1732 (O_1732,N_17495,N_19780);
and UO_1733 (O_1733,N_16225,N_19298);
xnor UO_1734 (O_1734,N_17905,N_18412);
nor UO_1735 (O_1735,N_19038,N_19016);
and UO_1736 (O_1736,N_19954,N_18208);
xnor UO_1737 (O_1737,N_17510,N_18601);
and UO_1738 (O_1738,N_17829,N_16474);
nor UO_1739 (O_1739,N_17168,N_19553);
nand UO_1740 (O_1740,N_18932,N_19521);
xnor UO_1741 (O_1741,N_17436,N_18648);
nand UO_1742 (O_1742,N_18827,N_18105);
nor UO_1743 (O_1743,N_18401,N_18911);
nor UO_1744 (O_1744,N_18833,N_19702);
nand UO_1745 (O_1745,N_16773,N_16155);
nor UO_1746 (O_1746,N_16093,N_19191);
nor UO_1747 (O_1747,N_16012,N_17964);
xnor UO_1748 (O_1748,N_19716,N_17913);
xor UO_1749 (O_1749,N_19461,N_19325);
xor UO_1750 (O_1750,N_17819,N_18661);
xor UO_1751 (O_1751,N_19062,N_16711);
or UO_1752 (O_1752,N_16159,N_19858);
and UO_1753 (O_1753,N_16653,N_17214);
nand UO_1754 (O_1754,N_19714,N_18403);
or UO_1755 (O_1755,N_17725,N_16836);
and UO_1756 (O_1756,N_16384,N_19683);
nand UO_1757 (O_1757,N_18939,N_16580);
nand UO_1758 (O_1758,N_18488,N_19506);
or UO_1759 (O_1759,N_17925,N_16605);
or UO_1760 (O_1760,N_16507,N_19654);
or UO_1761 (O_1761,N_16266,N_18462);
or UO_1762 (O_1762,N_19501,N_19245);
xor UO_1763 (O_1763,N_16571,N_18953);
or UO_1764 (O_1764,N_19299,N_19314);
or UO_1765 (O_1765,N_17466,N_16393);
and UO_1766 (O_1766,N_17559,N_18855);
nand UO_1767 (O_1767,N_18434,N_18195);
and UO_1768 (O_1768,N_16509,N_16232);
or UO_1769 (O_1769,N_18133,N_19635);
or UO_1770 (O_1770,N_18787,N_16844);
nand UO_1771 (O_1771,N_18464,N_16086);
nor UO_1772 (O_1772,N_18453,N_18883);
and UO_1773 (O_1773,N_19484,N_16527);
nor UO_1774 (O_1774,N_19908,N_17805);
nor UO_1775 (O_1775,N_18902,N_16555);
and UO_1776 (O_1776,N_17551,N_18015);
or UO_1777 (O_1777,N_18147,N_19362);
nand UO_1778 (O_1778,N_19902,N_19710);
and UO_1779 (O_1779,N_16447,N_19126);
nor UO_1780 (O_1780,N_16068,N_16059);
nor UO_1781 (O_1781,N_18379,N_17505);
or UO_1782 (O_1782,N_17406,N_17536);
and UO_1783 (O_1783,N_16019,N_17131);
xnor UO_1784 (O_1784,N_18836,N_17747);
nor UO_1785 (O_1785,N_19649,N_17255);
xnor UO_1786 (O_1786,N_17640,N_19909);
or UO_1787 (O_1787,N_16876,N_17375);
nor UO_1788 (O_1788,N_18320,N_17723);
nand UO_1789 (O_1789,N_17101,N_18158);
nand UO_1790 (O_1790,N_19405,N_18405);
xnor UO_1791 (O_1791,N_18711,N_19070);
or UO_1792 (O_1792,N_17845,N_18870);
nand UO_1793 (O_1793,N_17772,N_16548);
and UO_1794 (O_1794,N_18969,N_19098);
nor UO_1795 (O_1795,N_18130,N_16164);
nand UO_1796 (O_1796,N_16330,N_19968);
and UO_1797 (O_1797,N_18292,N_18568);
or UO_1798 (O_1798,N_16537,N_19638);
nand UO_1799 (O_1799,N_19241,N_18685);
nor UO_1800 (O_1800,N_18477,N_19134);
and UO_1801 (O_1801,N_19935,N_17836);
and UO_1802 (O_1802,N_18557,N_16783);
nand UO_1803 (O_1803,N_16672,N_17890);
and UO_1804 (O_1804,N_16165,N_16151);
and UO_1805 (O_1805,N_16378,N_19773);
nor UO_1806 (O_1806,N_16109,N_17647);
and UO_1807 (O_1807,N_17666,N_16136);
nand UO_1808 (O_1808,N_19788,N_19173);
nor UO_1809 (O_1809,N_19659,N_17981);
xnor UO_1810 (O_1810,N_19574,N_16703);
nor UO_1811 (O_1811,N_17223,N_16119);
nand UO_1812 (O_1812,N_17399,N_17263);
or UO_1813 (O_1813,N_17521,N_19482);
xnor UO_1814 (O_1814,N_18521,N_19995);
and UO_1815 (O_1815,N_19399,N_19381);
nor UO_1816 (O_1816,N_17218,N_17740);
or UO_1817 (O_1817,N_18319,N_18607);
xnor UO_1818 (O_1818,N_19734,N_19450);
nor UO_1819 (O_1819,N_18475,N_19758);
and UO_1820 (O_1820,N_16885,N_17132);
xnor UO_1821 (O_1821,N_17326,N_17440);
or UO_1822 (O_1822,N_16216,N_18301);
or UO_1823 (O_1823,N_18736,N_16112);
and UO_1824 (O_1824,N_18631,N_16020);
nor UO_1825 (O_1825,N_16574,N_19904);
nand UO_1826 (O_1826,N_17465,N_19671);
nor UO_1827 (O_1827,N_19809,N_18900);
or UO_1828 (O_1828,N_16547,N_18065);
nand UO_1829 (O_1829,N_18032,N_16691);
xor UO_1830 (O_1830,N_16116,N_19789);
xnor UO_1831 (O_1831,N_18762,N_18080);
and UO_1832 (O_1832,N_17200,N_19084);
nand UO_1833 (O_1833,N_18835,N_18295);
xor UO_1834 (O_1834,N_18439,N_17310);
nor UO_1835 (O_1835,N_16990,N_18011);
nand UO_1836 (O_1836,N_16307,N_16623);
and UO_1837 (O_1837,N_19263,N_17308);
and UO_1838 (O_1838,N_19675,N_19188);
nand UO_1839 (O_1839,N_18277,N_16236);
nor UO_1840 (O_1840,N_17299,N_18410);
or UO_1841 (O_1841,N_17538,N_17785);
xnor UO_1842 (O_1842,N_18857,N_19326);
or UO_1843 (O_1843,N_18509,N_16678);
nor UO_1844 (O_1844,N_19398,N_17038);
nand UO_1845 (O_1845,N_18249,N_19470);
nor UO_1846 (O_1846,N_17933,N_16280);
nand UO_1847 (O_1847,N_16099,N_16241);
nand UO_1848 (O_1848,N_18356,N_16900);
and UO_1849 (O_1849,N_18899,N_19650);
nor UO_1850 (O_1850,N_17962,N_16624);
and UO_1851 (O_1851,N_18790,N_18756);
nor UO_1852 (O_1852,N_16023,N_18362);
nand UO_1853 (O_1853,N_16410,N_16244);
and UO_1854 (O_1854,N_17766,N_17121);
or UO_1855 (O_1855,N_17189,N_18500);
and UO_1856 (O_1856,N_17960,N_17607);
nor UO_1857 (O_1857,N_16098,N_19978);
and UO_1858 (O_1858,N_17378,N_18323);
or UO_1859 (O_1859,N_17635,N_19746);
nand UO_1860 (O_1860,N_17398,N_16283);
nand UO_1861 (O_1861,N_19764,N_18959);
and UO_1862 (O_1862,N_16489,N_17741);
or UO_1863 (O_1863,N_18898,N_17488);
nand UO_1864 (O_1864,N_16414,N_19053);
or UO_1865 (O_1865,N_19026,N_19110);
nand UO_1866 (O_1866,N_19532,N_16599);
nor UO_1867 (O_1867,N_16999,N_17969);
xnor UO_1868 (O_1868,N_19113,N_18169);
nor UO_1869 (O_1869,N_16357,N_18343);
or UO_1870 (O_1870,N_18364,N_16070);
nand UO_1871 (O_1871,N_17941,N_18013);
nor UO_1872 (O_1872,N_17498,N_17173);
or UO_1873 (O_1873,N_18411,N_16762);
nor UO_1874 (O_1874,N_16091,N_17593);
xnor UO_1875 (O_1875,N_19598,N_16640);
xnor UO_1876 (O_1876,N_18084,N_19744);
nor UO_1877 (O_1877,N_18056,N_16428);
xnor UO_1878 (O_1878,N_19279,N_18888);
or UO_1879 (O_1879,N_19421,N_19015);
nor UO_1880 (O_1880,N_19132,N_16449);
or UO_1881 (O_1881,N_17916,N_19919);
and UO_1882 (O_1882,N_17963,N_19803);
or UO_1883 (O_1883,N_16314,N_17411);
nand UO_1884 (O_1884,N_17986,N_19524);
nand UO_1885 (O_1885,N_16758,N_17004);
nor UO_1886 (O_1886,N_17400,N_17802);
nor UO_1887 (O_1887,N_19940,N_18108);
xor UO_1888 (O_1888,N_17691,N_16095);
xnor UO_1889 (O_1889,N_19631,N_19403);
and UO_1890 (O_1890,N_16803,N_17306);
nand UO_1891 (O_1891,N_19627,N_18182);
nor UO_1892 (O_1892,N_18047,N_17253);
or UO_1893 (O_1893,N_19215,N_18134);
nand UO_1894 (O_1894,N_19091,N_19096);
and UO_1895 (O_1895,N_16881,N_19536);
or UO_1896 (O_1896,N_16712,N_16857);
xor UO_1897 (O_1897,N_18455,N_19247);
nand UO_1898 (O_1898,N_16117,N_19225);
and UO_1899 (O_1899,N_19158,N_19676);
and UO_1900 (O_1900,N_17028,N_19953);
nand UO_1901 (O_1901,N_16795,N_17180);
or UO_1902 (O_1902,N_19560,N_16617);
nand UO_1903 (O_1903,N_17895,N_16339);
and UO_1904 (O_1904,N_17312,N_16663);
and UO_1905 (O_1905,N_17578,N_16670);
or UO_1906 (O_1906,N_19617,N_17690);
xnor UO_1907 (O_1907,N_17516,N_16522);
nor UO_1908 (O_1908,N_18849,N_17769);
and UO_1909 (O_1909,N_19387,N_19494);
nor UO_1910 (O_1910,N_18881,N_17002);
or UO_1911 (O_1911,N_18374,N_19417);
nor UO_1912 (O_1912,N_17661,N_16444);
nand UO_1913 (O_1913,N_17978,N_16995);
or UO_1914 (O_1914,N_17520,N_18232);
and UO_1915 (O_1915,N_17349,N_19735);
or UO_1916 (O_1916,N_19186,N_19811);
and UO_1917 (O_1917,N_19816,N_18803);
and UO_1918 (O_1918,N_19785,N_16813);
nand UO_1919 (O_1919,N_18691,N_17848);
nand UO_1920 (O_1920,N_16488,N_19108);
or UO_1921 (O_1921,N_16296,N_18526);
or UO_1922 (O_1922,N_18151,N_16542);
or UO_1923 (O_1923,N_18361,N_18621);
nor UO_1924 (O_1924,N_19021,N_16568);
nor UO_1925 (O_1925,N_16321,N_16664);
xor UO_1926 (O_1926,N_19831,N_18131);
or UO_1927 (O_1927,N_18432,N_16768);
and UO_1928 (O_1928,N_19392,N_17268);
xor UO_1929 (O_1929,N_17518,N_16057);
nand UO_1930 (O_1930,N_18709,N_19221);
or UO_1931 (O_1931,N_18717,N_18216);
or UO_1932 (O_1932,N_17357,N_19950);
xnor UO_1933 (O_1933,N_17948,N_16163);
xor UO_1934 (O_1934,N_17241,N_19842);
nand UO_1935 (O_1935,N_19149,N_18258);
nand UO_1936 (O_1936,N_19784,N_16088);
and UO_1937 (O_1937,N_18318,N_19001);
and UO_1938 (O_1938,N_17862,N_17457);
and UO_1939 (O_1939,N_19386,N_16964);
or UO_1940 (O_1940,N_19280,N_18298);
xor UO_1941 (O_1941,N_17293,N_18483);
and UO_1942 (O_1942,N_16486,N_19468);
xnor UO_1943 (O_1943,N_18413,N_18564);
xor UO_1944 (O_1944,N_16041,N_19111);
and UO_1945 (O_1945,N_18750,N_19235);
nor UO_1946 (O_1946,N_19400,N_17405);
xnor UO_1947 (O_1947,N_18309,N_18600);
and UO_1948 (O_1948,N_16504,N_16868);
and UO_1949 (O_1949,N_16487,N_16584);
xor UO_1950 (O_1950,N_19316,N_16801);
and UO_1951 (O_1951,N_17333,N_17066);
nand UO_1952 (O_1952,N_17507,N_16316);
xnor UO_1953 (O_1953,N_19335,N_17063);
nand UO_1954 (O_1954,N_16926,N_19446);
and UO_1955 (O_1955,N_18766,N_16942);
nand UO_1956 (O_1956,N_17794,N_17884);
and UO_1957 (O_1957,N_17928,N_18670);
and UO_1958 (O_1958,N_19304,N_18798);
xnor UO_1959 (O_1959,N_19881,N_18302);
nand UO_1960 (O_1960,N_16891,N_16638);
or UO_1961 (O_1961,N_18376,N_18269);
xnor UO_1962 (O_1962,N_17065,N_17587);
nor UO_1963 (O_1963,N_17809,N_18792);
xnor UO_1964 (O_1964,N_17235,N_17999);
nor UO_1965 (O_1965,N_18155,N_17921);
nor UO_1966 (O_1966,N_18435,N_17561);
nor UO_1967 (O_1967,N_16798,N_19549);
or UO_1968 (O_1968,N_18983,N_19267);
and UO_1969 (O_1969,N_17579,N_18611);
xor UO_1970 (O_1970,N_19760,N_18170);
nand UO_1971 (O_1971,N_18555,N_17685);
and UO_1972 (O_1972,N_19223,N_17324);
xor UO_1973 (O_1973,N_17678,N_18173);
or UO_1974 (O_1974,N_18441,N_16463);
or UO_1975 (O_1975,N_17169,N_16018);
nand UO_1976 (O_1976,N_18165,N_16394);
nor UO_1977 (O_1977,N_18206,N_16650);
nand UO_1978 (O_1978,N_16692,N_19164);
nand UO_1979 (O_1979,N_18007,N_17382);
xnor UO_1980 (O_1980,N_17037,N_19390);
nand UO_1981 (O_1981,N_17057,N_18850);
and UO_1982 (O_1982,N_17273,N_17891);
nand UO_1983 (O_1983,N_17874,N_17645);
or UO_1984 (O_1984,N_17048,N_19429);
xnor UO_1985 (O_1985,N_19420,N_19297);
xor UO_1986 (O_1986,N_17734,N_17894);
nor UO_1987 (O_1987,N_16226,N_18088);
nor UO_1988 (O_1988,N_19766,N_18152);
nor UO_1989 (O_1989,N_18700,N_16272);
or UO_1990 (O_1990,N_19848,N_18956);
or UO_1991 (O_1991,N_16124,N_19061);
nor UO_1992 (O_1992,N_17227,N_17229);
xnor UO_1993 (O_1993,N_16516,N_19452);
and UO_1994 (O_1994,N_19589,N_18244);
or UO_1995 (O_1995,N_16689,N_16075);
xnor UO_1996 (O_1996,N_16450,N_16687);
and UO_1997 (O_1997,N_18807,N_16986);
xnor UO_1998 (O_1998,N_17757,N_18018);
or UO_1999 (O_1999,N_19423,N_18513);
and UO_2000 (O_2000,N_18470,N_18188);
xor UO_2001 (O_2001,N_17077,N_19093);
xor UO_2002 (O_2002,N_17495,N_19347);
nor UO_2003 (O_2003,N_18270,N_16842);
xor UO_2004 (O_2004,N_16485,N_16283);
xnor UO_2005 (O_2005,N_16276,N_17777);
nand UO_2006 (O_2006,N_19167,N_18571);
xor UO_2007 (O_2007,N_17206,N_18509);
and UO_2008 (O_2008,N_18547,N_18869);
nor UO_2009 (O_2009,N_18930,N_17461);
xnor UO_2010 (O_2010,N_16064,N_16627);
and UO_2011 (O_2011,N_18428,N_18861);
nand UO_2012 (O_2012,N_18608,N_16107);
and UO_2013 (O_2013,N_16298,N_18715);
and UO_2014 (O_2014,N_19432,N_17321);
and UO_2015 (O_2015,N_18365,N_16464);
or UO_2016 (O_2016,N_16863,N_17734);
or UO_2017 (O_2017,N_18922,N_17385);
nor UO_2018 (O_2018,N_16201,N_17483);
nand UO_2019 (O_2019,N_19295,N_17110);
or UO_2020 (O_2020,N_16947,N_19778);
xnor UO_2021 (O_2021,N_17183,N_17572);
nor UO_2022 (O_2022,N_16670,N_16242);
and UO_2023 (O_2023,N_19494,N_19845);
xnor UO_2024 (O_2024,N_17781,N_18948);
nor UO_2025 (O_2025,N_19698,N_16521);
or UO_2026 (O_2026,N_19459,N_16908);
and UO_2027 (O_2027,N_18969,N_16324);
nand UO_2028 (O_2028,N_18958,N_18578);
or UO_2029 (O_2029,N_16842,N_17906);
nor UO_2030 (O_2030,N_18491,N_19375);
nor UO_2031 (O_2031,N_19908,N_18543);
nor UO_2032 (O_2032,N_17472,N_16581);
or UO_2033 (O_2033,N_19389,N_17538);
and UO_2034 (O_2034,N_19125,N_18761);
and UO_2035 (O_2035,N_18931,N_18735);
nor UO_2036 (O_2036,N_16154,N_16170);
xor UO_2037 (O_2037,N_19651,N_19804);
or UO_2038 (O_2038,N_19371,N_18025);
and UO_2039 (O_2039,N_16853,N_18639);
and UO_2040 (O_2040,N_17391,N_16668);
nor UO_2041 (O_2041,N_18557,N_16605);
nor UO_2042 (O_2042,N_17706,N_17904);
xor UO_2043 (O_2043,N_19141,N_18535);
or UO_2044 (O_2044,N_17277,N_18008);
and UO_2045 (O_2045,N_16608,N_17712);
nand UO_2046 (O_2046,N_16993,N_17620);
nand UO_2047 (O_2047,N_18482,N_18458);
xor UO_2048 (O_2048,N_17218,N_18162);
and UO_2049 (O_2049,N_17260,N_16522);
xnor UO_2050 (O_2050,N_16606,N_17192);
nor UO_2051 (O_2051,N_16306,N_19232);
or UO_2052 (O_2052,N_16664,N_19767);
xnor UO_2053 (O_2053,N_17541,N_19429);
xnor UO_2054 (O_2054,N_16880,N_19656);
and UO_2055 (O_2055,N_16369,N_16650);
xor UO_2056 (O_2056,N_19577,N_18518);
xor UO_2057 (O_2057,N_17604,N_17196);
and UO_2058 (O_2058,N_16059,N_16341);
and UO_2059 (O_2059,N_16370,N_17280);
nor UO_2060 (O_2060,N_16218,N_17510);
nor UO_2061 (O_2061,N_19547,N_17669);
xnor UO_2062 (O_2062,N_19070,N_19361);
or UO_2063 (O_2063,N_18160,N_18755);
xnor UO_2064 (O_2064,N_17521,N_17161);
nor UO_2065 (O_2065,N_17254,N_17883);
xor UO_2066 (O_2066,N_16740,N_17543);
nand UO_2067 (O_2067,N_19226,N_18738);
nor UO_2068 (O_2068,N_18902,N_17973);
and UO_2069 (O_2069,N_18036,N_19032);
or UO_2070 (O_2070,N_19324,N_18255);
or UO_2071 (O_2071,N_17181,N_18596);
or UO_2072 (O_2072,N_19546,N_18009);
xor UO_2073 (O_2073,N_19556,N_19488);
nor UO_2074 (O_2074,N_17144,N_19598);
or UO_2075 (O_2075,N_16455,N_19422);
nand UO_2076 (O_2076,N_16303,N_17689);
nor UO_2077 (O_2077,N_19193,N_19287);
and UO_2078 (O_2078,N_19980,N_19455);
nor UO_2079 (O_2079,N_17916,N_16692);
or UO_2080 (O_2080,N_18752,N_18946);
nor UO_2081 (O_2081,N_19260,N_17982);
nand UO_2082 (O_2082,N_19498,N_16270);
and UO_2083 (O_2083,N_16590,N_18364);
and UO_2084 (O_2084,N_19603,N_18753);
nand UO_2085 (O_2085,N_16161,N_17657);
nand UO_2086 (O_2086,N_19352,N_19685);
xnor UO_2087 (O_2087,N_17779,N_19233);
nor UO_2088 (O_2088,N_18573,N_19209);
xor UO_2089 (O_2089,N_19987,N_18530);
nand UO_2090 (O_2090,N_17024,N_19851);
xnor UO_2091 (O_2091,N_17360,N_17690);
xor UO_2092 (O_2092,N_17608,N_18191);
nand UO_2093 (O_2093,N_18621,N_19846);
xnor UO_2094 (O_2094,N_19584,N_19537);
nand UO_2095 (O_2095,N_19045,N_18739);
or UO_2096 (O_2096,N_16737,N_16579);
or UO_2097 (O_2097,N_18140,N_17146);
or UO_2098 (O_2098,N_19958,N_16343);
nor UO_2099 (O_2099,N_18137,N_18618);
and UO_2100 (O_2100,N_17503,N_19523);
nand UO_2101 (O_2101,N_16508,N_16057);
or UO_2102 (O_2102,N_18050,N_19966);
xor UO_2103 (O_2103,N_18205,N_16672);
or UO_2104 (O_2104,N_18757,N_17971);
nor UO_2105 (O_2105,N_19135,N_17844);
and UO_2106 (O_2106,N_17177,N_17352);
nand UO_2107 (O_2107,N_16343,N_17415);
nor UO_2108 (O_2108,N_16321,N_19681);
or UO_2109 (O_2109,N_17385,N_16191);
nand UO_2110 (O_2110,N_17840,N_16552);
nor UO_2111 (O_2111,N_19381,N_16272);
nand UO_2112 (O_2112,N_18314,N_17672);
and UO_2113 (O_2113,N_16650,N_17456);
nor UO_2114 (O_2114,N_18771,N_18075);
nor UO_2115 (O_2115,N_18762,N_18746);
nor UO_2116 (O_2116,N_16464,N_16036);
xnor UO_2117 (O_2117,N_17800,N_18013);
and UO_2118 (O_2118,N_18157,N_18556);
nor UO_2119 (O_2119,N_18512,N_19482);
or UO_2120 (O_2120,N_19389,N_18975);
nand UO_2121 (O_2121,N_16765,N_19555);
xor UO_2122 (O_2122,N_16307,N_16733);
nor UO_2123 (O_2123,N_16183,N_16931);
xor UO_2124 (O_2124,N_19584,N_16722);
xnor UO_2125 (O_2125,N_19451,N_18025);
or UO_2126 (O_2126,N_18066,N_16520);
nor UO_2127 (O_2127,N_18098,N_19921);
nor UO_2128 (O_2128,N_18474,N_18011);
nor UO_2129 (O_2129,N_16748,N_16827);
and UO_2130 (O_2130,N_19994,N_17697);
xnor UO_2131 (O_2131,N_17139,N_19488);
nor UO_2132 (O_2132,N_18526,N_19844);
nand UO_2133 (O_2133,N_18965,N_16255);
and UO_2134 (O_2134,N_18973,N_18627);
nor UO_2135 (O_2135,N_19288,N_19850);
nor UO_2136 (O_2136,N_18592,N_16767);
nand UO_2137 (O_2137,N_17350,N_18734);
or UO_2138 (O_2138,N_16941,N_17717);
nand UO_2139 (O_2139,N_16903,N_18556);
nor UO_2140 (O_2140,N_18120,N_18873);
or UO_2141 (O_2141,N_16819,N_18830);
and UO_2142 (O_2142,N_17843,N_18319);
nand UO_2143 (O_2143,N_19854,N_19970);
and UO_2144 (O_2144,N_18362,N_18222);
or UO_2145 (O_2145,N_19601,N_17281);
and UO_2146 (O_2146,N_17486,N_18785);
xor UO_2147 (O_2147,N_18887,N_18483);
or UO_2148 (O_2148,N_17143,N_18143);
or UO_2149 (O_2149,N_18948,N_16217);
xor UO_2150 (O_2150,N_19805,N_18247);
nand UO_2151 (O_2151,N_19839,N_18298);
and UO_2152 (O_2152,N_16603,N_18442);
xor UO_2153 (O_2153,N_19587,N_18527);
or UO_2154 (O_2154,N_19690,N_19574);
and UO_2155 (O_2155,N_18511,N_16325);
or UO_2156 (O_2156,N_18559,N_19713);
xor UO_2157 (O_2157,N_18722,N_18970);
and UO_2158 (O_2158,N_17194,N_16842);
xor UO_2159 (O_2159,N_19998,N_17732);
nand UO_2160 (O_2160,N_18385,N_19811);
and UO_2161 (O_2161,N_16628,N_16832);
and UO_2162 (O_2162,N_18797,N_17546);
nand UO_2163 (O_2163,N_17013,N_19965);
and UO_2164 (O_2164,N_19450,N_18246);
nor UO_2165 (O_2165,N_17551,N_19646);
xnor UO_2166 (O_2166,N_19581,N_16634);
and UO_2167 (O_2167,N_16554,N_17117);
and UO_2168 (O_2168,N_19586,N_19559);
xnor UO_2169 (O_2169,N_17925,N_16809);
or UO_2170 (O_2170,N_17604,N_16584);
and UO_2171 (O_2171,N_17539,N_19941);
or UO_2172 (O_2172,N_17888,N_17286);
and UO_2173 (O_2173,N_16935,N_16010);
nor UO_2174 (O_2174,N_19639,N_16719);
and UO_2175 (O_2175,N_18262,N_18130);
nor UO_2176 (O_2176,N_17073,N_19629);
or UO_2177 (O_2177,N_16777,N_18086);
xor UO_2178 (O_2178,N_18507,N_17657);
and UO_2179 (O_2179,N_18010,N_19383);
or UO_2180 (O_2180,N_16242,N_18873);
xor UO_2181 (O_2181,N_17536,N_19983);
nor UO_2182 (O_2182,N_18704,N_16444);
nor UO_2183 (O_2183,N_16787,N_18760);
nand UO_2184 (O_2184,N_17574,N_19205);
and UO_2185 (O_2185,N_19719,N_18698);
xor UO_2186 (O_2186,N_17403,N_16503);
nand UO_2187 (O_2187,N_17158,N_19455);
nor UO_2188 (O_2188,N_18908,N_17344);
nand UO_2189 (O_2189,N_18528,N_17339);
nor UO_2190 (O_2190,N_17713,N_17497);
and UO_2191 (O_2191,N_16429,N_16840);
nor UO_2192 (O_2192,N_18165,N_16587);
nor UO_2193 (O_2193,N_16389,N_19396);
nor UO_2194 (O_2194,N_16740,N_17165);
xor UO_2195 (O_2195,N_18778,N_18722);
and UO_2196 (O_2196,N_17812,N_19831);
nor UO_2197 (O_2197,N_19981,N_17240);
or UO_2198 (O_2198,N_17465,N_19855);
or UO_2199 (O_2199,N_18202,N_18204);
or UO_2200 (O_2200,N_18674,N_17399);
nor UO_2201 (O_2201,N_16620,N_18680);
xor UO_2202 (O_2202,N_17428,N_16730);
nand UO_2203 (O_2203,N_19857,N_18509);
nand UO_2204 (O_2204,N_18181,N_17624);
nor UO_2205 (O_2205,N_19657,N_18993);
and UO_2206 (O_2206,N_16167,N_18367);
nor UO_2207 (O_2207,N_16697,N_18112);
nand UO_2208 (O_2208,N_19912,N_18500);
or UO_2209 (O_2209,N_17498,N_17275);
xor UO_2210 (O_2210,N_18318,N_19804);
or UO_2211 (O_2211,N_19723,N_17798);
nand UO_2212 (O_2212,N_17154,N_16374);
or UO_2213 (O_2213,N_17621,N_19257);
xnor UO_2214 (O_2214,N_17835,N_18512);
xnor UO_2215 (O_2215,N_18747,N_18042);
or UO_2216 (O_2216,N_19862,N_17300);
and UO_2217 (O_2217,N_16977,N_18173);
or UO_2218 (O_2218,N_16779,N_19815);
and UO_2219 (O_2219,N_17232,N_18522);
nand UO_2220 (O_2220,N_18853,N_19507);
and UO_2221 (O_2221,N_16284,N_16810);
or UO_2222 (O_2222,N_19914,N_17402);
nor UO_2223 (O_2223,N_18743,N_19618);
nor UO_2224 (O_2224,N_18450,N_19829);
xor UO_2225 (O_2225,N_16591,N_17737);
nand UO_2226 (O_2226,N_17821,N_19376);
and UO_2227 (O_2227,N_16425,N_18518);
and UO_2228 (O_2228,N_18938,N_17714);
nor UO_2229 (O_2229,N_17277,N_16277);
and UO_2230 (O_2230,N_18034,N_16202);
and UO_2231 (O_2231,N_17907,N_18779);
nand UO_2232 (O_2232,N_19755,N_18331);
nand UO_2233 (O_2233,N_17179,N_19939);
nand UO_2234 (O_2234,N_16116,N_16099);
nand UO_2235 (O_2235,N_18667,N_18390);
and UO_2236 (O_2236,N_19075,N_17609);
xor UO_2237 (O_2237,N_18050,N_17270);
and UO_2238 (O_2238,N_17997,N_19353);
and UO_2239 (O_2239,N_18507,N_19556);
nand UO_2240 (O_2240,N_17068,N_16260);
xor UO_2241 (O_2241,N_16152,N_17284);
nand UO_2242 (O_2242,N_17488,N_18497);
nor UO_2243 (O_2243,N_19994,N_16539);
nand UO_2244 (O_2244,N_17014,N_17424);
nor UO_2245 (O_2245,N_16026,N_19489);
and UO_2246 (O_2246,N_16424,N_16428);
or UO_2247 (O_2247,N_17224,N_17273);
nand UO_2248 (O_2248,N_18876,N_17011);
nor UO_2249 (O_2249,N_18805,N_19984);
nand UO_2250 (O_2250,N_19168,N_17861);
xnor UO_2251 (O_2251,N_17094,N_16007);
or UO_2252 (O_2252,N_18602,N_19001);
or UO_2253 (O_2253,N_17083,N_19095);
xor UO_2254 (O_2254,N_19370,N_17529);
and UO_2255 (O_2255,N_19569,N_16980);
nor UO_2256 (O_2256,N_16097,N_18756);
and UO_2257 (O_2257,N_17997,N_18115);
xor UO_2258 (O_2258,N_18308,N_16795);
xnor UO_2259 (O_2259,N_19999,N_18451);
nand UO_2260 (O_2260,N_18171,N_17726);
and UO_2261 (O_2261,N_18091,N_16855);
nand UO_2262 (O_2262,N_18867,N_18641);
or UO_2263 (O_2263,N_19871,N_19603);
and UO_2264 (O_2264,N_16427,N_18701);
or UO_2265 (O_2265,N_17083,N_16824);
nor UO_2266 (O_2266,N_18874,N_17394);
nor UO_2267 (O_2267,N_17320,N_18037);
and UO_2268 (O_2268,N_16349,N_17215);
nand UO_2269 (O_2269,N_16768,N_19348);
and UO_2270 (O_2270,N_18352,N_17308);
and UO_2271 (O_2271,N_18614,N_16656);
nor UO_2272 (O_2272,N_17146,N_16826);
nand UO_2273 (O_2273,N_18971,N_19076);
nand UO_2274 (O_2274,N_18210,N_18483);
xor UO_2275 (O_2275,N_16610,N_16460);
nand UO_2276 (O_2276,N_17599,N_17417);
xnor UO_2277 (O_2277,N_16841,N_17117);
nand UO_2278 (O_2278,N_16292,N_18337);
nor UO_2279 (O_2279,N_16261,N_19766);
or UO_2280 (O_2280,N_18830,N_18820);
xor UO_2281 (O_2281,N_16053,N_19375);
nand UO_2282 (O_2282,N_17132,N_19863);
and UO_2283 (O_2283,N_19318,N_17357);
nor UO_2284 (O_2284,N_19899,N_17373);
nand UO_2285 (O_2285,N_16641,N_16138);
xnor UO_2286 (O_2286,N_19677,N_19859);
nor UO_2287 (O_2287,N_18780,N_16147);
or UO_2288 (O_2288,N_16185,N_18383);
xnor UO_2289 (O_2289,N_18303,N_19285);
nand UO_2290 (O_2290,N_18515,N_18058);
nand UO_2291 (O_2291,N_18312,N_19460);
and UO_2292 (O_2292,N_16917,N_17507);
and UO_2293 (O_2293,N_17329,N_18062);
or UO_2294 (O_2294,N_16566,N_17682);
xnor UO_2295 (O_2295,N_19327,N_18760);
and UO_2296 (O_2296,N_17343,N_16483);
and UO_2297 (O_2297,N_18031,N_18292);
nand UO_2298 (O_2298,N_16447,N_19641);
and UO_2299 (O_2299,N_18345,N_17666);
xor UO_2300 (O_2300,N_17767,N_19261);
nand UO_2301 (O_2301,N_17862,N_19826);
xor UO_2302 (O_2302,N_19474,N_18958);
nand UO_2303 (O_2303,N_16588,N_18195);
or UO_2304 (O_2304,N_19266,N_18903);
and UO_2305 (O_2305,N_18048,N_17088);
nor UO_2306 (O_2306,N_17086,N_18307);
nor UO_2307 (O_2307,N_16644,N_16041);
nor UO_2308 (O_2308,N_19201,N_17980);
nor UO_2309 (O_2309,N_19251,N_19262);
or UO_2310 (O_2310,N_18862,N_16935);
or UO_2311 (O_2311,N_18857,N_19003);
nor UO_2312 (O_2312,N_18939,N_17732);
or UO_2313 (O_2313,N_16731,N_16399);
nand UO_2314 (O_2314,N_18674,N_16292);
and UO_2315 (O_2315,N_17657,N_19385);
nor UO_2316 (O_2316,N_16928,N_17584);
nand UO_2317 (O_2317,N_19779,N_19839);
nor UO_2318 (O_2318,N_16564,N_19102);
and UO_2319 (O_2319,N_17612,N_16362);
or UO_2320 (O_2320,N_19597,N_16940);
nand UO_2321 (O_2321,N_16824,N_16370);
xor UO_2322 (O_2322,N_16026,N_18144);
and UO_2323 (O_2323,N_19111,N_19483);
xor UO_2324 (O_2324,N_19640,N_16867);
and UO_2325 (O_2325,N_18532,N_19124);
and UO_2326 (O_2326,N_16568,N_19046);
nand UO_2327 (O_2327,N_17374,N_19783);
and UO_2328 (O_2328,N_19206,N_18023);
xnor UO_2329 (O_2329,N_18837,N_17189);
or UO_2330 (O_2330,N_19658,N_16125);
nand UO_2331 (O_2331,N_19066,N_19970);
or UO_2332 (O_2332,N_18094,N_16185);
nand UO_2333 (O_2333,N_19952,N_16741);
and UO_2334 (O_2334,N_17684,N_19084);
nor UO_2335 (O_2335,N_17594,N_17415);
or UO_2336 (O_2336,N_17923,N_19388);
nor UO_2337 (O_2337,N_19260,N_16887);
or UO_2338 (O_2338,N_17752,N_19548);
xor UO_2339 (O_2339,N_18659,N_18986);
or UO_2340 (O_2340,N_16723,N_17285);
xor UO_2341 (O_2341,N_19286,N_19949);
nand UO_2342 (O_2342,N_18548,N_19323);
xor UO_2343 (O_2343,N_18029,N_19622);
and UO_2344 (O_2344,N_19405,N_16511);
nand UO_2345 (O_2345,N_19595,N_19729);
nand UO_2346 (O_2346,N_19551,N_19212);
or UO_2347 (O_2347,N_17574,N_18443);
nor UO_2348 (O_2348,N_17011,N_16280);
and UO_2349 (O_2349,N_16487,N_19211);
or UO_2350 (O_2350,N_17950,N_17516);
xnor UO_2351 (O_2351,N_16233,N_18212);
and UO_2352 (O_2352,N_18799,N_17888);
xnor UO_2353 (O_2353,N_18330,N_16926);
and UO_2354 (O_2354,N_18444,N_19973);
xnor UO_2355 (O_2355,N_18070,N_19668);
xnor UO_2356 (O_2356,N_18000,N_19086);
and UO_2357 (O_2357,N_18085,N_17777);
and UO_2358 (O_2358,N_16421,N_19441);
xor UO_2359 (O_2359,N_19179,N_16341);
and UO_2360 (O_2360,N_16691,N_17995);
xnor UO_2361 (O_2361,N_17280,N_19852);
or UO_2362 (O_2362,N_16973,N_16778);
and UO_2363 (O_2363,N_19519,N_16151);
xnor UO_2364 (O_2364,N_16288,N_19696);
nand UO_2365 (O_2365,N_18411,N_19115);
xnor UO_2366 (O_2366,N_17006,N_19255);
xor UO_2367 (O_2367,N_17189,N_17006);
nor UO_2368 (O_2368,N_19244,N_17810);
nand UO_2369 (O_2369,N_16690,N_18613);
and UO_2370 (O_2370,N_16935,N_16712);
or UO_2371 (O_2371,N_18384,N_17733);
and UO_2372 (O_2372,N_18001,N_16046);
nand UO_2373 (O_2373,N_16487,N_17801);
nor UO_2374 (O_2374,N_18392,N_16542);
nor UO_2375 (O_2375,N_19849,N_16410);
and UO_2376 (O_2376,N_17033,N_16115);
and UO_2377 (O_2377,N_17764,N_17329);
xor UO_2378 (O_2378,N_18574,N_16518);
nor UO_2379 (O_2379,N_19482,N_19899);
xnor UO_2380 (O_2380,N_17112,N_19178);
nand UO_2381 (O_2381,N_17365,N_17945);
and UO_2382 (O_2382,N_19127,N_18124);
or UO_2383 (O_2383,N_16335,N_18704);
nand UO_2384 (O_2384,N_18767,N_17938);
nand UO_2385 (O_2385,N_17852,N_17026);
and UO_2386 (O_2386,N_18035,N_16837);
and UO_2387 (O_2387,N_18258,N_17710);
or UO_2388 (O_2388,N_19257,N_17625);
or UO_2389 (O_2389,N_19617,N_17064);
nor UO_2390 (O_2390,N_18941,N_17824);
nor UO_2391 (O_2391,N_18354,N_18749);
or UO_2392 (O_2392,N_16056,N_16719);
and UO_2393 (O_2393,N_16867,N_18905);
nand UO_2394 (O_2394,N_17221,N_16513);
nor UO_2395 (O_2395,N_19777,N_18176);
nand UO_2396 (O_2396,N_19721,N_16667);
nand UO_2397 (O_2397,N_18869,N_16448);
xor UO_2398 (O_2398,N_18195,N_16343);
nor UO_2399 (O_2399,N_17869,N_17625);
nand UO_2400 (O_2400,N_18573,N_17134);
and UO_2401 (O_2401,N_17223,N_18225);
or UO_2402 (O_2402,N_16036,N_18174);
or UO_2403 (O_2403,N_18921,N_19159);
nor UO_2404 (O_2404,N_19342,N_17694);
xnor UO_2405 (O_2405,N_17444,N_16548);
or UO_2406 (O_2406,N_17993,N_19957);
nor UO_2407 (O_2407,N_16375,N_19505);
nor UO_2408 (O_2408,N_19069,N_19374);
nand UO_2409 (O_2409,N_19495,N_19919);
nor UO_2410 (O_2410,N_17375,N_18793);
or UO_2411 (O_2411,N_19549,N_17348);
or UO_2412 (O_2412,N_19346,N_19984);
nand UO_2413 (O_2413,N_18831,N_17400);
nor UO_2414 (O_2414,N_18959,N_19174);
and UO_2415 (O_2415,N_18279,N_17231);
xor UO_2416 (O_2416,N_18847,N_17226);
nor UO_2417 (O_2417,N_17355,N_17994);
xor UO_2418 (O_2418,N_19193,N_17330);
or UO_2419 (O_2419,N_16756,N_18151);
or UO_2420 (O_2420,N_18631,N_19702);
nand UO_2421 (O_2421,N_19925,N_17859);
or UO_2422 (O_2422,N_16496,N_17357);
nand UO_2423 (O_2423,N_19208,N_19056);
and UO_2424 (O_2424,N_17493,N_18828);
and UO_2425 (O_2425,N_16010,N_19903);
nor UO_2426 (O_2426,N_18163,N_18688);
nand UO_2427 (O_2427,N_18956,N_16137);
and UO_2428 (O_2428,N_16715,N_16078);
nand UO_2429 (O_2429,N_19786,N_16968);
xor UO_2430 (O_2430,N_17713,N_18278);
nor UO_2431 (O_2431,N_16661,N_16865);
xnor UO_2432 (O_2432,N_17558,N_17758);
and UO_2433 (O_2433,N_17634,N_19287);
and UO_2434 (O_2434,N_17040,N_17047);
nor UO_2435 (O_2435,N_19283,N_16911);
nor UO_2436 (O_2436,N_17759,N_17648);
nand UO_2437 (O_2437,N_19440,N_17255);
and UO_2438 (O_2438,N_16322,N_16477);
nand UO_2439 (O_2439,N_18182,N_19728);
nor UO_2440 (O_2440,N_17843,N_19764);
nand UO_2441 (O_2441,N_18615,N_16646);
or UO_2442 (O_2442,N_16065,N_19110);
and UO_2443 (O_2443,N_19163,N_17548);
nand UO_2444 (O_2444,N_16688,N_17118);
xnor UO_2445 (O_2445,N_17439,N_18393);
nor UO_2446 (O_2446,N_19935,N_16564);
and UO_2447 (O_2447,N_16546,N_17311);
nand UO_2448 (O_2448,N_19345,N_16021);
and UO_2449 (O_2449,N_18700,N_18218);
xnor UO_2450 (O_2450,N_19860,N_16062);
nor UO_2451 (O_2451,N_19787,N_17383);
and UO_2452 (O_2452,N_19950,N_19060);
and UO_2453 (O_2453,N_16376,N_18521);
xnor UO_2454 (O_2454,N_19645,N_17702);
and UO_2455 (O_2455,N_17587,N_19136);
or UO_2456 (O_2456,N_17400,N_19224);
nor UO_2457 (O_2457,N_19345,N_17244);
nand UO_2458 (O_2458,N_18593,N_19142);
nor UO_2459 (O_2459,N_16608,N_18290);
and UO_2460 (O_2460,N_18423,N_16102);
nand UO_2461 (O_2461,N_16466,N_16683);
xnor UO_2462 (O_2462,N_16018,N_18766);
or UO_2463 (O_2463,N_17833,N_19315);
or UO_2464 (O_2464,N_17914,N_18653);
nor UO_2465 (O_2465,N_16861,N_17622);
nand UO_2466 (O_2466,N_16412,N_17868);
or UO_2467 (O_2467,N_17263,N_16068);
nand UO_2468 (O_2468,N_18616,N_19915);
xnor UO_2469 (O_2469,N_16237,N_18008);
nand UO_2470 (O_2470,N_17557,N_19240);
or UO_2471 (O_2471,N_19589,N_19925);
and UO_2472 (O_2472,N_17612,N_17221);
xnor UO_2473 (O_2473,N_17732,N_17038);
nor UO_2474 (O_2474,N_18199,N_19407);
nor UO_2475 (O_2475,N_17807,N_19637);
nor UO_2476 (O_2476,N_16788,N_19733);
and UO_2477 (O_2477,N_18379,N_19273);
nand UO_2478 (O_2478,N_16119,N_19743);
and UO_2479 (O_2479,N_16259,N_17522);
xnor UO_2480 (O_2480,N_17069,N_16063);
nand UO_2481 (O_2481,N_16116,N_19241);
and UO_2482 (O_2482,N_17442,N_18671);
nand UO_2483 (O_2483,N_17837,N_16955);
and UO_2484 (O_2484,N_17506,N_16744);
or UO_2485 (O_2485,N_19548,N_17991);
or UO_2486 (O_2486,N_18643,N_19676);
xnor UO_2487 (O_2487,N_19072,N_17996);
xnor UO_2488 (O_2488,N_18898,N_19088);
and UO_2489 (O_2489,N_18975,N_18103);
or UO_2490 (O_2490,N_18491,N_17895);
xor UO_2491 (O_2491,N_17890,N_16273);
nand UO_2492 (O_2492,N_18747,N_17389);
nand UO_2493 (O_2493,N_17519,N_17267);
xor UO_2494 (O_2494,N_19914,N_18682);
or UO_2495 (O_2495,N_19979,N_19685);
and UO_2496 (O_2496,N_18801,N_18755);
nand UO_2497 (O_2497,N_19654,N_18894);
nand UO_2498 (O_2498,N_16178,N_17819);
and UO_2499 (O_2499,N_18688,N_19545);
endmodule